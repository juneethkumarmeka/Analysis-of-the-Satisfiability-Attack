module basic_3000_30000_3500_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_1357,In_620);
or U1 (N_1,In_2512,In_1053);
or U2 (N_2,In_2750,In_2073);
or U3 (N_3,In_1156,In_1421);
and U4 (N_4,In_1925,In_2204);
nor U5 (N_5,In_847,In_744);
nor U6 (N_6,In_2318,In_2738);
and U7 (N_7,In_2333,In_113);
and U8 (N_8,In_80,In_1687);
nor U9 (N_9,In_2595,In_795);
nand U10 (N_10,In_474,In_1581);
nor U11 (N_11,In_2896,In_2614);
nor U12 (N_12,In_96,In_2583);
nand U13 (N_13,In_2920,In_699);
nand U14 (N_14,In_1203,In_1928);
nor U15 (N_15,In_1834,In_2727);
nand U16 (N_16,In_2115,In_46);
and U17 (N_17,In_1532,In_2167);
nor U18 (N_18,In_2586,In_1645);
nor U19 (N_19,In_1153,In_1688);
xor U20 (N_20,In_1122,In_2615);
and U21 (N_21,In_2027,In_2916);
nor U22 (N_22,In_1046,In_641);
xor U23 (N_23,In_2867,In_693);
nor U24 (N_24,In_2224,In_457);
nand U25 (N_25,In_2078,In_2416);
xnor U26 (N_26,In_2732,In_887);
nand U27 (N_27,In_1367,In_966);
or U28 (N_28,In_1021,In_566);
nand U29 (N_29,In_537,In_184);
xnor U30 (N_30,In_2068,In_2638);
nand U31 (N_31,In_298,In_840);
nand U32 (N_32,In_318,In_825);
and U33 (N_33,In_62,In_1103);
nand U34 (N_34,In_741,In_1220);
or U35 (N_35,In_736,In_792);
or U36 (N_36,In_72,In_1691);
or U37 (N_37,In_619,In_2449);
nand U38 (N_38,In_2852,In_1467);
and U39 (N_39,In_544,In_1833);
xor U40 (N_40,In_2571,In_479);
and U41 (N_41,In_900,In_1383);
or U42 (N_42,In_1571,In_1978);
nor U43 (N_43,In_814,In_1698);
or U44 (N_44,In_2917,In_2069);
nor U45 (N_45,In_2108,In_2451);
and U46 (N_46,In_2533,In_1321);
nand U47 (N_47,In_2706,In_1546);
nor U48 (N_48,In_994,In_47);
and U49 (N_49,In_743,In_1128);
or U50 (N_50,In_1562,In_928);
or U51 (N_51,In_2754,In_2504);
xnor U52 (N_52,In_2822,In_2802);
or U53 (N_53,In_2551,In_289);
nor U54 (N_54,In_1629,In_297);
or U55 (N_55,In_2398,In_762);
xnor U56 (N_56,In_2966,In_453);
xor U57 (N_57,In_1118,In_2319);
and U58 (N_58,In_2400,In_2077);
nor U59 (N_59,In_1214,In_1719);
nand U60 (N_60,In_607,In_462);
xnor U61 (N_61,In_2976,In_2579);
nand U62 (N_62,In_456,In_821);
and U63 (N_63,In_2621,In_2532);
xnor U64 (N_64,In_1011,In_508);
and U65 (N_65,In_243,In_1152);
nor U66 (N_66,In_2019,In_2634);
or U67 (N_67,In_2662,In_2567);
nand U68 (N_68,In_734,In_2020);
nor U69 (N_69,In_341,In_2212);
nand U70 (N_70,In_2023,In_2182);
nand U71 (N_71,In_150,In_2796);
xnor U72 (N_72,In_2828,In_2274);
nand U73 (N_73,In_503,In_657);
nor U74 (N_74,In_956,In_1873);
nand U75 (N_75,In_28,In_1393);
xnor U76 (N_76,In_407,In_127);
xnor U77 (N_77,In_514,In_1548);
or U78 (N_78,In_1625,In_93);
and U79 (N_79,In_1588,In_2511);
xor U80 (N_80,In_1398,In_37);
nor U81 (N_81,In_991,In_173);
nor U82 (N_82,In_2798,In_2777);
xor U83 (N_83,In_1486,In_708);
nand U84 (N_84,In_1524,In_1644);
or U85 (N_85,In_1161,In_1353);
xor U86 (N_86,In_147,In_2229);
nor U87 (N_87,In_1423,In_1433);
and U88 (N_88,In_1222,In_2792);
nand U89 (N_89,In_258,In_2658);
nand U90 (N_90,In_2993,In_2900);
xor U91 (N_91,In_1198,In_2873);
or U92 (N_92,In_2158,In_123);
nor U93 (N_93,In_977,In_969);
xnor U94 (N_94,In_981,In_2813);
nand U95 (N_95,In_979,In_601);
nand U96 (N_96,In_141,In_1035);
nor U97 (N_97,In_1692,In_2098);
nor U98 (N_98,In_1980,In_2979);
nand U99 (N_99,In_39,In_749);
nor U100 (N_100,In_1074,In_1133);
nand U101 (N_101,In_2371,In_2779);
nand U102 (N_102,In_2506,In_1595);
or U103 (N_103,In_1759,In_1683);
nand U104 (N_104,In_2804,In_1263);
xor U105 (N_105,In_522,In_975);
or U106 (N_106,In_1494,In_2345);
xnor U107 (N_107,In_1662,In_2861);
or U108 (N_108,In_581,In_1374);
and U109 (N_109,In_1717,In_2847);
nand U110 (N_110,In_2965,In_2324);
nand U111 (N_111,In_65,In_2885);
xor U112 (N_112,In_628,In_1368);
or U113 (N_113,In_1530,In_475);
or U114 (N_114,In_1193,In_2559);
and U115 (N_115,In_2737,In_338);
and U116 (N_116,In_133,In_691);
xor U117 (N_117,In_2929,In_2924);
and U118 (N_118,In_142,In_2962);
nor U119 (N_119,In_550,In_2630);
nor U120 (N_120,In_904,In_1407);
nor U121 (N_121,In_2473,In_2940);
and U122 (N_122,In_2969,In_2017);
nor U123 (N_123,In_1885,In_712);
xnor U124 (N_124,In_73,In_1438);
xor U125 (N_125,In_2958,In_2139);
nor U126 (N_126,In_2679,In_1646);
xnor U127 (N_127,In_198,In_1617);
xor U128 (N_128,In_2650,In_871);
and U129 (N_129,In_1556,In_1937);
or U130 (N_130,In_53,In_1906);
nand U131 (N_131,In_2104,In_1224);
xor U132 (N_132,In_1750,In_40);
nand U133 (N_133,In_542,In_1129);
and U134 (N_134,In_2435,In_454);
xor U135 (N_135,In_1831,In_1130);
nand U136 (N_136,In_1138,In_590);
or U137 (N_137,In_107,In_1033);
nand U138 (N_138,In_9,In_1648);
nand U139 (N_139,In_1098,In_1057);
and U140 (N_140,In_835,In_1338);
and U141 (N_141,In_1446,In_696);
and U142 (N_142,In_1305,In_2629);
nor U143 (N_143,In_1682,In_355);
or U144 (N_144,In_2290,In_211);
xor U145 (N_145,In_1820,In_2056);
and U146 (N_146,In_1990,In_1345);
and U147 (N_147,In_2808,In_171);
nor U148 (N_148,In_756,In_167);
xnor U149 (N_149,In_1753,In_2233);
nor U150 (N_150,In_288,In_2838);
or U151 (N_151,In_2276,In_1196);
or U152 (N_152,In_1079,In_1848);
nand U153 (N_153,In_320,In_1694);
xor U154 (N_154,In_612,In_2692);
xnor U155 (N_155,In_399,In_667);
and U156 (N_156,In_1195,In_1815);
and U157 (N_157,In_264,In_247);
xnor U158 (N_158,In_2380,In_1481);
xor U159 (N_159,In_2013,In_1748);
nor U160 (N_160,In_159,In_913);
or U161 (N_161,In_1147,In_2100);
and U162 (N_162,In_1337,In_2384);
xnor U163 (N_163,In_2758,In_995);
and U164 (N_164,In_1081,In_721);
nand U165 (N_165,In_1487,In_1180);
nand U166 (N_166,In_2674,In_784);
nand U167 (N_167,In_2913,In_1000);
and U168 (N_168,In_812,In_1787);
and U169 (N_169,In_2087,In_724);
nand U170 (N_170,In_2067,In_2744);
nor U171 (N_171,In_1943,In_2112);
xnor U172 (N_172,In_2422,In_2074);
nand U173 (N_173,In_218,In_746);
nor U174 (N_174,In_2111,In_2684);
nor U175 (N_175,In_1096,In_1769);
or U176 (N_176,In_2482,In_1450);
and U177 (N_177,In_64,In_1477);
nor U178 (N_178,In_351,In_61);
or U179 (N_179,In_1356,In_2521);
nor U180 (N_180,In_1951,In_1778);
nor U181 (N_181,In_1823,In_2649);
or U182 (N_182,In_1510,In_1830);
or U183 (N_183,In_1522,In_1019);
nand U184 (N_184,In_1857,In_2654);
and U185 (N_185,In_400,In_914);
nand U186 (N_186,In_1593,In_1689);
nand U187 (N_187,In_91,In_116);
nand U188 (N_188,In_1893,In_2597);
and U189 (N_189,In_1061,In_1640);
or U190 (N_190,In_803,In_2519);
or U191 (N_191,In_1782,In_2010);
nand U192 (N_192,In_949,In_2240);
and U193 (N_193,In_1295,In_830);
and U194 (N_194,In_2460,In_1811);
or U195 (N_195,In_1836,In_2762);
nand U196 (N_196,In_1794,In_1630);
xnor U197 (N_197,In_1656,In_815);
nand U198 (N_198,In_1382,In_690);
or U199 (N_199,In_446,In_1067);
or U200 (N_200,In_2335,In_2529);
and U201 (N_201,In_1870,In_882);
and U202 (N_202,In_2316,In_2700);
or U203 (N_203,In_1696,In_2251);
nand U204 (N_204,In_2711,In_2315);
nand U205 (N_205,In_1140,In_2553);
or U206 (N_206,In_2222,In_511);
or U207 (N_207,In_2101,In_16);
xnor U208 (N_208,In_170,In_13);
xor U209 (N_209,In_1452,In_2547);
xor U210 (N_210,In_621,In_1297);
nand U211 (N_211,In_1669,In_1244);
and U212 (N_212,In_1235,In_458);
nor U213 (N_213,In_883,In_60);
and U214 (N_214,In_906,In_1786);
or U215 (N_215,In_953,In_263);
nand U216 (N_216,In_420,In_2877);
or U217 (N_217,In_910,In_1797);
or U218 (N_218,In_2036,In_2725);
or U219 (N_219,In_1049,In_1474);
nor U220 (N_220,In_2016,In_2573);
xnor U221 (N_221,In_1422,In_101);
nand U222 (N_222,In_1983,In_1790);
xnor U223 (N_223,In_1183,In_1852);
xor U224 (N_224,In_1217,In_2652);
nand U225 (N_225,In_2392,In_286);
nand U226 (N_226,In_233,In_2329);
or U227 (N_227,In_750,In_2983);
xnor U228 (N_228,In_556,In_839);
nand U229 (N_229,In_1547,In_2468);
or U230 (N_230,In_788,In_1953);
and U231 (N_231,In_1479,In_357);
nand U232 (N_232,In_1208,In_569);
nand U233 (N_233,In_941,In_1484);
or U234 (N_234,In_1955,In_1380);
nor U235 (N_235,In_2050,In_1724);
xnor U236 (N_236,In_2455,In_1904);
nor U237 (N_237,In_816,In_988);
and U238 (N_238,In_996,In_1829);
or U239 (N_239,In_559,In_2898);
nand U240 (N_240,In_1110,In_1563);
or U241 (N_241,In_1454,In_2456);
nand U242 (N_242,In_1229,In_1960);
xor U243 (N_243,In_1458,In_1417);
and U244 (N_244,In_1957,In_2642);
nor U245 (N_245,In_1435,In_1880);
or U246 (N_246,In_2569,In_2352);
xnor U247 (N_247,In_1589,In_412);
or U248 (N_248,In_411,In_1453);
and U249 (N_249,In_1862,In_483);
nor U250 (N_250,In_1974,In_707);
or U251 (N_251,In_2520,In_1525);
and U252 (N_252,In_95,In_2619);
and U253 (N_253,In_627,In_1206);
nand U254 (N_254,In_698,In_2611);
nor U255 (N_255,In_585,In_329);
or U256 (N_256,In_365,In_1250);
nor U257 (N_257,In_2783,In_2601);
xor U258 (N_258,In_2347,In_2492);
and U259 (N_259,In_1069,In_2374);
nor U260 (N_260,In_112,In_98);
and U261 (N_261,In_2285,In_2097);
or U262 (N_262,In_2496,In_1143);
nand U263 (N_263,In_54,In_940);
or U264 (N_264,In_854,In_2952);
nand U265 (N_265,In_2474,In_1959);
xnor U266 (N_266,In_2605,In_2193);
xnor U267 (N_267,In_448,In_881);
or U268 (N_268,In_2914,In_1997);
xnor U269 (N_269,In_2636,In_1392);
nor U270 (N_270,In_1285,In_1569);
or U271 (N_271,In_876,In_276);
nand U272 (N_272,In_2135,In_2218);
nand U273 (N_273,In_2912,In_134);
or U274 (N_274,In_2857,In_1164);
nor U275 (N_275,In_2800,In_600);
nand U276 (N_276,In_1419,In_796);
or U277 (N_277,In_1708,In_1213);
and U278 (N_278,In_524,In_498);
or U279 (N_279,In_248,In_1171);
xor U280 (N_280,In_2923,In_767);
nor U281 (N_281,In_1651,In_1958);
nor U282 (N_282,In_2063,In_2501);
nand U283 (N_283,In_2021,In_782);
and U284 (N_284,In_1238,In_2348);
xor U285 (N_285,In_1492,In_2685);
nor U286 (N_286,In_589,In_1329);
xnor U287 (N_287,In_1799,In_2438);
xnor U288 (N_288,In_2169,In_1888);
nand U289 (N_289,In_1853,In_1363);
xnor U290 (N_290,In_2517,In_965);
or U291 (N_291,In_2598,In_308);
xnor U292 (N_292,In_2498,In_2095);
nor U293 (N_293,In_1083,In_719);
or U294 (N_294,In_262,In_496);
nand U295 (N_295,In_2070,In_2973);
xor U296 (N_296,In_2411,In_747);
nor U297 (N_297,In_1056,In_493);
nor U298 (N_298,In_2357,In_119);
or U299 (N_299,In_126,In_516);
nor U300 (N_300,In_1080,In_2853);
or U301 (N_301,In_32,In_2221);
or U302 (N_302,In_669,In_2264);
xor U303 (N_303,In_1654,In_431);
nand U304 (N_304,In_2327,In_685);
or U305 (N_305,In_97,In_1058);
xor U306 (N_306,In_1760,In_445);
nor U307 (N_307,In_602,In_951);
nor U308 (N_308,In_2687,In_2015);
and U309 (N_309,In_1878,In_1791);
or U310 (N_310,In_2830,In_2234);
nor U311 (N_311,In_890,In_813);
xor U312 (N_312,In_149,In_434);
nand U313 (N_313,In_1298,In_1531);
and U314 (N_314,In_2927,In_1456);
nor U315 (N_315,In_1647,In_2465);
nand U316 (N_316,In_1896,In_662);
xnor U317 (N_317,In_1908,In_717);
and U318 (N_318,In_1894,In_517);
or U319 (N_319,In_44,In_939);
or U320 (N_320,In_1981,In_1875);
nor U321 (N_321,In_1041,In_1802);
nand U322 (N_322,In_2472,In_413);
nand U323 (N_323,In_2564,In_1535);
nand U324 (N_324,In_2541,In_5);
xor U325 (N_325,In_799,In_2382);
or U326 (N_326,In_1471,In_418);
and U327 (N_327,In_804,In_957);
nor U328 (N_328,In_1402,In_1408);
nor U329 (N_329,In_340,In_1695);
nor U330 (N_330,In_853,In_1386);
xor U331 (N_331,In_1844,In_2084);
nor U332 (N_332,In_2425,In_2591);
nand U333 (N_333,In_1642,In_34);
nor U334 (N_334,In_2849,In_2942);
nor U335 (N_335,In_947,In_2888);
or U336 (N_336,In_283,In_1668);
or U337 (N_337,In_2954,In_1362);
nand U338 (N_338,In_2255,In_834);
and U339 (N_339,In_1040,In_2186);
xor U340 (N_340,In_1023,In_1485);
or U341 (N_341,In_1371,In_2918);
and U342 (N_342,In_444,In_1723);
nand U343 (N_343,In_2386,In_2704);
or U344 (N_344,In_2809,In_972);
xnor U345 (N_345,In_1095,In_385);
and U346 (N_346,In_145,In_2887);
nand U347 (N_347,In_2820,In_199);
nand U348 (N_348,In_570,In_1350);
or U349 (N_349,In_2466,In_260);
and U350 (N_350,In_2042,In_765);
and U351 (N_351,In_2975,In_2265);
nand U352 (N_352,In_2275,In_2890);
nand U353 (N_353,In_2726,In_2360);
or U354 (N_354,In_358,In_2612);
and U355 (N_355,In_2933,In_2213);
or U356 (N_356,In_1863,In_1840);
xnor U357 (N_357,In_2493,In_285);
nand U358 (N_358,In_2844,In_1565);
and U359 (N_359,In_325,In_903);
xor U360 (N_360,In_964,In_1429);
or U361 (N_361,In_1734,In_868);
nor U362 (N_362,In_1464,In_1396);
and U363 (N_363,In_1861,In_501);
xor U364 (N_364,In_2944,In_2040);
nand U365 (N_365,In_128,In_1169);
nand U366 (N_366,In_1897,In_2870);
nand U367 (N_367,In_294,In_2593);
nor U368 (N_368,In_635,In_824);
nor U369 (N_369,In_1188,In_2041);
nor U370 (N_370,In_2279,In_715);
or U371 (N_371,In_791,In_2440);
nand U372 (N_372,In_292,In_1635);
or U373 (N_373,In_959,In_2176);
nand U374 (N_374,In_896,In_927);
nor U375 (N_375,In_1381,In_630);
nand U376 (N_376,In_1922,In_2842);
xnor U377 (N_377,In_801,In_1923);
or U378 (N_378,In_2724,In_2209);
xor U379 (N_379,In_689,In_1771);
nor U380 (N_380,In_1882,In_2344);
xnor U381 (N_381,In_1613,In_1762);
xnor U382 (N_382,In_168,In_2818);
nand U383 (N_383,In_1162,In_2833);
nand U384 (N_384,In_1817,In_538);
or U385 (N_385,In_1660,In_215);
or U386 (N_386,In_2986,In_2740);
nor U387 (N_387,In_2854,In_301);
nand U388 (N_388,In_486,In_1042);
nor U389 (N_389,In_1680,In_2977);
nor U390 (N_390,In_2153,In_1307);
nand U391 (N_391,In_23,In_2082);
nand U392 (N_392,In_1663,In_1520);
xor U393 (N_393,In_2280,In_2296);
nor U394 (N_394,In_352,In_611);
or U395 (N_395,In_789,In_2705);
nor U396 (N_396,In_1246,In_2831);
and U397 (N_397,In_380,In_1318);
nor U398 (N_398,In_1288,In_955);
xor U399 (N_399,In_778,In_1373);
or U400 (N_400,In_1555,In_1561);
nand U401 (N_401,In_1361,In_745);
xor U402 (N_402,In_2599,In_1059);
nand U403 (N_403,In_987,In_2079);
or U404 (N_404,In_2834,In_636);
xnor U405 (N_405,In_354,In_625);
or U406 (N_406,In_2781,In_1500);
and U407 (N_407,In_163,In_2281);
nor U408 (N_408,In_1966,In_1533);
xnor U409 (N_409,In_944,In_1043);
xor U410 (N_410,In_684,In_2930);
or U411 (N_411,In_1029,In_1031);
and U412 (N_412,In_557,In_2850);
xnor U413 (N_413,In_67,In_2075);
nor U414 (N_414,In_1239,In_2575);
and U415 (N_415,In_884,In_2215);
or U416 (N_416,In_1330,In_2159);
or U417 (N_417,In_878,In_838);
and U418 (N_418,In_2550,In_1993);
nand U419 (N_419,In_1131,In_1157);
and U420 (N_420,In_1843,In_1789);
xnor U421 (N_421,In_239,In_2478);
xnor U422 (N_422,In_936,In_2772);
nand U423 (N_423,In_737,In_1292);
xor U424 (N_424,In_2346,In_1247);
or U425 (N_425,In_459,In_2443);
xnor U426 (N_426,In_1254,In_2922);
nand U427 (N_427,In_1913,In_2062);
nand U428 (N_428,In_1512,In_2339);
and U429 (N_429,In_1720,In_2542);
or U430 (N_430,In_1742,In_1534);
and U431 (N_431,In_2117,In_1889);
nor U432 (N_432,In_1973,In_2355);
xor U433 (N_433,In_656,In_2058);
xnor U434 (N_434,In_1275,In_392);
xnor U435 (N_435,In_440,In_836);
and U436 (N_436,In_1952,In_2308);
nor U437 (N_437,In_2810,In_2089);
xor U438 (N_438,In_105,In_415);
and U439 (N_439,In_1168,In_402);
or U440 (N_440,In_1874,In_331);
and U441 (N_441,In_2590,In_1917);
nor U442 (N_442,In_2676,In_2856);
and U443 (N_443,In_1409,In_2765);
and U444 (N_444,In_195,In_382);
nor U445 (N_445,In_488,In_2247);
xor U446 (N_446,In_2091,In_552);
or U447 (N_447,In_2829,In_2168);
and U448 (N_448,In_802,In_327);
or U449 (N_449,In_397,In_608);
nand U450 (N_450,In_2710,In_2897);
nand U451 (N_451,In_560,In_309);
xor U452 (N_452,In_500,In_509);
nor U453 (N_453,In_1697,In_1397);
xnor U454 (N_454,In_1703,In_2407);
xnor U455 (N_455,In_2766,In_2814);
xor U456 (N_456,In_1470,In_702);
nand U457 (N_457,In_1804,In_1582);
xor U458 (N_458,In_1366,In_938);
nor U459 (N_459,In_870,In_2866);
and U460 (N_460,In_1657,In_2786);
nand U461 (N_461,In_2925,In_2723);
or U462 (N_462,In_1509,In_35);
and U463 (N_463,In_18,In_558);
or U464 (N_464,In_1100,In_2378);
or U465 (N_465,In_1015,In_848);
nor U466 (N_466,In_1800,In_2336);
nor U467 (N_467,In_565,In_1887);
and U468 (N_468,In_1544,In_564);
nor U469 (N_469,In_663,In_158);
nor U470 (N_470,In_2490,In_2513);
nand U471 (N_471,In_852,In_1113);
xnor U472 (N_472,In_1605,In_2033);
or U473 (N_473,In_2475,In_1030);
or U474 (N_474,In_506,In_332);
xor U475 (N_475,In_1347,In_1914);
or U476 (N_476,In_2263,In_257);
xor U477 (N_477,In_1226,In_907);
nand U478 (N_478,In_1792,In_729);
or U479 (N_479,In_671,In_2261);
and U480 (N_480,In_2165,In_2311);
or U481 (N_481,In_1219,In_1160);
nand U482 (N_482,In_2403,In_180);
and U483 (N_483,In_1681,In_2602);
and U484 (N_484,In_2447,In_1323);
nor U485 (N_485,In_980,In_1093);
or U486 (N_486,In_626,In_477);
xnor U487 (N_487,In_703,In_2409);
nand U488 (N_488,In_2670,In_109);
nand U489 (N_489,In_738,In_1664);
nor U490 (N_490,In_2049,In_322);
or U491 (N_491,In_1616,In_948);
nor U492 (N_492,In_654,In_1442);
or U493 (N_493,In_1210,In_2338);
nand U494 (N_494,In_1145,In_2552);
or U495 (N_495,In_265,In_1652);
xnor U496 (N_496,In_38,In_1949);
nand U497 (N_497,In_874,In_2714);
nand U498 (N_498,In_2841,In_2972);
nor U499 (N_499,In_1600,In_210);
xnor U500 (N_500,In_866,In_1835);
nand U501 (N_501,In_1892,In_615);
and U502 (N_502,In_1883,In_1364);
or U503 (N_503,In_1732,In_245);
nor U504 (N_504,In_1718,In_809);
or U505 (N_505,In_2470,In_2270);
or U506 (N_506,In_2878,In_794);
xnor U507 (N_507,In_1737,In_2127);
and U508 (N_508,In_609,In_2200);
and U509 (N_509,In_539,In_1094);
xnor U510 (N_510,In_678,In_1550);
and U511 (N_511,In_1735,In_1276);
xor U512 (N_512,In_2960,In_2776);
or U513 (N_513,In_2066,In_2886);
nor U514 (N_514,In_731,In_1060);
or U515 (N_515,In_424,In_2543);
xnor U516 (N_516,In_429,In_312);
nor U517 (N_517,In_1349,In_1260);
nand U518 (N_518,In_1225,In_916);
and U519 (N_519,In_2353,In_1249);
and U520 (N_520,In_293,In_1325);
and U521 (N_521,In_983,In_968);
nor U522 (N_522,In_534,In_1071);
nand U523 (N_523,In_1117,In_2982);
and U524 (N_524,In_1570,In_1803);
nor U525 (N_525,In_2163,In_2458);
or U526 (N_526,In_2022,In_1675);
nand U527 (N_527,In_1257,In_388);
nand U528 (N_528,In_2471,In_735);
xor U529 (N_529,In_2530,In_2092);
xor U530 (N_530,In_2194,In_2826);
nor U531 (N_531,In_249,In_2410);
nor U532 (N_532,In_2028,In_435);
nand U533 (N_533,In_2388,In_808);
nor U534 (N_534,In_250,In_2367);
nand U535 (N_535,In_208,In_2356);
nand U536 (N_536,In_2789,In_2915);
xor U537 (N_537,In_1930,In_2910);
xor U538 (N_538,In_686,In_648);
nand U539 (N_539,In_1776,In_1905);
or U540 (N_540,In_2052,In_943);
and U541 (N_541,In_1425,In_770);
nor U542 (N_542,In_1504,In_330);
xor U543 (N_543,In_2875,In_1701);
or U544 (N_544,In_1518,In_1462);
xnor U545 (N_545,In_31,In_2639);
xnor U546 (N_546,In_2437,In_1860);
and U547 (N_547,In_2026,In_640);
nor U548 (N_548,In_1954,In_2429);
nand U549 (N_549,In_253,In_2430);
and U550 (N_550,In_1359,In_1506);
nand U551 (N_551,In_1855,In_1969);
xnor U552 (N_552,In_1965,In_634);
and U553 (N_553,In_1559,In_1369);
xor U554 (N_554,In_182,In_2190);
or U555 (N_555,In_356,In_2769);
xor U556 (N_556,In_2701,In_1536);
xnor U557 (N_557,In_2528,In_2396);
nand U558 (N_558,In_2300,In_2081);
nand U559 (N_559,In_2625,In_1655);
xnor U560 (N_560,In_2978,In_468);
and U561 (N_561,In_469,In_181);
nand U562 (N_562,In_2370,In_2787);
and U563 (N_563,In_1447,In_679);
xnor U564 (N_564,In_754,In_2257);
nand U565 (N_565,In_350,In_1624);
or U566 (N_566,In_2664,In_2752);
nand U567 (N_567,In_1202,In_1673);
nand U568 (N_568,In_1064,In_631);
nor U569 (N_569,In_1667,In_492);
or U570 (N_570,In_2238,In_2749);
or U571 (N_571,In_1466,In_2282);
or U572 (N_572,In_1623,In_280);
or U573 (N_573,In_278,In_2297);
nor U574 (N_574,In_985,In_606);
nor U575 (N_575,In_138,In_701);
and U576 (N_576,In_370,In_1400);
or U577 (N_577,In_246,In_2303);
nand U578 (N_578,In_1666,In_807);
nor U579 (N_579,In_87,In_2256);
nor U580 (N_580,In_2561,In_1743);
xor U581 (N_581,In_1384,In_1856);
nor U582 (N_582,In_443,In_2170);
nand U583 (N_583,In_1932,In_2462);
xnor U584 (N_584,In_1612,In_1702);
nor U585 (N_585,In_2909,In_394);
nand U586 (N_586,In_2709,In_1076);
nor U587 (N_587,In_1166,In_1261);
nor U588 (N_588,In_2046,In_409);
xnor U589 (N_589,In_1399,In_2120);
nand U590 (N_590,In_1854,In_1335);
xor U591 (N_591,In_1228,In_2548);
and U592 (N_592,In_236,In_1410);
or U593 (N_593,In_637,In_1876);
and U594 (N_594,In_1401,In_919);
xor U595 (N_595,In_2034,In_2340);
nor U596 (N_596,In_572,In_992);
xor U597 (N_597,In_2061,In_1780);
or U598 (N_598,In_1716,In_1818);
nor U599 (N_599,In_2955,In_1503);
nor U600 (N_600,In_920,In_1967);
or U601 (N_601,In_1733,In_225);
or U602 (N_602,In_2006,In_2249);
nand U603 (N_603,In_2879,In_2373);
xnor U604 (N_604,In_2505,In_2819);
and U605 (N_605,In_1314,In_374);
nor U606 (N_606,In_505,In_1010);
nand U607 (N_607,In_63,In_3);
nand U608 (N_608,In_2269,In_1596);
nand U609 (N_609,In_1788,In_2996);
xor U610 (N_610,In_2242,In_1199);
xor U611 (N_611,In_2628,In_1391);
nand U612 (N_612,In_1432,In_1119);
xor U613 (N_613,In_1726,In_305);
xor U614 (N_614,In_114,In_555);
nand U615 (N_615,In_2354,In_677);
nand U616 (N_616,In_2051,In_2584);
nand U617 (N_617,In_2963,In_2503);
and U618 (N_618,In_387,In_700);
nor U619 (N_619,In_1197,In_1622);
or U620 (N_620,In_610,In_1252);
or U621 (N_621,In_1721,In_136);
xor U622 (N_622,In_2557,In_873);
nor U623 (N_623,In_1601,In_1112);
or U624 (N_624,In_2936,In_484);
nor U625 (N_625,In_2959,In_2119);
nand U626 (N_626,In_4,In_449);
nor U627 (N_627,In_213,In_2231);
xor U628 (N_628,In_2720,In_764);
nand U629 (N_629,In_1573,In_50);
nor U630 (N_630,In_2463,In_1333);
and U631 (N_631,In_1459,In_1813);
or U632 (N_632,In_974,In_1713);
or U633 (N_633,In_727,In_1457);
and U634 (N_634,In_2065,In_2495);
or U635 (N_635,In_725,In_1850);
nor U636 (N_636,In_688,In_216);
xnor U637 (N_637,In_108,In_732);
or U638 (N_638,In_1181,In_1016);
xor U639 (N_639,In_1389,In_895);
xnor U640 (N_640,In_90,In_472);
xor U641 (N_641,In_668,In_1977);
xor U642 (N_642,In_193,In_2735);
nor U643 (N_643,In_1312,In_1841);
nand U644 (N_644,In_2402,In_343);
and U645 (N_645,In_43,In_2232);
nor U646 (N_646,In_2871,In_19);
nor U647 (N_647,In_1267,In_942);
nand U648 (N_648,In_892,In_2489);
xor U649 (N_649,In_1137,In_1255);
and U650 (N_650,In_2372,In_2566);
and U651 (N_651,In_2659,In_638);
nand U652 (N_652,In_1572,In_1032);
xnor U653 (N_653,In_401,In_1837);
xnor U654 (N_654,In_632,In_2733);
nand U655 (N_655,In_2939,In_137);
nand U656 (N_656,In_1744,In_763);
xnor U657 (N_657,In_1628,In_2736);
or U658 (N_658,In_536,In_1475);
and U659 (N_659,In_2747,In_1483);
xnor U660 (N_660,In_275,In_1931);
or U661 (N_661,In_2361,In_277);
and U662 (N_662,In_818,In_183);
nor U663 (N_663,In_2855,In_926);
nand U664 (N_664,In_2461,In_1984);
nand U665 (N_665,In_1839,In_1440);
or U666 (N_666,In_1286,In_172);
and U667 (N_667,In_2990,In_1756);
and U668 (N_668,In_2540,In_2906);
xor U669 (N_669,In_823,In_1269);
xor U670 (N_670,In_1822,In_533);
xor U671 (N_671,In_2071,In_335);
or U672 (N_672,In_1944,In_1587);
nand U673 (N_673,In_21,In_2985);
nand U674 (N_674,In_872,In_2934);
xor U675 (N_675,In_2568,In_1236);
or U676 (N_676,In_2469,In_201);
nor U677 (N_677,In_202,In_2207);
and U678 (N_678,In_337,In_1764);
or U679 (N_679,In_2884,In_1300);
and U680 (N_680,In_1087,In_845);
and U681 (N_681,In_1832,In_2577);
xnor U682 (N_682,In_841,In_20);
and U683 (N_683,In_2860,In_2739);
and U684 (N_684,In_437,In_2405);
and U685 (N_685,In_1428,In_1476);
xnor U686 (N_686,In_978,In_425);
xnor U687 (N_687,In_2731,In_2309);
or U688 (N_688,In_2477,In_580);
nand U689 (N_689,In_571,In_2858);
xnor U690 (N_690,In_973,In_85);
xor U691 (N_691,In_176,In_83);
and U692 (N_692,In_178,In_1941);
and U693 (N_693,In_1927,In_935);
and U694 (N_694,In_404,In_1690);
xnor U695 (N_695,In_1879,In_1537);
and U696 (N_696,In_2487,In_470);
xnor U697 (N_697,In_2214,In_2730);
nand U698 (N_698,In_2531,In_2729);
or U699 (N_699,In_912,In_2341);
nor U700 (N_700,In_75,In_2394);
nand U701 (N_701,In_2,In_2572);
nand U702 (N_702,In_1607,In_2932);
and U703 (N_703,In_1938,In_1178);
or U704 (N_704,In_1620,In_2518);
and U705 (N_705,In_1678,In_1414);
or U706 (N_706,In_2287,In_797);
xnor U707 (N_707,In_1480,In_1747);
nand U708 (N_708,In_1551,In_2105);
or U709 (N_709,In_156,In_2208);
nand U710 (N_710,In_51,In_2574);
or U711 (N_711,In_2681,In_2620);
nor U712 (N_712,In_1496,In_14);
or U713 (N_713,In_1173,In_317);
xor U714 (N_714,In_837,In_489);
or U715 (N_715,In_2152,In_1999);
or U716 (N_716,In_2244,In_1631);
nor U717 (N_717,In_774,In_1772);
and U718 (N_718,In_1686,In_1436);
nand U719 (N_719,In_859,In_1158);
or U720 (N_720,In_1185,In_2417);
and U721 (N_721,In_1560,In_2130);
and U722 (N_722,In_933,In_1465);
xor U723 (N_723,In_1871,In_17);
and U724 (N_724,In_891,In_2272);
or U725 (N_725,In_197,In_646);
nand U726 (N_726,In_11,In_2031);
nor U727 (N_727,In_1731,In_768);
nand U728 (N_728,In_115,In_1528);
or U729 (N_729,In_368,In_2502);
and U730 (N_730,In_1271,In_2230);
xor U731 (N_731,In_428,In_6);
nor U732 (N_732,In_2608,In_281);
and U733 (N_733,In_2454,In_1146);
or U734 (N_734,In_1327,In_2780);
and U735 (N_735,In_1051,In_2734);
or U736 (N_736,In_578,In_2640);
and U737 (N_737,In_255,In_256);
or U738 (N_738,In_1727,In_775);
nand U739 (N_739,In_1890,In_1121);
xnor U740 (N_740,In_1519,In_1736);
or U741 (N_741,In_2656,In_92);
and U742 (N_742,In_241,In_1545);
nand U743 (N_743,In_1478,In_1405);
or U744 (N_744,In_682,In_1441);
nor U745 (N_745,In_1141,In_2797);
and U746 (N_746,In_1986,In_577);
nor U747 (N_747,In_575,In_645);
and U748 (N_748,In_595,In_94);
and U749 (N_749,In_2643,In_886);
or U750 (N_750,In_1821,In_174);
or U751 (N_751,In_805,In_1864);
xnor U752 (N_752,In_2246,In_1714);
or U753 (N_753,In_692,In_1413);
xor U754 (N_754,In_162,In_1634);
and U755 (N_755,In_647,In_683);
nand U756 (N_756,In_2988,In_2096);
nand U757 (N_757,In_2647,In_1976);
and U758 (N_758,In_2741,In_2266);
or U759 (N_759,In_2174,In_2172);
xnor U760 (N_760,In_2510,In_877);
nand U761 (N_761,In_526,In_1189);
nor U762 (N_762,In_1578,In_598);
nand U763 (N_763,In_1513,In_36);
nand U764 (N_764,In_333,In_1182);
xor U765 (N_765,In_2002,In_88);
nor U766 (N_766,In_1490,In_2423);
xnor U767 (N_767,In_2054,In_2997);
nor U768 (N_768,In_1526,In_952);
nand U769 (N_769,In_2162,In_2668);
and U770 (N_770,In_2651,In_1115);
and U771 (N_771,In_1026,In_244);
or U772 (N_772,In_2313,In_1992);
nand U773 (N_773,In_2483,In_2142);
nand U774 (N_774,In_1045,In_766);
nor U775 (N_775,In_2928,In_1916);
or U776 (N_776,In_152,In_652);
nor U777 (N_777,In_1637,In_2150);
and U778 (N_778,In_1167,In_2432);
nand U779 (N_779,In_1240,In_2072);
or U780 (N_780,In_1116,In_694);
or U781 (N_781,In_177,In_367);
xor U782 (N_782,In_2949,In_2514);
nand U783 (N_783,In_800,In_2024);
nand U784 (N_784,In_1370,In_2160);
and U785 (N_785,In_1289,In_742);
xnor U786 (N_786,In_2839,In_528);
and U787 (N_787,In_2554,In_1847);
nor U788 (N_788,In_1746,In_2099);
or U789 (N_789,In_1451,In_2931);
nor U790 (N_790,In_2334,In_2312);
nand U791 (N_791,In_272,In_2248);
nand U792 (N_792,In_1877,In_2774);
nor U793 (N_793,In_432,In_793);
or U794 (N_794,In_103,In_644);
xnor U795 (N_795,In_49,In_2406);
or U796 (N_796,In_1299,In_863);
nor U797 (N_797,In_596,In_2412);
xnor U798 (N_798,In_1282,In_1204);
or U799 (N_799,In_2807,In_1684);
and U800 (N_800,In_1092,In_2464);
nand U801 (N_801,In_41,In_2827);
or U802 (N_802,In_672,In_1109);
xor U803 (N_803,In_1963,In_1154);
nand U804 (N_804,In_2821,In_364);
and U805 (N_805,In_2424,In_2239);
nand U806 (N_806,In_30,In_2166);
nand U807 (N_807,In_377,In_922);
and U808 (N_808,In_2110,In_2603);
xor U809 (N_809,In_2522,In_1586);
and U810 (N_810,In_2707,In_2235);
xnor U811 (N_811,In_1174,In_771);
nand U812 (N_812,In_867,In_499);
or U813 (N_813,In_2785,In_706);
nor U814 (N_814,In_2721,In_485);
and U815 (N_815,In_545,In_850);
nor U816 (N_816,In_617,In_12);
and U817 (N_817,In_2951,In_2702);
nand U818 (N_818,In_2565,In_1427);
and U819 (N_819,In_1050,In_405);
nor U820 (N_820,In_2005,In_2921);
and U821 (N_821,In_1599,In_1626);
and U822 (N_822,In_10,In_56);
nor U823 (N_823,In_510,In_2359);
xnor U824 (N_824,In_2717,In_269);
nor U825 (N_825,In_476,In_2459);
nor U826 (N_826,In_2641,In_408);
nand U827 (N_827,In_1378,In_2206);
nand U828 (N_828,In_934,In_2480);
xor U829 (N_829,In_1403,In_315);
xnor U830 (N_830,In_494,In_1842);
nor U831 (N_831,In_2945,In_2499);
nand U832 (N_832,In_1209,In_1002);
nand U833 (N_833,In_597,In_2189);
nor U834 (N_834,In_1988,In_2895);
nor U835 (N_835,In_1426,In_2967);
nor U836 (N_836,In_826,In_2948);
and U837 (N_837,In_1670,In_1898);
and U838 (N_838,In_655,In_2157);
nand U839 (N_839,In_676,In_918);
and U840 (N_840,In_588,In_1343);
and U841 (N_841,In_1,In_2790);
nand U842 (N_842,In_2715,In_2880);
nand U843 (N_843,In_194,In_1558);
nand U844 (N_844,In_1712,In_1779);
nor U845 (N_845,In_79,In_781);
nor U846 (N_846,In_2236,In_2038);
nand U847 (N_847,In_1136,In_207);
xor U848 (N_848,In_1352,In_2728);
nand U849 (N_849,In_1745,In_1309);
or U850 (N_850,In_1473,In_1674);
nor U851 (N_851,In_2148,In_2332);
nand U852 (N_852,In_433,In_2673);
or U853 (N_853,In_1604,In_2648);
nand U854 (N_854,In_2795,In_1200);
or U855 (N_855,In_651,In_2549);
nor U856 (N_856,In_2134,In_344);
xnor U857 (N_857,In_2862,In_2136);
or U858 (N_858,In_455,In_1806);
and U859 (N_859,In_1676,In_334);
or U860 (N_860,In_1054,In_1048);
nand U861 (N_861,In_2784,In_899);
or U862 (N_862,In_366,In_849);
nor U863 (N_863,In_2507,In_2175);
or U864 (N_864,In_1028,In_1082);
nand U865 (N_865,In_2000,In_33);
nand U866 (N_866,In_855,In_1819);
nor U867 (N_867,In_1387,In_1920);
nand U868 (N_868,In_261,In_436);
nand U869 (N_869,In_2712,In_512);
nor U870 (N_870,In_1606,In_1590);
nand U871 (N_871,In_2420,In_2008);
nand U872 (N_872,In_2203,In_1348);
nand U873 (N_873,In_1705,In_1006);
xnor U874 (N_874,In_427,In_295);
nand U875 (N_875,In_2003,In_58);
nand U876 (N_876,In_1302,In_1499);
nand U877 (N_877,In_946,In_1482);
nand U878 (N_878,In_915,In_2421);
nand U879 (N_879,In_2210,In_2196);
xor U880 (N_880,In_954,In_2623);
nand U881 (N_881,In_2118,In_1165);
or U882 (N_882,In_1472,In_282);
nor U883 (N_883,In_2580,In_131);
nor U884 (N_884,In_2616,In_1948);
xnor U885 (N_885,In_709,In_504);
xor U886 (N_886,In_820,In_48);
and U887 (N_887,In_165,In_1542);
nand U888 (N_888,In_1935,In_2801);
nand U889 (N_889,In_894,In_1849);
and U890 (N_890,In_1207,In_889);
nor U891 (N_891,In_160,In_711);
or U892 (N_892,In_697,In_1598);
and U893 (N_893,In_1218,In_2748);
nand U894 (N_894,In_1120,In_1388);
nor U895 (N_895,In_908,In_1037);
or U896 (N_896,In_1929,In_1758);
nand U897 (N_897,In_2292,In_231);
xnor U898 (N_898,In_1017,In_2125);
or U899 (N_899,In_284,In_1242);
and U900 (N_900,In_2761,In_2581);
nor U901 (N_901,In_1406,In_2538);
xor U902 (N_902,In_2293,In_2337);
or U903 (N_903,In_324,In_1541);
nand U904 (N_904,In_2164,In_100);
and U905 (N_905,In_71,In_1615);
or U906 (N_906,In_1014,In_2587);
and U907 (N_907,In_2326,In_665);
nor U908 (N_908,In_773,In_924);
nand U909 (N_909,In_441,In_130);
or U910 (N_910,In_1728,In_2610);
nor U911 (N_911,In_1638,In_251);
nand U912 (N_912,In_1766,In_787);
nand U913 (N_913,In_643,In_204);
xor U914 (N_914,In_1296,In_1975);
nor U915 (N_915,In_2745,In_1968);
or U916 (N_916,In_2289,In_561);
nor U917 (N_917,In_1956,In_1084);
nor U918 (N_918,In_1310,In_2799);
nor U919 (N_919,In_2947,In_1704);
and U920 (N_920,In_553,In_1592);
nand U921 (N_921,In_2350,In_898);
nor U922 (N_922,In_1741,In_2788);
and U923 (N_923,In_2299,In_2385);
or U924 (N_924,In_618,In_2138);
or U925 (N_925,In_1099,In_579);
xor U926 (N_926,In_179,In_381);
nand U927 (N_927,In_2904,In_229);
nand U928 (N_928,In_649,In_2379);
nor U929 (N_929,In_1272,In_1424);
nor U930 (N_930,In_1700,In_2305);
and U931 (N_931,In_624,In_417);
nor U932 (N_932,In_2223,In_614);
or U933 (N_933,In_930,In_2250);
nand U934 (N_934,In_353,In_1303);
nor U935 (N_935,In_1996,In_2252);
nand U936 (N_936,In_1527,In_547);
and U937 (N_937,In_2404,In_2273);
or U938 (N_938,In_313,In_221);
nor U939 (N_939,In_345,In_120);
and U940 (N_940,In_2375,In_228);
nand U941 (N_941,In_2782,In_937);
nand U942 (N_942,In_1653,In_2794);
xor U943 (N_943,In_129,In_111);
xnor U944 (N_944,In_760,In_1773);
or U945 (N_945,In_2228,In_144);
and U946 (N_946,In_22,In_2812);
and U947 (N_947,In_226,In_541);
xnor U948 (N_948,In_1075,In_785);
or U949 (N_949,In_2322,In_1430);
or U950 (N_950,In_2307,In_2328);
xnor U951 (N_951,In_2607,In_1194);
and U952 (N_952,In_2563,In_398);
and U953 (N_953,In_2102,In_1073);
nor U954 (N_954,In_291,In_1679);
or U955 (N_955,In_761,In_1358);
nor U956 (N_956,In_1132,In_1749);
xor U957 (N_957,In_592,In_2645);
nand U958 (N_958,In_2080,In_1066);
nand U959 (N_959,In_2703,In_348);
and U960 (N_960,In_1175,In_2824);
and U961 (N_961,In_2562,In_89);
nand U962 (N_962,In_2773,In_2693);
and U963 (N_963,In_1947,In_2631);
and U964 (N_964,In_2383,In_1283);
or U965 (N_965,In_1671,In_2434);
or U966 (N_966,In_2211,In_1866);
nor U967 (N_967,In_982,In_829);
nand U968 (N_968,In_658,In_1699);
or U969 (N_969,In_1089,In_1434);
and U970 (N_970,In_2644,In_2516);
nor U971 (N_971,In_2393,In_2690);
nand U972 (N_972,In_1108,In_76);
nand U973 (N_973,In_1911,In_2718);
or U974 (N_974,In_2943,In_554);
or U975 (N_975,In_604,In_1306);
or U976 (N_976,In_1891,In_2484);
nor U977 (N_977,In_2064,In_1463);
or U978 (N_978,In_1259,In_223);
nor U979 (N_979,In_1774,In_2381);
nor U980 (N_980,In_2527,In_2260);
or U981 (N_981,In_1468,In_1761);
xnor U982 (N_982,In_2271,In_2185);
or U983 (N_983,In_1872,In_549);
nand U984 (N_984,In_1915,In_1557);
nor U985 (N_985,In_2863,In_1543);
or U986 (N_986,In_1564,In_1757);
xor U987 (N_987,In_993,In_673);
nand U988 (N_988,In_2414,In_185);
or U989 (N_989,In_2624,In_196);
and U990 (N_990,In_1961,In_846);
or U991 (N_991,In_143,In_2147);
nand U992 (N_992,In_1658,In_562);
nor U993 (N_993,In_2060,In_2476);
nand U994 (N_994,In_2399,In_2570);
nand U995 (N_995,In_1245,In_1317);
nor U996 (N_996,In_2600,In_1825);
or U997 (N_997,In_2791,In_1262);
or U998 (N_998,In_230,In_491);
and U999 (N_999,In_2039,In_1783);
nor U1000 (N_1000,In_346,In_1985);
or U1001 (N_1001,In_403,In_2803);
and U1002 (N_1002,In_777,In_2226);
xnor U1003 (N_1003,In_2446,In_2428);
nor U1004 (N_1004,In_339,In_1062);
nor U1005 (N_1005,In_1964,In_2155);
and U1006 (N_1006,In_2001,In_1411);
and U1007 (N_1007,In_2323,In_2901);
nand U1008 (N_1008,In_2321,In_287);
xor U1009 (N_1009,In_790,In_1970);
xor U1010 (N_1010,In_1237,In_971);
or U1011 (N_1011,In_310,In_1725);
nor U1012 (N_1012,In_2220,In_1594);
or U1013 (N_1013,In_77,In_1012);
and U1014 (N_1014,In_240,In_1768);
nand U1015 (N_1015,In_1777,In_1304);
xor U1016 (N_1016,In_2188,In_1291);
and U1017 (N_1017,In_389,In_1105);
xor U1018 (N_1018,In_2995,In_2678);
or U1019 (N_1019,In_2695,In_238);
nand U1020 (N_1020,In_2442,In_1311);
or U1021 (N_1021,In_2453,In_2698);
or U1022 (N_1022,In_1730,In_307);
and U1023 (N_1023,In_2151,In_2515);
or U1024 (N_1024,In_1796,In_2672);
and U1025 (N_1025,In_901,In_416);
or U1026 (N_1026,In_986,In_328);
nand U1027 (N_1027,In_819,In_862);
and U1028 (N_1028,In_1365,In_1319);
xnor U1029 (N_1029,In_2991,In_806);
and U1030 (N_1030,In_271,In_831);
and U1031 (N_1031,In_1277,In_1460);
nand U1032 (N_1032,In_1583,In_2876);
nor U1033 (N_1033,In_1212,In_1287);
xor U1034 (N_1034,In_59,In_2764);
nor U1035 (N_1035,In_1576,In_929);
and U1036 (N_1036,In_613,In_319);
or U1037 (N_1037,In_1994,In_2694);
xnor U1038 (N_1038,In_2146,In_661);
xor U1039 (N_1039,In_8,In_2713);
nand U1040 (N_1040,In_857,In_616);
nand U1041 (N_1041,In_1566,In_2768);
nor U1042 (N_1042,In_2004,In_1603);
and U1043 (N_1043,In_2926,In_78);
nor U1044 (N_1044,In_962,In_893);
nand U1045 (N_1045,In_2364,In_1070);
and U1046 (N_1046,In_2043,In_206);
nand U1047 (N_1047,In_1431,In_1900);
xor U1048 (N_1048,In_817,In_2179);
nand U1049 (N_1049,In_1332,In_2746);
nor U1050 (N_1050,In_2343,In_161);
and U1051 (N_1051,In_1144,In_2161);
xnor U1052 (N_1052,In_235,In_1502);
or U1053 (N_1053,In_2950,In_191);
xnor U1054 (N_1054,In_1633,In_1858);
xnor U1055 (N_1055,In_2588,In_576);
nand U1056 (N_1056,In_2667,In_718);
nor U1057 (N_1057,In_1785,In_1201);
or U1058 (N_1058,In_391,In_2298);
and U1059 (N_1059,In_2397,In_963);
xor U1060 (N_1060,In_209,In_2467);
and U1061 (N_1061,In_1610,In_1106);
nand U1062 (N_1062,In_753,In_1339);
or U1063 (N_1063,In_2771,In_148);
and U1064 (N_1064,In_2893,In_1602);
nand U1065 (N_1065,In_1022,In_1448);
nor U1066 (N_1066,In_714,In_1585);
xor U1067 (N_1067,In_755,In_1186);
xor U1068 (N_1068,In_2219,In_723);
nand U1069 (N_1069,In_410,In_2675);
xor U1070 (N_1070,In_546,In_1316);
xor U1071 (N_1071,In_856,In_2582);
or U1072 (N_1072,In_1627,In_2488);
xnor U1073 (N_1073,In_419,In_1775);
nor U1074 (N_1074,In_1577,In_2689);
or U1075 (N_1075,In_1135,In_660);
xnor U1076 (N_1076,In_2961,In_361);
or U1077 (N_1077,In_1123,In_1177);
and U1078 (N_1078,In_151,In_452);
nor U1079 (N_1079,In_426,In_675);
xor U1080 (N_1080,In_2145,In_1097);
and U1081 (N_1081,In_1685,In_1461);
nand U1082 (N_1082,In_2088,In_2030);
and U1083 (N_1083,In_2660,In_406);
nand U1084 (N_1084,In_1107,In_2408);
and U1085 (N_1085,In_471,In_1007);
and U1086 (N_1086,In_798,In_1151);
nor U1087 (N_1087,In_2957,In_2415);
xnor U1088 (N_1088,In_2377,In_1672);
and U1089 (N_1089,In_2365,In_591);
and U1090 (N_1090,In_99,In_518);
xor U1091 (N_1091,In_2864,In_521);
nor U1092 (N_1092,In_1340,In_1379);
or U1093 (N_1093,In_102,In_375);
nand U1094 (N_1094,In_2665,In_594);
or U1095 (N_1095,In_373,In_1584);
or U1096 (N_1096,In_487,In_1580);
or U1097 (N_1097,In_1025,In_2535);
or U1098 (N_1098,In_1416,In_2419);
and U1099 (N_1099,In_1579,In_1517);
nand U1100 (N_1100,In_2555,In_480);
nor U1101 (N_1101,In_758,In_2376);
nor U1102 (N_1102,In_2661,In_1643);
and U1103 (N_1103,In_460,In_1867);
nand U1104 (N_1104,In_704,In_222);
nor U1105 (N_1105,In_1385,In_2902);
or U1106 (N_1106,In_342,In_2816);
xor U1107 (N_1107,In_1521,In_2680);
xor U1108 (N_1108,In_132,In_217);
or U1109 (N_1109,In_2055,In_495);
nor U1110 (N_1110,In_1415,In_2832);
nor U1111 (N_1111,In_1940,In_1808);
and U1112 (N_1112,In_82,In_52);
nor U1113 (N_1113,In_642,In_279);
or U1114 (N_1114,In_1505,In_1065);
and U1115 (N_1115,In_2450,In_1611);
nor U1116 (N_1116,In_989,In_2525);
and U1117 (N_1117,In_2216,In_135);
or U1118 (N_1118,In_1326,In_2989);
and U1119 (N_1119,In_2342,In_2971);
nand U1120 (N_1120,In_748,In_1232);
nor U1121 (N_1121,In_2722,In_363);
xor U1122 (N_1122,In_2903,In_2286);
nand U1123 (N_1123,In_465,In_582);
nor U1124 (N_1124,In_2872,In_1614);
or U1125 (N_1125,In_2546,In_2390);
nand U1126 (N_1126,In_326,In_961);
xor U1127 (N_1127,In_2626,In_740);
nand U1128 (N_1128,In_2882,In_1278);
nor U1129 (N_1129,In_2500,In_2937);
xnor U1130 (N_1130,In_2094,In_439);
xor U1131 (N_1131,In_623,In_1706);
or U1132 (N_1132,In_2627,In_2699);
nor U1133 (N_1133,In_1812,In_1187);
nor U1134 (N_1134,In_786,In_2613);
nor U1135 (N_1135,In_2441,In_1104);
nand U1136 (N_1136,In_2288,In_1568);
xor U1137 (N_1137,In_2753,In_2558);
xor U1138 (N_1138,In_970,In_393);
xnor U1139 (N_1139,In_2199,In_822);
nand U1140 (N_1140,In_2485,In_1418);
nor U1141 (N_1141,In_2045,In_2325);
xnor U1142 (N_1142,In_2301,In_2556);
nor U1143 (N_1143,In_188,In_759);
nor U1144 (N_1144,In_395,In_2044);
xnor U1145 (N_1145,In_2294,In_1553);
nand U1146 (N_1146,In_2198,In_376);
and U1147 (N_1147,In_1412,In_2126);
or U1148 (N_1148,In_1895,In_386);
or U1149 (N_1149,In_827,In_7);
xnor U1150 (N_1150,In_527,In_1223);
and U1151 (N_1151,In_2941,In_2691);
nor U1152 (N_1152,In_2848,In_2032);
and U1153 (N_1153,In_2770,In_1609);
nand U1154 (N_1154,In_2793,In_2141);
and U1155 (N_1155,In_2113,In_998);
nand U1156 (N_1156,In_1036,In_442);
xnor U1157 (N_1157,In_1540,In_1619);
nand U1158 (N_1158,In_880,In_2320);
nand U1159 (N_1159,In_2486,In_674);
or U1160 (N_1160,In_55,In_121);
nand U1161 (N_1161,In_1443,In_2953);
xnor U1162 (N_1162,In_2304,In_175);
nand U1163 (N_1163,In_450,In_629);
nor U1164 (N_1164,In_1221,In_2144);
and U1165 (N_1165,In_2653,In_1989);
xnor U1166 (N_1166,In_2609,In_2756);
xor U1167 (N_1167,In_1024,In_1126);
or U1168 (N_1168,In_169,In_1995);
and U1169 (N_1169,In_1793,In_2537);
xnor U1170 (N_1170,In_86,In_2837);
xor U1171 (N_1171,In_273,In_2090);
and U1172 (N_1172,In_166,In_1290);
nand U1173 (N_1173,In_593,In_2992);
xnor U1174 (N_1174,In_2202,In_1234);
nor U1175 (N_1175,In_833,In_396);
nor U1176 (N_1176,In_1918,In_653);
nor U1177 (N_1177,In_302,In_1845);
and U1178 (N_1178,In_2427,In_1375);
or U1179 (N_1179,In_1677,In_917);
or U1180 (N_1180,In_733,In_1523);
xor U1181 (N_1181,In_2413,In_967);
nand U1182 (N_1182,In_2835,In_1574);
and U1183 (N_1183,In_925,In_2180);
and U1184 (N_1184,In_192,In_220);
and U1185 (N_1185,In_1102,In_2823);
and U1186 (N_1186,In_1936,In_2594);
nor U1187 (N_1187,In_1376,In_2278);
or U1188 (N_1188,In_2401,In_15);
nor U1189 (N_1189,In_212,In_2716);
nor U1190 (N_1190,In_29,In_154);
or U1191 (N_1191,In_1814,In_945);
xnor U1192 (N_1192,In_2217,In_2205);
nand U1193 (N_1193,In_2682,In_254);
and U1194 (N_1194,In_2178,In_252);
xnor U1195 (N_1195,In_2596,In_1881);
xnor U1196 (N_1196,In_27,In_2362);
nand U1197 (N_1197,In_290,In_1754);
and U1198 (N_1198,In_1227,In_1192);
or U1199 (N_1199,In_2633,In_2122);
xor U1200 (N_1200,In_2655,In_728);
nand U1201 (N_1201,In_1495,In_1394);
nand U1202 (N_1202,In_2846,In_1395);
nand U1203 (N_1203,In_1336,In_1341);
and U1204 (N_1204,In_960,In_2539);
xnor U1205 (N_1205,In_515,In_2938);
or U1206 (N_1206,In_810,In_2245);
nand U1207 (N_1207,In_2935,In_2622);
xnor U1208 (N_1208,In_2173,In_769);
and U1209 (N_1209,In_2868,In_2494);
and U1210 (N_1210,In_1155,In_2606);
and U1211 (N_1211,In_1280,In_1215);
or U1212 (N_1212,In_1331,In_2007);
nand U1213 (N_1213,In_605,In_2589);
or U1214 (N_1214,In_1148,In_2851);
xnor U1215 (N_1215,In_730,In_1739);
and U1216 (N_1216,In_2836,In_466);
xor U1217 (N_1217,In_422,In_1538);
nor U1218 (N_1218,In_447,In_205);
xor U1219 (N_1219,In_1205,In_2604);
xor U1220 (N_1220,In_1004,In_633);
nor U1221 (N_1221,In_1324,In_828);
xor U1222 (N_1222,In_1608,In_2268);
xnor U1223 (N_1223,In_1013,In_2592);
or U1224 (N_1224,In_2369,In_2181);
nor U1225 (N_1225,In_1910,In_1884);
nor U1226 (N_1226,In_117,In_1859);
nand U1227 (N_1227,In_423,In_520);
nor U1228 (N_1228,In_1507,In_1270);
or U1229 (N_1229,In_1149,In_70);
xor U1230 (N_1230,In_2391,In_490);
nand U1231 (N_1231,In_74,In_259);
or U1232 (N_1232,In_1090,In_2187);
nor U1233 (N_1233,In_1575,In_2677);
or U1234 (N_1234,In_2197,In_2869);
nand U1235 (N_1235,In_1816,In_299);
and U1236 (N_1236,In_1661,In_349);
or U1237 (N_1237,In_1740,In_2805);
nor U1238 (N_1238,In_659,In_523);
xnor U1239 (N_1239,In_1444,In_1907);
or U1240 (N_1240,In_710,In_1265);
nor U1241 (N_1241,In_1945,In_1597);
nor U1242 (N_1242,In_153,In_371);
or U1243 (N_1243,In_2047,In_563);
xnor U1244 (N_1244,In_1170,In_1489);
xnor U1245 (N_1245,In_414,In_2743);
nand U1246 (N_1246,In_2751,In_481);
and U1247 (N_1247,In_2129,In_1567);
nor U1248 (N_1248,In_268,In_1233);
xor U1249 (N_1249,In_1909,In_1809);
nand U1250 (N_1250,In_1824,In_843);
xor U1251 (N_1251,In_2666,In_2132);
xnor U1252 (N_1252,In_1636,In_2968);
or U1253 (N_1253,In_2984,In_1134);
or U1254 (N_1254,In_2306,In_2014);
xnor U1255 (N_1255,In_507,In_622);
xnor U1256 (N_1256,In_921,In_1552);
and U1257 (N_1257,In_1072,In_540);
or U1258 (N_1258,In_463,In_586);
xor U1259 (N_1259,In_1693,In_670);
and U1260 (N_1260,In_2201,In_1784);
xor U1261 (N_1261,In_347,In_2057);
and U1262 (N_1262,In_2883,In_1868);
xnor U1263 (N_1263,In_875,In_2974);
xor U1264 (N_1264,In_1991,In_783);
xor U1265 (N_1265,In_267,In_2237);
nand U1266 (N_1266,In_2526,In_1063);
or U1267 (N_1267,In_1253,In_532);
and U1268 (N_1268,In_2907,In_2225);
and U1269 (N_1269,In_2426,In_1038);
xnor U1270 (N_1270,In_390,In_2585);
nand U1271 (N_1271,In_548,In_2980);
nand U1272 (N_1272,In_1497,In_869);
or U1273 (N_1273,In_1508,In_2137);
nor U1274 (N_1274,In_383,In_2184);
xor U1275 (N_1275,In_186,In_1342);
or U1276 (N_1276,In_2128,In_858);
nor U1277 (N_1277,In_1176,In_911);
xor U1278 (N_1278,In_306,In_864);
and U1279 (N_1279,In_203,In_1085);
nand U1280 (N_1280,In_567,In_2970);
or U1281 (N_1281,In_2114,In_2366);
and U1282 (N_1282,In_45,In_1933);
nor U1283 (N_1283,In_2349,In_879);
xnor U1284 (N_1284,In_1301,In_2183);
nor U1285 (N_1285,In_2669,In_1281);
and U1286 (N_1286,In_2618,In_513);
and U1287 (N_1287,In_296,In_2009);
or U1288 (N_1288,In_1111,In_2908);
nand U1289 (N_1289,In_1738,In_2840);
and U1290 (N_1290,In_772,In_2657);
or U1291 (N_1291,In_2267,In_2018);
nor U1292 (N_1292,In_2241,In_1279);
or U1293 (N_1293,In_1709,In_2999);
nor U1294 (N_1294,In_1826,In_1179);
and U1295 (N_1295,In_525,In_573);
nand U1296 (N_1296,In_2508,In_780);
or U1297 (N_1297,In_2436,In_2258);
and U1298 (N_1298,In_42,In_1554);
nand U1299 (N_1299,In_1190,In_1230);
nand U1300 (N_1300,In_976,In_551);
nand U1301 (N_1301,In_84,In_1514);
and U1302 (N_1302,In_316,In_2284);
xnor U1303 (N_1303,In_336,In_1827);
nand U1304 (N_1304,In_1711,In_1346);
and U1305 (N_1305,In_2994,In_68);
nor U1306 (N_1306,In_2433,In_2107);
xnor U1307 (N_1307,In_2509,In_1902);
xnor U1308 (N_1308,In_2919,In_57);
nand U1309 (N_1309,In_25,In_1039);
and U1310 (N_1310,In_1360,In_997);
xor U1311 (N_1311,In_1707,In_266);
and U1312 (N_1312,In_2534,In_932);
nand U1313 (N_1313,In_2663,In_2881);
nor U1314 (N_1314,In_1268,In_2697);
xnor U1315 (N_1315,In_2544,In_237);
or U1316 (N_1316,In_2536,In_214);
nor U1317 (N_1317,In_811,In_1191);
xor U1318 (N_1318,In_713,In_1828);
nor U1319 (N_1319,In_2439,In_2560);
or U1320 (N_1320,In_303,In_1869);
xnor U1321 (N_1321,In_1077,In_1632);
nor U1322 (N_1322,In_2905,In_1320);
and U1323 (N_1323,In_1801,In_2892);
and U1324 (N_1324,In_1114,In_2637);
or U1325 (N_1325,In_2760,In_666);
xnor U1326 (N_1326,In_66,In_1924);
nand U1327 (N_1327,In_1449,In_1851);
xnor U1328 (N_1328,In_2124,In_2946);
nor U1329 (N_1329,In_1539,In_1184);
xor U1330 (N_1330,In_2389,In_1729);
and U1331 (N_1331,In_1001,In_2859);
and U1332 (N_1332,In_323,In_122);
and U1333 (N_1333,In_599,In_2479);
or U1334 (N_1334,In_680,In_224);
xor U1335 (N_1335,In_118,In_2894);
nand U1336 (N_1336,In_2671,In_1163);
nor U1337 (N_1337,In_1912,In_1998);
nand U1338 (N_1338,In_461,In_1055);
nor U1339 (N_1339,In_2330,In_2011);
xnor U1340 (N_1340,In_2109,In_726);
xnor U1341 (N_1341,In_362,In_1498);
nand U1342 (N_1342,In_716,In_2302);
or U1343 (N_1343,In_603,In_2843);
nand U1344 (N_1344,In_2368,In_1795);
nor U1345 (N_1345,In_842,In_2775);
nor U1346 (N_1346,In_923,In_2195);
or U1347 (N_1347,In_451,In_274);
nand U1348 (N_1348,In_2025,In_584);
nand U1349 (N_1349,In_2576,In_1127);
xor U1350 (N_1350,In_360,In_26);
and U1351 (N_1351,In_497,In_1294);
and U1352 (N_1352,In_695,In_2140);
xor U1353 (N_1353,In_421,In_888);
xor U1354 (N_1354,In_1798,In_378);
nor U1355 (N_1355,In_1256,In_187);
or U1356 (N_1356,In_139,In_529);
xnor U1357 (N_1357,In_1770,In_311);
xor U1358 (N_1358,In_2767,In_321);
or U1359 (N_1359,In_189,In_865);
xnor U1360 (N_1360,In_1919,In_950);
xnor U1361 (N_1361,In_2763,In_1765);
and U1362 (N_1362,In_2243,In_2116);
and U1363 (N_1363,In_1501,In_1216);
nand U1364 (N_1364,In_2177,In_1390);
xor U1365 (N_1365,In_430,In_905);
or U1366 (N_1366,In_2759,In_2683);
xnor U1367 (N_1367,In_1710,In_2351);
nor U1368 (N_1368,In_1946,In_2632);
and U1369 (N_1369,In_270,In_146);
xnor U1370 (N_1370,In_1355,In_1715);
xnor U1371 (N_1371,In_314,In_2156);
or U1372 (N_1372,In_2171,In_69);
and U1373 (N_1373,In_1751,In_2523);
xnor U1374 (N_1374,In_1763,In_2085);
or U1375 (N_1375,In_2363,In_1020);
nand U1376 (N_1376,In_1404,In_2987);
or U1377 (N_1377,In_2998,In_104);
xnor U1378 (N_1378,In_1979,In_2154);
and U1379 (N_1379,In_140,In_1124);
or U1380 (N_1380,In_219,In_587);
or U1381 (N_1381,In_1274,In_2358);
nor U1382 (N_1382,In_190,In_1437);
xor U1383 (N_1383,In_2192,In_776);
xor U1384 (N_1384,In_110,In_1241);
nor U1385 (N_1385,In_2037,In_2874);
or U1386 (N_1386,In_2889,In_2817);
and U1387 (N_1387,In_1971,In_2059);
nand U1388 (N_1388,In_2481,In_2545);
nand U1389 (N_1389,In_1511,In_227);
and U1390 (N_1390,In_757,In_1328);
and U1391 (N_1391,In_1650,In_574);
nand U1392 (N_1392,In_1068,In_2865);
nor U1393 (N_1393,In_2891,In_2149);
nor U1394 (N_1394,In_1018,In_535);
nand U1395 (N_1395,In_751,In_1962);
nor U1396 (N_1396,In_2811,In_2778);
or U1397 (N_1397,In_2845,In_990);
nand U1398 (N_1398,In_300,In_1982);
xnor U1399 (N_1399,In_1044,In_832);
xnor U1400 (N_1400,In_2696,In_1052);
xor U1401 (N_1401,In_359,In_379);
xor U1402 (N_1402,In_369,In_530);
nor U1403 (N_1403,In_568,In_2317);
nor U1404 (N_1404,In_2708,In_720);
and U1405 (N_1405,In_1939,In_639);
nor U1406 (N_1406,In_583,In_2452);
nor U1407 (N_1407,In_1243,In_1591);
xnor U1408 (N_1408,In_999,In_543);
or U1409 (N_1409,In_1248,In_1047);
nand U1410 (N_1410,In_1899,In_1088);
and U1411 (N_1411,In_664,In_1807);
or U1412 (N_1412,In_1251,In_2331);
nor U1413 (N_1413,In_0,In_1172);
nand U1414 (N_1414,In_1752,In_1009);
and U1415 (N_1415,In_1344,In_2524);
and U1416 (N_1416,In_1284,In_2445);
and U1417 (N_1417,In_372,In_909);
and U1418 (N_1418,In_1264,In_1659);
or U1419 (N_1419,In_482,In_897);
or U1420 (N_1420,In_2121,In_531);
xnor U1421 (N_1421,In_1621,In_2815);
or U1422 (N_1422,In_779,In_124);
nand U1423 (N_1423,In_384,In_1649);
nand U1424 (N_1424,In_1515,In_1125);
nand U1425 (N_1425,In_1003,In_2131);
or U1426 (N_1426,In_232,In_1838);
nor U1427 (N_1427,In_860,In_1722);
and U1428 (N_1428,In_1445,In_2431);
nand U1429 (N_1429,In_1942,In_722);
nand U1430 (N_1430,In_2444,In_687);
or U1431 (N_1431,In_2035,In_2291);
xnor U1432 (N_1432,In_2262,In_2254);
nor U1433 (N_1433,In_164,In_2048);
or U1434 (N_1434,In_502,In_1334);
xor U1435 (N_1435,In_473,In_1488);
and U1436 (N_1436,In_2106,In_1618);
xnor U1437 (N_1437,In_1639,In_2093);
nand U1438 (N_1438,In_1231,In_81);
and U1439 (N_1439,In_2076,In_1101);
nor U1440 (N_1440,In_1091,In_2806);
and U1441 (N_1441,In_2448,In_1903);
nor U1442 (N_1442,In_2719,In_1027);
nor U1443 (N_1443,In_1322,In_2191);
xor U1444 (N_1444,In_519,In_844);
or U1445 (N_1445,In_1008,In_1273);
nand U1446 (N_1446,In_1493,In_1972);
nand U1447 (N_1447,In_1921,In_1313);
xnor U1448 (N_1448,In_200,In_885);
and U1449 (N_1449,In_2825,In_1926);
nor U1450 (N_1450,In_24,In_2283);
or U1451 (N_1451,In_1372,In_1315);
xnor U1452 (N_1452,In_2387,In_1150);
and U1453 (N_1453,In_2083,In_2686);
and U1454 (N_1454,In_2757,In_155);
and U1455 (N_1455,In_1034,In_2491);
or U1456 (N_1456,In_1781,In_1987);
or U1457 (N_1457,In_1767,In_2755);
or U1458 (N_1458,In_2295,In_1665);
xnor U1459 (N_1459,In_2029,In_752);
xor U1460 (N_1460,In_2899,In_2133);
and U1461 (N_1461,In_1377,In_1549);
and U1462 (N_1462,In_931,In_2956);
xor U1463 (N_1463,In_2617,In_851);
xnor U1464 (N_1464,In_1641,In_739);
and U1465 (N_1465,In_2310,In_2012);
xnor U1466 (N_1466,In_242,In_1901);
nand U1467 (N_1467,In_2742,In_478);
nor U1468 (N_1468,In_1755,In_2086);
nor U1469 (N_1469,In_1491,In_2227);
and U1470 (N_1470,In_2314,In_1351);
and U1471 (N_1471,In_2395,In_1805);
nand U1472 (N_1472,In_861,In_2103);
or U1473 (N_1473,In_1078,In_1308);
or U1474 (N_1474,In_1139,In_234);
xnor U1475 (N_1475,In_2053,In_1354);
nor U1476 (N_1476,In_2253,In_1455);
or U1477 (N_1477,In_2277,In_1516);
and U1478 (N_1478,In_681,In_2143);
and U1479 (N_1479,In_2646,In_2964);
xor U1480 (N_1480,In_467,In_1469);
nor U1481 (N_1481,In_1142,In_106);
nand U1482 (N_1482,In_1934,In_1420);
nand U1483 (N_1483,In_464,In_2457);
and U1484 (N_1484,In_2259,In_650);
or U1485 (N_1485,In_2497,In_902);
nor U1486 (N_1486,In_1950,In_1211);
and U1487 (N_1487,In_1293,In_157);
or U1488 (N_1488,In_1086,In_1529);
nor U1489 (N_1489,In_1005,In_1258);
or U1490 (N_1490,In_2418,In_304);
and U1491 (N_1491,In_1846,In_1886);
and U1492 (N_1492,In_2635,In_1439);
or U1493 (N_1493,In_2578,In_2688);
nand U1494 (N_1494,In_2123,In_1159);
nor U1495 (N_1495,In_958,In_984);
xor U1496 (N_1496,In_2981,In_705);
nand U1497 (N_1497,In_1266,In_125);
nor U1498 (N_1498,In_1865,In_438);
nand U1499 (N_1499,In_2911,In_1810);
and U1500 (N_1500,In_458,In_153);
nand U1501 (N_1501,In_2166,In_2268);
xnor U1502 (N_1502,In_263,In_882);
and U1503 (N_1503,In_6,In_1841);
nor U1504 (N_1504,In_1452,In_84);
nand U1505 (N_1505,In_2274,In_2091);
nand U1506 (N_1506,In_2306,In_1890);
or U1507 (N_1507,In_1250,In_2521);
xnor U1508 (N_1508,In_869,In_2360);
nand U1509 (N_1509,In_1402,In_2502);
nand U1510 (N_1510,In_2209,In_1139);
nand U1511 (N_1511,In_2103,In_1928);
and U1512 (N_1512,In_79,In_2312);
xnor U1513 (N_1513,In_396,In_1451);
and U1514 (N_1514,In_83,In_1839);
nand U1515 (N_1515,In_1662,In_471);
or U1516 (N_1516,In_2667,In_2060);
xnor U1517 (N_1517,In_1367,In_177);
nor U1518 (N_1518,In_2201,In_2014);
nand U1519 (N_1519,In_887,In_1419);
nor U1520 (N_1520,In_745,In_1432);
or U1521 (N_1521,In_1352,In_2996);
nand U1522 (N_1522,In_484,In_2913);
nor U1523 (N_1523,In_2715,In_2545);
xnor U1524 (N_1524,In_2097,In_2989);
nor U1525 (N_1525,In_1903,In_1645);
nor U1526 (N_1526,In_2774,In_2381);
xor U1527 (N_1527,In_1330,In_1684);
and U1528 (N_1528,In_43,In_1742);
and U1529 (N_1529,In_436,In_2139);
xnor U1530 (N_1530,In_1930,In_2991);
nand U1531 (N_1531,In_1923,In_2719);
and U1532 (N_1532,In_46,In_1060);
and U1533 (N_1533,In_833,In_152);
and U1534 (N_1534,In_1754,In_1261);
nor U1535 (N_1535,In_2436,In_2003);
nor U1536 (N_1536,In_2322,In_1059);
xnor U1537 (N_1537,In_2968,In_628);
nor U1538 (N_1538,In_726,In_2001);
nor U1539 (N_1539,In_2210,In_2701);
or U1540 (N_1540,In_625,In_1717);
xor U1541 (N_1541,In_379,In_2640);
nor U1542 (N_1542,In_374,In_1366);
nand U1543 (N_1543,In_651,In_756);
nor U1544 (N_1544,In_2503,In_1787);
nor U1545 (N_1545,In_2648,In_2099);
and U1546 (N_1546,In_333,In_266);
and U1547 (N_1547,In_2321,In_1948);
nor U1548 (N_1548,In_697,In_1017);
and U1549 (N_1549,In_268,In_1625);
or U1550 (N_1550,In_955,In_2122);
xnor U1551 (N_1551,In_1811,In_2540);
nand U1552 (N_1552,In_2418,In_2733);
and U1553 (N_1553,In_654,In_2859);
or U1554 (N_1554,In_13,In_1696);
nand U1555 (N_1555,In_969,In_460);
nor U1556 (N_1556,In_736,In_1928);
nor U1557 (N_1557,In_12,In_2414);
or U1558 (N_1558,In_1943,In_300);
nand U1559 (N_1559,In_2221,In_1396);
xnor U1560 (N_1560,In_1548,In_726);
or U1561 (N_1561,In_722,In_278);
nand U1562 (N_1562,In_866,In_1032);
or U1563 (N_1563,In_1375,In_27);
or U1564 (N_1564,In_2958,In_1708);
or U1565 (N_1565,In_2458,In_528);
and U1566 (N_1566,In_1487,In_1916);
and U1567 (N_1567,In_1550,In_2174);
or U1568 (N_1568,In_2451,In_512);
or U1569 (N_1569,In_315,In_201);
or U1570 (N_1570,In_2475,In_984);
nor U1571 (N_1571,In_1472,In_932);
nor U1572 (N_1572,In_2810,In_405);
nor U1573 (N_1573,In_2627,In_118);
and U1574 (N_1574,In_1915,In_2968);
xnor U1575 (N_1575,In_92,In_1940);
and U1576 (N_1576,In_2428,In_1551);
nand U1577 (N_1577,In_2667,In_715);
nor U1578 (N_1578,In_2605,In_531);
xor U1579 (N_1579,In_729,In_1565);
nor U1580 (N_1580,In_817,In_611);
nand U1581 (N_1581,In_1663,In_1544);
nor U1582 (N_1582,In_139,In_315);
and U1583 (N_1583,In_460,In_278);
or U1584 (N_1584,In_2198,In_2013);
or U1585 (N_1585,In_148,In_1592);
nand U1586 (N_1586,In_1058,In_152);
or U1587 (N_1587,In_661,In_1768);
nand U1588 (N_1588,In_431,In_1088);
or U1589 (N_1589,In_71,In_1971);
xnor U1590 (N_1590,In_1560,In_2056);
xnor U1591 (N_1591,In_1607,In_2977);
nand U1592 (N_1592,In_1468,In_425);
nand U1593 (N_1593,In_153,In_315);
xnor U1594 (N_1594,In_1289,In_757);
xnor U1595 (N_1595,In_789,In_2916);
nand U1596 (N_1596,In_2720,In_571);
nand U1597 (N_1597,In_1600,In_97);
nand U1598 (N_1598,In_2087,In_2401);
nand U1599 (N_1599,In_1164,In_748);
xnor U1600 (N_1600,In_342,In_2987);
nor U1601 (N_1601,In_1534,In_2529);
or U1602 (N_1602,In_145,In_998);
nor U1603 (N_1603,In_2596,In_983);
nor U1604 (N_1604,In_983,In_2710);
nand U1605 (N_1605,In_376,In_605);
and U1606 (N_1606,In_295,In_1974);
and U1607 (N_1607,In_1358,In_2645);
and U1608 (N_1608,In_2101,In_510);
xor U1609 (N_1609,In_2984,In_362);
and U1610 (N_1610,In_1362,In_1009);
xnor U1611 (N_1611,In_1758,In_360);
and U1612 (N_1612,In_352,In_535);
nor U1613 (N_1613,In_1568,In_2785);
nor U1614 (N_1614,In_2046,In_1462);
nand U1615 (N_1615,In_557,In_2262);
xor U1616 (N_1616,In_2410,In_1936);
or U1617 (N_1617,In_1727,In_2853);
or U1618 (N_1618,In_2422,In_983);
or U1619 (N_1619,In_2685,In_2379);
xnor U1620 (N_1620,In_1220,In_2349);
nor U1621 (N_1621,In_1910,In_2712);
nor U1622 (N_1622,In_159,In_2065);
xor U1623 (N_1623,In_1255,In_2178);
nand U1624 (N_1624,In_1284,In_1575);
xor U1625 (N_1625,In_1459,In_2639);
and U1626 (N_1626,In_2643,In_2141);
and U1627 (N_1627,In_1850,In_2786);
or U1628 (N_1628,In_727,In_433);
nand U1629 (N_1629,In_139,In_318);
or U1630 (N_1630,In_2076,In_2886);
and U1631 (N_1631,In_1034,In_1123);
and U1632 (N_1632,In_454,In_1292);
nor U1633 (N_1633,In_716,In_2920);
xnor U1634 (N_1634,In_221,In_1976);
or U1635 (N_1635,In_782,In_101);
nor U1636 (N_1636,In_1510,In_958);
or U1637 (N_1637,In_2746,In_2863);
and U1638 (N_1638,In_374,In_2287);
or U1639 (N_1639,In_2646,In_1245);
or U1640 (N_1640,In_1147,In_437);
and U1641 (N_1641,In_118,In_2561);
xor U1642 (N_1642,In_674,In_893);
xor U1643 (N_1643,In_2218,In_1829);
or U1644 (N_1644,In_2436,In_1568);
nor U1645 (N_1645,In_2830,In_96);
and U1646 (N_1646,In_1568,In_3);
xnor U1647 (N_1647,In_2549,In_1952);
nand U1648 (N_1648,In_2681,In_2926);
xor U1649 (N_1649,In_1308,In_2184);
nand U1650 (N_1650,In_1331,In_894);
nor U1651 (N_1651,In_2254,In_1988);
nand U1652 (N_1652,In_8,In_1410);
xnor U1653 (N_1653,In_25,In_1546);
nor U1654 (N_1654,In_1280,In_2458);
and U1655 (N_1655,In_598,In_1703);
nor U1656 (N_1656,In_114,In_1230);
and U1657 (N_1657,In_1922,In_2764);
or U1658 (N_1658,In_1743,In_2703);
nand U1659 (N_1659,In_1018,In_2958);
nor U1660 (N_1660,In_1229,In_1246);
and U1661 (N_1661,In_1620,In_2754);
xnor U1662 (N_1662,In_854,In_1073);
nor U1663 (N_1663,In_1304,In_464);
nor U1664 (N_1664,In_1523,In_2562);
or U1665 (N_1665,In_167,In_2554);
or U1666 (N_1666,In_1233,In_572);
and U1667 (N_1667,In_601,In_593);
or U1668 (N_1668,In_141,In_674);
nor U1669 (N_1669,In_1665,In_1657);
or U1670 (N_1670,In_1041,In_972);
or U1671 (N_1671,In_230,In_550);
xnor U1672 (N_1672,In_594,In_1412);
nand U1673 (N_1673,In_591,In_2939);
and U1674 (N_1674,In_723,In_427);
xor U1675 (N_1675,In_1468,In_910);
nor U1676 (N_1676,In_153,In_644);
and U1677 (N_1677,In_1068,In_2406);
nor U1678 (N_1678,In_2828,In_1264);
and U1679 (N_1679,In_208,In_2556);
xnor U1680 (N_1680,In_1108,In_2326);
or U1681 (N_1681,In_393,In_1641);
nand U1682 (N_1682,In_259,In_2512);
nor U1683 (N_1683,In_1725,In_2963);
or U1684 (N_1684,In_164,In_2943);
nor U1685 (N_1685,In_386,In_2159);
nor U1686 (N_1686,In_2463,In_2667);
or U1687 (N_1687,In_1202,In_1678);
and U1688 (N_1688,In_680,In_2328);
or U1689 (N_1689,In_2005,In_1327);
and U1690 (N_1690,In_829,In_987);
xnor U1691 (N_1691,In_2489,In_632);
or U1692 (N_1692,In_782,In_970);
nor U1693 (N_1693,In_1547,In_735);
nor U1694 (N_1694,In_2174,In_1379);
nand U1695 (N_1695,In_2956,In_1625);
xnor U1696 (N_1696,In_427,In_2637);
or U1697 (N_1697,In_2566,In_2865);
or U1698 (N_1698,In_1848,In_1976);
nor U1699 (N_1699,In_2139,In_2566);
or U1700 (N_1700,In_822,In_2887);
xnor U1701 (N_1701,In_1080,In_50);
and U1702 (N_1702,In_1045,In_1832);
nand U1703 (N_1703,In_1328,In_2028);
xnor U1704 (N_1704,In_2965,In_402);
and U1705 (N_1705,In_2558,In_2386);
nor U1706 (N_1706,In_2731,In_1754);
and U1707 (N_1707,In_1271,In_1735);
nand U1708 (N_1708,In_61,In_462);
nor U1709 (N_1709,In_948,In_1708);
or U1710 (N_1710,In_411,In_933);
nor U1711 (N_1711,In_1453,In_2647);
nor U1712 (N_1712,In_1971,In_866);
nor U1713 (N_1713,In_162,In_300);
and U1714 (N_1714,In_666,In_766);
nand U1715 (N_1715,In_1441,In_1252);
xor U1716 (N_1716,In_1561,In_1103);
xnor U1717 (N_1717,In_2732,In_397);
nor U1718 (N_1718,In_709,In_2612);
nand U1719 (N_1719,In_970,In_2420);
xor U1720 (N_1720,In_196,In_509);
nand U1721 (N_1721,In_1082,In_361);
and U1722 (N_1722,In_2873,In_1766);
xnor U1723 (N_1723,In_1063,In_783);
or U1724 (N_1724,In_2128,In_502);
nor U1725 (N_1725,In_1695,In_1291);
nand U1726 (N_1726,In_1751,In_2584);
nand U1727 (N_1727,In_2260,In_1544);
xor U1728 (N_1728,In_1585,In_1896);
nand U1729 (N_1729,In_927,In_773);
xor U1730 (N_1730,In_2675,In_1807);
xor U1731 (N_1731,In_2617,In_1033);
nand U1732 (N_1732,In_970,In_2161);
nand U1733 (N_1733,In_1819,In_853);
nand U1734 (N_1734,In_484,In_2454);
or U1735 (N_1735,In_2360,In_126);
nor U1736 (N_1736,In_811,In_716);
nand U1737 (N_1737,In_2093,In_2289);
nor U1738 (N_1738,In_2561,In_9);
xor U1739 (N_1739,In_1644,In_504);
xnor U1740 (N_1740,In_2298,In_2041);
or U1741 (N_1741,In_492,In_2377);
nor U1742 (N_1742,In_1256,In_379);
nand U1743 (N_1743,In_2237,In_1623);
xor U1744 (N_1744,In_2405,In_1213);
nand U1745 (N_1745,In_1425,In_1177);
xnor U1746 (N_1746,In_2601,In_2677);
nor U1747 (N_1747,In_956,In_2088);
xor U1748 (N_1748,In_2254,In_1237);
xnor U1749 (N_1749,In_2035,In_2523);
xnor U1750 (N_1750,In_2846,In_2534);
xnor U1751 (N_1751,In_1756,In_2425);
xor U1752 (N_1752,In_878,In_1867);
nor U1753 (N_1753,In_762,In_2092);
and U1754 (N_1754,In_485,In_2328);
and U1755 (N_1755,In_1385,In_1226);
xor U1756 (N_1756,In_1090,In_2196);
xnor U1757 (N_1757,In_2537,In_174);
and U1758 (N_1758,In_2326,In_917);
xnor U1759 (N_1759,In_1316,In_1072);
or U1760 (N_1760,In_2713,In_2158);
xor U1761 (N_1761,In_1326,In_1968);
or U1762 (N_1762,In_544,In_1359);
or U1763 (N_1763,In_1719,In_2113);
xnor U1764 (N_1764,In_2286,In_2367);
and U1765 (N_1765,In_1163,In_2772);
and U1766 (N_1766,In_1700,In_874);
nor U1767 (N_1767,In_370,In_674);
and U1768 (N_1768,In_2037,In_2741);
nor U1769 (N_1769,In_711,In_2672);
nor U1770 (N_1770,In_219,In_148);
nand U1771 (N_1771,In_2451,In_2067);
or U1772 (N_1772,In_1610,In_2160);
and U1773 (N_1773,In_1549,In_718);
xor U1774 (N_1774,In_429,In_1063);
and U1775 (N_1775,In_2157,In_1436);
or U1776 (N_1776,In_525,In_2488);
xor U1777 (N_1777,In_2576,In_1156);
xor U1778 (N_1778,In_13,In_2643);
nand U1779 (N_1779,In_549,In_2120);
xor U1780 (N_1780,In_1446,In_2342);
and U1781 (N_1781,In_2713,In_2367);
or U1782 (N_1782,In_2660,In_1539);
nor U1783 (N_1783,In_1069,In_2262);
or U1784 (N_1784,In_2561,In_340);
xor U1785 (N_1785,In_2783,In_670);
xnor U1786 (N_1786,In_1967,In_2463);
or U1787 (N_1787,In_45,In_52);
xor U1788 (N_1788,In_1765,In_1473);
or U1789 (N_1789,In_418,In_2457);
xor U1790 (N_1790,In_1923,In_2806);
or U1791 (N_1791,In_278,In_599);
or U1792 (N_1792,In_2580,In_639);
nand U1793 (N_1793,In_1299,In_741);
nor U1794 (N_1794,In_2261,In_2221);
nand U1795 (N_1795,In_156,In_857);
and U1796 (N_1796,In_2571,In_2952);
nor U1797 (N_1797,In_798,In_522);
xnor U1798 (N_1798,In_1969,In_2569);
or U1799 (N_1799,In_515,In_578);
or U1800 (N_1800,In_1613,In_850);
or U1801 (N_1801,In_138,In_2987);
or U1802 (N_1802,In_2935,In_1272);
nor U1803 (N_1803,In_441,In_2862);
or U1804 (N_1804,In_2757,In_1321);
xnor U1805 (N_1805,In_2924,In_1651);
nand U1806 (N_1806,In_1378,In_1384);
nand U1807 (N_1807,In_2002,In_1168);
or U1808 (N_1808,In_2503,In_1195);
nor U1809 (N_1809,In_2090,In_799);
nand U1810 (N_1810,In_2023,In_2528);
xnor U1811 (N_1811,In_2580,In_457);
nand U1812 (N_1812,In_2836,In_2522);
or U1813 (N_1813,In_2568,In_2523);
nor U1814 (N_1814,In_2839,In_49);
and U1815 (N_1815,In_1487,In_20);
nor U1816 (N_1816,In_2680,In_1158);
and U1817 (N_1817,In_1197,In_1975);
xor U1818 (N_1818,In_455,In_50);
and U1819 (N_1819,In_2035,In_888);
nand U1820 (N_1820,In_1441,In_660);
or U1821 (N_1821,In_1452,In_115);
xor U1822 (N_1822,In_2999,In_2417);
xnor U1823 (N_1823,In_70,In_686);
xnor U1824 (N_1824,In_699,In_2722);
or U1825 (N_1825,In_1598,In_1579);
nor U1826 (N_1826,In_1232,In_1607);
and U1827 (N_1827,In_1461,In_604);
or U1828 (N_1828,In_674,In_939);
nand U1829 (N_1829,In_945,In_776);
nor U1830 (N_1830,In_1797,In_699);
xor U1831 (N_1831,In_2231,In_2833);
nor U1832 (N_1832,In_2295,In_2999);
xor U1833 (N_1833,In_2061,In_2977);
and U1834 (N_1834,In_2968,In_1384);
xor U1835 (N_1835,In_2573,In_907);
and U1836 (N_1836,In_370,In_815);
or U1837 (N_1837,In_1236,In_1938);
xnor U1838 (N_1838,In_664,In_30);
nand U1839 (N_1839,In_2981,In_277);
nand U1840 (N_1840,In_1116,In_2441);
nor U1841 (N_1841,In_1974,In_836);
xnor U1842 (N_1842,In_1702,In_2771);
xnor U1843 (N_1843,In_1266,In_1601);
nand U1844 (N_1844,In_1666,In_224);
or U1845 (N_1845,In_665,In_467);
or U1846 (N_1846,In_2712,In_2070);
nor U1847 (N_1847,In_510,In_1270);
or U1848 (N_1848,In_2717,In_2317);
nor U1849 (N_1849,In_1032,In_935);
nor U1850 (N_1850,In_595,In_2058);
nand U1851 (N_1851,In_476,In_291);
or U1852 (N_1852,In_2826,In_1022);
nand U1853 (N_1853,In_1938,In_2808);
xnor U1854 (N_1854,In_942,In_1763);
xor U1855 (N_1855,In_1318,In_1889);
nor U1856 (N_1856,In_147,In_2916);
nor U1857 (N_1857,In_2873,In_383);
nor U1858 (N_1858,In_215,In_2703);
nor U1859 (N_1859,In_423,In_2579);
nand U1860 (N_1860,In_1345,In_2558);
and U1861 (N_1861,In_1922,In_461);
xor U1862 (N_1862,In_2763,In_57);
and U1863 (N_1863,In_803,In_1624);
xor U1864 (N_1864,In_162,In_1051);
or U1865 (N_1865,In_767,In_2162);
nor U1866 (N_1866,In_2699,In_2018);
and U1867 (N_1867,In_190,In_1797);
nor U1868 (N_1868,In_378,In_903);
nand U1869 (N_1869,In_2215,In_228);
nor U1870 (N_1870,In_531,In_1953);
and U1871 (N_1871,In_1404,In_2893);
nand U1872 (N_1872,In_1699,In_2462);
xnor U1873 (N_1873,In_1117,In_2791);
or U1874 (N_1874,In_1512,In_2636);
and U1875 (N_1875,In_571,In_2869);
nor U1876 (N_1876,In_806,In_1489);
xnor U1877 (N_1877,In_1871,In_2681);
nor U1878 (N_1878,In_1972,In_2485);
xnor U1879 (N_1879,In_591,In_628);
xnor U1880 (N_1880,In_1143,In_832);
or U1881 (N_1881,In_125,In_1898);
or U1882 (N_1882,In_265,In_2527);
nand U1883 (N_1883,In_543,In_502);
nor U1884 (N_1884,In_230,In_1512);
nor U1885 (N_1885,In_869,In_1217);
nand U1886 (N_1886,In_2463,In_1082);
and U1887 (N_1887,In_1002,In_1951);
xor U1888 (N_1888,In_70,In_531);
or U1889 (N_1889,In_527,In_2029);
nor U1890 (N_1890,In_2434,In_203);
and U1891 (N_1891,In_2730,In_2710);
xnor U1892 (N_1892,In_817,In_678);
nand U1893 (N_1893,In_2345,In_1890);
or U1894 (N_1894,In_487,In_1402);
xnor U1895 (N_1895,In_1310,In_2956);
xnor U1896 (N_1896,In_751,In_399);
or U1897 (N_1897,In_2886,In_457);
and U1898 (N_1898,In_2244,In_1451);
or U1899 (N_1899,In_517,In_931);
nor U1900 (N_1900,In_2543,In_2922);
nand U1901 (N_1901,In_518,In_1893);
nand U1902 (N_1902,In_1968,In_1300);
and U1903 (N_1903,In_2847,In_272);
nand U1904 (N_1904,In_2844,In_277);
nor U1905 (N_1905,In_2003,In_2577);
or U1906 (N_1906,In_1713,In_1463);
nand U1907 (N_1907,In_2954,In_2804);
and U1908 (N_1908,In_2732,In_1801);
nor U1909 (N_1909,In_1544,In_244);
nor U1910 (N_1910,In_21,In_249);
and U1911 (N_1911,In_2932,In_480);
or U1912 (N_1912,In_557,In_762);
xor U1913 (N_1913,In_217,In_2431);
nand U1914 (N_1914,In_1039,In_598);
or U1915 (N_1915,In_413,In_2349);
nand U1916 (N_1916,In_2927,In_2983);
nor U1917 (N_1917,In_2915,In_1399);
and U1918 (N_1918,In_1967,In_2107);
nand U1919 (N_1919,In_442,In_87);
or U1920 (N_1920,In_2145,In_1898);
xor U1921 (N_1921,In_2243,In_2216);
nor U1922 (N_1922,In_2649,In_2315);
or U1923 (N_1923,In_2093,In_759);
xor U1924 (N_1924,In_2149,In_1412);
nand U1925 (N_1925,In_2964,In_1609);
xnor U1926 (N_1926,In_362,In_1206);
xnor U1927 (N_1927,In_485,In_2882);
or U1928 (N_1928,In_368,In_1808);
xnor U1929 (N_1929,In_848,In_366);
nand U1930 (N_1930,In_2369,In_156);
xor U1931 (N_1931,In_265,In_946);
xor U1932 (N_1932,In_161,In_1277);
nand U1933 (N_1933,In_443,In_892);
and U1934 (N_1934,In_954,In_2500);
and U1935 (N_1935,In_1705,In_2758);
or U1936 (N_1936,In_923,In_1951);
and U1937 (N_1937,In_1319,In_360);
and U1938 (N_1938,In_183,In_858);
and U1939 (N_1939,In_2802,In_2020);
nand U1940 (N_1940,In_187,In_1175);
and U1941 (N_1941,In_1497,In_739);
nand U1942 (N_1942,In_2291,In_582);
and U1943 (N_1943,In_1456,In_200);
nand U1944 (N_1944,In_729,In_2092);
nand U1945 (N_1945,In_2860,In_1345);
and U1946 (N_1946,In_819,In_167);
xnor U1947 (N_1947,In_763,In_1683);
xor U1948 (N_1948,In_1128,In_222);
or U1949 (N_1949,In_1110,In_322);
xor U1950 (N_1950,In_108,In_7);
nand U1951 (N_1951,In_2140,In_1877);
nor U1952 (N_1952,In_12,In_1391);
nor U1953 (N_1953,In_1898,In_1051);
nor U1954 (N_1954,In_1475,In_1758);
nand U1955 (N_1955,In_1886,In_1495);
xor U1956 (N_1956,In_1234,In_580);
or U1957 (N_1957,In_448,In_1919);
nand U1958 (N_1958,In_1953,In_302);
nand U1959 (N_1959,In_1469,In_1985);
nand U1960 (N_1960,In_1155,In_2450);
xor U1961 (N_1961,In_2881,In_542);
nor U1962 (N_1962,In_1064,In_1219);
nand U1963 (N_1963,In_224,In_2054);
nor U1964 (N_1964,In_1158,In_380);
xor U1965 (N_1965,In_1195,In_2969);
or U1966 (N_1966,In_2201,In_2667);
and U1967 (N_1967,In_66,In_1605);
nand U1968 (N_1968,In_734,In_2840);
nand U1969 (N_1969,In_1099,In_1551);
and U1970 (N_1970,In_2586,In_1036);
nand U1971 (N_1971,In_23,In_1160);
nor U1972 (N_1972,In_568,In_333);
nor U1973 (N_1973,In_2574,In_559);
nand U1974 (N_1974,In_2561,In_2679);
nor U1975 (N_1975,In_2873,In_769);
nor U1976 (N_1976,In_945,In_1134);
nand U1977 (N_1977,In_664,In_489);
nor U1978 (N_1978,In_951,In_583);
nor U1979 (N_1979,In_529,In_2507);
xor U1980 (N_1980,In_471,In_2326);
nand U1981 (N_1981,In_933,In_1239);
or U1982 (N_1982,In_140,In_1872);
xnor U1983 (N_1983,In_2086,In_295);
xor U1984 (N_1984,In_2826,In_1438);
nor U1985 (N_1985,In_752,In_677);
nor U1986 (N_1986,In_1069,In_1411);
nand U1987 (N_1987,In_1900,In_685);
or U1988 (N_1988,In_664,In_761);
or U1989 (N_1989,In_1637,In_1957);
and U1990 (N_1990,In_1094,In_2354);
and U1991 (N_1991,In_1425,In_108);
or U1992 (N_1992,In_684,In_2575);
and U1993 (N_1993,In_906,In_742);
nand U1994 (N_1994,In_2487,In_1253);
or U1995 (N_1995,In_2764,In_2337);
nor U1996 (N_1996,In_2901,In_1917);
nor U1997 (N_1997,In_2181,In_1190);
nor U1998 (N_1998,In_459,In_2429);
and U1999 (N_1999,In_1357,In_377);
nor U2000 (N_2000,In_598,In_2530);
nor U2001 (N_2001,In_507,In_2455);
xor U2002 (N_2002,In_1636,In_1420);
nor U2003 (N_2003,In_1894,In_1507);
nand U2004 (N_2004,In_1449,In_2428);
and U2005 (N_2005,In_297,In_264);
xnor U2006 (N_2006,In_2228,In_835);
nand U2007 (N_2007,In_2535,In_2720);
nand U2008 (N_2008,In_1057,In_2990);
nor U2009 (N_2009,In_2509,In_2096);
or U2010 (N_2010,In_1844,In_1769);
or U2011 (N_2011,In_2984,In_855);
or U2012 (N_2012,In_1261,In_1154);
or U2013 (N_2013,In_283,In_2008);
nor U2014 (N_2014,In_2360,In_829);
nand U2015 (N_2015,In_1733,In_2548);
nor U2016 (N_2016,In_21,In_2817);
nor U2017 (N_2017,In_1215,In_1684);
or U2018 (N_2018,In_504,In_2707);
nor U2019 (N_2019,In_433,In_760);
nor U2020 (N_2020,In_1051,In_2688);
nand U2021 (N_2021,In_1141,In_1957);
nor U2022 (N_2022,In_2377,In_1438);
nor U2023 (N_2023,In_1318,In_1898);
and U2024 (N_2024,In_1579,In_1879);
xor U2025 (N_2025,In_25,In_238);
nand U2026 (N_2026,In_867,In_2411);
xnor U2027 (N_2027,In_1252,In_166);
and U2028 (N_2028,In_541,In_2342);
nor U2029 (N_2029,In_2738,In_749);
nand U2030 (N_2030,In_2855,In_2327);
xor U2031 (N_2031,In_2291,In_949);
nand U2032 (N_2032,In_2280,In_2143);
xnor U2033 (N_2033,In_277,In_1296);
xnor U2034 (N_2034,In_1601,In_793);
nor U2035 (N_2035,In_2601,In_666);
nor U2036 (N_2036,In_797,In_1048);
xnor U2037 (N_2037,In_654,In_1329);
or U2038 (N_2038,In_2150,In_1888);
nor U2039 (N_2039,In_1434,In_1034);
or U2040 (N_2040,In_284,In_957);
xnor U2041 (N_2041,In_1861,In_21);
and U2042 (N_2042,In_1336,In_2942);
and U2043 (N_2043,In_241,In_1264);
xnor U2044 (N_2044,In_2459,In_558);
or U2045 (N_2045,In_1287,In_112);
nor U2046 (N_2046,In_1143,In_2225);
xor U2047 (N_2047,In_1483,In_228);
xor U2048 (N_2048,In_985,In_2747);
and U2049 (N_2049,In_1467,In_604);
nor U2050 (N_2050,In_681,In_2752);
xnor U2051 (N_2051,In_2594,In_966);
xnor U2052 (N_2052,In_2064,In_2031);
or U2053 (N_2053,In_1956,In_947);
nor U2054 (N_2054,In_1003,In_1875);
xnor U2055 (N_2055,In_2184,In_653);
or U2056 (N_2056,In_2968,In_1209);
xor U2057 (N_2057,In_561,In_1914);
nand U2058 (N_2058,In_320,In_506);
and U2059 (N_2059,In_1070,In_2313);
nor U2060 (N_2060,In_1125,In_1155);
nand U2061 (N_2061,In_95,In_1382);
or U2062 (N_2062,In_1392,In_1769);
xnor U2063 (N_2063,In_2969,In_2318);
xnor U2064 (N_2064,In_2047,In_2432);
nand U2065 (N_2065,In_486,In_1783);
or U2066 (N_2066,In_1344,In_269);
and U2067 (N_2067,In_135,In_1285);
nand U2068 (N_2068,In_938,In_1569);
xor U2069 (N_2069,In_319,In_2697);
and U2070 (N_2070,In_2074,In_627);
nor U2071 (N_2071,In_2528,In_2211);
xnor U2072 (N_2072,In_630,In_946);
xnor U2073 (N_2073,In_1558,In_2609);
and U2074 (N_2074,In_2458,In_887);
and U2075 (N_2075,In_1545,In_2807);
or U2076 (N_2076,In_1573,In_2778);
nand U2077 (N_2077,In_1039,In_108);
and U2078 (N_2078,In_626,In_1249);
and U2079 (N_2079,In_669,In_1024);
xnor U2080 (N_2080,In_937,In_2574);
xnor U2081 (N_2081,In_2412,In_991);
or U2082 (N_2082,In_252,In_2493);
and U2083 (N_2083,In_872,In_2617);
nand U2084 (N_2084,In_2993,In_480);
nor U2085 (N_2085,In_968,In_1947);
and U2086 (N_2086,In_1295,In_91);
or U2087 (N_2087,In_1116,In_965);
nor U2088 (N_2088,In_1038,In_2270);
nor U2089 (N_2089,In_1796,In_1391);
nor U2090 (N_2090,In_2140,In_2275);
or U2091 (N_2091,In_308,In_2217);
nand U2092 (N_2092,In_2418,In_276);
or U2093 (N_2093,In_2194,In_2331);
or U2094 (N_2094,In_1223,In_1784);
and U2095 (N_2095,In_627,In_214);
nor U2096 (N_2096,In_1292,In_769);
xor U2097 (N_2097,In_2918,In_524);
nand U2098 (N_2098,In_1247,In_2636);
nand U2099 (N_2099,In_2441,In_1810);
nor U2100 (N_2100,In_2567,In_1976);
and U2101 (N_2101,In_2022,In_2053);
xor U2102 (N_2102,In_475,In_2714);
or U2103 (N_2103,In_2165,In_843);
and U2104 (N_2104,In_1730,In_1115);
and U2105 (N_2105,In_924,In_1152);
or U2106 (N_2106,In_1068,In_2409);
nor U2107 (N_2107,In_335,In_1077);
xnor U2108 (N_2108,In_564,In_2825);
nor U2109 (N_2109,In_2461,In_1273);
nand U2110 (N_2110,In_397,In_2946);
and U2111 (N_2111,In_256,In_1642);
xor U2112 (N_2112,In_1329,In_694);
or U2113 (N_2113,In_1602,In_496);
nand U2114 (N_2114,In_1590,In_333);
xor U2115 (N_2115,In_915,In_2618);
nor U2116 (N_2116,In_457,In_780);
xnor U2117 (N_2117,In_1696,In_320);
and U2118 (N_2118,In_1526,In_456);
nor U2119 (N_2119,In_1683,In_2164);
and U2120 (N_2120,In_2724,In_928);
nand U2121 (N_2121,In_686,In_1005);
nor U2122 (N_2122,In_937,In_1823);
nand U2123 (N_2123,In_867,In_1328);
nand U2124 (N_2124,In_1966,In_1962);
nor U2125 (N_2125,In_2375,In_2131);
and U2126 (N_2126,In_1390,In_679);
nor U2127 (N_2127,In_723,In_2247);
xor U2128 (N_2128,In_85,In_458);
xnor U2129 (N_2129,In_2023,In_567);
or U2130 (N_2130,In_875,In_2176);
or U2131 (N_2131,In_1663,In_814);
and U2132 (N_2132,In_1731,In_380);
and U2133 (N_2133,In_71,In_1735);
nor U2134 (N_2134,In_874,In_202);
and U2135 (N_2135,In_1297,In_2039);
xnor U2136 (N_2136,In_1069,In_1793);
xnor U2137 (N_2137,In_1955,In_406);
nor U2138 (N_2138,In_1652,In_1483);
nor U2139 (N_2139,In_1094,In_2347);
or U2140 (N_2140,In_235,In_593);
nor U2141 (N_2141,In_1312,In_2698);
or U2142 (N_2142,In_166,In_1927);
nor U2143 (N_2143,In_2745,In_1448);
nand U2144 (N_2144,In_2833,In_904);
and U2145 (N_2145,In_2991,In_1462);
and U2146 (N_2146,In_2482,In_2484);
or U2147 (N_2147,In_2335,In_424);
and U2148 (N_2148,In_1319,In_899);
nand U2149 (N_2149,In_1917,In_815);
and U2150 (N_2150,In_2541,In_2882);
or U2151 (N_2151,In_2929,In_399);
and U2152 (N_2152,In_1251,In_2705);
xor U2153 (N_2153,In_1716,In_2486);
and U2154 (N_2154,In_2783,In_582);
xor U2155 (N_2155,In_2839,In_2258);
and U2156 (N_2156,In_513,In_1890);
nor U2157 (N_2157,In_1466,In_2051);
nand U2158 (N_2158,In_453,In_1758);
nand U2159 (N_2159,In_1812,In_1680);
and U2160 (N_2160,In_595,In_125);
nor U2161 (N_2161,In_2469,In_2114);
nor U2162 (N_2162,In_1728,In_2338);
nand U2163 (N_2163,In_1025,In_513);
or U2164 (N_2164,In_2643,In_561);
nor U2165 (N_2165,In_2608,In_308);
nand U2166 (N_2166,In_418,In_260);
xor U2167 (N_2167,In_711,In_2849);
nor U2168 (N_2168,In_1716,In_1951);
nor U2169 (N_2169,In_417,In_1769);
nand U2170 (N_2170,In_1778,In_1265);
xnor U2171 (N_2171,In_2220,In_2569);
and U2172 (N_2172,In_1443,In_2961);
and U2173 (N_2173,In_2736,In_682);
and U2174 (N_2174,In_501,In_2526);
xnor U2175 (N_2175,In_2823,In_905);
nand U2176 (N_2176,In_575,In_1696);
xnor U2177 (N_2177,In_2137,In_2835);
nor U2178 (N_2178,In_168,In_2815);
and U2179 (N_2179,In_2709,In_860);
or U2180 (N_2180,In_2624,In_1609);
nand U2181 (N_2181,In_1324,In_1910);
xnor U2182 (N_2182,In_943,In_2029);
nor U2183 (N_2183,In_2733,In_724);
and U2184 (N_2184,In_738,In_88);
xor U2185 (N_2185,In_2688,In_2505);
nand U2186 (N_2186,In_1899,In_435);
nor U2187 (N_2187,In_494,In_2511);
nor U2188 (N_2188,In_2589,In_2995);
nand U2189 (N_2189,In_2075,In_2694);
xor U2190 (N_2190,In_1693,In_1959);
nor U2191 (N_2191,In_2442,In_2868);
nor U2192 (N_2192,In_1236,In_2820);
and U2193 (N_2193,In_1360,In_202);
or U2194 (N_2194,In_1143,In_783);
and U2195 (N_2195,In_165,In_760);
and U2196 (N_2196,In_680,In_1860);
nand U2197 (N_2197,In_1851,In_815);
and U2198 (N_2198,In_2401,In_2640);
nand U2199 (N_2199,In_1321,In_1573);
or U2200 (N_2200,In_1392,In_981);
or U2201 (N_2201,In_1969,In_943);
xor U2202 (N_2202,In_278,In_1036);
nor U2203 (N_2203,In_597,In_2673);
or U2204 (N_2204,In_1722,In_1458);
xnor U2205 (N_2205,In_1065,In_2204);
and U2206 (N_2206,In_2559,In_1618);
nor U2207 (N_2207,In_2236,In_2073);
or U2208 (N_2208,In_1337,In_1358);
or U2209 (N_2209,In_1113,In_2982);
xnor U2210 (N_2210,In_403,In_2567);
nor U2211 (N_2211,In_2965,In_2689);
nand U2212 (N_2212,In_442,In_2786);
nor U2213 (N_2213,In_2664,In_893);
nand U2214 (N_2214,In_2478,In_264);
nor U2215 (N_2215,In_2300,In_2779);
and U2216 (N_2216,In_2274,In_909);
xnor U2217 (N_2217,In_2209,In_994);
nor U2218 (N_2218,In_296,In_2642);
and U2219 (N_2219,In_1823,In_1463);
xor U2220 (N_2220,In_1263,In_470);
nor U2221 (N_2221,In_367,In_966);
nand U2222 (N_2222,In_1183,In_515);
nor U2223 (N_2223,In_1125,In_628);
or U2224 (N_2224,In_417,In_2905);
or U2225 (N_2225,In_2891,In_2189);
or U2226 (N_2226,In_2032,In_1889);
nor U2227 (N_2227,In_983,In_1265);
nor U2228 (N_2228,In_1879,In_2407);
nand U2229 (N_2229,In_1456,In_1689);
and U2230 (N_2230,In_2493,In_1051);
xnor U2231 (N_2231,In_642,In_1202);
nand U2232 (N_2232,In_2736,In_1264);
xor U2233 (N_2233,In_714,In_1569);
nand U2234 (N_2234,In_155,In_2682);
and U2235 (N_2235,In_2013,In_2851);
and U2236 (N_2236,In_834,In_1145);
and U2237 (N_2237,In_119,In_2723);
xor U2238 (N_2238,In_2505,In_912);
nor U2239 (N_2239,In_708,In_2333);
nor U2240 (N_2240,In_2908,In_2773);
nand U2241 (N_2241,In_2858,In_302);
or U2242 (N_2242,In_470,In_2506);
nand U2243 (N_2243,In_444,In_2512);
xor U2244 (N_2244,In_2268,In_1098);
and U2245 (N_2245,In_2459,In_361);
xnor U2246 (N_2246,In_2750,In_1230);
and U2247 (N_2247,In_1057,In_1586);
xnor U2248 (N_2248,In_1144,In_725);
xor U2249 (N_2249,In_144,In_1954);
nor U2250 (N_2250,In_1681,In_1648);
xnor U2251 (N_2251,In_2628,In_243);
xnor U2252 (N_2252,In_1955,In_2906);
xnor U2253 (N_2253,In_179,In_2493);
nor U2254 (N_2254,In_244,In_420);
and U2255 (N_2255,In_829,In_1092);
xnor U2256 (N_2256,In_1649,In_0);
nand U2257 (N_2257,In_848,In_2654);
nand U2258 (N_2258,In_998,In_1186);
xnor U2259 (N_2259,In_351,In_757);
nand U2260 (N_2260,In_1661,In_1483);
xor U2261 (N_2261,In_1604,In_247);
xor U2262 (N_2262,In_1277,In_1701);
xnor U2263 (N_2263,In_2776,In_2645);
and U2264 (N_2264,In_427,In_1095);
nor U2265 (N_2265,In_366,In_332);
and U2266 (N_2266,In_519,In_2377);
or U2267 (N_2267,In_1284,In_1724);
or U2268 (N_2268,In_2395,In_2892);
nor U2269 (N_2269,In_920,In_964);
or U2270 (N_2270,In_128,In_2923);
nand U2271 (N_2271,In_465,In_1125);
nor U2272 (N_2272,In_1785,In_785);
nand U2273 (N_2273,In_482,In_397);
and U2274 (N_2274,In_543,In_1428);
and U2275 (N_2275,In_442,In_1844);
xnor U2276 (N_2276,In_2709,In_2014);
and U2277 (N_2277,In_2399,In_2762);
or U2278 (N_2278,In_2531,In_2446);
nor U2279 (N_2279,In_105,In_2854);
nor U2280 (N_2280,In_2433,In_540);
and U2281 (N_2281,In_554,In_747);
nor U2282 (N_2282,In_1601,In_717);
and U2283 (N_2283,In_1965,In_475);
or U2284 (N_2284,In_433,In_2564);
or U2285 (N_2285,In_15,In_315);
or U2286 (N_2286,In_1320,In_2044);
or U2287 (N_2287,In_2190,In_2426);
or U2288 (N_2288,In_539,In_1054);
and U2289 (N_2289,In_1780,In_2679);
nand U2290 (N_2290,In_1109,In_1707);
xor U2291 (N_2291,In_885,In_1739);
xnor U2292 (N_2292,In_1015,In_1011);
or U2293 (N_2293,In_1329,In_2673);
and U2294 (N_2294,In_436,In_2051);
or U2295 (N_2295,In_1071,In_1045);
nand U2296 (N_2296,In_1324,In_2451);
xor U2297 (N_2297,In_1135,In_2241);
nor U2298 (N_2298,In_2588,In_1117);
nand U2299 (N_2299,In_51,In_1984);
nand U2300 (N_2300,In_952,In_2918);
nor U2301 (N_2301,In_866,In_1945);
and U2302 (N_2302,In_968,In_2976);
nand U2303 (N_2303,In_822,In_2107);
and U2304 (N_2304,In_2572,In_600);
nand U2305 (N_2305,In_1270,In_2099);
or U2306 (N_2306,In_2557,In_97);
xor U2307 (N_2307,In_1201,In_462);
or U2308 (N_2308,In_1038,In_2313);
xor U2309 (N_2309,In_478,In_2632);
or U2310 (N_2310,In_1314,In_1253);
nor U2311 (N_2311,In_1345,In_2496);
nor U2312 (N_2312,In_2080,In_656);
xor U2313 (N_2313,In_1941,In_1235);
nand U2314 (N_2314,In_1642,In_219);
nand U2315 (N_2315,In_2915,In_1688);
nand U2316 (N_2316,In_2466,In_235);
nor U2317 (N_2317,In_2483,In_2273);
nor U2318 (N_2318,In_2951,In_348);
or U2319 (N_2319,In_2403,In_817);
nor U2320 (N_2320,In_987,In_1044);
and U2321 (N_2321,In_1931,In_447);
nand U2322 (N_2322,In_2063,In_1802);
nand U2323 (N_2323,In_2821,In_2591);
and U2324 (N_2324,In_2051,In_1976);
nor U2325 (N_2325,In_1950,In_82);
and U2326 (N_2326,In_1077,In_1110);
or U2327 (N_2327,In_905,In_1900);
and U2328 (N_2328,In_7,In_113);
xnor U2329 (N_2329,In_1242,In_494);
nor U2330 (N_2330,In_1754,In_2226);
and U2331 (N_2331,In_1802,In_684);
nor U2332 (N_2332,In_1283,In_2262);
xnor U2333 (N_2333,In_1711,In_357);
xor U2334 (N_2334,In_2077,In_1079);
or U2335 (N_2335,In_2000,In_2630);
nand U2336 (N_2336,In_1531,In_2930);
and U2337 (N_2337,In_2777,In_2896);
nor U2338 (N_2338,In_554,In_906);
and U2339 (N_2339,In_1692,In_1450);
and U2340 (N_2340,In_1903,In_1243);
and U2341 (N_2341,In_267,In_1374);
and U2342 (N_2342,In_2830,In_220);
nand U2343 (N_2343,In_588,In_2672);
and U2344 (N_2344,In_1938,In_2539);
xnor U2345 (N_2345,In_445,In_1045);
or U2346 (N_2346,In_2336,In_2653);
or U2347 (N_2347,In_1035,In_1551);
and U2348 (N_2348,In_1015,In_1328);
xor U2349 (N_2349,In_2224,In_1890);
xor U2350 (N_2350,In_2270,In_472);
nor U2351 (N_2351,In_1548,In_2191);
xnor U2352 (N_2352,In_1812,In_1106);
and U2353 (N_2353,In_2373,In_258);
or U2354 (N_2354,In_2715,In_489);
and U2355 (N_2355,In_136,In_2922);
and U2356 (N_2356,In_1018,In_2395);
and U2357 (N_2357,In_552,In_897);
xor U2358 (N_2358,In_1582,In_2868);
and U2359 (N_2359,In_2663,In_462);
nor U2360 (N_2360,In_2569,In_662);
xor U2361 (N_2361,In_2531,In_2136);
nand U2362 (N_2362,In_50,In_1596);
or U2363 (N_2363,In_1436,In_1634);
xnor U2364 (N_2364,In_448,In_932);
nand U2365 (N_2365,In_1586,In_1702);
nor U2366 (N_2366,In_1524,In_105);
or U2367 (N_2367,In_53,In_146);
or U2368 (N_2368,In_295,In_1530);
nand U2369 (N_2369,In_700,In_2589);
nand U2370 (N_2370,In_2262,In_1826);
and U2371 (N_2371,In_437,In_1663);
xnor U2372 (N_2372,In_1353,In_706);
and U2373 (N_2373,In_1826,In_1902);
or U2374 (N_2374,In_2459,In_2173);
xor U2375 (N_2375,In_2530,In_1133);
or U2376 (N_2376,In_744,In_1078);
or U2377 (N_2377,In_660,In_1980);
or U2378 (N_2378,In_2095,In_2966);
or U2379 (N_2379,In_1262,In_1343);
nand U2380 (N_2380,In_97,In_325);
or U2381 (N_2381,In_587,In_2939);
xor U2382 (N_2382,In_2972,In_1185);
nand U2383 (N_2383,In_2117,In_1671);
or U2384 (N_2384,In_2308,In_2259);
xor U2385 (N_2385,In_1532,In_727);
and U2386 (N_2386,In_2865,In_2316);
nor U2387 (N_2387,In_67,In_1420);
and U2388 (N_2388,In_1045,In_2283);
or U2389 (N_2389,In_1427,In_1315);
xor U2390 (N_2390,In_1916,In_2756);
and U2391 (N_2391,In_2255,In_2095);
nor U2392 (N_2392,In_1930,In_2483);
xnor U2393 (N_2393,In_1809,In_1551);
and U2394 (N_2394,In_2112,In_1291);
and U2395 (N_2395,In_181,In_2743);
xor U2396 (N_2396,In_582,In_2225);
xor U2397 (N_2397,In_2365,In_292);
or U2398 (N_2398,In_1589,In_92);
nor U2399 (N_2399,In_787,In_2211);
and U2400 (N_2400,In_2381,In_136);
nand U2401 (N_2401,In_367,In_2245);
and U2402 (N_2402,In_592,In_892);
or U2403 (N_2403,In_2498,In_82);
xnor U2404 (N_2404,In_2357,In_1270);
nor U2405 (N_2405,In_1638,In_2495);
nor U2406 (N_2406,In_762,In_2950);
nor U2407 (N_2407,In_1512,In_50);
xor U2408 (N_2408,In_2220,In_1443);
xnor U2409 (N_2409,In_2912,In_382);
and U2410 (N_2410,In_2428,In_281);
xor U2411 (N_2411,In_2863,In_1986);
nor U2412 (N_2412,In_948,In_328);
xor U2413 (N_2413,In_1062,In_266);
or U2414 (N_2414,In_2132,In_1483);
or U2415 (N_2415,In_2839,In_1321);
nor U2416 (N_2416,In_1504,In_1536);
nand U2417 (N_2417,In_890,In_1200);
nand U2418 (N_2418,In_1306,In_59);
or U2419 (N_2419,In_2065,In_117);
or U2420 (N_2420,In_1633,In_2059);
nand U2421 (N_2421,In_1381,In_177);
xor U2422 (N_2422,In_959,In_863);
or U2423 (N_2423,In_2912,In_218);
or U2424 (N_2424,In_248,In_36);
nand U2425 (N_2425,In_1465,In_555);
nand U2426 (N_2426,In_2095,In_2243);
and U2427 (N_2427,In_607,In_76);
nor U2428 (N_2428,In_1259,In_2154);
nor U2429 (N_2429,In_1060,In_1878);
and U2430 (N_2430,In_1176,In_88);
xor U2431 (N_2431,In_2553,In_594);
xor U2432 (N_2432,In_2511,In_2991);
and U2433 (N_2433,In_2621,In_1038);
nand U2434 (N_2434,In_1426,In_570);
nand U2435 (N_2435,In_2613,In_2410);
nand U2436 (N_2436,In_386,In_2012);
nand U2437 (N_2437,In_715,In_288);
and U2438 (N_2438,In_1723,In_786);
nor U2439 (N_2439,In_530,In_1138);
nand U2440 (N_2440,In_1711,In_1771);
or U2441 (N_2441,In_109,In_2163);
nand U2442 (N_2442,In_1207,In_1813);
and U2443 (N_2443,In_2401,In_370);
nand U2444 (N_2444,In_170,In_2494);
xnor U2445 (N_2445,In_1132,In_2966);
xor U2446 (N_2446,In_2656,In_2672);
xnor U2447 (N_2447,In_577,In_747);
nor U2448 (N_2448,In_1290,In_715);
nor U2449 (N_2449,In_1305,In_441);
or U2450 (N_2450,In_2806,In_2499);
xor U2451 (N_2451,In_1337,In_733);
and U2452 (N_2452,In_1939,In_1504);
nor U2453 (N_2453,In_1528,In_52);
nor U2454 (N_2454,In_1063,In_358);
xnor U2455 (N_2455,In_539,In_2632);
and U2456 (N_2456,In_2032,In_445);
nor U2457 (N_2457,In_1480,In_2359);
and U2458 (N_2458,In_2644,In_1189);
or U2459 (N_2459,In_2400,In_598);
and U2460 (N_2460,In_305,In_2160);
and U2461 (N_2461,In_294,In_1748);
xnor U2462 (N_2462,In_2502,In_2731);
nand U2463 (N_2463,In_2435,In_2732);
xnor U2464 (N_2464,In_1982,In_1957);
xor U2465 (N_2465,In_2107,In_1422);
nor U2466 (N_2466,In_1267,In_2562);
nor U2467 (N_2467,In_686,In_2285);
and U2468 (N_2468,In_2817,In_1459);
nor U2469 (N_2469,In_209,In_2830);
xnor U2470 (N_2470,In_1176,In_528);
nor U2471 (N_2471,In_2418,In_2682);
and U2472 (N_2472,In_1338,In_695);
nand U2473 (N_2473,In_2648,In_904);
or U2474 (N_2474,In_2359,In_1672);
nand U2475 (N_2475,In_941,In_1574);
xnor U2476 (N_2476,In_1961,In_2490);
or U2477 (N_2477,In_824,In_647);
nand U2478 (N_2478,In_1301,In_2289);
nor U2479 (N_2479,In_2145,In_1963);
xnor U2480 (N_2480,In_2939,In_1597);
nor U2481 (N_2481,In_2903,In_859);
nand U2482 (N_2482,In_2335,In_255);
xnor U2483 (N_2483,In_1946,In_1786);
or U2484 (N_2484,In_377,In_1467);
and U2485 (N_2485,In_1955,In_1529);
or U2486 (N_2486,In_2304,In_1267);
xor U2487 (N_2487,In_727,In_1724);
xnor U2488 (N_2488,In_104,In_1812);
or U2489 (N_2489,In_2163,In_1983);
or U2490 (N_2490,In_959,In_1064);
nand U2491 (N_2491,In_1518,In_390);
or U2492 (N_2492,In_1113,In_922);
xnor U2493 (N_2493,In_2564,In_1803);
nor U2494 (N_2494,In_80,In_1237);
and U2495 (N_2495,In_674,In_999);
nor U2496 (N_2496,In_2240,In_2805);
nand U2497 (N_2497,In_2620,In_1988);
or U2498 (N_2498,In_80,In_2848);
nor U2499 (N_2499,In_1161,In_385);
and U2500 (N_2500,In_2183,In_378);
nor U2501 (N_2501,In_2293,In_1992);
or U2502 (N_2502,In_2693,In_2533);
or U2503 (N_2503,In_123,In_2590);
or U2504 (N_2504,In_2837,In_1342);
nand U2505 (N_2505,In_1594,In_1502);
xor U2506 (N_2506,In_1307,In_518);
nor U2507 (N_2507,In_2940,In_1349);
nand U2508 (N_2508,In_1697,In_1103);
or U2509 (N_2509,In_373,In_245);
and U2510 (N_2510,In_120,In_2334);
or U2511 (N_2511,In_2789,In_275);
and U2512 (N_2512,In_965,In_1006);
and U2513 (N_2513,In_253,In_2808);
xor U2514 (N_2514,In_1708,In_1795);
nand U2515 (N_2515,In_526,In_2713);
nand U2516 (N_2516,In_930,In_1415);
and U2517 (N_2517,In_476,In_306);
nor U2518 (N_2518,In_1452,In_2970);
or U2519 (N_2519,In_2709,In_796);
xnor U2520 (N_2520,In_1533,In_1922);
or U2521 (N_2521,In_1213,In_1235);
and U2522 (N_2522,In_378,In_2741);
xor U2523 (N_2523,In_2118,In_2784);
xor U2524 (N_2524,In_2772,In_2353);
or U2525 (N_2525,In_646,In_1582);
or U2526 (N_2526,In_1297,In_854);
nor U2527 (N_2527,In_2646,In_2339);
and U2528 (N_2528,In_195,In_275);
and U2529 (N_2529,In_2295,In_882);
nand U2530 (N_2530,In_847,In_2426);
xnor U2531 (N_2531,In_748,In_273);
or U2532 (N_2532,In_1092,In_1499);
xor U2533 (N_2533,In_377,In_898);
and U2534 (N_2534,In_1104,In_1433);
or U2535 (N_2535,In_1995,In_1238);
or U2536 (N_2536,In_865,In_2095);
nor U2537 (N_2537,In_1712,In_2370);
nand U2538 (N_2538,In_2891,In_1532);
xor U2539 (N_2539,In_874,In_2481);
nand U2540 (N_2540,In_586,In_2467);
and U2541 (N_2541,In_2923,In_91);
nor U2542 (N_2542,In_386,In_923);
xor U2543 (N_2543,In_407,In_1215);
xnor U2544 (N_2544,In_1093,In_1661);
and U2545 (N_2545,In_735,In_2828);
nand U2546 (N_2546,In_751,In_833);
xor U2547 (N_2547,In_318,In_2122);
or U2548 (N_2548,In_190,In_176);
nor U2549 (N_2549,In_1473,In_1608);
nand U2550 (N_2550,In_1922,In_1459);
and U2551 (N_2551,In_1035,In_2442);
or U2552 (N_2552,In_996,In_1518);
nand U2553 (N_2553,In_1533,In_47);
and U2554 (N_2554,In_1682,In_1999);
nand U2555 (N_2555,In_2986,In_1941);
or U2556 (N_2556,In_443,In_841);
and U2557 (N_2557,In_2008,In_2343);
and U2558 (N_2558,In_2179,In_2708);
nand U2559 (N_2559,In_943,In_162);
and U2560 (N_2560,In_1031,In_353);
and U2561 (N_2561,In_699,In_1223);
and U2562 (N_2562,In_1767,In_2170);
nor U2563 (N_2563,In_43,In_689);
and U2564 (N_2564,In_2669,In_2264);
nand U2565 (N_2565,In_1484,In_2342);
xor U2566 (N_2566,In_1671,In_1084);
or U2567 (N_2567,In_1742,In_520);
nand U2568 (N_2568,In_448,In_2337);
and U2569 (N_2569,In_284,In_1212);
nand U2570 (N_2570,In_106,In_2885);
nand U2571 (N_2571,In_2874,In_1602);
nor U2572 (N_2572,In_852,In_2603);
xor U2573 (N_2573,In_661,In_1577);
and U2574 (N_2574,In_1069,In_47);
xor U2575 (N_2575,In_2994,In_598);
or U2576 (N_2576,In_2998,In_2819);
or U2577 (N_2577,In_1260,In_1640);
and U2578 (N_2578,In_1640,In_448);
or U2579 (N_2579,In_2817,In_1900);
nor U2580 (N_2580,In_2832,In_1103);
or U2581 (N_2581,In_1783,In_2435);
nor U2582 (N_2582,In_2986,In_1796);
nand U2583 (N_2583,In_2871,In_77);
and U2584 (N_2584,In_1074,In_912);
xor U2585 (N_2585,In_2335,In_665);
nor U2586 (N_2586,In_1321,In_1878);
and U2587 (N_2587,In_708,In_679);
and U2588 (N_2588,In_2830,In_1892);
xnor U2589 (N_2589,In_565,In_4);
xor U2590 (N_2590,In_1368,In_878);
nand U2591 (N_2591,In_2962,In_423);
or U2592 (N_2592,In_1490,In_2039);
xnor U2593 (N_2593,In_1983,In_1985);
nand U2594 (N_2594,In_1705,In_2106);
xor U2595 (N_2595,In_2344,In_2184);
xor U2596 (N_2596,In_2285,In_11);
and U2597 (N_2597,In_1715,In_2462);
or U2598 (N_2598,In_908,In_2322);
nand U2599 (N_2599,In_1467,In_2442);
and U2600 (N_2600,In_1278,In_1157);
or U2601 (N_2601,In_2455,In_466);
nand U2602 (N_2602,In_2546,In_204);
nor U2603 (N_2603,In_2121,In_2557);
or U2604 (N_2604,In_201,In_2838);
nor U2605 (N_2605,In_340,In_918);
and U2606 (N_2606,In_2599,In_918);
and U2607 (N_2607,In_43,In_234);
nand U2608 (N_2608,In_950,In_2614);
nand U2609 (N_2609,In_2434,In_285);
or U2610 (N_2610,In_536,In_506);
and U2611 (N_2611,In_598,In_2574);
nand U2612 (N_2612,In_687,In_624);
nor U2613 (N_2613,In_1499,In_900);
and U2614 (N_2614,In_2083,In_1917);
or U2615 (N_2615,In_665,In_2669);
and U2616 (N_2616,In_798,In_1000);
xor U2617 (N_2617,In_273,In_1365);
xor U2618 (N_2618,In_739,In_1731);
xnor U2619 (N_2619,In_1799,In_620);
and U2620 (N_2620,In_1003,In_2967);
xnor U2621 (N_2621,In_70,In_390);
or U2622 (N_2622,In_1869,In_1583);
or U2623 (N_2623,In_2586,In_1311);
nand U2624 (N_2624,In_894,In_2231);
nand U2625 (N_2625,In_645,In_2872);
nand U2626 (N_2626,In_174,In_2337);
xnor U2627 (N_2627,In_1597,In_984);
and U2628 (N_2628,In_1928,In_698);
nor U2629 (N_2629,In_1036,In_261);
nor U2630 (N_2630,In_1217,In_1140);
nand U2631 (N_2631,In_1366,In_448);
nor U2632 (N_2632,In_623,In_2692);
xor U2633 (N_2633,In_1834,In_1941);
and U2634 (N_2634,In_2871,In_223);
or U2635 (N_2635,In_131,In_1920);
and U2636 (N_2636,In_2525,In_52);
xor U2637 (N_2637,In_2310,In_1912);
or U2638 (N_2638,In_622,In_2816);
and U2639 (N_2639,In_2853,In_212);
nor U2640 (N_2640,In_165,In_243);
and U2641 (N_2641,In_2662,In_2303);
nor U2642 (N_2642,In_1030,In_2891);
and U2643 (N_2643,In_963,In_1986);
nand U2644 (N_2644,In_18,In_654);
and U2645 (N_2645,In_686,In_103);
xor U2646 (N_2646,In_2527,In_2695);
xor U2647 (N_2647,In_217,In_2742);
and U2648 (N_2648,In_2879,In_2609);
nand U2649 (N_2649,In_1724,In_2870);
xor U2650 (N_2650,In_868,In_1185);
and U2651 (N_2651,In_1318,In_2020);
nor U2652 (N_2652,In_2804,In_119);
nand U2653 (N_2653,In_801,In_2852);
nor U2654 (N_2654,In_1273,In_2081);
xnor U2655 (N_2655,In_2839,In_1151);
and U2656 (N_2656,In_1968,In_2682);
and U2657 (N_2657,In_23,In_1399);
or U2658 (N_2658,In_1101,In_382);
and U2659 (N_2659,In_645,In_2373);
nand U2660 (N_2660,In_754,In_1003);
and U2661 (N_2661,In_357,In_2231);
nor U2662 (N_2662,In_2384,In_53);
nor U2663 (N_2663,In_2466,In_897);
nand U2664 (N_2664,In_1107,In_2676);
nor U2665 (N_2665,In_2842,In_188);
or U2666 (N_2666,In_677,In_2745);
xnor U2667 (N_2667,In_1519,In_591);
nor U2668 (N_2668,In_1527,In_2056);
and U2669 (N_2669,In_1999,In_554);
and U2670 (N_2670,In_623,In_2629);
or U2671 (N_2671,In_2183,In_752);
or U2672 (N_2672,In_1245,In_1352);
nand U2673 (N_2673,In_1265,In_2545);
nand U2674 (N_2674,In_1081,In_658);
nand U2675 (N_2675,In_1581,In_966);
and U2676 (N_2676,In_2948,In_2231);
and U2677 (N_2677,In_969,In_2523);
nand U2678 (N_2678,In_2770,In_1102);
and U2679 (N_2679,In_1545,In_2578);
and U2680 (N_2680,In_1641,In_2751);
nor U2681 (N_2681,In_1205,In_1973);
xor U2682 (N_2682,In_1460,In_1096);
and U2683 (N_2683,In_1507,In_2376);
and U2684 (N_2684,In_1982,In_829);
nand U2685 (N_2685,In_163,In_44);
xor U2686 (N_2686,In_2749,In_142);
xor U2687 (N_2687,In_2276,In_1102);
or U2688 (N_2688,In_227,In_1839);
nand U2689 (N_2689,In_2118,In_530);
nand U2690 (N_2690,In_2632,In_879);
and U2691 (N_2691,In_842,In_338);
nand U2692 (N_2692,In_75,In_1502);
xor U2693 (N_2693,In_516,In_1063);
and U2694 (N_2694,In_2931,In_2802);
nor U2695 (N_2695,In_2143,In_1381);
and U2696 (N_2696,In_1918,In_62);
and U2697 (N_2697,In_2202,In_2864);
and U2698 (N_2698,In_183,In_2514);
and U2699 (N_2699,In_2700,In_507);
nand U2700 (N_2700,In_2068,In_963);
nand U2701 (N_2701,In_1892,In_1101);
nor U2702 (N_2702,In_1218,In_2309);
or U2703 (N_2703,In_2289,In_680);
and U2704 (N_2704,In_2284,In_2624);
and U2705 (N_2705,In_2194,In_659);
or U2706 (N_2706,In_2997,In_918);
or U2707 (N_2707,In_2439,In_676);
nand U2708 (N_2708,In_1861,In_1358);
nor U2709 (N_2709,In_240,In_2744);
xnor U2710 (N_2710,In_1130,In_2228);
and U2711 (N_2711,In_1650,In_528);
and U2712 (N_2712,In_443,In_1901);
nor U2713 (N_2713,In_1121,In_802);
or U2714 (N_2714,In_368,In_2115);
nor U2715 (N_2715,In_2014,In_1983);
nor U2716 (N_2716,In_1588,In_1380);
xnor U2717 (N_2717,In_1830,In_915);
nor U2718 (N_2718,In_1749,In_1699);
nand U2719 (N_2719,In_645,In_201);
and U2720 (N_2720,In_2757,In_1266);
nand U2721 (N_2721,In_1355,In_1477);
xor U2722 (N_2722,In_2518,In_735);
and U2723 (N_2723,In_1629,In_2090);
xor U2724 (N_2724,In_1910,In_197);
nand U2725 (N_2725,In_2820,In_115);
nor U2726 (N_2726,In_2374,In_1594);
xor U2727 (N_2727,In_1678,In_36);
nor U2728 (N_2728,In_2712,In_705);
nand U2729 (N_2729,In_2672,In_1383);
and U2730 (N_2730,In_459,In_741);
nor U2731 (N_2731,In_1862,In_1102);
nand U2732 (N_2732,In_1446,In_2759);
nand U2733 (N_2733,In_33,In_957);
or U2734 (N_2734,In_1841,In_247);
nand U2735 (N_2735,In_2989,In_463);
nand U2736 (N_2736,In_1845,In_1878);
nor U2737 (N_2737,In_2737,In_2693);
and U2738 (N_2738,In_1627,In_2299);
nor U2739 (N_2739,In_1427,In_2418);
or U2740 (N_2740,In_1560,In_1393);
or U2741 (N_2741,In_757,In_1864);
nand U2742 (N_2742,In_1918,In_2078);
xor U2743 (N_2743,In_2452,In_11);
nor U2744 (N_2744,In_387,In_1419);
xor U2745 (N_2745,In_482,In_1736);
or U2746 (N_2746,In_626,In_2341);
or U2747 (N_2747,In_2859,In_968);
and U2748 (N_2748,In_2052,In_1270);
or U2749 (N_2749,In_2502,In_1764);
or U2750 (N_2750,In_2414,In_1933);
nand U2751 (N_2751,In_2123,In_2292);
or U2752 (N_2752,In_2969,In_2045);
and U2753 (N_2753,In_1662,In_442);
and U2754 (N_2754,In_936,In_1019);
and U2755 (N_2755,In_1737,In_460);
or U2756 (N_2756,In_1340,In_645);
or U2757 (N_2757,In_1340,In_431);
nand U2758 (N_2758,In_2970,In_2004);
nor U2759 (N_2759,In_457,In_2620);
or U2760 (N_2760,In_815,In_1112);
and U2761 (N_2761,In_1291,In_2591);
nor U2762 (N_2762,In_885,In_2621);
nor U2763 (N_2763,In_2580,In_888);
and U2764 (N_2764,In_1363,In_2449);
or U2765 (N_2765,In_2070,In_422);
and U2766 (N_2766,In_1127,In_2279);
nand U2767 (N_2767,In_2209,In_1960);
xor U2768 (N_2768,In_545,In_277);
or U2769 (N_2769,In_2710,In_2093);
nand U2770 (N_2770,In_400,In_883);
or U2771 (N_2771,In_811,In_1195);
nand U2772 (N_2772,In_1492,In_881);
nor U2773 (N_2773,In_465,In_850);
nand U2774 (N_2774,In_900,In_1723);
nand U2775 (N_2775,In_1090,In_2785);
nand U2776 (N_2776,In_1977,In_317);
nor U2777 (N_2777,In_1544,In_1478);
and U2778 (N_2778,In_298,In_853);
and U2779 (N_2779,In_2384,In_976);
nand U2780 (N_2780,In_757,In_1540);
nor U2781 (N_2781,In_1961,In_217);
nor U2782 (N_2782,In_1861,In_218);
and U2783 (N_2783,In_1753,In_1010);
nor U2784 (N_2784,In_1023,In_2046);
or U2785 (N_2785,In_2510,In_1888);
xor U2786 (N_2786,In_2668,In_342);
and U2787 (N_2787,In_301,In_2343);
xnor U2788 (N_2788,In_2721,In_2123);
and U2789 (N_2789,In_1839,In_1449);
or U2790 (N_2790,In_582,In_19);
or U2791 (N_2791,In_2309,In_2096);
and U2792 (N_2792,In_2748,In_2281);
nand U2793 (N_2793,In_518,In_1717);
and U2794 (N_2794,In_939,In_2807);
xor U2795 (N_2795,In_2231,In_354);
nor U2796 (N_2796,In_1613,In_1412);
nor U2797 (N_2797,In_635,In_154);
and U2798 (N_2798,In_1225,In_649);
xor U2799 (N_2799,In_681,In_2045);
and U2800 (N_2800,In_2802,In_2666);
nor U2801 (N_2801,In_360,In_2021);
and U2802 (N_2802,In_528,In_1177);
nand U2803 (N_2803,In_2607,In_2370);
nand U2804 (N_2804,In_2819,In_660);
xnor U2805 (N_2805,In_745,In_2687);
or U2806 (N_2806,In_2523,In_1169);
nand U2807 (N_2807,In_1720,In_1070);
nand U2808 (N_2808,In_2373,In_23);
nor U2809 (N_2809,In_1971,In_2814);
nand U2810 (N_2810,In_43,In_2948);
nor U2811 (N_2811,In_2160,In_2563);
nand U2812 (N_2812,In_288,In_965);
or U2813 (N_2813,In_1503,In_1441);
xor U2814 (N_2814,In_2561,In_2213);
and U2815 (N_2815,In_2050,In_1439);
nor U2816 (N_2816,In_1544,In_2509);
or U2817 (N_2817,In_781,In_1291);
and U2818 (N_2818,In_2093,In_69);
nand U2819 (N_2819,In_2121,In_2567);
and U2820 (N_2820,In_1654,In_1568);
xor U2821 (N_2821,In_397,In_548);
nand U2822 (N_2822,In_2108,In_974);
or U2823 (N_2823,In_2592,In_2442);
nand U2824 (N_2824,In_2829,In_2125);
nor U2825 (N_2825,In_2286,In_75);
or U2826 (N_2826,In_2598,In_1876);
xnor U2827 (N_2827,In_2556,In_2472);
nor U2828 (N_2828,In_2877,In_1946);
and U2829 (N_2829,In_1006,In_8);
xor U2830 (N_2830,In_2843,In_916);
or U2831 (N_2831,In_2512,In_1420);
and U2832 (N_2832,In_1740,In_2000);
nand U2833 (N_2833,In_1630,In_1669);
nand U2834 (N_2834,In_477,In_1712);
nand U2835 (N_2835,In_1330,In_2465);
xor U2836 (N_2836,In_630,In_1884);
or U2837 (N_2837,In_2349,In_678);
nor U2838 (N_2838,In_2640,In_1072);
nor U2839 (N_2839,In_2949,In_2527);
nand U2840 (N_2840,In_1583,In_2105);
nor U2841 (N_2841,In_1706,In_1065);
xor U2842 (N_2842,In_303,In_82);
or U2843 (N_2843,In_2843,In_628);
nor U2844 (N_2844,In_2129,In_1113);
nand U2845 (N_2845,In_2683,In_2896);
and U2846 (N_2846,In_1933,In_1102);
and U2847 (N_2847,In_1918,In_2515);
nor U2848 (N_2848,In_326,In_661);
xor U2849 (N_2849,In_2831,In_865);
or U2850 (N_2850,In_2519,In_89);
or U2851 (N_2851,In_2010,In_2441);
or U2852 (N_2852,In_649,In_1838);
xor U2853 (N_2853,In_2749,In_2616);
and U2854 (N_2854,In_1436,In_1675);
nor U2855 (N_2855,In_1974,In_2973);
nand U2856 (N_2856,In_2138,In_678);
or U2857 (N_2857,In_2836,In_1483);
and U2858 (N_2858,In_2653,In_931);
xor U2859 (N_2859,In_1083,In_380);
and U2860 (N_2860,In_1276,In_1037);
or U2861 (N_2861,In_2509,In_930);
nand U2862 (N_2862,In_1304,In_1482);
xor U2863 (N_2863,In_2045,In_1060);
nor U2864 (N_2864,In_2548,In_2381);
xnor U2865 (N_2865,In_440,In_1959);
xor U2866 (N_2866,In_1139,In_847);
xor U2867 (N_2867,In_2344,In_210);
nor U2868 (N_2868,In_1541,In_996);
nor U2869 (N_2869,In_1297,In_1577);
xnor U2870 (N_2870,In_2721,In_1912);
nand U2871 (N_2871,In_1375,In_2658);
nand U2872 (N_2872,In_1280,In_980);
xnor U2873 (N_2873,In_1415,In_428);
xnor U2874 (N_2874,In_806,In_49);
or U2875 (N_2875,In_988,In_730);
nand U2876 (N_2876,In_396,In_1653);
or U2877 (N_2877,In_1244,In_2994);
or U2878 (N_2878,In_592,In_2402);
nand U2879 (N_2879,In_745,In_1127);
nand U2880 (N_2880,In_2963,In_2172);
and U2881 (N_2881,In_594,In_291);
xnor U2882 (N_2882,In_2079,In_2552);
or U2883 (N_2883,In_290,In_2682);
or U2884 (N_2884,In_2671,In_680);
nor U2885 (N_2885,In_2838,In_1743);
nor U2886 (N_2886,In_451,In_1320);
nor U2887 (N_2887,In_2119,In_1297);
nor U2888 (N_2888,In_1328,In_1209);
and U2889 (N_2889,In_1999,In_1310);
or U2890 (N_2890,In_1094,In_415);
xor U2891 (N_2891,In_2086,In_1307);
xor U2892 (N_2892,In_1831,In_1685);
or U2893 (N_2893,In_874,In_2776);
nor U2894 (N_2894,In_597,In_686);
xnor U2895 (N_2895,In_2765,In_542);
nand U2896 (N_2896,In_509,In_1861);
nand U2897 (N_2897,In_2125,In_2461);
xor U2898 (N_2898,In_808,In_2413);
nor U2899 (N_2899,In_1920,In_1344);
or U2900 (N_2900,In_1939,In_1371);
nand U2901 (N_2901,In_2578,In_917);
or U2902 (N_2902,In_2035,In_1253);
nand U2903 (N_2903,In_2986,In_2887);
xnor U2904 (N_2904,In_1323,In_1451);
xor U2905 (N_2905,In_461,In_423);
and U2906 (N_2906,In_157,In_1823);
and U2907 (N_2907,In_398,In_2534);
xor U2908 (N_2908,In_1881,In_1092);
nand U2909 (N_2909,In_167,In_2443);
or U2910 (N_2910,In_135,In_2103);
xnor U2911 (N_2911,In_585,In_1216);
nand U2912 (N_2912,In_2018,In_2023);
or U2913 (N_2913,In_2422,In_820);
nand U2914 (N_2914,In_1617,In_1784);
xnor U2915 (N_2915,In_2312,In_807);
or U2916 (N_2916,In_2504,In_2094);
xor U2917 (N_2917,In_919,In_2813);
and U2918 (N_2918,In_0,In_2388);
and U2919 (N_2919,In_1537,In_668);
or U2920 (N_2920,In_1340,In_2988);
nand U2921 (N_2921,In_1089,In_2818);
and U2922 (N_2922,In_738,In_205);
xnor U2923 (N_2923,In_2515,In_2807);
nor U2924 (N_2924,In_1253,In_1648);
xor U2925 (N_2925,In_738,In_775);
xnor U2926 (N_2926,In_219,In_189);
nand U2927 (N_2927,In_247,In_2186);
nor U2928 (N_2928,In_1103,In_1096);
nand U2929 (N_2929,In_2727,In_996);
nor U2930 (N_2930,In_2903,In_2556);
or U2931 (N_2931,In_1667,In_2449);
nand U2932 (N_2932,In_2382,In_2475);
nand U2933 (N_2933,In_156,In_2943);
xnor U2934 (N_2934,In_2958,In_958);
or U2935 (N_2935,In_1269,In_2355);
and U2936 (N_2936,In_987,In_1756);
and U2937 (N_2937,In_1465,In_2474);
or U2938 (N_2938,In_20,In_2804);
or U2939 (N_2939,In_2703,In_2290);
and U2940 (N_2940,In_811,In_79);
and U2941 (N_2941,In_2616,In_298);
nand U2942 (N_2942,In_2883,In_2705);
xnor U2943 (N_2943,In_940,In_17);
nor U2944 (N_2944,In_1461,In_2730);
nor U2945 (N_2945,In_1647,In_967);
nand U2946 (N_2946,In_680,In_2335);
nor U2947 (N_2947,In_810,In_2423);
nor U2948 (N_2948,In_1059,In_1378);
nor U2949 (N_2949,In_1623,In_1871);
and U2950 (N_2950,In_1523,In_1882);
nor U2951 (N_2951,In_2795,In_384);
nor U2952 (N_2952,In_2551,In_1245);
nand U2953 (N_2953,In_2051,In_1574);
nand U2954 (N_2954,In_771,In_879);
nand U2955 (N_2955,In_1449,In_300);
xnor U2956 (N_2956,In_2771,In_1254);
and U2957 (N_2957,In_2869,In_476);
or U2958 (N_2958,In_46,In_743);
nor U2959 (N_2959,In_2487,In_831);
or U2960 (N_2960,In_2757,In_1382);
or U2961 (N_2961,In_2453,In_2576);
or U2962 (N_2962,In_31,In_316);
and U2963 (N_2963,In_1787,In_1386);
nand U2964 (N_2964,In_1949,In_1237);
or U2965 (N_2965,In_2454,In_522);
nand U2966 (N_2966,In_884,In_2202);
or U2967 (N_2967,In_2083,In_39);
nand U2968 (N_2968,In_1907,In_2725);
and U2969 (N_2969,In_481,In_1261);
or U2970 (N_2970,In_21,In_333);
nand U2971 (N_2971,In_2028,In_1682);
or U2972 (N_2972,In_581,In_2522);
xnor U2973 (N_2973,In_572,In_624);
and U2974 (N_2974,In_2100,In_1059);
xor U2975 (N_2975,In_1054,In_1664);
nand U2976 (N_2976,In_2595,In_982);
nand U2977 (N_2977,In_2890,In_585);
xor U2978 (N_2978,In_1181,In_365);
xor U2979 (N_2979,In_1965,In_633);
or U2980 (N_2980,In_1007,In_1106);
and U2981 (N_2981,In_1222,In_2211);
xor U2982 (N_2982,In_2271,In_1376);
nand U2983 (N_2983,In_2683,In_2425);
and U2984 (N_2984,In_965,In_1282);
and U2985 (N_2985,In_404,In_2553);
and U2986 (N_2986,In_968,In_1804);
xnor U2987 (N_2987,In_150,In_1327);
nor U2988 (N_2988,In_1488,In_2374);
or U2989 (N_2989,In_2682,In_2869);
xor U2990 (N_2990,In_2335,In_682);
xnor U2991 (N_2991,In_1650,In_179);
nand U2992 (N_2992,In_2362,In_230);
and U2993 (N_2993,In_1119,In_2299);
nor U2994 (N_2994,In_340,In_2701);
xnor U2995 (N_2995,In_2608,In_122);
nor U2996 (N_2996,In_2519,In_1713);
and U2997 (N_2997,In_209,In_2304);
or U2998 (N_2998,In_232,In_751);
nand U2999 (N_2999,In_335,In_814);
and U3000 (N_3000,N_961,N_271);
nor U3001 (N_3001,N_2911,N_597);
nand U3002 (N_3002,N_149,N_377);
nor U3003 (N_3003,N_53,N_669);
xnor U3004 (N_3004,N_978,N_2521);
and U3005 (N_3005,N_902,N_2003);
and U3006 (N_3006,N_2691,N_1769);
nor U3007 (N_3007,N_1990,N_550);
nand U3008 (N_3008,N_3,N_2327);
nor U3009 (N_3009,N_60,N_716);
or U3010 (N_3010,N_1106,N_952);
nand U3011 (N_3011,N_2436,N_1784);
xor U3012 (N_3012,N_861,N_1817);
or U3013 (N_3013,N_1068,N_1157);
or U3014 (N_3014,N_2405,N_1995);
or U3015 (N_3015,N_705,N_1028);
xor U3016 (N_3016,N_1668,N_2996);
and U3017 (N_3017,N_521,N_228);
or U3018 (N_3018,N_695,N_2273);
xor U3019 (N_3019,N_427,N_2696);
nor U3020 (N_3020,N_549,N_1021);
or U3021 (N_3021,N_1249,N_2675);
xnor U3022 (N_3022,N_691,N_1334);
nand U3023 (N_3023,N_1502,N_912);
nor U3024 (N_3024,N_706,N_1416);
xnor U3025 (N_3025,N_1494,N_816);
and U3026 (N_3026,N_115,N_268);
nor U3027 (N_3027,N_1159,N_433);
and U3028 (N_3028,N_100,N_163);
or U3029 (N_3029,N_2444,N_402);
nor U3030 (N_3030,N_2517,N_261);
and U3031 (N_3031,N_2113,N_958);
nand U3032 (N_3032,N_1713,N_857);
xnor U3033 (N_3033,N_1798,N_1103);
nor U3034 (N_3034,N_1257,N_1577);
nor U3035 (N_3035,N_910,N_1179);
xnor U3036 (N_3036,N_353,N_2950);
nand U3037 (N_3037,N_859,N_131);
nand U3038 (N_3038,N_47,N_890);
nor U3039 (N_3039,N_1617,N_2751);
and U3040 (N_3040,N_2447,N_293);
or U3041 (N_3041,N_394,N_317);
xor U3042 (N_3042,N_193,N_2154);
nor U3043 (N_3043,N_2046,N_1481);
or U3044 (N_3044,N_1055,N_309);
xnor U3045 (N_3045,N_1391,N_2101);
nor U3046 (N_3046,N_2352,N_2432);
nand U3047 (N_3047,N_1174,N_2940);
or U3048 (N_3048,N_230,N_791);
nand U3049 (N_3049,N_324,N_2822);
nor U3050 (N_3050,N_1581,N_1210);
or U3051 (N_3051,N_365,N_1946);
nand U3052 (N_3052,N_1357,N_238);
nand U3053 (N_3053,N_2491,N_2093);
xnor U3054 (N_3054,N_251,N_658);
and U3055 (N_3055,N_1310,N_2644);
nor U3056 (N_3056,N_959,N_1892);
xnor U3057 (N_3057,N_2633,N_165);
nand U3058 (N_3058,N_465,N_332);
or U3059 (N_3059,N_1402,N_2485);
nand U3060 (N_3060,N_2642,N_345);
or U3061 (N_3061,N_1065,N_2133);
nand U3062 (N_3062,N_130,N_2587);
xnor U3063 (N_3063,N_2823,N_1992);
nor U3064 (N_3064,N_1187,N_1156);
or U3065 (N_3065,N_1533,N_1653);
nor U3066 (N_3066,N_2657,N_1183);
nor U3067 (N_3067,N_2858,N_1927);
nand U3068 (N_3068,N_322,N_1666);
nor U3069 (N_3069,N_1478,N_1604);
or U3070 (N_3070,N_1690,N_2064);
nor U3071 (N_3071,N_141,N_2178);
nand U3072 (N_3072,N_1501,N_2254);
xor U3073 (N_3073,N_828,N_1611);
or U3074 (N_3074,N_1619,N_2719);
or U3075 (N_3075,N_2208,N_1601);
and U3076 (N_3076,N_35,N_2130);
xor U3077 (N_3077,N_1925,N_1823);
nand U3078 (N_3078,N_1796,N_2762);
nor U3079 (N_3079,N_1462,N_2140);
or U3080 (N_3080,N_1936,N_1412);
and U3081 (N_3081,N_1994,N_2588);
nand U3082 (N_3082,N_2532,N_1772);
or U3083 (N_3083,N_2928,N_1909);
xnor U3084 (N_3084,N_1410,N_583);
or U3085 (N_3085,N_1589,N_2699);
and U3086 (N_3086,N_2129,N_1050);
or U3087 (N_3087,N_1813,N_1913);
or U3088 (N_3088,N_657,N_2209);
or U3089 (N_3089,N_1506,N_506);
nor U3090 (N_3090,N_2877,N_1778);
nand U3091 (N_3091,N_2744,N_540);
nand U3092 (N_3092,N_2780,N_2802);
nor U3093 (N_3093,N_1976,N_75);
or U3094 (N_3094,N_187,N_2036);
and U3095 (N_3095,N_43,N_2157);
xor U3096 (N_3096,N_2037,N_652);
nor U3097 (N_3097,N_2071,N_2278);
nor U3098 (N_3098,N_2776,N_2362);
xor U3099 (N_3099,N_288,N_1133);
xnor U3100 (N_3100,N_1023,N_1192);
or U3101 (N_3101,N_2285,N_2593);
xor U3102 (N_3102,N_1010,N_932);
nor U3103 (N_3103,N_325,N_605);
nor U3104 (N_3104,N_2239,N_2302);
and U3105 (N_3105,N_477,N_869);
xor U3106 (N_3106,N_2164,N_2769);
nor U3107 (N_3107,N_2002,N_1258);
xnor U3108 (N_3108,N_320,N_2553);
nor U3109 (N_3109,N_2516,N_2537);
nor U3110 (N_3110,N_779,N_2736);
nor U3111 (N_3111,N_1298,N_1836);
nor U3112 (N_3112,N_630,N_2793);
and U3113 (N_3113,N_732,N_782);
nand U3114 (N_3114,N_2812,N_1684);
nand U3115 (N_3115,N_1742,N_2323);
nor U3116 (N_3116,N_2507,N_2547);
nand U3117 (N_3117,N_2555,N_96);
or U3118 (N_3118,N_360,N_395);
nor U3119 (N_3119,N_2925,N_1180);
and U3120 (N_3120,N_397,N_2543);
or U3121 (N_3121,N_969,N_2032);
xor U3122 (N_3122,N_687,N_931);
xnor U3123 (N_3123,N_1614,N_425);
nor U3124 (N_3124,N_613,N_1255);
or U3125 (N_3125,N_1264,N_1962);
nor U3126 (N_3126,N_2333,N_1038);
nand U3127 (N_3127,N_2216,N_2722);
or U3128 (N_3128,N_1809,N_1736);
or U3129 (N_3129,N_2427,N_572);
nor U3130 (N_3130,N_1880,N_837);
and U3131 (N_3131,N_1514,N_254);
nor U3132 (N_3132,N_44,N_2042);
or U3133 (N_3133,N_1429,N_626);
nor U3134 (N_3134,N_849,N_2045);
nor U3135 (N_3135,N_528,N_1726);
xnor U3136 (N_3136,N_556,N_1094);
or U3137 (N_3137,N_2887,N_1779);
nor U3138 (N_3138,N_1718,N_432);
nor U3139 (N_3139,N_2471,N_2057);
nand U3140 (N_3140,N_1337,N_2685);
nor U3141 (N_3141,N_388,N_2550);
nand U3142 (N_3142,N_1590,N_945);
xor U3143 (N_3143,N_265,N_2635);
nand U3144 (N_3144,N_2372,N_410);
xnor U3145 (N_3145,N_984,N_1761);
xnor U3146 (N_3146,N_748,N_198);
and U3147 (N_3147,N_1168,N_1679);
or U3148 (N_3148,N_29,N_2929);
or U3149 (N_3149,N_666,N_1582);
nand U3150 (N_3150,N_1363,N_2712);
and U3151 (N_3151,N_2402,N_314);
xnor U3152 (N_3152,N_962,N_792);
xor U3153 (N_3153,N_1250,N_595);
nor U3154 (N_3154,N_2941,N_832);
nand U3155 (N_3155,N_2538,N_2167);
or U3156 (N_3156,N_2956,N_2321);
nor U3157 (N_3157,N_781,N_643);
and U3158 (N_3158,N_2655,N_1715);
nand U3159 (N_3159,N_2143,N_741);
nor U3160 (N_3160,N_2843,N_169);
nor U3161 (N_3161,N_1985,N_1007);
or U3162 (N_3162,N_2438,N_994);
or U3163 (N_3163,N_951,N_318);
xor U3164 (N_3164,N_1982,N_2827);
nor U3165 (N_3165,N_1491,N_2609);
and U3166 (N_3166,N_2185,N_560);
nor U3167 (N_3167,N_1943,N_2945);
nor U3168 (N_3168,N_1579,N_137);
or U3169 (N_3169,N_279,N_2369);
or U3170 (N_3170,N_1495,N_2189);
xnor U3171 (N_3171,N_2206,N_127);
or U3172 (N_3172,N_278,N_439);
or U3173 (N_3173,N_372,N_1868);
xnor U3174 (N_3174,N_111,N_1767);
xor U3175 (N_3175,N_2968,N_1522);
xnor U3176 (N_3176,N_1591,N_2639);
or U3177 (N_3177,N_1153,N_102);
and U3178 (N_3178,N_1548,N_97);
xnor U3179 (N_3179,N_2415,N_2999);
nand U3180 (N_3180,N_128,N_2374);
or U3181 (N_3181,N_1259,N_236);
and U3182 (N_3182,N_64,N_9);
nand U3183 (N_3183,N_686,N_1035);
nor U3184 (N_3184,N_2295,N_382);
xor U3185 (N_3185,N_2778,N_2282);
xor U3186 (N_3186,N_2456,N_1528);
nor U3187 (N_3187,N_2307,N_2612);
nand U3188 (N_3188,N_2431,N_510);
or U3189 (N_3189,N_775,N_2605);
or U3190 (N_3190,N_257,N_1236);
nor U3191 (N_3191,N_898,N_1170);
or U3192 (N_3192,N_2473,N_876);
or U3193 (N_3193,N_766,N_2775);
nand U3194 (N_3194,N_1562,N_2406);
or U3195 (N_3195,N_1015,N_589);
nand U3196 (N_3196,N_2747,N_2397);
and U3197 (N_3197,N_239,N_2294);
xor U3198 (N_3198,N_2418,N_2052);
and U3199 (N_3199,N_2370,N_2579);
xnor U3200 (N_3200,N_1698,N_724);
nand U3201 (N_3201,N_1573,N_2753);
and U3202 (N_3202,N_2081,N_1375);
or U3203 (N_3203,N_2790,N_408);
or U3204 (N_3204,N_466,N_1191);
nor U3205 (N_3205,N_2868,N_2669);
or U3206 (N_3206,N_168,N_462);
nor U3207 (N_3207,N_2810,N_1025);
and U3208 (N_3208,N_1887,N_500);
nor U3209 (N_3209,N_424,N_281);
nand U3210 (N_3210,N_2048,N_2331);
nand U3211 (N_3211,N_2760,N_569);
and U3212 (N_3212,N_1919,N_2451);
nor U3213 (N_3213,N_1006,N_1659);
and U3214 (N_3214,N_1359,N_1696);
nand U3215 (N_3215,N_303,N_1847);
and U3216 (N_3216,N_1876,N_2180);
or U3217 (N_3217,N_2009,N_2492);
or U3218 (N_3218,N_1320,N_1711);
nor U3219 (N_3219,N_1443,N_979);
and U3220 (N_3220,N_1871,N_1161);
nand U3221 (N_3221,N_2236,N_2872);
or U3222 (N_3222,N_443,N_78);
nor U3223 (N_3223,N_1881,N_1903);
nand U3224 (N_3224,N_2151,N_2342);
and U3225 (N_3225,N_2698,N_420);
and U3226 (N_3226,N_2661,N_2224);
or U3227 (N_3227,N_380,N_2572);
nand U3228 (N_3228,N_335,N_2092);
nor U3229 (N_3229,N_1929,N_2390);
xnor U3230 (N_3230,N_520,N_1801);
nand U3231 (N_3231,N_2155,N_206);
nor U3232 (N_3232,N_1643,N_1398);
nor U3233 (N_3233,N_161,N_2566);
nor U3234 (N_3234,N_2934,N_2256);
nand U3235 (N_3235,N_921,N_618);
xnor U3236 (N_3236,N_157,N_757);
nor U3237 (N_3237,N_457,N_177);
and U3238 (N_3238,N_374,N_923);
or U3239 (N_3239,N_2797,N_1444);
nor U3240 (N_3240,N_2548,N_1154);
or U3241 (N_3241,N_2924,N_545);
nand U3242 (N_3242,N_112,N_2690);
nand U3243 (N_3243,N_2643,N_216);
nor U3244 (N_3244,N_2275,N_1327);
nor U3245 (N_3245,N_1474,N_640);
nor U3246 (N_3246,N_1704,N_689);
xor U3247 (N_3247,N_1353,N_863);
and U3248 (N_3248,N_2580,N_1692);
xor U3249 (N_3249,N_1907,N_2560);
nor U3250 (N_3250,N_1189,N_1268);
nor U3251 (N_3251,N_488,N_1722);
and U3252 (N_3252,N_366,N_693);
or U3253 (N_3253,N_1143,N_999);
nand U3254 (N_3254,N_207,N_2463);
and U3255 (N_3255,N_2668,N_2920);
nand U3256 (N_3256,N_81,N_1200);
xor U3257 (N_3257,N_1596,N_2804);
nand U3258 (N_3258,N_787,N_2330);
xnor U3259 (N_3259,N_1012,N_31);
nand U3260 (N_3260,N_2735,N_1541);
nor U3261 (N_3261,N_1126,N_707);
or U3262 (N_3262,N_1821,N_1476);
and U3263 (N_3263,N_2611,N_179);
xor U3264 (N_3264,N_2198,N_373);
and U3265 (N_3265,N_134,N_1561);
nand U3266 (N_3266,N_2297,N_1140);
or U3267 (N_3267,N_2512,N_1669);
nand U3268 (N_3268,N_2475,N_1859);
and U3269 (N_3269,N_1656,N_296);
and U3270 (N_3270,N_761,N_644);
nand U3271 (N_3271,N_944,N_722);
xor U3272 (N_3272,N_2761,N_1063);
or U3273 (N_3273,N_480,N_1487);
and U3274 (N_3274,N_2030,N_2839);
nand U3275 (N_3275,N_52,N_610);
or U3276 (N_3276,N_2077,N_516);
and U3277 (N_3277,N_2146,N_449);
or U3278 (N_3278,N_525,N_2477);
nor U3279 (N_3279,N_284,N_2878);
nor U3280 (N_3280,N_1017,N_2708);
nand U3281 (N_3281,N_1266,N_20);
nor U3282 (N_3282,N_80,N_1875);
or U3283 (N_3283,N_1479,N_1745);
or U3284 (N_3284,N_2523,N_0);
nor U3285 (N_3285,N_1505,N_1751);
nand U3286 (N_3286,N_762,N_1229);
xor U3287 (N_3287,N_2375,N_1307);
nand U3288 (N_3288,N_1234,N_189);
or U3289 (N_3289,N_809,N_844);
or U3290 (N_3290,N_2862,N_2099);
xor U3291 (N_3291,N_246,N_2774);
and U3292 (N_3292,N_2695,N_412);
nand U3293 (N_3293,N_2479,N_1555);
nand U3294 (N_3294,N_1701,N_1922);
nor U3295 (N_3295,N_37,N_1734);
and U3296 (N_3296,N_1741,N_2047);
nand U3297 (N_3297,N_2671,N_270);
xnor U3298 (N_3298,N_1077,N_594);
xnor U3299 (N_3299,N_574,N_1246);
nor U3300 (N_3300,N_1475,N_1109);
and U3301 (N_3301,N_1630,N_2309);
and U3302 (N_3302,N_2453,N_2994);
xnor U3303 (N_3303,N_1197,N_585);
xor U3304 (N_3304,N_2808,N_248);
xnor U3305 (N_3305,N_2900,N_147);
or U3306 (N_3306,N_2384,N_1401);
nor U3307 (N_3307,N_865,N_2662);
and U3308 (N_3308,N_70,N_68);
nand U3309 (N_3309,N_767,N_1703);
or U3310 (N_3310,N_400,N_2090);
or U3311 (N_3311,N_1648,N_769);
xor U3312 (N_3312,N_609,N_153);
and U3313 (N_3313,N_2905,N_1584);
or U3314 (N_3314,N_411,N_838);
nand U3315 (N_3315,N_2087,N_328);
and U3316 (N_3316,N_2651,N_1660);
or U3317 (N_3317,N_1981,N_2065);
xnor U3318 (N_3318,N_2656,N_1790);
nand U3319 (N_3319,N_1697,N_6);
nor U3320 (N_3320,N_641,N_843);
and U3321 (N_3321,N_1276,N_1305);
nor U3322 (N_3322,N_13,N_1542);
xnor U3323 (N_3323,N_2345,N_1647);
xor U3324 (N_3324,N_2739,N_1317);
or U3325 (N_3325,N_2450,N_1111);
nor U3326 (N_3326,N_708,N_874);
and U3327 (N_3327,N_2970,N_2325);
and U3328 (N_3328,N_1289,N_2788);
and U3329 (N_3329,N_2422,N_2335);
xnor U3330 (N_3330,N_34,N_2184);
or U3331 (N_3331,N_2589,N_2715);
xor U3332 (N_3332,N_1001,N_329);
nand U3333 (N_3333,N_879,N_2292);
nor U3334 (N_3334,N_702,N_1040);
nand U3335 (N_3335,N_36,N_1540);
nand U3336 (N_3336,N_1862,N_1271);
nand U3337 (N_3337,N_2368,N_2895);
and U3338 (N_3338,N_2926,N_2287);
nor U3339 (N_3339,N_2494,N_2931);
or U3340 (N_3340,N_1944,N_231);
xor U3341 (N_3341,N_2896,N_1912);
and U3342 (N_3342,N_1685,N_2365);
and U3343 (N_3343,N_1843,N_1378);
or U3344 (N_3344,N_2781,N_530);
nand U3345 (N_3345,N_1553,N_2076);
nand U3346 (N_3346,N_2684,N_2001);
nor U3347 (N_3347,N_604,N_1732);
nand U3348 (N_3348,N_2314,N_593);
or U3349 (N_3349,N_1480,N_1196);
and U3350 (N_3350,N_1245,N_185);
nor U3351 (N_3351,N_1355,N_286);
or U3352 (N_3352,N_343,N_135);
and U3353 (N_3353,N_1404,N_1804);
nand U3354 (N_3354,N_888,N_1112);
and U3355 (N_3355,N_1177,N_2435);
and U3356 (N_3356,N_896,N_955);
or U3357 (N_3357,N_1997,N_765);
and U3358 (N_3358,N_1516,N_2203);
xnor U3359 (N_3359,N_62,N_1938);
nand U3360 (N_3360,N_262,N_785);
xnor U3361 (N_3361,N_1664,N_2546);
nand U3362 (N_3362,N_160,N_2876);
or U3363 (N_3363,N_2414,N_2952);
and U3364 (N_3364,N_1607,N_1338);
and U3365 (N_3365,N_1631,N_1184);
nor U3366 (N_3366,N_1543,N_2595);
or U3367 (N_3367,N_311,N_1729);
and U3368 (N_3368,N_2569,N_224);
and U3369 (N_3369,N_2764,N_836);
nor U3370 (N_3370,N_918,N_2906);
xnor U3371 (N_3371,N_877,N_636);
or U3372 (N_3372,N_2854,N_1534);
nor U3373 (N_3373,N_2623,N_1445);
and U3374 (N_3374,N_65,N_1058);
and U3375 (N_3375,N_1625,N_1332);
or U3376 (N_3376,N_2391,N_2179);
nor U3377 (N_3377,N_612,N_1004);
nand U3378 (N_3378,N_649,N_2304);
and U3379 (N_3379,N_295,N_1110);
and U3380 (N_3380,N_565,N_1822);
nor U3381 (N_3381,N_2062,N_1477);
nor U3382 (N_3382,N_805,N_76);
and U3383 (N_3383,N_2551,N_772);
nand U3384 (N_3384,N_2361,N_2652);
and U3385 (N_3385,N_1400,N_2540);
nand U3386 (N_3386,N_754,N_1118);
or U3387 (N_3387,N_2205,N_1303);
or U3388 (N_3388,N_562,N_2267);
or U3389 (N_3389,N_2288,N_1996);
nor U3390 (N_3390,N_1343,N_2161);
and U3391 (N_3391,N_2409,N_1865);
nor U3392 (N_3392,N_2211,N_2412);
nor U3393 (N_3393,N_1531,N_1615);
and U3394 (N_3394,N_2128,N_1673);
nor U3395 (N_3395,N_2503,N_2981);
nor U3396 (N_3396,N_2654,N_853);
or U3397 (N_3397,N_1567,N_2752);
nand U3398 (N_3398,N_2653,N_2059);
nand U3399 (N_3399,N_1854,N_555);
nand U3400 (N_3400,N_976,N_2613);
nor U3401 (N_3401,N_205,N_1757);
and U3402 (N_3402,N_2104,N_868);
xnor U3403 (N_3403,N_508,N_194);
and U3404 (N_3404,N_1688,N_659);
or U3405 (N_3405,N_2734,N_992);
xor U3406 (N_3406,N_2413,N_1978);
or U3407 (N_3407,N_2069,N_2913);
and U3408 (N_3408,N_1473,N_2571);
or U3409 (N_3409,N_1965,N_1764);
nor U3410 (N_3410,N_1014,N_2883);
or U3411 (N_3411,N_2226,N_1488);
nor U3412 (N_3412,N_2681,N_1454);
xor U3413 (N_3413,N_1248,N_2933);
nor U3414 (N_3414,N_2350,N_698);
nor U3415 (N_3415,N_1,N_2201);
or U3416 (N_3416,N_2541,N_2756);
nor U3417 (N_3417,N_2227,N_1634);
or U3418 (N_3418,N_1242,N_1674);
nand U3419 (N_3419,N_470,N_276);
xnor U3420 (N_3420,N_1213,N_2443);
or U3421 (N_3421,N_2056,N_671);
or U3422 (N_3422,N_2094,N_2828);
or U3423 (N_3423,N_875,N_934);
nor U3424 (N_3424,N_2937,N_2306);
or U3425 (N_3425,N_2219,N_1309);
nand U3426 (N_3426,N_2332,N_25);
nor U3427 (N_3427,N_615,N_358);
xor U3428 (N_3428,N_906,N_2944);
and U3429 (N_3429,N_1629,N_1889);
nand U3430 (N_3430,N_2863,N_2581);
and U3431 (N_3431,N_2768,N_1933);
nand U3432 (N_3432,N_1975,N_2253);
xnor U3433 (N_3433,N_813,N_1721);
xor U3434 (N_3434,N_229,N_1991);
and U3435 (N_3435,N_1294,N_592);
and U3436 (N_3436,N_448,N_202);
xnor U3437 (N_3437,N_1870,N_1850);
nor U3438 (N_3438,N_1424,N_1906);
xnor U3439 (N_3439,N_2486,N_1037);
and U3440 (N_3440,N_267,N_654);
and U3441 (N_3441,N_1831,N_2482);
xnor U3442 (N_3442,N_653,N_263);
and U3443 (N_3443,N_2108,N_2274);
and U3444 (N_3444,N_798,N_2890);
and U3445 (N_3445,N_2529,N_1252);
and U3446 (N_3446,N_222,N_1786);
and U3447 (N_3447,N_1597,N_1792);
and U3448 (N_3448,N_1665,N_2844);
or U3449 (N_3449,N_2618,N_1527);
nand U3450 (N_3450,N_1951,N_2799);
and U3451 (N_3451,N_2680,N_2039);
xnor U3452 (N_3452,N_1420,N_1439);
xnor U3453 (N_3453,N_2316,N_419);
or U3454 (N_3454,N_1115,N_88);
or U3455 (N_3455,N_2015,N_498);
nand U3456 (N_3456,N_421,N_2918);
nor U3457 (N_3457,N_983,N_1535);
or U3458 (N_3458,N_783,N_252);
and U3459 (N_3459,N_1418,N_2085);
or U3460 (N_3460,N_1090,N_2531);
nor U3461 (N_3461,N_1760,N_2586);
nor U3462 (N_3462,N_2242,N_1820);
and U3463 (N_3463,N_2634,N_2711);
and U3464 (N_3464,N_2499,N_734);
or U3465 (N_3465,N_1848,N_367);
or U3466 (N_3466,N_2930,N_1998);
xor U3467 (N_3467,N_2935,N_1867);
xor U3468 (N_3468,N_2337,N_2648);
and U3469 (N_3469,N_848,N_897);
xor U3470 (N_3470,N_873,N_2942);
or U3471 (N_3471,N_2923,N_710);
xnor U3472 (N_3472,N_2676,N_1536);
nor U3473 (N_3473,N_2955,N_83);
or U3474 (N_3474,N_2770,N_2962);
nor U3475 (N_3475,N_2658,N_2496);
nand U3476 (N_3476,N_450,N_905);
or U3477 (N_3477,N_1485,N_2842);
and U3478 (N_3478,N_2312,N_1563);
and U3479 (N_3479,N_1286,N_2136);
nor U3480 (N_3480,N_399,N_1190);
xnor U3481 (N_3481,N_777,N_726);
or U3482 (N_3482,N_829,N_2483);
xor U3483 (N_3483,N_2212,N_244);
and U3484 (N_3484,N_499,N_784);
xor U3485 (N_3485,N_1059,N_2826);
nand U3486 (N_3486,N_1336,N_1222);
xor U3487 (N_3487,N_2795,N_2213);
or U3488 (N_3488,N_826,N_1915);
and U3489 (N_3489,N_176,N_527);
xor U3490 (N_3490,N_2440,N_234);
nor U3491 (N_3491,N_2106,N_720);
or U3492 (N_3492,N_622,N_1509);
xor U3493 (N_3493,N_2221,N_1879);
and U3494 (N_3494,N_2959,N_1451);
xnor U3495 (N_3495,N_2504,N_1135);
nor U3496 (N_3496,N_617,N_662);
nor U3497 (N_3497,N_2986,N_518);
or U3498 (N_3498,N_2582,N_1735);
xor U3499 (N_3499,N_2520,N_11);
nand U3500 (N_3500,N_110,N_1304);
nor U3501 (N_3501,N_2196,N_192);
nand U3502 (N_3502,N_1815,N_1254);
and U3503 (N_3503,N_2907,N_2286);
or U3504 (N_3504,N_1149,N_1041);
nand U3505 (N_3505,N_2351,N_1104);
xnor U3506 (N_3506,N_1139,N_2272);
nor U3507 (N_3507,N_831,N_747);
xnor U3508 (N_3508,N_243,N_2053);
nand U3509 (N_3509,N_2054,N_486);
nor U3510 (N_3510,N_2441,N_1193);
nand U3511 (N_3511,N_1073,N_2423);
nand U3512 (N_3512,N_298,N_1387);
or U3513 (N_3513,N_1830,N_2552);
xor U3514 (N_3514,N_1728,N_1176);
or U3515 (N_3515,N_1856,N_2720);
or U3516 (N_3516,N_517,N_158);
nor U3517 (N_3517,N_2783,N_818);
xnor U3518 (N_3518,N_2019,N_715);
nand U3519 (N_3519,N_342,N_2055);
nand U3520 (N_3520,N_2112,N_645);
and U3521 (N_3521,N_603,N_1221);
nor U3522 (N_3522,N_305,N_2336);
nand U3523 (N_3523,N_124,N_1651);
and U3524 (N_3524,N_1306,N_908);
or U3525 (N_3525,N_2565,N_886);
nand U3526 (N_3526,N_2299,N_733);
or U3527 (N_3527,N_108,N_2220);
nand U3528 (N_3528,N_582,N_2488);
nor U3529 (N_3529,N_2258,N_1194);
or U3530 (N_3530,N_940,N_2892);
xnor U3531 (N_3531,N_1861,N_1747);
xnor U3532 (N_3532,N_2117,N_7);
nand U3533 (N_3533,N_800,N_21);
or U3534 (N_3534,N_2249,N_2266);
nor U3535 (N_3535,N_2462,N_2660);
nand U3536 (N_3536,N_2577,N_681);
nor U3537 (N_3537,N_2789,N_2419);
xor U3538 (N_3538,N_1529,N_2506);
or U3539 (N_3539,N_1484,N_2915);
nor U3540 (N_3540,N_967,N_2366);
xnor U3541 (N_3541,N_370,N_2574);
or U3542 (N_3542,N_2544,N_1845);
and U3543 (N_3543,N_2040,N_2465);
xnor U3544 (N_3544,N_422,N_1763);
nor U3545 (N_3545,N_2976,N_2244);
nand U3546 (N_3546,N_2111,N_77);
xor U3547 (N_3547,N_2710,N_2951);
nand U3548 (N_3548,N_680,N_2755);
xor U3549 (N_3549,N_2058,N_1661);
xnor U3550 (N_3550,N_1832,N_2721);
xor U3551 (N_3551,N_2207,N_409);
nand U3552 (N_3552,N_2888,N_810);
nand U3553 (N_3553,N_633,N_114);
nand U3554 (N_3554,N_1326,N_1608);
nand U3555 (N_3555,N_362,N_344);
xor U3556 (N_3556,N_218,N_1287);
and U3557 (N_3557,N_349,N_1595);
nor U3558 (N_3558,N_2919,N_1539);
nand U3559 (N_3559,N_209,N_122);
xor U3560 (N_3560,N_1062,N_2647);
nand U3561 (N_3561,N_1564,N_1873);
or U3562 (N_3562,N_1240,N_1612);
or U3563 (N_3563,N_2014,N_1671);
and U3564 (N_3564,N_1455,N_1613);
xor U3565 (N_3565,N_1574,N_2387);
xnor U3566 (N_3566,N_1273,N_434);
or U3567 (N_3567,N_755,N_1211);
and U3568 (N_3568,N_139,N_203);
xor U3569 (N_3569,N_1279,N_1970);
and U3570 (N_3570,N_1942,N_2943);
or U3571 (N_3571,N_1162,N_1829);
nand U3572 (N_3572,N_2562,N_847);
and U3573 (N_3573,N_1081,N_1803);
and U3574 (N_3574,N_1884,N_1447);
nand U3575 (N_3575,N_1609,N_1839);
or U3576 (N_3576,N_2199,N_18);
nor U3577 (N_3577,N_1349,N_2998);
xor U3578 (N_3578,N_1945,N_428);
or U3579 (N_3579,N_2105,N_2530);
xor U3580 (N_3580,N_1750,N_2277);
and U3581 (N_3581,N_2169,N_452);
nor U3582 (N_3582,N_889,N_2188);
nor U3583 (N_3583,N_171,N_1030);
nand U3584 (N_3584,N_2694,N_2792);
xnor U3585 (N_3585,N_1136,N_155);
and U3586 (N_3586,N_1275,N_352);
nor U3587 (N_3587,N_2086,N_2355);
nand U3588 (N_3588,N_1493,N_956);
nand U3589 (N_3589,N_225,N_1948);
and U3590 (N_3590,N_1931,N_2276);
nand U3591 (N_3591,N_2992,N_824);
or U3592 (N_3592,N_738,N_1201);
nand U3593 (N_3593,N_1550,N_986);
nor U3594 (N_3594,N_974,N_893);
nor U3595 (N_3595,N_2319,N_371);
nand U3596 (N_3596,N_1566,N_405);
and U3597 (N_3597,N_2771,N_283);
xor U3598 (N_3598,N_580,N_162);
xnor U3599 (N_3599,N_629,N_1247);
and U3600 (N_3600,N_1409,N_227);
nand U3601 (N_3601,N_1947,N_1800);
or U3602 (N_3602,N_164,N_1377);
xor U3603 (N_3603,N_2706,N_505);
nor U3604 (N_3604,N_1069,N_1681);
nor U3605 (N_3605,N_1042,N_2689);
nand U3606 (N_3606,N_1319,N_2757);
nand U3607 (N_3607,N_512,N_175);
nor U3608 (N_3608,N_1780,N_2987);
or U3609 (N_3609,N_1770,N_247);
or U3610 (N_3610,N_1383,N_1834);
nand U3611 (N_3611,N_2746,N_1797);
and U3612 (N_3612,N_1755,N_459);
or U3613 (N_3613,N_2811,N_1393);
nor U3614 (N_3614,N_242,N_1503);
or U3615 (N_3615,N_1325,N_670);
nand U3616 (N_3616,N_55,N_1583);
nand U3617 (N_3617,N_188,N_2966);
and U3618 (N_3618,N_1899,N_1186);
or U3619 (N_3619,N_472,N_1432);
nor U3620 (N_3620,N_1565,N_2524);
nor U3621 (N_3621,N_359,N_2882);
nand U3622 (N_3622,N_1144,N_914);
xnor U3623 (N_3623,N_1178,N_1733);
nand U3624 (N_3624,N_839,N_1756);
xnor U3625 (N_3625,N_1470,N_1278);
nor U3626 (N_3626,N_808,N_1606);
xor U3627 (N_3627,N_1148,N_416);
xor U3628 (N_3628,N_1890,N_677);
nor U3629 (N_3629,N_91,N_347);
nand U3630 (N_3630,N_749,N_447);
and U3631 (N_3631,N_154,N_985);
xor U3632 (N_3632,N_1743,N_49);
xor U3633 (N_3633,N_173,N_2853);
and U3634 (N_3634,N_73,N_2468);
xnor U3635 (N_3635,N_1926,N_543);
nor U3636 (N_3636,N_2794,N_581);
nand U3637 (N_3637,N_2233,N_993);
and U3638 (N_3638,N_1497,N_1623);
xor U3639 (N_3639,N_1637,N_1739);
or U3640 (N_3640,N_1026,N_1003);
and U3641 (N_3641,N_990,N_1605);
xnor U3642 (N_3642,N_1683,N_2079);
and U3643 (N_3643,N_968,N_2013);
and U3644 (N_3644,N_1013,N_2310);
and U3645 (N_3645,N_2396,N_1407);
or U3646 (N_3646,N_2237,N_1905);
and U3647 (N_3647,N_1600,N_1882);
nor U3648 (N_3648,N_2766,N_338);
nand U3649 (N_3649,N_2988,N_182);
nor U3650 (N_3650,N_1341,N_301);
nor U3651 (N_3651,N_256,N_2425);
xnor U3652 (N_3652,N_2599,N_1074);
nand U3653 (N_3653,N_1672,N_2979);
or U3654 (N_3654,N_5,N_2960);
xnor U3655 (N_3655,N_1056,N_2518);
nand U3656 (N_3656,N_1819,N_935);
and U3657 (N_3657,N_2005,N_2313);
and U3658 (N_3658,N_501,N_1675);
nor U3659 (N_3659,N_1123,N_1072);
nand U3660 (N_3660,N_1622,N_217);
xnor U3661 (N_3661,N_1097,N_1414);
or U3662 (N_3662,N_120,N_201);
nor U3663 (N_3663,N_804,N_950);
and U3664 (N_3664,N_1864,N_1362);
or U3665 (N_3665,N_1483,N_1091);
and U3666 (N_3666,N_2025,N_599);
or U3667 (N_3667,N_675,N_2210);
nand U3668 (N_3668,N_2478,N_93);
xor U3669 (N_3669,N_541,N_2874);
nand U3670 (N_3670,N_2973,N_361);
or U3671 (N_3671,N_485,N_2156);
nor U3672 (N_3672,N_95,N_2851);
or U3673 (N_3673,N_2119,N_1598);
nor U3674 (N_3674,N_2324,N_2601);
and U3675 (N_3675,N_1435,N_2204);
and U3676 (N_3676,N_142,N_1419);
or U3677 (N_3677,N_1237,N_1095);
nand U3678 (N_3678,N_2329,N_378);
nor U3679 (N_3679,N_2107,N_1442);
nand U3680 (N_3680,N_1917,N_464);
xor U3681 (N_3681,N_1987,N_2291);
or U3682 (N_3682,N_2814,N_2215);
xor U3683 (N_3683,N_392,N_1841);
xor U3684 (N_3684,N_144,N_1496);
nor U3685 (N_3685,N_166,N_2693);
xnor U3686 (N_3686,N_2176,N_33);
nor U3687 (N_3687,N_2125,N_41);
nand U3688 (N_3688,N_1712,N_1709);
nor U3689 (N_3689,N_2016,N_494);
xor U3690 (N_3690,N_1374,N_814);
nor U3691 (N_3691,N_2673,N_2026);
xor U3692 (N_3692,N_2270,N_1101);
or U3693 (N_3693,N_2784,N_2773);
nand U3694 (N_3694,N_1100,N_415);
and U3695 (N_3695,N_1482,N_1195);
or U3696 (N_3696,N_821,N_1269);
and U3697 (N_3697,N_2311,N_2697);
and U3698 (N_3698,N_2265,N_881);
or U3699 (N_3699,N_1350,N_2455);
nor U3700 (N_3700,N_223,N_1152);
nor U3701 (N_3701,N_2869,N_1067);
and U3702 (N_3702,N_1061,N_1045);
or U3703 (N_3703,N_2864,N_966);
and U3704 (N_3704,N_39,N_2367);
xnor U3705 (N_3705,N_1667,N_567);
or U3706 (N_3706,N_503,N_753);
and U3707 (N_3707,N_2782,N_1434);
and U3708 (N_3708,N_364,N_2763);
nand U3709 (N_3709,N_1243,N_576);
xor U3710 (N_3710,N_2263,N_479);
and U3711 (N_3711,N_469,N_1762);
xor U3712 (N_3712,N_272,N_513);
and U3713 (N_3713,N_2038,N_1345);
or U3714 (N_3714,N_854,N_1046);
or U3715 (N_3715,N_2078,N_1205);
xor U3716 (N_3716,N_1092,N_183);
xor U3717 (N_3717,N_1235,N_2411);
or U3718 (N_3718,N_867,N_2912);
nand U3719 (N_3719,N_23,N_1638);
nand U3720 (N_3720,N_2539,N_458);
nor U3721 (N_3721,N_2339,N_998);
and U3722 (N_3722,N_947,N_2262);
nor U3723 (N_3723,N_2982,N_1935);
xor U3724 (N_3724,N_2289,N_403);
nor U3725 (N_3725,N_2600,N_1738);
nand U3726 (N_3726,N_2554,N_2222);
nand U3727 (N_3727,N_949,N_2031);
or U3728 (N_3728,N_2232,N_2305);
and U3729 (N_3729,N_778,N_1039);
nor U3730 (N_3730,N_1198,N_212);
and U3731 (N_3731,N_1585,N_2398);
xor U3732 (N_3732,N_178,N_1358);
xor U3733 (N_3733,N_2731,N_942);
and U3734 (N_3734,N_1686,N_737);
nor U3735 (N_3735,N_237,N_1620);
and U3736 (N_3736,N_1920,N_2141);
xor U3737 (N_3737,N_2103,N_731);
xor U3738 (N_3738,N_2963,N_289);
xor U3739 (N_3739,N_2279,N_815);
nor U3740 (N_3740,N_2832,N_152);
or U3741 (N_3741,N_953,N_2223);
and U3742 (N_3742,N_336,N_2495);
nor U3743 (N_3743,N_1908,N_2448);
nand U3744 (N_3744,N_1241,N_2502);
and U3745 (N_3745,N_339,N_2195);
xor U3746 (N_3746,N_752,N_1807);
and U3747 (N_3747,N_1165,N_2255);
and U3748 (N_3748,N_2909,N_2386);
and U3749 (N_3749,N_919,N_290);
nand U3750 (N_3750,N_1633,N_2991);
xor U3751 (N_3751,N_2303,N_2777);
or U3752 (N_3752,N_2261,N_758);
or U3753 (N_3753,N_2949,N_1989);
xnor U3754 (N_3754,N_770,N_2526);
xnor U3755 (N_3755,N_1385,N_988);
or U3756 (N_3756,N_1024,N_1217);
nor U3757 (N_3757,N_1508,N_1900);
nor U3758 (N_3758,N_2407,N_2743);
or U3759 (N_3759,N_884,N_315);
nor U3760 (N_3760,N_872,N_1523);
nand U3761 (N_3761,N_2732,N_845);
xor U3762 (N_3762,N_197,N_1492);
nand U3763 (N_3763,N_2964,N_2118);
and U3764 (N_3764,N_1723,N_2231);
nand U3765 (N_3765,N_682,N_2363);
or U3766 (N_3766,N_692,N_12);
or U3767 (N_3767,N_602,N_199);
nand U3768 (N_3768,N_117,N_1893);
nand U3769 (N_3769,N_684,N_1085);
xnor U3770 (N_3770,N_1145,N_2114);
and U3771 (N_3771,N_1265,N_954);
and U3772 (N_3772,N_2393,N_1096);
nand U3773 (N_3773,N_2426,N_2452);
xor U3774 (N_3774,N_2446,N_509);
xor U3775 (N_3775,N_1315,N_773);
nor U3776 (N_3776,N_1710,N_827);
nor U3777 (N_3777,N_789,N_2664);
nor U3778 (N_3778,N_2904,N_1285);
xor U3779 (N_3779,N_909,N_2857);
and U3780 (N_3780,N_2142,N_885);
and U3781 (N_3781,N_195,N_1251);
nand U3782 (N_3782,N_1966,N_2625);
xnor U3783 (N_3783,N_407,N_1525);
and U3784 (N_3784,N_2097,N_2750);
xor U3785 (N_3785,N_1281,N_66);
nand U3786 (N_3786,N_2044,N_2604);
and U3787 (N_3787,N_2457,N_2663);
nor U3788 (N_3788,N_2975,N_1087);
xor U3789 (N_3789,N_1616,N_704);
and U3790 (N_3790,N_1397,N_191);
and U3791 (N_3791,N_774,N_788);
and U3792 (N_3792,N_126,N_564);
and U3793 (N_3793,N_987,N_2837);
nand U3794 (N_3794,N_1471,N_2283);
nor U3795 (N_3795,N_444,N_2383);
xor U3796 (N_3796,N_1777,N_619);
nor U3797 (N_3797,N_98,N_2598);
and U3798 (N_3798,N_46,N_2122);
xor U3799 (N_3799,N_181,N_2377);
and U3800 (N_3800,N_2894,N_1852);
xnor U3801 (N_3801,N_2590,N_319);
xor U3802 (N_3802,N_930,N_48);
or U3803 (N_3803,N_982,N_14);
or U3804 (N_3804,N_2358,N_2378);
and U3805 (N_3805,N_260,N_1427);
nand U3806 (N_3806,N_891,N_624);
xnor U3807 (N_3807,N_24,N_938);
xor U3808 (N_3808,N_467,N_89);
or U3809 (N_3809,N_1708,N_1340);
or U3810 (N_3810,N_431,N_856);
nand U3811 (N_3811,N_1918,N_1175);
and U3812 (N_3812,N_1228,N_475);
nand U3813 (N_3813,N_190,N_823);
nand U3814 (N_3814,N_1226,N_2072);
and U3815 (N_3815,N_1532,N_1047);
nor U3816 (N_3816,N_38,N_2728);
xnor U3817 (N_3817,N_729,N_2800);
and U3818 (N_3818,N_2729,N_2381);
nand U3819 (N_3819,N_948,N_1720);
and U3820 (N_3820,N_186,N_1370);
and U3821 (N_3821,N_294,N_1993);
nand U3822 (N_3822,N_423,N_2880);
nand U3823 (N_3823,N_1678,N_1206);
and U3824 (N_3824,N_1468,N_1440);
xor U3825 (N_3825,N_2326,N_2424);
xor U3826 (N_3826,N_728,N_2985);
and U3827 (N_3827,N_1498,N_381);
nand U3828 (N_3828,N_1066,N_1849);
nand U3829 (N_3829,N_1967,N_883);
and U3830 (N_3830,N_997,N_2260);
xor U3831 (N_3831,N_1043,N_2603);
xor U3832 (N_3832,N_2860,N_2672);
and U3833 (N_3833,N_2649,N_648);
xor U3834 (N_3834,N_750,N_1799);
nand U3835 (N_3835,N_2022,N_1964);
or U3836 (N_3836,N_1640,N_1979);
and U3837 (N_3837,N_1898,N_1699);
or U3838 (N_3838,N_2767,N_2724);
nor U3839 (N_3839,N_1811,N_442);
nand U3840 (N_3840,N_2144,N_30);
nand U3841 (N_3841,N_2123,N_2631);
nand U3842 (N_3842,N_2051,N_1544);
xnor U3843 (N_3843,N_1022,N_623);
nor U3844 (N_3844,N_2489,N_393);
nor U3845 (N_3845,N_1344,N_1768);
nor U3846 (N_3846,N_285,N_1940);
nor U3847 (N_3847,N_2830,N_326);
or U3848 (N_3848,N_2801,N_1125);
or U3849 (N_3849,N_2505,N_2461);
or U3850 (N_3850,N_22,N_1578);
or U3851 (N_3851,N_2300,N_2192);
nor U3852 (N_3852,N_2029,N_2967);
nand U3853 (N_3853,N_1172,N_59);
and U3854 (N_3854,N_1270,N_1552);
or U3855 (N_3855,N_1983,N_709);
and U3856 (N_3856,N_1980,N_507);
or U3857 (N_3857,N_1417,N_2395);
nor U3858 (N_3858,N_2610,N_1449);
or U3859 (N_3859,N_455,N_1376);
nand U3860 (N_3860,N_2807,N_2439);
and U3861 (N_3861,N_794,N_2251);
or U3862 (N_3862,N_1075,N_685);
or U3863 (N_3863,N_99,N_2315);
and U3864 (N_3864,N_1639,N_1117);
nor U3865 (N_3865,N_2779,N_2308);
and U3866 (N_3866,N_2120,N_1430);
xor U3867 (N_3867,N_482,N_2645);
nand U3868 (N_3868,N_927,N_743);
xor U3869 (N_3869,N_2158,N_404);
nor U3870 (N_3870,N_334,N_577);
nand U3871 (N_3871,N_1971,N_321);
or U3872 (N_3872,N_297,N_269);
and U3873 (N_3873,N_4,N_1891);
or U3874 (N_3874,N_1331,N_588);
nor U3875 (N_3875,N_2131,N_1885);
nand U3876 (N_3876,N_1208,N_140);
or U3877 (N_3877,N_2677,N_718);
and U3878 (N_3878,N_714,N_1737);
xor U3879 (N_3879,N_1347,N_1628);
and U3880 (N_3880,N_2472,N_2437);
and U3881 (N_3881,N_584,N_172);
and U3882 (N_3882,N_2594,N_2796);
nand U3883 (N_3883,N_598,N_1260);
nand U3884 (N_3884,N_2983,N_1089);
and U3885 (N_3885,N_390,N_756);
xor U3886 (N_3886,N_911,N_275);
nor U3887 (N_3887,N_2740,N_2214);
xor U3888 (N_3888,N_316,N_143);
nand U3889 (N_3889,N_323,N_1299);
nand U3890 (N_3890,N_1663,N_116);
nor U3891 (N_3891,N_2153,N_1517);
and U3892 (N_3892,N_240,N_790);
or U3893 (N_3893,N_970,N_376);
nand U3894 (N_3894,N_575,N_2401);
or U3895 (N_3895,N_1846,N_258);
or U3896 (N_3896,N_1389,N_1082);
nand U3897 (N_3897,N_1121,N_803);
nor U3898 (N_3898,N_398,N_1599);
and U3899 (N_3899,N_1446,N_493);
nor U3900 (N_3900,N_2687,N_551);
or U3901 (N_3901,N_878,N_2513);
or U3902 (N_3902,N_1610,N_2990);
nand U3903 (N_3903,N_356,N_2191);
and U3904 (N_3904,N_2536,N_1318);
xor U3905 (N_3905,N_1181,N_451);
xnor U3906 (N_3906,N_2946,N_1137);
nand U3907 (N_3907,N_679,N_2247);
or U3908 (N_3908,N_1654,N_2050);
xnor U3909 (N_3909,N_1282,N_1973);
nand U3910 (N_3910,N_1957,N_614);
nor U3911 (N_3911,N_1182,N_870);
and U3912 (N_3912,N_1953,N_2011);
xor U3913 (N_3913,N_694,N_2567);
or U3914 (N_3914,N_2269,N_2596);
nor U3915 (N_3915,N_2813,N_2459);
nand U3916 (N_3916,N_2392,N_730);
or U3917 (N_3917,N_2127,N_621);
or U3918 (N_3918,N_2021,N_2727);
or U3919 (N_3919,N_1052,N_1388);
xnor U3920 (N_3920,N_497,N_554);
nor U3921 (N_3921,N_2514,N_2202);
or U3922 (N_3922,N_2152,N_2527);
nor U3923 (N_3923,N_1203,N_625);
and U3924 (N_3924,N_1894,N_904);
or U3925 (N_3925,N_632,N_2674);
xor U3926 (N_3926,N_2230,N_2126);
and U3927 (N_3927,N_2717,N_1171);
xor U3928 (N_3928,N_1650,N_2346);
xnor U3929 (N_3929,N_2182,N_8);
xor U3930 (N_3930,N_797,N_2971);
nor U3931 (N_3931,N_711,N_2338);
nand U3932 (N_3932,N_430,N_2328);
nor U3933 (N_3933,N_2831,N_2284);
nor U3934 (N_3934,N_2932,N_907);
nand U3935 (N_3935,N_2641,N_2958);
nand U3936 (N_3936,N_1490,N_900);
and U3937 (N_3937,N_1874,N_1911);
or U3938 (N_3938,N_2873,N_1108);
nor U3939 (N_3939,N_1405,N_1033);
and U3940 (N_3940,N_308,N_2379);
nand U3941 (N_3941,N_2866,N_1048);
or U3942 (N_3942,N_522,N_287);
nor U3943 (N_3943,N_2819,N_1771);
nor U3944 (N_3944,N_1670,N_87);
xor U3945 (N_3945,N_2961,N_2173);
nand U3946 (N_3946,N_1253,N_1725);
nand U3947 (N_3947,N_1057,N_2682);
nor U3948 (N_3948,N_2583,N_184);
or U3949 (N_3949,N_56,N_1524);
nand U3950 (N_3950,N_2493,N_1380);
nand U3951 (N_3951,N_1163,N_1627);
or U3952 (N_3952,N_1386,N_1694);
xnor U3953 (N_3953,N_2089,N_2893);
or U3954 (N_3954,N_302,N_17);
xnor U3955 (N_3955,N_855,N_2608);
and U3956 (N_3956,N_946,N_2557);
or U3957 (N_3957,N_807,N_1689);
xnor U3958 (N_3958,N_2836,N_1421);
or U3959 (N_3959,N_2476,N_2716);
nor U3960 (N_3960,N_1314,N_1450);
or U3961 (N_3961,N_1308,N_759);
or U3962 (N_3962,N_739,N_1593);
nand U3963 (N_3963,N_2229,N_697);
nand U3964 (N_3964,N_515,N_156);
and U3965 (N_3965,N_2891,N_2620);
or U3966 (N_3966,N_2791,N_1886);
and U3967 (N_3967,N_2068,N_2578);
or U3968 (N_3968,N_1415,N_2922);
xnor U3969 (N_3969,N_786,N_174);
nand U3970 (N_3970,N_972,N_2322);
xnor U3971 (N_3971,N_1897,N_2838);
nor U3972 (N_3972,N_1138,N_313);
and U3973 (N_3973,N_1373,N_1438);
xor U3974 (N_3974,N_1924,N_894);
or U3975 (N_3975,N_1695,N_1204);
xor U3976 (N_3976,N_850,N_642);
or U3977 (N_3977,N_1961,N_1185);
xor U3978 (N_3978,N_1923,N_2879);
or U3979 (N_3979,N_1132,N_2908);
and U3980 (N_3980,N_330,N_84);
xor U3981 (N_3981,N_717,N_2980);
nor U3982 (N_3982,N_2573,N_1895);
nor U3983 (N_3983,N_1549,N_1765);
xnor U3984 (N_3984,N_1705,N_2268);
xnor U3985 (N_3985,N_1857,N_215);
nand U3986 (N_3986,N_2559,N_559);
nand U3987 (N_3987,N_2404,N_548);
nor U3988 (N_3988,N_1456,N_2816);
xor U3989 (N_3989,N_1000,N_241);
and U3990 (N_3990,N_1569,N_1858);
and U3991 (N_3991,N_1956,N_2995);
nor U3992 (N_3992,N_2829,N_899);
nor U3993 (N_3993,N_2701,N_151);
xnor U3994 (N_3994,N_1588,N_2748);
and U3995 (N_3995,N_1207,N_700);
and U3996 (N_3996,N_1215,N_744);
nor U3997 (N_3997,N_1645,N_123);
nand U3998 (N_3998,N_943,N_2429);
or U3999 (N_3999,N_2174,N_2745);
nor U4000 (N_4000,N_573,N_341);
or U4001 (N_4001,N_2852,N_1576);
or U4002 (N_4002,N_929,N_1437);
nand U4003 (N_4003,N_456,N_1825);
and U4004 (N_4004,N_2145,N_1877);
nand U4005 (N_4005,N_1130,N_977);
and U4006 (N_4006,N_1291,N_1422);
xor U4007 (N_4007,N_1934,N_2187);
xnor U4008 (N_4008,N_351,N_806);
nor U4009 (N_4009,N_1321,N_2382);
and U4010 (N_4010,N_570,N_1869);
xnor U4011 (N_4011,N_2027,N_1960);
nand U4012 (N_4012,N_2290,N_922);
or U4013 (N_4013,N_2786,N_1263);
and U4014 (N_4014,N_2993,N_2885);
xnor U4015 (N_4015,N_822,N_1379);
xnor U4016 (N_4016,N_1518,N_1520);
nand U4017 (N_4017,N_474,N_2841);
nand U4018 (N_4018,N_1107,N_1706);
nand U4019 (N_4019,N_2442,N_2264);
nor U4020 (N_4020,N_2714,N_2373);
xor U4021 (N_4021,N_713,N_639);
xor U4022 (N_4022,N_996,N_2510);
nor U4023 (N_4023,N_1356,N_463);
nor U4024 (N_4024,N_620,N_544);
xnor U4025 (N_4025,N_1826,N_534);
nand U4026 (N_4026,N_484,N_1348);
nand U4027 (N_4027,N_655,N_1754);
nand U4028 (N_4028,N_586,N_1950);
nand U4029 (N_4029,N_2197,N_2238);
xnor U4030 (N_4030,N_473,N_1624);
or U4031 (N_4031,N_1371,N_2487);
or U4032 (N_4032,N_121,N_1300);
or U4033 (N_4033,N_1301,N_2041);
nor U4034 (N_4034,N_1810,N_2508);
and U4035 (N_4035,N_1618,N_2349);
nand U4036 (N_4036,N_2098,N_1312);
nor U4037 (N_4037,N_2467,N_1088);
nor U4038 (N_4038,N_1500,N_557);
nand U4039 (N_4039,N_213,N_991);
and U4040 (N_4040,N_1354,N_628);
and U4041 (N_4041,N_2190,N_2954);
xor U4042 (N_4042,N_1360,N_27);
or U4043 (N_4043,N_1448,N_768);
nand U4044 (N_4044,N_159,N_2606);
and U4045 (N_4045,N_2870,N_2166);
and U4046 (N_4046,N_1272,N_1521);
nand U4047 (N_4047,N_1969,N_1594);
and U4048 (N_4048,N_2394,N_2584);
and U4049 (N_4049,N_491,N_1632);
nand U4050 (N_4050,N_15,N_1774);
nand U4051 (N_4051,N_210,N_561);
nor U4052 (N_4052,N_1526,N_2181);
xor U4053 (N_4053,N_1134,N_1572);
xor U4054 (N_4054,N_2561,N_1511);
or U4055 (N_4055,N_1368,N_2034);
or U4056 (N_4056,N_2035,N_1833);
nand U4057 (N_4057,N_2805,N_1717);
or U4058 (N_4058,N_145,N_1127);
and U4059 (N_4059,N_235,N_2978);
nand U4060 (N_4060,N_1436,N_2165);
and U4061 (N_4061,N_1776,N_1212);
nor U4062 (N_4062,N_611,N_2194);
nor U4063 (N_4063,N_426,N_406);
xnor U4064 (N_4064,N_701,N_2012);
and U4065 (N_4065,N_2241,N_2525);
xnor U4066 (N_4066,N_2132,N_552);
or U4067 (N_4067,N_1649,N_558);
nand U4068 (N_4068,N_801,N_980);
nand U4069 (N_4069,N_1545,N_746);
nand U4070 (N_4070,N_1232,N_840);
or U4071 (N_4071,N_401,N_2248);
nand U4072 (N_4072,N_862,N_106);
and U4073 (N_4073,N_1411,N_2522);
nor U4074 (N_4074,N_1458,N_740);
nor U4075 (N_4075,N_1642,N_1510);
nand U4076 (N_4076,N_1339,N_2558);
and U4077 (N_4077,N_1802,N_1116);
nor U4078 (N_4078,N_104,N_664);
nand U4079 (N_4079,N_331,N_2096);
or U4080 (N_4080,N_2637,N_1693);
xnor U4081 (N_4081,N_2997,N_2886);
nor U4082 (N_4082,N_496,N_2257);
nand U4083 (N_4083,N_1658,N_901);
and U4084 (N_4084,N_1431,N_1173);
nand U4085 (N_4085,N_1219,N_2785);
nand U4086 (N_4086,N_2856,N_1863);
nand U4087 (N_4087,N_1731,N_1230);
and U4088 (N_4088,N_578,N_1662);
nor U4089 (N_4089,N_928,N_2134);
nor U4090 (N_4090,N_1702,N_2281);
or U4091 (N_4091,N_1333,N_1972);
or U4092 (N_4092,N_1844,N_2389);
xnor U4093 (N_4093,N_2088,N_438);
or U4094 (N_4094,N_2686,N_563);
nor U4095 (N_4095,N_300,N_2357);
nor U4096 (N_4096,N_760,N_1031);
or U4097 (N_4097,N_1766,N_1793);
and U4098 (N_4098,N_211,N_2259);
or U4099 (N_4099,N_1952,N_2850);
xnor U4100 (N_4100,N_1621,N_1636);
nand U4101 (N_4101,N_1719,N_1244);
nor U4102 (N_4102,N_2061,N_440);
xor U4103 (N_4103,N_476,N_1169);
and U4104 (N_4104,N_2840,N_1453);
nor U4105 (N_4105,N_1949,N_333);
and U4106 (N_4106,N_536,N_1395);
xor U4107 (N_4107,N_1113,N_1866);
or U4108 (N_4108,N_133,N_936);
and U4109 (N_4109,N_1328,N_1323);
and U4110 (N_4110,N_858,N_1461);
nor U4111 (N_4111,N_2063,N_2334);
nor U4112 (N_4112,N_2650,N_1324);
nor U4113 (N_4113,N_2458,N_835);
nor U4114 (N_4114,N_2591,N_2665);
and U4115 (N_4115,N_2400,N_2464);
nand U4116 (N_4116,N_660,N_2250);
and U4117 (N_4117,N_2825,N_656);
nand U4118 (N_4118,N_417,N_1167);
nor U4119 (N_4119,N_688,N_2602);
xor U4120 (N_4120,N_487,N_846);
nor U4121 (N_4121,N_2759,N_1746);
xor U4122 (N_4122,N_42,N_2177);
xnor U4123 (N_4123,N_119,N_1910);
xor U4124 (N_4124,N_1426,N_2617);
and U4125 (N_4125,N_2124,N_1224);
xnor U4126 (N_4126,N_1958,N_1872);
and U4127 (N_4127,N_2803,N_418);
and U4128 (N_4128,N_1816,N_1655);
nor U4129 (N_4129,N_2867,N_663);
and U4130 (N_4130,N_2163,N_2614);
nor U4131 (N_4131,N_699,N_2360);
or U4132 (N_4132,N_2416,N_2320);
or U4133 (N_4133,N_2430,N_2910);
or U4134 (N_4134,N_1806,N_396);
and U4135 (N_4135,N_435,N_913);
xor U4136 (N_4136,N_745,N_414);
xnor U4137 (N_4137,N_2678,N_2200);
xnor U4138 (N_4138,N_1977,N_2008);
or U4139 (N_4139,N_2082,N_107);
and U4140 (N_4140,N_2576,N_2271);
or U4141 (N_4141,N_2080,N_245);
nor U4142 (N_4142,N_2515,N_820);
nand U4143 (N_4143,N_2460,N_2449);
nand U4144 (N_4144,N_2861,N_1406);
nor U4145 (N_4145,N_2545,N_1781);
xnor U4146 (N_4146,N_2344,N_391);
and U4147 (N_4147,N_306,N_971);
nand U4148 (N_4148,N_2921,N_1963);
nor U4149 (N_4149,N_2017,N_1558);
nor U4150 (N_4150,N_634,N_1551);
nand U4151 (N_4151,N_1423,N_354);
and U4152 (N_4152,N_1290,N_1489);
nor U4153 (N_4153,N_1568,N_842);
xor U4154 (N_4154,N_468,N_2707);
or U4155 (N_4155,N_1808,N_1146);
or U4156 (N_4156,N_519,N_1261);
nand U4157 (N_4157,N_249,N_2341);
and U4158 (N_4158,N_2692,N_1974);
xnor U4159 (N_4159,N_764,N_2528);
or U4160 (N_4160,N_735,N_1840);
nor U4161 (N_4161,N_492,N_531);
nor U4162 (N_4162,N_57,N_719);
xor U4163 (N_4163,N_2159,N_819);
or U4164 (N_4164,N_232,N_1114);
nor U4165 (N_4165,N_1752,N_915);
nand U4166 (N_4166,N_2004,N_136);
xor U4167 (N_4167,N_2018,N_1851);
xor U4168 (N_4168,N_82,N_2121);
nand U4169 (N_4169,N_71,N_616);
and U4170 (N_4170,N_2234,N_90);
and U4171 (N_4171,N_1805,N_1700);
xnor U4172 (N_4172,N_637,N_2754);
or U4173 (N_4173,N_94,N_1005);
nor U4174 (N_4174,N_2622,N_2298);
xor U4175 (N_4175,N_1223,N_1463);
nor U4176 (N_4176,N_2074,N_58);
and U4177 (N_4177,N_712,N_1218);
or U4178 (N_4178,N_1020,N_2359);
and U4179 (N_4179,N_2835,N_368);
nand U4180 (N_4180,N_2938,N_502);
nand U4181 (N_4181,N_1302,N_1687);
nand U4182 (N_4182,N_2659,N_2737);
nand U4183 (N_4183,N_266,N_2730);
or U4184 (N_4184,N_2481,N_1284);
xor U4185 (N_4185,N_1335,N_2939);
xor U4186 (N_4186,N_478,N_903);
nand U4187 (N_4187,N_437,N_2903);
and U4188 (N_4188,N_2741,N_917);
nor U4189 (N_4189,N_532,N_2354);
nand U4190 (N_4190,N_1827,N_833);
xor U4191 (N_4191,N_2758,N_2408);
nand U4192 (N_4192,N_208,N_2738);
and U4193 (N_4193,N_2630,N_129);
nand U4194 (N_4194,N_2095,N_1855);
and U4195 (N_4195,N_1392,N_871);
nand U4196 (N_4196,N_1791,N_1160);
nor U4197 (N_4197,N_631,N_233);
nand U4198 (N_4198,N_2700,N_387);
or U4199 (N_4199,N_2947,N_866);
nand U4200 (N_4200,N_2845,N_2388);
nor U4201 (N_4201,N_1408,N_1365);
nand U4202 (N_4202,N_1098,N_571);
nand U4203 (N_4203,N_981,N_939);
nand U4204 (N_4204,N_2160,N_1716);
or U4205 (N_4205,N_125,N_1691);
xnor U4206 (N_4206,N_941,N_2043);
nor U4207 (N_4207,N_916,N_1441);
and U4208 (N_4208,N_2709,N_54);
xnor U4209 (N_4209,N_2640,N_1016);
nor U4210 (N_4210,N_1466,N_1381);
nand U4211 (N_4211,N_727,N_1515);
or U4212 (N_4212,N_1128,N_1602);
nand U4213 (N_4213,N_2965,N_1122);
nor U4214 (N_4214,N_2725,N_751);
xnor U4215 (N_4215,N_511,N_2713);
nor U4216 (N_4216,N_2989,N_1888);
and U4217 (N_4217,N_1070,N_2296);
nand U4218 (N_4218,N_2718,N_776);
nor U4219 (N_4219,N_1837,N_101);
and U4220 (N_4220,N_2417,N_2702);
nand U4221 (N_4221,N_2977,N_453);
xnor U4222 (N_4222,N_92,N_1256);
nor U4223 (N_4223,N_167,N_118);
xnor U4224 (N_4224,N_2899,N_2809);
xor U4225 (N_4225,N_2246,N_1932);
and U4226 (N_4226,N_1054,N_436);
and U4227 (N_4227,N_1433,N_1227);
nor U4228 (N_4228,N_2356,N_2217);
nor U4229 (N_4229,N_250,N_2917);
nor U4230 (N_4230,N_495,N_441);
nand U4231 (N_4231,N_2847,N_2147);
nor U4232 (N_4232,N_2240,N_606);
nor U4233 (N_4233,N_2817,N_1530);
and U4234 (N_4234,N_1084,N_357);
nand U4235 (N_4235,N_72,N_1928);
and U4236 (N_4236,N_568,N_2511);
nand U4237 (N_4237,N_975,N_1202);
or U4238 (N_4238,N_566,N_2626);
or U4239 (N_4239,N_638,N_1220);
nand U4240 (N_4240,N_1019,N_105);
nor U4241 (N_4241,N_1835,N_85);
and U4242 (N_4242,N_2726,N_2445);
nand U4243 (N_4243,N_1396,N_2704);
xor U4244 (N_4244,N_2621,N_2243);
and U4245 (N_4245,N_2168,N_2006);
and U4246 (N_4246,N_1233,N_1773);
and U4247 (N_4247,N_646,N_1032);
xor U4248 (N_4248,N_2000,N_2497);
and U4249 (N_4249,N_1789,N_1274);
and U4250 (N_4250,N_299,N_1939);
and U4251 (N_4251,N_742,N_74);
nor U4252 (N_4252,N_2615,N_1027);
xor U4253 (N_4253,N_2193,N_973);
nor U4254 (N_4254,N_1586,N_16);
and U4255 (N_4255,N_273,N_1079);
xor U4256 (N_4256,N_1080,N_2542);
xor U4257 (N_4257,N_2172,N_1044);
or U4258 (N_4258,N_383,N_2084);
and U4259 (N_4259,N_1547,N_1188);
nor U4260 (N_4260,N_1860,N_1102);
nor U4261 (N_4261,N_1785,N_460);
nand U4262 (N_4262,N_1842,N_1457);
and U4263 (N_4263,N_2575,N_2646);
or U4264 (N_4264,N_2969,N_2916);
or U4265 (N_4265,N_690,N_1394);
nor U4266 (N_4266,N_1076,N_667);
nor U4267 (N_4267,N_673,N_461);
xor U4268 (N_4268,N_1794,N_538);
nor U4269 (N_4269,N_2235,N_2549);
or U4270 (N_4270,N_933,N_1384);
and U4271 (N_4271,N_547,N_363);
and U4272 (N_4272,N_1682,N_50);
xor U4273 (N_4273,N_2948,N_385);
and U4274 (N_4274,N_1214,N_2723);
or U4275 (N_4275,N_1071,N_1120);
or U4276 (N_4276,N_1262,N_2927);
nand U4277 (N_4277,N_86,N_1199);
nor U4278 (N_4278,N_1984,N_2060);
nor U4279 (N_4279,N_2433,N_483);
and U4280 (N_4280,N_1099,N_860);
nor U4281 (N_4281,N_1537,N_937);
nor U4282 (N_4282,N_340,N_1295);
or U4283 (N_4283,N_795,N_19);
xor U4284 (N_4284,N_2616,N_1954);
nor U4285 (N_4285,N_2116,N_259);
and U4286 (N_4286,N_1740,N_864);
nand U4287 (N_4287,N_1231,N_523);
xor U4288 (N_4288,N_220,N_219);
nor U4289 (N_4289,N_1787,N_2110);
or U4290 (N_4290,N_1916,N_1519);
nor U4291 (N_4291,N_1554,N_587);
or U4292 (N_4292,N_526,N_1147);
xor U4293 (N_4293,N_1580,N_375);
nor U4294 (N_4294,N_2818,N_1225);
nor U4295 (N_4295,N_255,N_2175);
nand U4296 (N_4296,N_2568,N_1053);
nor U4297 (N_4297,N_10,N_2070);
or U4298 (N_4298,N_841,N_307);
and U4299 (N_4299,N_1676,N_2109);
or U4300 (N_4300,N_2218,N_146);
xor U4301 (N_4301,N_2897,N_796);
nor U4302 (N_4302,N_1782,N_647);
or U4303 (N_4303,N_2535,N_348);
xor U4304 (N_4304,N_2585,N_2007);
nand U4305 (N_4305,N_892,N_2343);
nor U4306 (N_4306,N_965,N_292);
xnor U4307 (N_4307,N_2833,N_924);
nand U4308 (N_4308,N_763,N_1986);
nand U4309 (N_4309,N_672,N_45);
xnor U4310 (N_4310,N_2403,N_2186);
or U4311 (N_4311,N_2466,N_1239);
nor U4312 (N_4312,N_1277,N_2075);
nand U4313 (N_4313,N_1049,N_2347);
and U4314 (N_4314,N_635,N_1413);
nand U4315 (N_4315,N_539,N_481);
or U4316 (N_4316,N_1351,N_1853);
or U4317 (N_4317,N_310,N_1292);
or U4318 (N_4318,N_1727,N_1425);
xnor U4319 (N_4319,N_2148,N_1238);
and U4320 (N_4320,N_1968,N_2556);
xor U4321 (N_4321,N_2469,N_138);
or U4322 (N_4322,N_2293,N_1818);
nor U4323 (N_4323,N_2519,N_1680);
xnor U4324 (N_4324,N_2619,N_1902);
or U4325 (N_4325,N_1346,N_1034);
nor U4326 (N_4326,N_214,N_490);
nand U4327 (N_4327,N_2073,N_1795);
nand U4328 (N_4328,N_291,N_132);
or U4329 (N_4329,N_1930,N_2953);
and U4330 (N_4330,N_1216,N_26);
nor U4331 (N_4331,N_1775,N_1267);
or U4332 (N_4332,N_2301,N_1029);
xnor U4333 (N_4333,N_170,N_537);
xnor U4334 (N_4334,N_2150,N_920);
xor U4335 (N_4335,N_2162,N_2020);
xnor U4336 (N_4336,N_1838,N_1051);
xnor U4337 (N_4337,N_1124,N_1288);
nand U4338 (N_4338,N_627,N_2765);
and U4339 (N_4339,N_1209,N_1372);
xnor U4340 (N_4340,N_668,N_2138);
and U4341 (N_4341,N_2592,N_2798);
or U4342 (N_4342,N_277,N_608);
and U4343 (N_4343,N_1707,N_1828);
xor U4344 (N_4344,N_346,N_2787);
nor U4345 (N_4345,N_882,N_180);
nand U4346 (N_4346,N_2597,N_2859);
nor U4347 (N_4347,N_1538,N_1592);
nand U4348 (N_4348,N_2636,N_2170);
or U4349 (N_4349,N_1105,N_1060);
nand U4350 (N_4350,N_2010,N_683);
nor U4351 (N_4351,N_2280,N_67);
xor U4352 (N_4352,N_1011,N_109);
or U4353 (N_4353,N_1129,N_2703);
nor U4354 (N_4354,N_1759,N_825);
nor U4355 (N_4355,N_780,N_852);
and U4356 (N_4356,N_2815,N_1018);
and U4357 (N_4357,N_2632,N_2);
nand U4358 (N_4358,N_1959,N_2974);
nand U4359 (N_4359,N_1814,N_1293);
and U4360 (N_4360,N_1093,N_2474);
nand U4361 (N_4361,N_579,N_1342);
or U4362 (N_4362,N_1570,N_1556);
xor U4363 (N_4363,N_1382,N_2824);
and U4364 (N_4364,N_2024,N_1364);
nor U4365 (N_4365,N_696,N_989);
or U4366 (N_4366,N_79,N_2881);
or U4367 (N_4367,N_2139,N_1921);
or U4368 (N_4368,N_471,N_2049);
and U4369 (N_4369,N_676,N_925);
xnor U4370 (N_4370,N_2846,N_2957);
and U4371 (N_4371,N_1603,N_2149);
or U4372 (N_4372,N_2849,N_895);
xor U4373 (N_4373,N_2820,N_678);
or U4374 (N_4374,N_2498,N_2340);
xor U4375 (N_4375,N_386,N_69);
nand U4376 (N_4376,N_2067,N_834);
nand U4377 (N_4377,N_607,N_2225);
nand U4378 (N_4378,N_2348,N_887);
nand U4379 (N_4379,N_2638,N_723);
xor U4380 (N_4380,N_1546,N_2484);
nand U4381 (N_4381,N_113,N_2490);
and U4382 (N_4382,N_600,N_337);
nand U4383 (N_4383,N_1283,N_1141);
and U4384 (N_4384,N_1571,N_2670);
xnor U4385 (N_4385,N_1366,N_2091);
and U4386 (N_4386,N_1730,N_2607);
xor U4387 (N_4387,N_1753,N_384);
and U4388 (N_4388,N_504,N_830);
or U4389 (N_4389,N_596,N_1083);
xnor U4390 (N_4390,N_1151,N_1507);
xor U4391 (N_4391,N_880,N_1329);
nor U4392 (N_4392,N_2772,N_2252);
xor U4393 (N_4393,N_204,N_793);
xnor U4394 (N_4394,N_817,N_1399);
nand U4395 (N_4395,N_1641,N_1403);
or U4396 (N_4396,N_1635,N_369);
and U4397 (N_4397,N_1646,N_1352);
nand U4398 (N_4398,N_1499,N_1158);
nand U4399 (N_4399,N_61,N_148);
nand U4400 (N_4400,N_1078,N_1955);
xor U4401 (N_4401,N_1361,N_2428);
and U4402 (N_4402,N_1469,N_40);
nand U4403 (N_4403,N_553,N_2066);
xnor U4404 (N_4404,N_2421,N_1486);
xor U4405 (N_4405,N_1131,N_429);
xnor U4406 (N_4406,N_2318,N_2353);
nand U4407 (N_4407,N_2245,N_1313);
and U4408 (N_4408,N_2629,N_1988);
nor U4409 (N_4409,N_1164,N_1644);
or U4410 (N_4410,N_2102,N_2501);
nor U4411 (N_4411,N_2137,N_304);
or U4412 (N_4412,N_2984,N_327);
and U4413 (N_4413,N_1316,N_2480);
nand U4414 (N_4414,N_2083,N_1824);
and U4415 (N_4415,N_812,N_2848);
nor U4416 (N_4416,N_274,N_2399);
nor U4417 (N_4417,N_2183,N_1452);
or U4418 (N_4418,N_2570,N_282);
or U4419 (N_4419,N_1783,N_1390);
and U4420 (N_4420,N_591,N_2364);
nor U4421 (N_4421,N_2749,N_1036);
nor U4422 (N_4422,N_535,N_280);
nor U4423 (N_4423,N_2688,N_2972);
nor U4424 (N_4424,N_28,N_2865);
and U4425 (N_4425,N_2171,N_2679);
xnor U4426 (N_4426,N_851,N_2385);
nor U4427 (N_4427,N_2028,N_1896);
and U4428 (N_4428,N_1941,N_2901);
nand U4429 (N_4429,N_1512,N_1369);
and U4430 (N_4430,N_226,N_150);
or U4431 (N_4431,N_1714,N_1465);
nand U4432 (N_4432,N_1166,N_1155);
or U4433 (N_4433,N_703,N_2834);
nand U4434 (N_4434,N_389,N_650);
and U4435 (N_4435,N_63,N_2821);
nand U4436 (N_4436,N_32,N_1086);
nor U4437 (N_4437,N_1460,N_103);
nand U4438 (N_4438,N_2563,N_590);
nor U4439 (N_4439,N_2683,N_2666);
xor U4440 (N_4440,N_964,N_1330);
xor U4441 (N_4441,N_1652,N_1513);
or U4442 (N_4442,N_2500,N_1064);
nor U4443 (N_4443,N_489,N_264);
nand U4444 (N_4444,N_995,N_1999);
and U4445 (N_4445,N_2871,N_2855);
or U4446 (N_4446,N_963,N_651);
nor U4447 (N_4447,N_200,N_1428);
nor U4448 (N_4448,N_2884,N_2033);
nand U4449 (N_4449,N_736,N_379);
and U4450 (N_4450,N_926,N_2380);
nor U4451 (N_4451,N_253,N_529);
nand U4452 (N_4452,N_721,N_601);
or U4453 (N_4453,N_454,N_196);
nor U4454 (N_4454,N_2628,N_51);
nand U4455 (N_4455,N_445,N_2742);
nand U4456 (N_4456,N_1297,N_1280);
xor U4457 (N_4457,N_2624,N_533);
nor U4458 (N_4458,N_355,N_1812);
nand U4459 (N_4459,N_2806,N_2564);
and U4460 (N_4460,N_2317,N_1788);
and U4461 (N_4461,N_1744,N_1901);
nand U4462 (N_4462,N_2705,N_2875);
xnor U4463 (N_4463,N_1467,N_811);
xnor U4464 (N_4464,N_1587,N_2420);
xnor U4465 (N_4465,N_2936,N_1464);
xnor U4466 (N_4466,N_957,N_2410);
nor U4467 (N_4467,N_2534,N_665);
or U4468 (N_4468,N_2371,N_514);
nor U4469 (N_4469,N_1904,N_546);
and U4470 (N_4470,N_1758,N_1296);
and U4471 (N_4471,N_1311,N_2135);
and U4472 (N_4472,N_1749,N_2627);
nor U4473 (N_4473,N_1322,N_1008);
xor U4474 (N_4474,N_2533,N_1575);
nand U4475 (N_4475,N_2023,N_1150);
nor U4476 (N_4476,N_2100,N_2889);
nand U4477 (N_4477,N_1119,N_1937);
xor U4478 (N_4478,N_1560,N_2376);
nand U4479 (N_4479,N_799,N_413);
xnor U4480 (N_4480,N_446,N_1504);
or U4481 (N_4481,N_1009,N_725);
or U4482 (N_4482,N_1559,N_2434);
xor U4483 (N_4483,N_1557,N_2115);
nand U4484 (N_4484,N_2733,N_221);
nand U4485 (N_4485,N_1657,N_1367);
or U4486 (N_4486,N_1883,N_1724);
nor U4487 (N_4487,N_350,N_542);
nand U4488 (N_4488,N_1748,N_1878);
nand U4489 (N_4489,N_2914,N_2509);
nand U4490 (N_4490,N_1626,N_2898);
or U4491 (N_4491,N_674,N_661);
or U4492 (N_4492,N_524,N_2667);
or U4493 (N_4493,N_2454,N_1677);
nor U4494 (N_4494,N_771,N_2902);
nand U4495 (N_4495,N_1472,N_1002);
or U4496 (N_4496,N_312,N_2228);
and U4497 (N_4497,N_960,N_1142);
xnor U4498 (N_4498,N_802,N_2470);
or U4499 (N_4499,N_1459,N_1914);
nor U4500 (N_4500,N_363,N_2371);
nor U4501 (N_4501,N_1668,N_1430);
and U4502 (N_4502,N_2343,N_1473);
and U4503 (N_4503,N_2793,N_2682);
or U4504 (N_4504,N_779,N_1047);
nor U4505 (N_4505,N_2906,N_1346);
xor U4506 (N_4506,N_2564,N_2639);
or U4507 (N_4507,N_1874,N_183);
nand U4508 (N_4508,N_2918,N_1766);
or U4509 (N_4509,N_1633,N_2603);
xnor U4510 (N_4510,N_1601,N_265);
and U4511 (N_4511,N_363,N_2757);
nor U4512 (N_4512,N_102,N_1160);
or U4513 (N_4513,N_1439,N_643);
or U4514 (N_4514,N_124,N_959);
and U4515 (N_4515,N_2056,N_2129);
or U4516 (N_4516,N_1264,N_1927);
and U4517 (N_4517,N_2662,N_1520);
xnor U4518 (N_4518,N_1225,N_2560);
or U4519 (N_4519,N_2450,N_163);
xor U4520 (N_4520,N_190,N_2050);
nor U4521 (N_4521,N_2618,N_432);
nand U4522 (N_4522,N_207,N_1230);
and U4523 (N_4523,N_163,N_119);
nand U4524 (N_4524,N_2860,N_2017);
nand U4525 (N_4525,N_2531,N_1875);
xor U4526 (N_4526,N_669,N_1964);
nand U4527 (N_4527,N_1209,N_2041);
and U4528 (N_4528,N_1465,N_129);
nand U4529 (N_4529,N_623,N_1908);
and U4530 (N_4530,N_1597,N_2455);
nand U4531 (N_4531,N_424,N_1829);
nor U4532 (N_4532,N_1016,N_1814);
nand U4533 (N_4533,N_1831,N_2160);
xnor U4534 (N_4534,N_2485,N_1508);
nor U4535 (N_4535,N_103,N_100);
nor U4536 (N_4536,N_2455,N_381);
and U4537 (N_4537,N_858,N_259);
or U4538 (N_4538,N_1825,N_1108);
xor U4539 (N_4539,N_2816,N_2902);
or U4540 (N_4540,N_1012,N_1617);
and U4541 (N_4541,N_1093,N_460);
nand U4542 (N_4542,N_2730,N_1245);
xor U4543 (N_4543,N_715,N_1802);
xor U4544 (N_4544,N_1793,N_2008);
nand U4545 (N_4545,N_1796,N_399);
and U4546 (N_4546,N_1106,N_770);
nand U4547 (N_4547,N_2051,N_2698);
and U4548 (N_4548,N_358,N_1820);
and U4549 (N_4549,N_1039,N_1088);
nand U4550 (N_4550,N_1719,N_1234);
and U4551 (N_4551,N_2989,N_2740);
nand U4552 (N_4552,N_2856,N_811);
nor U4553 (N_4553,N_2765,N_578);
xnor U4554 (N_4554,N_628,N_2005);
or U4555 (N_4555,N_1071,N_1708);
nor U4556 (N_4556,N_281,N_2020);
and U4557 (N_4557,N_905,N_1817);
or U4558 (N_4558,N_756,N_1791);
xnor U4559 (N_4559,N_585,N_1696);
and U4560 (N_4560,N_2143,N_1347);
and U4561 (N_4561,N_585,N_607);
nor U4562 (N_4562,N_1616,N_2474);
nor U4563 (N_4563,N_664,N_2330);
and U4564 (N_4564,N_2185,N_390);
xor U4565 (N_4565,N_2816,N_267);
or U4566 (N_4566,N_2427,N_2807);
nor U4567 (N_4567,N_2403,N_2214);
nand U4568 (N_4568,N_55,N_2243);
and U4569 (N_4569,N_1515,N_973);
nor U4570 (N_4570,N_1573,N_458);
or U4571 (N_4571,N_1527,N_2998);
or U4572 (N_4572,N_91,N_1892);
nand U4573 (N_4573,N_370,N_2685);
nor U4574 (N_4574,N_1808,N_2069);
nand U4575 (N_4575,N_746,N_1117);
or U4576 (N_4576,N_2583,N_126);
and U4577 (N_4577,N_823,N_833);
and U4578 (N_4578,N_2950,N_75);
and U4579 (N_4579,N_2421,N_104);
and U4580 (N_4580,N_2006,N_2504);
nand U4581 (N_4581,N_1488,N_720);
xor U4582 (N_4582,N_1664,N_2108);
nor U4583 (N_4583,N_2320,N_2801);
and U4584 (N_4584,N_262,N_442);
nand U4585 (N_4585,N_2347,N_716);
or U4586 (N_4586,N_1181,N_531);
xor U4587 (N_4587,N_2292,N_194);
and U4588 (N_4588,N_2830,N_878);
nor U4589 (N_4589,N_2054,N_63);
xor U4590 (N_4590,N_30,N_1287);
nor U4591 (N_4591,N_173,N_2860);
and U4592 (N_4592,N_483,N_1090);
nand U4593 (N_4593,N_1762,N_1639);
xnor U4594 (N_4594,N_1541,N_696);
and U4595 (N_4595,N_940,N_911);
or U4596 (N_4596,N_606,N_977);
nor U4597 (N_4597,N_2042,N_2957);
nand U4598 (N_4598,N_2232,N_2781);
nand U4599 (N_4599,N_1144,N_289);
xnor U4600 (N_4600,N_1777,N_90);
nor U4601 (N_4601,N_788,N_142);
xnor U4602 (N_4602,N_535,N_2087);
nand U4603 (N_4603,N_1306,N_2119);
xor U4604 (N_4604,N_1712,N_1966);
nand U4605 (N_4605,N_533,N_2429);
and U4606 (N_4606,N_2749,N_1734);
nand U4607 (N_4607,N_2772,N_2702);
xor U4608 (N_4608,N_1774,N_2012);
xnor U4609 (N_4609,N_2739,N_2096);
nand U4610 (N_4610,N_2883,N_1347);
nor U4611 (N_4611,N_1146,N_2121);
nor U4612 (N_4612,N_2285,N_1944);
nor U4613 (N_4613,N_1363,N_555);
and U4614 (N_4614,N_1191,N_659);
or U4615 (N_4615,N_478,N_1833);
xnor U4616 (N_4616,N_851,N_1761);
or U4617 (N_4617,N_1060,N_2239);
or U4618 (N_4618,N_1996,N_99);
xnor U4619 (N_4619,N_2930,N_2230);
xnor U4620 (N_4620,N_2568,N_63);
nand U4621 (N_4621,N_1195,N_520);
nand U4622 (N_4622,N_1322,N_588);
xnor U4623 (N_4623,N_269,N_1848);
or U4624 (N_4624,N_2956,N_928);
nand U4625 (N_4625,N_2364,N_1145);
and U4626 (N_4626,N_841,N_788);
nor U4627 (N_4627,N_2204,N_501);
nor U4628 (N_4628,N_1068,N_1783);
nand U4629 (N_4629,N_124,N_2715);
nor U4630 (N_4630,N_1666,N_663);
nand U4631 (N_4631,N_1322,N_2920);
and U4632 (N_4632,N_1444,N_1747);
and U4633 (N_4633,N_884,N_2624);
nor U4634 (N_4634,N_2797,N_730);
nand U4635 (N_4635,N_709,N_466);
xnor U4636 (N_4636,N_945,N_2885);
or U4637 (N_4637,N_496,N_2995);
xor U4638 (N_4638,N_771,N_138);
or U4639 (N_4639,N_2840,N_1581);
or U4640 (N_4640,N_1658,N_1398);
xnor U4641 (N_4641,N_1454,N_953);
nor U4642 (N_4642,N_1257,N_2167);
or U4643 (N_4643,N_432,N_2480);
and U4644 (N_4644,N_2735,N_243);
nor U4645 (N_4645,N_2572,N_1504);
nor U4646 (N_4646,N_1006,N_1169);
nand U4647 (N_4647,N_323,N_1472);
nor U4648 (N_4648,N_172,N_2047);
and U4649 (N_4649,N_2759,N_241);
nor U4650 (N_4650,N_671,N_2694);
nand U4651 (N_4651,N_157,N_876);
nor U4652 (N_4652,N_2056,N_708);
nor U4653 (N_4653,N_1018,N_2846);
xor U4654 (N_4654,N_1332,N_2688);
nor U4655 (N_4655,N_1312,N_1415);
nand U4656 (N_4656,N_1834,N_1515);
nor U4657 (N_4657,N_2524,N_2129);
nand U4658 (N_4658,N_1806,N_1943);
nand U4659 (N_4659,N_659,N_1334);
nand U4660 (N_4660,N_1956,N_2919);
or U4661 (N_4661,N_1127,N_2914);
and U4662 (N_4662,N_2985,N_353);
nor U4663 (N_4663,N_10,N_351);
or U4664 (N_4664,N_847,N_108);
and U4665 (N_4665,N_2982,N_1481);
and U4666 (N_4666,N_1408,N_708);
nand U4667 (N_4667,N_342,N_1924);
or U4668 (N_4668,N_69,N_230);
nand U4669 (N_4669,N_1160,N_2297);
xnor U4670 (N_4670,N_2004,N_2520);
nor U4671 (N_4671,N_2067,N_2663);
xor U4672 (N_4672,N_1872,N_2959);
xor U4673 (N_4673,N_377,N_2072);
xor U4674 (N_4674,N_2385,N_1884);
nor U4675 (N_4675,N_104,N_600);
nand U4676 (N_4676,N_33,N_2031);
nor U4677 (N_4677,N_1777,N_2651);
nand U4678 (N_4678,N_804,N_1612);
xor U4679 (N_4679,N_2688,N_1799);
and U4680 (N_4680,N_1395,N_1432);
or U4681 (N_4681,N_406,N_876);
and U4682 (N_4682,N_1948,N_2995);
or U4683 (N_4683,N_567,N_2859);
nor U4684 (N_4684,N_1984,N_2738);
nand U4685 (N_4685,N_2376,N_2322);
and U4686 (N_4686,N_1674,N_2996);
or U4687 (N_4687,N_16,N_117);
and U4688 (N_4688,N_521,N_238);
nor U4689 (N_4689,N_1352,N_89);
xor U4690 (N_4690,N_2945,N_395);
or U4691 (N_4691,N_57,N_1801);
and U4692 (N_4692,N_1749,N_2419);
nor U4693 (N_4693,N_1829,N_627);
nor U4694 (N_4694,N_1622,N_945);
xor U4695 (N_4695,N_229,N_2613);
xor U4696 (N_4696,N_2713,N_2404);
nor U4697 (N_4697,N_2366,N_571);
or U4698 (N_4698,N_1132,N_1419);
nor U4699 (N_4699,N_2080,N_2128);
xnor U4700 (N_4700,N_2070,N_2343);
xnor U4701 (N_4701,N_352,N_849);
nor U4702 (N_4702,N_1637,N_2572);
nor U4703 (N_4703,N_1346,N_1699);
nand U4704 (N_4704,N_1184,N_1836);
xor U4705 (N_4705,N_305,N_1019);
and U4706 (N_4706,N_596,N_2643);
xor U4707 (N_4707,N_1742,N_535);
nor U4708 (N_4708,N_2318,N_1398);
nor U4709 (N_4709,N_675,N_27);
or U4710 (N_4710,N_410,N_2891);
nor U4711 (N_4711,N_40,N_1184);
or U4712 (N_4712,N_2354,N_2426);
or U4713 (N_4713,N_1466,N_702);
nor U4714 (N_4714,N_169,N_650);
nor U4715 (N_4715,N_295,N_529);
xnor U4716 (N_4716,N_111,N_2407);
and U4717 (N_4717,N_2778,N_660);
xor U4718 (N_4718,N_845,N_2017);
and U4719 (N_4719,N_2450,N_148);
and U4720 (N_4720,N_901,N_1449);
nor U4721 (N_4721,N_2229,N_555);
or U4722 (N_4722,N_2330,N_1997);
nor U4723 (N_4723,N_1557,N_257);
or U4724 (N_4724,N_282,N_2412);
nor U4725 (N_4725,N_2431,N_2239);
nand U4726 (N_4726,N_146,N_1064);
and U4727 (N_4727,N_945,N_544);
xnor U4728 (N_4728,N_2815,N_1377);
nand U4729 (N_4729,N_860,N_810);
nor U4730 (N_4730,N_919,N_1353);
or U4731 (N_4731,N_712,N_2452);
xor U4732 (N_4732,N_1747,N_1555);
nor U4733 (N_4733,N_0,N_1287);
xor U4734 (N_4734,N_1440,N_2075);
and U4735 (N_4735,N_2207,N_2473);
xor U4736 (N_4736,N_1266,N_391);
nand U4737 (N_4737,N_2984,N_2729);
xor U4738 (N_4738,N_2372,N_2412);
or U4739 (N_4739,N_1709,N_188);
xnor U4740 (N_4740,N_2522,N_1866);
nor U4741 (N_4741,N_1697,N_1761);
and U4742 (N_4742,N_386,N_1619);
xnor U4743 (N_4743,N_2488,N_2037);
nand U4744 (N_4744,N_1095,N_628);
nand U4745 (N_4745,N_1758,N_2678);
xor U4746 (N_4746,N_854,N_2461);
or U4747 (N_4747,N_1486,N_2971);
or U4748 (N_4748,N_1310,N_1790);
xor U4749 (N_4749,N_2011,N_1215);
xnor U4750 (N_4750,N_673,N_1217);
and U4751 (N_4751,N_2314,N_1423);
or U4752 (N_4752,N_1899,N_2601);
and U4753 (N_4753,N_1936,N_2441);
nor U4754 (N_4754,N_472,N_176);
nand U4755 (N_4755,N_182,N_1863);
nor U4756 (N_4756,N_619,N_1217);
xnor U4757 (N_4757,N_392,N_257);
nand U4758 (N_4758,N_182,N_1299);
nor U4759 (N_4759,N_1777,N_157);
or U4760 (N_4760,N_1776,N_2420);
nor U4761 (N_4761,N_919,N_1338);
nor U4762 (N_4762,N_493,N_2596);
nand U4763 (N_4763,N_982,N_2520);
xor U4764 (N_4764,N_2946,N_86);
xnor U4765 (N_4765,N_2258,N_2268);
xor U4766 (N_4766,N_591,N_683);
and U4767 (N_4767,N_2568,N_2522);
or U4768 (N_4768,N_597,N_1191);
nand U4769 (N_4769,N_1876,N_1797);
nor U4770 (N_4770,N_2485,N_2140);
nor U4771 (N_4771,N_1373,N_2977);
xnor U4772 (N_4772,N_2669,N_906);
nor U4773 (N_4773,N_210,N_2165);
nand U4774 (N_4774,N_2651,N_336);
or U4775 (N_4775,N_696,N_137);
nand U4776 (N_4776,N_1197,N_2563);
or U4777 (N_4777,N_739,N_2467);
and U4778 (N_4778,N_769,N_1486);
and U4779 (N_4779,N_2768,N_465);
nor U4780 (N_4780,N_1162,N_98);
xnor U4781 (N_4781,N_994,N_2522);
nand U4782 (N_4782,N_1956,N_2350);
and U4783 (N_4783,N_6,N_964);
nor U4784 (N_4784,N_1937,N_373);
nand U4785 (N_4785,N_768,N_710);
and U4786 (N_4786,N_2127,N_92);
nand U4787 (N_4787,N_968,N_1587);
nor U4788 (N_4788,N_2593,N_725);
or U4789 (N_4789,N_591,N_1630);
nor U4790 (N_4790,N_627,N_541);
xnor U4791 (N_4791,N_490,N_2140);
nand U4792 (N_4792,N_2964,N_2645);
nand U4793 (N_4793,N_1015,N_2947);
xor U4794 (N_4794,N_1669,N_2166);
nor U4795 (N_4795,N_1097,N_2460);
nand U4796 (N_4796,N_1400,N_1131);
xor U4797 (N_4797,N_1053,N_2782);
nand U4798 (N_4798,N_750,N_791);
and U4799 (N_4799,N_667,N_551);
and U4800 (N_4800,N_2918,N_2557);
nand U4801 (N_4801,N_142,N_2821);
and U4802 (N_4802,N_61,N_965);
nor U4803 (N_4803,N_2406,N_528);
nor U4804 (N_4804,N_2684,N_873);
xnor U4805 (N_4805,N_1678,N_471);
nand U4806 (N_4806,N_1007,N_1834);
nand U4807 (N_4807,N_609,N_1472);
or U4808 (N_4808,N_1532,N_2381);
or U4809 (N_4809,N_1259,N_947);
nand U4810 (N_4810,N_1230,N_880);
xnor U4811 (N_4811,N_1019,N_1768);
nand U4812 (N_4812,N_43,N_2641);
and U4813 (N_4813,N_1436,N_127);
nor U4814 (N_4814,N_483,N_1474);
xor U4815 (N_4815,N_791,N_1410);
and U4816 (N_4816,N_859,N_2185);
nor U4817 (N_4817,N_2903,N_644);
nand U4818 (N_4818,N_1323,N_1180);
nand U4819 (N_4819,N_851,N_1930);
xor U4820 (N_4820,N_632,N_1954);
nand U4821 (N_4821,N_513,N_1);
nand U4822 (N_4822,N_2144,N_1533);
nor U4823 (N_4823,N_1536,N_2139);
nor U4824 (N_4824,N_1171,N_662);
xor U4825 (N_4825,N_2504,N_534);
nor U4826 (N_4826,N_2393,N_167);
or U4827 (N_4827,N_1166,N_1250);
or U4828 (N_4828,N_866,N_1721);
or U4829 (N_4829,N_645,N_1489);
nand U4830 (N_4830,N_900,N_2381);
xnor U4831 (N_4831,N_375,N_169);
xor U4832 (N_4832,N_1646,N_423);
nor U4833 (N_4833,N_1354,N_868);
or U4834 (N_4834,N_1935,N_2788);
or U4835 (N_4835,N_2239,N_1479);
and U4836 (N_4836,N_2844,N_1702);
or U4837 (N_4837,N_212,N_347);
or U4838 (N_4838,N_1426,N_361);
nor U4839 (N_4839,N_810,N_1803);
nand U4840 (N_4840,N_2799,N_960);
or U4841 (N_4841,N_2109,N_1262);
or U4842 (N_4842,N_388,N_2108);
nor U4843 (N_4843,N_1713,N_2864);
or U4844 (N_4844,N_487,N_1011);
nor U4845 (N_4845,N_1215,N_541);
or U4846 (N_4846,N_1101,N_955);
nor U4847 (N_4847,N_1799,N_248);
nand U4848 (N_4848,N_757,N_1316);
xnor U4849 (N_4849,N_2737,N_2600);
or U4850 (N_4850,N_614,N_915);
nand U4851 (N_4851,N_713,N_1972);
nand U4852 (N_4852,N_405,N_772);
or U4853 (N_4853,N_2190,N_2396);
nand U4854 (N_4854,N_2443,N_1951);
and U4855 (N_4855,N_2875,N_1425);
xor U4856 (N_4856,N_2051,N_65);
and U4857 (N_4857,N_1244,N_2882);
nor U4858 (N_4858,N_458,N_2927);
and U4859 (N_4859,N_1889,N_2564);
xor U4860 (N_4860,N_2109,N_2073);
nor U4861 (N_4861,N_2217,N_2296);
and U4862 (N_4862,N_2185,N_2858);
nor U4863 (N_4863,N_818,N_2240);
xor U4864 (N_4864,N_1774,N_2908);
and U4865 (N_4865,N_976,N_1733);
nor U4866 (N_4866,N_1279,N_152);
nand U4867 (N_4867,N_2699,N_1355);
or U4868 (N_4868,N_2866,N_2463);
nand U4869 (N_4869,N_2743,N_2296);
xor U4870 (N_4870,N_1692,N_1710);
xor U4871 (N_4871,N_2696,N_1935);
xor U4872 (N_4872,N_1563,N_1871);
xor U4873 (N_4873,N_1942,N_919);
and U4874 (N_4874,N_1010,N_1327);
or U4875 (N_4875,N_592,N_490);
xnor U4876 (N_4876,N_146,N_2298);
nor U4877 (N_4877,N_2941,N_425);
nor U4878 (N_4878,N_2361,N_2364);
and U4879 (N_4879,N_1702,N_1767);
nand U4880 (N_4880,N_2187,N_1994);
nand U4881 (N_4881,N_1977,N_2091);
nor U4882 (N_4882,N_2045,N_2644);
xnor U4883 (N_4883,N_2067,N_2668);
and U4884 (N_4884,N_610,N_2305);
and U4885 (N_4885,N_1682,N_645);
nand U4886 (N_4886,N_1400,N_1516);
nor U4887 (N_4887,N_1188,N_2968);
nor U4888 (N_4888,N_397,N_899);
nor U4889 (N_4889,N_2345,N_1312);
or U4890 (N_4890,N_2658,N_1211);
nand U4891 (N_4891,N_2435,N_2707);
or U4892 (N_4892,N_2871,N_1394);
and U4893 (N_4893,N_2275,N_67);
xor U4894 (N_4894,N_2979,N_136);
xnor U4895 (N_4895,N_358,N_1389);
xnor U4896 (N_4896,N_411,N_651);
and U4897 (N_4897,N_606,N_2382);
nand U4898 (N_4898,N_704,N_2496);
nor U4899 (N_4899,N_194,N_831);
or U4900 (N_4900,N_1747,N_1752);
or U4901 (N_4901,N_2437,N_2685);
nor U4902 (N_4902,N_1879,N_1171);
nor U4903 (N_4903,N_1186,N_950);
and U4904 (N_4904,N_2353,N_716);
xnor U4905 (N_4905,N_1074,N_206);
nand U4906 (N_4906,N_372,N_33);
nand U4907 (N_4907,N_1714,N_339);
nand U4908 (N_4908,N_2366,N_2086);
xor U4909 (N_4909,N_1624,N_1413);
xor U4910 (N_4910,N_1244,N_1400);
nor U4911 (N_4911,N_2384,N_530);
nand U4912 (N_4912,N_1734,N_2);
xor U4913 (N_4913,N_601,N_1990);
nand U4914 (N_4914,N_1232,N_156);
or U4915 (N_4915,N_1186,N_1413);
nand U4916 (N_4916,N_1512,N_1764);
and U4917 (N_4917,N_735,N_1446);
xor U4918 (N_4918,N_1026,N_2640);
nor U4919 (N_4919,N_1102,N_2703);
nor U4920 (N_4920,N_663,N_1869);
and U4921 (N_4921,N_2096,N_691);
or U4922 (N_4922,N_918,N_31);
and U4923 (N_4923,N_1133,N_33);
or U4924 (N_4924,N_2631,N_2420);
or U4925 (N_4925,N_2556,N_2146);
or U4926 (N_4926,N_2083,N_2951);
nor U4927 (N_4927,N_418,N_1285);
xor U4928 (N_4928,N_1130,N_866);
xor U4929 (N_4929,N_1134,N_1537);
xnor U4930 (N_4930,N_1742,N_116);
nand U4931 (N_4931,N_2900,N_170);
nor U4932 (N_4932,N_513,N_2167);
or U4933 (N_4933,N_2150,N_1599);
nor U4934 (N_4934,N_2331,N_1704);
nor U4935 (N_4935,N_1482,N_16);
and U4936 (N_4936,N_1533,N_2776);
or U4937 (N_4937,N_1675,N_533);
nand U4938 (N_4938,N_1159,N_910);
or U4939 (N_4939,N_1671,N_963);
or U4940 (N_4940,N_52,N_231);
or U4941 (N_4941,N_1733,N_743);
nand U4942 (N_4942,N_1047,N_2068);
nand U4943 (N_4943,N_1278,N_638);
xnor U4944 (N_4944,N_1009,N_1611);
nand U4945 (N_4945,N_1089,N_1883);
or U4946 (N_4946,N_103,N_2304);
and U4947 (N_4947,N_1414,N_2364);
nand U4948 (N_4948,N_1294,N_2966);
and U4949 (N_4949,N_1540,N_505);
nand U4950 (N_4950,N_2521,N_1670);
nand U4951 (N_4951,N_1621,N_668);
nor U4952 (N_4952,N_614,N_1310);
nand U4953 (N_4953,N_1524,N_1147);
and U4954 (N_4954,N_1550,N_2168);
and U4955 (N_4955,N_2781,N_901);
or U4956 (N_4956,N_2813,N_2325);
nor U4957 (N_4957,N_1791,N_1021);
nand U4958 (N_4958,N_981,N_809);
and U4959 (N_4959,N_853,N_1411);
and U4960 (N_4960,N_416,N_2822);
xor U4961 (N_4961,N_1437,N_1345);
and U4962 (N_4962,N_2886,N_1406);
and U4963 (N_4963,N_785,N_2334);
xor U4964 (N_4964,N_1069,N_1924);
nor U4965 (N_4965,N_2399,N_272);
xnor U4966 (N_4966,N_1456,N_26);
nor U4967 (N_4967,N_2390,N_2068);
xor U4968 (N_4968,N_2957,N_2839);
nand U4969 (N_4969,N_1624,N_1197);
or U4970 (N_4970,N_23,N_171);
and U4971 (N_4971,N_1185,N_1829);
nand U4972 (N_4972,N_2422,N_2442);
xnor U4973 (N_4973,N_2356,N_739);
nand U4974 (N_4974,N_2394,N_348);
nor U4975 (N_4975,N_451,N_1805);
nor U4976 (N_4976,N_809,N_1092);
and U4977 (N_4977,N_1531,N_583);
and U4978 (N_4978,N_2870,N_540);
xor U4979 (N_4979,N_2151,N_2931);
or U4980 (N_4980,N_184,N_1334);
or U4981 (N_4981,N_230,N_559);
xor U4982 (N_4982,N_2922,N_2496);
nand U4983 (N_4983,N_855,N_199);
nor U4984 (N_4984,N_131,N_67);
nand U4985 (N_4985,N_1019,N_2321);
nor U4986 (N_4986,N_2163,N_78);
xor U4987 (N_4987,N_685,N_1094);
or U4988 (N_4988,N_2119,N_2943);
nor U4989 (N_4989,N_838,N_2829);
nand U4990 (N_4990,N_556,N_1143);
or U4991 (N_4991,N_657,N_301);
nor U4992 (N_4992,N_1486,N_1528);
nand U4993 (N_4993,N_852,N_114);
or U4994 (N_4994,N_1177,N_2591);
and U4995 (N_4995,N_1164,N_2711);
xor U4996 (N_4996,N_2973,N_696);
nor U4997 (N_4997,N_1852,N_1679);
and U4998 (N_4998,N_2314,N_1570);
nand U4999 (N_4999,N_476,N_2444);
or U5000 (N_5000,N_1084,N_2238);
xor U5001 (N_5001,N_2073,N_592);
nor U5002 (N_5002,N_745,N_1505);
or U5003 (N_5003,N_60,N_2242);
and U5004 (N_5004,N_2455,N_316);
and U5005 (N_5005,N_957,N_1860);
and U5006 (N_5006,N_1788,N_1865);
or U5007 (N_5007,N_1712,N_1155);
or U5008 (N_5008,N_1536,N_966);
nand U5009 (N_5009,N_2021,N_72);
xnor U5010 (N_5010,N_37,N_2126);
xnor U5011 (N_5011,N_966,N_2954);
or U5012 (N_5012,N_1271,N_1809);
nand U5013 (N_5013,N_1320,N_614);
nor U5014 (N_5014,N_1524,N_2901);
or U5015 (N_5015,N_2564,N_1830);
or U5016 (N_5016,N_296,N_2951);
or U5017 (N_5017,N_738,N_2037);
nor U5018 (N_5018,N_528,N_363);
and U5019 (N_5019,N_107,N_2517);
xnor U5020 (N_5020,N_1256,N_1644);
nand U5021 (N_5021,N_681,N_708);
or U5022 (N_5022,N_2892,N_779);
nand U5023 (N_5023,N_2812,N_949);
or U5024 (N_5024,N_2991,N_93);
and U5025 (N_5025,N_1571,N_1028);
nand U5026 (N_5026,N_2670,N_1463);
nor U5027 (N_5027,N_2151,N_2257);
xor U5028 (N_5028,N_335,N_1333);
xnor U5029 (N_5029,N_663,N_1308);
xnor U5030 (N_5030,N_55,N_125);
or U5031 (N_5031,N_690,N_213);
nand U5032 (N_5032,N_2822,N_290);
nor U5033 (N_5033,N_2089,N_2383);
nor U5034 (N_5034,N_2710,N_70);
nor U5035 (N_5035,N_1694,N_1051);
xnor U5036 (N_5036,N_1934,N_852);
nand U5037 (N_5037,N_1155,N_2031);
nand U5038 (N_5038,N_215,N_172);
nand U5039 (N_5039,N_1915,N_2223);
nand U5040 (N_5040,N_478,N_2161);
and U5041 (N_5041,N_357,N_1263);
nor U5042 (N_5042,N_615,N_2478);
or U5043 (N_5043,N_620,N_2188);
xor U5044 (N_5044,N_2980,N_2143);
and U5045 (N_5045,N_2490,N_1247);
nor U5046 (N_5046,N_994,N_2609);
nor U5047 (N_5047,N_2278,N_1289);
and U5048 (N_5048,N_1611,N_1189);
or U5049 (N_5049,N_195,N_2066);
or U5050 (N_5050,N_768,N_2136);
nand U5051 (N_5051,N_1881,N_894);
xor U5052 (N_5052,N_2502,N_995);
nor U5053 (N_5053,N_1632,N_2698);
or U5054 (N_5054,N_2563,N_2708);
xor U5055 (N_5055,N_2403,N_1008);
or U5056 (N_5056,N_815,N_1475);
or U5057 (N_5057,N_2306,N_1010);
nor U5058 (N_5058,N_2667,N_2535);
or U5059 (N_5059,N_662,N_1067);
nor U5060 (N_5060,N_2217,N_2078);
and U5061 (N_5061,N_691,N_1153);
xor U5062 (N_5062,N_395,N_1914);
nand U5063 (N_5063,N_1535,N_1801);
nor U5064 (N_5064,N_78,N_479);
or U5065 (N_5065,N_1247,N_1367);
xnor U5066 (N_5066,N_2306,N_2921);
and U5067 (N_5067,N_2416,N_206);
or U5068 (N_5068,N_2336,N_375);
nand U5069 (N_5069,N_2640,N_1886);
xor U5070 (N_5070,N_2995,N_2401);
xnor U5071 (N_5071,N_899,N_2220);
and U5072 (N_5072,N_966,N_1187);
nand U5073 (N_5073,N_1198,N_1136);
nand U5074 (N_5074,N_1938,N_1763);
nand U5075 (N_5075,N_2961,N_1435);
and U5076 (N_5076,N_2928,N_1745);
nor U5077 (N_5077,N_1212,N_1114);
or U5078 (N_5078,N_1580,N_1144);
or U5079 (N_5079,N_100,N_109);
nor U5080 (N_5080,N_1845,N_1987);
or U5081 (N_5081,N_158,N_2256);
or U5082 (N_5082,N_192,N_1958);
nand U5083 (N_5083,N_2152,N_1742);
nand U5084 (N_5084,N_456,N_2943);
and U5085 (N_5085,N_2279,N_2501);
nor U5086 (N_5086,N_2700,N_399);
xnor U5087 (N_5087,N_2856,N_2019);
nor U5088 (N_5088,N_2012,N_1292);
nor U5089 (N_5089,N_2910,N_208);
and U5090 (N_5090,N_1092,N_1734);
xor U5091 (N_5091,N_1147,N_868);
xnor U5092 (N_5092,N_2719,N_428);
nor U5093 (N_5093,N_2240,N_2000);
nor U5094 (N_5094,N_1224,N_1201);
or U5095 (N_5095,N_622,N_2358);
or U5096 (N_5096,N_104,N_1358);
xor U5097 (N_5097,N_220,N_1694);
xnor U5098 (N_5098,N_1321,N_359);
xnor U5099 (N_5099,N_2738,N_2358);
or U5100 (N_5100,N_64,N_451);
nand U5101 (N_5101,N_2007,N_1873);
nand U5102 (N_5102,N_2224,N_905);
xor U5103 (N_5103,N_2516,N_2671);
and U5104 (N_5104,N_2392,N_82);
or U5105 (N_5105,N_2921,N_715);
xor U5106 (N_5106,N_1579,N_2633);
xnor U5107 (N_5107,N_2586,N_2);
nand U5108 (N_5108,N_427,N_507);
nor U5109 (N_5109,N_191,N_2169);
xnor U5110 (N_5110,N_784,N_1857);
nor U5111 (N_5111,N_1105,N_2965);
nor U5112 (N_5112,N_1622,N_2730);
and U5113 (N_5113,N_1186,N_1439);
nand U5114 (N_5114,N_890,N_167);
nand U5115 (N_5115,N_2827,N_2385);
or U5116 (N_5116,N_2262,N_527);
xor U5117 (N_5117,N_2838,N_2157);
xnor U5118 (N_5118,N_1039,N_2852);
nor U5119 (N_5119,N_2752,N_1426);
nor U5120 (N_5120,N_2875,N_2824);
nand U5121 (N_5121,N_1172,N_825);
nor U5122 (N_5122,N_2456,N_379);
nor U5123 (N_5123,N_176,N_1062);
nand U5124 (N_5124,N_1605,N_2590);
nor U5125 (N_5125,N_367,N_762);
or U5126 (N_5126,N_2507,N_1059);
or U5127 (N_5127,N_736,N_2169);
or U5128 (N_5128,N_711,N_2880);
nand U5129 (N_5129,N_1030,N_822);
nand U5130 (N_5130,N_215,N_1606);
or U5131 (N_5131,N_1542,N_1470);
and U5132 (N_5132,N_2680,N_158);
and U5133 (N_5133,N_2890,N_319);
nand U5134 (N_5134,N_1939,N_1995);
nor U5135 (N_5135,N_2361,N_214);
xor U5136 (N_5136,N_2349,N_532);
and U5137 (N_5137,N_1041,N_868);
nand U5138 (N_5138,N_635,N_1008);
nor U5139 (N_5139,N_1141,N_207);
nand U5140 (N_5140,N_2118,N_2712);
and U5141 (N_5141,N_2663,N_1930);
or U5142 (N_5142,N_2065,N_1133);
or U5143 (N_5143,N_828,N_2147);
and U5144 (N_5144,N_1307,N_1701);
xor U5145 (N_5145,N_546,N_2386);
nand U5146 (N_5146,N_1919,N_358);
nand U5147 (N_5147,N_597,N_1614);
and U5148 (N_5148,N_2253,N_436);
and U5149 (N_5149,N_853,N_44);
and U5150 (N_5150,N_92,N_715);
or U5151 (N_5151,N_1335,N_603);
nor U5152 (N_5152,N_671,N_2318);
xor U5153 (N_5153,N_300,N_731);
nand U5154 (N_5154,N_285,N_2438);
nand U5155 (N_5155,N_972,N_1600);
xor U5156 (N_5156,N_2120,N_1545);
and U5157 (N_5157,N_2471,N_414);
or U5158 (N_5158,N_2688,N_978);
nand U5159 (N_5159,N_1252,N_1504);
and U5160 (N_5160,N_1207,N_2299);
nand U5161 (N_5161,N_767,N_1725);
xnor U5162 (N_5162,N_1993,N_1208);
xor U5163 (N_5163,N_1151,N_561);
xor U5164 (N_5164,N_462,N_644);
nor U5165 (N_5165,N_1207,N_1270);
nor U5166 (N_5166,N_2502,N_1175);
nor U5167 (N_5167,N_447,N_2028);
nor U5168 (N_5168,N_2976,N_1257);
and U5169 (N_5169,N_2931,N_788);
or U5170 (N_5170,N_1345,N_1016);
nor U5171 (N_5171,N_2270,N_291);
and U5172 (N_5172,N_1966,N_1107);
nand U5173 (N_5173,N_2112,N_1095);
and U5174 (N_5174,N_1235,N_1389);
nand U5175 (N_5175,N_1863,N_2887);
and U5176 (N_5176,N_1380,N_973);
nor U5177 (N_5177,N_2584,N_1600);
and U5178 (N_5178,N_832,N_1996);
xnor U5179 (N_5179,N_900,N_2809);
or U5180 (N_5180,N_2033,N_2585);
and U5181 (N_5181,N_209,N_2816);
nor U5182 (N_5182,N_2221,N_2432);
and U5183 (N_5183,N_2549,N_2716);
and U5184 (N_5184,N_2775,N_783);
xnor U5185 (N_5185,N_2737,N_746);
nor U5186 (N_5186,N_2020,N_1617);
nand U5187 (N_5187,N_2680,N_446);
nand U5188 (N_5188,N_1908,N_2600);
or U5189 (N_5189,N_342,N_1896);
or U5190 (N_5190,N_2898,N_2342);
or U5191 (N_5191,N_171,N_181);
or U5192 (N_5192,N_726,N_1715);
xnor U5193 (N_5193,N_44,N_1748);
nor U5194 (N_5194,N_2891,N_2957);
nor U5195 (N_5195,N_2349,N_1059);
or U5196 (N_5196,N_498,N_1113);
nand U5197 (N_5197,N_2080,N_1506);
nand U5198 (N_5198,N_1945,N_708);
nand U5199 (N_5199,N_618,N_1299);
or U5200 (N_5200,N_276,N_918);
or U5201 (N_5201,N_131,N_2206);
or U5202 (N_5202,N_2087,N_2710);
nand U5203 (N_5203,N_681,N_2791);
nor U5204 (N_5204,N_1167,N_2963);
xor U5205 (N_5205,N_2090,N_0);
and U5206 (N_5206,N_7,N_792);
nor U5207 (N_5207,N_461,N_2572);
or U5208 (N_5208,N_65,N_1756);
nand U5209 (N_5209,N_1429,N_968);
and U5210 (N_5210,N_1672,N_1020);
xnor U5211 (N_5211,N_2864,N_2074);
and U5212 (N_5212,N_41,N_1494);
xnor U5213 (N_5213,N_2042,N_2500);
and U5214 (N_5214,N_1109,N_2909);
or U5215 (N_5215,N_1337,N_1946);
nand U5216 (N_5216,N_274,N_1951);
xor U5217 (N_5217,N_2958,N_1353);
nor U5218 (N_5218,N_689,N_1249);
nor U5219 (N_5219,N_1956,N_2820);
nor U5220 (N_5220,N_746,N_171);
nand U5221 (N_5221,N_376,N_2198);
nand U5222 (N_5222,N_2032,N_1480);
nand U5223 (N_5223,N_2186,N_2394);
nor U5224 (N_5224,N_1303,N_2578);
nor U5225 (N_5225,N_914,N_2476);
nor U5226 (N_5226,N_95,N_1401);
or U5227 (N_5227,N_1035,N_1709);
and U5228 (N_5228,N_532,N_1677);
and U5229 (N_5229,N_1929,N_665);
and U5230 (N_5230,N_2391,N_2610);
or U5231 (N_5231,N_2770,N_2241);
or U5232 (N_5232,N_901,N_656);
nand U5233 (N_5233,N_452,N_2893);
and U5234 (N_5234,N_616,N_965);
and U5235 (N_5235,N_2715,N_2667);
and U5236 (N_5236,N_1438,N_1702);
xor U5237 (N_5237,N_2851,N_2666);
or U5238 (N_5238,N_2751,N_2529);
or U5239 (N_5239,N_1181,N_2488);
xnor U5240 (N_5240,N_920,N_2742);
xor U5241 (N_5241,N_580,N_234);
or U5242 (N_5242,N_903,N_2614);
nand U5243 (N_5243,N_1492,N_341);
nor U5244 (N_5244,N_2364,N_623);
nand U5245 (N_5245,N_1244,N_1565);
xnor U5246 (N_5246,N_1895,N_1520);
or U5247 (N_5247,N_412,N_1757);
nand U5248 (N_5248,N_1088,N_1962);
or U5249 (N_5249,N_492,N_1686);
or U5250 (N_5250,N_2152,N_2507);
xor U5251 (N_5251,N_289,N_2663);
nor U5252 (N_5252,N_507,N_1906);
nand U5253 (N_5253,N_778,N_1148);
or U5254 (N_5254,N_1835,N_1508);
xnor U5255 (N_5255,N_2156,N_2888);
nand U5256 (N_5256,N_711,N_2816);
nand U5257 (N_5257,N_2157,N_1191);
or U5258 (N_5258,N_1164,N_2075);
and U5259 (N_5259,N_2679,N_1588);
xor U5260 (N_5260,N_587,N_2879);
xnor U5261 (N_5261,N_1953,N_1118);
or U5262 (N_5262,N_809,N_2503);
or U5263 (N_5263,N_2851,N_529);
nor U5264 (N_5264,N_2735,N_2233);
and U5265 (N_5265,N_2740,N_1164);
and U5266 (N_5266,N_1773,N_1207);
or U5267 (N_5267,N_2707,N_1046);
nand U5268 (N_5268,N_2029,N_2083);
and U5269 (N_5269,N_156,N_385);
and U5270 (N_5270,N_345,N_367);
xnor U5271 (N_5271,N_2040,N_2808);
xnor U5272 (N_5272,N_695,N_2606);
and U5273 (N_5273,N_2980,N_1649);
nand U5274 (N_5274,N_2996,N_2581);
or U5275 (N_5275,N_1682,N_1402);
nand U5276 (N_5276,N_473,N_1151);
nor U5277 (N_5277,N_2923,N_609);
xnor U5278 (N_5278,N_957,N_1567);
xor U5279 (N_5279,N_757,N_788);
and U5280 (N_5280,N_2395,N_156);
xor U5281 (N_5281,N_20,N_676);
or U5282 (N_5282,N_2544,N_2257);
nand U5283 (N_5283,N_2862,N_1782);
and U5284 (N_5284,N_409,N_1964);
and U5285 (N_5285,N_2459,N_2750);
nand U5286 (N_5286,N_876,N_1320);
nand U5287 (N_5287,N_2484,N_1300);
and U5288 (N_5288,N_1917,N_92);
or U5289 (N_5289,N_1872,N_2682);
xnor U5290 (N_5290,N_2502,N_11);
nand U5291 (N_5291,N_1626,N_2425);
nor U5292 (N_5292,N_2765,N_1062);
nand U5293 (N_5293,N_1814,N_2843);
or U5294 (N_5294,N_2454,N_222);
nor U5295 (N_5295,N_1054,N_2151);
or U5296 (N_5296,N_819,N_1664);
or U5297 (N_5297,N_2676,N_48);
xnor U5298 (N_5298,N_1541,N_593);
xor U5299 (N_5299,N_1036,N_236);
nor U5300 (N_5300,N_210,N_2655);
nor U5301 (N_5301,N_1966,N_2683);
xnor U5302 (N_5302,N_1427,N_2796);
or U5303 (N_5303,N_435,N_2501);
or U5304 (N_5304,N_702,N_1333);
nor U5305 (N_5305,N_2686,N_231);
nand U5306 (N_5306,N_405,N_557);
xnor U5307 (N_5307,N_155,N_1062);
or U5308 (N_5308,N_2738,N_55);
xor U5309 (N_5309,N_1731,N_2395);
or U5310 (N_5310,N_1501,N_2116);
nand U5311 (N_5311,N_841,N_791);
or U5312 (N_5312,N_34,N_1015);
and U5313 (N_5313,N_296,N_295);
and U5314 (N_5314,N_258,N_2900);
nand U5315 (N_5315,N_1473,N_397);
nor U5316 (N_5316,N_1683,N_2771);
nor U5317 (N_5317,N_2340,N_2244);
xnor U5318 (N_5318,N_1471,N_683);
nor U5319 (N_5319,N_2719,N_1189);
xnor U5320 (N_5320,N_640,N_1462);
xor U5321 (N_5321,N_1434,N_504);
xor U5322 (N_5322,N_1135,N_2625);
xor U5323 (N_5323,N_2971,N_157);
xnor U5324 (N_5324,N_2451,N_2217);
or U5325 (N_5325,N_651,N_1644);
nor U5326 (N_5326,N_108,N_1293);
and U5327 (N_5327,N_957,N_554);
and U5328 (N_5328,N_2283,N_368);
or U5329 (N_5329,N_1450,N_1639);
or U5330 (N_5330,N_156,N_2738);
or U5331 (N_5331,N_2748,N_2444);
or U5332 (N_5332,N_1630,N_2396);
or U5333 (N_5333,N_1202,N_2539);
or U5334 (N_5334,N_1710,N_2620);
xnor U5335 (N_5335,N_1335,N_579);
nand U5336 (N_5336,N_774,N_1730);
nor U5337 (N_5337,N_1663,N_95);
or U5338 (N_5338,N_1150,N_2120);
or U5339 (N_5339,N_1875,N_2988);
xor U5340 (N_5340,N_1847,N_945);
nor U5341 (N_5341,N_1227,N_52);
nor U5342 (N_5342,N_1496,N_2064);
nand U5343 (N_5343,N_895,N_599);
and U5344 (N_5344,N_1666,N_586);
nor U5345 (N_5345,N_2159,N_1032);
and U5346 (N_5346,N_1738,N_836);
xnor U5347 (N_5347,N_236,N_948);
and U5348 (N_5348,N_1457,N_1498);
nand U5349 (N_5349,N_2435,N_24);
and U5350 (N_5350,N_2745,N_2704);
nor U5351 (N_5351,N_2135,N_2708);
nor U5352 (N_5352,N_2063,N_2804);
nor U5353 (N_5353,N_562,N_19);
or U5354 (N_5354,N_332,N_1852);
or U5355 (N_5355,N_1680,N_2605);
and U5356 (N_5356,N_649,N_740);
nor U5357 (N_5357,N_2645,N_2762);
nor U5358 (N_5358,N_34,N_1961);
and U5359 (N_5359,N_2564,N_70);
nor U5360 (N_5360,N_411,N_1599);
nand U5361 (N_5361,N_2684,N_576);
nor U5362 (N_5362,N_1088,N_431);
and U5363 (N_5363,N_475,N_1932);
xnor U5364 (N_5364,N_13,N_856);
xnor U5365 (N_5365,N_301,N_997);
nand U5366 (N_5366,N_1699,N_880);
and U5367 (N_5367,N_2643,N_1282);
nor U5368 (N_5368,N_324,N_2837);
nand U5369 (N_5369,N_2258,N_1718);
and U5370 (N_5370,N_2962,N_150);
or U5371 (N_5371,N_187,N_595);
and U5372 (N_5372,N_2473,N_1578);
and U5373 (N_5373,N_1407,N_923);
or U5374 (N_5374,N_106,N_2565);
nand U5375 (N_5375,N_287,N_281);
and U5376 (N_5376,N_2419,N_2930);
or U5377 (N_5377,N_1455,N_2595);
and U5378 (N_5378,N_2006,N_1299);
xnor U5379 (N_5379,N_212,N_755);
xnor U5380 (N_5380,N_2132,N_262);
nand U5381 (N_5381,N_1847,N_2065);
nand U5382 (N_5382,N_276,N_793);
xnor U5383 (N_5383,N_1719,N_1385);
nand U5384 (N_5384,N_1087,N_1139);
xnor U5385 (N_5385,N_757,N_2561);
and U5386 (N_5386,N_691,N_610);
nor U5387 (N_5387,N_2989,N_2851);
and U5388 (N_5388,N_1614,N_835);
xor U5389 (N_5389,N_2685,N_607);
and U5390 (N_5390,N_2199,N_2156);
and U5391 (N_5391,N_2166,N_1946);
nand U5392 (N_5392,N_2582,N_136);
nor U5393 (N_5393,N_2609,N_1803);
and U5394 (N_5394,N_1575,N_967);
nor U5395 (N_5395,N_1060,N_1228);
or U5396 (N_5396,N_1598,N_2187);
nand U5397 (N_5397,N_2326,N_620);
nor U5398 (N_5398,N_1139,N_1014);
nand U5399 (N_5399,N_349,N_2910);
xnor U5400 (N_5400,N_2553,N_1708);
nor U5401 (N_5401,N_2770,N_2520);
nor U5402 (N_5402,N_749,N_2794);
or U5403 (N_5403,N_1805,N_819);
or U5404 (N_5404,N_2716,N_2948);
nor U5405 (N_5405,N_2034,N_1307);
nor U5406 (N_5406,N_1886,N_2544);
or U5407 (N_5407,N_184,N_2820);
and U5408 (N_5408,N_2837,N_1937);
nor U5409 (N_5409,N_1467,N_2764);
nand U5410 (N_5410,N_167,N_1304);
nor U5411 (N_5411,N_879,N_860);
and U5412 (N_5412,N_1079,N_2489);
nand U5413 (N_5413,N_22,N_1332);
or U5414 (N_5414,N_2237,N_17);
xnor U5415 (N_5415,N_2562,N_2179);
or U5416 (N_5416,N_1195,N_714);
xnor U5417 (N_5417,N_698,N_1629);
xnor U5418 (N_5418,N_2389,N_1148);
nor U5419 (N_5419,N_969,N_2890);
or U5420 (N_5420,N_2705,N_1377);
or U5421 (N_5421,N_2871,N_371);
nor U5422 (N_5422,N_317,N_638);
nor U5423 (N_5423,N_2338,N_2799);
nor U5424 (N_5424,N_2674,N_2065);
nand U5425 (N_5425,N_1924,N_1391);
and U5426 (N_5426,N_2739,N_1605);
or U5427 (N_5427,N_2016,N_2088);
xor U5428 (N_5428,N_1521,N_372);
nand U5429 (N_5429,N_1334,N_1278);
or U5430 (N_5430,N_2381,N_1530);
xor U5431 (N_5431,N_1266,N_93);
nand U5432 (N_5432,N_155,N_2577);
nand U5433 (N_5433,N_726,N_1618);
nand U5434 (N_5434,N_2826,N_2141);
nand U5435 (N_5435,N_2973,N_1772);
xor U5436 (N_5436,N_1982,N_923);
and U5437 (N_5437,N_2104,N_1032);
nor U5438 (N_5438,N_1639,N_2216);
and U5439 (N_5439,N_1130,N_85);
xor U5440 (N_5440,N_2099,N_41);
xnor U5441 (N_5441,N_684,N_1005);
nor U5442 (N_5442,N_389,N_2677);
or U5443 (N_5443,N_1152,N_161);
or U5444 (N_5444,N_2266,N_982);
nand U5445 (N_5445,N_2102,N_265);
nand U5446 (N_5446,N_1058,N_1501);
or U5447 (N_5447,N_1773,N_1401);
nor U5448 (N_5448,N_2239,N_1664);
nor U5449 (N_5449,N_2061,N_1202);
nand U5450 (N_5450,N_928,N_1321);
nor U5451 (N_5451,N_2222,N_1050);
nand U5452 (N_5452,N_2920,N_1396);
or U5453 (N_5453,N_1797,N_1829);
nand U5454 (N_5454,N_1153,N_1393);
nand U5455 (N_5455,N_2371,N_939);
xor U5456 (N_5456,N_1132,N_1317);
nor U5457 (N_5457,N_2003,N_1987);
and U5458 (N_5458,N_2869,N_927);
xor U5459 (N_5459,N_2507,N_291);
and U5460 (N_5460,N_1772,N_2185);
nor U5461 (N_5461,N_1089,N_1203);
or U5462 (N_5462,N_1693,N_976);
nand U5463 (N_5463,N_1340,N_915);
or U5464 (N_5464,N_1844,N_2493);
and U5465 (N_5465,N_2591,N_734);
xnor U5466 (N_5466,N_956,N_1045);
nand U5467 (N_5467,N_2993,N_2865);
or U5468 (N_5468,N_1212,N_323);
nor U5469 (N_5469,N_1793,N_2254);
nand U5470 (N_5470,N_1367,N_1835);
nand U5471 (N_5471,N_45,N_1560);
xnor U5472 (N_5472,N_247,N_2999);
nor U5473 (N_5473,N_816,N_769);
nor U5474 (N_5474,N_2475,N_2830);
nand U5475 (N_5475,N_2485,N_728);
nor U5476 (N_5476,N_1514,N_642);
nand U5477 (N_5477,N_665,N_2902);
nand U5478 (N_5478,N_2511,N_529);
and U5479 (N_5479,N_1974,N_434);
nand U5480 (N_5480,N_1358,N_1550);
or U5481 (N_5481,N_2259,N_2565);
and U5482 (N_5482,N_509,N_1232);
and U5483 (N_5483,N_1298,N_180);
nor U5484 (N_5484,N_2734,N_729);
xnor U5485 (N_5485,N_2163,N_670);
xnor U5486 (N_5486,N_99,N_1064);
nor U5487 (N_5487,N_1001,N_2959);
xnor U5488 (N_5488,N_1860,N_2707);
xor U5489 (N_5489,N_2940,N_545);
nand U5490 (N_5490,N_1699,N_1495);
and U5491 (N_5491,N_336,N_1648);
and U5492 (N_5492,N_1740,N_1781);
nand U5493 (N_5493,N_1895,N_2038);
nand U5494 (N_5494,N_286,N_2410);
xnor U5495 (N_5495,N_530,N_1235);
and U5496 (N_5496,N_1373,N_426);
and U5497 (N_5497,N_1495,N_2570);
nor U5498 (N_5498,N_1305,N_1549);
xor U5499 (N_5499,N_1846,N_1135);
xor U5500 (N_5500,N_2828,N_788);
and U5501 (N_5501,N_2998,N_122);
xor U5502 (N_5502,N_2715,N_2303);
and U5503 (N_5503,N_2005,N_1687);
nor U5504 (N_5504,N_698,N_235);
xnor U5505 (N_5505,N_1040,N_2604);
xor U5506 (N_5506,N_614,N_590);
and U5507 (N_5507,N_2764,N_2804);
nand U5508 (N_5508,N_152,N_136);
xor U5509 (N_5509,N_1516,N_2648);
nand U5510 (N_5510,N_1917,N_915);
nor U5511 (N_5511,N_2365,N_1206);
and U5512 (N_5512,N_32,N_1437);
xor U5513 (N_5513,N_2511,N_1624);
and U5514 (N_5514,N_55,N_281);
xor U5515 (N_5515,N_1208,N_2820);
nor U5516 (N_5516,N_2839,N_1367);
and U5517 (N_5517,N_651,N_114);
xor U5518 (N_5518,N_421,N_766);
nand U5519 (N_5519,N_1738,N_1672);
nor U5520 (N_5520,N_2785,N_2231);
nand U5521 (N_5521,N_1336,N_285);
nand U5522 (N_5522,N_543,N_2834);
or U5523 (N_5523,N_726,N_2443);
nor U5524 (N_5524,N_1844,N_2564);
or U5525 (N_5525,N_1443,N_931);
nand U5526 (N_5526,N_1887,N_312);
and U5527 (N_5527,N_216,N_1282);
xnor U5528 (N_5528,N_1704,N_983);
and U5529 (N_5529,N_244,N_965);
nand U5530 (N_5530,N_1612,N_2491);
xnor U5531 (N_5531,N_449,N_1369);
nand U5532 (N_5532,N_1320,N_2942);
or U5533 (N_5533,N_2617,N_754);
and U5534 (N_5534,N_1934,N_536);
and U5535 (N_5535,N_93,N_1751);
xnor U5536 (N_5536,N_925,N_2919);
and U5537 (N_5537,N_1957,N_1737);
nor U5538 (N_5538,N_1174,N_1680);
nor U5539 (N_5539,N_1658,N_1688);
nor U5540 (N_5540,N_814,N_2955);
nor U5541 (N_5541,N_2323,N_1394);
and U5542 (N_5542,N_2843,N_2150);
nand U5543 (N_5543,N_1663,N_432);
nor U5544 (N_5544,N_1715,N_415);
nand U5545 (N_5545,N_1699,N_2869);
xnor U5546 (N_5546,N_2734,N_1783);
xor U5547 (N_5547,N_996,N_2806);
xor U5548 (N_5548,N_2890,N_1278);
xnor U5549 (N_5549,N_1107,N_1834);
nand U5550 (N_5550,N_2698,N_2812);
nand U5551 (N_5551,N_1846,N_906);
nor U5552 (N_5552,N_1969,N_254);
or U5553 (N_5553,N_2211,N_1277);
and U5554 (N_5554,N_1097,N_2551);
nor U5555 (N_5555,N_613,N_1965);
xor U5556 (N_5556,N_2101,N_1511);
nor U5557 (N_5557,N_822,N_926);
nand U5558 (N_5558,N_444,N_1665);
nor U5559 (N_5559,N_2380,N_144);
xor U5560 (N_5560,N_591,N_857);
nor U5561 (N_5561,N_2275,N_116);
xor U5562 (N_5562,N_1389,N_2063);
nand U5563 (N_5563,N_323,N_2798);
xnor U5564 (N_5564,N_1892,N_296);
xor U5565 (N_5565,N_755,N_2239);
xor U5566 (N_5566,N_1701,N_1539);
and U5567 (N_5567,N_356,N_2357);
xnor U5568 (N_5568,N_1487,N_1901);
nand U5569 (N_5569,N_735,N_2534);
nor U5570 (N_5570,N_591,N_2446);
and U5571 (N_5571,N_2747,N_2913);
and U5572 (N_5572,N_1066,N_1233);
or U5573 (N_5573,N_1146,N_481);
and U5574 (N_5574,N_2644,N_2707);
nor U5575 (N_5575,N_476,N_1763);
nor U5576 (N_5576,N_1051,N_2859);
and U5577 (N_5577,N_742,N_927);
or U5578 (N_5578,N_2341,N_1929);
nor U5579 (N_5579,N_1997,N_2832);
nor U5580 (N_5580,N_2704,N_1539);
nand U5581 (N_5581,N_998,N_2591);
nor U5582 (N_5582,N_2823,N_539);
xor U5583 (N_5583,N_21,N_198);
or U5584 (N_5584,N_1254,N_2505);
xor U5585 (N_5585,N_2881,N_699);
nor U5586 (N_5586,N_1751,N_1476);
or U5587 (N_5587,N_620,N_1304);
or U5588 (N_5588,N_107,N_80);
xor U5589 (N_5589,N_1201,N_1016);
xor U5590 (N_5590,N_1826,N_1825);
xnor U5591 (N_5591,N_459,N_722);
nor U5592 (N_5592,N_1526,N_2099);
nor U5593 (N_5593,N_1769,N_2032);
and U5594 (N_5594,N_750,N_603);
and U5595 (N_5595,N_1729,N_441);
and U5596 (N_5596,N_388,N_2833);
nor U5597 (N_5597,N_739,N_2318);
nand U5598 (N_5598,N_2034,N_458);
and U5599 (N_5599,N_2252,N_1387);
and U5600 (N_5600,N_2902,N_652);
nor U5601 (N_5601,N_1969,N_1815);
nand U5602 (N_5602,N_35,N_2376);
xor U5603 (N_5603,N_520,N_1174);
and U5604 (N_5604,N_1665,N_2183);
and U5605 (N_5605,N_1723,N_463);
or U5606 (N_5606,N_2690,N_169);
nor U5607 (N_5607,N_2018,N_946);
and U5608 (N_5608,N_2818,N_2140);
or U5609 (N_5609,N_649,N_2536);
nand U5610 (N_5610,N_2080,N_1034);
nor U5611 (N_5611,N_999,N_1394);
and U5612 (N_5612,N_935,N_2067);
xor U5613 (N_5613,N_1777,N_2260);
nor U5614 (N_5614,N_1818,N_62);
and U5615 (N_5615,N_182,N_2268);
xor U5616 (N_5616,N_712,N_990);
nor U5617 (N_5617,N_1997,N_1396);
nand U5618 (N_5618,N_2972,N_1897);
or U5619 (N_5619,N_441,N_2196);
xnor U5620 (N_5620,N_2506,N_145);
and U5621 (N_5621,N_85,N_1767);
or U5622 (N_5622,N_2304,N_317);
nand U5623 (N_5623,N_872,N_1508);
and U5624 (N_5624,N_497,N_2672);
xnor U5625 (N_5625,N_1958,N_1174);
and U5626 (N_5626,N_1499,N_1049);
nor U5627 (N_5627,N_1865,N_2286);
and U5628 (N_5628,N_1832,N_1555);
nand U5629 (N_5629,N_2253,N_2044);
and U5630 (N_5630,N_387,N_1571);
nand U5631 (N_5631,N_1054,N_65);
nor U5632 (N_5632,N_2876,N_1336);
xor U5633 (N_5633,N_1425,N_2553);
or U5634 (N_5634,N_1622,N_565);
or U5635 (N_5635,N_2961,N_452);
and U5636 (N_5636,N_678,N_673);
xor U5637 (N_5637,N_1893,N_819);
nor U5638 (N_5638,N_1707,N_1539);
nand U5639 (N_5639,N_2159,N_1872);
xor U5640 (N_5640,N_2448,N_13);
nand U5641 (N_5641,N_136,N_934);
and U5642 (N_5642,N_1062,N_2847);
nor U5643 (N_5643,N_467,N_975);
and U5644 (N_5644,N_2058,N_840);
nor U5645 (N_5645,N_2952,N_2332);
xor U5646 (N_5646,N_1187,N_2184);
nor U5647 (N_5647,N_1863,N_725);
or U5648 (N_5648,N_1020,N_1705);
nor U5649 (N_5649,N_594,N_856);
and U5650 (N_5650,N_1797,N_278);
and U5651 (N_5651,N_90,N_2014);
xor U5652 (N_5652,N_916,N_2412);
nand U5653 (N_5653,N_1706,N_1484);
nand U5654 (N_5654,N_1538,N_903);
xnor U5655 (N_5655,N_1227,N_2718);
and U5656 (N_5656,N_1397,N_93);
nor U5657 (N_5657,N_480,N_1520);
nor U5658 (N_5658,N_238,N_1314);
or U5659 (N_5659,N_2084,N_2330);
and U5660 (N_5660,N_1908,N_2350);
nand U5661 (N_5661,N_2456,N_2010);
nand U5662 (N_5662,N_1319,N_487);
xnor U5663 (N_5663,N_1548,N_1288);
and U5664 (N_5664,N_1799,N_2209);
xnor U5665 (N_5665,N_666,N_1053);
nand U5666 (N_5666,N_1296,N_1496);
nor U5667 (N_5667,N_2223,N_2298);
xor U5668 (N_5668,N_2637,N_1322);
nor U5669 (N_5669,N_2076,N_663);
or U5670 (N_5670,N_2672,N_897);
or U5671 (N_5671,N_321,N_1413);
xor U5672 (N_5672,N_2804,N_719);
or U5673 (N_5673,N_765,N_1505);
nor U5674 (N_5674,N_2323,N_1556);
or U5675 (N_5675,N_114,N_1847);
nor U5676 (N_5676,N_2954,N_1471);
or U5677 (N_5677,N_1933,N_1129);
or U5678 (N_5678,N_1494,N_2212);
or U5679 (N_5679,N_2311,N_1863);
nor U5680 (N_5680,N_69,N_2716);
nor U5681 (N_5681,N_756,N_1145);
xnor U5682 (N_5682,N_1220,N_407);
or U5683 (N_5683,N_656,N_154);
nand U5684 (N_5684,N_309,N_1211);
or U5685 (N_5685,N_831,N_161);
or U5686 (N_5686,N_2086,N_1154);
nor U5687 (N_5687,N_1092,N_2212);
xor U5688 (N_5688,N_800,N_218);
nor U5689 (N_5689,N_1319,N_2040);
nor U5690 (N_5690,N_2164,N_1132);
nor U5691 (N_5691,N_1676,N_295);
nand U5692 (N_5692,N_711,N_1384);
nand U5693 (N_5693,N_1283,N_1899);
nand U5694 (N_5694,N_528,N_1880);
xnor U5695 (N_5695,N_514,N_666);
and U5696 (N_5696,N_2036,N_2350);
and U5697 (N_5697,N_2934,N_2433);
xnor U5698 (N_5698,N_1001,N_2247);
and U5699 (N_5699,N_1852,N_1585);
nor U5700 (N_5700,N_610,N_1276);
and U5701 (N_5701,N_1696,N_1188);
and U5702 (N_5702,N_366,N_104);
and U5703 (N_5703,N_1058,N_2743);
nor U5704 (N_5704,N_2269,N_1872);
xnor U5705 (N_5705,N_462,N_220);
nor U5706 (N_5706,N_966,N_1949);
xor U5707 (N_5707,N_2936,N_477);
nor U5708 (N_5708,N_191,N_603);
xnor U5709 (N_5709,N_2582,N_2862);
or U5710 (N_5710,N_347,N_2896);
nand U5711 (N_5711,N_1883,N_102);
nand U5712 (N_5712,N_1510,N_312);
xnor U5713 (N_5713,N_2697,N_282);
or U5714 (N_5714,N_2241,N_1561);
xor U5715 (N_5715,N_506,N_2642);
nand U5716 (N_5716,N_947,N_2203);
xnor U5717 (N_5717,N_2305,N_2644);
nor U5718 (N_5718,N_2925,N_862);
nor U5719 (N_5719,N_2447,N_25);
nor U5720 (N_5720,N_1443,N_1343);
nor U5721 (N_5721,N_2865,N_1481);
nand U5722 (N_5722,N_2836,N_2281);
nor U5723 (N_5723,N_350,N_1676);
and U5724 (N_5724,N_1225,N_1030);
or U5725 (N_5725,N_1740,N_1426);
xnor U5726 (N_5726,N_954,N_1522);
and U5727 (N_5727,N_1900,N_657);
or U5728 (N_5728,N_731,N_822);
and U5729 (N_5729,N_2614,N_2658);
nand U5730 (N_5730,N_2891,N_2870);
or U5731 (N_5731,N_2064,N_2191);
nand U5732 (N_5732,N_1815,N_116);
nand U5733 (N_5733,N_1835,N_130);
and U5734 (N_5734,N_573,N_39);
xnor U5735 (N_5735,N_1083,N_497);
nor U5736 (N_5736,N_1104,N_2370);
nand U5737 (N_5737,N_264,N_1981);
nand U5738 (N_5738,N_19,N_2265);
or U5739 (N_5739,N_1051,N_761);
and U5740 (N_5740,N_1441,N_2189);
nor U5741 (N_5741,N_2287,N_953);
and U5742 (N_5742,N_1546,N_2343);
and U5743 (N_5743,N_2513,N_1303);
or U5744 (N_5744,N_82,N_87);
and U5745 (N_5745,N_1899,N_1697);
or U5746 (N_5746,N_2823,N_1418);
and U5747 (N_5747,N_1231,N_2977);
nor U5748 (N_5748,N_948,N_2283);
and U5749 (N_5749,N_1842,N_2571);
xor U5750 (N_5750,N_1880,N_2139);
nand U5751 (N_5751,N_1775,N_2975);
nand U5752 (N_5752,N_1717,N_2769);
xnor U5753 (N_5753,N_1140,N_1027);
nand U5754 (N_5754,N_411,N_716);
and U5755 (N_5755,N_2684,N_2396);
or U5756 (N_5756,N_361,N_2200);
or U5757 (N_5757,N_2199,N_1137);
xnor U5758 (N_5758,N_2067,N_819);
and U5759 (N_5759,N_1598,N_1324);
xnor U5760 (N_5760,N_1607,N_158);
and U5761 (N_5761,N_1808,N_565);
nand U5762 (N_5762,N_2518,N_854);
and U5763 (N_5763,N_2262,N_2992);
nor U5764 (N_5764,N_538,N_2189);
and U5765 (N_5765,N_2095,N_808);
xor U5766 (N_5766,N_2924,N_1040);
and U5767 (N_5767,N_2191,N_700);
xor U5768 (N_5768,N_1099,N_1394);
and U5769 (N_5769,N_2566,N_2390);
nand U5770 (N_5770,N_2352,N_895);
or U5771 (N_5771,N_93,N_1137);
or U5772 (N_5772,N_1884,N_838);
nand U5773 (N_5773,N_1127,N_2928);
nand U5774 (N_5774,N_836,N_2567);
or U5775 (N_5775,N_1884,N_1013);
xor U5776 (N_5776,N_2898,N_573);
nor U5777 (N_5777,N_2509,N_1630);
or U5778 (N_5778,N_1080,N_1954);
or U5779 (N_5779,N_1006,N_2542);
and U5780 (N_5780,N_2894,N_1576);
nor U5781 (N_5781,N_2513,N_568);
xor U5782 (N_5782,N_1025,N_2727);
and U5783 (N_5783,N_229,N_172);
or U5784 (N_5784,N_2208,N_2798);
nor U5785 (N_5785,N_1233,N_604);
or U5786 (N_5786,N_704,N_2775);
nand U5787 (N_5787,N_2966,N_1443);
nor U5788 (N_5788,N_619,N_979);
nor U5789 (N_5789,N_799,N_1485);
xnor U5790 (N_5790,N_1214,N_2855);
nor U5791 (N_5791,N_605,N_911);
xor U5792 (N_5792,N_2580,N_1376);
and U5793 (N_5793,N_2546,N_1572);
nand U5794 (N_5794,N_2003,N_138);
and U5795 (N_5795,N_2929,N_2516);
or U5796 (N_5796,N_1696,N_504);
nor U5797 (N_5797,N_2977,N_1624);
xnor U5798 (N_5798,N_1878,N_1842);
nand U5799 (N_5799,N_1144,N_2052);
nand U5800 (N_5800,N_450,N_700);
or U5801 (N_5801,N_21,N_788);
and U5802 (N_5802,N_1716,N_1293);
xor U5803 (N_5803,N_345,N_1187);
or U5804 (N_5804,N_685,N_2246);
nand U5805 (N_5805,N_1168,N_171);
nor U5806 (N_5806,N_601,N_2334);
nor U5807 (N_5807,N_406,N_865);
or U5808 (N_5808,N_145,N_521);
nand U5809 (N_5809,N_978,N_188);
and U5810 (N_5810,N_33,N_2280);
nor U5811 (N_5811,N_2976,N_1717);
or U5812 (N_5812,N_2631,N_1207);
nand U5813 (N_5813,N_743,N_588);
nand U5814 (N_5814,N_644,N_2092);
or U5815 (N_5815,N_1456,N_2926);
or U5816 (N_5816,N_508,N_2921);
nor U5817 (N_5817,N_1581,N_2401);
nand U5818 (N_5818,N_2016,N_854);
and U5819 (N_5819,N_2381,N_1458);
nand U5820 (N_5820,N_1477,N_2887);
or U5821 (N_5821,N_1101,N_972);
nand U5822 (N_5822,N_2594,N_1611);
xnor U5823 (N_5823,N_484,N_400);
or U5824 (N_5824,N_1412,N_478);
nand U5825 (N_5825,N_2947,N_148);
xor U5826 (N_5826,N_251,N_1621);
and U5827 (N_5827,N_1627,N_1671);
nor U5828 (N_5828,N_2934,N_2475);
and U5829 (N_5829,N_1186,N_354);
nor U5830 (N_5830,N_2033,N_2892);
nor U5831 (N_5831,N_1235,N_1363);
and U5832 (N_5832,N_1777,N_372);
and U5833 (N_5833,N_2841,N_2220);
xnor U5834 (N_5834,N_2548,N_1172);
or U5835 (N_5835,N_252,N_2875);
xnor U5836 (N_5836,N_2578,N_466);
and U5837 (N_5837,N_1654,N_971);
nor U5838 (N_5838,N_460,N_2440);
nand U5839 (N_5839,N_1775,N_581);
nor U5840 (N_5840,N_593,N_2933);
xor U5841 (N_5841,N_1447,N_2922);
nand U5842 (N_5842,N_246,N_929);
or U5843 (N_5843,N_1415,N_1178);
nor U5844 (N_5844,N_825,N_2572);
and U5845 (N_5845,N_1708,N_1189);
and U5846 (N_5846,N_1531,N_2685);
and U5847 (N_5847,N_1270,N_39);
xor U5848 (N_5848,N_788,N_22);
or U5849 (N_5849,N_2281,N_378);
nand U5850 (N_5850,N_2378,N_2718);
nor U5851 (N_5851,N_2059,N_1211);
nor U5852 (N_5852,N_1373,N_1408);
nand U5853 (N_5853,N_2774,N_992);
and U5854 (N_5854,N_954,N_174);
or U5855 (N_5855,N_2341,N_2378);
and U5856 (N_5856,N_1733,N_2580);
xor U5857 (N_5857,N_1832,N_2815);
and U5858 (N_5858,N_398,N_1862);
or U5859 (N_5859,N_1116,N_1218);
nor U5860 (N_5860,N_2301,N_1311);
and U5861 (N_5861,N_1653,N_127);
nor U5862 (N_5862,N_210,N_2967);
xnor U5863 (N_5863,N_2804,N_628);
xnor U5864 (N_5864,N_1239,N_186);
nand U5865 (N_5865,N_2509,N_2678);
or U5866 (N_5866,N_1824,N_2213);
nand U5867 (N_5867,N_1455,N_233);
or U5868 (N_5868,N_2891,N_141);
and U5869 (N_5869,N_907,N_2849);
and U5870 (N_5870,N_1227,N_2205);
nand U5871 (N_5871,N_1015,N_1684);
xnor U5872 (N_5872,N_1878,N_2833);
and U5873 (N_5873,N_622,N_2791);
nor U5874 (N_5874,N_2022,N_2301);
xor U5875 (N_5875,N_2887,N_1012);
and U5876 (N_5876,N_1427,N_194);
and U5877 (N_5877,N_296,N_80);
nand U5878 (N_5878,N_1126,N_1573);
or U5879 (N_5879,N_882,N_491);
or U5880 (N_5880,N_396,N_1117);
nand U5881 (N_5881,N_1176,N_691);
nand U5882 (N_5882,N_353,N_2018);
xor U5883 (N_5883,N_142,N_306);
and U5884 (N_5884,N_509,N_253);
xor U5885 (N_5885,N_2027,N_2736);
xnor U5886 (N_5886,N_2257,N_1437);
and U5887 (N_5887,N_1176,N_926);
xor U5888 (N_5888,N_995,N_2626);
and U5889 (N_5889,N_2706,N_1743);
and U5890 (N_5890,N_2205,N_991);
nor U5891 (N_5891,N_550,N_1676);
or U5892 (N_5892,N_1951,N_620);
nand U5893 (N_5893,N_2915,N_1282);
nor U5894 (N_5894,N_2456,N_2919);
or U5895 (N_5895,N_341,N_1434);
or U5896 (N_5896,N_1642,N_410);
nand U5897 (N_5897,N_117,N_2587);
and U5898 (N_5898,N_2036,N_1446);
xnor U5899 (N_5899,N_900,N_2073);
xnor U5900 (N_5900,N_2250,N_1197);
xnor U5901 (N_5901,N_2571,N_889);
and U5902 (N_5902,N_60,N_2574);
and U5903 (N_5903,N_401,N_2033);
xor U5904 (N_5904,N_966,N_442);
xnor U5905 (N_5905,N_2674,N_2053);
or U5906 (N_5906,N_2016,N_741);
nor U5907 (N_5907,N_1651,N_1164);
nand U5908 (N_5908,N_912,N_2012);
or U5909 (N_5909,N_2269,N_1124);
or U5910 (N_5910,N_593,N_1057);
or U5911 (N_5911,N_2366,N_1526);
nor U5912 (N_5912,N_2535,N_1246);
and U5913 (N_5913,N_676,N_926);
xnor U5914 (N_5914,N_1643,N_1616);
or U5915 (N_5915,N_2877,N_1342);
and U5916 (N_5916,N_435,N_2745);
xor U5917 (N_5917,N_2582,N_111);
xor U5918 (N_5918,N_736,N_2422);
or U5919 (N_5919,N_2496,N_228);
and U5920 (N_5920,N_2564,N_2501);
and U5921 (N_5921,N_2892,N_729);
xnor U5922 (N_5922,N_1828,N_1699);
nor U5923 (N_5923,N_1916,N_811);
xor U5924 (N_5924,N_737,N_2613);
and U5925 (N_5925,N_2453,N_2442);
nand U5926 (N_5926,N_1004,N_253);
nand U5927 (N_5927,N_2418,N_2694);
nor U5928 (N_5928,N_1876,N_1743);
xor U5929 (N_5929,N_276,N_1711);
xor U5930 (N_5930,N_1316,N_2067);
or U5931 (N_5931,N_1598,N_808);
nor U5932 (N_5932,N_715,N_1937);
nand U5933 (N_5933,N_1836,N_2058);
nand U5934 (N_5934,N_2471,N_2390);
or U5935 (N_5935,N_1160,N_1526);
nand U5936 (N_5936,N_41,N_2843);
and U5937 (N_5937,N_1357,N_2143);
nor U5938 (N_5938,N_87,N_965);
or U5939 (N_5939,N_1206,N_2050);
or U5940 (N_5940,N_2565,N_354);
or U5941 (N_5941,N_2800,N_1085);
or U5942 (N_5942,N_1876,N_1178);
xor U5943 (N_5943,N_755,N_1811);
or U5944 (N_5944,N_968,N_2608);
and U5945 (N_5945,N_466,N_889);
xor U5946 (N_5946,N_2843,N_915);
and U5947 (N_5947,N_1667,N_1160);
and U5948 (N_5948,N_1798,N_1775);
nor U5949 (N_5949,N_1650,N_301);
or U5950 (N_5950,N_2468,N_293);
and U5951 (N_5951,N_1714,N_1009);
and U5952 (N_5952,N_2502,N_224);
or U5953 (N_5953,N_1148,N_1022);
xnor U5954 (N_5954,N_2676,N_2611);
nor U5955 (N_5955,N_2453,N_2353);
nand U5956 (N_5956,N_2470,N_2109);
nor U5957 (N_5957,N_2751,N_584);
and U5958 (N_5958,N_1945,N_518);
and U5959 (N_5959,N_2558,N_2466);
nand U5960 (N_5960,N_1424,N_649);
nor U5961 (N_5961,N_2014,N_967);
xor U5962 (N_5962,N_367,N_1831);
xnor U5963 (N_5963,N_2528,N_1640);
or U5964 (N_5964,N_1007,N_1382);
or U5965 (N_5965,N_2052,N_1854);
xor U5966 (N_5966,N_1491,N_666);
xor U5967 (N_5967,N_296,N_686);
nand U5968 (N_5968,N_2193,N_2784);
or U5969 (N_5969,N_2119,N_2983);
nand U5970 (N_5970,N_2842,N_2484);
xnor U5971 (N_5971,N_2095,N_273);
or U5972 (N_5972,N_2425,N_787);
nand U5973 (N_5973,N_1955,N_1670);
and U5974 (N_5974,N_1909,N_1942);
and U5975 (N_5975,N_412,N_1063);
and U5976 (N_5976,N_2145,N_2160);
xnor U5977 (N_5977,N_501,N_964);
or U5978 (N_5978,N_2555,N_1077);
xor U5979 (N_5979,N_115,N_1977);
nand U5980 (N_5980,N_2093,N_2424);
or U5981 (N_5981,N_1496,N_1284);
nand U5982 (N_5982,N_587,N_488);
nor U5983 (N_5983,N_955,N_76);
and U5984 (N_5984,N_58,N_508);
nor U5985 (N_5985,N_2572,N_1227);
nor U5986 (N_5986,N_1430,N_1204);
and U5987 (N_5987,N_2935,N_2899);
or U5988 (N_5988,N_2845,N_1541);
and U5989 (N_5989,N_2457,N_1447);
xor U5990 (N_5990,N_476,N_2581);
and U5991 (N_5991,N_1174,N_1756);
and U5992 (N_5992,N_363,N_1938);
and U5993 (N_5993,N_2130,N_498);
nand U5994 (N_5994,N_2170,N_414);
nor U5995 (N_5995,N_2821,N_476);
or U5996 (N_5996,N_1299,N_2002);
xor U5997 (N_5997,N_746,N_1056);
or U5998 (N_5998,N_924,N_1677);
or U5999 (N_5999,N_329,N_1618);
nor U6000 (N_6000,N_3631,N_4292);
nor U6001 (N_6001,N_5578,N_4200);
and U6002 (N_6002,N_3223,N_4401);
nand U6003 (N_6003,N_3646,N_3471);
or U6004 (N_6004,N_3448,N_4156);
nor U6005 (N_6005,N_3781,N_4398);
nand U6006 (N_6006,N_3245,N_5191);
nand U6007 (N_6007,N_4034,N_4120);
xor U6008 (N_6008,N_5563,N_5463);
xnor U6009 (N_6009,N_4744,N_3578);
nand U6010 (N_6010,N_3357,N_3704);
and U6011 (N_6011,N_3052,N_3869);
xor U6012 (N_6012,N_4041,N_3279);
xor U6013 (N_6013,N_4122,N_4070);
and U6014 (N_6014,N_4348,N_5949);
xnor U6015 (N_6015,N_3932,N_3118);
nand U6016 (N_6016,N_4805,N_5217);
nor U6017 (N_6017,N_5828,N_5484);
nor U6018 (N_6018,N_3626,N_4087);
or U6019 (N_6019,N_3572,N_3666);
and U6020 (N_6020,N_4172,N_5928);
nand U6021 (N_6021,N_5438,N_5332);
nor U6022 (N_6022,N_3239,N_4620);
nand U6023 (N_6023,N_4884,N_5729);
xor U6024 (N_6024,N_5140,N_4365);
or U6025 (N_6025,N_3622,N_3660);
nand U6026 (N_6026,N_4972,N_5870);
or U6027 (N_6027,N_4747,N_3332);
nor U6028 (N_6028,N_5139,N_5104);
nor U6029 (N_6029,N_3485,N_3066);
or U6030 (N_6030,N_4859,N_5344);
xor U6031 (N_6031,N_3679,N_4947);
nand U6032 (N_6032,N_3786,N_5397);
xor U6033 (N_6033,N_4180,N_4424);
xnor U6034 (N_6034,N_3888,N_4425);
nand U6035 (N_6035,N_4066,N_3136);
and U6036 (N_6036,N_4831,N_5406);
nand U6037 (N_6037,N_4223,N_3717);
or U6038 (N_6038,N_4691,N_4543);
and U6039 (N_6039,N_4104,N_3008);
or U6040 (N_6040,N_4519,N_5527);
and U6041 (N_6041,N_4073,N_5181);
or U6042 (N_6042,N_4832,N_5437);
and U6043 (N_6043,N_4042,N_5877);
and U6044 (N_6044,N_5070,N_3913);
nand U6045 (N_6045,N_5500,N_3397);
xnor U6046 (N_6046,N_3810,N_5987);
and U6047 (N_6047,N_4731,N_5162);
and U6048 (N_6048,N_3518,N_3460);
xor U6049 (N_6049,N_4265,N_5091);
or U6050 (N_6050,N_3632,N_5557);
nand U6051 (N_6051,N_3105,N_5746);
nand U6052 (N_6052,N_5316,N_5938);
nor U6053 (N_6053,N_4175,N_3647);
or U6054 (N_6054,N_5416,N_3957);
and U6055 (N_6055,N_3442,N_4804);
nand U6056 (N_6056,N_3431,N_4877);
and U6057 (N_6057,N_3723,N_5363);
or U6058 (N_6058,N_5743,N_3211);
or U6059 (N_6059,N_3251,N_3944);
xor U6060 (N_6060,N_3611,N_3173);
nand U6061 (N_6061,N_4726,N_5808);
or U6062 (N_6062,N_3589,N_5055);
nand U6063 (N_6063,N_3979,N_3090);
and U6064 (N_6064,N_3691,N_5822);
or U6065 (N_6065,N_5999,N_5408);
and U6066 (N_6066,N_4625,N_3829);
xor U6067 (N_6067,N_3734,N_4355);
nand U6068 (N_6068,N_3452,N_5932);
and U6069 (N_6069,N_3694,N_5710);
or U6070 (N_6070,N_3686,N_4976);
nand U6071 (N_6071,N_4513,N_3566);
nand U6072 (N_6072,N_5789,N_4289);
and U6073 (N_6073,N_4718,N_4719);
xnor U6074 (N_6074,N_4183,N_3182);
nor U6075 (N_6075,N_5208,N_5649);
and U6076 (N_6076,N_4422,N_4141);
nand U6077 (N_6077,N_3100,N_4126);
nor U6078 (N_6078,N_4303,N_4944);
or U6079 (N_6079,N_5769,N_3721);
nand U6080 (N_6080,N_4908,N_5741);
xor U6081 (N_6081,N_3826,N_3109);
nor U6082 (N_6082,N_3355,N_4788);
or U6083 (N_6083,N_5018,N_3633);
and U6084 (N_6084,N_3127,N_5414);
xor U6085 (N_6085,N_3305,N_5767);
xor U6086 (N_6086,N_3583,N_5687);
or U6087 (N_6087,N_4338,N_3492);
and U6088 (N_6088,N_4394,N_4538);
nand U6089 (N_6089,N_4190,N_3561);
or U6090 (N_6090,N_3710,N_4678);
xnor U6091 (N_6091,N_5155,N_4061);
or U6092 (N_6092,N_4294,N_4400);
or U6093 (N_6093,N_4351,N_4517);
and U6094 (N_6094,N_3901,N_3338);
and U6095 (N_6095,N_3454,N_3013);
nor U6096 (N_6096,N_5787,N_4943);
xnor U6097 (N_6097,N_4373,N_4029);
and U6098 (N_6098,N_3068,N_5977);
nor U6099 (N_6099,N_5296,N_4453);
and U6100 (N_6100,N_3994,N_5176);
or U6101 (N_6101,N_5660,N_5528);
and U6102 (N_6102,N_3323,N_3653);
xor U6103 (N_6103,N_5967,N_3837);
and U6104 (N_6104,N_3814,N_5809);
xor U6105 (N_6105,N_4282,N_5841);
nor U6106 (N_6106,N_5616,N_5830);
and U6107 (N_6107,N_4579,N_5412);
or U6108 (N_6108,N_5177,N_4015);
nand U6109 (N_6109,N_3474,N_4550);
or U6110 (N_6110,N_5538,N_4032);
nand U6111 (N_6111,N_3522,N_4497);
xnor U6112 (N_6112,N_3190,N_4562);
nand U6113 (N_6113,N_3123,N_5756);
nand U6114 (N_6114,N_4802,N_3639);
and U6115 (N_6115,N_5119,N_4433);
or U6116 (N_6116,N_3350,N_3965);
nand U6117 (N_6117,N_4227,N_3387);
nand U6118 (N_6118,N_3733,N_3379);
xnor U6119 (N_6119,N_4336,N_5387);
and U6120 (N_6120,N_4257,N_4464);
xnor U6121 (N_6121,N_4876,N_4926);
and U6122 (N_6122,N_3648,N_5219);
and U6123 (N_6123,N_5936,N_5630);
xor U6124 (N_6124,N_3971,N_4417);
and U6125 (N_6125,N_4815,N_3069);
and U6126 (N_6126,N_5546,N_3946);
xnor U6127 (N_6127,N_3416,N_5613);
xor U6128 (N_6128,N_3549,N_4604);
or U6129 (N_6129,N_3598,N_4060);
nor U6130 (N_6130,N_5581,N_3966);
and U6131 (N_6131,N_3226,N_4954);
nand U6132 (N_6132,N_5835,N_4885);
xnor U6133 (N_6133,N_4165,N_3497);
xnor U6134 (N_6134,N_4164,N_5714);
and U6135 (N_6135,N_5893,N_3865);
or U6136 (N_6136,N_5206,N_3158);
or U6137 (N_6137,N_3774,N_3699);
xor U6138 (N_6138,N_5591,N_5167);
nand U6139 (N_6139,N_3800,N_4204);
xor U6140 (N_6140,N_3895,N_5939);
xor U6141 (N_6141,N_5873,N_3914);
xnor U6142 (N_6142,N_3541,N_4529);
or U6143 (N_6143,N_4749,N_3651);
and U6144 (N_6144,N_4912,N_3010);
xor U6145 (N_6145,N_5857,N_4046);
nor U6146 (N_6146,N_3712,N_4423);
nor U6147 (N_6147,N_3934,N_5313);
xnor U6148 (N_6148,N_3511,N_5816);
or U6149 (N_6149,N_5554,N_4784);
nor U6150 (N_6150,N_3358,N_4961);
xnor U6151 (N_6151,N_3517,N_5106);
xor U6152 (N_6152,N_4469,N_4866);
nor U6153 (N_6153,N_4897,N_3117);
or U6154 (N_6154,N_3614,N_4629);
or U6155 (N_6155,N_5559,N_4710);
xnor U6156 (N_6156,N_5023,N_3879);
nor U6157 (N_6157,N_3726,N_4331);
nor U6158 (N_6158,N_4531,N_4483);
xnor U6159 (N_6159,N_4435,N_5671);
xnor U6160 (N_6160,N_5537,N_5573);
xor U6161 (N_6161,N_3303,N_3619);
nor U6162 (N_6162,N_3976,N_3991);
xnor U6163 (N_6163,N_5876,N_5282);
or U6164 (N_6164,N_3907,N_3133);
nand U6165 (N_6165,N_3776,N_3748);
or U6166 (N_6166,N_5589,N_5317);
and U6167 (N_6167,N_3186,N_4794);
nand U6168 (N_6168,N_3390,N_5024);
nand U6169 (N_6169,N_5829,N_4148);
nor U6170 (N_6170,N_4411,N_4219);
and U6171 (N_6171,N_5275,N_4632);
and U6172 (N_6172,N_3145,N_3084);
nand U6173 (N_6173,N_5824,N_4208);
xnor U6174 (N_6174,N_4369,N_4430);
or U6175 (N_6175,N_4891,N_5742);
nor U6176 (N_6176,N_4623,N_3533);
and U6177 (N_6177,N_3669,N_5233);
or U6178 (N_6178,N_3828,N_3571);
and U6179 (N_6179,N_3709,N_3176);
or U6180 (N_6180,N_4648,N_5389);
nor U6181 (N_6181,N_5585,N_5875);
nand U6182 (N_6182,N_4697,N_5226);
nor U6183 (N_6183,N_5855,N_5840);
or U6184 (N_6184,N_3366,N_5530);
nor U6185 (N_6185,N_5518,N_3846);
nand U6186 (N_6186,N_4198,N_5436);
nor U6187 (N_6187,N_5636,N_3383);
nor U6188 (N_6188,N_5600,N_3349);
nand U6189 (N_6189,N_5948,N_3085);
nand U6190 (N_6190,N_3188,N_4651);
nand U6191 (N_6191,N_3806,N_4935);
or U6192 (N_6192,N_4207,N_4149);
xnor U6193 (N_6193,N_3220,N_5187);
and U6194 (N_6194,N_5804,N_4268);
and U6195 (N_6195,N_4048,N_5826);
or U6196 (N_6196,N_3322,N_4676);
nand U6197 (N_6197,N_3247,N_5066);
nand U6198 (N_6198,N_5077,N_4192);
nor U6199 (N_6199,N_3335,N_4978);
and U6200 (N_6200,N_5593,N_5674);
nand U6201 (N_6201,N_4572,N_3990);
nor U6202 (N_6202,N_4376,N_5921);
nor U6203 (N_6203,N_3419,N_5166);
or U6204 (N_6204,N_4037,N_5353);
or U6205 (N_6205,N_5516,N_4386);
and U6206 (N_6206,N_3667,N_3797);
nor U6207 (N_6207,N_5421,N_4931);
nor U6208 (N_6208,N_5862,N_3071);
or U6209 (N_6209,N_4594,N_4283);
nor U6210 (N_6210,N_5307,N_3605);
nand U6211 (N_6211,N_4459,N_5793);
nand U6212 (N_6212,N_4610,N_4526);
nor U6213 (N_6213,N_4793,N_5844);
nor U6214 (N_6214,N_5570,N_5485);
nand U6215 (N_6215,N_3447,N_5403);
nand U6216 (N_6216,N_3627,N_3317);
nor U6217 (N_6217,N_3843,N_3097);
xnor U6218 (N_6218,N_4184,N_3370);
and U6219 (N_6219,N_3139,N_4878);
or U6220 (N_6220,N_4515,N_3036);
nand U6221 (N_6221,N_3950,N_4635);
xor U6222 (N_6222,N_5053,N_4860);
and U6223 (N_6223,N_5293,N_4672);
nand U6224 (N_6224,N_3925,N_3249);
nand U6225 (N_6225,N_4704,N_5638);
nor U6226 (N_6226,N_4335,N_3181);
or U6227 (N_6227,N_3854,N_5618);
and U6228 (N_6228,N_3293,N_5280);
xor U6229 (N_6229,N_5254,N_4468);
xnor U6230 (N_6230,N_4687,N_3311);
nand U6231 (N_6231,N_5351,N_5452);
xnor U6232 (N_6232,N_3902,N_3830);
and U6233 (N_6233,N_4103,N_3201);
xnor U6234 (N_6234,N_4232,N_3009);
xor U6235 (N_6235,N_4450,N_5846);
nand U6236 (N_6236,N_5654,N_4605);
xor U6237 (N_6237,N_5045,N_3987);
nor U6238 (N_6238,N_3788,N_4167);
nor U6239 (N_6239,N_4668,N_3599);
nand U6240 (N_6240,N_5776,N_5161);
or U6241 (N_6241,N_4174,N_4383);
or U6242 (N_6242,N_5080,N_3006);
xnor U6243 (N_6243,N_3132,N_5134);
and U6244 (N_6244,N_5805,N_3369);
or U6245 (N_6245,N_3114,N_4153);
nor U6246 (N_6246,N_5661,N_4746);
and U6247 (N_6247,N_4823,N_5821);
xnor U6248 (N_6248,N_5605,N_4843);
and U6249 (N_6249,N_5614,N_3345);
xor U6250 (N_6250,N_5922,N_5553);
xor U6251 (N_6251,N_5994,N_3574);
nor U6252 (N_6252,N_5050,N_3267);
and U6253 (N_6253,N_5243,N_4218);
nand U6254 (N_6254,N_3041,N_3790);
and U6255 (N_6255,N_3138,N_3412);
nor U6256 (N_6256,N_4317,N_5753);
xor U6257 (N_6257,N_5791,N_5272);
or U6258 (N_6258,N_3628,N_5175);
nor U6259 (N_6259,N_4662,N_3894);
or U6260 (N_6260,N_4762,N_5951);
nor U6261 (N_6261,N_4086,N_3656);
nor U6262 (N_6262,N_4052,N_5825);
nand U6263 (N_6263,N_4770,N_4503);
or U6264 (N_6264,N_4971,N_3706);
or U6265 (N_6265,N_5321,N_4500);
and U6266 (N_6266,N_5642,N_5146);
or U6267 (N_6267,N_4911,N_4124);
xor U6268 (N_6268,N_4945,N_5298);
xor U6269 (N_6269,N_3001,N_3613);
xnor U6270 (N_6270,N_4764,N_3811);
nand U6271 (N_6271,N_3343,N_4590);
and U6272 (N_6272,N_3764,N_3450);
xnor U6273 (N_6273,N_4627,N_4110);
or U6274 (N_6274,N_5330,N_5535);
and U6275 (N_6275,N_4301,N_3867);
xor U6276 (N_6276,N_5430,N_4137);
nand U6277 (N_6277,N_5702,N_5078);
nor U6278 (N_6278,N_4688,N_5690);
and U6279 (N_6279,N_3208,N_5507);
nand U6280 (N_6280,N_5428,N_5035);
xor U6281 (N_6281,N_4951,N_4785);
and U6282 (N_6282,N_3803,N_5878);
nand U6283 (N_6283,N_5964,N_3877);
and U6284 (N_6284,N_4119,N_3047);
nand U6285 (N_6285,N_4895,N_3889);
nand U6286 (N_6286,N_3883,N_3844);
xnor U6287 (N_6287,N_5902,N_3773);
nand U6288 (N_6288,N_3584,N_4454);
xor U6289 (N_6289,N_4616,N_4963);
nor U6290 (N_6290,N_3213,N_4980);
and U6291 (N_6291,N_4089,N_3935);
nand U6292 (N_6292,N_4892,N_4291);
nor U6293 (N_6293,N_4559,N_3972);
and U6294 (N_6294,N_5465,N_5621);
nand U6295 (N_6295,N_3853,N_5195);
and U6296 (N_6296,N_5668,N_3791);
and U6297 (N_6297,N_3489,N_5739);
xor U6298 (N_6298,N_5099,N_3552);
and U6299 (N_6299,N_4750,N_4899);
or U6300 (N_6300,N_4660,N_4667);
or U6301 (N_6301,N_4161,N_4131);
nand U6302 (N_6302,N_4539,N_3559);
or U6303 (N_6303,N_5314,N_4979);
xor U6304 (N_6304,N_4838,N_3775);
xnor U6305 (N_6305,N_3538,N_5092);
xnor U6306 (N_6306,N_4690,N_4281);
nand U6307 (N_6307,N_5192,N_5283);
and U6308 (N_6308,N_3816,N_4603);
xor U6309 (N_6309,N_4756,N_5622);
nor U6310 (N_6310,N_4540,N_4202);
xor U6311 (N_6311,N_4998,N_5235);
and U6312 (N_6312,N_5634,N_4679);
nand U6313 (N_6313,N_4507,N_4363);
nor U6314 (N_6314,N_3250,N_5026);
nor U6315 (N_6315,N_3556,N_5778);
nand U6316 (N_6316,N_4178,N_3785);
nand U6317 (N_6317,N_4906,N_3360);
or U6318 (N_6318,N_3286,N_5407);
nand U6319 (N_6319,N_4845,N_5189);
or U6320 (N_6320,N_5856,N_3600);
or U6321 (N_6321,N_5108,N_4134);
nand U6322 (N_6322,N_4206,N_4587);
and U6323 (N_6323,N_3755,N_5497);
nor U6324 (N_6324,N_3595,N_3000);
or U6325 (N_6325,N_3752,N_3103);
nand U6326 (N_6326,N_3858,N_4914);
nand U6327 (N_6327,N_4586,N_3168);
nand U6328 (N_6328,N_5366,N_5914);
xnor U6329 (N_6329,N_4533,N_5980);
and U6330 (N_6330,N_4229,N_5502);
and U6331 (N_6331,N_3253,N_5960);
nor U6332 (N_6332,N_4220,N_4777);
and U6333 (N_6333,N_3409,N_4921);
nor U6334 (N_6334,N_4506,N_4534);
or U6335 (N_6335,N_5717,N_4846);
nor U6336 (N_6336,N_3104,N_4732);
and U6337 (N_6337,N_5771,N_4078);
nand U6338 (N_6338,N_5115,N_5594);
nor U6339 (N_6339,N_5700,N_5576);
and U6340 (N_6340,N_5625,N_3062);
nand U6341 (N_6341,N_5451,N_3662);
nand U6342 (N_6342,N_5820,N_5101);
xor U6343 (N_6343,N_4693,N_5386);
nand U6344 (N_6344,N_3840,N_3420);
and U6345 (N_6345,N_3608,N_3822);
or U6346 (N_6346,N_5764,N_5168);
nor U6347 (N_6347,N_5394,N_5063);
xnor U6348 (N_6348,N_3418,N_5874);
and U6349 (N_6349,N_5505,N_4551);
nand U6350 (N_6350,N_3098,N_4940);
nor U6351 (N_6351,N_4640,N_4495);
xor U6352 (N_6352,N_3330,N_3524);
and U6353 (N_6353,N_3316,N_4946);
or U6354 (N_6354,N_5940,N_3274);
nor U6355 (N_6355,N_5930,N_5385);
xnor U6356 (N_6356,N_3607,N_4847);
nor U6357 (N_6357,N_4484,N_5650);
nand U6358 (N_6358,N_4905,N_4695);
xor U6359 (N_6359,N_5443,N_4582);
and U6360 (N_6360,N_4498,N_3027);
nand U6361 (N_6361,N_3967,N_4516);
nor U6362 (N_6362,N_3546,N_4669);
xnor U6363 (N_6363,N_4372,N_3737);
nor U6364 (N_6364,N_3807,N_3273);
nand U6365 (N_6365,N_4439,N_3378);
xor U6366 (N_6366,N_5477,N_3395);
nand U6367 (N_6367,N_3348,N_4353);
nand U6368 (N_6368,N_3093,N_4983);
xnor U6369 (N_6369,N_4975,N_5689);
and U6370 (N_6370,N_3164,N_5584);
nand U6371 (N_6371,N_3729,N_4340);
or U6372 (N_6372,N_5496,N_4647);
and U6373 (N_6373,N_4556,N_5383);
nor U6374 (N_6374,N_3727,N_4739);
nand U6375 (N_6375,N_4377,N_5399);
nand U6376 (N_6376,N_5304,N_5241);
nand U6377 (N_6377,N_3445,N_3115);
xor U6378 (N_6378,N_5229,N_3714);
nor U6379 (N_6379,N_4478,N_4269);
nand U6380 (N_6380,N_5453,N_5464);
xor U6381 (N_6381,N_4729,N_3024);
nor U6382 (N_6382,N_3403,N_5694);
and U6383 (N_6383,N_3232,N_5072);
and U6384 (N_6384,N_4033,N_5156);
xor U6385 (N_6385,N_4828,N_3275);
xor U6386 (N_6386,N_5785,N_5046);
or U6387 (N_6387,N_3570,N_3421);
xor U6388 (N_6388,N_4881,N_3515);
xnor U6389 (N_6389,N_4001,N_3495);
nor U6390 (N_6390,N_3095,N_4112);
nand U6391 (N_6391,N_4460,N_3096);
nand U6392 (N_6392,N_5815,N_4455);
xor U6393 (N_6393,N_5564,N_5112);
and U6394 (N_6394,N_5867,N_3110);
or U6395 (N_6395,N_5807,N_3030);
xnor U6396 (N_6396,N_3212,N_5864);
nand U6397 (N_6397,N_4284,N_3745);
xnor U6398 (N_6398,N_4028,N_5398);
xor U6399 (N_6399,N_3149,N_5409);
nor U6400 (N_6400,N_5923,N_3225);
xor U6401 (N_6401,N_3540,N_3817);
nand U6402 (N_6402,N_4090,N_5952);
nand U6403 (N_6403,N_4391,N_4548);
and U6404 (N_6404,N_3494,N_3684);
nor U6405 (N_6405,N_4673,N_3919);
or U6406 (N_6406,N_5655,N_3028);
nor U6407 (N_6407,N_5747,N_4263);
nor U6408 (N_6408,N_3077,N_3405);
nand U6409 (N_6409,N_5859,N_4054);
nand U6410 (N_6410,N_5277,N_4143);
or U6411 (N_6411,N_3962,N_3458);
nand U6412 (N_6412,N_4482,N_5014);
or U6413 (N_6413,N_4151,N_5598);
xor U6414 (N_6414,N_5185,N_4308);
nor U6415 (N_6415,N_5542,N_5531);
xnor U6416 (N_6416,N_3980,N_3500);
or U6417 (N_6417,N_4009,N_5419);
nand U6418 (N_6418,N_5456,N_5377);
or U6419 (N_6419,N_4922,N_5944);
xor U6420 (N_6420,N_5138,N_3683);
xor U6421 (N_6421,N_4395,N_3779);
nor U6422 (N_6422,N_4321,N_3525);
nand U6423 (N_6423,N_4129,N_3059);
xnor U6424 (N_6424,N_3736,N_3368);
and U6425 (N_6425,N_4545,N_5849);
or U6426 (N_6426,N_3798,N_3038);
or U6427 (N_6427,N_4871,N_5757);
nand U6428 (N_6428,N_4212,N_3411);
xnor U6429 (N_6429,N_5211,N_5222);
and U6430 (N_6430,N_4343,N_3528);
nor U6431 (N_6431,N_5560,N_4795);
nor U6432 (N_6432,N_3342,N_3918);
and U6433 (N_6433,N_5918,N_5094);
nand U6434 (N_6434,N_5699,N_3490);
or U6435 (N_6435,N_5533,N_3986);
and U6436 (N_6436,N_3591,N_4707);
or U6437 (N_6437,N_5567,N_4547);
and U6438 (N_6438,N_5462,N_4568);
nand U6439 (N_6439,N_5566,N_4599);
nor U6440 (N_6440,N_3695,N_3820);
nor U6441 (N_6441,N_5262,N_4168);
nand U6442 (N_6442,N_4230,N_5020);
nand U6443 (N_6443,N_5736,N_4532);
and U6444 (N_6444,N_4201,N_3526);
xnor U6445 (N_6445,N_3380,N_4919);
nor U6446 (N_6446,N_3917,N_3464);
nor U6447 (N_6447,N_3657,N_3292);
nor U6448 (N_6448,N_3262,N_3496);
nand U6449 (N_6449,N_5240,N_4243);
nor U6450 (N_6450,N_5693,N_5158);
nor U6451 (N_6451,N_5904,N_4924);
and U6452 (N_6452,N_4580,N_4622);
nand U6453 (N_6453,N_3429,N_3997);
nand U6454 (N_6454,N_5360,N_4682);
nand U6455 (N_6455,N_5220,N_3417);
or U6456 (N_6456,N_5556,N_4114);
and U6457 (N_6457,N_5745,N_3032);
xor U6458 (N_6458,N_4182,N_3285);
nor U6459 (N_6459,N_3243,N_5149);
and U6460 (N_6460,N_4988,N_5637);
or U6461 (N_6461,N_4789,N_3111);
or U6462 (N_6462,N_4297,N_5684);
nor U6463 (N_6463,N_3277,N_5039);
nor U6464 (N_6464,N_4790,N_3831);
nor U6465 (N_6465,N_4237,N_5534);
nand U6466 (N_6466,N_4479,N_5439);
nor U6467 (N_6467,N_5632,N_3075);
nor U6468 (N_6468,N_3035,N_5494);
and U6469 (N_6469,N_5415,N_5706);
xnor U6470 (N_6470,N_4609,N_3824);
and U6471 (N_6471,N_3446,N_4429);
and U6472 (N_6472,N_3943,N_3931);
nand U6473 (N_6473,N_5230,N_4489);
and U6474 (N_6474,N_4684,N_5881);
nor U6475 (N_6475,N_3007,N_5264);
xor U6476 (N_6476,N_5159,N_4159);
or U6477 (N_6477,N_4990,N_5482);
or U6478 (N_6478,N_5052,N_4490);
nand U6479 (N_6479,N_5998,N_5544);
xnor U6480 (N_6480,N_3762,N_5603);
nand U6481 (N_6481,N_5498,N_3839);
nand U6482 (N_6482,N_4442,N_3542);
nor U6483 (N_6483,N_3473,N_3974);
nand U6484 (N_6484,N_4366,N_3080);
xnor U6485 (N_6485,N_4014,N_3851);
xnor U6486 (N_6486,N_4638,N_4653);
nand U6487 (N_6487,N_4840,N_3025);
nand U6488 (N_6488,N_5493,N_4325);
or U6489 (N_6489,N_5312,N_5459);
xnor U6490 (N_6490,N_5044,N_5562);
or U6491 (N_6491,N_3910,N_5906);
or U6492 (N_6492,N_4819,N_4745);
xor U6493 (N_6493,N_5431,N_4318);
and U6494 (N_6494,N_3823,N_3716);
nor U6495 (N_6495,N_4867,N_4007);
or U6496 (N_6496,N_3166,N_4967);
or U6497 (N_6497,N_5629,N_5597);
nor U6498 (N_6498,N_3969,N_4592);
and U6499 (N_6499,N_5157,N_4520);
xnor U6500 (N_6500,N_3845,N_5688);
nand U6501 (N_6501,N_3711,N_4743);
or U6502 (N_6502,N_4692,N_5708);
nand U6503 (N_6503,N_4407,N_3558);
nand U6504 (N_6504,N_3470,N_4512);
or U6505 (N_6505,N_4862,N_5255);
and U6506 (N_6506,N_3198,N_4728);
or U6507 (N_6507,N_5372,N_3904);
nand U6508 (N_6508,N_3941,N_4277);
xor U6509 (N_6509,N_3240,N_5996);
xnor U6510 (N_6510,N_5267,N_3119);
xnor U6511 (N_6511,N_5132,N_4140);
or U6512 (N_6512,N_3655,N_4476);
xor U6513 (N_6513,N_4511,N_4494);
and U6514 (N_6514,N_5579,N_5961);
and U6515 (N_6515,N_3328,N_4273);
nand U6516 (N_6516,N_3685,N_5810);
xor U6517 (N_6517,N_5338,N_5733);
xor U6518 (N_6518,N_3909,N_4522);
nor U6519 (N_6519,N_4071,N_3406);
and U6520 (N_6520,N_5958,N_4013);
nor U6521 (N_6521,N_3720,N_4549);
xor U6522 (N_6522,N_5997,N_4286);
nor U6523 (N_6523,N_5448,N_3521);
nor U6524 (N_6524,N_3017,N_5354);
or U6525 (N_6525,N_5165,N_5768);
and U6526 (N_6526,N_3926,N_5201);
and U6527 (N_6527,N_4820,N_3058);
nand U6528 (N_6528,N_3064,N_3433);
and U6529 (N_6529,N_5216,N_5551);
nand U6530 (N_6530,N_4280,N_3270);
nand U6531 (N_6531,N_3435,N_5691);
and U6532 (N_6532,N_4896,N_3130);
nand U6533 (N_6533,N_5631,N_3386);
and U6534 (N_6534,N_5574,N_4199);
or U6535 (N_6535,N_4863,N_3291);
xor U6536 (N_6536,N_4446,N_5853);
nor U6537 (N_6537,N_3805,N_4600);
and U6538 (N_6538,N_4157,N_5831);
xor U6539 (N_6539,N_5225,N_4583);
nand U6540 (N_6540,N_5607,N_5141);
or U6541 (N_6541,N_4960,N_3165);
nor U6542 (N_6542,N_4397,N_3863);
nand U6543 (N_6543,N_3012,N_5111);
nand U6544 (N_6544,N_5103,N_5990);
nand U6545 (N_6545,N_4171,N_5885);
or U6546 (N_6546,N_5107,N_3057);
nor U6547 (N_6547,N_4613,N_3930);
nor U6548 (N_6548,N_5966,N_4855);
xor U6549 (N_6549,N_5117,N_3361);
nor U6550 (N_6550,N_5400,N_4894);
and U6551 (N_6551,N_4883,N_4527);
xor U6552 (N_6552,N_4345,N_4426);
and U6553 (N_6553,N_5009,N_5775);
nand U6554 (N_6554,N_4072,N_3134);
and U6555 (N_6555,N_4510,N_3276);
xor U6556 (N_6556,N_3048,N_4671);
or U6557 (N_6557,N_3185,N_5889);
and U6558 (N_6558,N_3441,N_4518);
and U6559 (N_6559,N_4771,N_5483);
and U6560 (N_6560,N_4864,N_3738);
or U6561 (N_6561,N_3638,N_3229);
nand U6562 (N_6562,N_5954,N_4188);
and U6563 (N_6563,N_3271,N_3975);
or U6564 (N_6564,N_4323,N_3650);
or U6565 (N_6565,N_5118,N_3642);
xor U6566 (N_6566,N_4231,N_3749);
or U6567 (N_6567,N_5268,N_3604);
nand U6568 (N_6568,N_3258,N_5210);
nor U6569 (N_6569,N_3167,N_3312);
xor U6570 (N_6570,N_3880,N_5982);
and U6571 (N_6571,N_5059,N_3688);
nor U6572 (N_6572,N_5539,N_5334);
nor U6573 (N_6573,N_3857,N_3766);
xnor U6574 (N_6574,N_5279,N_3743);
nand U6575 (N_6575,N_4370,N_4637);
nand U6576 (N_6576,N_4965,N_3767);
nand U6577 (N_6577,N_5879,N_4062);
and U6578 (N_6578,N_4711,N_4696);
xnor U6579 (N_6579,N_3227,N_5510);
or U6580 (N_6580,N_5418,N_4093);
xnor U6581 (N_6581,N_5989,N_5646);
or U6582 (N_6582,N_3480,N_4514);
and U6583 (N_6583,N_3375,N_4456);
nor U6584 (N_6584,N_4999,N_3537);
nand U6585 (N_6585,N_4560,N_3278);
and U6586 (N_6586,N_4591,N_3915);
and U6587 (N_6587,N_4251,N_4923);
and U6588 (N_6588,N_4111,N_3875);
nor U6589 (N_6589,N_3970,N_3770);
xor U6590 (N_6590,N_4984,N_5281);
xnor U6591 (N_6591,N_4239,N_3757);
nor U6592 (N_6592,N_5350,N_4578);
xnor U6593 (N_6593,N_5900,N_4385);
or U6594 (N_6594,N_5405,N_5340);
and U6595 (N_6595,N_5790,N_4630);
xor U6596 (N_6596,N_5703,N_5325);
nor U6597 (N_6597,N_4612,N_4333);
and U6598 (N_6598,N_4811,N_5152);
nor U6599 (N_6599,N_4026,N_3183);
nand U6600 (N_6600,N_4933,N_5899);
xor U6601 (N_6601,N_4856,N_5081);
xor U6602 (N_6602,N_4374,N_4160);
nor U6603 (N_6603,N_3206,N_4035);
and U6604 (N_6604,N_4589,N_4689);
xor U6605 (N_6605,N_5223,N_3750);
or U6606 (N_6606,N_4368,N_4234);
xor U6607 (N_6607,N_5097,N_4387);
nor U6608 (N_6608,N_3624,N_4102);
or U6609 (N_6609,N_5937,N_4403);
xor U6610 (N_6610,N_5170,N_4974);
nand U6611 (N_6611,N_5988,N_5772);
nand U6612 (N_6612,N_5147,N_5365);
nand U6613 (N_6613,N_4705,N_5245);
xnor U6614 (N_6614,N_3550,N_3725);
and U6615 (N_6615,N_5752,N_4523);
nand U6616 (N_6616,N_3488,N_3801);
and U6617 (N_6617,N_5411,N_3512);
nor U6618 (N_6618,N_5858,N_4741);
xnor U6619 (N_6619,N_4763,N_4631);
xnor U6620 (N_6620,N_5737,N_4108);
nand U6621 (N_6621,N_3299,N_5872);
nor U6622 (N_6622,N_3649,N_3177);
nand U6623 (N_6623,N_3324,N_3336);
xnor U6624 (N_6624,N_4169,N_3087);
nor U6625 (N_6625,N_3477,N_3171);
nor U6626 (N_6626,N_4939,N_4886);
nor U6627 (N_6627,N_4065,N_3437);
xnor U6628 (N_6628,N_3681,N_3841);
nor U6629 (N_6629,N_5120,N_3590);
or U6630 (N_6630,N_3783,N_5818);
or U6631 (N_6631,N_3596,N_3180);
nand U6632 (N_6632,N_4909,N_4727);
xnor U6633 (N_6633,N_3754,N_4044);
or U6634 (N_6634,N_5367,N_3548);
or U6635 (N_6635,N_5231,N_4278);
nor U6636 (N_6636,N_5586,N_4851);
and U6637 (N_6637,N_4247,N_3099);
nor U6638 (N_6638,N_5588,N_4787);
or U6639 (N_6639,N_3881,N_4782);
nand U6640 (N_6640,N_3760,N_4964);
xnor U6641 (N_6641,N_5315,N_5543);
and U6642 (N_6642,N_5817,N_3493);
or U6643 (N_6643,N_5123,N_5643);
or U6644 (N_6644,N_5049,N_4197);
and U6645 (N_6645,N_5190,N_4254);
xor U6646 (N_6646,N_5273,N_4057);
nor U6647 (N_6647,N_4493,N_5524);
xnor U6648 (N_6648,N_3959,N_5200);
xor U6649 (N_6649,N_5128,N_5532);
xnor U6650 (N_6650,N_5204,N_5547);
and U6651 (N_6651,N_3415,N_4448);
nand U6652 (N_6652,N_5883,N_5186);
nand U6653 (N_6653,N_5748,N_5374);
or U6654 (N_6654,N_4786,N_3155);
and U6655 (N_6655,N_4869,N_4712);
nand U6656 (N_6656,N_3900,N_5555);
nand U6657 (N_6657,N_3731,N_4958);
or U6658 (N_6658,N_5056,N_5865);
or U6659 (N_6659,N_3742,N_3426);
nand U6660 (N_6660,N_5326,N_4393);
nand U6661 (N_6661,N_3664,N_3189);
or U6662 (N_6662,N_3116,N_5184);
nand U6663 (N_6663,N_5343,N_5796);
or U6664 (N_6664,N_5641,N_3992);
or U6665 (N_6665,N_5012,N_5331);
nand U6666 (N_6666,N_3718,N_5188);
nor U6667 (N_6667,N_4738,N_4101);
xnor U6668 (N_6668,N_3995,N_4723);
or U6669 (N_6669,N_5628,N_3923);
and U6670 (N_6670,N_4618,N_3313);
nor U6671 (N_6671,N_5011,N_3268);
xnor U6672 (N_6672,N_5000,N_3836);
nor U6673 (N_6673,N_5004,N_3623);
and U6674 (N_6674,N_4181,N_5067);
and U6675 (N_6675,N_5221,N_4991);
or U6676 (N_6676,N_4737,N_4801);
nor U6677 (N_6677,N_3234,N_3150);
xor U6678 (N_6678,N_3091,N_5721);
or U6679 (N_6679,N_3408,N_3385);
nand U6680 (N_6680,N_3747,N_3506);
nand U6681 (N_6681,N_3898,N_4275);
nor U6682 (N_6682,N_3389,N_3937);
nand U6683 (N_6683,N_4203,N_3351);
nor U6684 (N_6684,N_4959,N_5427);
and U6685 (N_6685,N_3086,N_4115);
nor U6686 (N_6686,N_3359,N_5725);
nor U6687 (N_6687,N_3294,N_5651);
xnor U6688 (N_6688,N_4887,N_4132);
nor U6689 (N_6689,N_5866,N_4434);
nor U6690 (N_6690,N_4818,N_3963);
and U6691 (N_6691,N_5986,N_5475);
nand U6692 (N_6692,N_3771,N_5583);
xnor U6693 (N_6693,N_4162,N_4038);
or U6694 (N_6694,N_5782,N_3238);
nor U6695 (N_6695,N_4722,N_4879);
and U6696 (N_6696,N_4797,N_5976);
nor U6697 (N_6697,N_4058,N_4621);
or U6698 (N_6698,N_3367,N_5238);
nand U6699 (N_6699,N_3510,N_3031);
nand U6700 (N_6700,N_4501,N_3033);
nand U6701 (N_6701,N_5461,N_3661);
and U6702 (N_6702,N_5234,N_4296);
nand U6703 (N_6703,N_5754,N_3475);
nor U6704 (N_6704,N_3698,N_5991);
xnor U6705 (N_6705,N_5288,N_5718);
and U6706 (N_6706,N_4177,N_4069);
nor U6707 (N_6707,N_5795,N_3159);
xor U6708 (N_6708,N_4643,N_4917);
nand U6709 (N_6709,N_3532,N_5837);
or U6710 (N_6710,N_5565,N_5309);
nand U6711 (N_6711,N_3265,N_5037);
or U6712 (N_6712,N_3065,N_5662);
xnor U6713 (N_6713,N_4270,N_3531);
or U6714 (N_6714,N_3719,N_5734);
nand U6715 (N_6715,N_5455,N_4463);
nor U6716 (N_6716,N_3434,N_4196);
and U6717 (N_6717,N_4814,N_5420);
nand U6718 (N_6718,N_5972,N_5061);
and U6719 (N_6719,N_5029,N_3353);
xor U6720 (N_6720,N_3670,N_3654);
nand U6721 (N_6721,N_3778,N_5709);
nand U6722 (N_6722,N_3248,N_4698);
nor U6723 (N_6723,N_5765,N_5890);
nor U6724 (N_6724,N_5569,N_5911);
or U6725 (N_6725,N_3363,N_4367);
nor U6726 (N_6726,N_5738,N_5263);
or U6727 (N_6727,N_5558,N_4626);
nor U6728 (N_6728,N_4903,N_4274);
or U6729 (N_6729,N_5898,N_3364);
and U6730 (N_6730,N_3592,N_5623);
nor U6731 (N_6731,N_3060,N_5571);
or U6732 (N_6732,N_3219,N_4299);
nand U6733 (N_6733,N_3874,N_3257);
and U6734 (N_6734,N_3847,N_5730);
nand U6735 (N_6735,N_3878,N_4645);
nor U6736 (N_6736,N_5143,N_3832);
or U6737 (N_6737,N_3061,N_5683);
nand U6738 (N_6738,N_4304,N_3621);
nand U6739 (N_6739,N_3451,N_4272);
nand U6740 (N_6740,N_3740,N_4019);
and U6741 (N_6741,N_4018,N_4077);
xor U6742 (N_6742,N_5968,N_5376);
nand U6743 (N_6743,N_4993,N_3281);
nor U6744 (N_6744,N_5287,N_4890);
and U6745 (N_6745,N_5659,N_4416);
nor U6746 (N_6746,N_4615,N_4471);
nor U6747 (N_6747,N_3214,N_5203);
or U6748 (N_6748,N_5673,N_4880);
or U6749 (N_6749,N_4873,N_3005);
or U6750 (N_6750,N_3465,N_4261);
nor U6751 (N_6751,N_4406,N_3905);
nor U6752 (N_6752,N_4870,N_4287);
nor U6753 (N_6753,N_4680,N_5017);
xnor U6754 (N_6754,N_4807,N_4195);
and U6755 (N_6755,N_5301,N_5347);
nand U6756 (N_6756,N_3516,N_3326);
nand U6757 (N_6757,N_5068,N_5740);
and U6758 (N_6758,N_4238,N_3637);
nand U6759 (N_6759,N_5919,N_4039);
nor U6760 (N_6760,N_5323,N_5575);
nor U6761 (N_6761,N_4686,N_5144);
or U6762 (N_6762,N_3050,N_3172);
nor U6763 (N_6763,N_4049,N_4106);
xnor U6764 (N_6764,N_4083,N_5148);
nor U6765 (N_6765,N_5511,N_4761);
nor U6766 (N_6766,N_4359,N_5060);
nand U6767 (N_6767,N_3019,N_3866);
and U6768 (N_6768,N_5062,N_4210);
or U6769 (N_6769,N_3308,N_5015);
xor U6770 (N_6770,N_5006,N_5744);
or U6771 (N_6771,N_5441,N_3112);
nand U6772 (N_6772,N_3302,N_5308);
or U6773 (N_6773,N_3479,N_3056);
or U6774 (N_6774,N_4295,N_4255);
and U6775 (N_6775,N_5252,N_4205);
or U6776 (N_6776,N_3301,N_5606);
nor U6777 (N_6777,N_5300,N_5154);
or U6778 (N_6778,N_4608,N_3588);
nand U6779 (N_6779,N_3453,N_3400);
nor U6780 (N_6780,N_3819,N_4258);
or U6781 (N_6781,N_5758,N_5031);
xor U6782 (N_6782,N_4409,N_5424);
nor U6783 (N_6783,N_5568,N_5897);
and U6784 (N_6784,N_3802,N_3241);
and U6785 (N_6785,N_3125,N_3565);
nor U6786 (N_6786,N_5665,N_4088);
xor U6787 (N_6787,N_4734,N_5085);
xnor U6788 (N_6788,N_3671,N_5652);
and U6789 (N_6789,N_4717,N_3722);
and U6790 (N_6790,N_4379,N_3759);
and U6791 (N_6791,N_4561,N_3481);
xor U6792 (N_6792,N_3947,N_5457);
or U6793 (N_6793,N_3427,N_3787);
nand U6794 (N_6794,N_3472,N_3668);
nand U6795 (N_6795,N_3751,N_3884);
xnor U6796 (N_6796,N_3443,N_3414);
xor U6797 (N_6797,N_3795,N_5695);
nand U6798 (N_6798,N_5054,N_3297);
and U6799 (N_6799,N_5269,N_5472);
and U6800 (N_6800,N_3088,N_5512);
and U6801 (N_6801,N_5292,N_5337);
xnor U6802 (N_6802,N_4155,N_3153);
and U6803 (N_6803,N_5611,N_5413);
xnor U6804 (N_6804,N_3612,N_3269);
or U6805 (N_6805,N_5032,N_4852);
and U6806 (N_6806,N_3993,N_4224);
or U6807 (N_6807,N_3804,N_5322);
and U6808 (N_6808,N_4027,N_4700);
xnor U6809 (N_6809,N_5202,N_3067);
nor U6810 (N_6810,N_3231,N_4607);
and U6811 (N_6811,N_3543,N_4384);
xnor U6812 (N_6812,N_3461,N_4328);
xor U6813 (N_6813,N_4339,N_5349);
nand U6814 (N_6814,N_4766,N_3491);
or U6815 (N_6815,N_5962,N_3978);
nor U6816 (N_6816,N_4185,N_5087);
or U6817 (N_6817,N_4721,N_5692);
or U6818 (N_6818,N_3659,N_3692);
xnor U6819 (N_6819,N_3021,N_5125);
xnor U6820 (N_6820,N_3004,N_5040);
nand U6821 (N_6821,N_5953,N_3424);
nor U6822 (N_6822,N_4674,N_4584);
and U6823 (N_6823,N_4043,N_3121);
nor U6824 (N_6824,N_3673,N_3053);
xnor U6825 (N_6825,N_4228,N_4146);
and U6826 (N_6826,N_3394,N_4012);
nor U6827 (N_6827,N_5514,N_4817);
xnor U6828 (N_6828,N_5719,N_5113);
and U6829 (N_6829,N_4798,N_5247);
xor U6830 (N_6830,N_3217,N_3794);
and U6831 (N_6831,N_4312,N_4096);
nor U6832 (N_6832,N_3161,N_5894);
nand U6833 (N_6833,N_4252,N_5284);
xnor U6834 (N_6834,N_5947,N_5712);
nand U6835 (N_6835,N_5069,N_5432);
nor U6836 (N_6836,N_5368,N_4213);
nor U6837 (N_6837,N_5100,N_5342);
nand U6838 (N_6838,N_4474,N_5871);
nand U6839 (N_6839,N_5978,N_5802);
or U6840 (N_6840,N_3676,N_5888);
xor U6841 (N_6841,N_5523,N_4677);
nand U6842 (N_6842,N_3911,N_5845);
or U6843 (N_6843,N_3184,N_3693);
nand U6844 (N_6844,N_4260,N_4715);
and U6845 (N_6845,N_5388,N_5207);
nand U6846 (N_6846,N_5716,N_4681);
nor U6847 (N_6847,N_4992,N_3896);
and U6848 (N_6848,N_4346,N_4542);
nand U6849 (N_6849,N_3428,N_5008);
nor U6850 (N_6850,N_3892,N_5028);
and U6851 (N_6851,N_3199,N_3499);
or U6852 (N_6852,N_5955,N_4822);
and U6853 (N_6853,N_5370,N_5848);
xor U6854 (N_6854,N_5329,N_4461);
xor U6855 (N_6855,N_3371,N_4389);
nor U6856 (N_6856,N_4068,N_5178);
and U6857 (N_6857,N_3306,N_4492);
nand U6858 (N_6858,N_3331,N_3523);
or U6859 (N_6859,N_5595,N_5811);
nor U6860 (N_6860,N_3929,N_4242);
nand U6861 (N_6861,N_4868,N_5380);
xnor U6862 (N_6862,N_4857,N_5965);
or U6863 (N_6863,N_3266,N_5929);
and U6864 (N_6864,N_5927,N_3401);
xor U6865 (N_6865,N_3746,N_4074);
xor U6866 (N_6866,N_5663,N_3603);
nand U6867 (N_6867,N_3527,N_5173);
xor U6868 (N_6868,N_4565,N_3756);
nor U6869 (N_6869,N_4315,N_4611);
or U6870 (N_6870,N_3634,N_4298);
and U6871 (N_6871,N_5895,N_4438);
and U6872 (N_6872,N_5615,N_3074);
xnor U6873 (N_6873,N_4349,N_5763);
and U6874 (N_6874,N_3347,N_4441);
nand U6875 (N_6875,N_5766,N_3903);
and U6876 (N_6876,N_3484,N_3782);
xor U6877 (N_6877,N_5781,N_5318);
and U6878 (N_6878,N_4186,N_4842);
and U6879 (N_6879,N_4769,N_5812);
nand U6880 (N_6880,N_5352,N_3885);
and U6881 (N_6881,N_5022,N_5256);
nand U6882 (N_6882,N_5854,N_5096);
or U6883 (N_6883,N_4701,N_4730);
nor U6884 (N_6884,N_4829,N_3289);
nand U6885 (N_6885,N_5130,N_3044);
xnor U6886 (N_6886,N_4193,N_4021);
nor U6887 (N_6887,N_5601,N_4428);
nor U6888 (N_6888,N_3715,N_4226);
and U6889 (N_6889,N_4853,N_4850);
nor U6890 (N_6890,N_4563,N_4316);
nor U6891 (N_6891,N_3852,N_4036);
or U6892 (N_6892,N_4176,N_4285);
xor U6893 (N_6893,N_5098,N_3730);
xor U6894 (N_6894,N_4699,N_4792);
and U6895 (N_6895,N_5290,N_3697);
or U6896 (N_6896,N_3587,N_5036);
and U6897 (N_6897,N_3402,N_3856);
nand U6898 (N_6898,N_3083,N_5517);
and U6899 (N_6899,N_4970,N_5838);
nand U6900 (N_6900,N_4758,N_4152);
or U6901 (N_6901,N_5707,N_3179);
and U6902 (N_6902,N_5102,N_4222);
or U6903 (N_6903,N_4830,N_5842);
or U6904 (N_6904,N_3625,N_3081);
or U6905 (N_6905,N_5667,N_4412);
and U6906 (N_6906,N_3796,N_5504);
or U6907 (N_6907,N_4005,N_4553);
xnor U6908 (N_6908,N_4685,N_5289);
xnor U6909 (N_6909,N_3629,N_4740);
or U6910 (N_6910,N_4938,N_4326);
nand U6911 (N_6911,N_5488,N_5850);
nor U6912 (N_6912,N_4874,N_5666);
xor U6913 (N_6913,N_3256,N_3861);
or U6914 (N_6914,N_5792,N_4451);
nand U6915 (N_6915,N_5679,N_4415);
or U6916 (N_6916,N_3107,N_3140);
xor U6917 (N_6917,N_3610,N_4803);
nor U6918 (N_6918,N_5525,N_5800);
nor U6919 (N_6919,N_4981,N_5105);
xnor U6920 (N_6920,N_5541,N_3601);
nand U6921 (N_6921,N_4045,N_5345);
or U6922 (N_6922,N_3063,N_3630);
and U6923 (N_6923,N_4447,N_4356);
or U6924 (N_6924,N_5909,N_5760);
xnor U6925 (N_6925,N_3393,N_5713);
nor U6926 (N_6926,N_3422,N_3777);
and U6927 (N_6927,N_5442,N_3151);
or U6928 (N_6928,N_5449,N_4396);
and U6929 (N_6929,N_3713,N_5058);
nor U6930 (N_6930,N_3576,N_5214);
and U6931 (N_6931,N_3799,N_4989);
nand U6932 (N_6932,N_3459,N_4810);
xor U6933 (N_6933,N_3162,N_4121);
nor U6934 (N_6934,N_3079,N_4310);
nand U6935 (N_6935,N_5305,N_5073);
xor U6936 (N_6936,N_3054,N_4982);
nor U6937 (N_6937,N_3055,N_3202);
and U6938 (N_6938,N_5306,N_4619);
or U6939 (N_6939,N_4521,N_5924);
and U6940 (N_6940,N_3842,N_4916);
or U6941 (N_6941,N_5794,N_4163);
nor U6942 (N_6942,N_4759,N_5896);
xnor U6943 (N_6943,N_4779,N_5508);
nor U6944 (N_6944,N_4655,N_5095);
nand U6945 (N_6945,N_3658,N_5382);
nand U6946 (N_6946,N_4329,N_4431);
and U6947 (N_6947,N_4941,N_3872);
xnor U6948 (N_6948,N_4486,N_5458);
nor U6949 (N_6949,N_5410,N_4528);
nand U6950 (N_6950,N_3761,N_3813);
nand U6951 (N_6951,N_3545,N_4187);
xor U6952 (N_6952,N_3131,N_5355);
and U6953 (N_6953,N_4996,N_3961);
and U6954 (N_6954,N_4646,N_3732);
and U6955 (N_6955,N_4307,N_3502);
nand U6956 (N_6956,N_3689,N_5362);
xnor U6957 (N_6957,N_4311,N_4929);
nor U6958 (N_6958,N_4378,N_3029);
nor U6959 (N_6959,N_4920,N_4091);
xnor U6960 (N_6960,N_3042,N_3101);
and U6961 (N_6961,N_5246,N_3928);
nor U6962 (N_6962,N_5797,N_5664);
and U6963 (N_6963,N_5346,N_3128);
or U6964 (N_6964,N_5596,N_3260);
nor U6965 (N_6965,N_3333,N_4443);
nand U6966 (N_6966,N_4889,N_3373);
xor U6967 (N_6967,N_3890,N_3772);
xnor U6968 (N_6968,N_3141,N_3672);
nor U6969 (N_6969,N_4342,N_5250);
nor U6970 (N_6970,N_5519,N_4948);
and U6971 (N_6971,N_5887,N_5209);
nand U6972 (N_6972,N_3708,N_4392);
and U6973 (N_6973,N_4708,N_4371);
nand U6974 (N_6974,N_5644,N_5599);
nor U6975 (N_6975,N_4320,N_5970);
and U6976 (N_6976,N_4457,N_4440);
and U6977 (N_6977,N_3618,N_4574);
nand U6978 (N_6978,N_5806,N_4658);
nand U6979 (N_6979,N_4735,N_5194);
or U6980 (N_6980,N_4957,N_4569);
xnor U6981 (N_6981,N_5869,N_3554);
and U6982 (N_6982,N_4898,N_5860);
and U6983 (N_6983,N_3675,N_5057);
nor U6984 (N_6984,N_3780,N_3868);
and U6985 (N_6985,N_4650,N_5434);
xnor U6986 (N_6986,N_3882,N_3924);
nor U6987 (N_6987,N_3037,N_3547);
or U6988 (N_6988,N_3339,N_4341);
nand U6989 (N_6989,N_4930,N_3825);
xor U6990 (N_6990,N_5974,N_4105);
nor U6991 (N_6991,N_5480,N_3244);
xnor U6992 (N_6992,N_4421,N_3620);
nor U6993 (N_6993,N_3020,N_3504);
xnor U6994 (N_6994,N_5973,N_4432);
or U6995 (N_6995,N_5925,N_5422);
nor U6996 (N_6996,N_3871,N_4973);
nand U6997 (N_6997,N_4834,N_4150);
xnor U6998 (N_6998,N_3120,N_3954);
nand U6999 (N_6999,N_4246,N_3985);
nand U7000 (N_7000,N_4390,N_5645);
and U7001 (N_7001,N_4598,N_4437);
xor U7002 (N_7002,N_4577,N_3187);
or U7003 (N_7003,N_3520,N_3254);
xnor U7004 (N_7004,N_4225,N_5552);
nor U7005 (N_7005,N_4781,N_5653);
nand U7006 (N_7006,N_5124,N_4020);
nand U7007 (N_7007,N_5799,N_3821);
nor U7008 (N_7008,N_3148,N_3912);
and U7009 (N_7009,N_4109,N_5227);
nor U7010 (N_7010,N_3462,N_5336);
or U7011 (N_7011,N_4768,N_4113);
nand U7012 (N_7012,N_3505,N_5487);
nor U7013 (N_7013,N_3530,N_3678);
xnor U7014 (N_7014,N_4347,N_4418);
or U7015 (N_7015,N_3376,N_3870);
nand U7016 (N_7016,N_4360,N_4010);
and U7017 (N_7017,N_5823,N_5843);
nand U7018 (N_7018,N_3864,N_5698);
and U7019 (N_7019,N_4900,N_4449);
and U7020 (N_7020,N_5359,N_4634);
xor U7021 (N_7021,N_3144,N_3082);
nor U7022 (N_7022,N_4714,N_4404);
or U7023 (N_7023,N_3812,N_5847);
or U7024 (N_7024,N_5393,N_4985);
xnor U7025 (N_7025,N_5770,N_4955);
nand U7026 (N_7026,N_5657,N_5722);
nor U7027 (N_7027,N_5460,N_5619);
or U7028 (N_7028,N_5813,N_3113);
nand U7029 (N_7029,N_5381,N_3739);
or U7030 (N_7030,N_5468,N_3315);
or U7031 (N_7031,N_4306,N_4773);
and U7032 (N_7032,N_3325,N_4465);
xnor U7033 (N_7033,N_4127,N_3014);
and U7034 (N_7034,N_3196,N_5476);
or U7035 (N_7035,N_5311,N_3597);
nand U7036 (N_7036,N_5620,N_5260);
nor U7037 (N_7037,N_5274,N_4470);
and U7038 (N_7038,N_3536,N_4067);
nor U7039 (N_7039,N_4666,N_3690);
xor U7040 (N_7040,N_5361,N_3951);
and U7041 (N_7041,N_5627,N_4191);
nand U7042 (N_7042,N_3002,N_5153);
xnor U7043 (N_7043,N_4952,N_3555);
nor U7044 (N_7044,N_3508,N_4844);
and U7045 (N_7045,N_5979,N_4824);
nor U7046 (N_7046,N_4079,N_4530);
or U7047 (N_7047,N_4288,N_5884);
nand U7048 (N_7048,N_4240,N_3236);
nand U7049 (N_7049,N_4011,N_5521);
or U7050 (N_7050,N_4117,N_4663);
xor U7051 (N_7051,N_4772,N_3899);
nor U7052 (N_7052,N_3513,N_5592);
nand U7053 (N_7053,N_3272,N_4791);
xnor U7054 (N_7054,N_5429,N_3444);
or U7055 (N_7055,N_5910,N_3958);
and U7056 (N_7056,N_4080,N_5696);
and U7057 (N_7057,N_5086,N_3939);
or U7058 (N_7058,N_5319,N_5851);
xor U7059 (N_7059,N_3998,N_4444);
xor U7060 (N_7060,N_5236,N_5832);
xnor U7061 (N_7061,N_4554,N_5258);
nand U7062 (N_7062,N_5941,N_4003);
and U7063 (N_7063,N_5013,N_4816);
xor U7064 (N_7064,N_5261,N_5711);
and U7065 (N_7065,N_3129,N_5265);
or U7066 (N_7066,N_5064,N_5450);
or U7067 (N_7067,N_5005,N_5486);
nor U7068 (N_7068,N_4030,N_4928);
xnor U7069 (N_7069,N_3594,N_5561);
or U7070 (N_7070,N_4402,N_5602);
nor U7071 (N_7071,N_5390,N_3204);
xor U7072 (N_7072,N_5145,N_3936);
xnor U7073 (N_7073,N_4664,N_3808);
nor U7074 (N_7074,N_5075,N_4508);
nand U7075 (N_7075,N_4375,N_3224);
nor U7076 (N_7076,N_5950,N_3557);
xnor U7077 (N_7077,N_3252,N_5784);
xor U7078 (N_7078,N_3076,N_5467);
nand U7079 (N_7079,N_4445,N_4827);
nor U7080 (N_7080,N_4614,N_4576);
and U7081 (N_7081,N_4050,N_5423);
nor U7082 (N_7082,N_4557,N_3160);
and U7083 (N_7083,N_3261,N_5174);
or U7084 (N_7084,N_3124,N_3674);
and U7085 (N_7085,N_4290,N_5704);
nor U7086 (N_7086,N_5682,N_3949);
xor U7087 (N_7087,N_4139,N_5116);
and U7088 (N_7088,N_5648,N_5271);
and U7089 (N_7089,N_3665,N_5218);
and U7090 (N_7090,N_4436,N_3968);
nand U7091 (N_7091,N_5433,N_5935);
and U7092 (N_7092,N_4084,N_4570);
xnor U7093 (N_7093,N_5788,N_3135);
xor U7094 (N_7094,N_3977,N_4913);
xor U7095 (N_7095,N_4267,N_5681);
and U7096 (N_7096,N_3147,N_3298);
and U7097 (N_7097,N_5224,N_5276);
nor U7098 (N_7098,N_3983,N_3953);
and U7099 (N_7099,N_3960,N_5526);
or U7100 (N_7100,N_4055,N_5658);
xor U7101 (N_7101,N_4915,N_5248);
nor U7102 (N_7102,N_5160,N_3615);
nor U7103 (N_7103,N_3449,N_3585);
or U7104 (N_7104,N_3906,N_4327);
nor U7105 (N_7105,N_4821,N_3388);
xnor U7106 (N_7106,N_4097,N_4942);
nor U7107 (N_7107,N_3580,N_3163);
or U7108 (N_7108,N_5310,N_5723);
or U7109 (N_7109,N_5339,N_4170);
or U7110 (N_7110,N_3707,N_3982);
and U7111 (N_7111,N_4854,N_3455);
nand U7112 (N_7112,N_5199,N_4189);
or U7113 (N_7113,N_5786,N_4987);
nand U7114 (N_7114,N_5577,N_3593);
nor U7115 (N_7115,N_5384,N_5356);
or U7116 (N_7116,N_5129,N_3242);
and U7117 (N_7117,N_4765,N_5945);
or U7118 (N_7118,N_5126,N_4128);
or U7119 (N_7119,N_5299,N_4361);
and U7120 (N_7120,N_4496,N_5444);
nor U7121 (N_7121,N_4606,N_4799);
or U7122 (N_7122,N_4573,N_3157);
or U7123 (N_7123,N_3263,N_5047);
xnor U7124 (N_7124,N_4427,N_5545);
xor U7125 (N_7125,N_3404,N_4617);
and U7126 (N_7126,N_3964,N_5506);
and U7127 (N_7127,N_5076,N_4597);
nand U7128 (N_7128,N_4997,N_4233);
nor U7129 (N_7129,N_5724,N_4888);
or U7130 (N_7130,N_5490,N_5612);
or U7131 (N_7131,N_4241,N_4138);
nand U7132 (N_7132,N_3483,N_3582);
and U7133 (N_7133,N_5868,N_4505);
nor U7134 (N_7134,N_3175,N_3310);
or U7135 (N_7135,N_4452,N_3049);
xor U7136 (N_7136,N_4487,N_4808);
and U7137 (N_7137,N_5626,N_4249);
or U7138 (N_7138,N_3137,N_5920);
nand U7139 (N_7139,N_3356,N_3146);
xor U7140 (N_7140,N_4601,N_4706);
or U7141 (N_7141,N_3838,N_4535);
and U7142 (N_7142,N_3216,N_5196);
and U7143 (N_7143,N_3372,N_3606);
nor U7144 (N_7144,N_4656,N_3026);
and U7145 (N_7145,N_3765,N_4596);
or U7146 (N_7146,N_5916,N_5395);
and U7147 (N_7147,N_4825,N_3235);
and U7148 (N_7148,N_3320,N_4812);
nor U7149 (N_7149,N_5401,N_3046);
or U7150 (N_7150,N_3560,N_3309);
nand U7151 (N_7151,N_4053,N_5232);
nand U7152 (N_7152,N_4313,N_3126);
nor U7153 (N_7153,N_5705,N_5548);
and U7154 (N_7154,N_5913,N_3284);
nand U7155 (N_7155,N_5981,N_4966);
or U7156 (N_7156,N_5926,N_5198);
or U7157 (N_7157,N_4075,N_5943);
and U7158 (N_7158,N_4624,N_5169);
nor U7159 (N_7159,N_5110,N_3468);
or U7160 (N_7160,N_4555,N_3534);
nand U7161 (N_7161,N_5774,N_4593);
nor U7162 (N_7162,N_5931,N_3259);
nor U7163 (N_7163,N_3564,N_3933);
or U7164 (N_7164,N_3996,N_4016);
and U7165 (N_7165,N_4865,N_3089);
xnor U7166 (N_7166,N_3015,N_5863);
nand U7167 (N_7167,N_4702,N_5172);
nand U7168 (N_7168,N_5992,N_4000);
nor U7169 (N_7169,N_4092,N_3108);
nand U7170 (N_7170,N_5697,N_4305);
xnor U7171 (N_7171,N_5328,N_4472);
nand U7172 (N_7172,N_4849,N_3700);
nand U7173 (N_7173,N_5907,N_5294);
and U7174 (N_7174,N_5213,N_4552);
xnor U7175 (N_7175,N_3938,N_3078);
and U7176 (N_7176,N_5079,N_4130);
and U7177 (N_7177,N_5348,N_4956);
nand U7178 (N_7178,N_5065,N_5819);
xor U7179 (N_7179,N_3321,N_4399);
xor U7180 (N_7180,N_4994,N_3156);
and U7181 (N_7181,N_5635,N_4757);
xnor U7182 (N_7182,N_3391,N_4602);
xor U7183 (N_7183,N_3392,N_3509);
nor U7184 (N_7184,N_5358,N_3478);
nand U7185 (N_7185,N_4969,N_3922);
or U7186 (N_7186,N_4925,N_5435);
nor U7187 (N_7187,N_5489,N_3034);
and U7188 (N_7188,N_3296,N_5291);
and U7189 (N_7189,N_4642,N_5975);
and U7190 (N_7190,N_5007,N_5002);
and U7191 (N_7191,N_5373,N_4566);
or U7192 (N_7192,N_4410,N_4099);
nand U7193 (N_7193,N_3094,N_4800);
or U7194 (N_7194,N_5375,N_5446);
xor U7195 (N_7195,N_4541,N_4809);
xor U7196 (N_7196,N_3043,N_5183);
xnor U7197 (N_7197,N_5933,N_5122);
nand U7198 (N_7198,N_5136,N_3793);
and U7199 (N_7199,N_4217,N_5852);
nor U7200 (N_7200,N_3102,N_5720);
or U7201 (N_7201,N_4661,N_3784);
or U7202 (N_7202,N_5750,N_5529);
nand U7203 (N_7203,N_5278,N_3955);
and U7204 (N_7204,N_3439,N_3702);
xnor U7205 (N_7205,N_5016,N_4352);
nor U7206 (N_7206,N_5364,N_4546);
or U7207 (N_7207,N_4221,N_4748);
xor U7208 (N_7208,N_3300,N_4271);
and U7209 (N_7209,N_4882,N_3346);
nor U7210 (N_7210,N_4525,N_4094);
xor U7211 (N_7211,N_4293,N_4778);
and U7212 (N_7212,N_4659,N_5957);
xor U7213 (N_7213,N_4504,N_4564);
xnor U7214 (N_7214,N_4725,N_3307);
and U7215 (N_7215,N_5640,N_3230);
nand U7216 (N_7216,N_3365,N_3815);
xor U7217 (N_7217,N_3413,N_4264);
nor U7218 (N_7218,N_4907,N_5253);
or U7219 (N_7219,N_4414,N_3169);
nand U7220 (N_7220,N_4575,N_4473);
nand U7221 (N_7221,N_4937,N_5675);
nor U7222 (N_7222,N_4953,N_5520);
nand U7223 (N_7223,N_3644,N_4362);
nor U7224 (N_7224,N_4125,N_4968);
or U7225 (N_7225,N_3246,N_4491);
nor U7226 (N_7226,N_3663,N_4780);
nand U7227 (N_7227,N_5735,N_5237);
nand U7228 (N_7228,N_3070,N_5901);
nor U7229 (N_7229,N_4839,N_4244);
nand U7230 (N_7230,N_4100,N_4709);
and U7231 (N_7231,N_5286,N_5335);
and U7232 (N_7232,N_4040,N_4031);
nor U7233 (N_7233,N_3908,N_3423);
or U7234 (N_7234,N_5137,N_5333);
nor U7235 (N_7235,N_3362,N_4716);
nand U7236 (N_7236,N_5912,N_5780);
nand U7237 (N_7237,N_5882,N_3003);
nand U7238 (N_7238,N_3282,N_4154);
nor U7239 (N_7239,N_4025,N_4002);
xor U7240 (N_7240,N_5685,N_3430);
and U7241 (N_7241,N_5266,N_4136);
nand U7242 (N_7242,N_4901,N_4502);
nand U7243 (N_7243,N_4259,N_5151);
and U7244 (N_7244,N_4215,N_5880);
and U7245 (N_7245,N_5025,N_3640);
nor U7246 (N_7246,N_4194,N_4147);
or U7247 (N_7247,N_3848,N_3341);
nor U7248 (N_7248,N_5043,N_5084);
and U7249 (N_7249,N_3469,N_4022);
and U7250 (N_7250,N_5773,N_3381);
nand U7251 (N_7251,N_3194,N_5582);
nand U7252 (N_7252,N_4848,N_5019);
or U7253 (N_7253,N_5549,N_4475);
nand U7254 (N_7254,N_5083,N_3396);
xnor U7255 (N_7255,N_3228,N_4344);
xor U7256 (N_7256,N_5131,N_4524);
and U7257 (N_7257,N_5956,N_4950);
and U7258 (N_7258,N_3205,N_4253);
xor U7259 (N_7259,N_4235,N_4302);
nor U7260 (N_7260,N_5777,N_4670);
nor U7261 (N_7261,N_3519,N_4861);
xor U7262 (N_7262,N_5127,N_5470);
nor U7263 (N_7263,N_4076,N_4358);
and U7264 (N_7264,N_3789,N_4588);
nor U7265 (N_7265,N_5445,N_5759);
nor U7266 (N_7266,N_4544,N_5515);
nor U7267 (N_7267,N_3873,N_5715);
nor U7268 (N_7268,N_3503,N_5071);
and U7269 (N_7269,N_5701,N_3314);
nand U7270 (N_7270,N_4008,N_3022);
and U7271 (N_7271,N_4872,N_5391);
nor U7272 (N_7272,N_4466,N_3973);
xor U7273 (N_7273,N_4462,N_3407);
nand U7274 (N_7274,N_5357,N_5993);
nor U7275 (N_7275,N_4644,N_5402);
xnor U7276 (N_7276,N_3569,N_5670);
xnor U7277 (N_7277,N_3753,N_3178);
or U7278 (N_7278,N_5491,N_4675);
xnor U7279 (N_7279,N_3529,N_5946);
nor U7280 (N_7280,N_4334,N_5580);
and U7281 (N_7281,N_5133,N_3200);
nand U7282 (N_7282,N_3476,N_4236);
nand U7283 (N_7283,N_5647,N_5473);
or U7284 (N_7284,N_3410,N_3581);
or U7285 (N_7285,N_3617,N_3501);
nand U7286 (N_7286,N_4755,N_4932);
and U7287 (N_7287,N_4633,N_4949);
and U7288 (N_7288,N_4995,N_5686);
or U7289 (N_7289,N_3643,N_5762);
nor U7290 (N_7290,N_4837,N_3860);
and U7291 (N_7291,N_4144,N_3191);
xnor U7292 (N_7292,N_5341,N_4107);
and U7293 (N_7293,N_3255,N_3835);
nand U7294 (N_7294,N_3768,N_3763);
and U7295 (N_7295,N_3834,N_4135);
and U7296 (N_7296,N_5656,N_4324);
and U7297 (N_7297,N_4419,N_3142);
or U7298 (N_7298,N_4082,N_5827);
nand U7299 (N_7299,N_5984,N_5051);
and U7300 (N_7300,N_4322,N_5142);
xor U7301 (N_7301,N_5164,N_5639);
and U7302 (N_7302,N_4703,N_3687);
or U7303 (N_7303,N_5492,N_5495);
nand U7304 (N_7304,N_3106,N_3382);
and U7305 (N_7305,N_5327,N_5001);
and U7306 (N_7306,N_4751,N_3575);
nand U7307 (N_7307,N_5726,N_5303);
xnor U7308 (N_7308,N_3233,N_4796);
xor U7309 (N_7309,N_5215,N_5798);
nand U7310 (N_7310,N_4485,N_4636);
xnor U7311 (N_7311,N_3897,N_3264);
and U7312 (N_7312,N_3827,N_4380);
xnor U7313 (N_7313,N_3337,N_5379);
nor U7314 (N_7314,N_3398,N_3463);
nand U7315 (N_7315,N_3384,N_3018);
nor U7316 (N_7316,N_4902,N_4458);
and U7317 (N_7317,N_4382,N_4116);
or U7318 (N_7318,N_3143,N_4641);
and U7319 (N_7319,N_5608,N_5550);
and U7320 (N_7320,N_3999,N_4388);
nor U7321 (N_7321,N_4179,N_4833);
or U7322 (N_7322,N_5839,N_3573);
xor U7323 (N_7323,N_5509,N_3237);
nand U7324 (N_7324,N_5834,N_5680);
nand U7325 (N_7325,N_4581,N_4017);
or U7326 (N_7326,N_4910,N_4133);
nand U7327 (N_7327,N_3318,N_5917);
or U7328 (N_7328,N_4742,N_3327);
nand U7329 (N_7329,N_5963,N_3514);
xor U7330 (N_7330,N_5088,N_5587);
nand U7331 (N_7331,N_3891,N_4753);
nor U7332 (N_7332,N_5801,N_4266);
nand U7333 (N_7333,N_5803,N_5995);
nor U7334 (N_7334,N_4006,N_5469);
nand U7335 (N_7335,N_3952,N_5135);
or U7336 (N_7336,N_4173,N_4357);
and U7337 (N_7337,N_4276,N_3988);
xnor U7338 (N_7338,N_5093,N_3122);
or U7339 (N_7339,N_3425,N_3288);
or U7340 (N_7340,N_3945,N_3862);
nor U7341 (N_7341,N_5471,N_4499);
or U7342 (N_7342,N_5257,N_3641);
nor U7343 (N_7343,N_4209,N_3280);
xor U7344 (N_7344,N_3701,N_3051);
xor U7345 (N_7345,N_5378,N_3221);
nand U7346 (N_7346,N_3741,N_5985);
nand U7347 (N_7347,N_3283,N_4250);
nand U7348 (N_7348,N_4381,N_3792);
xor U7349 (N_7349,N_3507,N_3567);
xor U7350 (N_7350,N_4064,N_3579);
or U7351 (N_7351,N_5320,N_5540);
nor U7352 (N_7352,N_3568,N_5481);
and U7353 (N_7353,N_3680,N_3927);
xnor U7354 (N_7354,N_4628,N_4537);
nor U7355 (N_7355,N_3609,N_3040);
nor U7356 (N_7356,N_5836,N_3192);
xor U7357 (N_7357,N_5915,N_3092);
nand U7358 (N_7358,N_5959,N_5302);
or U7359 (N_7359,N_4585,N_4639);
and U7360 (N_7360,N_4211,N_3645);
xnor U7361 (N_7361,N_5474,N_3152);
or U7362 (N_7362,N_5239,N_3956);
and U7363 (N_7363,N_5478,N_4420);
nor U7364 (N_7364,N_5228,N_4063);
nand U7365 (N_7365,N_3818,N_5082);
or U7366 (N_7366,N_5251,N_3432);
nand U7367 (N_7367,N_3304,N_4142);
and U7368 (N_7368,N_3344,N_4166);
nand U7369 (N_7369,N_3466,N_4319);
xor U7370 (N_7370,N_5180,N_4934);
xnor U7371 (N_7371,N_4724,N_3039);
or U7372 (N_7372,N_4477,N_3023);
nand U7373 (N_7373,N_5934,N_4977);
xnor U7374 (N_7374,N_3769,N_3174);
nor U7375 (N_7375,N_3893,N_5501);
and U7376 (N_7376,N_3577,N_5903);
nand U7377 (N_7377,N_3586,N_3482);
nand U7378 (N_7378,N_4567,N_5417);
and U7379 (N_7379,N_4649,N_5034);
xnor U7380 (N_7380,N_3535,N_3602);
and U7381 (N_7381,N_5861,N_3916);
xor U7382 (N_7382,N_5814,N_3859);
nand U7383 (N_7383,N_3438,N_5179);
nor U7384 (N_7384,N_5447,N_4123);
xnor U7385 (N_7385,N_4056,N_4118);
nor U7386 (N_7386,N_3319,N_4245);
xnor U7387 (N_7387,N_3374,N_5672);
or U7388 (N_7388,N_4051,N_4536);
nor U7389 (N_7389,N_3551,N_5297);
nor U7390 (N_7390,N_3849,N_5969);
nor U7391 (N_7391,N_4309,N_4158);
or U7392 (N_7392,N_4248,N_4657);
and U7393 (N_7393,N_3809,N_5905);
or U7394 (N_7394,N_5295,N_5021);
nand U7395 (N_7395,N_3920,N_5513);
xnor U7396 (N_7396,N_4767,N_4813);
and U7397 (N_7397,N_5270,N_5633);
xor U7398 (N_7398,N_5779,N_4858);
nand U7399 (N_7399,N_3744,N_5205);
or U7400 (N_7400,N_3487,N_5003);
or U7401 (N_7401,N_4986,N_4047);
nor U7402 (N_7402,N_3636,N_4354);
nand U7403 (N_7403,N_5150,N_5522);
xor U7404 (N_7404,N_4558,N_3616);
or U7405 (N_7405,N_5371,N_4216);
nand U7406 (N_7406,N_3981,N_5182);
or U7407 (N_7407,N_5259,N_3399);
and U7408 (N_7408,N_4350,N_4467);
nand U7409 (N_7409,N_3340,N_5604);
or U7410 (N_7410,N_5197,N_4405);
and U7411 (N_7411,N_5609,N_3334);
and U7412 (N_7412,N_4962,N_5503);
xnor U7413 (N_7413,N_5109,N_4918);
or U7414 (N_7414,N_3170,N_5983);
nand U7415 (N_7415,N_5749,N_4023);
xor U7416 (N_7416,N_5536,N_5392);
nand U7417 (N_7417,N_4760,N_3677);
xor U7418 (N_7418,N_5369,N_3940);
xor U7419 (N_7419,N_3377,N_3045);
nand U7420 (N_7420,N_5751,N_3682);
or U7421 (N_7421,N_3724,N_4413);
xnor U7422 (N_7422,N_4145,N_5027);
or U7423 (N_7423,N_4754,N_3735);
and U7424 (N_7424,N_5678,N_4488);
xnor U7425 (N_7425,N_5761,N_5677);
xor U7426 (N_7426,N_4652,N_3544);
nor U7427 (N_7427,N_5089,N_3073);
xnor U7428 (N_7428,N_5010,N_5033);
or U7429 (N_7429,N_3467,N_5285);
or U7430 (N_7430,N_5572,N_5971);
xor U7431 (N_7431,N_5038,N_3562);
nor U7432 (N_7432,N_3652,N_4841);
nand U7433 (N_7433,N_5193,N_4875);
or U7434 (N_7434,N_4904,N_4665);
nor U7435 (N_7435,N_3295,N_3287);
nor U7436 (N_7436,N_3218,N_4004);
or U7437 (N_7437,N_5942,N_5732);
or U7438 (N_7438,N_3833,N_4098);
and U7439 (N_7439,N_3329,N_4752);
or U7440 (N_7440,N_5440,N_5244);
nor U7441 (N_7441,N_4836,N_5886);
and U7442 (N_7442,N_5425,N_5171);
and U7443 (N_7443,N_4776,N_3635);
or U7444 (N_7444,N_4480,N_4774);
xnor U7445 (N_7445,N_3855,N_4059);
nand U7446 (N_7446,N_5212,N_5114);
and U7447 (N_7447,N_5731,N_3290);
xor U7448 (N_7448,N_3215,N_3352);
and U7449 (N_7449,N_5499,N_3193);
xnor U7450 (N_7450,N_4364,N_4571);
nand U7451 (N_7451,N_5074,N_5728);
and U7452 (N_7452,N_3498,N_4337);
or U7453 (N_7453,N_5479,N_4733);
and U7454 (N_7454,N_5042,N_4936);
and U7455 (N_7455,N_5833,N_3197);
nand U7456 (N_7456,N_5324,N_5891);
and U7457 (N_7457,N_3195,N_3948);
and U7458 (N_7458,N_3354,N_5783);
and U7459 (N_7459,N_3210,N_5048);
nand U7460 (N_7460,N_5163,N_3876);
nor U7461 (N_7461,N_4835,N_5396);
or U7462 (N_7462,N_5755,N_4081);
or U7463 (N_7463,N_3072,N_4783);
nor U7464 (N_7464,N_5090,N_5669);
nand U7465 (N_7465,N_5466,N_4683);
and U7466 (N_7466,N_4654,N_3758);
nand U7467 (N_7467,N_4262,N_5404);
nand U7468 (N_7468,N_5610,N_5426);
nor U7469 (N_7469,N_3728,N_4736);
or U7470 (N_7470,N_3457,N_5617);
xnor U7471 (N_7471,N_4927,N_5892);
nand U7472 (N_7472,N_3222,N_4893);
nor U7473 (N_7473,N_3207,N_5624);
or U7474 (N_7474,N_5030,N_3436);
or U7475 (N_7475,N_3989,N_3703);
nor U7476 (N_7476,N_3696,N_4775);
and U7477 (N_7477,N_3539,N_5676);
or U7478 (N_7478,N_4481,N_5454);
nand U7479 (N_7479,N_4095,N_4826);
or U7480 (N_7480,N_3942,N_5908);
xor U7481 (N_7481,N_4332,N_4300);
nand U7482 (N_7482,N_3486,N_5121);
and U7483 (N_7483,N_4214,N_4713);
or U7484 (N_7484,N_3886,N_3440);
or U7485 (N_7485,N_5727,N_3850);
and U7486 (N_7486,N_4085,N_3705);
or U7487 (N_7487,N_3921,N_4720);
nand U7488 (N_7488,N_4314,N_3456);
xnor U7489 (N_7489,N_5249,N_4330);
nand U7490 (N_7490,N_3203,N_4509);
xnor U7491 (N_7491,N_3553,N_5242);
xor U7492 (N_7492,N_4024,N_5590);
and U7493 (N_7493,N_4806,N_5041);
and U7494 (N_7494,N_3563,N_3016);
or U7495 (N_7495,N_3011,N_3984);
or U7496 (N_7496,N_4279,N_4694);
or U7497 (N_7497,N_4408,N_4256);
and U7498 (N_7498,N_4595,N_3209);
xnor U7499 (N_7499,N_3887,N_3154);
and U7500 (N_7500,N_4325,N_5151);
and U7501 (N_7501,N_5671,N_4925);
nand U7502 (N_7502,N_4583,N_3644);
nand U7503 (N_7503,N_3972,N_4121);
nand U7504 (N_7504,N_5326,N_3770);
and U7505 (N_7505,N_3011,N_3280);
xnor U7506 (N_7506,N_5648,N_3663);
and U7507 (N_7507,N_5494,N_4453);
or U7508 (N_7508,N_5203,N_5960);
nor U7509 (N_7509,N_3840,N_3882);
xor U7510 (N_7510,N_3464,N_5077);
nor U7511 (N_7511,N_4947,N_5603);
and U7512 (N_7512,N_5874,N_4403);
nand U7513 (N_7513,N_3635,N_4997);
or U7514 (N_7514,N_4170,N_3116);
and U7515 (N_7515,N_5728,N_3544);
nor U7516 (N_7516,N_5403,N_5737);
nor U7517 (N_7517,N_4822,N_3625);
and U7518 (N_7518,N_4150,N_5941);
and U7519 (N_7519,N_3375,N_3666);
or U7520 (N_7520,N_3988,N_4592);
and U7521 (N_7521,N_4732,N_3012);
nor U7522 (N_7522,N_3156,N_3319);
or U7523 (N_7523,N_4726,N_5161);
nand U7524 (N_7524,N_3910,N_5581);
nor U7525 (N_7525,N_3755,N_3415);
xor U7526 (N_7526,N_3666,N_5129);
nand U7527 (N_7527,N_4342,N_5663);
and U7528 (N_7528,N_4324,N_5707);
and U7529 (N_7529,N_3527,N_3084);
or U7530 (N_7530,N_4483,N_5854);
xnor U7531 (N_7531,N_5320,N_5558);
nor U7532 (N_7532,N_5123,N_4597);
nor U7533 (N_7533,N_5497,N_4458);
and U7534 (N_7534,N_3533,N_4480);
nor U7535 (N_7535,N_5468,N_4729);
nand U7536 (N_7536,N_4258,N_5233);
nand U7537 (N_7537,N_5948,N_4422);
xnor U7538 (N_7538,N_4181,N_4172);
and U7539 (N_7539,N_5561,N_4285);
and U7540 (N_7540,N_4921,N_3537);
nand U7541 (N_7541,N_4429,N_5097);
nor U7542 (N_7542,N_4564,N_4802);
nand U7543 (N_7543,N_3413,N_5657);
or U7544 (N_7544,N_4728,N_4254);
xnor U7545 (N_7545,N_4339,N_4903);
nand U7546 (N_7546,N_4975,N_5446);
or U7547 (N_7547,N_3355,N_3257);
nor U7548 (N_7548,N_5833,N_4848);
nor U7549 (N_7549,N_3256,N_4133);
or U7550 (N_7550,N_5730,N_5644);
and U7551 (N_7551,N_3866,N_3356);
xor U7552 (N_7552,N_5391,N_5191);
xnor U7553 (N_7553,N_3938,N_5774);
and U7554 (N_7554,N_3614,N_5896);
and U7555 (N_7555,N_5459,N_5972);
xnor U7556 (N_7556,N_5435,N_3552);
nor U7557 (N_7557,N_4785,N_4563);
nor U7558 (N_7558,N_4709,N_3135);
nor U7559 (N_7559,N_3038,N_4780);
and U7560 (N_7560,N_5511,N_4473);
xnor U7561 (N_7561,N_5981,N_5803);
and U7562 (N_7562,N_4143,N_4189);
nand U7563 (N_7563,N_4724,N_3294);
xor U7564 (N_7564,N_4742,N_4248);
or U7565 (N_7565,N_4588,N_3847);
and U7566 (N_7566,N_5487,N_5315);
and U7567 (N_7567,N_3289,N_3991);
nor U7568 (N_7568,N_3841,N_5595);
nor U7569 (N_7569,N_4757,N_4467);
and U7570 (N_7570,N_5308,N_5802);
nor U7571 (N_7571,N_3043,N_4897);
or U7572 (N_7572,N_3520,N_5671);
nor U7573 (N_7573,N_3499,N_4737);
xnor U7574 (N_7574,N_5125,N_4946);
nand U7575 (N_7575,N_5802,N_4284);
or U7576 (N_7576,N_5635,N_3828);
and U7577 (N_7577,N_3370,N_3041);
nor U7578 (N_7578,N_4492,N_3914);
xnor U7579 (N_7579,N_3181,N_5039);
nor U7580 (N_7580,N_4651,N_3477);
and U7581 (N_7581,N_4646,N_3052);
nor U7582 (N_7582,N_5473,N_3346);
and U7583 (N_7583,N_4596,N_3691);
or U7584 (N_7584,N_5453,N_4983);
and U7585 (N_7585,N_5909,N_4521);
xnor U7586 (N_7586,N_3173,N_5336);
or U7587 (N_7587,N_4034,N_4736);
nor U7588 (N_7588,N_5798,N_5718);
or U7589 (N_7589,N_4602,N_3402);
xnor U7590 (N_7590,N_3630,N_5606);
nor U7591 (N_7591,N_4866,N_3791);
nand U7592 (N_7592,N_5122,N_3446);
nand U7593 (N_7593,N_3602,N_4037);
nor U7594 (N_7594,N_3282,N_4354);
nand U7595 (N_7595,N_5664,N_3486);
or U7596 (N_7596,N_4447,N_4328);
and U7597 (N_7597,N_5023,N_4179);
or U7598 (N_7598,N_5638,N_4782);
xor U7599 (N_7599,N_5187,N_4906);
nor U7600 (N_7600,N_4413,N_3791);
xor U7601 (N_7601,N_3114,N_3370);
nand U7602 (N_7602,N_3117,N_5409);
nor U7603 (N_7603,N_3591,N_4802);
and U7604 (N_7604,N_3285,N_3182);
nand U7605 (N_7605,N_3333,N_5939);
xnor U7606 (N_7606,N_4901,N_3207);
and U7607 (N_7607,N_5402,N_5134);
and U7608 (N_7608,N_4335,N_3418);
xor U7609 (N_7609,N_3753,N_4060);
nand U7610 (N_7610,N_5390,N_4486);
nor U7611 (N_7611,N_5682,N_4614);
and U7612 (N_7612,N_3654,N_4449);
or U7613 (N_7613,N_3617,N_5965);
or U7614 (N_7614,N_4595,N_4111);
nor U7615 (N_7615,N_4071,N_4417);
nor U7616 (N_7616,N_3960,N_5116);
nor U7617 (N_7617,N_5606,N_5821);
or U7618 (N_7618,N_5222,N_5156);
nand U7619 (N_7619,N_5460,N_4361);
and U7620 (N_7620,N_3060,N_5421);
or U7621 (N_7621,N_5998,N_4063);
and U7622 (N_7622,N_3568,N_4628);
or U7623 (N_7623,N_3019,N_5365);
xor U7624 (N_7624,N_3075,N_5929);
nor U7625 (N_7625,N_3530,N_4435);
nor U7626 (N_7626,N_3329,N_5407);
nand U7627 (N_7627,N_3527,N_4141);
xnor U7628 (N_7628,N_5811,N_3490);
or U7629 (N_7629,N_3195,N_4497);
nand U7630 (N_7630,N_5675,N_3409);
nor U7631 (N_7631,N_5435,N_5293);
xnor U7632 (N_7632,N_4123,N_4380);
nand U7633 (N_7633,N_5951,N_4773);
xnor U7634 (N_7634,N_3949,N_5567);
and U7635 (N_7635,N_5971,N_4872);
and U7636 (N_7636,N_5447,N_5180);
nand U7637 (N_7637,N_3109,N_5526);
nor U7638 (N_7638,N_5100,N_3298);
nor U7639 (N_7639,N_4582,N_5056);
nand U7640 (N_7640,N_3446,N_4536);
nand U7641 (N_7641,N_4820,N_4797);
or U7642 (N_7642,N_3966,N_5597);
or U7643 (N_7643,N_4634,N_3533);
or U7644 (N_7644,N_4296,N_3850);
or U7645 (N_7645,N_4305,N_4824);
or U7646 (N_7646,N_5174,N_3301);
and U7647 (N_7647,N_5763,N_5540);
nor U7648 (N_7648,N_3403,N_4026);
and U7649 (N_7649,N_4817,N_3355);
xnor U7650 (N_7650,N_5317,N_3035);
xor U7651 (N_7651,N_4762,N_5719);
nand U7652 (N_7652,N_5423,N_5611);
or U7653 (N_7653,N_4613,N_4189);
nor U7654 (N_7654,N_5900,N_5246);
or U7655 (N_7655,N_3319,N_4561);
nor U7656 (N_7656,N_5099,N_4471);
nor U7657 (N_7657,N_4461,N_5359);
xor U7658 (N_7658,N_4845,N_4334);
or U7659 (N_7659,N_3957,N_5832);
nand U7660 (N_7660,N_5273,N_4204);
nor U7661 (N_7661,N_5189,N_4678);
or U7662 (N_7662,N_4186,N_4349);
nand U7663 (N_7663,N_4652,N_3995);
nand U7664 (N_7664,N_5129,N_4400);
or U7665 (N_7665,N_4484,N_3100);
nand U7666 (N_7666,N_3225,N_5793);
or U7667 (N_7667,N_3424,N_3464);
or U7668 (N_7668,N_3750,N_4174);
nand U7669 (N_7669,N_4218,N_4450);
or U7670 (N_7670,N_4676,N_5956);
or U7671 (N_7671,N_3204,N_4413);
or U7672 (N_7672,N_3478,N_5994);
or U7673 (N_7673,N_3745,N_5456);
nand U7674 (N_7674,N_3392,N_4944);
and U7675 (N_7675,N_3410,N_5092);
or U7676 (N_7676,N_4330,N_3969);
nor U7677 (N_7677,N_3157,N_3074);
xnor U7678 (N_7678,N_4030,N_5148);
nand U7679 (N_7679,N_4997,N_4268);
nor U7680 (N_7680,N_3364,N_3675);
or U7681 (N_7681,N_5971,N_5816);
or U7682 (N_7682,N_4683,N_5796);
and U7683 (N_7683,N_3398,N_3479);
nand U7684 (N_7684,N_4051,N_5957);
nor U7685 (N_7685,N_5059,N_4667);
and U7686 (N_7686,N_3797,N_3090);
nand U7687 (N_7687,N_5390,N_5973);
or U7688 (N_7688,N_5066,N_3226);
nand U7689 (N_7689,N_4937,N_4668);
xnor U7690 (N_7690,N_5850,N_4644);
xor U7691 (N_7691,N_4763,N_5841);
nor U7692 (N_7692,N_4217,N_5424);
and U7693 (N_7693,N_4570,N_3488);
nor U7694 (N_7694,N_4232,N_3946);
nand U7695 (N_7695,N_4711,N_5954);
nor U7696 (N_7696,N_4658,N_3993);
or U7697 (N_7697,N_4875,N_3294);
and U7698 (N_7698,N_3379,N_4688);
xnor U7699 (N_7699,N_4482,N_3998);
and U7700 (N_7700,N_3332,N_4573);
nor U7701 (N_7701,N_4877,N_3415);
or U7702 (N_7702,N_3772,N_5063);
xnor U7703 (N_7703,N_3568,N_4064);
nor U7704 (N_7704,N_4262,N_3175);
or U7705 (N_7705,N_3417,N_4124);
nand U7706 (N_7706,N_4990,N_3033);
and U7707 (N_7707,N_5568,N_5209);
and U7708 (N_7708,N_4139,N_3268);
and U7709 (N_7709,N_3791,N_5564);
and U7710 (N_7710,N_5845,N_4440);
or U7711 (N_7711,N_5964,N_3912);
and U7712 (N_7712,N_4886,N_5235);
xnor U7713 (N_7713,N_5152,N_4630);
xnor U7714 (N_7714,N_3373,N_4308);
nor U7715 (N_7715,N_3597,N_3336);
and U7716 (N_7716,N_3708,N_5747);
nand U7717 (N_7717,N_4135,N_4882);
or U7718 (N_7718,N_3954,N_5137);
or U7719 (N_7719,N_5314,N_5756);
xnor U7720 (N_7720,N_5231,N_3327);
and U7721 (N_7721,N_5149,N_5344);
and U7722 (N_7722,N_5719,N_4526);
nor U7723 (N_7723,N_5763,N_5006);
nor U7724 (N_7724,N_3005,N_5943);
xnor U7725 (N_7725,N_3251,N_4919);
nand U7726 (N_7726,N_3133,N_5470);
nor U7727 (N_7727,N_5674,N_3439);
xor U7728 (N_7728,N_3738,N_5837);
nor U7729 (N_7729,N_3801,N_3733);
or U7730 (N_7730,N_5895,N_3782);
or U7731 (N_7731,N_5868,N_4742);
and U7732 (N_7732,N_5472,N_4407);
nand U7733 (N_7733,N_3278,N_5393);
xor U7734 (N_7734,N_4817,N_3995);
or U7735 (N_7735,N_4736,N_3196);
and U7736 (N_7736,N_4063,N_5072);
and U7737 (N_7737,N_5913,N_4636);
or U7738 (N_7738,N_5196,N_3822);
nor U7739 (N_7739,N_4798,N_5102);
nand U7740 (N_7740,N_3005,N_4631);
nand U7741 (N_7741,N_3051,N_4861);
xnor U7742 (N_7742,N_5658,N_5343);
nand U7743 (N_7743,N_4921,N_3027);
or U7744 (N_7744,N_4819,N_5539);
and U7745 (N_7745,N_5745,N_5990);
and U7746 (N_7746,N_3092,N_4735);
nor U7747 (N_7747,N_4788,N_4521);
and U7748 (N_7748,N_5985,N_3641);
nand U7749 (N_7749,N_3347,N_5656);
xnor U7750 (N_7750,N_5361,N_4162);
or U7751 (N_7751,N_3310,N_5896);
nor U7752 (N_7752,N_4734,N_3007);
nand U7753 (N_7753,N_5289,N_5104);
or U7754 (N_7754,N_5610,N_3209);
xor U7755 (N_7755,N_3394,N_3842);
and U7756 (N_7756,N_3116,N_4206);
or U7757 (N_7757,N_4000,N_4395);
nor U7758 (N_7758,N_3861,N_4791);
and U7759 (N_7759,N_5590,N_5214);
or U7760 (N_7760,N_5880,N_5733);
nor U7761 (N_7761,N_3276,N_5723);
xnor U7762 (N_7762,N_3530,N_3964);
and U7763 (N_7763,N_5939,N_3318);
nand U7764 (N_7764,N_5244,N_4449);
or U7765 (N_7765,N_3836,N_4523);
and U7766 (N_7766,N_3581,N_3572);
nand U7767 (N_7767,N_5608,N_5801);
or U7768 (N_7768,N_4741,N_5657);
xnor U7769 (N_7769,N_5132,N_5805);
and U7770 (N_7770,N_4904,N_5355);
nand U7771 (N_7771,N_3159,N_4722);
or U7772 (N_7772,N_5780,N_3738);
or U7773 (N_7773,N_5098,N_5830);
or U7774 (N_7774,N_4746,N_4319);
or U7775 (N_7775,N_4106,N_5831);
and U7776 (N_7776,N_3135,N_3158);
nand U7777 (N_7777,N_5834,N_4286);
xor U7778 (N_7778,N_3097,N_4145);
nor U7779 (N_7779,N_5448,N_5541);
xnor U7780 (N_7780,N_4646,N_3677);
or U7781 (N_7781,N_4974,N_4021);
or U7782 (N_7782,N_3591,N_3365);
nand U7783 (N_7783,N_5597,N_3655);
nor U7784 (N_7784,N_5859,N_4978);
xnor U7785 (N_7785,N_4287,N_4100);
xor U7786 (N_7786,N_3250,N_3098);
or U7787 (N_7787,N_4918,N_3313);
nand U7788 (N_7788,N_3598,N_4075);
xor U7789 (N_7789,N_4645,N_5809);
nor U7790 (N_7790,N_5119,N_4644);
nand U7791 (N_7791,N_5620,N_4316);
or U7792 (N_7792,N_4574,N_4885);
or U7793 (N_7793,N_5557,N_5842);
and U7794 (N_7794,N_5036,N_3764);
and U7795 (N_7795,N_3464,N_5213);
nor U7796 (N_7796,N_4962,N_5042);
or U7797 (N_7797,N_5141,N_4742);
nand U7798 (N_7798,N_3316,N_3880);
nand U7799 (N_7799,N_3024,N_4676);
or U7800 (N_7800,N_5505,N_3596);
nand U7801 (N_7801,N_5160,N_3209);
and U7802 (N_7802,N_4322,N_4371);
xnor U7803 (N_7803,N_3655,N_4619);
and U7804 (N_7804,N_4401,N_5462);
nor U7805 (N_7805,N_5058,N_5707);
xnor U7806 (N_7806,N_3455,N_4394);
xnor U7807 (N_7807,N_5693,N_3146);
or U7808 (N_7808,N_4809,N_4370);
nand U7809 (N_7809,N_4876,N_4700);
xnor U7810 (N_7810,N_3805,N_5380);
nand U7811 (N_7811,N_3520,N_3872);
and U7812 (N_7812,N_5696,N_3276);
nand U7813 (N_7813,N_4432,N_3734);
xor U7814 (N_7814,N_3198,N_3626);
and U7815 (N_7815,N_4695,N_3532);
nor U7816 (N_7816,N_3283,N_4084);
nand U7817 (N_7817,N_4381,N_3882);
xnor U7818 (N_7818,N_5578,N_3816);
and U7819 (N_7819,N_3017,N_3696);
xnor U7820 (N_7820,N_4871,N_4966);
nor U7821 (N_7821,N_3345,N_5555);
xor U7822 (N_7822,N_4848,N_3663);
xor U7823 (N_7823,N_4702,N_4106);
and U7824 (N_7824,N_5000,N_5572);
nor U7825 (N_7825,N_3547,N_4308);
or U7826 (N_7826,N_5937,N_5460);
and U7827 (N_7827,N_5654,N_4545);
nor U7828 (N_7828,N_3561,N_5002);
and U7829 (N_7829,N_3897,N_5019);
xnor U7830 (N_7830,N_5091,N_4643);
xor U7831 (N_7831,N_5345,N_5232);
nand U7832 (N_7832,N_3909,N_4296);
xor U7833 (N_7833,N_4991,N_4997);
and U7834 (N_7834,N_4958,N_4687);
xor U7835 (N_7835,N_3657,N_5242);
and U7836 (N_7836,N_3309,N_4717);
or U7837 (N_7837,N_5356,N_5812);
and U7838 (N_7838,N_5539,N_3967);
xor U7839 (N_7839,N_5956,N_5446);
xor U7840 (N_7840,N_5919,N_4125);
xnor U7841 (N_7841,N_5943,N_3253);
nor U7842 (N_7842,N_3705,N_3684);
nor U7843 (N_7843,N_3942,N_5619);
xnor U7844 (N_7844,N_3979,N_4850);
and U7845 (N_7845,N_3143,N_5331);
nand U7846 (N_7846,N_5660,N_3655);
xor U7847 (N_7847,N_3507,N_5730);
xor U7848 (N_7848,N_4488,N_5176);
nor U7849 (N_7849,N_5166,N_4161);
xor U7850 (N_7850,N_5756,N_5038);
xnor U7851 (N_7851,N_5316,N_4914);
xor U7852 (N_7852,N_3236,N_3719);
or U7853 (N_7853,N_5835,N_3843);
and U7854 (N_7854,N_4532,N_4744);
nand U7855 (N_7855,N_5846,N_3295);
xor U7856 (N_7856,N_5638,N_3219);
or U7857 (N_7857,N_3372,N_3745);
nand U7858 (N_7858,N_5895,N_5930);
nor U7859 (N_7859,N_5805,N_5787);
nand U7860 (N_7860,N_3808,N_5264);
xnor U7861 (N_7861,N_3495,N_5669);
or U7862 (N_7862,N_4450,N_4211);
nor U7863 (N_7863,N_5234,N_3250);
and U7864 (N_7864,N_4079,N_3623);
nor U7865 (N_7865,N_4388,N_5870);
nand U7866 (N_7866,N_4515,N_5979);
or U7867 (N_7867,N_5859,N_3894);
xnor U7868 (N_7868,N_4152,N_3199);
or U7869 (N_7869,N_3322,N_4244);
nand U7870 (N_7870,N_5920,N_3775);
nor U7871 (N_7871,N_5547,N_5041);
nand U7872 (N_7872,N_3579,N_4937);
xnor U7873 (N_7873,N_4572,N_5286);
nand U7874 (N_7874,N_4361,N_3298);
nand U7875 (N_7875,N_4008,N_3159);
xnor U7876 (N_7876,N_3999,N_3955);
or U7877 (N_7877,N_4783,N_5461);
nor U7878 (N_7878,N_5892,N_3425);
and U7879 (N_7879,N_4100,N_4542);
xnor U7880 (N_7880,N_4718,N_4844);
xor U7881 (N_7881,N_5139,N_4463);
or U7882 (N_7882,N_5620,N_3888);
and U7883 (N_7883,N_4269,N_5672);
nor U7884 (N_7884,N_3017,N_5869);
or U7885 (N_7885,N_4430,N_5661);
nor U7886 (N_7886,N_5214,N_3151);
and U7887 (N_7887,N_5002,N_3109);
nor U7888 (N_7888,N_4004,N_3517);
xor U7889 (N_7889,N_5280,N_4012);
xor U7890 (N_7890,N_5041,N_4742);
or U7891 (N_7891,N_5763,N_3060);
and U7892 (N_7892,N_4816,N_5680);
nand U7893 (N_7893,N_3065,N_5416);
and U7894 (N_7894,N_4663,N_3931);
nand U7895 (N_7895,N_3639,N_3509);
nor U7896 (N_7896,N_4585,N_5112);
or U7897 (N_7897,N_4758,N_4702);
nand U7898 (N_7898,N_3772,N_4892);
nand U7899 (N_7899,N_4932,N_3184);
nand U7900 (N_7900,N_3161,N_5887);
nor U7901 (N_7901,N_5940,N_5235);
and U7902 (N_7902,N_3203,N_4545);
xnor U7903 (N_7903,N_4302,N_5356);
and U7904 (N_7904,N_3482,N_3113);
xor U7905 (N_7905,N_4208,N_3037);
nor U7906 (N_7906,N_4442,N_3445);
xor U7907 (N_7907,N_3297,N_3293);
and U7908 (N_7908,N_3902,N_4756);
nand U7909 (N_7909,N_4247,N_4903);
and U7910 (N_7910,N_4315,N_4444);
xor U7911 (N_7911,N_3124,N_4985);
xor U7912 (N_7912,N_4856,N_3891);
and U7913 (N_7913,N_3334,N_3355);
xnor U7914 (N_7914,N_4021,N_3447);
nor U7915 (N_7915,N_5428,N_3295);
and U7916 (N_7916,N_3974,N_4951);
and U7917 (N_7917,N_5503,N_3979);
or U7918 (N_7918,N_5667,N_4189);
xnor U7919 (N_7919,N_3989,N_4666);
and U7920 (N_7920,N_3671,N_4912);
nor U7921 (N_7921,N_3688,N_3108);
xor U7922 (N_7922,N_5462,N_3844);
or U7923 (N_7923,N_3928,N_4959);
nor U7924 (N_7924,N_5601,N_5702);
and U7925 (N_7925,N_5870,N_3145);
or U7926 (N_7926,N_5587,N_5204);
and U7927 (N_7927,N_3262,N_4402);
xnor U7928 (N_7928,N_5409,N_3097);
and U7929 (N_7929,N_5522,N_3863);
or U7930 (N_7930,N_5058,N_5808);
xnor U7931 (N_7931,N_4211,N_3666);
and U7932 (N_7932,N_5192,N_5678);
nor U7933 (N_7933,N_5060,N_5780);
nand U7934 (N_7934,N_4106,N_3819);
xnor U7935 (N_7935,N_5135,N_4720);
or U7936 (N_7936,N_4007,N_5401);
xnor U7937 (N_7937,N_4850,N_5433);
nor U7938 (N_7938,N_5595,N_3914);
nor U7939 (N_7939,N_4535,N_3858);
nor U7940 (N_7940,N_4085,N_5681);
and U7941 (N_7941,N_3904,N_3111);
or U7942 (N_7942,N_5793,N_3604);
xnor U7943 (N_7943,N_5971,N_4965);
xnor U7944 (N_7944,N_4725,N_5441);
xnor U7945 (N_7945,N_5708,N_4283);
or U7946 (N_7946,N_3494,N_3461);
nand U7947 (N_7947,N_4744,N_5664);
nor U7948 (N_7948,N_3573,N_4714);
or U7949 (N_7949,N_5023,N_4796);
nor U7950 (N_7950,N_3139,N_5932);
nor U7951 (N_7951,N_5973,N_5599);
or U7952 (N_7952,N_5318,N_3796);
or U7953 (N_7953,N_4975,N_3955);
and U7954 (N_7954,N_5507,N_3199);
xor U7955 (N_7955,N_3624,N_4100);
or U7956 (N_7956,N_5221,N_4863);
xor U7957 (N_7957,N_4396,N_4250);
xnor U7958 (N_7958,N_4252,N_4256);
nor U7959 (N_7959,N_5815,N_3083);
and U7960 (N_7960,N_4722,N_3398);
nor U7961 (N_7961,N_3177,N_4872);
and U7962 (N_7962,N_4210,N_4623);
nor U7963 (N_7963,N_5389,N_5977);
and U7964 (N_7964,N_3441,N_4312);
xor U7965 (N_7965,N_5663,N_5058);
xnor U7966 (N_7966,N_3825,N_4387);
nor U7967 (N_7967,N_3750,N_3718);
xnor U7968 (N_7968,N_3747,N_3504);
and U7969 (N_7969,N_4027,N_3237);
nand U7970 (N_7970,N_3203,N_5974);
and U7971 (N_7971,N_3120,N_4396);
and U7972 (N_7972,N_5969,N_4885);
nand U7973 (N_7973,N_3434,N_4489);
nor U7974 (N_7974,N_5873,N_4278);
nand U7975 (N_7975,N_4054,N_5509);
or U7976 (N_7976,N_4637,N_4587);
or U7977 (N_7977,N_4607,N_5372);
or U7978 (N_7978,N_3154,N_5379);
or U7979 (N_7979,N_3795,N_5516);
and U7980 (N_7980,N_5792,N_4044);
and U7981 (N_7981,N_3239,N_5375);
xor U7982 (N_7982,N_4466,N_5492);
xnor U7983 (N_7983,N_4374,N_5353);
nand U7984 (N_7984,N_4839,N_4985);
and U7985 (N_7985,N_4276,N_4893);
nand U7986 (N_7986,N_4959,N_4215);
or U7987 (N_7987,N_4494,N_4180);
and U7988 (N_7988,N_3381,N_3157);
xnor U7989 (N_7989,N_5912,N_4975);
and U7990 (N_7990,N_5608,N_4476);
nand U7991 (N_7991,N_3079,N_4403);
and U7992 (N_7992,N_4168,N_5970);
or U7993 (N_7993,N_4425,N_5385);
and U7994 (N_7994,N_3859,N_5285);
nor U7995 (N_7995,N_5138,N_3450);
and U7996 (N_7996,N_4690,N_5649);
xnor U7997 (N_7997,N_3706,N_5038);
nand U7998 (N_7998,N_5017,N_5181);
nand U7999 (N_7999,N_5731,N_3139);
or U8000 (N_8000,N_3943,N_5110);
and U8001 (N_8001,N_5022,N_4846);
nand U8002 (N_8002,N_5511,N_4563);
xor U8003 (N_8003,N_3950,N_5788);
or U8004 (N_8004,N_5009,N_4658);
nor U8005 (N_8005,N_4064,N_3739);
nand U8006 (N_8006,N_5978,N_5386);
and U8007 (N_8007,N_3446,N_5124);
xnor U8008 (N_8008,N_3911,N_4265);
or U8009 (N_8009,N_5974,N_5596);
or U8010 (N_8010,N_5499,N_4164);
or U8011 (N_8011,N_4624,N_3254);
and U8012 (N_8012,N_4277,N_3239);
xor U8013 (N_8013,N_3929,N_3642);
and U8014 (N_8014,N_5476,N_3765);
or U8015 (N_8015,N_3767,N_5960);
nand U8016 (N_8016,N_5874,N_5983);
nor U8017 (N_8017,N_5488,N_5457);
xnor U8018 (N_8018,N_5367,N_5998);
xnor U8019 (N_8019,N_4151,N_3472);
or U8020 (N_8020,N_5296,N_5090);
or U8021 (N_8021,N_4401,N_5793);
nand U8022 (N_8022,N_5109,N_5374);
and U8023 (N_8023,N_4021,N_3557);
or U8024 (N_8024,N_4781,N_5465);
and U8025 (N_8025,N_5722,N_3306);
xor U8026 (N_8026,N_4067,N_3721);
and U8027 (N_8027,N_5101,N_5357);
or U8028 (N_8028,N_3860,N_4912);
nand U8029 (N_8029,N_4569,N_3423);
nand U8030 (N_8030,N_5006,N_4927);
nand U8031 (N_8031,N_5262,N_5220);
nand U8032 (N_8032,N_5581,N_5254);
nor U8033 (N_8033,N_4882,N_5004);
nor U8034 (N_8034,N_4291,N_4451);
nand U8035 (N_8035,N_5748,N_5018);
or U8036 (N_8036,N_3888,N_4929);
or U8037 (N_8037,N_4746,N_5105);
and U8038 (N_8038,N_4208,N_3767);
and U8039 (N_8039,N_3398,N_4089);
or U8040 (N_8040,N_4599,N_4878);
and U8041 (N_8041,N_3249,N_5344);
or U8042 (N_8042,N_5558,N_5461);
nor U8043 (N_8043,N_3052,N_5107);
or U8044 (N_8044,N_5457,N_3488);
nand U8045 (N_8045,N_5812,N_5439);
or U8046 (N_8046,N_3285,N_3364);
nand U8047 (N_8047,N_3297,N_3434);
xor U8048 (N_8048,N_3871,N_4564);
nor U8049 (N_8049,N_5967,N_3864);
nand U8050 (N_8050,N_4892,N_4747);
nor U8051 (N_8051,N_4574,N_4668);
nand U8052 (N_8052,N_4563,N_5603);
or U8053 (N_8053,N_4444,N_3723);
nor U8054 (N_8054,N_4812,N_4271);
nor U8055 (N_8055,N_3819,N_5318);
nand U8056 (N_8056,N_5273,N_4435);
nand U8057 (N_8057,N_4438,N_3017);
nand U8058 (N_8058,N_4891,N_3398);
and U8059 (N_8059,N_4352,N_3327);
nand U8060 (N_8060,N_5442,N_3428);
and U8061 (N_8061,N_4861,N_5305);
nand U8062 (N_8062,N_3202,N_5613);
xor U8063 (N_8063,N_5607,N_4412);
or U8064 (N_8064,N_4234,N_5392);
or U8065 (N_8065,N_5600,N_5013);
nor U8066 (N_8066,N_5501,N_3282);
xnor U8067 (N_8067,N_3277,N_5781);
or U8068 (N_8068,N_3433,N_3323);
nand U8069 (N_8069,N_4694,N_5937);
and U8070 (N_8070,N_4895,N_4285);
and U8071 (N_8071,N_5674,N_3433);
nor U8072 (N_8072,N_5074,N_4631);
xnor U8073 (N_8073,N_5408,N_4186);
and U8074 (N_8074,N_4037,N_5070);
nand U8075 (N_8075,N_4217,N_5147);
xnor U8076 (N_8076,N_4058,N_5872);
or U8077 (N_8077,N_4244,N_5726);
and U8078 (N_8078,N_5315,N_3379);
or U8079 (N_8079,N_5834,N_5166);
and U8080 (N_8080,N_4928,N_5873);
xor U8081 (N_8081,N_5438,N_3272);
xor U8082 (N_8082,N_5843,N_3811);
nand U8083 (N_8083,N_4580,N_5285);
or U8084 (N_8084,N_4287,N_5156);
xnor U8085 (N_8085,N_5165,N_4091);
xnor U8086 (N_8086,N_3616,N_4524);
xor U8087 (N_8087,N_5257,N_4115);
nor U8088 (N_8088,N_5060,N_4345);
nor U8089 (N_8089,N_5487,N_5273);
nor U8090 (N_8090,N_3212,N_4322);
nor U8091 (N_8091,N_3230,N_3467);
nand U8092 (N_8092,N_4139,N_3719);
nand U8093 (N_8093,N_3581,N_5692);
nand U8094 (N_8094,N_3216,N_3224);
xnor U8095 (N_8095,N_4409,N_4967);
and U8096 (N_8096,N_3607,N_3370);
nor U8097 (N_8097,N_5917,N_3978);
and U8098 (N_8098,N_4565,N_4490);
nand U8099 (N_8099,N_4016,N_4430);
or U8100 (N_8100,N_4138,N_3282);
or U8101 (N_8101,N_3257,N_4788);
nand U8102 (N_8102,N_4366,N_5221);
xor U8103 (N_8103,N_4741,N_3278);
or U8104 (N_8104,N_3956,N_4512);
and U8105 (N_8105,N_4315,N_4920);
nor U8106 (N_8106,N_3086,N_4563);
xnor U8107 (N_8107,N_3686,N_3563);
nand U8108 (N_8108,N_5133,N_3398);
or U8109 (N_8109,N_4976,N_3763);
nor U8110 (N_8110,N_3733,N_4633);
nor U8111 (N_8111,N_5257,N_5535);
nand U8112 (N_8112,N_3526,N_4939);
nand U8113 (N_8113,N_4767,N_4170);
and U8114 (N_8114,N_3197,N_4021);
nand U8115 (N_8115,N_3350,N_5838);
and U8116 (N_8116,N_3476,N_5989);
nor U8117 (N_8117,N_4487,N_3692);
or U8118 (N_8118,N_5590,N_3365);
and U8119 (N_8119,N_4109,N_3646);
and U8120 (N_8120,N_5399,N_4883);
nand U8121 (N_8121,N_5363,N_3127);
and U8122 (N_8122,N_3054,N_5116);
or U8123 (N_8123,N_5095,N_3421);
and U8124 (N_8124,N_4078,N_4169);
nand U8125 (N_8125,N_5858,N_3997);
nor U8126 (N_8126,N_4440,N_5979);
xnor U8127 (N_8127,N_3301,N_5409);
xor U8128 (N_8128,N_4309,N_3653);
xnor U8129 (N_8129,N_4460,N_4153);
or U8130 (N_8130,N_3832,N_4266);
or U8131 (N_8131,N_4152,N_5303);
nor U8132 (N_8132,N_4102,N_4168);
xnor U8133 (N_8133,N_5016,N_3199);
nand U8134 (N_8134,N_3367,N_5597);
nor U8135 (N_8135,N_3128,N_3212);
xnor U8136 (N_8136,N_4176,N_5842);
nor U8137 (N_8137,N_3716,N_5719);
or U8138 (N_8138,N_5978,N_5761);
or U8139 (N_8139,N_4879,N_4370);
nand U8140 (N_8140,N_3625,N_3783);
or U8141 (N_8141,N_5827,N_4911);
nand U8142 (N_8142,N_3321,N_4430);
and U8143 (N_8143,N_3468,N_3773);
xnor U8144 (N_8144,N_4365,N_3422);
and U8145 (N_8145,N_5120,N_5311);
and U8146 (N_8146,N_4289,N_4526);
or U8147 (N_8147,N_3961,N_4297);
nand U8148 (N_8148,N_5609,N_5614);
or U8149 (N_8149,N_3676,N_5420);
nor U8150 (N_8150,N_3481,N_4744);
nor U8151 (N_8151,N_3335,N_3285);
and U8152 (N_8152,N_5653,N_3939);
nand U8153 (N_8153,N_4669,N_5262);
or U8154 (N_8154,N_5407,N_3558);
nor U8155 (N_8155,N_4653,N_3759);
nand U8156 (N_8156,N_3822,N_3324);
nor U8157 (N_8157,N_4399,N_3021);
nand U8158 (N_8158,N_5671,N_5726);
and U8159 (N_8159,N_4692,N_5372);
or U8160 (N_8160,N_3499,N_3707);
nand U8161 (N_8161,N_5088,N_3861);
or U8162 (N_8162,N_4183,N_5377);
nor U8163 (N_8163,N_3560,N_5948);
and U8164 (N_8164,N_4264,N_4963);
xor U8165 (N_8165,N_5022,N_5891);
or U8166 (N_8166,N_4610,N_4252);
nand U8167 (N_8167,N_5767,N_5625);
nor U8168 (N_8168,N_3473,N_4155);
nor U8169 (N_8169,N_5963,N_5306);
nand U8170 (N_8170,N_5302,N_5239);
and U8171 (N_8171,N_5644,N_5670);
xor U8172 (N_8172,N_3470,N_3933);
nand U8173 (N_8173,N_4484,N_3115);
and U8174 (N_8174,N_3898,N_4503);
xor U8175 (N_8175,N_4278,N_5830);
or U8176 (N_8176,N_5384,N_4503);
and U8177 (N_8177,N_3278,N_4159);
and U8178 (N_8178,N_4172,N_5464);
and U8179 (N_8179,N_4920,N_3338);
nor U8180 (N_8180,N_5560,N_5096);
nor U8181 (N_8181,N_4695,N_3271);
or U8182 (N_8182,N_4870,N_3116);
or U8183 (N_8183,N_4938,N_4742);
xor U8184 (N_8184,N_3192,N_5759);
nand U8185 (N_8185,N_4644,N_4391);
or U8186 (N_8186,N_4400,N_3551);
nor U8187 (N_8187,N_4418,N_5393);
and U8188 (N_8188,N_3045,N_4799);
xnor U8189 (N_8189,N_4988,N_5252);
xor U8190 (N_8190,N_5408,N_4060);
or U8191 (N_8191,N_5592,N_5255);
xor U8192 (N_8192,N_5449,N_5651);
nand U8193 (N_8193,N_4853,N_4147);
nor U8194 (N_8194,N_4295,N_4688);
and U8195 (N_8195,N_3934,N_4687);
and U8196 (N_8196,N_3483,N_3237);
nor U8197 (N_8197,N_4566,N_4994);
and U8198 (N_8198,N_3162,N_5698);
nand U8199 (N_8199,N_5934,N_5395);
xor U8200 (N_8200,N_5753,N_3173);
xnor U8201 (N_8201,N_5702,N_4829);
and U8202 (N_8202,N_5991,N_4378);
nor U8203 (N_8203,N_5199,N_4526);
nor U8204 (N_8204,N_4553,N_3102);
nand U8205 (N_8205,N_5070,N_4703);
xnor U8206 (N_8206,N_3530,N_4283);
xor U8207 (N_8207,N_5461,N_5065);
and U8208 (N_8208,N_4756,N_5969);
xnor U8209 (N_8209,N_4849,N_3703);
nand U8210 (N_8210,N_4886,N_4969);
xor U8211 (N_8211,N_5372,N_5125);
xor U8212 (N_8212,N_4438,N_3242);
or U8213 (N_8213,N_5337,N_4836);
nand U8214 (N_8214,N_5463,N_3116);
or U8215 (N_8215,N_4522,N_5622);
or U8216 (N_8216,N_3624,N_4508);
nand U8217 (N_8217,N_3454,N_5216);
nor U8218 (N_8218,N_3365,N_5625);
nand U8219 (N_8219,N_4631,N_5825);
xor U8220 (N_8220,N_5480,N_3407);
xor U8221 (N_8221,N_3213,N_5815);
xnor U8222 (N_8222,N_4184,N_5309);
or U8223 (N_8223,N_4336,N_5971);
and U8224 (N_8224,N_4897,N_4316);
nand U8225 (N_8225,N_4411,N_3084);
nand U8226 (N_8226,N_5446,N_5634);
or U8227 (N_8227,N_4697,N_4924);
and U8228 (N_8228,N_5344,N_4604);
or U8229 (N_8229,N_5027,N_5140);
or U8230 (N_8230,N_3163,N_4630);
and U8231 (N_8231,N_3815,N_4960);
nor U8232 (N_8232,N_3029,N_4405);
and U8233 (N_8233,N_4491,N_5382);
nand U8234 (N_8234,N_3927,N_3236);
nand U8235 (N_8235,N_5832,N_4453);
nor U8236 (N_8236,N_4167,N_3011);
or U8237 (N_8237,N_3729,N_4051);
and U8238 (N_8238,N_3319,N_5160);
or U8239 (N_8239,N_4474,N_5498);
nor U8240 (N_8240,N_4705,N_3539);
and U8241 (N_8241,N_3338,N_4910);
and U8242 (N_8242,N_4253,N_4036);
and U8243 (N_8243,N_4618,N_5839);
nor U8244 (N_8244,N_5708,N_5795);
and U8245 (N_8245,N_3224,N_3945);
or U8246 (N_8246,N_5460,N_4509);
nor U8247 (N_8247,N_4726,N_3117);
xor U8248 (N_8248,N_4883,N_5065);
and U8249 (N_8249,N_5815,N_3006);
nor U8250 (N_8250,N_5984,N_4413);
xor U8251 (N_8251,N_3865,N_5033);
nand U8252 (N_8252,N_5794,N_4882);
nand U8253 (N_8253,N_5407,N_4968);
or U8254 (N_8254,N_3729,N_3206);
nor U8255 (N_8255,N_5956,N_3042);
or U8256 (N_8256,N_3916,N_4265);
and U8257 (N_8257,N_3603,N_5394);
xnor U8258 (N_8258,N_4604,N_5506);
nor U8259 (N_8259,N_4363,N_5826);
xor U8260 (N_8260,N_5343,N_3669);
nand U8261 (N_8261,N_3884,N_5703);
nand U8262 (N_8262,N_3437,N_5626);
and U8263 (N_8263,N_4446,N_4147);
and U8264 (N_8264,N_4273,N_5317);
and U8265 (N_8265,N_4132,N_3928);
xnor U8266 (N_8266,N_3105,N_5495);
or U8267 (N_8267,N_4153,N_4840);
or U8268 (N_8268,N_4055,N_4998);
and U8269 (N_8269,N_4059,N_4619);
and U8270 (N_8270,N_4666,N_5885);
xor U8271 (N_8271,N_5226,N_5353);
nand U8272 (N_8272,N_3391,N_3535);
or U8273 (N_8273,N_3935,N_3187);
and U8274 (N_8274,N_5708,N_4203);
xor U8275 (N_8275,N_3497,N_5974);
nor U8276 (N_8276,N_4756,N_5968);
xor U8277 (N_8277,N_5304,N_4057);
and U8278 (N_8278,N_3944,N_3311);
nand U8279 (N_8279,N_5762,N_3671);
and U8280 (N_8280,N_3631,N_5048);
or U8281 (N_8281,N_4990,N_3636);
and U8282 (N_8282,N_3238,N_4458);
and U8283 (N_8283,N_4267,N_5530);
and U8284 (N_8284,N_3424,N_3719);
nor U8285 (N_8285,N_3308,N_4259);
xnor U8286 (N_8286,N_3503,N_3697);
or U8287 (N_8287,N_5701,N_5274);
xnor U8288 (N_8288,N_4886,N_3215);
or U8289 (N_8289,N_5013,N_3374);
nor U8290 (N_8290,N_4603,N_5308);
nor U8291 (N_8291,N_3010,N_3888);
xor U8292 (N_8292,N_3711,N_5316);
or U8293 (N_8293,N_5352,N_4308);
and U8294 (N_8294,N_5604,N_5048);
and U8295 (N_8295,N_4116,N_5143);
or U8296 (N_8296,N_4219,N_5017);
or U8297 (N_8297,N_4999,N_5922);
nand U8298 (N_8298,N_5363,N_4620);
nor U8299 (N_8299,N_4724,N_4764);
nor U8300 (N_8300,N_5555,N_4966);
and U8301 (N_8301,N_4333,N_3060);
xor U8302 (N_8302,N_3747,N_5182);
or U8303 (N_8303,N_5000,N_5960);
xor U8304 (N_8304,N_5663,N_3226);
xnor U8305 (N_8305,N_5225,N_3348);
xnor U8306 (N_8306,N_3382,N_4209);
and U8307 (N_8307,N_3185,N_4828);
xnor U8308 (N_8308,N_5623,N_4097);
xor U8309 (N_8309,N_4863,N_5570);
nor U8310 (N_8310,N_4953,N_3498);
or U8311 (N_8311,N_3907,N_5479);
nor U8312 (N_8312,N_3555,N_5514);
nand U8313 (N_8313,N_3895,N_4477);
xor U8314 (N_8314,N_4901,N_5513);
and U8315 (N_8315,N_4871,N_5589);
nor U8316 (N_8316,N_3451,N_3031);
and U8317 (N_8317,N_5394,N_4099);
xor U8318 (N_8318,N_4881,N_3422);
or U8319 (N_8319,N_4309,N_3349);
or U8320 (N_8320,N_3962,N_4559);
nand U8321 (N_8321,N_3979,N_5048);
nand U8322 (N_8322,N_4930,N_5900);
nand U8323 (N_8323,N_3105,N_3239);
xor U8324 (N_8324,N_5530,N_4128);
and U8325 (N_8325,N_4638,N_3414);
or U8326 (N_8326,N_3167,N_3779);
and U8327 (N_8327,N_3565,N_4680);
or U8328 (N_8328,N_4425,N_4429);
xnor U8329 (N_8329,N_4853,N_4646);
or U8330 (N_8330,N_3281,N_3929);
and U8331 (N_8331,N_5069,N_5129);
or U8332 (N_8332,N_3303,N_3635);
xnor U8333 (N_8333,N_4360,N_5317);
nand U8334 (N_8334,N_5019,N_3666);
or U8335 (N_8335,N_5887,N_5985);
or U8336 (N_8336,N_5057,N_4758);
nand U8337 (N_8337,N_5504,N_5560);
xnor U8338 (N_8338,N_3403,N_3600);
and U8339 (N_8339,N_4001,N_5852);
nand U8340 (N_8340,N_3861,N_5272);
or U8341 (N_8341,N_3470,N_4327);
nand U8342 (N_8342,N_5737,N_5892);
nor U8343 (N_8343,N_5755,N_3510);
nand U8344 (N_8344,N_4911,N_4229);
and U8345 (N_8345,N_4013,N_5784);
xor U8346 (N_8346,N_5071,N_3315);
nand U8347 (N_8347,N_3834,N_3958);
nand U8348 (N_8348,N_5580,N_4005);
xor U8349 (N_8349,N_3922,N_3623);
nand U8350 (N_8350,N_5949,N_4967);
nor U8351 (N_8351,N_4278,N_4618);
and U8352 (N_8352,N_5272,N_5403);
nand U8353 (N_8353,N_4475,N_3776);
and U8354 (N_8354,N_4404,N_5385);
nor U8355 (N_8355,N_3492,N_3718);
or U8356 (N_8356,N_4955,N_4575);
nand U8357 (N_8357,N_3662,N_4474);
or U8358 (N_8358,N_4344,N_4467);
and U8359 (N_8359,N_5046,N_4484);
or U8360 (N_8360,N_3363,N_5824);
nand U8361 (N_8361,N_3070,N_5026);
and U8362 (N_8362,N_5916,N_5428);
nor U8363 (N_8363,N_4981,N_5598);
nor U8364 (N_8364,N_3961,N_3050);
nor U8365 (N_8365,N_5307,N_5948);
xor U8366 (N_8366,N_3572,N_5322);
xor U8367 (N_8367,N_5085,N_3163);
xnor U8368 (N_8368,N_4796,N_4998);
and U8369 (N_8369,N_4058,N_3542);
nand U8370 (N_8370,N_5181,N_4665);
or U8371 (N_8371,N_3357,N_3321);
or U8372 (N_8372,N_3465,N_5513);
and U8373 (N_8373,N_5707,N_3931);
nand U8374 (N_8374,N_3627,N_4063);
or U8375 (N_8375,N_4333,N_5978);
nor U8376 (N_8376,N_5897,N_5130);
and U8377 (N_8377,N_5501,N_5156);
or U8378 (N_8378,N_4043,N_3490);
nand U8379 (N_8379,N_4456,N_4773);
and U8380 (N_8380,N_3369,N_5906);
and U8381 (N_8381,N_3733,N_3592);
or U8382 (N_8382,N_4978,N_3844);
and U8383 (N_8383,N_3404,N_5052);
and U8384 (N_8384,N_3957,N_3488);
xor U8385 (N_8385,N_3078,N_4310);
nor U8386 (N_8386,N_3780,N_3756);
or U8387 (N_8387,N_5630,N_3938);
and U8388 (N_8388,N_4725,N_5914);
nand U8389 (N_8389,N_3562,N_3069);
xor U8390 (N_8390,N_4568,N_3533);
or U8391 (N_8391,N_3470,N_5414);
and U8392 (N_8392,N_3347,N_3645);
and U8393 (N_8393,N_5830,N_3669);
nor U8394 (N_8394,N_3760,N_4869);
nand U8395 (N_8395,N_4356,N_4635);
nor U8396 (N_8396,N_4423,N_4467);
xor U8397 (N_8397,N_5276,N_3435);
nand U8398 (N_8398,N_5863,N_3069);
nand U8399 (N_8399,N_3781,N_3514);
and U8400 (N_8400,N_3132,N_3300);
or U8401 (N_8401,N_4082,N_3490);
xnor U8402 (N_8402,N_5315,N_3793);
xor U8403 (N_8403,N_4256,N_4845);
and U8404 (N_8404,N_4057,N_4616);
and U8405 (N_8405,N_5584,N_5100);
xnor U8406 (N_8406,N_4773,N_5474);
and U8407 (N_8407,N_3223,N_3925);
or U8408 (N_8408,N_4611,N_5892);
and U8409 (N_8409,N_3943,N_3178);
nor U8410 (N_8410,N_5015,N_3734);
nand U8411 (N_8411,N_5972,N_4926);
nor U8412 (N_8412,N_5125,N_5437);
xor U8413 (N_8413,N_4938,N_4563);
nor U8414 (N_8414,N_3762,N_5798);
xor U8415 (N_8415,N_4746,N_5982);
xnor U8416 (N_8416,N_4308,N_4437);
xnor U8417 (N_8417,N_3412,N_4143);
or U8418 (N_8418,N_3441,N_5543);
and U8419 (N_8419,N_5132,N_3086);
and U8420 (N_8420,N_4589,N_4767);
and U8421 (N_8421,N_5415,N_5332);
and U8422 (N_8422,N_3046,N_5139);
nand U8423 (N_8423,N_5620,N_3306);
xnor U8424 (N_8424,N_5295,N_4274);
nor U8425 (N_8425,N_4738,N_4284);
xor U8426 (N_8426,N_5557,N_4206);
nor U8427 (N_8427,N_5087,N_3573);
or U8428 (N_8428,N_3443,N_5994);
nor U8429 (N_8429,N_4205,N_4059);
nor U8430 (N_8430,N_5524,N_5459);
xnor U8431 (N_8431,N_3497,N_5399);
nor U8432 (N_8432,N_3063,N_5970);
xnor U8433 (N_8433,N_5008,N_5070);
nand U8434 (N_8434,N_5824,N_3730);
nor U8435 (N_8435,N_5221,N_4983);
nor U8436 (N_8436,N_5651,N_5654);
nor U8437 (N_8437,N_5452,N_3813);
nand U8438 (N_8438,N_5777,N_4012);
or U8439 (N_8439,N_4346,N_4826);
and U8440 (N_8440,N_3751,N_5268);
nand U8441 (N_8441,N_5825,N_5235);
or U8442 (N_8442,N_3434,N_5768);
and U8443 (N_8443,N_5964,N_3736);
or U8444 (N_8444,N_4317,N_3450);
or U8445 (N_8445,N_3555,N_4590);
xor U8446 (N_8446,N_3673,N_5558);
nand U8447 (N_8447,N_3639,N_5896);
nand U8448 (N_8448,N_5700,N_4043);
nand U8449 (N_8449,N_4403,N_5272);
nor U8450 (N_8450,N_3631,N_4316);
and U8451 (N_8451,N_5720,N_5613);
nand U8452 (N_8452,N_4204,N_4410);
or U8453 (N_8453,N_4678,N_5334);
nor U8454 (N_8454,N_5007,N_3524);
nand U8455 (N_8455,N_5288,N_3573);
nand U8456 (N_8456,N_4446,N_5326);
nor U8457 (N_8457,N_3649,N_3496);
or U8458 (N_8458,N_3815,N_4531);
and U8459 (N_8459,N_3275,N_3958);
or U8460 (N_8460,N_4650,N_4210);
or U8461 (N_8461,N_4019,N_5861);
and U8462 (N_8462,N_3875,N_3244);
or U8463 (N_8463,N_4763,N_4383);
nand U8464 (N_8464,N_4905,N_5196);
nor U8465 (N_8465,N_4199,N_4072);
and U8466 (N_8466,N_3611,N_3801);
or U8467 (N_8467,N_5312,N_4637);
or U8468 (N_8468,N_5412,N_3041);
and U8469 (N_8469,N_4007,N_3652);
or U8470 (N_8470,N_5897,N_5017);
and U8471 (N_8471,N_4566,N_4370);
or U8472 (N_8472,N_5541,N_4786);
or U8473 (N_8473,N_3582,N_4437);
xor U8474 (N_8474,N_5635,N_5986);
xnor U8475 (N_8475,N_3830,N_3179);
or U8476 (N_8476,N_3228,N_3540);
nor U8477 (N_8477,N_5600,N_4821);
nand U8478 (N_8478,N_4948,N_5685);
xor U8479 (N_8479,N_4006,N_5743);
or U8480 (N_8480,N_4901,N_3037);
nand U8481 (N_8481,N_3143,N_5351);
nand U8482 (N_8482,N_3616,N_4515);
xor U8483 (N_8483,N_4486,N_3448);
xnor U8484 (N_8484,N_5497,N_5902);
xnor U8485 (N_8485,N_3101,N_5138);
and U8486 (N_8486,N_3295,N_5786);
nand U8487 (N_8487,N_3971,N_4438);
xor U8488 (N_8488,N_3631,N_3098);
nor U8489 (N_8489,N_3520,N_3844);
or U8490 (N_8490,N_3932,N_5148);
nand U8491 (N_8491,N_5345,N_3116);
or U8492 (N_8492,N_3271,N_4394);
xnor U8493 (N_8493,N_3494,N_5290);
xnor U8494 (N_8494,N_5126,N_3894);
xnor U8495 (N_8495,N_3142,N_5321);
nand U8496 (N_8496,N_5103,N_5854);
or U8497 (N_8497,N_3969,N_5195);
or U8498 (N_8498,N_5792,N_5919);
xor U8499 (N_8499,N_4206,N_4395);
nor U8500 (N_8500,N_4374,N_5710);
nor U8501 (N_8501,N_3155,N_4791);
nand U8502 (N_8502,N_4858,N_3224);
nand U8503 (N_8503,N_5783,N_4445);
xor U8504 (N_8504,N_4942,N_4900);
or U8505 (N_8505,N_5401,N_4163);
xnor U8506 (N_8506,N_4163,N_3604);
and U8507 (N_8507,N_3244,N_5787);
or U8508 (N_8508,N_3946,N_3667);
nand U8509 (N_8509,N_4966,N_5911);
and U8510 (N_8510,N_4452,N_3440);
nand U8511 (N_8511,N_4718,N_4988);
nand U8512 (N_8512,N_3045,N_3917);
or U8513 (N_8513,N_3690,N_5978);
and U8514 (N_8514,N_5120,N_5036);
nand U8515 (N_8515,N_5022,N_3706);
and U8516 (N_8516,N_3447,N_5515);
nor U8517 (N_8517,N_3693,N_3708);
nand U8518 (N_8518,N_3507,N_3542);
or U8519 (N_8519,N_3347,N_3966);
nand U8520 (N_8520,N_4343,N_4054);
nor U8521 (N_8521,N_3291,N_5278);
or U8522 (N_8522,N_4818,N_5949);
and U8523 (N_8523,N_5986,N_3614);
nand U8524 (N_8524,N_4771,N_4707);
and U8525 (N_8525,N_4258,N_3401);
nand U8526 (N_8526,N_4519,N_5213);
and U8527 (N_8527,N_3518,N_5931);
xnor U8528 (N_8528,N_4938,N_4550);
or U8529 (N_8529,N_4789,N_3386);
xor U8530 (N_8530,N_5065,N_3405);
xnor U8531 (N_8531,N_5330,N_3413);
or U8532 (N_8532,N_4515,N_5931);
or U8533 (N_8533,N_3729,N_4729);
or U8534 (N_8534,N_5389,N_4681);
and U8535 (N_8535,N_5136,N_5313);
or U8536 (N_8536,N_4216,N_3965);
nor U8537 (N_8537,N_5756,N_5103);
and U8538 (N_8538,N_4813,N_3996);
and U8539 (N_8539,N_4718,N_3406);
and U8540 (N_8540,N_4260,N_4297);
or U8541 (N_8541,N_3770,N_3662);
or U8542 (N_8542,N_3813,N_3802);
or U8543 (N_8543,N_3929,N_3195);
and U8544 (N_8544,N_4311,N_3716);
or U8545 (N_8545,N_3321,N_4539);
xnor U8546 (N_8546,N_3516,N_3515);
and U8547 (N_8547,N_5231,N_3727);
nor U8548 (N_8548,N_5394,N_4165);
and U8549 (N_8549,N_3093,N_4247);
xor U8550 (N_8550,N_3087,N_5526);
nor U8551 (N_8551,N_4284,N_4085);
and U8552 (N_8552,N_3876,N_4676);
nand U8553 (N_8553,N_3302,N_3639);
xnor U8554 (N_8554,N_5200,N_3917);
nor U8555 (N_8555,N_5392,N_3555);
nand U8556 (N_8556,N_4252,N_5988);
nor U8557 (N_8557,N_5035,N_5016);
and U8558 (N_8558,N_5868,N_3517);
or U8559 (N_8559,N_5438,N_3431);
nand U8560 (N_8560,N_4015,N_5074);
nor U8561 (N_8561,N_3463,N_5849);
or U8562 (N_8562,N_3979,N_3189);
nand U8563 (N_8563,N_3371,N_3986);
xnor U8564 (N_8564,N_5298,N_3457);
nor U8565 (N_8565,N_4041,N_5595);
nor U8566 (N_8566,N_5505,N_5709);
nand U8567 (N_8567,N_4841,N_4792);
nor U8568 (N_8568,N_3234,N_3802);
or U8569 (N_8569,N_4056,N_5197);
or U8570 (N_8570,N_5291,N_3815);
nor U8571 (N_8571,N_5432,N_3563);
nand U8572 (N_8572,N_4487,N_5035);
and U8573 (N_8573,N_5251,N_4298);
nand U8574 (N_8574,N_4216,N_4196);
and U8575 (N_8575,N_3040,N_4462);
nand U8576 (N_8576,N_3145,N_4931);
nand U8577 (N_8577,N_3027,N_3153);
or U8578 (N_8578,N_4067,N_5749);
or U8579 (N_8579,N_3552,N_3024);
and U8580 (N_8580,N_3378,N_3077);
nand U8581 (N_8581,N_4921,N_5060);
nand U8582 (N_8582,N_3955,N_3251);
xnor U8583 (N_8583,N_5048,N_4789);
or U8584 (N_8584,N_5795,N_5344);
nor U8585 (N_8585,N_5958,N_5582);
nor U8586 (N_8586,N_4276,N_4617);
or U8587 (N_8587,N_5460,N_3556);
nand U8588 (N_8588,N_4285,N_3409);
or U8589 (N_8589,N_4164,N_5838);
or U8590 (N_8590,N_5371,N_5780);
and U8591 (N_8591,N_5961,N_5736);
xor U8592 (N_8592,N_5389,N_5019);
nand U8593 (N_8593,N_3700,N_5093);
nand U8594 (N_8594,N_4862,N_4181);
xor U8595 (N_8595,N_4887,N_5673);
nand U8596 (N_8596,N_3438,N_4120);
nand U8597 (N_8597,N_4064,N_3197);
or U8598 (N_8598,N_4110,N_4086);
nand U8599 (N_8599,N_5041,N_4123);
xor U8600 (N_8600,N_3901,N_3752);
xnor U8601 (N_8601,N_3186,N_5532);
xor U8602 (N_8602,N_5513,N_3368);
nand U8603 (N_8603,N_5591,N_4884);
or U8604 (N_8604,N_5865,N_4689);
and U8605 (N_8605,N_5513,N_5796);
nor U8606 (N_8606,N_4432,N_5591);
nand U8607 (N_8607,N_5608,N_4071);
or U8608 (N_8608,N_4111,N_4945);
nand U8609 (N_8609,N_4976,N_4085);
xor U8610 (N_8610,N_4320,N_3131);
nand U8611 (N_8611,N_5266,N_5066);
and U8612 (N_8612,N_3724,N_5718);
nor U8613 (N_8613,N_4242,N_3377);
xnor U8614 (N_8614,N_4255,N_3349);
nand U8615 (N_8615,N_5956,N_4338);
nor U8616 (N_8616,N_4880,N_3779);
nand U8617 (N_8617,N_4662,N_4220);
nand U8618 (N_8618,N_5535,N_3546);
xor U8619 (N_8619,N_3060,N_5765);
xnor U8620 (N_8620,N_4032,N_4828);
nand U8621 (N_8621,N_5647,N_4606);
nor U8622 (N_8622,N_4890,N_4873);
xnor U8623 (N_8623,N_4204,N_4352);
and U8624 (N_8624,N_5328,N_3817);
and U8625 (N_8625,N_3568,N_4435);
xor U8626 (N_8626,N_4752,N_4645);
nand U8627 (N_8627,N_5922,N_5269);
or U8628 (N_8628,N_5872,N_3649);
or U8629 (N_8629,N_4504,N_5712);
and U8630 (N_8630,N_5570,N_4557);
nor U8631 (N_8631,N_4380,N_3704);
or U8632 (N_8632,N_5674,N_5085);
and U8633 (N_8633,N_3362,N_3686);
nand U8634 (N_8634,N_5593,N_5265);
nand U8635 (N_8635,N_4465,N_4836);
xor U8636 (N_8636,N_5967,N_3176);
nand U8637 (N_8637,N_5551,N_4067);
xnor U8638 (N_8638,N_4452,N_5756);
and U8639 (N_8639,N_5007,N_4059);
or U8640 (N_8640,N_5417,N_3302);
nand U8641 (N_8641,N_4453,N_3874);
xor U8642 (N_8642,N_5937,N_3706);
or U8643 (N_8643,N_4297,N_5003);
nand U8644 (N_8644,N_3821,N_5149);
nand U8645 (N_8645,N_4537,N_5001);
or U8646 (N_8646,N_3485,N_4580);
or U8647 (N_8647,N_3035,N_4513);
and U8648 (N_8648,N_4692,N_3310);
nand U8649 (N_8649,N_4030,N_5892);
nand U8650 (N_8650,N_5820,N_4432);
and U8651 (N_8651,N_4312,N_5167);
and U8652 (N_8652,N_3757,N_4739);
nor U8653 (N_8653,N_5706,N_5817);
nor U8654 (N_8654,N_4838,N_4806);
nand U8655 (N_8655,N_4165,N_3771);
or U8656 (N_8656,N_4058,N_4023);
and U8657 (N_8657,N_4809,N_4080);
nor U8658 (N_8658,N_5337,N_4789);
and U8659 (N_8659,N_4485,N_5957);
nor U8660 (N_8660,N_5245,N_3123);
or U8661 (N_8661,N_5489,N_4521);
nand U8662 (N_8662,N_4493,N_4393);
nand U8663 (N_8663,N_3330,N_5767);
nand U8664 (N_8664,N_3950,N_5340);
and U8665 (N_8665,N_4805,N_5939);
nor U8666 (N_8666,N_4324,N_3486);
xnor U8667 (N_8667,N_4932,N_3634);
nor U8668 (N_8668,N_5457,N_3231);
nand U8669 (N_8669,N_5138,N_5628);
xnor U8670 (N_8670,N_3594,N_5090);
xor U8671 (N_8671,N_5184,N_5988);
nor U8672 (N_8672,N_4743,N_5504);
and U8673 (N_8673,N_3597,N_5860);
nand U8674 (N_8674,N_3108,N_4268);
xor U8675 (N_8675,N_5963,N_5804);
and U8676 (N_8676,N_5051,N_3505);
nand U8677 (N_8677,N_5587,N_3888);
or U8678 (N_8678,N_3341,N_4245);
nor U8679 (N_8679,N_3401,N_3003);
or U8680 (N_8680,N_5898,N_4029);
xor U8681 (N_8681,N_5641,N_4659);
or U8682 (N_8682,N_5104,N_4934);
xnor U8683 (N_8683,N_4339,N_3036);
nand U8684 (N_8684,N_4342,N_3181);
and U8685 (N_8685,N_4759,N_5865);
and U8686 (N_8686,N_4433,N_3468);
and U8687 (N_8687,N_3291,N_5640);
nor U8688 (N_8688,N_3080,N_4876);
or U8689 (N_8689,N_4259,N_3417);
nand U8690 (N_8690,N_4289,N_5324);
xnor U8691 (N_8691,N_4061,N_4507);
xnor U8692 (N_8692,N_4455,N_4914);
xnor U8693 (N_8693,N_4244,N_5547);
and U8694 (N_8694,N_5334,N_5944);
or U8695 (N_8695,N_4795,N_5834);
and U8696 (N_8696,N_5983,N_4353);
or U8697 (N_8697,N_5299,N_5690);
xnor U8698 (N_8698,N_4525,N_3710);
xor U8699 (N_8699,N_3018,N_3489);
and U8700 (N_8700,N_4688,N_5372);
xor U8701 (N_8701,N_5443,N_3795);
nand U8702 (N_8702,N_5749,N_3512);
and U8703 (N_8703,N_3174,N_5127);
and U8704 (N_8704,N_4666,N_5417);
and U8705 (N_8705,N_5188,N_5138);
nand U8706 (N_8706,N_5700,N_3993);
xnor U8707 (N_8707,N_4766,N_3297);
or U8708 (N_8708,N_3570,N_5615);
xnor U8709 (N_8709,N_3852,N_5638);
nor U8710 (N_8710,N_3909,N_3387);
or U8711 (N_8711,N_4040,N_4686);
nor U8712 (N_8712,N_5022,N_3943);
nand U8713 (N_8713,N_3658,N_3446);
nor U8714 (N_8714,N_3515,N_4539);
and U8715 (N_8715,N_5214,N_5137);
or U8716 (N_8716,N_4347,N_5999);
or U8717 (N_8717,N_4944,N_3605);
nand U8718 (N_8718,N_5546,N_5103);
and U8719 (N_8719,N_4868,N_5134);
nand U8720 (N_8720,N_4130,N_3493);
xor U8721 (N_8721,N_5389,N_3697);
and U8722 (N_8722,N_5994,N_4691);
xor U8723 (N_8723,N_5652,N_3644);
xor U8724 (N_8724,N_4656,N_5404);
nor U8725 (N_8725,N_3179,N_3211);
nor U8726 (N_8726,N_4503,N_4723);
and U8727 (N_8727,N_4616,N_3299);
xor U8728 (N_8728,N_4463,N_5366);
nor U8729 (N_8729,N_3799,N_3540);
nor U8730 (N_8730,N_4360,N_4946);
and U8731 (N_8731,N_5733,N_5098);
nand U8732 (N_8732,N_3645,N_4879);
or U8733 (N_8733,N_3142,N_5961);
or U8734 (N_8734,N_3794,N_5180);
and U8735 (N_8735,N_5169,N_3901);
xnor U8736 (N_8736,N_5463,N_3593);
and U8737 (N_8737,N_3308,N_5449);
nand U8738 (N_8738,N_5479,N_4396);
nand U8739 (N_8739,N_5307,N_4503);
nand U8740 (N_8740,N_5881,N_4670);
xnor U8741 (N_8741,N_3006,N_4013);
or U8742 (N_8742,N_4514,N_4221);
and U8743 (N_8743,N_3450,N_3930);
nor U8744 (N_8744,N_4290,N_5471);
nand U8745 (N_8745,N_5242,N_5659);
xnor U8746 (N_8746,N_5176,N_3895);
nor U8747 (N_8747,N_4102,N_4816);
nor U8748 (N_8748,N_4436,N_5446);
xor U8749 (N_8749,N_4558,N_3922);
nor U8750 (N_8750,N_5749,N_5222);
nand U8751 (N_8751,N_3249,N_5534);
and U8752 (N_8752,N_3624,N_3110);
nand U8753 (N_8753,N_3451,N_3487);
nor U8754 (N_8754,N_4486,N_4473);
nand U8755 (N_8755,N_4085,N_4933);
nor U8756 (N_8756,N_5857,N_3733);
and U8757 (N_8757,N_4040,N_4007);
or U8758 (N_8758,N_5213,N_5349);
nor U8759 (N_8759,N_3601,N_3369);
and U8760 (N_8760,N_5852,N_4530);
nor U8761 (N_8761,N_5587,N_3500);
or U8762 (N_8762,N_3124,N_3229);
and U8763 (N_8763,N_4976,N_5755);
or U8764 (N_8764,N_5585,N_4965);
nor U8765 (N_8765,N_3685,N_4164);
and U8766 (N_8766,N_5638,N_3065);
nor U8767 (N_8767,N_3645,N_4967);
or U8768 (N_8768,N_4026,N_5497);
nand U8769 (N_8769,N_4647,N_4111);
nand U8770 (N_8770,N_5626,N_4807);
and U8771 (N_8771,N_3019,N_5072);
nor U8772 (N_8772,N_4342,N_4764);
nor U8773 (N_8773,N_5232,N_5731);
nor U8774 (N_8774,N_4390,N_5157);
or U8775 (N_8775,N_4259,N_5261);
xnor U8776 (N_8776,N_3674,N_4240);
or U8777 (N_8777,N_3501,N_3653);
xor U8778 (N_8778,N_3284,N_5691);
nor U8779 (N_8779,N_4342,N_5754);
nor U8780 (N_8780,N_4455,N_3314);
or U8781 (N_8781,N_4968,N_3831);
and U8782 (N_8782,N_4669,N_4290);
and U8783 (N_8783,N_3826,N_4792);
and U8784 (N_8784,N_5930,N_5353);
xnor U8785 (N_8785,N_5105,N_5408);
nand U8786 (N_8786,N_4168,N_4714);
and U8787 (N_8787,N_5876,N_4100);
xor U8788 (N_8788,N_3473,N_4824);
nand U8789 (N_8789,N_4654,N_4618);
xor U8790 (N_8790,N_4808,N_5167);
and U8791 (N_8791,N_3756,N_4325);
xor U8792 (N_8792,N_4412,N_3051);
or U8793 (N_8793,N_3425,N_5796);
and U8794 (N_8794,N_3283,N_5597);
and U8795 (N_8795,N_4222,N_5711);
nand U8796 (N_8796,N_5666,N_4233);
xnor U8797 (N_8797,N_5537,N_5895);
xnor U8798 (N_8798,N_3282,N_3565);
xnor U8799 (N_8799,N_3652,N_5394);
or U8800 (N_8800,N_3927,N_5452);
nand U8801 (N_8801,N_3549,N_4936);
xor U8802 (N_8802,N_4338,N_5738);
or U8803 (N_8803,N_3752,N_3949);
or U8804 (N_8804,N_4596,N_3000);
and U8805 (N_8805,N_3850,N_5977);
xnor U8806 (N_8806,N_3919,N_4705);
xor U8807 (N_8807,N_5718,N_4903);
nor U8808 (N_8808,N_5703,N_3971);
or U8809 (N_8809,N_5557,N_5985);
xnor U8810 (N_8810,N_5179,N_5900);
or U8811 (N_8811,N_3162,N_3477);
and U8812 (N_8812,N_4357,N_5629);
xor U8813 (N_8813,N_4266,N_4347);
nand U8814 (N_8814,N_4936,N_3490);
xor U8815 (N_8815,N_4569,N_5008);
nor U8816 (N_8816,N_5571,N_4724);
nand U8817 (N_8817,N_5184,N_5287);
or U8818 (N_8818,N_4105,N_3977);
xor U8819 (N_8819,N_3344,N_5292);
nand U8820 (N_8820,N_3566,N_4671);
and U8821 (N_8821,N_3132,N_5450);
xnor U8822 (N_8822,N_4949,N_3228);
or U8823 (N_8823,N_3391,N_3833);
or U8824 (N_8824,N_5438,N_5614);
xnor U8825 (N_8825,N_5555,N_4670);
nor U8826 (N_8826,N_3516,N_3597);
nand U8827 (N_8827,N_4685,N_5505);
nor U8828 (N_8828,N_3295,N_5703);
xnor U8829 (N_8829,N_3711,N_5149);
or U8830 (N_8830,N_5675,N_3592);
nand U8831 (N_8831,N_5399,N_4296);
nor U8832 (N_8832,N_5766,N_4472);
or U8833 (N_8833,N_5230,N_4622);
xor U8834 (N_8834,N_3008,N_3604);
or U8835 (N_8835,N_4469,N_5549);
nand U8836 (N_8836,N_4463,N_5808);
nor U8837 (N_8837,N_4545,N_3496);
or U8838 (N_8838,N_4716,N_3336);
nand U8839 (N_8839,N_4514,N_5354);
or U8840 (N_8840,N_3656,N_3125);
nand U8841 (N_8841,N_4757,N_5086);
and U8842 (N_8842,N_5331,N_4686);
xor U8843 (N_8843,N_5326,N_3622);
nand U8844 (N_8844,N_5337,N_3121);
nor U8845 (N_8845,N_4635,N_5453);
and U8846 (N_8846,N_5874,N_5995);
nor U8847 (N_8847,N_4953,N_3191);
and U8848 (N_8848,N_3206,N_5913);
nand U8849 (N_8849,N_4679,N_3048);
xnor U8850 (N_8850,N_3865,N_3116);
and U8851 (N_8851,N_4326,N_5316);
xnor U8852 (N_8852,N_3610,N_5958);
xor U8853 (N_8853,N_5762,N_5691);
and U8854 (N_8854,N_5240,N_3957);
or U8855 (N_8855,N_5549,N_3130);
or U8856 (N_8856,N_4843,N_4199);
and U8857 (N_8857,N_3748,N_5803);
and U8858 (N_8858,N_3949,N_3058);
or U8859 (N_8859,N_4936,N_3285);
and U8860 (N_8860,N_5442,N_5137);
and U8861 (N_8861,N_4217,N_4790);
or U8862 (N_8862,N_4294,N_4697);
and U8863 (N_8863,N_3643,N_4968);
xor U8864 (N_8864,N_5697,N_4567);
nor U8865 (N_8865,N_3301,N_5321);
nor U8866 (N_8866,N_3599,N_4222);
xor U8867 (N_8867,N_5007,N_3922);
nor U8868 (N_8868,N_4536,N_3166);
and U8869 (N_8869,N_3307,N_5693);
xor U8870 (N_8870,N_5666,N_4823);
nand U8871 (N_8871,N_4575,N_5580);
xor U8872 (N_8872,N_5700,N_3512);
or U8873 (N_8873,N_5380,N_3249);
and U8874 (N_8874,N_5311,N_3115);
or U8875 (N_8875,N_3307,N_3226);
and U8876 (N_8876,N_3760,N_5929);
xnor U8877 (N_8877,N_5687,N_4844);
or U8878 (N_8878,N_4635,N_5134);
nor U8879 (N_8879,N_3171,N_3537);
nor U8880 (N_8880,N_3470,N_4684);
and U8881 (N_8881,N_4038,N_4914);
xor U8882 (N_8882,N_5819,N_5007);
and U8883 (N_8883,N_4842,N_3004);
nor U8884 (N_8884,N_4714,N_3964);
xnor U8885 (N_8885,N_3496,N_3267);
or U8886 (N_8886,N_4433,N_3831);
or U8887 (N_8887,N_5644,N_3072);
and U8888 (N_8888,N_3337,N_4487);
and U8889 (N_8889,N_3226,N_4395);
nand U8890 (N_8890,N_5329,N_4190);
nor U8891 (N_8891,N_4675,N_3493);
or U8892 (N_8892,N_3110,N_5738);
nor U8893 (N_8893,N_5817,N_3242);
or U8894 (N_8894,N_4535,N_5734);
nand U8895 (N_8895,N_5293,N_5212);
or U8896 (N_8896,N_3231,N_5024);
or U8897 (N_8897,N_4566,N_4104);
nand U8898 (N_8898,N_4318,N_4379);
xnor U8899 (N_8899,N_5070,N_5007);
xnor U8900 (N_8900,N_4510,N_3692);
xor U8901 (N_8901,N_5207,N_5246);
nand U8902 (N_8902,N_5792,N_5688);
and U8903 (N_8903,N_3796,N_4407);
nand U8904 (N_8904,N_3956,N_3359);
nor U8905 (N_8905,N_5593,N_4311);
xor U8906 (N_8906,N_5401,N_4170);
xnor U8907 (N_8907,N_5235,N_5437);
nand U8908 (N_8908,N_3428,N_5167);
and U8909 (N_8909,N_3334,N_3428);
nor U8910 (N_8910,N_3054,N_3142);
nor U8911 (N_8911,N_3440,N_5738);
nand U8912 (N_8912,N_3943,N_3274);
and U8913 (N_8913,N_4352,N_3364);
or U8914 (N_8914,N_5349,N_3467);
nor U8915 (N_8915,N_5819,N_3234);
and U8916 (N_8916,N_5469,N_4949);
or U8917 (N_8917,N_4377,N_3402);
nor U8918 (N_8918,N_5333,N_4275);
xor U8919 (N_8919,N_5976,N_3464);
or U8920 (N_8920,N_5674,N_3326);
and U8921 (N_8921,N_4088,N_4181);
and U8922 (N_8922,N_3459,N_3787);
nor U8923 (N_8923,N_3516,N_5260);
and U8924 (N_8924,N_4394,N_3406);
or U8925 (N_8925,N_5605,N_3582);
xnor U8926 (N_8926,N_4850,N_5782);
or U8927 (N_8927,N_5541,N_5813);
or U8928 (N_8928,N_5588,N_4050);
nor U8929 (N_8929,N_3001,N_5687);
or U8930 (N_8930,N_3784,N_3589);
and U8931 (N_8931,N_5772,N_5754);
nand U8932 (N_8932,N_3542,N_5031);
xnor U8933 (N_8933,N_5839,N_5118);
xnor U8934 (N_8934,N_3407,N_3176);
nor U8935 (N_8935,N_3600,N_3605);
and U8936 (N_8936,N_5716,N_4268);
xor U8937 (N_8937,N_4100,N_3691);
or U8938 (N_8938,N_5740,N_3341);
or U8939 (N_8939,N_3916,N_4451);
xor U8940 (N_8940,N_4038,N_4231);
nor U8941 (N_8941,N_4761,N_5326);
or U8942 (N_8942,N_3229,N_5004);
nand U8943 (N_8943,N_4507,N_4183);
and U8944 (N_8944,N_4432,N_5233);
or U8945 (N_8945,N_4026,N_5706);
and U8946 (N_8946,N_5367,N_4387);
nand U8947 (N_8947,N_5335,N_4803);
and U8948 (N_8948,N_3392,N_5681);
or U8949 (N_8949,N_3810,N_5766);
nand U8950 (N_8950,N_4785,N_5048);
nor U8951 (N_8951,N_4618,N_5174);
and U8952 (N_8952,N_5657,N_5518);
or U8953 (N_8953,N_5750,N_3767);
xnor U8954 (N_8954,N_5912,N_5290);
nand U8955 (N_8955,N_5796,N_5770);
and U8956 (N_8956,N_4177,N_4123);
nand U8957 (N_8957,N_5818,N_3514);
nor U8958 (N_8958,N_5589,N_4124);
xor U8959 (N_8959,N_5099,N_5411);
or U8960 (N_8960,N_3411,N_4937);
nor U8961 (N_8961,N_3389,N_4886);
or U8962 (N_8962,N_5771,N_3795);
or U8963 (N_8963,N_3759,N_4154);
nor U8964 (N_8964,N_5752,N_5666);
nor U8965 (N_8965,N_3072,N_4416);
nor U8966 (N_8966,N_4471,N_4295);
xor U8967 (N_8967,N_4355,N_5575);
and U8968 (N_8968,N_3957,N_5170);
xnor U8969 (N_8969,N_4481,N_5408);
and U8970 (N_8970,N_5502,N_5545);
or U8971 (N_8971,N_4429,N_5072);
nand U8972 (N_8972,N_3880,N_4168);
nor U8973 (N_8973,N_4955,N_4007);
or U8974 (N_8974,N_4329,N_3421);
nor U8975 (N_8975,N_4521,N_5116);
nand U8976 (N_8976,N_3238,N_3650);
or U8977 (N_8977,N_4672,N_3258);
xor U8978 (N_8978,N_5339,N_5930);
nand U8979 (N_8979,N_4714,N_5015);
nand U8980 (N_8980,N_5797,N_3331);
xor U8981 (N_8981,N_4151,N_4928);
or U8982 (N_8982,N_4289,N_3707);
and U8983 (N_8983,N_4910,N_5487);
nor U8984 (N_8984,N_4435,N_4161);
nor U8985 (N_8985,N_4345,N_5155);
or U8986 (N_8986,N_3460,N_4856);
or U8987 (N_8987,N_5813,N_5803);
and U8988 (N_8988,N_4821,N_5947);
and U8989 (N_8989,N_4634,N_5022);
or U8990 (N_8990,N_5353,N_4621);
nor U8991 (N_8991,N_5330,N_3245);
or U8992 (N_8992,N_5252,N_3846);
nand U8993 (N_8993,N_4331,N_4046);
nand U8994 (N_8994,N_3153,N_5928);
and U8995 (N_8995,N_4251,N_4344);
or U8996 (N_8996,N_5376,N_5607);
and U8997 (N_8997,N_3766,N_5150);
or U8998 (N_8998,N_4178,N_5041);
nand U8999 (N_8999,N_5962,N_3480);
nand U9000 (N_9000,N_7663,N_6131);
nor U9001 (N_9001,N_7306,N_6332);
nor U9002 (N_9002,N_7360,N_6691);
and U9003 (N_9003,N_7469,N_8606);
or U9004 (N_9004,N_8819,N_7685);
or U9005 (N_9005,N_7666,N_6046);
and U9006 (N_9006,N_7283,N_8007);
or U9007 (N_9007,N_6783,N_8969);
nand U9008 (N_9008,N_7697,N_6922);
nand U9009 (N_9009,N_8982,N_6883);
nand U9010 (N_9010,N_8126,N_8146);
nand U9011 (N_9011,N_8476,N_8540);
nor U9012 (N_9012,N_8639,N_7181);
or U9013 (N_9013,N_7783,N_8313);
or U9014 (N_9014,N_6649,N_6190);
and U9015 (N_9015,N_8907,N_7852);
xor U9016 (N_9016,N_7453,N_6802);
nand U9017 (N_9017,N_6152,N_8110);
and U9018 (N_9018,N_8025,N_8227);
nor U9019 (N_9019,N_7098,N_8478);
or U9020 (N_9020,N_6757,N_6610);
or U9021 (N_9021,N_6684,N_8927);
xor U9022 (N_9022,N_7848,N_8243);
and U9023 (N_9023,N_6565,N_6656);
xnor U9024 (N_9024,N_7352,N_8936);
nand U9025 (N_9025,N_7755,N_8895);
nor U9026 (N_9026,N_8270,N_8168);
and U9027 (N_9027,N_6384,N_8665);
and U9028 (N_9028,N_6873,N_8357);
or U9029 (N_9029,N_6737,N_6365);
xnor U9030 (N_9030,N_6837,N_8296);
and U9031 (N_9031,N_6741,N_6180);
and U9032 (N_9032,N_8721,N_6943);
xnor U9033 (N_9033,N_8348,N_7792);
nor U9034 (N_9034,N_6371,N_6990);
nor U9035 (N_9035,N_7737,N_8125);
or U9036 (N_9036,N_7325,N_8866);
xor U9037 (N_9037,N_6731,N_6683);
nand U9038 (N_9038,N_6538,N_7738);
nor U9039 (N_9039,N_7412,N_6506);
nand U9040 (N_9040,N_6675,N_6653);
nor U9041 (N_9041,N_6315,N_8507);
xnor U9042 (N_9042,N_6426,N_7134);
xnor U9043 (N_9043,N_8720,N_7950);
nand U9044 (N_9044,N_8477,N_6673);
and U9045 (N_9045,N_7732,N_8200);
nand U9046 (N_9046,N_8998,N_8953);
xnor U9047 (N_9047,N_6068,N_6339);
and U9048 (N_9048,N_8663,N_7119);
or U9049 (N_9049,N_7121,N_7856);
nor U9050 (N_9050,N_6167,N_8627);
nand U9051 (N_9051,N_6377,N_8411);
xnor U9052 (N_9052,N_6210,N_7772);
nand U9053 (N_9053,N_8383,N_8382);
or U9054 (N_9054,N_8643,N_7545);
nand U9055 (N_9055,N_6334,N_8656);
and U9056 (N_9056,N_8033,N_7553);
nand U9057 (N_9057,N_6651,N_6844);
and U9058 (N_9058,N_7384,N_8582);
or U9059 (N_9059,N_6230,N_6824);
or U9060 (N_9060,N_8701,N_6056);
nor U9061 (N_9061,N_7049,N_6055);
nor U9062 (N_9062,N_6630,N_7541);
nor U9063 (N_9063,N_6009,N_7809);
nor U9064 (N_9064,N_6976,N_6957);
nand U9065 (N_9065,N_6027,N_6963);
nor U9066 (N_9066,N_8324,N_8752);
xnor U9067 (N_9067,N_7735,N_6306);
nand U9068 (N_9068,N_6408,N_8696);
xnor U9069 (N_9069,N_7235,N_8824);
and U9070 (N_9070,N_6671,N_7152);
and U9071 (N_9071,N_8799,N_8236);
nor U9072 (N_9072,N_7803,N_7122);
and U9073 (N_9073,N_8750,N_8899);
xor U9074 (N_9074,N_8737,N_8743);
xnor U9075 (N_9075,N_7934,N_7835);
nand U9076 (N_9076,N_7350,N_6289);
nor U9077 (N_9077,N_6387,N_8961);
xor U9078 (N_9078,N_6081,N_7303);
nand U9079 (N_9079,N_6667,N_7226);
nor U9080 (N_9080,N_7000,N_6109);
and U9081 (N_9081,N_7425,N_6359);
nor U9082 (N_9082,N_6747,N_7632);
and U9083 (N_9083,N_8307,N_6602);
nor U9084 (N_9084,N_8305,N_6601);
nand U9085 (N_9085,N_8727,N_7232);
or U9086 (N_9086,N_8523,N_8091);
xor U9087 (N_9087,N_8816,N_7896);
xnor U9088 (N_9088,N_8249,N_7679);
nor U9089 (N_9089,N_6712,N_8553);
or U9090 (N_9090,N_8617,N_6607);
and U9091 (N_9091,N_6380,N_6717);
or U9092 (N_9092,N_7689,N_6744);
or U9093 (N_9093,N_8369,N_7954);
xnor U9094 (N_9094,N_8707,N_6617);
or U9095 (N_9095,N_6382,N_8822);
and U9096 (N_9096,N_6498,N_6924);
nor U9097 (N_9097,N_8492,N_6202);
and U9098 (N_9098,N_8043,N_7702);
and U9099 (N_9099,N_7734,N_6257);
xor U9100 (N_9100,N_7429,N_7006);
or U9101 (N_9101,N_8371,N_6150);
or U9102 (N_9102,N_6204,N_8848);
nor U9103 (N_9103,N_7505,N_8865);
xor U9104 (N_9104,N_8437,N_8003);
nor U9105 (N_9105,N_8744,N_7536);
or U9106 (N_9106,N_8855,N_8511);
and U9107 (N_9107,N_6518,N_7806);
nor U9108 (N_9108,N_7643,N_6142);
nand U9109 (N_9109,N_7642,N_8287);
nand U9110 (N_9110,N_6608,N_6448);
xnor U9111 (N_9111,N_7272,N_8378);
nor U9112 (N_9112,N_7515,N_8263);
or U9113 (N_9113,N_6887,N_6777);
xnor U9114 (N_9114,N_7867,N_6154);
nor U9115 (N_9115,N_8195,N_8475);
nand U9116 (N_9116,N_7568,N_7647);
nand U9117 (N_9117,N_6907,N_6329);
and U9118 (N_9118,N_8127,N_6214);
and U9119 (N_9119,N_7510,N_7354);
nand U9120 (N_9120,N_8712,N_8144);
nor U9121 (N_9121,N_6096,N_8558);
or U9122 (N_9122,N_8714,N_7840);
nand U9123 (N_9123,N_6156,N_8930);
and U9124 (N_9124,N_8254,N_8487);
and U9125 (N_9125,N_7489,N_7364);
or U9126 (N_9126,N_6889,N_6369);
or U9127 (N_9127,N_8856,N_7047);
and U9128 (N_9128,N_8757,N_7095);
nor U9129 (N_9129,N_7458,N_8370);
xor U9130 (N_9130,N_8578,N_7111);
and U9131 (N_9131,N_8271,N_6195);
nor U9132 (N_9132,N_6842,N_8622);
or U9133 (N_9133,N_7317,N_8648);
or U9134 (N_9134,N_6533,N_6241);
xor U9135 (N_9135,N_8657,N_8916);
or U9136 (N_9136,N_7795,N_6423);
nand U9137 (N_9137,N_8049,N_8465);
nand U9138 (N_9138,N_8039,N_8248);
nor U9139 (N_9139,N_7514,N_8864);
and U9140 (N_9140,N_7854,N_6102);
or U9141 (N_9141,N_7258,N_6571);
or U9142 (N_9142,N_6422,N_7129);
xnor U9143 (N_9143,N_8420,N_8684);
and U9144 (N_9144,N_7634,N_8600);
and U9145 (N_9145,N_8000,N_7842);
and U9146 (N_9146,N_6599,N_6762);
xor U9147 (N_9147,N_8801,N_7508);
nand U9148 (N_9148,N_6268,N_7929);
and U9149 (N_9149,N_7436,N_6012);
xor U9150 (N_9150,N_6934,N_6999);
or U9151 (N_9151,N_7951,N_7736);
nand U9152 (N_9152,N_8191,N_7378);
nand U9153 (N_9153,N_7748,N_7316);
nor U9154 (N_9154,N_8967,N_7447);
xnor U9155 (N_9155,N_7296,N_7542);
xnor U9156 (N_9156,N_7424,N_8229);
and U9157 (N_9157,N_8242,N_7752);
nand U9158 (N_9158,N_8745,N_6120);
or U9159 (N_9159,N_6255,N_7699);
nand U9160 (N_9160,N_8527,N_7940);
or U9161 (N_9161,N_6300,N_6531);
nor U9162 (N_9162,N_7361,N_6967);
xnor U9163 (N_9163,N_6079,N_7312);
and U9164 (N_9164,N_6028,N_7112);
nor U9165 (N_9165,N_8180,N_7494);
or U9166 (N_9166,N_6211,N_6185);
nand U9167 (N_9167,N_6988,N_8516);
nand U9168 (N_9168,N_8970,N_8497);
xnor U9169 (N_9169,N_6301,N_7266);
nor U9170 (N_9170,N_7673,N_7033);
or U9171 (N_9171,N_6458,N_8404);
nand U9172 (N_9172,N_6413,N_6926);
and U9173 (N_9173,N_8532,N_8213);
and U9174 (N_9174,N_7713,N_8048);
nor U9175 (N_9175,N_7847,N_7986);
or U9176 (N_9176,N_7259,N_6789);
or U9177 (N_9177,N_7547,N_7426);
or U9178 (N_9178,N_7063,N_7869);
xor U9179 (N_9179,N_7428,N_7930);
and U9180 (N_9180,N_7749,N_7089);
nand U9181 (N_9181,N_7766,N_8100);
nand U9182 (N_9182,N_7830,N_8055);
and U9183 (N_9183,N_7440,N_6856);
nand U9184 (N_9184,N_7725,N_6494);
and U9185 (N_9185,N_7837,N_7273);
and U9186 (N_9186,N_6295,N_8652);
nor U9187 (N_9187,N_7348,N_6828);
and U9188 (N_9188,N_6445,N_7926);
nor U9189 (N_9189,N_7765,N_6393);
or U9190 (N_9190,N_7516,N_8449);
and U9191 (N_9191,N_7786,N_6778);
and U9192 (N_9192,N_6863,N_8001);
nand U9193 (N_9193,N_7800,N_7621);
or U9194 (N_9194,N_8767,N_8047);
and U9195 (N_9195,N_7747,N_6949);
or U9196 (N_9196,N_6266,N_7292);
and U9197 (N_9197,N_8005,N_8624);
xnor U9198 (N_9198,N_8379,N_7641);
and U9199 (N_9199,N_7216,N_8786);
xor U9200 (N_9200,N_8211,N_7889);
and U9201 (N_9201,N_6435,N_8060);
nor U9202 (N_9202,N_6388,N_8289);
nor U9203 (N_9203,N_8891,N_8932);
and U9204 (N_9204,N_7903,N_7041);
nand U9205 (N_9205,N_8027,N_8823);
nand U9206 (N_9206,N_6430,N_8362);
or U9207 (N_9207,N_7802,N_6327);
and U9208 (N_9208,N_8247,N_8835);
and U9209 (N_9209,N_7654,N_7085);
and U9210 (N_9210,N_8356,N_6414);
xnor U9211 (N_9211,N_8674,N_6196);
nor U9212 (N_9212,N_7608,N_8159);
nor U9213 (N_9213,N_6094,N_7276);
nor U9214 (N_9214,N_8447,N_8610);
xor U9215 (N_9215,N_6584,N_6360);
nand U9216 (N_9216,N_8154,N_6921);
xnor U9217 (N_9217,N_6010,N_8124);
nand U9218 (N_9218,N_7556,N_7966);
and U9219 (N_9219,N_6901,N_8469);
xor U9220 (N_9220,N_7572,N_7864);
xnor U9221 (N_9221,N_6491,N_7297);
xor U9222 (N_9222,N_7318,N_6194);
nand U9223 (N_9223,N_8590,N_7177);
nor U9224 (N_9224,N_8851,N_6972);
or U9225 (N_9225,N_8235,N_6766);
or U9226 (N_9226,N_7512,N_6823);
and U9227 (N_9227,N_8679,N_6112);
xor U9228 (N_9228,N_8978,N_8011);
xor U9229 (N_9229,N_8253,N_6585);
xnor U9230 (N_9230,N_6383,N_7114);
or U9231 (N_9231,N_6818,N_8295);
and U9232 (N_9232,N_6349,N_7876);
or U9233 (N_9233,N_8323,N_6875);
nand U9234 (N_9234,N_8580,N_8708);
and U9235 (N_9235,N_8002,N_8813);
and U9236 (N_9236,N_7845,N_7970);
nand U9237 (N_9237,N_8547,N_7020);
and U9238 (N_9238,N_7154,N_6239);
xnor U9239 (N_9239,N_6184,N_8607);
nand U9240 (N_9240,N_7922,N_6544);
and U9241 (N_9241,N_7885,N_6455);
nor U9242 (N_9242,N_8741,N_7636);
or U9243 (N_9243,N_8833,N_6583);
xor U9244 (N_9244,N_8638,N_7157);
nor U9245 (N_9245,N_7454,N_7288);
xor U9246 (N_9246,N_6016,N_7200);
nand U9247 (N_9247,N_6070,N_7075);
nor U9248 (N_9248,N_8350,N_6704);
xnor U9249 (N_9249,N_8148,N_6089);
nor U9250 (N_9250,N_6222,N_8075);
and U9251 (N_9251,N_7956,N_7298);
or U9252 (N_9252,N_8203,N_7392);
xnor U9253 (N_9253,N_8418,N_7282);
or U9254 (N_9254,N_7849,N_7964);
nor U9255 (N_9255,N_8642,N_6501);
and U9256 (N_9256,N_8424,N_6718);
nand U9257 (N_9257,N_8141,N_8973);
xnor U9258 (N_9258,N_7186,N_6475);
or U9259 (N_9259,N_7141,N_6471);
xnor U9260 (N_9260,N_6172,N_8777);
and U9261 (N_9261,N_6786,N_7592);
or U9262 (N_9262,N_6740,N_6362);
nor U9263 (N_9263,N_7761,N_8680);
nand U9264 (N_9264,N_6956,N_8059);
xnor U9265 (N_9265,N_6946,N_6902);
or U9266 (N_9266,N_7594,N_8640);
or U9267 (N_9267,N_7180,N_6272);
xnor U9268 (N_9268,N_7832,N_7865);
xor U9269 (N_9269,N_7328,N_6293);
nor U9270 (N_9270,N_6345,N_6997);
or U9271 (N_9271,N_7045,N_6636);
nor U9272 (N_9272,N_8343,N_6451);
xnor U9273 (N_9273,N_8104,N_6140);
or U9274 (N_9274,N_6376,N_7070);
xnor U9275 (N_9275,N_8985,N_8083);
xnor U9276 (N_9276,N_8302,N_8935);
or U9277 (N_9277,N_6661,N_7637);
and U9278 (N_9278,N_6570,N_6427);
and U9279 (N_9279,N_6466,N_8053);
xor U9280 (N_9280,N_7919,N_7910);
nand U9281 (N_9281,N_7402,N_6419);
nor U9282 (N_9282,N_7196,N_7880);
xor U9283 (N_9283,N_7231,N_7058);
and U9284 (N_9284,N_8765,N_8056);
nand U9285 (N_9285,N_6253,N_8987);
nor U9286 (N_9286,N_7787,N_8837);
nand U9287 (N_9287,N_7714,N_8219);
and U9288 (N_9288,N_7758,N_6892);
or U9289 (N_9289,N_8206,N_8603);
nor U9290 (N_9290,N_8883,N_6912);
and U9291 (N_9291,N_7548,N_8790);
xnor U9292 (N_9292,N_7341,N_7579);
and U9293 (N_9293,N_6611,N_6839);
or U9294 (N_9294,N_6868,N_7182);
nand U9295 (N_9295,N_8337,N_6219);
nand U9296 (N_9296,N_6994,N_6078);
nand U9297 (N_9297,N_6951,N_7135);
or U9298 (N_9298,N_7413,N_8114);
and U9299 (N_9299,N_7976,N_7819);
or U9300 (N_9300,N_7340,N_6311);
nand U9301 (N_9301,N_6303,N_8115);
xor U9302 (N_9302,N_8029,N_6898);
and U9303 (N_9303,N_6054,N_8692);
or U9304 (N_9304,N_7385,N_6524);
nand U9305 (N_9305,N_7895,N_6952);
and U9306 (N_9306,N_8836,N_7343);
nand U9307 (N_9307,N_7882,N_7473);
or U9308 (N_9308,N_8421,N_8291);
nand U9309 (N_9309,N_8804,N_8064);
or U9310 (N_9310,N_7016,N_6159);
or U9311 (N_9311,N_6637,N_8861);
and U9312 (N_9312,N_8258,N_6291);
nand U9313 (N_9313,N_6625,N_6274);
nor U9314 (N_9314,N_6929,N_6342);
nor U9315 (N_9315,N_8699,N_8294);
xnor U9316 (N_9316,N_6198,N_8441);
nand U9317 (N_9317,N_6790,N_7031);
nor U9318 (N_9318,N_8746,N_8564);
xor U9319 (N_9319,N_7060,N_6011);
xnor U9320 (N_9320,N_6605,N_8858);
and U9321 (N_9321,N_8901,N_7339);
xnor U9322 (N_9322,N_8502,N_6572);
nor U9323 (N_9323,N_8332,N_7081);
nor U9324 (N_9324,N_6795,N_6125);
and U9325 (N_9325,N_8283,N_8522);
xnor U9326 (N_9326,N_6805,N_7815);
nor U9327 (N_9327,N_8041,N_8782);
and U9328 (N_9328,N_8175,N_8890);
xor U9329 (N_9329,N_8647,N_7238);
xor U9330 (N_9330,N_6550,N_6647);
or U9331 (N_9331,N_7941,N_6650);
xor U9332 (N_9332,N_7859,N_6288);
xnor U9333 (N_9333,N_7433,N_6192);
and U9334 (N_9334,N_8538,N_6064);
xnor U9335 (N_9335,N_8192,N_6385);
or U9336 (N_9336,N_7086,N_7295);
nand U9337 (N_9337,N_7323,N_7390);
nand U9338 (N_9338,N_8923,N_7255);
nor U9339 (N_9339,N_6394,N_6203);
and U9340 (N_9340,N_6631,N_7301);
nand U9341 (N_9341,N_6294,N_6048);
and U9342 (N_9342,N_6779,N_8251);
or U9343 (N_9343,N_8595,N_6804);
nand U9344 (N_9344,N_6940,N_6310);
nor U9345 (N_9345,N_7038,N_7018);
or U9346 (N_9346,N_8798,N_6725);
nand U9347 (N_9347,N_6793,N_6258);
or U9348 (N_9348,N_7486,N_6250);
nor U9349 (N_9349,N_8090,N_6846);
nand U9350 (N_9350,N_7423,N_7683);
or U9351 (N_9351,N_7836,N_8887);
nor U9352 (N_9352,N_7708,N_8694);
nor U9353 (N_9353,N_7496,N_7136);
nor U9354 (N_9354,N_7243,N_7500);
or U9355 (N_9355,N_8493,N_7582);
xor U9356 (N_9356,N_6044,N_7932);
or U9357 (N_9357,N_8228,N_6206);
and U9358 (N_9358,N_6093,N_7746);
xnor U9359 (N_9359,N_8396,N_7978);
nor U9360 (N_9360,N_6254,N_6076);
nor U9361 (N_9361,N_7219,N_7788);
xor U9362 (N_9362,N_7814,N_8215);
xor U9363 (N_9363,N_6568,N_8417);
and U9364 (N_9364,N_8281,N_6259);
nand U9365 (N_9365,N_6654,N_7529);
xnor U9366 (N_9366,N_7899,N_7291);
and U9367 (N_9367,N_8473,N_6233);
and U9368 (N_9368,N_6987,N_6453);
and U9369 (N_9369,N_6030,N_6621);
xor U9370 (N_9370,N_8136,N_7630);
nor U9371 (N_9371,N_7872,N_6316);
nand U9372 (N_9372,N_7957,N_6304);
nand U9373 (N_9373,N_8474,N_7228);
nor U9374 (N_9374,N_8943,N_6928);
xnor U9375 (N_9375,N_6886,N_8036);
xor U9376 (N_9376,N_7150,N_7530);
or U9377 (N_9377,N_8984,N_6791);
and U9378 (N_9378,N_7427,N_7550);
nand U9379 (N_9379,N_8410,N_7771);
and U9380 (N_9380,N_7274,N_8894);
and U9381 (N_9381,N_8586,N_6908);
nand U9382 (N_9382,N_7503,N_6539);
nand U9383 (N_9383,N_8808,N_7731);
xor U9384 (N_9384,N_6622,N_7333);
xor U9385 (N_9385,N_8483,N_7712);
nand U9386 (N_9386,N_6454,N_8499);
or U9387 (N_9387,N_7064,N_7344);
nand U9388 (N_9388,N_8700,N_8884);
nand U9389 (N_9389,N_7422,N_7199);
or U9390 (N_9390,N_7088,N_6827);
nand U9391 (N_9391,N_6026,N_8664);
xor U9392 (N_9392,N_8810,N_6105);
nor U9393 (N_9393,N_7399,N_6439);
nor U9394 (N_9394,N_8314,N_8140);
nand U9395 (N_9395,N_8014,N_7798);
nand U9396 (N_9396,N_6769,N_6520);
nor U9397 (N_9397,N_6399,N_8122);
nor U9398 (N_9398,N_8990,N_6344);
xnor U9399 (N_9399,N_6982,N_6017);
xnor U9400 (N_9400,N_8071,N_7993);
or U9401 (N_9401,N_8150,N_8724);
or U9402 (N_9402,N_8065,N_7332);
and U9403 (N_9403,N_8852,N_7879);
and U9404 (N_9404,N_8086,N_7353);
xor U9405 (N_9405,N_7294,N_7096);
xnor U9406 (N_9406,N_8019,N_8769);
or U9407 (N_9407,N_7195,N_6396);
and U9408 (N_9408,N_6756,N_7523);
nand U9409 (N_9409,N_7946,N_6700);
or U9410 (N_9410,N_6136,N_6496);
or U9411 (N_9411,N_6124,N_8004);
nand U9412 (N_9412,N_7831,N_7797);
nor U9413 (N_9413,N_6472,N_8885);
or U9414 (N_9414,N_8467,N_6465);
nand U9415 (N_9415,N_7140,N_7604);
or U9416 (N_9416,N_7552,N_6504);
xnor U9417 (N_9417,N_6042,N_6603);
xnor U9418 (N_9418,N_7054,N_8625);
or U9419 (N_9419,N_8905,N_7314);
nor U9420 (N_9420,N_8366,N_7662);
nor U9421 (N_9421,N_6226,N_7227);
or U9422 (N_9422,N_7275,N_6041);
nand U9423 (N_9423,N_8246,N_8376);
or U9424 (N_9424,N_6216,N_8162);
and U9425 (N_9425,N_8933,N_8035);
nand U9426 (N_9426,N_6169,N_8385);
or U9427 (N_9427,N_8119,N_6151);
and U9428 (N_9428,N_6593,N_7420);
nand U9429 (N_9429,N_8549,N_6270);
nand U9430 (N_9430,N_7789,N_8874);
nor U9431 (N_9431,N_7942,N_6881);
xnor U9432 (N_9432,N_6002,N_6275);
and U9433 (N_9433,N_7445,N_8335);
or U9434 (N_9434,N_7696,N_6559);
xnor U9435 (N_9435,N_7709,N_6586);
nand U9436 (N_9436,N_6177,N_7935);
xnor U9437 (N_9437,N_8020,N_8878);
nor U9438 (N_9438,N_7464,N_7822);
nor U9439 (N_9439,N_7452,N_7796);
nor U9440 (N_9440,N_7076,N_7569);
or U9441 (N_9441,N_8755,N_8530);
nand U9442 (N_9442,N_8193,N_7753);
nor U9443 (N_9443,N_7206,N_7271);
xor U9444 (N_9444,N_8189,N_8685);
nand U9445 (N_9445,N_6476,N_6407);
nor U9446 (N_9446,N_6090,N_7495);
xnor U9447 (N_9447,N_7260,N_8304);
nand U9448 (N_9448,N_7061,N_6083);
and U9449 (N_9449,N_8108,N_7640);
nor U9450 (N_9450,N_8649,N_6375);
or U9451 (N_9451,N_8194,N_7825);
and U9452 (N_9452,N_7212,N_7967);
nand U9453 (N_9453,N_7600,N_7442);
or U9454 (N_9454,N_8120,N_8186);
or U9455 (N_9455,N_6745,N_7980);
and U9456 (N_9456,N_7717,N_6225);
nand U9457 (N_9457,N_8422,N_7706);
xor U9458 (N_9458,N_6681,N_6911);
and U9459 (N_9459,N_7931,N_7381);
xnor U9460 (N_9460,N_8871,N_8466);
or U9461 (N_9461,N_6950,N_7262);
nor U9462 (N_9462,N_6995,N_6662);
xor U9463 (N_9463,N_7287,N_6244);
or U9464 (N_9464,N_7048,N_7370);
xnor U9465 (N_9465,N_7912,N_7205);
or U9466 (N_9466,N_8570,N_7193);
and U9467 (N_9467,N_6983,N_6428);
or U9468 (N_9468,N_7599,N_8412);
xor U9469 (N_9469,N_8960,N_7633);
and U9470 (N_9470,N_6264,N_6733);
nand U9471 (N_9471,N_7393,N_7403);
or U9472 (N_9472,N_7624,N_7408);
xor U9473 (N_9473,N_7011,N_7818);
nand U9474 (N_9474,N_7389,N_6449);
and U9475 (N_9475,N_8089,N_8407);
nor U9476 (N_9476,N_6227,N_6488);
or U9477 (N_9477,N_8695,N_7590);
xnor U9478 (N_9478,N_8130,N_6245);
xnor U9479 (N_9479,N_6734,N_8037);
or U9480 (N_9480,N_7234,N_6566);
or U9481 (N_9481,N_7457,N_6758);
or U9482 (N_9482,N_7520,N_6900);
nor U9483 (N_9483,N_6841,N_7337);
or U9484 (N_9484,N_8662,N_8443);
nand U9485 (N_9485,N_7664,N_6200);
or U9486 (N_9486,N_8999,N_7742);
or U9487 (N_9487,N_7862,N_6635);
and U9488 (N_9488,N_6354,N_8456);
xnor U9489 (N_9489,N_6271,N_6395);
xnor U9490 (N_9490,N_8952,N_7077);
and U9491 (N_9491,N_7278,N_8028);
and U9492 (N_9492,N_7511,N_6925);
and U9493 (N_9493,N_7625,N_7578);
nand U9494 (N_9494,N_7091,N_8317);
or U9495 (N_9495,N_7943,N_6098);
nor U9496 (N_9496,N_7261,N_7628);
or U9497 (N_9497,N_8903,N_8983);
or U9498 (N_9498,N_8044,N_8859);
and U9499 (N_9499,N_7451,N_6087);
xor U9500 (N_9500,N_8448,N_8311);
or U9501 (N_9501,N_6708,N_6147);
and U9502 (N_9502,N_8063,N_7277);
xor U9503 (N_9503,N_8391,N_7502);
xnor U9504 (N_9504,N_6859,N_7462);
or U9505 (N_9505,N_8872,N_7558);
xor U9506 (N_9506,N_7358,N_8346);
or U9507 (N_9507,N_6187,N_6594);
nor U9508 (N_9508,N_8135,N_6173);
and U9509 (N_9509,N_7877,N_7720);
xnor U9510 (N_9510,N_6050,N_7581);
xnor U9511 (N_9511,N_7913,N_8980);
nor U9512 (N_9512,N_8430,N_7770);
and U9513 (N_9513,N_7249,N_6317);
or U9514 (N_9514,N_7554,N_6975);
xor U9515 (N_9515,N_6181,N_8085);
nor U9516 (N_9516,N_7911,N_8626);
nand U9517 (N_9517,N_7069,N_6265);
xnor U9518 (N_9518,N_6378,N_8628);
nor U9519 (N_9519,N_8515,N_7546);
xnor U9520 (N_9520,N_8481,N_8128);
nand U9521 (N_9521,N_6318,N_7705);
nor U9522 (N_9522,N_8879,N_6052);
nand U9523 (N_9523,N_8536,N_6980);
and U9524 (N_9524,N_7053,N_6961);
xor U9525 (N_9525,N_6057,N_8659);
xor U9526 (N_9526,N_8653,N_7841);
or U9527 (N_9527,N_8948,N_6469);
nor U9528 (N_9528,N_6699,N_7133);
nand U9529 (N_9529,N_7593,N_6687);
nand U9530 (N_9530,N_7165,N_8658);
nand U9531 (N_9531,N_7302,N_6138);
nor U9532 (N_9532,N_6598,N_8429);
or U9533 (N_9533,N_8264,N_7855);
nor U9534 (N_9534,N_7431,N_7214);
or U9535 (N_9535,N_6364,N_8177);
or U9536 (N_9536,N_7540,N_6843);
and U9537 (N_9537,N_6024,N_7694);
and U9538 (N_9538,N_6073,N_8187);
or U9539 (N_9539,N_6854,N_6459);
or U9540 (N_9540,N_8524,N_6486);
nor U9541 (N_9541,N_7887,N_8454);
nand U9542 (N_9542,N_8514,N_7118);
nand U9543 (N_9543,N_8926,N_7844);
nand U9544 (N_9544,N_8419,N_7767);
nand U9545 (N_9545,N_8157,N_6545);
and U9546 (N_9546,N_8214,N_6965);
or U9547 (N_9547,N_8636,N_6979);
nor U9548 (N_9548,N_7577,N_8330);
nand U9549 (N_9549,N_7019,N_7857);
and U9550 (N_9550,N_7338,N_8543);
nand U9551 (N_9551,N_7521,N_7359);
xor U9552 (N_9552,N_8170,N_7101);
xor U9553 (N_9553,N_7345,N_6450);
or U9554 (N_9554,N_7588,N_6556);
xnor U9555 (N_9555,N_6106,N_6861);
or U9556 (N_9556,N_8276,N_6003);
nand U9557 (N_9557,N_8612,N_6197);
nor U9558 (N_9558,N_8078,N_8797);
and U9559 (N_9559,N_8273,N_8959);
nand U9560 (N_9560,N_8839,N_8102);
or U9561 (N_9561,N_6474,N_6082);
or U9562 (N_9562,N_6515,N_8779);
nand U9563 (N_9563,N_7997,N_7382);
nand U9564 (N_9564,N_7925,N_7952);
or U9565 (N_9565,N_7597,N_7242);
nand U9566 (N_9566,N_6401,N_8734);
nor U9567 (N_9567,N_7607,N_8809);
nor U9568 (N_9568,N_7678,N_6348);
and U9569 (N_9569,N_8269,N_7890);
xor U9570 (N_9570,N_7080,N_6484);
nand U9571 (N_9571,N_8849,N_7892);
nand U9572 (N_9572,N_7470,N_7490);
nor U9573 (N_9573,N_8439,N_7914);
and U9574 (N_9574,N_6962,N_8921);
nand U9575 (N_9575,N_8435,N_7388);
and U9576 (N_9576,N_7349,N_6020);
and U9577 (N_9577,N_8220,N_7146);
xnor U9578 (N_9578,N_8197,N_7656);
nand U9579 (N_9579,N_7466,N_6467);
nor U9580 (N_9580,N_6909,N_8537);
nand U9581 (N_9581,N_6890,N_8829);
and U9582 (N_9582,N_8842,N_8359);
nor U9583 (N_9583,N_7998,N_6405);
nand U9584 (N_9584,N_7991,N_8199);
xnor U9585 (N_9585,N_8444,N_8597);
nor U9586 (N_9586,N_7769,N_6537);
and U9587 (N_9587,N_6217,N_6797);
or U9588 (N_9588,N_8678,N_7253);
or U9589 (N_9589,N_8325,N_8641);
nand U9590 (N_9590,N_8613,N_7387);
xnor U9591 (N_9591,N_7900,N_6153);
xor U9592 (N_9592,N_6981,N_7573);
xor U9593 (N_9593,N_7959,N_6481);
nor U9594 (N_9594,N_8318,N_6960);
or U9595 (N_9595,N_6640,N_7410);
or U9596 (N_9596,N_6452,N_8225);
or U9597 (N_9597,N_6416,N_7740);
nor U9598 (N_9598,N_8277,N_7023);
xnor U9599 (N_9599,N_8218,N_6074);
nand U9600 (N_9600,N_8900,N_7777);
xnor U9601 (N_9601,N_6510,N_7838);
xnor U9602 (N_9602,N_6903,N_6328);
nand U9603 (N_9603,N_8468,N_7404);
and U9604 (N_9604,N_6563,N_8929);
xnor U9605 (N_9605,N_8726,N_8761);
and U9606 (N_9606,N_6267,N_8986);
and U9607 (N_9607,N_6668,N_7194);
xnor U9608 (N_9608,N_7644,N_6256);
or U9609 (N_9609,N_6308,N_8103);
or U9610 (N_9610,N_7775,N_7179);
xor U9611 (N_9611,N_6330,N_7124);
and U9612 (N_9612,N_8946,N_8898);
xnor U9613 (N_9613,N_7620,N_6785);
or U9614 (N_9614,N_8736,N_6977);
xor U9615 (N_9615,N_6193,N_7866);
or U9616 (N_9616,N_8426,N_6281);
and U9617 (N_9617,N_6726,N_6592);
or U9618 (N_9618,N_6224,N_8517);
nand U9619 (N_9619,N_6672,N_6292);
or U9620 (N_9620,N_7151,N_7863);
and U9621 (N_9621,N_6871,N_6632);
nor U9622 (N_9622,N_7860,N_6006);
nand U9623 (N_9623,N_6324,N_7610);
or U9624 (N_9624,N_7534,N_8205);
nor U9625 (N_9625,N_7237,N_8563);
nor U9626 (N_9626,N_8531,N_6867);
xnor U9627 (N_9627,N_6806,N_8132);
xor U9628 (N_9628,N_7421,N_7396);
or U9629 (N_9629,N_7651,N_8955);
and U9630 (N_9630,N_7477,N_7627);
and U9631 (N_9631,N_8482,N_6534);
nor U9632 (N_9632,N_8630,N_8344);
and U9633 (N_9633,N_6812,N_6551);
and U9634 (N_9634,N_7022,N_6670);
or U9635 (N_9635,N_7589,N_6335);
nand U9636 (N_9636,N_7040,N_8644);
and U9637 (N_9637,N_7071,N_6337);
xor U9638 (N_9638,N_6088,N_7208);
xnor U9639 (N_9639,N_6280,N_8181);
nand U9640 (N_9640,N_8796,N_7439);
and U9641 (N_9641,N_6526,N_7975);
or U9642 (N_9642,N_6512,N_6884);
nand U9643 (N_9643,N_6996,N_6511);
xor U9644 (N_9644,N_7667,N_7960);
xnor U9645 (N_9645,N_8908,N_8738);
xor U9646 (N_9646,N_6508,N_7504);
xor U9647 (N_9647,N_7638,N_7072);
nor U9648 (N_9648,N_8245,N_6894);
and U9649 (N_9649,N_8886,N_7355);
nand U9650 (N_9650,N_7861,N_8691);
or U9651 (N_9651,N_8024,N_6163);
nor U9652 (N_9652,N_7733,N_6992);
or U9653 (N_9653,N_7263,N_6590);
nand U9654 (N_9654,N_7025,N_6803);
and U9655 (N_9655,N_7741,N_7517);
xor U9656 (N_9656,N_7368,N_7304);
or U9657 (N_9657,N_6155,N_8576);
nand U9658 (N_9658,N_6855,N_7106);
xor U9659 (N_9659,N_8751,N_6792);
nor U9660 (N_9660,N_8166,N_6927);
and U9661 (N_9661,N_8408,N_8331);
xor U9662 (N_9662,N_8771,N_6836);
nand U9663 (N_9663,N_8529,N_8749);
and U9664 (N_9664,N_7012,N_6305);
and U9665 (N_9665,N_8403,N_6249);
and U9666 (N_9666,N_8096,N_6693);
or U9667 (N_9667,N_8730,N_7616);
nand U9668 (N_9668,N_6130,N_6015);
and U9669 (N_9669,N_6236,N_6312);
nor U9670 (N_9670,N_8974,N_8768);
and U9671 (N_9671,N_6953,N_6893);
nand U9672 (N_9672,N_6208,N_8095);
xor U9673 (N_9673,N_6609,N_8334);
nor U9674 (N_9674,N_7584,N_6974);
and U9675 (N_9675,N_7528,N_7026);
and U9676 (N_9676,N_7245,N_7042);
nor U9677 (N_9677,N_8094,N_8794);
xnor U9678 (N_9678,N_8689,N_6493);
and U9679 (N_9679,N_7472,N_6221);
nor U9680 (N_9680,N_8676,N_8081);
or U9681 (N_9681,N_8116,N_6763);
xor U9682 (N_9682,N_6477,N_7149);
nand U9683 (N_9683,N_7677,N_8840);
nand U9684 (N_9684,N_6536,N_6959);
nor U9685 (N_9685,N_6008,N_8485);
and U9686 (N_9686,N_7779,N_7108);
and U9687 (N_9687,N_6059,N_6589);
xnor U9688 (N_9688,N_6800,N_8042);
xnor U9689 (N_9689,N_6495,N_8315);
and U9690 (N_9690,N_7051,N_6817);
and U9691 (N_9691,N_7805,N_7973);
and U9692 (N_9692,N_7598,N_7813);
and U9693 (N_9693,N_6528,N_6558);
and U9694 (N_9694,N_8423,N_7221);
and U9695 (N_9695,N_7917,N_6220);
and U9696 (N_9696,N_6897,N_6352);
and U9697 (N_9697,N_8284,N_6092);
xor U9698 (N_9698,N_8282,N_7225);
and U9699 (N_9699,N_7014,N_8778);
and U9700 (N_9700,N_6379,N_7563);
nand U9701 (N_9701,N_7246,N_7468);
xor U9702 (N_9702,N_6004,N_8598);
xor U9703 (N_9703,N_8462,N_6860);
nor U9704 (N_9704,N_6366,N_6132);
nand U9705 (N_9705,N_6829,N_6606);
nand U9706 (N_9706,N_8950,N_8562);
nand U9707 (N_9707,N_6424,N_8131);
and U9708 (N_9708,N_8239,N_6418);
nor U9709 (N_9709,N_7961,N_6851);
nor U9710 (N_9710,N_7603,N_7475);
nand U9711 (N_9711,N_8588,N_7366);
nor U9712 (N_9712,N_6135,N_7904);
xor U9713 (N_9713,N_8888,N_8087);
and U9714 (N_9714,N_8262,N_7092);
nand U9715 (N_9715,N_6845,N_6989);
xor U9716 (N_9716,N_8329,N_6034);
nor U9717 (N_9717,N_6229,N_7596);
or U9718 (N_9718,N_7591,N_6916);
and U9719 (N_9719,N_6546,N_6355);
or U9720 (N_9720,N_6935,N_7418);
or U9721 (N_9721,N_6904,N_6040);
and U9722 (N_9722,N_7223,N_6331);
and U9723 (N_9723,N_7794,N_6497);
nand U9724 (N_9724,N_6358,N_7990);
xor U9725 (N_9725,N_7538,N_6037);
xor U9726 (N_9726,N_8068,N_7251);
xnor U9727 (N_9727,N_7927,N_6513);
nor U9728 (N_9728,N_8748,N_8428);
or U9729 (N_9729,N_8756,N_7972);
and U9730 (N_9730,N_7315,N_6788);
and U9731 (N_9731,N_6444,N_7097);
and U9732 (N_9732,N_7921,N_8587);
nand U9733 (N_9733,N_8208,N_7126);
nor U9734 (N_9734,N_8919,N_7132);
nor U9735 (N_9735,N_6021,N_6343);
and U9736 (N_9736,N_7102,N_8179);
or U9737 (N_9737,N_6463,N_7873);
nor U9738 (N_9738,N_6822,N_7988);
and U9739 (N_9739,N_7982,N_8693);
and U9740 (N_9740,N_6666,N_8683);
nand U9741 (N_9741,N_8139,N_7826);
xor U9742 (N_9742,N_6085,N_6732);
nor U9743 (N_9743,N_6062,N_8240);
nor U9744 (N_9744,N_7460,N_7005);
and U9745 (N_9745,N_6703,N_7479);
xnor U9746 (N_9746,N_6205,N_7650);
and U9747 (N_9747,N_6122,N_7675);
xor U9748 (N_9748,N_6525,N_6547);
or U9749 (N_9749,N_7169,N_8398);
nand U9750 (N_9750,N_7992,N_8012);
xor U9751 (N_9751,N_7331,N_7918);
nand U9752 (N_9752,N_7897,N_8544);
xnor U9753 (N_9753,N_8204,N_8328);
or U9754 (N_9754,N_8605,N_8066);
nor U9755 (N_9755,N_8023,N_8280);
or U9756 (N_9756,N_6429,N_7583);
nand U9757 (N_9757,N_8964,N_7307);
nand U9758 (N_9758,N_7113,N_6071);
nand U9759 (N_9759,N_7834,N_6910);
or U9760 (N_9760,N_6223,N_6646);
nand U9761 (N_9761,N_7760,N_7405);
nor U9762 (N_9762,N_8237,N_7028);
and U9763 (N_9763,N_8052,N_6391);
nand U9764 (N_9764,N_7004,N_7670);
and U9765 (N_9765,N_7724,N_8666);
and U9766 (N_9766,N_8399,N_6677);
and U9767 (N_9767,N_7909,N_7509);
and U9768 (N_9768,N_8844,N_7432);
nor U9769 (N_9769,N_8080,N_7719);
and U9770 (N_9770,N_6434,N_8963);
nand U9771 (N_9771,N_7833,N_7728);
nor U9772 (N_9772,N_7888,N_8133);
xnor U9773 (N_9773,N_6658,N_6619);
nand U9774 (N_9774,N_6319,N_7373);
or U9775 (N_9775,N_8875,N_8413);
or U9776 (N_9776,N_7293,N_8575);
and U9777 (N_9777,N_8355,N_8690);
or U9778 (N_9778,N_6938,N_6392);
or U9779 (N_9779,N_7409,N_7166);
xor U9780 (N_9780,N_6019,N_8484);
nand U9781 (N_9781,N_6047,N_7631);
nor U9782 (N_9782,N_8893,N_8728);
xor U9783 (N_9783,N_7184,N_7374);
xnor U9784 (N_9784,N_7394,N_8300);
nand U9785 (N_9785,N_7711,N_7974);
nand U9786 (N_9786,N_7730,N_7827);
xor U9787 (N_9787,N_7562,N_8533);
xor U9788 (N_9788,N_6038,N_8566);
xor U9789 (N_9789,N_6532,N_7414);
xnor U9790 (N_9790,N_8062,N_7491);
or U9791 (N_9791,N_8106,N_7958);
nand U9792 (N_9792,N_6492,N_6914);
xnor U9793 (N_9793,N_6891,N_6489);
nor U9794 (N_9794,N_8846,N_6698);
and U9795 (N_9795,N_7560,N_7419);
nand U9796 (N_9796,N_8158,N_6752);
nand U9797 (N_9797,N_7371,N_8814);
nand U9798 (N_9798,N_8336,N_7125);
nand U9799 (N_9799,N_7367,N_6410);
xor U9800 (N_9800,N_8671,N_6273);
xor U9801 (N_9801,N_8807,N_6696);
xor U9802 (N_9802,N_7778,N_6754);
and U9803 (N_9803,N_7984,N_7175);
or U9804 (N_9804,N_8572,N_6751);
nand U9805 (N_9805,N_8850,N_6032);
nor U9806 (N_9806,N_7372,N_8184);
xnor U9807 (N_9807,N_7220,N_7551);
xor U9808 (N_9808,N_8257,N_8098);
xnor U9809 (N_9809,N_8631,N_7127);
and U9810 (N_9810,N_8989,N_7804);
or U9811 (N_9811,N_6013,N_8160);
nand U9812 (N_9812,N_7799,N_8285);
xnor U9813 (N_9813,N_6523,N_6199);
nor U9814 (N_9814,N_6748,N_6134);
nor U9815 (N_9815,N_6674,N_6660);
and U9816 (N_9816,N_8224,N_8754);
nor U9817 (N_9817,N_7537,N_7290);
or U9818 (N_9818,N_8137,N_7281);
nand U9819 (N_9819,N_6314,N_8508);
nand U9820 (N_9820,N_6237,N_7784);
nand U9821 (N_9821,N_7557,N_7672);
or U9822 (N_9822,N_6749,N_8142);
or U9823 (N_9823,N_8256,N_7883);
xor U9824 (N_9824,N_6286,N_8445);
or U9825 (N_9825,N_6262,N_6260);
nor U9826 (N_9826,N_8913,N_7082);
nand U9827 (N_9827,N_8207,N_6833);
xor U9828 (N_9828,N_7626,N_8363);
and U9829 (N_9829,N_8512,N_8032);
xnor U9830 (N_9830,N_7104,N_7612);
xnor U9831 (N_9831,N_8780,N_8845);
xor U9832 (N_9832,N_8722,N_8968);
nor U9833 (N_9833,N_8167,N_7003);
or U9834 (N_9834,N_6587,N_8821);
nand U9835 (N_9835,N_6865,N_8975);
or U9836 (N_9836,N_6007,N_8753);
nand U9837 (N_9837,N_8288,N_7893);
nand U9838 (N_9838,N_8773,N_6022);
nor U9839 (N_9839,N_6460,N_6397);
nand U9840 (N_9840,N_7093,N_8993);
xor U9841 (N_9841,N_6582,N_8389);
and U9842 (N_9842,N_8489,N_8742);
xor U9843 (N_9843,N_8494,N_8397);
and U9844 (N_9844,N_6564,N_8581);
nand U9845 (N_9845,N_8503,N_6772);
xnor U9846 (N_9846,N_7660,N_6575);
or U9847 (N_9847,N_7655,N_8076);
xnor U9848 (N_9848,N_6971,N_6014);
nand U9849 (N_9849,N_8480,N_7224);
or U9850 (N_9850,N_7250,N_8279);
xnor U9851 (N_9851,N_6189,N_8414);
and U9852 (N_9852,N_7722,N_7908);
nand U9853 (N_9853,N_8675,N_7055);
nand U9854 (N_9854,N_7481,N_8268);
and U9855 (N_9855,N_6171,N_6578);
or U9856 (N_9856,N_8021,N_7191);
nand U9857 (N_9857,N_7383,N_6560);
nand U9858 (N_9858,N_7078,N_7902);
xor U9859 (N_9859,N_6905,N_7174);
xor U9860 (N_9860,N_8278,N_6796);
and U9861 (N_9861,N_7870,N_6179);
and U9862 (N_9862,N_6906,N_6645);
or U9863 (N_9863,N_6277,N_8009);
xor U9864 (N_9864,N_7068,N_8682);
or U9865 (N_9865,N_8713,N_7617);
nor U9866 (N_9866,N_8112,N_6885);
xnor U9867 (N_9867,N_8897,N_7635);
xnor U9868 (N_9868,N_7213,N_7605);
or U9869 (N_9869,N_8367,N_8555);
nand U9870 (N_9870,N_7233,N_8509);
or U9871 (N_9871,N_8994,N_8358);
nor U9872 (N_9872,N_8446,N_6107);
nand U9873 (N_9873,N_8107,N_6954);
and U9874 (N_9874,N_7718,N_7639);
nand U9875 (N_9875,N_8541,N_7032);
or U9876 (N_9876,N_7692,N_6097);
nand U9877 (N_9877,N_6299,N_6768);
or U9878 (N_9878,N_8817,N_7347);
or U9879 (N_9879,N_7280,N_8941);
nand U9880 (N_9880,N_6690,N_6655);
or U9881 (N_9881,N_8010,N_6509);
or U9882 (N_9882,N_8013,N_7401);
nand U9883 (N_9883,N_8997,N_6326);
or U9884 (N_9884,N_8016,N_8956);
or U9885 (N_9885,N_8645,N_8386);
and U9886 (N_9886,N_7821,N_7416);
nor U9887 (N_9887,N_8633,N_7211);
nor U9888 (N_9888,N_7485,N_7652);
nand U9889 (N_9889,N_8951,N_8301);
nand U9890 (N_9890,N_6577,N_7782);
and U9891 (N_9891,N_8433,N_6462);
or U9892 (N_9892,N_7207,N_7172);
and U9893 (N_9893,N_8099,N_7492);
nor U9894 (N_9894,N_7171,N_6128);
xor U9895 (N_9895,N_7543,N_6629);
or U9896 (N_9896,N_6191,N_8111);
nor U9897 (N_9897,N_6862,N_8395);
nor U9898 (N_9898,N_6679,N_6810);
nor U9899 (N_9899,N_8226,N_6065);
nor U9900 (N_9900,N_8971,N_7222);
or U9901 (N_9901,N_8711,N_8518);
and U9902 (N_9902,N_6158,N_6473);
or U9903 (N_9903,N_7823,N_6023);
xor U9904 (N_9904,N_7614,N_8787);
nor U9905 (N_9905,N_6931,N_6648);
nand U9906 (N_9906,N_7100,N_8793);
xor U9907 (N_9907,N_6641,N_8352);
nor U9908 (N_9908,N_6386,N_7571);
nor U9909 (N_9909,N_8486,N_8781);
nor U9910 (N_9910,N_8117,N_6058);
and U9911 (N_9911,N_7937,N_7131);
and U9912 (N_9912,N_8740,N_6573);
or U9913 (N_9913,N_8589,N_8155);
and U9914 (N_9914,N_8697,N_7886);
nor U9915 (N_9915,N_6659,N_6742);
xor U9916 (N_9916,N_8364,N_6175);
nor U9917 (N_9917,N_7322,N_7963);
and U9918 (N_9918,N_6882,N_8015);
or U9919 (N_9919,N_6320,N_8299);
xor U9920 (N_9920,N_7342,N_7907);
nand U9921 (N_9921,N_8008,N_8869);
nor U9922 (N_9922,N_8149,N_7891);
nor U9923 (N_9923,N_6433,N_6715);
or U9924 (N_9924,N_7501,N_7906);
nand U9925 (N_9925,N_7776,N_7197);
nor U9926 (N_9926,N_6919,N_7858);
or U9927 (N_9927,N_8702,N_6665);
xor U9928 (N_9928,N_7035,N_7449);
nor U9929 (N_9929,N_6984,N_6080);
xor U9930 (N_9930,N_6652,N_8962);
or U9931 (N_9931,N_8040,N_8673);
or U9932 (N_9932,N_8298,N_8552);
and U9933 (N_9933,N_8401,N_7356);
xor U9934 (N_9934,N_6247,N_6505);
nand U9935 (N_9935,N_7763,N_8910);
and U9936 (N_9936,N_7483,N_8290);
nand U9937 (N_9937,N_8272,N_8054);
nor U9938 (N_9938,N_8834,N_7757);
or U9939 (N_9939,N_6168,N_8938);
or U9940 (N_9940,N_6139,N_6176);
or U9941 (N_9941,N_8716,N_6049);
nor U9942 (N_9942,N_7665,N_8805);
nor U9943 (N_9943,N_8847,N_7532);
nand U9944 (N_9944,N_8451,N_8762);
xnor U9945 (N_9945,N_8405,N_8725);
nor U9946 (N_9946,N_8601,N_8873);
nand U9947 (N_9947,N_6000,N_6031);
nand U9948 (N_9948,N_7319,N_6743);
or U9949 (N_9949,N_8188,N_6709);
and U9950 (N_9950,N_6767,N_8618);
and U9951 (N_9951,N_6530,N_8594);
and U9952 (N_9952,N_7916,N_7324);
nand U9953 (N_9953,N_7311,N_6061);
nand U9954 (N_9954,N_7185,N_8365);
or U9955 (N_9955,N_8650,N_6985);
and U9956 (N_9956,N_6213,N_6947);
nor U9957 (N_9957,N_8450,N_8723);
or U9958 (N_9958,N_6799,N_6998);
nor U9959 (N_9959,N_6719,N_8459);
nor U9960 (N_9960,N_7601,N_8217);
xor U9961 (N_9961,N_7139,N_6421);
or U9962 (N_9962,N_8372,N_7284);
nor U9963 (N_9963,N_7363,N_8375);
nand U9964 (N_9964,N_6722,N_6826);
nor U9965 (N_9965,N_6933,N_8942);
xnor U9966 (N_9966,N_8567,N_6634);
xor U9967 (N_9967,N_6831,N_8792);
or U9968 (N_9968,N_8488,N_7875);
nand U9969 (N_9969,N_8088,N_8604);
nor U9970 (N_9970,N_7682,N_6285);
or U9971 (N_9971,N_7681,N_8109);
and U9972 (N_9972,N_7441,N_6479);
nor U9973 (N_9973,N_6595,N_6333);
xor U9974 (N_9974,N_8718,N_7116);
nor U9975 (N_9975,N_7817,N_8841);
nand U9976 (N_9976,N_6437,N_8457);
nand U9977 (N_9977,N_6600,N_8453);
or U9978 (N_9978,N_7933,N_7109);
xor U9979 (N_9979,N_7878,N_7727);
and U9980 (N_9980,N_7210,N_7120);
or U9981 (N_9981,N_6005,N_8791);
or U9982 (N_9982,N_8620,N_7217);
nand U9983 (N_9983,N_6870,N_6552);
and U9984 (N_9984,N_6261,N_6942);
and U9985 (N_9985,N_6440,N_6166);
or U9986 (N_9986,N_8686,N_8361);
xnor U9987 (N_9987,N_6403,N_8902);
and U9988 (N_9988,N_6798,N_8046);
nand U9989 (N_9989,N_8735,N_8267);
xor U9990 (N_9990,N_7456,N_7566);
nand U9991 (N_9991,N_8185,N_6527);
or U9992 (N_9992,N_8093,N_7979);
xnor U9993 (N_9993,N_6157,N_6899);
or U9994 (N_9994,N_7117,N_6626);
nor U9995 (N_9995,N_6069,N_6540);
xor U9996 (N_9996,N_8934,N_8812);
and U9997 (N_9997,N_6639,N_8917);
xor U9998 (N_9998,N_6170,N_6212);
or U9999 (N_9999,N_6436,N_8705);
or U10000 (N_10000,N_7999,N_8303);
xnor U10001 (N_10001,N_8381,N_7240);
nor U10002 (N_10002,N_6615,N_7335);
xnor U10003 (N_10003,N_8223,N_8635);
or U10004 (N_10004,N_8981,N_6442);
nand U10005 (N_10005,N_6516,N_8766);
or U10006 (N_10006,N_8319,N_6149);
and U10007 (N_10007,N_6468,N_6869);
xnor U10008 (N_10008,N_6251,N_8151);
xnor U10009 (N_10009,N_6263,N_7168);
nor U10010 (N_10010,N_8803,N_6108);
and U10011 (N_10011,N_7478,N_7905);
nor U10012 (N_10012,N_7687,N_6464);
nand U10013 (N_10013,N_6781,N_8828);
or U10014 (N_10014,N_8806,N_6809);
xnor U10015 (N_10015,N_8145,N_7187);
nand U10016 (N_10016,N_7507,N_7286);
xor U10017 (N_10017,N_7920,N_8914);
or U10018 (N_10018,N_8067,N_7484);
xnor U10019 (N_10019,N_7204,N_8925);
nand U10020 (N_10020,N_6642,N_6133);
nor U10021 (N_10021,N_6389,N_7066);
and U10022 (N_10022,N_7128,N_8763);
or U10023 (N_10023,N_6182,N_6773);
nor U10024 (N_10024,N_8360,N_7839);
xor U10025 (N_10025,N_7661,N_8472);
xnor U10026 (N_10026,N_6457,N_6143);
nor U10027 (N_10027,N_6321,N_6678);
nand U10028 (N_10028,N_7995,N_6104);
and U10029 (N_10029,N_6045,N_6018);
or U10030 (N_10030,N_8402,N_8202);
xor U10031 (N_10031,N_7241,N_7762);
xnor U10032 (N_10032,N_6764,N_7693);
xor U10033 (N_10033,N_8173,N_6067);
or U10034 (N_10034,N_7123,N_8862);
nand U10035 (N_10035,N_8668,N_6357);
nor U10036 (N_10036,N_7658,N_6784);
xor U10037 (N_10037,N_6483,N_6759);
xnor U10038 (N_10038,N_8863,N_8551);
xor U10039 (N_10039,N_6669,N_6148);
or U10040 (N_10040,N_7928,N_7824);
nand U10041 (N_10041,N_6562,N_7046);
xor U10042 (N_10042,N_8602,N_7622);
or U10043 (N_10043,N_6776,N_6680);
or U10044 (N_10044,N_8018,N_8230);
nand U10045 (N_10045,N_8731,N_6688);
or U10046 (N_10046,N_7729,N_8853);
or U10047 (N_10047,N_7015,N_8526);
nor U10048 (N_10048,N_6692,N_8030);
and U10049 (N_10049,N_7461,N_8255);
nand U10050 (N_10050,N_7039,N_7406);
nand U10051 (N_10051,N_8672,N_6234);
and U10052 (N_10052,N_8561,N_6706);
nor U10053 (N_10053,N_6302,N_6402);
or U10054 (N_10054,N_8338,N_6351);
nand U10055 (N_10055,N_8579,N_8169);
nand U10056 (N_10056,N_7279,N_6944);
and U10057 (N_10057,N_8309,N_6819);
nand U10058 (N_10058,N_8940,N_7555);
and U10059 (N_10059,N_8802,N_7145);
and U10060 (N_10060,N_8525,N_8949);
nand U10061 (N_10061,N_7450,N_8918);
or U10062 (N_10062,N_8118,N_6086);
nor U10063 (N_10063,N_6480,N_8101);
nand U10064 (N_10064,N_7565,N_7499);
and U10065 (N_10065,N_6490,N_7488);
nand U10066 (N_10066,N_8510,N_6770);
nand U10067 (N_10067,N_6579,N_8390);
and U10068 (N_10068,N_7202,N_8614);
and U10069 (N_10069,N_6215,N_6807);
or U10070 (N_10070,N_7159,N_8870);
and U10071 (N_10071,N_8860,N_8629);
or U10072 (N_10072,N_6235,N_6830);
and U10073 (N_10073,N_8991,N_7595);
or U10074 (N_10074,N_7407,N_7606);
nor U10075 (N_10075,N_7369,N_7522);
and U10076 (N_10076,N_7267,N_6676);
nor U10077 (N_10077,N_6367,N_7024);
and U10078 (N_10078,N_6478,N_6941);
or U10079 (N_10079,N_6356,N_7269);
or U10080 (N_10080,N_6633,N_6446);
or U10081 (N_10081,N_7110,N_6129);
nand U10082 (N_10082,N_8776,N_7531);
nand U10083 (N_10083,N_8504,N_6853);
or U10084 (N_10084,N_8548,N_6101);
nand U10085 (N_10085,N_7768,N_6441);
nor U10086 (N_10086,N_8593,N_7320);
or U10087 (N_10087,N_7493,N_8129);
nor U10088 (N_10088,N_8432,N_8800);
and U10089 (N_10089,N_6309,N_7268);
nor U10090 (N_10090,N_6425,N_6284);
nand U10091 (N_10091,N_7785,N_7482);
or U10092 (N_10092,N_8368,N_7379);
nor U10093 (N_10093,N_8795,N_8788);
or U10094 (N_10094,N_8698,N_6456);
nand U10095 (N_10095,N_7203,N_8232);
nor U10096 (N_10096,N_7518,N_6937);
nand U10097 (N_10097,N_8733,N_8425);
and U10098 (N_10098,N_8084,N_7334);
and U10099 (N_10099,N_7989,N_8571);
and U10100 (N_10100,N_8783,N_6541);
or U10101 (N_10101,N_6127,N_6567);
or U10102 (N_10102,N_7270,N_8221);
or U10103 (N_10103,N_7198,N_6341);
xnor U10104 (N_10104,N_8143,N_6123);
nand U10105 (N_10105,N_6517,N_7417);
or U10106 (N_10106,N_8495,N_8216);
xnor U10107 (N_10107,N_6162,N_7257);
and U10108 (N_10108,N_6721,N_8320);
and U10109 (N_10109,N_6115,N_8409);
nor U10110 (N_10110,N_8535,N_7448);
and U10111 (N_10111,N_7153,N_8832);
or U10112 (N_10112,N_7774,N_6485);
and U10113 (N_10113,N_8966,N_7285);
and U10114 (N_10114,N_8316,N_7820);
or U10115 (N_10115,N_7915,N_8321);
nor U10116 (N_10116,N_8274,N_6232);
nand U10117 (N_10117,N_8965,N_6832);
nand U10118 (N_10118,N_6313,N_6420);
xnor U10119 (N_10119,N_6053,N_8545);
xnor U10120 (N_10120,N_6543,N_7525);
nand U10121 (N_10121,N_8619,N_8546);
nor U10122 (N_10122,N_6820,N_8297);
and U10123 (N_10123,N_7021,N_7463);
and U10124 (N_10124,N_6461,N_7947);
nor U10125 (N_10125,N_6874,N_7002);
nor U10126 (N_10126,N_7264,N_7535);
or U10127 (N_10127,N_8073,N_6487);
nor U10128 (N_10128,N_8565,N_8715);
nand U10129 (N_10129,N_8669,N_8670);
and U10130 (N_10130,N_7619,N_7346);
xor U10131 (N_10131,N_6296,N_8954);
nor U10132 (N_10132,N_6144,N_8400);
and U10133 (N_10133,N_7252,N_7674);
nor U10134 (N_10134,N_7065,N_8340);
or U10135 (N_10135,N_8231,N_6580);
or U10136 (N_10136,N_6913,N_8491);
and U10137 (N_10137,N_7057,N_8661);
or U10138 (N_10138,N_7690,N_7438);
and U10139 (N_10139,N_8772,N_6697);
xnor U10140 (N_10140,N_7008,N_8924);
nand U10141 (N_10141,N_7236,N_7618);
or U10142 (N_10142,N_6287,N_6269);
nor U10143 (N_10143,N_8758,N_6955);
xnor U10144 (N_10144,N_6409,N_8265);
nand U10145 (N_10145,N_8770,N_8825);
or U10146 (N_10146,N_6978,N_6141);
and U10147 (N_10147,N_7506,N_6381);
nor U10148 (N_10148,N_8354,N_7602);
or U10149 (N_10149,N_7657,N_6529);
nor U10150 (N_10150,N_7526,N_8709);
nor U10151 (N_10151,N_6876,N_6279);
or U10152 (N_10152,N_6243,N_6735);
nand U10153 (N_10153,N_6519,N_8006);
or U10154 (N_10154,N_7007,N_8342);
nand U10155 (N_10155,N_8471,N_7142);
nand U10156 (N_10156,N_7309,N_6711);
or U10157 (N_10157,N_6099,N_8609);
xor U10158 (N_10158,N_8079,N_7646);
nand U10159 (N_10159,N_7079,N_7715);
xor U10160 (N_10160,N_7944,N_8550);
or U10161 (N_10161,N_7050,N_6821);
nand U10162 (N_10162,N_6612,N_7533);
or U10163 (N_10163,N_7327,N_6616);
and U10164 (N_10164,N_6346,N_6548);
or U10165 (N_10165,N_7156,N_8556);
and U10166 (N_10166,N_8171,N_6596);
or U10167 (N_10167,N_6276,N_8038);
nand U10168 (N_10168,N_8992,N_7467);
and U10169 (N_10169,N_7653,N_6438);
or U10170 (N_10170,N_8393,N_6066);
or U10171 (N_10171,N_8568,N_7056);
or U10172 (N_10172,N_8345,N_8904);
nor U10173 (N_10173,N_7812,N_6283);
nor U10174 (N_10174,N_7996,N_6431);
nand U10175 (N_10175,N_6404,N_8573);
nand U10176 (N_10176,N_8651,N_8557);
nor U10177 (N_10177,N_6623,N_8138);
nand U10178 (N_10178,N_8881,N_6624);
and U10179 (N_10179,N_6145,N_6724);
nor U10180 (N_10180,N_7377,N_6025);
xnor U10181 (N_10181,N_7781,N_6664);
nor U10182 (N_10182,N_8539,N_8880);
or U10183 (N_10183,N_7138,N_6322);
nor U10184 (N_10184,N_7985,N_8937);
nand U10185 (N_10185,N_7094,N_8438);
xor U10186 (N_10186,N_7716,N_6713);
nand U10187 (N_10187,N_6970,N_6500);
and U10188 (N_10188,N_8496,N_7034);
xnor U10189 (N_10189,N_8045,N_8945);
nor U10190 (N_10190,N_8584,N_8719);
and U10191 (N_10191,N_7801,N_6825);
and U10192 (N_10192,N_8569,N_6412);
nand U10193 (N_10193,N_6373,N_8178);
and U10194 (N_10194,N_6597,N_6787);
nand U10195 (N_10195,N_6729,N_8764);
or U10196 (N_10196,N_8074,N_7487);
and U10197 (N_10197,N_8174,N_7575);
and U10198 (N_10198,N_6361,N_7759);
nor U10199 (N_10199,N_6561,N_8222);
nor U10200 (N_10200,N_8906,N_8416);
nand U10201 (N_10201,N_8196,N_7629);
or U10202 (N_10202,N_7155,N_8703);
nor U10203 (N_10203,N_8373,N_6973);
nor U10204 (N_10204,N_8542,N_7688);
xor U10205 (N_10205,N_6969,N_8931);
and U10206 (N_10206,N_8826,N_8616);
or U10207 (N_10207,N_8293,N_7587);
or U10208 (N_10208,N_6755,N_7700);
and U10209 (N_10209,N_8238,N_6739);
and U10210 (N_10210,N_7137,N_7793);
nor U10211 (N_10211,N_8351,N_7254);
nor U10212 (N_10212,N_7300,N_8500);
xor U10213 (N_10213,N_7868,N_6029);
or U10214 (N_10214,N_8596,N_7923);
nand U10215 (N_10215,N_6864,N_8165);
or U10216 (N_10216,N_8646,N_6218);
and U10217 (N_10217,N_7539,N_7397);
and U10218 (N_10218,N_8915,N_7201);
nand U10219 (N_10219,N_7160,N_6390);
nor U10220 (N_10220,N_7435,N_8574);
nand U10221 (N_10221,N_6406,N_7953);
xor U10222 (N_10222,N_8717,N_8818);
nand U10223 (N_10223,N_6895,N_6350);
nor U10224 (N_10224,N_8830,N_6771);
nor U10225 (N_10225,N_7229,N_6036);
or U10226 (N_10226,N_6613,N_6702);
xor U10227 (N_10227,N_8498,N_6858);
or U10228 (N_10228,N_7497,N_7780);
xor U10229 (N_10229,N_6535,N_7476);
nand U10230 (N_10230,N_7365,N_6238);
nand U10231 (N_10231,N_7465,N_6372);
xor U10232 (N_10232,N_8017,N_8460);
and U10233 (N_10233,N_7164,N_7816);
or U10234 (N_10234,N_7707,N_6618);
and U10235 (N_10235,N_7668,N_6174);
and U10236 (N_10236,N_8440,N_7977);
nand U10237 (N_10237,N_8912,N_8326);
xnor U10238 (N_10238,N_6638,N_6964);
nand U10239 (N_10239,N_7669,N_8275);
nor U10240 (N_10240,N_7062,N_8585);
or U10241 (N_10241,N_7648,N_6470);
xnor U10242 (N_10242,N_7443,N_6001);
nand U10243 (N_10243,N_8241,N_8501);
xnor U10244 (N_10244,N_6432,N_7750);
xor U10245 (N_10245,N_7147,N_8827);
xor U10246 (N_10246,N_7351,N_8031);
nor U10247 (N_10247,N_6091,N_7704);
or U10248 (N_10248,N_7745,N_8183);
and U10249 (N_10249,N_6968,N_8406);
nand U10250 (N_10250,N_7391,N_7881);
or U10251 (N_10251,N_8152,N_7987);
xor U10252 (N_10252,N_7544,N_8513);
nand U10253 (N_10253,N_7218,N_8854);
nand U10254 (N_10254,N_6077,N_8789);
or U10255 (N_10255,N_7430,N_7945);
or U10256 (N_10256,N_6282,N_8347);
nand U10257 (N_10257,N_8161,N_8972);
nor U10258 (N_10258,N_6137,N_8775);
and U10259 (N_10259,N_8022,N_7519);
xnor U10260 (N_10260,N_8667,N_6110);
nor U10261 (N_10261,N_7459,N_7570);
or U10262 (N_10262,N_7609,N_7811);
or U10263 (N_10263,N_7192,N_7574);
or U10264 (N_10264,N_7756,N_7676);
xnor U10265 (N_10265,N_6750,N_6848);
or U10266 (N_10266,N_6411,N_7103);
nand U10267 (N_10267,N_7726,N_7567);
or U10268 (N_10268,N_8341,N_7009);
or U10269 (N_10269,N_6936,N_6231);
nand U10270 (N_10270,N_7471,N_6710);
xor U10271 (N_10271,N_7209,N_6682);
xor U10272 (N_10272,N_7962,N_6278);
nand U10273 (N_10273,N_7580,N_6554);
or U10274 (N_10274,N_7949,N_7739);
nand U10275 (N_10275,N_7994,N_7871);
nand U10276 (N_10276,N_8920,N_7894);
xnor U10277 (N_10277,N_8072,N_8815);
nand U10278 (N_10278,N_8163,N_7559);
nor U10279 (N_10279,N_6415,N_7044);
nand U10280 (N_10280,N_8388,N_8322);
or U10281 (N_10281,N_8261,N_7936);
xnor U10282 (N_10282,N_6920,N_7190);
xnor U10283 (N_10283,N_6736,N_6323);
nor U10284 (N_10284,N_6336,N_6694);
nor U10285 (N_10285,N_7524,N_7807);
or U10286 (N_10286,N_8164,N_8266);
xnor U10287 (N_10287,N_8615,N_8233);
or U10288 (N_10288,N_8947,N_6986);
nand U10289 (N_10289,N_7764,N_6966);
and U10290 (N_10290,N_7744,N_7163);
and U10291 (N_10291,N_8327,N_6872);
and U10292 (N_10292,N_7939,N_6507);
xor U10293 (N_10293,N_8838,N_6723);
and U10294 (N_10294,N_8153,N_7170);
or U10295 (N_10295,N_7969,N_6248);
or U10296 (N_10296,N_8876,N_8312);
nand U10297 (N_10297,N_6298,N_7850);
xor U10298 (N_10298,N_8260,N_7968);
and U10299 (N_10299,N_7386,N_6878);
nor U10300 (N_10300,N_6761,N_6443);
and U10301 (N_10301,N_8070,N_7611);
xnor U10302 (N_10302,N_8123,N_6502);
nand U10303 (N_10303,N_8528,N_7981);
xnor U10304 (N_10304,N_6542,N_6574);
and U10305 (N_10305,N_8479,N_6307);
or U10306 (N_10306,N_8250,N_7791);
nand U10307 (N_10307,N_7955,N_6695);
nor U10308 (N_10308,N_8599,N_7027);
nand U10309 (N_10309,N_8176,N_7143);
and U10310 (N_10310,N_6297,N_8660);
and U10311 (N_10311,N_6103,N_8455);
and U10312 (N_10312,N_6714,N_7248);
nor U10313 (N_10313,N_8710,N_7527);
and U10314 (N_10314,N_8458,N_6084);
nand U10315 (N_10315,N_8505,N_6207);
or U10316 (N_10316,N_8681,N_7437);
nor U10317 (N_10317,N_8057,N_7884);
and U10318 (N_10318,N_7265,N_6765);
xnor U10319 (N_10319,N_6557,N_7395);
or U10320 (N_10320,N_6126,N_8583);
and U10321 (N_10321,N_6100,N_7846);
xnor U10322 (N_10322,N_6146,N_7189);
or U10323 (N_10323,N_8979,N_6917);
or U10324 (N_10324,N_8156,N_8427);
nand U10325 (N_10325,N_6252,N_8292);
nand U10326 (N_10326,N_6801,N_6813);
or U10327 (N_10327,N_8026,N_8333);
nor U10328 (N_10328,N_7161,N_6753);
nand U10329 (N_10329,N_7898,N_8212);
nor U10330 (N_10330,N_7010,N_6834);
nor U10331 (N_10331,N_8431,N_7721);
xnor U10332 (N_10332,N_6794,N_6576);
xor U10333 (N_10333,N_8634,N_6930);
nand U10334 (N_10334,N_6663,N_7924);
nor U10335 (N_10335,N_6614,N_7376);
or U10336 (N_10336,N_8621,N_7645);
xnor U10337 (N_10337,N_7613,N_6240);
nor U10338 (N_10338,N_7183,N_7965);
nand U10339 (N_10339,N_6918,N_8182);
xnor U10340 (N_10340,N_7851,N_6119);
xnor U10341 (N_10341,N_8461,N_6398);
and U10342 (N_10342,N_6780,N_8928);
and U10343 (N_10343,N_8490,N_6746);
or U10344 (N_10344,N_6835,N_6338);
nor U10345 (N_10345,N_8623,N_8190);
nor U10346 (N_10346,N_8506,N_7400);
nor U10347 (N_10347,N_6880,N_7321);
nand U10348 (N_10348,N_8922,N_8706);
xnor U10349 (N_10349,N_8349,N_7144);
and U10350 (N_10350,N_6183,N_7828);
or U10351 (N_10351,N_8560,N_7671);
nor U10352 (N_10352,N_8380,N_8353);
xnor U10353 (N_10353,N_8739,N_7017);
nand U10354 (N_10354,N_6347,N_8996);
and U10355 (N_10355,N_6738,N_8857);
nand U10356 (N_10356,N_7691,N_8097);
nor U10357 (N_10357,N_7375,N_6716);
and U10358 (N_10358,N_7087,N_6847);
and U10359 (N_10359,N_6374,N_7698);
nand U10360 (N_10360,N_6340,N_6161);
nand U10361 (N_10361,N_7305,N_7043);
or U10362 (N_10362,N_6201,N_6774);
nor U10363 (N_10363,N_8939,N_7686);
or U10364 (N_10364,N_6164,N_7561);
xnor U10365 (N_10365,N_6353,N_7680);
nand U10366 (N_10366,N_7239,N_6644);
and U10367 (N_10367,N_8889,N_6095);
and U10368 (N_10368,N_8521,N_8896);
and U10369 (N_10369,N_8201,N_6072);
and U10370 (N_10370,N_8077,N_7710);
and U10371 (N_10371,N_8784,N_6588);
xor U10372 (N_10372,N_7444,N_7615);
nor U10373 (N_10373,N_6368,N_7743);
xor U10374 (N_10374,N_7244,N_6628);
nand U10375 (N_10375,N_6569,N_8811);
and U10376 (N_10376,N_6075,N_7130);
or U10377 (N_10377,N_8592,N_8415);
or U10378 (N_10378,N_6417,N_8591);
nand U10379 (N_10379,N_7474,N_6689);
nand U10380 (N_10380,N_7513,N_8121);
nor U10381 (N_10381,N_8210,N_7938);
and U10382 (N_10382,N_8306,N_7411);
nand U10383 (N_10383,N_6363,N_6553);
nor U10384 (N_10384,N_7455,N_6117);
and U10385 (N_10385,N_8520,N_7703);
nor U10386 (N_10386,N_7052,N_8732);
or U10387 (N_10387,N_7215,N_8377);
nand U10388 (N_10388,N_6521,N_8820);
nor U10389 (N_10389,N_8534,N_6782);
and U10390 (N_10390,N_8747,N_8209);
or U10391 (N_10391,N_6035,N_6246);
and U10392 (N_10392,N_6879,N_8339);
xnor U10393 (N_10393,N_6114,N_8611);
or U10394 (N_10394,N_8082,N_7810);
nor U10395 (N_10395,N_7162,N_6705);
and U10396 (N_10396,N_7983,N_7829);
nand U10397 (N_10397,N_7623,N_6043);
or U10398 (N_10398,N_8843,N_8310);
and U10399 (N_10399,N_6877,N_6857);
or U10400 (N_10400,N_7415,N_7230);
xor U10401 (N_10401,N_7099,N_8172);
nand U10402 (N_10402,N_7853,N_8147);
xnor U10403 (N_10403,N_6888,N_8882);
and U10404 (N_10404,N_7549,N_7380);
or U10405 (N_10405,N_6993,N_6915);
nor U10406 (N_10406,N_8384,N_6188);
nor U10407 (N_10407,N_6811,N_6814);
nand U10408 (N_10408,N_6657,N_8909);
nand U10409 (N_10409,N_7701,N_6727);
xnor U10410 (N_10410,N_8868,N_6370);
xor U10411 (N_10411,N_6178,N_8988);
xnor U10412 (N_10412,N_6522,N_7176);
xnor U10413 (N_10413,N_7167,N_7173);
nor U10414 (N_10414,N_6720,N_6945);
and U10415 (N_10415,N_7329,N_7586);
or U10416 (N_10416,N_8452,N_8944);
or U10417 (N_10417,N_7037,N_6923);
nor U10418 (N_10418,N_8677,N_7434);
xnor U10419 (N_10419,N_8470,N_7971);
nand U10420 (N_10420,N_8759,N_8051);
or U10421 (N_10421,N_8374,N_7843);
nand U10422 (N_10422,N_7188,N_7029);
and U10423 (N_10423,N_7564,N_6816);
nand U10424 (N_10424,N_7107,N_6400);
xnor U10425 (N_10425,N_7948,N_6627);
and U10426 (N_10426,N_8637,N_7874);
nand U10427 (N_10427,N_7754,N_7649);
xnor U10428 (N_10428,N_8892,N_8394);
nand U10429 (N_10429,N_7773,N_6063);
nand U10430 (N_10430,N_7808,N_6118);
or U10431 (N_10431,N_6290,N_7115);
and U10432 (N_10432,N_7362,N_7576);
xor U10433 (N_10433,N_7336,N_8655);
nand U10434 (N_10434,N_7446,N_6165);
xnor U10435 (N_10435,N_6499,N_6116);
nor U10436 (N_10436,N_8654,N_6728);
and U10437 (N_10437,N_6686,N_8877);
nand U10438 (N_10438,N_7330,N_7247);
or U10439 (N_10439,N_8259,N_8050);
nand U10440 (N_10440,N_7073,N_8608);
nand U10441 (N_10441,N_7067,N_6896);
or U10442 (N_10442,N_8434,N_8785);
and U10443 (N_10443,N_6591,N_7256);
nor U10444 (N_10444,N_7083,N_7308);
nor U10445 (N_10445,N_6060,N_6760);
nand U10446 (N_10446,N_6620,N_8069);
xor U10447 (N_10447,N_6514,N_7059);
or U10448 (N_10448,N_7001,N_6051);
or U10449 (N_10449,N_7498,N_8867);
xnor U10450 (N_10450,N_6838,N_8977);
nand U10451 (N_10451,N_8252,N_8774);
xor U10452 (N_10452,N_7158,N_6447);
nor U10453 (N_10453,N_6685,N_6242);
and U10454 (N_10454,N_6815,N_8554);
nor U10455 (N_10455,N_7148,N_6325);
xor U10456 (N_10456,N_8729,N_8463);
xnor U10457 (N_10457,N_7357,N_8995);
and U10458 (N_10458,N_6643,N_7178);
xnor U10459 (N_10459,N_7398,N_8519);
xor U10460 (N_10460,N_8034,N_7289);
and U10461 (N_10461,N_6958,N_6707);
or U10462 (N_10462,N_7751,N_7790);
and U10463 (N_10463,N_8688,N_8092);
or U10464 (N_10464,N_8958,N_6840);
and U10465 (N_10465,N_8308,N_8244);
and U10466 (N_10466,N_8577,N_8704);
nand U10467 (N_10467,N_7585,N_6850);
nor U10468 (N_10468,N_8831,N_6948);
nand U10469 (N_10469,N_6121,N_7684);
or U10470 (N_10470,N_7723,N_7695);
xor U10471 (N_10471,N_6111,N_7901);
xnor U10472 (N_10472,N_7036,N_6160);
and U10473 (N_10473,N_6932,N_6555);
or U10474 (N_10474,N_8911,N_8113);
or U10475 (N_10475,N_6228,N_7299);
or U10476 (N_10476,N_6730,N_8760);
nor U10477 (N_10477,N_7105,N_7326);
nand U10478 (N_10478,N_7013,N_7090);
nand U10479 (N_10479,N_8387,N_6866);
nor U10480 (N_10480,N_6186,N_7480);
and U10481 (N_10481,N_8976,N_7313);
xnor U10482 (N_10482,N_6849,N_6701);
nand U10483 (N_10483,N_8464,N_8442);
or U10484 (N_10484,N_8286,N_7310);
or U10485 (N_10485,N_6549,N_8687);
and U10486 (N_10486,N_6482,N_8061);
or U10487 (N_10487,N_7074,N_6581);
nor U10488 (N_10488,N_8436,N_6939);
xor U10489 (N_10489,N_8105,N_8134);
nor U10490 (N_10490,N_7030,N_8234);
and U10491 (N_10491,N_8957,N_6775);
nor U10492 (N_10492,N_6604,N_8559);
and U10493 (N_10493,N_8392,N_7659);
or U10494 (N_10494,N_6503,N_6991);
xnor U10495 (N_10495,N_8632,N_6852);
nand U10496 (N_10496,N_7084,N_8198);
or U10497 (N_10497,N_6033,N_6039);
nor U10498 (N_10498,N_8058,N_6209);
nor U10499 (N_10499,N_6808,N_6113);
xor U10500 (N_10500,N_6672,N_8106);
xnor U10501 (N_10501,N_6579,N_8578);
and U10502 (N_10502,N_8049,N_6209);
and U10503 (N_10503,N_7014,N_6169);
and U10504 (N_10504,N_7433,N_6596);
or U10505 (N_10505,N_7886,N_8584);
xnor U10506 (N_10506,N_6375,N_6582);
nand U10507 (N_10507,N_6082,N_6743);
nand U10508 (N_10508,N_8562,N_8310);
and U10509 (N_10509,N_8126,N_7903);
nand U10510 (N_10510,N_6487,N_7082);
or U10511 (N_10511,N_7714,N_8260);
xnor U10512 (N_10512,N_8988,N_6016);
or U10513 (N_10513,N_6023,N_7364);
or U10514 (N_10514,N_6477,N_7613);
or U10515 (N_10515,N_8891,N_8943);
xnor U10516 (N_10516,N_8213,N_7860);
nor U10517 (N_10517,N_6295,N_8060);
or U10518 (N_10518,N_8817,N_7327);
xor U10519 (N_10519,N_7318,N_6280);
nor U10520 (N_10520,N_7153,N_6093);
nand U10521 (N_10521,N_7007,N_8881);
nor U10522 (N_10522,N_7326,N_6863);
or U10523 (N_10523,N_6467,N_6777);
or U10524 (N_10524,N_7603,N_8602);
or U10525 (N_10525,N_6634,N_6363);
and U10526 (N_10526,N_6740,N_6313);
or U10527 (N_10527,N_6734,N_7135);
or U10528 (N_10528,N_7561,N_8417);
or U10529 (N_10529,N_8863,N_6649);
and U10530 (N_10530,N_8604,N_6450);
nand U10531 (N_10531,N_8060,N_7881);
xor U10532 (N_10532,N_8476,N_7602);
nand U10533 (N_10533,N_6439,N_7325);
nand U10534 (N_10534,N_8798,N_7767);
nor U10535 (N_10535,N_6068,N_8112);
and U10536 (N_10536,N_6923,N_6896);
or U10537 (N_10537,N_7751,N_6462);
xnor U10538 (N_10538,N_8702,N_7792);
nor U10539 (N_10539,N_8315,N_8213);
nor U10540 (N_10540,N_8391,N_6414);
xor U10541 (N_10541,N_6362,N_6237);
nand U10542 (N_10542,N_8146,N_6066);
nand U10543 (N_10543,N_7914,N_7094);
or U10544 (N_10544,N_8022,N_6638);
nand U10545 (N_10545,N_6803,N_7506);
nor U10546 (N_10546,N_7272,N_7501);
or U10547 (N_10547,N_8666,N_6443);
nor U10548 (N_10548,N_6704,N_6920);
nor U10549 (N_10549,N_7717,N_8538);
nand U10550 (N_10550,N_6920,N_7219);
and U10551 (N_10551,N_6790,N_7501);
nor U10552 (N_10552,N_8587,N_7887);
or U10553 (N_10553,N_6895,N_8911);
nand U10554 (N_10554,N_6989,N_8254);
nand U10555 (N_10555,N_6328,N_8095);
or U10556 (N_10556,N_6798,N_6867);
and U10557 (N_10557,N_7860,N_6778);
or U10558 (N_10558,N_7254,N_6524);
or U10559 (N_10559,N_7250,N_7377);
xnor U10560 (N_10560,N_8795,N_8583);
or U10561 (N_10561,N_8061,N_7384);
and U10562 (N_10562,N_6521,N_7965);
nand U10563 (N_10563,N_6378,N_8558);
xnor U10564 (N_10564,N_8941,N_8621);
and U10565 (N_10565,N_6203,N_6233);
and U10566 (N_10566,N_7719,N_8801);
nor U10567 (N_10567,N_6335,N_7667);
nand U10568 (N_10568,N_8382,N_8088);
nand U10569 (N_10569,N_7442,N_7268);
or U10570 (N_10570,N_6040,N_6546);
nand U10571 (N_10571,N_7341,N_7615);
or U10572 (N_10572,N_6083,N_7384);
and U10573 (N_10573,N_6032,N_6395);
and U10574 (N_10574,N_6361,N_7199);
and U10575 (N_10575,N_7709,N_6684);
or U10576 (N_10576,N_6217,N_6826);
nor U10577 (N_10577,N_6799,N_8150);
and U10578 (N_10578,N_6211,N_8439);
nor U10579 (N_10579,N_7728,N_7806);
nor U10580 (N_10580,N_7337,N_6162);
nor U10581 (N_10581,N_7231,N_8494);
or U10582 (N_10582,N_8606,N_6376);
xor U10583 (N_10583,N_8923,N_8016);
and U10584 (N_10584,N_7986,N_8603);
xnor U10585 (N_10585,N_6526,N_7311);
and U10586 (N_10586,N_8842,N_6421);
or U10587 (N_10587,N_7876,N_6159);
or U10588 (N_10588,N_7245,N_6595);
nand U10589 (N_10589,N_6292,N_7509);
nand U10590 (N_10590,N_6340,N_6617);
nor U10591 (N_10591,N_8846,N_6365);
or U10592 (N_10592,N_6489,N_6953);
nor U10593 (N_10593,N_7203,N_6747);
or U10594 (N_10594,N_8507,N_8165);
nand U10595 (N_10595,N_6729,N_7049);
xnor U10596 (N_10596,N_8303,N_7245);
and U10597 (N_10597,N_7284,N_7566);
xor U10598 (N_10598,N_7788,N_7614);
or U10599 (N_10599,N_8396,N_7851);
or U10600 (N_10600,N_8163,N_6110);
xnor U10601 (N_10601,N_8636,N_8172);
xnor U10602 (N_10602,N_8105,N_8926);
or U10603 (N_10603,N_6486,N_8432);
xnor U10604 (N_10604,N_8466,N_8301);
or U10605 (N_10605,N_6038,N_7107);
or U10606 (N_10606,N_6701,N_7383);
and U10607 (N_10607,N_7289,N_7284);
and U10608 (N_10608,N_7992,N_6561);
nand U10609 (N_10609,N_8413,N_7577);
xnor U10610 (N_10610,N_6568,N_8481);
nand U10611 (N_10611,N_8389,N_7181);
xnor U10612 (N_10612,N_7290,N_8201);
or U10613 (N_10613,N_6891,N_6100);
or U10614 (N_10614,N_8578,N_6637);
or U10615 (N_10615,N_8818,N_7260);
nor U10616 (N_10616,N_7067,N_6616);
nand U10617 (N_10617,N_6797,N_7528);
nor U10618 (N_10618,N_7422,N_8766);
and U10619 (N_10619,N_7562,N_7326);
and U10620 (N_10620,N_8919,N_7813);
xor U10621 (N_10621,N_8230,N_8990);
and U10622 (N_10622,N_6713,N_7348);
and U10623 (N_10623,N_6957,N_8589);
nand U10624 (N_10624,N_6525,N_8363);
and U10625 (N_10625,N_7761,N_8574);
nand U10626 (N_10626,N_6120,N_8355);
or U10627 (N_10627,N_8460,N_7586);
and U10628 (N_10628,N_6912,N_8392);
nor U10629 (N_10629,N_8807,N_7033);
nor U10630 (N_10630,N_6118,N_8655);
nor U10631 (N_10631,N_8772,N_8165);
and U10632 (N_10632,N_6979,N_8964);
nor U10633 (N_10633,N_7811,N_7161);
xor U10634 (N_10634,N_7935,N_6459);
xnor U10635 (N_10635,N_7268,N_8010);
or U10636 (N_10636,N_7334,N_7162);
nor U10637 (N_10637,N_8274,N_7793);
or U10638 (N_10638,N_6440,N_7113);
nand U10639 (N_10639,N_7332,N_6356);
nand U10640 (N_10640,N_6300,N_8103);
xor U10641 (N_10641,N_7075,N_7871);
and U10642 (N_10642,N_7127,N_7034);
or U10643 (N_10643,N_8392,N_8370);
xnor U10644 (N_10644,N_6794,N_7153);
nor U10645 (N_10645,N_6349,N_6634);
and U10646 (N_10646,N_6735,N_7648);
nor U10647 (N_10647,N_6336,N_6003);
nand U10648 (N_10648,N_6851,N_7610);
nand U10649 (N_10649,N_6693,N_8713);
nor U10650 (N_10650,N_8676,N_8501);
nand U10651 (N_10651,N_8656,N_8332);
nand U10652 (N_10652,N_7037,N_6612);
nor U10653 (N_10653,N_6687,N_6199);
or U10654 (N_10654,N_7832,N_8021);
nor U10655 (N_10655,N_7991,N_8733);
or U10656 (N_10656,N_6245,N_7082);
and U10657 (N_10657,N_7114,N_7434);
nor U10658 (N_10658,N_6882,N_7860);
nand U10659 (N_10659,N_6080,N_8940);
xor U10660 (N_10660,N_7368,N_6774);
or U10661 (N_10661,N_7283,N_7348);
nor U10662 (N_10662,N_8837,N_8119);
nand U10663 (N_10663,N_8243,N_6527);
xnor U10664 (N_10664,N_6054,N_8327);
or U10665 (N_10665,N_8772,N_8254);
xnor U10666 (N_10666,N_6024,N_7753);
xnor U10667 (N_10667,N_8634,N_8884);
nor U10668 (N_10668,N_7832,N_8275);
or U10669 (N_10669,N_6853,N_7771);
nand U10670 (N_10670,N_7165,N_7194);
nor U10671 (N_10671,N_7439,N_7875);
and U10672 (N_10672,N_6978,N_7613);
nor U10673 (N_10673,N_8603,N_6941);
and U10674 (N_10674,N_8058,N_7024);
or U10675 (N_10675,N_8567,N_7719);
nor U10676 (N_10676,N_8739,N_8026);
xnor U10677 (N_10677,N_7332,N_7821);
nand U10678 (N_10678,N_8126,N_8474);
xor U10679 (N_10679,N_7614,N_7543);
and U10680 (N_10680,N_8689,N_7623);
xor U10681 (N_10681,N_8421,N_8155);
nor U10682 (N_10682,N_7557,N_6864);
and U10683 (N_10683,N_6333,N_7944);
nor U10684 (N_10684,N_6069,N_7849);
nor U10685 (N_10685,N_8132,N_6947);
nand U10686 (N_10686,N_8286,N_8703);
nor U10687 (N_10687,N_7771,N_7795);
and U10688 (N_10688,N_6435,N_6290);
and U10689 (N_10689,N_8654,N_6629);
and U10690 (N_10690,N_8862,N_8917);
nand U10691 (N_10691,N_7871,N_7577);
nand U10692 (N_10692,N_7776,N_7354);
nor U10693 (N_10693,N_8024,N_8226);
nor U10694 (N_10694,N_8602,N_6562);
or U10695 (N_10695,N_7576,N_6687);
xnor U10696 (N_10696,N_6035,N_7014);
xor U10697 (N_10697,N_8243,N_6221);
nand U10698 (N_10698,N_6171,N_8327);
and U10699 (N_10699,N_7277,N_7388);
nand U10700 (N_10700,N_7603,N_8748);
nor U10701 (N_10701,N_6315,N_8789);
xnor U10702 (N_10702,N_6442,N_7358);
and U10703 (N_10703,N_8102,N_6868);
xnor U10704 (N_10704,N_8860,N_7340);
xnor U10705 (N_10705,N_7877,N_7339);
or U10706 (N_10706,N_7186,N_6233);
and U10707 (N_10707,N_6829,N_7831);
nor U10708 (N_10708,N_6944,N_6676);
and U10709 (N_10709,N_8112,N_8418);
xnor U10710 (N_10710,N_6118,N_7290);
xnor U10711 (N_10711,N_8529,N_7259);
nand U10712 (N_10712,N_6007,N_8192);
and U10713 (N_10713,N_7080,N_6933);
nand U10714 (N_10714,N_6195,N_6244);
and U10715 (N_10715,N_8791,N_6640);
xor U10716 (N_10716,N_8368,N_6674);
xor U10717 (N_10717,N_6242,N_8607);
nand U10718 (N_10718,N_6263,N_6603);
nor U10719 (N_10719,N_6057,N_8053);
nand U10720 (N_10720,N_8170,N_8400);
nand U10721 (N_10721,N_7464,N_7856);
or U10722 (N_10722,N_7245,N_8974);
nor U10723 (N_10723,N_6850,N_8856);
nand U10724 (N_10724,N_7781,N_7478);
or U10725 (N_10725,N_7910,N_7547);
xnor U10726 (N_10726,N_8710,N_6267);
nor U10727 (N_10727,N_6182,N_6358);
or U10728 (N_10728,N_8652,N_6908);
nor U10729 (N_10729,N_7571,N_6572);
nand U10730 (N_10730,N_8414,N_8389);
nor U10731 (N_10731,N_8190,N_6438);
xnor U10732 (N_10732,N_8792,N_6133);
nor U10733 (N_10733,N_6424,N_6142);
and U10734 (N_10734,N_6894,N_6977);
or U10735 (N_10735,N_7958,N_6087);
nand U10736 (N_10736,N_6437,N_6320);
or U10737 (N_10737,N_6007,N_7091);
xor U10738 (N_10738,N_8704,N_8527);
xnor U10739 (N_10739,N_7995,N_8275);
or U10740 (N_10740,N_8001,N_8139);
nor U10741 (N_10741,N_8771,N_8596);
and U10742 (N_10742,N_8393,N_7508);
or U10743 (N_10743,N_8590,N_7638);
or U10744 (N_10744,N_6185,N_7367);
nand U10745 (N_10745,N_7058,N_8623);
nor U10746 (N_10746,N_7213,N_6782);
nand U10747 (N_10747,N_7786,N_8537);
nand U10748 (N_10748,N_6705,N_6117);
and U10749 (N_10749,N_8971,N_8411);
nor U10750 (N_10750,N_7638,N_8656);
xnor U10751 (N_10751,N_7363,N_8275);
xnor U10752 (N_10752,N_6983,N_6059);
nand U10753 (N_10753,N_7103,N_8080);
and U10754 (N_10754,N_6507,N_6872);
and U10755 (N_10755,N_8188,N_6722);
xnor U10756 (N_10756,N_6053,N_6334);
and U10757 (N_10757,N_6321,N_6007);
or U10758 (N_10758,N_8304,N_6275);
nor U10759 (N_10759,N_7380,N_7936);
xnor U10760 (N_10760,N_6338,N_6158);
or U10761 (N_10761,N_6932,N_7215);
or U10762 (N_10762,N_7604,N_6899);
or U10763 (N_10763,N_8309,N_6730);
or U10764 (N_10764,N_6409,N_8996);
and U10765 (N_10765,N_8466,N_6928);
or U10766 (N_10766,N_8716,N_7711);
xor U10767 (N_10767,N_6836,N_8149);
and U10768 (N_10768,N_8961,N_7144);
xor U10769 (N_10769,N_6859,N_6913);
nor U10770 (N_10770,N_8396,N_6088);
xnor U10771 (N_10771,N_6823,N_6275);
xor U10772 (N_10772,N_8030,N_7846);
xnor U10773 (N_10773,N_7090,N_7153);
or U10774 (N_10774,N_7936,N_8954);
xor U10775 (N_10775,N_7960,N_6567);
nor U10776 (N_10776,N_7838,N_8738);
nor U10777 (N_10777,N_8135,N_8392);
and U10778 (N_10778,N_7251,N_6542);
nand U10779 (N_10779,N_8423,N_6572);
nand U10780 (N_10780,N_8219,N_6241);
nor U10781 (N_10781,N_8956,N_7021);
nand U10782 (N_10782,N_6477,N_6701);
nor U10783 (N_10783,N_8508,N_6010);
xnor U10784 (N_10784,N_8868,N_7059);
nand U10785 (N_10785,N_8469,N_7460);
and U10786 (N_10786,N_6657,N_8041);
or U10787 (N_10787,N_7604,N_6869);
xor U10788 (N_10788,N_7759,N_6233);
xnor U10789 (N_10789,N_8632,N_8965);
nand U10790 (N_10790,N_8381,N_8263);
xnor U10791 (N_10791,N_8711,N_6410);
and U10792 (N_10792,N_7941,N_7381);
xor U10793 (N_10793,N_7403,N_7717);
nand U10794 (N_10794,N_7295,N_6906);
nor U10795 (N_10795,N_8079,N_6063);
xor U10796 (N_10796,N_8365,N_8458);
xor U10797 (N_10797,N_8728,N_7555);
nand U10798 (N_10798,N_8167,N_7118);
nor U10799 (N_10799,N_8209,N_7535);
and U10800 (N_10800,N_7537,N_7049);
xnor U10801 (N_10801,N_6673,N_8523);
xor U10802 (N_10802,N_8608,N_8542);
nor U10803 (N_10803,N_8303,N_7817);
or U10804 (N_10804,N_6571,N_6487);
and U10805 (N_10805,N_7083,N_7340);
nor U10806 (N_10806,N_7855,N_6469);
or U10807 (N_10807,N_8552,N_6130);
nand U10808 (N_10808,N_7024,N_6658);
nor U10809 (N_10809,N_8280,N_6995);
xnor U10810 (N_10810,N_8756,N_8920);
and U10811 (N_10811,N_8980,N_6761);
or U10812 (N_10812,N_6480,N_7052);
or U10813 (N_10813,N_6211,N_8522);
nand U10814 (N_10814,N_6448,N_8727);
nand U10815 (N_10815,N_6272,N_7104);
and U10816 (N_10816,N_7678,N_6643);
nand U10817 (N_10817,N_6911,N_8222);
nor U10818 (N_10818,N_7508,N_8741);
nand U10819 (N_10819,N_6586,N_6901);
xor U10820 (N_10820,N_6596,N_8177);
nor U10821 (N_10821,N_6316,N_6380);
nand U10822 (N_10822,N_6568,N_6703);
or U10823 (N_10823,N_8872,N_8472);
xor U10824 (N_10824,N_8802,N_6959);
nor U10825 (N_10825,N_8420,N_8618);
and U10826 (N_10826,N_8032,N_7078);
xor U10827 (N_10827,N_8654,N_6156);
nor U10828 (N_10828,N_7877,N_6687);
or U10829 (N_10829,N_7448,N_7306);
nand U10830 (N_10830,N_8284,N_7647);
nor U10831 (N_10831,N_8992,N_8059);
xnor U10832 (N_10832,N_7830,N_8667);
nand U10833 (N_10833,N_6554,N_6539);
and U10834 (N_10834,N_7393,N_6838);
or U10835 (N_10835,N_6167,N_8412);
or U10836 (N_10836,N_7906,N_6399);
xnor U10837 (N_10837,N_7228,N_6504);
nand U10838 (N_10838,N_7978,N_6582);
nor U10839 (N_10839,N_7041,N_7991);
xnor U10840 (N_10840,N_8121,N_7922);
xnor U10841 (N_10841,N_8784,N_7476);
xor U10842 (N_10842,N_6191,N_7873);
xor U10843 (N_10843,N_6693,N_8605);
nand U10844 (N_10844,N_7261,N_7599);
and U10845 (N_10845,N_6801,N_6195);
or U10846 (N_10846,N_8261,N_8974);
xor U10847 (N_10847,N_8542,N_6214);
or U10848 (N_10848,N_8391,N_8045);
and U10849 (N_10849,N_6250,N_7530);
nor U10850 (N_10850,N_8148,N_7999);
nor U10851 (N_10851,N_6738,N_6653);
or U10852 (N_10852,N_8857,N_6111);
and U10853 (N_10853,N_6148,N_8229);
and U10854 (N_10854,N_8161,N_8879);
nor U10855 (N_10855,N_6622,N_7103);
xor U10856 (N_10856,N_6888,N_8698);
nor U10857 (N_10857,N_6602,N_6749);
or U10858 (N_10858,N_7739,N_6426);
xnor U10859 (N_10859,N_8651,N_8798);
xor U10860 (N_10860,N_6877,N_8747);
and U10861 (N_10861,N_6632,N_7015);
xor U10862 (N_10862,N_7820,N_8600);
nor U10863 (N_10863,N_6155,N_6124);
nand U10864 (N_10864,N_7345,N_7782);
or U10865 (N_10865,N_6521,N_6308);
nand U10866 (N_10866,N_8441,N_7072);
or U10867 (N_10867,N_8052,N_6756);
nor U10868 (N_10868,N_6624,N_7731);
nor U10869 (N_10869,N_6016,N_7793);
nor U10870 (N_10870,N_7745,N_8755);
nand U10871 (N_10871,N_7809,N_6483);
and U10872 (N_10872,N_6540,N_8539);
xor U10873 (N_10873,N_7635,N_7685);
xor U10874 (N_10874,N_6617,N_6957);
nand U10875 (N_10875,N_6330,N_6820);
nor U10876 (N_10876,N_7078,N_8592);
and U10877 (N_10877,N_7554,N_8328);
or U10878 (N_10878,N_7821,N_7097);
or U10879 (N_10879,N_7080,N_6837);
nand U10880 (N_10880,N_8466,N_8129);
and U10881 (N_10881,N_8558,N_7670);
nand U10882 (N_10882,N_6245,N_6804);
nand U10883 (N_10883,N_7666,N_6279);
and U10884 (N_10884,N_7364,N_8145);
and U10885 (N_10885,N_6305,N_6281);
nor U10886 (N_10886,N_6426,N_8602);
nor U10887 (N_10887,N_8371,N_8271);
or U10888 (N_10888,N_8583,N_8928);
nand U10889 (N_10889,N_8160,N_7749);
xnor U10890 (N_10890,N_8212,N_6923);
xnor U10891 (N_10891,N_6662,N_6056);
or U10892 (N_10892,N_7609,N_7339);
nor U10893 (N_10893,N_6551,N_7637);
nor U10894 (N_10894,N_6536,N_7473);
xor U10895 (N_10895,N_7956,N_8116);
or U10896 (N_10896,N_7577,N_7047);
and U10897 (N_10897,N_8179,N_7909);
or U10898 (N_10898,N_7650,N_6263);
nor U10899 (N_10899,N_7732,N_8792);
and U10900 (N_10900,N_7066,N_6379);
nor U10901 (N_10901,N_6487,N_6691);
or U10902 (N_10902,N_7231,N_6570);
xor U10903 (N_10903,N_7846,N_8389);
xor U10904 (N_10904,N_8626,N_7996);
and U10905 (N_10905,N_6903,N_7715);
and U10906 (N_10906,N_8343,N_6937);
or U10907 (N_10907,N_7553,N_8899);
and U10908 (N_10908,N_8238,N_6788);
xor U10909 (N_10909,N_7746,N_6753);
or U10910 (N_10910,N_7160,N_8871);
and U10911 (N_10911,N_7490,N_6055);
xnor U10912 (N_10912,N_7503,N_7472);
nor U10913 (N_10913,N_7904,N_8504);
and U10914 (N_10914,N_7320,N_6871);
and U10915 (N_10915,N_8233,N_7887);
or U10916 (N_10916,N_7605,N_7586);
nor U10917 (N_10917,N_7254,N_6471);
or U10918 (N_10918,N_7060,N_6072);
xnor U10919 (N_10919,N_6347,N_8478);
or U10920 (N_10920,N_8522,N_6821);
nor U10921 (N_10921,N_6738,N_7796);
xnor U10922 (N_10922,N_6960,N_8419);
xnor U10923 (N_10923,N_6794,N_7853);
nor U10924 (N_10924,N_8138,N_7716);
nor U10925 (N_10925,N_6611,N_8421);
xor U10926 (N_10926,N_8260,N_8939);
nand U10927 (N_10927,N_6436,N_7761);
xor U10928 (N_10928,N_6767,N_7460);
nand U10929 (N_10929,N_6773,N_8703);
nor U10930 (N_10930,N_6659,N_6840);
and U10931 (N_10931,N_8495,N_7018);
or U10932 (N_10932,N_8638,N_6335);
and U10933 (N_10933,N_7917,N_6551);
nand U10934 (N_10934,N_7948,N_7016);
or U10935 (N_10935,N_7533,N_6602);
nor U10936 (N_10936,N_7321,N_8182);
nand U10937 (N_10937,N_8480,N_7585);
xor U10938 (N_10938,N_6194,N_6740);
and U10939 (N_10939,N_6132,N_8466);
xor U10940 (N_10940,N_8114,N_6311);
or U10941 (N_10941,N_7810,N_8766);
and U10942 (N_10942,N_8894,N_6494);
nand U10943 (N_10943,N_7841,N_7872);
and U10944 (N_10944,N_6376,N_6429);
nand U10945 (N_10945,N_6205,N_7527);
xor U10946 (N_10946,N_8967,N_7119);
or U10947 (N_10947,N_6227,N_6797);
nand U10948 (N_10948,N_7943,N_8649);
nor U10949 (N_10949,N_7286,N_7315);
xor U10950 (N_10950,N_6017,N_8640);
xor U10951 (N_10951,N_7047,N_7414);
nand U10952 (N_10952,N_7272,N_7707);
and U10953 (N_10953,N_8877,N_6913);
or U10954 (N_10954,N_8570,N_6834);
nand U10955 (N_10955,N_6100,N_7623);
xnor U10956 (N_10956,N_6749,N_8808);
and U10957 (N_10957,N_8512,N_8912);
and U10958 (N_10958,N_7211,N_7294);
or U10959 (N_10959,N_7579,N_8476);
nor U10960 (N_10960,N_8409,N_8544);
xnor U10961 (N_10961,N_6784,N_6102);
nand U10962 (N_10962,N_6358,N_7930);
or U10963 (N_10963,N_8129,N_6635);
and U10964 (N_10964,N_6870,N_6816);
nor U10965 (N_10965,N_7903,N_7013);
or U10966 (N_10966,N_7185,N_8662);
xor U10967 (N_10967,N_6795,N_7482);
nand U10968 (N_10968,N_6037,N_7099);
nor U10969 (N_10969,N_8255,N_6698);
and U10970 (N_10970,N_8275,N_7724);
and U10971 (N_10971,N_7536,N_6129);
nand U10972 (N_10972,N_8234,N_8847);
xnor U10973 (N_10973,N_6299,N_7584);
or U10974 (N_10974,N_8430,N_8023);
and U10975 (N_10975,N_7283,N_7972);
nand U10976 (N_10976,N_6793,N_8025);
or U10977 (N_10977,N_6103,N_6921);
nor U10978 (N_10978,N_8661,N_6205);
xnor U10979 (N_10979,N_6431,N_8133);
nor U10980 (N_10980,N_7248,N_7884);
nor U10981 (N_10981,N_7314,N_6182);
nor U10982 (N_10982,N_8219,N_6554);
and U10983 (N_10983,N_7902,N_7254);
nand U10984 (N_10984,N_8595,N_7781);
or U10985 (N_10985,N_7778,N_8833);
and U10986 (N_10986,N_7078,N_6241);
nand U10987 (N_10987,N_7393,N_6052);
or U10988 (N_10988,N_6441,N_6660);
or U10989 (N_10989,N_7434,N_7060);
and U10990 (N_10990,N_6315,N_7899);
nor U10991 (N_10991,N_7758,N_6304);
nor U10992 (N_10992,N_7968,N_7564);
xnor U10993 (N_10993,N_8121,N_8086);
xor U10994 (N_10994,N_8117,N_6165);
or U10995 (N_10995,N_8954,N_8673);
and U10996 (N_10996,N_6817,N_8900);
and U10997 (N_10997,N_6609,N_6584);
nor U10998 (N_10998,N_7197,N_6795);
nand U10999 (N_10999,N_7184,N_8547);
nand U11000 (N_11000,N_7786,N_7366);
nand U11001 (N_11001,N_8837,N_7690);
xor U11002 (N_11002,N_8736,N_7675);
xor U11003 (N_11003,N_6854,N_8078);
nand U11004 (N_11004,N_7951,N_7804);
nand U11005 (N_11005,N_8364,N_7185);
xor U11006 (N_11006,N_8800,N_8806);
and U11007 (N_11007,N_8487,N_6521);
xnor U11008 (N_11008,N_7954,N_8069);
and U11009 (N_11009,N_6975,N_6085);
nand U11010 (N_11010,N_6782,N_7838);
nor U11011 (N_11011,N_8822,N_6031);
xnor U11012 (N_11012,N_6789,N_8365);
xnor U11013 (N_11013,N_8272,N_7953);
and U11014 (N_11014,N_6460,N_8370);
nand U11015 (N_11015,N_8363,N_7476);
nand U11016 (N_11016,N_8075,N_6577);
nand U11017 (N_11017,N_6740,N_8437);
nand U11018 (N_11018,N_8242,N_6089);
nor U11019 (N_11019,N_6184,N_8660);
nor U11020 (N_11020,N_7444,N_7943);
and U11021 (N_11021,N_8432,N_8295);
nand U11022 (N_11022,N_6682,N_7388);
xor U11023 (N_11023,N_7400,N_7011);
nand U11024 (N_11024,N_7909,N_6766);
and U11025 (N_11025,N_8026,N_6773);
nor U11026 (N_11026,N_7683,N_6131);
or U11027 (N_11027,N_8727,N_6556);
and U11028 (N_11028,N_7278,N_7406);
nand U11029 (N_11029,N_8365,N_8638);
and U11030 (N_11030,N_8399,N_7609);
or U11031 (N_11031,N_8997,N_6786);
nand U11032 (N_11032,N_8872,N_8878);
or U11033 (N_11033,N_8841,N_7568);
or U11034 (N_11034,N_8092,N_8564);
nor U11035 (N_11035,N_7850,N_7158);
and U11036 (N_11036,N_6768,N_6362);
or U11037 (N_11037,N_6926,N_8586);
nor U11038 (N_11038,N_6259,N_8148);
and U11039 (N_11039,N_7741,N_7299);
xnor U11040 (N_11040,N_7072,N_7764);
or U11041 (N_11041,N_8900,N_7222);
or U11042 (N_11042,N_8184,N_6246);
nand U11043 (N_11043,N_8322,N_7040);
and U11044 (N_11044,N_8080,N_7644);
nand U11045 (N_11045,N_7579,N_6872);
and U11046 (N_11046,N_7428,N_7430);
or U11047 (N_11047,N_6472,N_8854);
xnor U11048 (N_11048,N_6171,N_6317);
nand U11049 (N_11049,N_6925,N_6776);
nand U11050 (N_11050,N_6383,N_6747);
nor U11051 (N_11051,N_6761,N_7752);
xnor U11052 (N_11052,N_7123,N_6438);
nand U11053 (N_11053,N_8092,N_8832);
or U11054 (N_11054,N_6570,N_8010);
or U11055 (N_11055,N_8741,N_8802);
nor U11056 (N_11056,N_8180,N_6760);
nor U11057 (N_11057,N_8466,N_8035);
xnor U11058 (N_11058,N_8702,N_7872);
or U11059 (N_11059,N_6855,N_8409);
xor U11060 (N_11060,N_7158,N_7578);
xor U11061 (N_11061,N_7485,N_6738);
and U11062 (N_11062,N_6088,N_7682);
nand U11063 (N_11063,N_7438,N_7251);
nand U11064 (N_11064,N_7994,N_7438);
nand U11065 (N_11065,N_8508,N_7215);
and U11066 (N_11066,N_8415,N_8744);
xnor U11067 (N_11067,N_7486,N_8661);
xnor U11068 (N_11068,N_7952,N_7667);
nor U11069 (N_11069,N_7142,N_6745);
nor U11070 (N_11070,N_7152,N_7068);
or U11071 (N_11071,N_6444,N_7732);
nand U11072 (N_11072,N_8590,N_7483);
nor U11073 (N_11073,N_6132,N_6439);
and U11074 (N_11074,N_6491,N_7245);
nor U11075 (N_11075,N_8889,N_7816);
nand U11076 (N_11076,N_6687,N_7467);
or U11077 (N_11077,N_6003,N_6202);
nand U11078 (N_11078,N_7055,N_6621);
xnor U11079 (N_11079,N_6023,N_7849);
nand U11080 (N_11080,N_7520,N_7414);
xnor U11081 (N_11081,N_7814,N_6266);
or U11082 (N_11082,N_6205,N_7719);
or U11083 (N_11083,N_6698,N_7111);
and U11084 (N_11084,N_6139,N_7107);
xor U11085 (N_11085,N_7717,N_8456);
and U11086 (N_11086,N_8619,N_8278);
and U11087 (N_11087,N_8026,N_6540);
and U11088 (N_11088,N_7463,N_8452);
or U11089 (N_11089,N_7163,N_7754);
nand U11090 (N_11090,N_6708,N_8108);
nand U11091 (N_11091,N_6623,N_7171);
and U11092 (N_11092,N_8168,N_6384);
xnor U11093 (N_11093,N_7241,N_8411);
xor U11094 (N_11094,N_8444,N_7630);
and U11095 (N_11095,N_8464,N_6402);
xnor U11096 (N_11096,N_6445,N_8534);
nand U11097 (N_11097,N_7510,N_8115);
nor U11098 (N_11098,N_8396,N_7345);
and U11099 (N_11099,N_6534,N_6117);
or U11100 (N_11100,N_7860,N_8544);
nand U11101 (N_11101,N_6067,N_8995);
nor U11102 (N_11102,N_7605,N_6935);
and U11103 (N_11103,N_7376,N_7469);
or U11104 (N_11104,N_7413,N_8671);
nor U11105 (N_11105,N_8374,N_7371);
xor U11106 (N_11106,N_6896,N_8248);
xnor U11107 (N_11107,N_8402,N_7468);
and U11108 (N_11108,N_7258,N_8557);
nand U11109 (N_11109,N_7319,N_8980);
nand U11110 (N_11110,N_7188,N_6673);
nor U11111 (N_11111,N_6837,N_6811);
and U11112 (N_11112,N_6337,N_7471);
nor U11113 (N_11113,N_8397,N_7934);
nor U11114 (N_11114,N_8999,N_8019);
nand U11115 (N_11115,N_6019,N_7932);
nor U11116 (N_11116,N_7845,N_7293);
nor U11117 (N_11117,N_7225,N_6003);
and U11118 (N_11118,N_8534,N_8643);
or U11119 (N_11119,N_8297,N_6542);
and U11120 (N_11120,N_8297,N_6832);
nand U11121 (N_11121,N_6893,N_6415);
nand U11122 (N_11122,N_7684,N_7517);
or U11123 (N_11123,N_7724,N_7802);
and U11124 (N_11124,N_7838,N_6363);
xor U11125 (N_11125,N_6242,N_8698);
or U11126 (N_11126,N_6281,N_7240);
and U11127 (N_11127,N_7142,N_7489);
and U11128 (N_11128,N_8616,N_8163);
or U11129 (N_11129,N_7780,N_6473);
nand U11130 (N_11130,N_8916,N_8209);
xor U11131 (N_11131,N_7644,N_7235);
nor U11132 (N_11132,N_7134,N_6207);
xor U11133 (N_11133,N_8686,N_8000);
and U11134 (N_11134,N_7897,N_8274);
or U11135 (N_11135,N_8215,N_8138);
and U11136 (N_11136,N_7756,N_6609);
or U11137 (N_11137,N_8404,N_7148);
xor U11138 (N_11138,N_8515,N_8403);
nor U11139 (N_11139,N_7460,N_8763);
xor U11140 (N_11140,N_6777,N_7090);
and U11141 (N_11141,N_8070,N_8621);
or U11142 (N_11142,N_8272,N_8193);
nor U11143 (N_11143,N_6615,N_8340);
nor U11144 (N_11144,N_6075,N_6891);
nor U11145 (N_11145,N_7509,N_7981);
and U11146 (N_11146,N_8447,N_8761);
nand U11147 (N_11147,N_6503,N_6599);
and U11148 (N_11148,N_7312,N_7904);
xnor U11149 (N_11149,N_7508,N_6467);
nor U11150 (N_11150,N_6237,N_7467);
and U11151 (N_11151,N_7633,N_6019);
or U11152 (N_11152,N_8228,N_8582);
nand U11153 (N_11153,N_6295,N_6701);
nand U11154 (N_11154,N_7766,N_8527);
and U11155 (N_11155,N_6055,N_6165);
nand U11156 (N_11156,N_6461,N_7051);
and U11157 (N_11157,N_7293,N_7760);
and U11158 (N_11158,N_7773,N_8585);
nand U11159 (N_11159,N_7972,N_8954);
xnor U11160 (N_11160,N_7265,N_6214);
xnor U11161 (N_11161,N_6194,N_6965);
nand U11162 (N_11162,N_8720,N_8908);
xnor U11163 (N_11163,N_6675,N_7597);
xnor U11164 (N_11164,N_7294,N_7273);
nand U11165 (N_11165,N_6501,N_8435);
xnor U11166 (N_11166,N_7731,N_8765);
nand U11167 (N_11167,N_8454,N_7997);
nor U11168 (N_11168,N_6955,N_7424);
xor U11169 (N_11169,N_8299,N_7045);
nand U11170 (N_11170,N_7713,N_6032);
or U11171 (N_11171,N_6501,N_8203);
xnor U11172 (N_11172,N_6598,N_6272);
nor U11173 (N_11173,N_6226,N_6555);
xnor U11174 (N_11174,N_8819,N_7484);
nor U11175 (N_11175,N_6194,N_7552);
nor U11176 (N_11176,N_8954,N_8687);
xor U11177 (N_11177,N_7274,N_6747);
nor U11178 (N_11178,N_8880,N_6406);
or U11179 (N_11179,N_8614,N_8435);
and U11180 (N_11180,N_7021,N_6820);
and U11181 (N_11181,N_8940,N_6409);
or U11182 (N_11182,N_7034,N_7147);
nand U11183 (N_11183,N_8255,N_8404);
nand U11184 (N_11184,N_8372,N_6927);
nor U11185 (N_11185,N_6580,N_8240);
nor U11186 (N_11186,N_7629,N_8530);
nor U11187 (N_11187,N_6926,N_7439);
nor U11188 (N_11188,N_8076,N_6159);
nor U11189 (N_11189,N_8720,N_6771);
nor U11190 (N_11190,N_8033,N_8436);
xor U11191 (N_11191,N_6852,N_8580);
and U11192 (N_11192,N_6049,N_7575);
or U11193 (N_11193,N_8347,N_8548);
xnor U11194 (N_11194,N_8482,N_8995);
and U11195 (N_11195,N_8061,N_8372);
nand U11196 (N_11196,N_6041,N_8676);
and U11197 (N_11197,N_8228,N_6452);
and U11198 (N_11198,N_7502,N_7573);
nor U11199 (N_11199,N_8278,N_6540);
and U11200 (N_11200,N_8846,N_8713);
and U11201 (N_11201,N_8359,N_8545);
nand U11202 (N_11202,N_7477,N_8132);
nor U11203 (N_11203,N_7681,N_6676);
and U11204 (N_11204,N_6878,N_7172);
nor U11205 (N_11205,N_6988,N_6609);
and U11206 (N_11206,N_6698,N_8601);
or U11207 (N_11207,N_7127,N_8485);
nor U11208 (N_11208,N_8423,N_7038);
or U11209 (N_11209,N_8198,N_6169);
and U11210 (N_11210,N_7046,N_6378);
nor U11211 (N_11211,N_8229,N_8508);
nor U11212 (N_11212,N_7832,N_7248);
and U11213 (N_11213,N_6767,N_8296);
nor U11214 (N_11214,N_6923,N_6463);
and U11215 (N_11215,N_6178,N_6430);
nor U11216 (N_11216,N_6512,N_8887);
and U11217 (N_11217,N_6190,N_7729);
or U11218 (N_11218,N_8055,N_8250);
and U11219 (N_11219,N_8751,N_6513);
xor U11220 (N_11220,N_8272,N_7437);
or U11221 (N_11221,N_8320,N_8861);
or U11222 (N_11222,N_8498,N_8967);
or U11223 (N_11223,N_8511,N_6686);
xnor U11224 (N_11224,N_8411,N_6595);
xnor U11225 (N_11225,N_7607,N_6155);
nand U11226 (N_11226,N_7824,N_7550);
xnor U11227 (N_11227,N_6680,N_7724);
nand U11228 (N_11228,N_7602,N_7151);
nor U11229 (N_11229,N_8110,N_6522);
xnor U11230 (N_11230,N_7329,N_8755);
nand U11231 (N_11231,N_7851,N_6094);
nor U11232 (N_11232,N_7623,N_6284);
nor U11233 (N_11233,N_6143,N_8903);
and U11234 (N_11234,N_6070,N_8075);
nor U11235 (N_11235,N_7329,N_6147);
xnor U11236 (N_11236,N_8571,N_7516);
or U11237 (N_11237,N_7414,N_7104);
nor U11238 (N_11238,N_6397,N_6315);
xnor U11239 (N_11239,N_7865,N_8122);
xor U11240 (N_11240,N_6303,N_6929);
xnor U11241 (N_11241,N_6705,N_7047);
and U11242 (N_11242,N_7981,N_6960);
nand U11243 (N_11243,N_7742,N_7641);
or U11244 (N_11244,N_8975,N_7159);
nor U11245 (N_11245,N_8618,N_6374);
nor U11246 (N_11246,N_8958,N_7720);
nand U11247 (N_11247,N_7821,N_7091);
and U11248 (N_11248,N_8510,N_7847);
xor U11249 (N_11249,N_6653,N_6623);
nand U11250 (N_11250,N_8745,N_8776);
xnor U11251 (N_11251,N_7131,N_8618);
or U11252 (N_11252,N_8865,N_8002);
and U11253 (N_11253,N_6324,N_6823);
nor U11254 (N_11254,N_6184,N_7295);
nand U11255 (N_11255,N_8951,N_8056);
and U11256 (N_11256,N_8292,N_6395);
xor U11257 (N_11257,N_8885,N_7791);
xor U11258 (N_11258,N_8094,N_6937);
nor U11259 (N_11259,N_6344,N_6213);
nand U11260 (N_11260,N_6190,N_6186);
and U11261 (N_11261,N_7357,N_6327);
xnor U11262 (N_11262,N_7410,N_6386);
and U11263 (N_11263,N_8203,N_6811);
nand U11264 (N_11264,N_8388,N_6195);
xnor U11265 (N_11265,N_8182,N_8754);
nor U11266 (N_11266,N_8275,N_6304);
and U11267 (N_11267,N_8190,N_7362);
xnor U11268 (N_11268,N_6506,N_8811);
or U11269 (N_11269,N_7758,N_7744);
nor U11270 (N_11270,N_6670,N_6824);
and U11271 (N_11271,N_7428,N_7703);
nor U11272 (N_11272,N_6017,N_6498);
xnor U11273 (N_11273,N_8207,N_7673);
and U11274 (N_11274,N_7773,N_7026);
nor U11275 (N_11275,N_7315,N_8850);
or U11276 (N_11276,N_6639,N_8595);
and U11277 (N_11277,N_8161,N_7166);
nand U11278 (N_11278,N_6884,N_7679);
nand U11279 (N_11279,N_7744,N_8744);
and U11280 (N_11280,N_8375,N_7953);
xor U11281 (N_11281,N_8575,N_8978);
and U11282 (N_11282,N_6024,N_6713);
or U11283 (N_11283,N_8232,N_8984);
xnor U11284 (N_11284,N_8829,N_6036);
nor U11285 (N_11285,N_8152,N_6895);
xor U11286 (N_11286,N_6132,N_7702);
xor U11287 (N_11287,N_7352,N_6623);
nor U11288 (N_11288,N_7304,N_8080);
nand U11289 (N_11289,N_8138,N_7335);
nor U11290 (N_11290,N_6442,N_7988);
and U11291 (N_11291,N_8061,N_6502);
nand U11292 (N_11292,N_6825,N_6357);
nand U11293 (N_11293,N_8797,N_6059);
xnor U11294 (N_11294,N_6456,N_8230);
and U11295 (N_11295,N_8827,N_7435);
and U11296 (N_11296,N_7574,N_8703);
nand U11297 (N_11297,N_6585,N_8656);
xnor U11298 (N_11298,N_6731,N_8930);
xnor U11299 (N_11299,N_6452,N_8998);
nor U11300 (N_11300,N_7488,N_7517);
xnor U11301 (N_11301,N_6473,N_6225);
xnor U11302 (N_11302,N_7748,N_6630);
or U11303 (N_11303,N_7098,N_8152);
and U11304 (N_11304,N_7022,N_6410);
and U11305 (N_11305,N_6231,N_7627);
xor U11306 (N_11306,N_8924,N_6405);
and U11307 (N_11307,N_6192,N_6185);
nor U11308 (N_11308,N_6467,N_6393);
or U11309 (N_11309,N_7251,N_7643);
xnor U11310 (N_11310,N_8481,N_8879);
nor U11311 (N_11311,N_8856,N_7679);
and U11312 (N_11312,N_7636,N_8484);
or U11313 (N_11313,N_7160,N_8255);
and U11314 (N_11314,N_7552,N_6997);
or U11315 (N_11315,N_7856,N_7900);
or U11316 (N_11316,N_7237,N_7808);
nand U11317 (N_11317,N_7359,N_7928);
nor U11318 (N_11318,N_7732,N_6242);
or U11319 (N_11319,N_8711,N_6917);
nand U11320 (N_11320,N_6629,N_7657);
and U11321 (N_11321,N_6107,N_8843);
and U11322 (N_11322,N_8983,N_6155);
nand U11323 (N_11323,N_6187,N_7428);
xor U11324 (N_11324,N_8382,N_8175);
nor U11325 (N_11325,N_8342,N_7368);
nand U11326 (N_11326,N_8316,N_6868);
nor U11327 (N_11327,N_7235,N_6439);
nand U11328 (N_11328,N_8951,N_7083);
and U11329 (N_11329,N_6389,N_7057);
nand U11330 (N_11330,N_6002,N_6398);
nor U11331 (N_11331,N_7846,N_8052);
and U11332 (N_11332,N_6903,N_7837);
nor U11333 (N_11333,N_6132,N_7988);
xor U11334 (N_11334,N_6061,N_8228);
xnor U11335 (N_11335,N_6702,N_6315);
nor U11336 (N_11336,N_6954,N_7673);
xnor U11337 (N_11337,N_6979,N_8772);
nand U11338 (N_11338,N_7731,N_7347);
or U11339 (N_11339,N_8097,N_7346);
and U11340 (N_11340,N_8803,N_6729);
nand U11341 (N_11341,N_8566,N_8073);
and U11342 (N_11342,N_7058,N_6179);
nand U11343 (N_11343,N_6201,N_7745);
xor U11344 (N_11344,N_6030,N_6396);
and U11345 (N_11345,N_7916,N_7083);
and U11346 (N_11346,N_8115,N_7820);
or U11347 (N_11347,N_8401,N_7325);
and U11348 (N_11348,N_7271,N_8805);
xnor U11349 (N_11349,N_6491,N_6841);
xor U11350 (N_11350,N_8364,N_7688);
xnor U11351 (N_11351,N_6179,N_6369);
xnor U11352 (N_11352,N_6841,N_7166);
xor U11353 (N_11353,N_7971,N_6496);
xor U11354 (N_11354,N_8651,N_7540);
xnor U11355 (N_11355,N_6969,N_6280);
or U11356 (N_11356,N_6321,N_7612);
and U11357 (N_11357,N_6423,N_7461);
nand U11358 (N_11358,N_7233,N_7395);
nand U11359 (N_11359,N_7958,N_7010);
xor U11360 (N_11360,N_7134,N_7792);
xor U11361 (N_11361,N_8714,N_6085);
or U11362 (N_11362,N_6182,N_8686);
nand U11363 (N_11363,N_6753,N_8850);
xnor U11364 (N_11364,N_7302,N_8544);
nor U11365 (N_11365,N_6132,N_8276);
or U11366 (N_11366,N_6770,N_8674);
nor U11367 (N_11367,N_7612,N_6163);
nand U11368 (N_11368,N_7375,N_8801);
nor U11369 (N_11369,N_6451,N_8922);
xnor U11370 (N_11370,N_6996,N_8586);
or U11371 (N_11371,N_8212,N_6250);
and U11372 (N_11372,N_7150,N_8501);
or U11373 (N_11373,N_8995,N_7266);
or U11374 (N_11374,N_6700,N_7383);
or U11375 (N_11375,N_7785,N_6443);
xor U11376 (N_11376,N_8148,N_8917);
and U11377 (N_11377,N_6635,N_8193);
xnor U11378 (N_11378,N_8458,N_7331);
or U11379 (N_11379,N_6241,N_8585);
and U11380 (N_11380,N_7587,N_7784);
or U11381 (N_11381,N_7106,N_7376);
or U11382 (N_11382,N_7679,N_8248);
nor U11383 (N_11383,N_8422,N_8949);
xnor U11384 (N_11384,N_6455,N_7308);
nor U11385 (N_11385,N_7387,N_6390);
xnor U11386 (N_11386,N_7741,N_6522);
nand U11387 (N_11387,N_6620,N_6458);
xor U11388 (N_11388,N_6540,N_8463);
nand U11389 (N_11389,N_6288,N_7243);
nand U11390 (N_11390,N_7792,N_6891);
xnor U11391 (N_11391,N_7696,N_7440);
and U11392 (N_11392,N_6021,N_7131);
xor U11393 (N_11393,N_8033,N_6020);
nor U11394 (N_11394,N_6102,N_8305);
nand U11395 (N_11395,N_6629,N_7565);
or U11396 (N_11396,N_7313,N_7587);
or U11397 (N_11397,N_6754,N_6174);
or U11398 (N_11398,N_6005,N_8788);
xnor U11399 (N_11399,N_6842,N_7125);
nor U11400 (N_11400,N_7103,N_8241);
and U11401 (N_11401,N_6198,N_8857);
nor U11402 (N_11402,N_8044,N_8122);
xnor U11403 (N_11403,N_7918,N_6370);
and U11404 (N_11404,N_8315,N_6131);
nor U11405 (N_11405,N_6138,N_6252);
or U11406 (N_11406,N_8099,N_6660);
or U11407 (N_11407,N_6492,N_8820);
xnor U11408 (N_11408,N_8519,N_6772);
nand U11409 (N_11409,N_8496,N_7446);
nor U11410 (N_11410,N_6944,N_7833);
nor U11411 (N_11411,N_8322,N_6283);
nor U11412 (N_11412,N_7618,N_8854);
and U11413 (N_11413,N_7926,N_6032);
xor U11414 (N_11414,N_7086,N_8645);
nor U11415 (N_11415,N_8483,N_7274);
nor U11416 (N_11416,N_7655,N_7053);
or U11417 (N_11417,N_7456,N_6387);
or U11418 (N_11418,N_6064,N_8104);
or U11419 (N_11419,N_7007,N_6355);
or U11420 (N_11420,N_8243,N_7248);
nand U11421 (N_11421,N_7661,N_8967);
nor U11422 (N_11422,N_6757,N_8614);
nor U11423 (N_11423,N_7978,N_7732);
xnor U11424 (N_11424,N_7275,N_7734);
xor U11425 (N_11425,N_7769,N_8461);
xnor U11426 (N_11426,N_6311,N_8046);
xor U11427 (N_11427,N_7236,N_7462);
nor U11428 (N_11428,N_7264,N_8092);
xor U11429 (N_11429,N_8629,N_8161);
nor U11430 (N_11430,N_8928,N_6394);
xnor U11431 (N_11431,N_7378,N_7109);
xor U11432 (N_11432,N_8528,N_6625);
or U11433 (N_11433,N_8767,N_7143);
nand U11434 (N_11434,N_8122,N_6182);
nor U11435 (N_11435,N_7279,N_8274);
nor U11436 (N_11436,N_6745,N_8870);
or U11437 (N_11437,N_7198,N_8679);
xnor U11438 (N_11438,N_7593,N_6691);
or U11439 (N_11439,N_7338,N_6855);
nand U11440 (N_11440,N_7218,N_7591);
nand U11441 (N_11441,N_7861,N_8805);
nor U11442 (N_11442,N_8086,N_7397);
or U11443 (N_11443,N_7568,N_8495);
or U11444 (N_11444,N_7173,N_7702);
or U11445 (N_11445,N_7306,N_6108);
nand U11446 (N_11446,N_8066,N_8964);
and U11447 (N_11447,N_6404,N_8974);
nand U11448 (N_11448,N_8323,N_6391);
or U11449 (N_11449,N_7267,N_7500);
xor U11450 (N_11450,N_8998,N_7999);
nor U11451 (N_11451,N_7696,N_8204);
nor U11452 (N_11452,N_8420,N_8796);
xnor U11453 (N_11453,N_6849,N_8320);
nand U11454 (N_11454,N_6144,N_7933);
nand U11455 (N_11455,N_6140,N_7911);
nand U11456 (N_11456,N_6021,N_6044);
nor U11457 (N_11457,N_7679,N_6670);
and U11458 (N_11458,N_6437,N_7963);
xnor U11459 (N_11459,N_8124,N_6677);
nor U11460 (N_11460,N_8560,N_7481);
or U11461 (N_11461,N_8818,N_7537);
nor U11462 (N_11462,N_7449,N_8620);
xnor U11463 (N_11463,N_8083,N_6932);
or U11464 (N_11464,N_7010,N_6170);
nand U11465 (N_11465,N_7846,N_7468);
nand U11466 (N_11466,N_6587,N_8606);
and U11467 (N_11467,N_8981,N_7956);
xnor U11468 (N_11468,N_8985,N_6293);
nor U11469 (N_11469,N_8107,N_7354);
and U11470 (N_11470,N_8098,N_8144);
xor U11471 (N_11471,N_8597,N_6353);
xnor U11472 (N_11472,N_6958,N_8621);
or U11473 (N_11473,N_7598,N_6470);
nand U11474 (N_11474,N_8033,N_7873);
and U11475 (N_11475,N_7718,N_8185);
and U11476 (N_11476,N_6085,N_7758);
and U11477 (N_11477,N_7627,N_7301);
xor U11478 (N_11478,N_6503,N_6786);
nor U11479 (N_11479,N_6970,N_7206);
nand U11480 (N_11480,N_8633,N_7216);
or U11481 (N_11481,N_6745,N_8474);
xnor U11482 (N_11482,N_7532,N_6542);
or U11483 (N_11483,N_6716,N_7690);
nor U11484 (N_11484,N_6936,N_7310);
and U11485 (N_11485,N_6009,N_7907);
nor U11486 (N_11486,N_8571,N_8637);
or U11487 (N_11487,N_6699,N_8478);
or U11488 (N_11488,N_8681,N_8782);
and U11489 (N_11489,N_6366,N_6906);
and U11490 (N_11490,N_6085,N_7379);
and U11491 (N_11491,N_6973,N_7041);
xor U11492 (N_11492,N_6514,N_8737);
or U11493 (N_11493,N_7466,N_6671);
or U11494 (N_11494,N_7389,N_7534);
nor U11495 (N_11495,N_8230,N_7639);
xnor U11496 (N_11496,N_6428,N_6368);
nand U11497 (N_11497,N_8495,N_8455);
and U11498 (N_11498,N_6172,N_8382);
and U11499 (N_11499,N_8028,N_8676);
xnor U11500 (N_11500,N_6469,N_8916);
nand U11501 (N_11501,N_7036,N_8037);
and U11502 (N_11502,N_7754,N_6327);
nor U11503 (N_11503,N_8700,N_8933);
nor U11504 (N_11504,N_7580,N_7974);
xor U11505 (N_11505,N_6178,N_8116);
nor U11506 (N_11506,N_7778,N_7270);
and U11507 (N_11507,N_8682,N_6813);
and U11508 (N_11508,N_8669,N_7853);
nor U11509 (N_11509,N_7711,N_6891);
and U11510 (N_11510,N_7609,N_8953);
xnor U11511 (N_11511,N_8268,N_7375);
or U11512 (N_11512,N_8775,N_7806);
nor U11513 (N_11513,N_7284,N_6879);
nor U11514 (N_11514,N_7496,N_7823);
nand U11515 (N_11515,N_8729,N_7770);
nor U11516 (N_11516,N_6039,N_8203);
xor U11517 (N_11517,N_8699,N_6327);
or U11518 (N_11518,N_6591,N_8164);
or U11519 (N_11519,N_8758,N_8321);
xnor U11520 (N_11520,N_7622,N_6703);
nand U11521 (N_11521,N_7164,N_8260);
nor U11522 (N_11522,N_6392,N_6595);
xnor U11523 (N_11523,N_8213,N_7965);
nor U11524 (N_11524,N_8972,N_6892);
xor U11525 (N_11525,N_7401,N_8801);
and U11526 (N_11526,N_8612,N_6475);
or U11527 (N_11527,N_7273,N_7765);
nand U11528 (N_11528,N_7778,N_8079);
or U11529 (N_11529,N_8749,N_6280);
and U11530 (N_11530,N_7049,N_6441);
xnor U11531 (N_11531,N_8549,N_8995);
or U11532 (N_11532,N_8726,N_7480);
or U11533 (N_11533,N_7493,N_6558);
or U11534 (N_11534,N_6861,N_6343);
nor U11535 (N_11535,N_6363,N_8579);
or U11536 (N_11536,N_7214,N_8659);
xor U11537 (N_11537,N_8630,N_8754);
and U11538 (N_11538,N_7101,N_8378);
and U11539 (N_11539,N_8011,N_6923);
nor U11540 (N_11540,N_6130,N_6335);
nand U11541 (N_11541,N_8460,N_8975);
nor U11542 (N_11542,N_6078,N_6629);
xnor U11543 (N_11543,N_8778,N_6087);
xnor U11544 (N_11544,N_6481,N_6180);
nand U11545 (N_11545,N_7298,N_6321);
and U11546 (N_11546,N_7974,N_7796);
nand U11547 (N_11547,N_7899,N_6244);
or U11548 (N_11548,N_8817,N_7644);
and U11549 (N_11549,N_7960,N_7501);
nand U11550 (N_11550,N_6255,N_7405);
nor U11551 (N_11551,N_7355,N_7771);
nand U11552 (N_11552,N_7326,N_7788);
nand U11553 (N_11553,N_6366,N_6837);
nand U11554 (N_11554,N_7702,N_8654);
nor U11555 (N_11555,N_6729,N_6039);
nand U11556 (N_11556,N_7465,N_6513);
and U11557 (N_11557,N_6061,N_8877);
xnor U11558 (N_11558,N_6426,N_7896);
xnor U11559 (N_11559,N_7614,N_7856);
xor U11560 (N_11560,N_8302,N_6300);
and U11561 (N_11561,N_6846,N_6999);
and U11562 (N_11562,N_6121,N_8998);
xnor U11563 (N_11563,N_6927,N_6228);
nand U11564 (N_11564,N_7175,N_6113);
nand U11565 (N_11565,N_7001,N_7814);
nand U11566 (N_11566,N_8379,N_8021);
nor U11567 (N_11567,N_6328,N_7048);
nand U11568 (N_11568,N_7268,N_7024);
nor U11569 (N_11569,N_7413,N_6464);
nand U11570 (N_11570,N_7714,N_7466);
xor U11571 (N_11571,N_7776,N_8737);
or U11572 (N_11572,N_6110,N_6086);
nand U11573 (N_11573,N_8136,N_7321);
xor U11574 (N_11574,N_6619,N_8988);
and U11575 (N_11575,N_7476,N_8746);
nand U11576 (N_11576,N_7086,N_6284);
nor U11577 (N_11577,N_6499,N_7490);
xnor U11578 (N_11578,N_8587,N_7215);
or U11579 (N_11579,N_8733,N_6942);
xnor U11580 (N_11580,N_6988,N_6250);
or U11581 (N_11581,N_6355,N_6687);
and U11582 (N_11582,N_6930,N_7738);
nor U11583 (N_11583,N_8803,N_8684);
nand U11584 (N_11584,N_6872,N_7610);
and U11585 (N_11585,N_6444,N_8920);
or U11586 (N_11586,N_7384,N_8129);
nor U11587 (N_11587,N_8660,N_8568);
nor U11588 (N_11588,N_8670,N_8276);
nor U11589 (N_11589,N_8710,N_8588);
or U11590 (N_11590,N_6738,N_6343);
nand U11591 (N_11591,N_7470,N_7860);
and U11592 (N_11592,N_8084,N_8495);
or U11593 (N_11593,N_7058,N_6319);
or U11594 (N_11594,N_7547,N_7012);
nand U11595 (N_11595,N_8254,N_8221);
or U11596 (N_11596,N_6040,N_8872);
nand U11597 (N_11597,N_8490,N_6136);
nand U11598 (N_11598,N_8350,N_6629);
or U11599 (N_11599,N_6006,N_6237);
nor U11600 (N_11600,N_6932,N_6242);
and U11601 (N_11601,N_7187,N_7799);
xor U11602 (N_11602,N_8163,N_6098);
nor U11603 (N_11603,N_6187,N_7847);
nor U11604 (N_11604,N_6322,N_8701);
xnor U11605 (N_11605,N_8769,N_7621);
xor U11606 (N_11606,N_7760,N_6204);
nor U11607 (N_11607,N_8681,N_8191);
xor U11608 (N_11608,N_7270,N_8287);
nor U11609 (N_11609,N_6038,N_8978);
nor U11610 (N_11610,N_7494,N_8996);
nand U11611 (N_11611,N_8808,N_8414);
and U11612 (N_11612,N_8993,N_7245);
and U11613 (N_11613,N_7603,N_8628);
xor U11614 (N_11614,N_7825,N_6074);
xnor U11615 (N_11615,N_7110,N_6591);
or U11616 (N_11616,N_7394,N_8765);
nor U11617 (N_11617,N_6850,N_7528);
or U11618 (N_11618,N_7671,N_7866);
nand U11619 (N_11619,N_8004,N_7610);
and U11620 (N_11620,N_7328,N_6897);
xnor U11621 (N_11621,N_7394,N_7972);
nand U11622 (N_11622,N_6101,N_6787);
xor U11623 (N_11623,N_8328,N_6237);
xor U11624 (N_11624,N_8178,N_8903);
or U11625 (N_11625,N_7425,N_7114);
xnor U11626 (N_11626,N_7341,N_8240);
nand U11627 (N_11627,N_6423,N_7003);
nand U11628 (N_11628,N_7858,N_8025);
or U11629 (N_11629,N_8360,N_7813);
or U11630 (N_11630,N_6109,N_7567);
nand U11631 (N_11631,N_6956,N_8526);
or U11632 (N_11632,N_7726,N_6219);
or U11633 (N_11633,N_6968,N_7047);
or U11634 (N_11634,N_7006,N_6747);
xor U11635 (N_11635,N_8768,N_7053);
nand U11636 (N_11636,N_8000,N_8882);
nand U11637 (N_11637,N_6974,N_6381);
or U11638 (N_11638,N_7313,N_8156);
nor U11639 (N_11639,N_8017,N_6793);
or U11640 (N_11640,N_8042,N_7386);
xor U11641 (N_11641,N_7966,N_7412);
nor U11642 (N_11642,N_8254,N_6368);
nand U11643 (N_11643,N_7578,N_7867);
nor U11644 (N_11644,N_7894,N_7154);
and U11645 (N_11645,N_7008,N_7055);
nor U11646 (N_11646,N_6933,N_7347);
or U11647 (N_11647,N_8340,N_6783);
xnor U11648 (N_11648,N_8593,N_7937);
nor U11649 (N_11649,N_8898,N_7761);
and U11650 (N_11650,N_8070,N_8383);
or U11651 (N_11651,N_8786,N_8455);
xnor U11652 (N_11652,N_8184,N_7945);
nor U11653 (N_11653,N_8730,N_6507);
xnor U11654 (N_11654,N_7019,N_7286);
or U11655 (N_11655,N_6944,N_7937);
nand U11656 (N_11656,N_6371,N_7065);
and U11657 (N_11657,N_6379,N_6412);
nor U11658 (N_11658,N_6894,N_7935);
nand U11659 (N_11659,N_8096,N_8292);
and U11660 (N_11660,N_8521,N_8134);
or U11661 (N_11661,N_8821,N_7873);
xnor U11662 (N_11662,N_7971,N_6277);
xor U11663 (N_11663,N_6574,N_7688);
and U11664 (N_11664,N_6970,N_8207);
and U11665 (N_11665,N_6406,N_7136);
and U11666 (N_11666,N_7058,N_8905);
nor U11667 (N_11667,N_8351,N_6664);
nor U11668 (N_11668,N_7555,N_7362);
or U11669 (N_11669,N_7901,N_6328);
or U11670 (N_11670,N_6208,N_7993);
nor U11671 (N_11671,N_6741,N_6447);
xnor U11672 (N_11672,N_8176,N_7349);
and U11673 (N_11673,N_6946,N_7900);
or U11674 (N_11674,N_7206,N_8543);
and U11675 (N_11675,N_6677,N_7132);
or U11676 (N_11676,N_8893,N_7274);
xnor U11677 (N_11677,N_8157,N_8076);
or U11678 (N_11678,N_8842,N_8568);
nor U11679 (N_11679,N_8608,N_7052);
or U11680 (N_11680,N_8437,N_7778);
or U11681 (N_11681,N_7576,N_8994);
xor U11682 (N_11682,N_6834,N_8067);
xnor U11683 (N_11683,N_6015,N_6878);
nand U11684 (N_11684,N_6238,N_6705);
xor U11685 (N_11685,N_7713,N_6761);
and U11686 (N_11686,N_6145,N_7259);
or U11687 (N_11687,N_8637,N_6981);
nand U11688 (N_11688,N_6009,N_8984);
and U11689 (N_11689,N_6907,N_7259);
and U11690 (N_11690,N_6609,N_6381);
or U11691 (N_11691,N_8400,N_8527);
and U11692 (N_11692,N_8201,N_7218);
or U11693 (N_11693,N_6150,N_8328);
or U11694 (N_11694,N_8685,N_6875);
nor U11695 (N_11695,N_7732,N_6916);
nor U11696 (N_11696,N_8109,N_7421);
or U11697 (N_11697,N_8228,N_8032);
nor U11698 (N_11698,N_8257,N_7271);
and U11699 (N_11699,N_6392,N_6795);
or U11700 (N_11700,N_7226,N_7177);
and U11701 (N_11701,N_7346,N_7523);
xnor U11702 (N_11702,N_7443,N_6134);
nor U11703 (N_11703,N_7932,N_6661);
xor U11704 (N_11704,N_6979,N_7970);
and U11705 (N_11705,N_8267,N_6230);
nand U11706 (N_11706,N_8168,N_7992);
xnor U11707 (N_11707,N_8490,N_8832);
and U11708 (N_11708,N_8978,N_7205);
or U11709 (N_11709,N_8451,N_8358);
or U11710 (N_11710,N_6038,N_8616);
and U11711 (N_11711,N_7600,N_8575);
and U11712 (N_11712,N_6553,N_8296);
or U11713 (N_11713,N_7759,N_7160);
and U11714 (N_11714,N_6681,N_8375);
xnor U11715 (N_11715,N_6273,N_7458);
nand U11716 (N_11716,N_7990,N_8408);
xnor U11717 (N_11717,N_6546,N_6336);
and U11718 (N_11718,N_7908,N_8560);
or U11719 (N_11719,N_6699,N_6629);
nor U11720 (N_11720,N_7214,N_6156);
nor U11721 (N_11721,N_7990,N_7947);
nand U11722 (N_11722,N_6729,N_6021);
and U11723 (N_11723,N_7587,N_8948);
xor U11724 (N_11724,N_7264,N_7417);
nor U11725 (N_11725,N_8174,N_8912);
nor U11726 (N_11726,N_8833,N_8619);
xnor U11727 (N_11727,N_6902,N_8984);
nor U11728 (N_11728,N_6614,N_8283);
and U11729 (N_11729,N_6214,N_6314);
and U11730 (N_11730,N_8377,N_6236);
xnor U11731 (N_11731,N_7946,N_7306);
xnor U11732 (N_11732,N_8712,N_6578);
nor U11733 (N_11733,N_6131,N_6026);
and U11734 (N_11734,N_8952,N_7129);
xor U11735 (N_11735,N_6433,N_7186);
xor U11736 (N_11736,N_6754,N_6573);
nand U11737 (N_11737,N_7163,N_7719);
or U11738 (N_11738,N_7605,N_8652);
and U11739 (N_11739,N_6263,N_7424);
and U11740 (N_11740,N_6177,N_7382);
nor U11741 (N_11741,N_7951,N_7329);
nor U11742 (N_11742,N_8734,N_7549);
xor U11743 (N_11743,N_8164,N_6242);
xor U11744 (N_11744,N_7220,N_6909);
nor U11745 (N_11745,N_7362,N_8779);
or U11746 (N_11746,N_6593,N_8271);
nor U11747 (N_11747,N_8396,N_8139);
or U11748 (N_11748,N_8717,N_8090);
or U11749 (N_11749,N_8805,N_8631);
nand U11750 (N_11750,N_7682,N_8663);
and U11751 (N_11751,N_8296,N_8916);
xnor U11752 (N_11752,N_6435,N_8734);
or U11753 (N_11753,N_7977,N_6798);
xor U11754 (N_11754,N_7246,N_8852);
or U11755 (N_11755,N_8882,N_6000);
or U11756 (N_11756,N_8105,N_8098);
nand U11757 (N_11757,N_6283,N_6435);
nor U11758 (N_11758,N_6415,N_6472);
nand U11759 (N_11759,N_8866,N_6759);
nand U11760 (N_11760,N_6071,N_8321);
or U11761 (N_11761,N_7062,N_8462);
nand U11762 (N_11762,N_8893,N_8194);
nand U11763 (N_11763,N_6623,N_8656);
nand U11764 (N_11764,N_6633,N_6626);
and U11765 (N_11765,N_8900,N_7383);
xor U11766 (N_11766,N_6085,N_8110);
or U11767 (N_11767,N_7701,N_8489);
or U11768 (N_11768,N_6367,N_8358);
nand U11769 (N_11769,N_7523,N_8173);
and U11770 (N_11770,N_8387,N_6809);
nand U11771 (N_11771,N_8680,N_6745);
nand U11772 (N_11772,N_7832,N_6403);
xnor U11773 (N_11773,N_6242,N_7507);
or U11774 (N_11774,N_8163,N_8149);
nand U11775 (N_11775,N_7137,N_8609);
xor U11776 (N_11776,N_8924,N_6594);
nor U11777 (N_11777,N_6048,N_8452);
or U11778 (N_11778,N_8594,N_7930);
nand U11779 (N_11779,N_6689,N_6091);
xnor U11780 (N_11780,N_7751,N_8112);
and U11781 (N_11781,N_8651,N_6964);
or U11782 (N_11782,N_7633,N_6662);
or U11783 (N_11783,N_7958,N_8370);
nor U11784 (N_11784,N_6065,N_8781);
nor U11785 (N_11785,N_8918,N_6379);
xor U11786 (N_11786,N_7080,N_7040);
nand U11787 (N_11787,N_8643,N_8673);
and U11788 (N_11788,N_6158,N_8099);
nand U11789 (N_11789,N_7211,N_8490);
nor U11790 (N_11790,N_8970,N_7738);
or U11791 (N_11791,N_8256,N_8356);
nand U11792 (N_11792,N_6841,N_7506);
xnor U11793 (N_11793,N_6908,N_6511);
nand U11794 (N_11794,N_6622,N_7230);
nand U11795 (N_11795,N_7913,N_6866);
or U11796 (N_11796,N_6354,N_6721);
or U11797 (N_11797,N_8311,N_8082);
and U11798 (N_11798,N_8708,N_6133);
nor U11799 (N_11799,N_7645,N_6890);
xnor U11800 (N_11800,N_8309,N_7627);
and U11801 (N_11801,N_6488,N_7464);
nor U11802 (N_11802,N_6772,N_8511);
xnor U11803 (N_11803,N_8036,N_8644);
or U11804 (N_11804,N_6809,N_6194);
and U11805 (N_11805,N_7326,N_6054);
nand U11806 (N_11806,N_8727,N_7084);
nand U11807 (N_11807,N_8195,N_8295);
or U11808 (N_11808,N_8705,N_6621);
and U11809 (N_11809,N_6277,N_7414);
and U11810 (N_11810,N_6988,N_6892);
or U11811 (N_11811,N_8802,N_7096);
xor U11812 (N_11812,N_7743,N_7860);
nand U11813 (N_11813,N_7567,N_8895);
nor U11814 (N_11814,N_8448,N_6329);
and U11815 (N_11815,N_8462,N_6794);
xor U11816 (N_11816,N_8391,N_8788);
nor U11817 (N_11817,N_7705,N_6037);
nor U11818 (N_11818,N_7861,N_7854);
xnor U11819 (N_11819,N_7559,N_7972);
nand U11820 (N_11820,N_7445,N_6757);
or U11821 (N_11821,N_7012,N_8014);
and U11822 (N_11822,N_8395,N_6507);
and U11823 (N_11823,N_8161,N_7730);
nand U11824 (N_11824,N_8500,N_8221);
xor U11825 (N_11825,N_7273,N_6122);
nand U11826 (N_11826,N_8109,N_7332);
nor U11827 (N_11827,N_6504,N_8177);
nand U11828 (N_11828,N_7681,N_6231);
nor U11829 (N_11829,N_8232,N_8303);
xnor U11830 (N_11830,N_7553,N_8473);
and U11831 (N_11831,N_6542,N_6107);
nor U11832 (N_11832,N_7615,N_6100);
xnor U11833 (N_11833,N_7651,N_8030);
and U11834 (N_11834,N_8617,N_8635);
nor U11835 (N_11835,N_6128,N_7619);
or U11836 (N_11836,N_6496,N_7353);
nor U11837 (N_11837,N_6461,N_8532);
nand U11838 (N_11838,N_7137,N_7450);
xnor U11839 (N_11839,N_6065,N_6134);
and U11840 (N_11840,N_8033,N_8640);
nor U11841 (N_11841,N_7370,N_7457);
xor U11842 (N_11842,N_7258,N_7460);
and U11843 (N_11843,N_8525,N_7523);
and U11844 (N_11844,N_7727,N_6898);
xnor U11845 (N_11845,N_7957,N_6881);
nand U11846 (N_11846,N_8663,N_7368);
and U11847 (N_11847,N_7167,N_7625);
nand U11848 (N_11848,N_8627,N_7367);
nor U11849 (N_11849,N_8542,N_7941);
and U11850 (N_11850,N_6700,N_6842);
nand U11851 (N_11851,N_8203,N_6982);
xnor U11852 (N_11852,N_6005,N_8219);
and U11853 (N_11853,N_6416,N_6620);
nor U11854 (N_11854,N_6869,N_7570);
nand U11855 (N_11855,N_7637,N_8296);
nor U11856 (N_11856,N_6998,N_8560);
and U11857 (N_11857,N_8464,N_7261);
xor U11858 (N_11858,N_7653,N_7807);
nor U11859 (N_11859,N_7627,N_8211);
nand U11860 (N_11860,N_7187,N_7340);
nor U11861 (N_11861,N_8656,N_8892);
or U11862 (N_11862,N_6977,N_8681);
and U11863 (N_11863,N_8301,N_8036);
and U11864 (N_11864,N_7144,N_8758);
nand U11865 (N_11865,N_8859,N_8963);
and U11866 (N_11866,N_6770,N_8027);
nand U11867 (N_11867,N_7482,N_6965);
nor U11868 (N_11868,N_6622,N_6406);
and U11869 (N_11869,N_8168,N_8740);
nand U11870 (N_11870,N_7872,N_6303);
xnor U11871 (N_11871,N_8058,N_6266);
and U11872 (N_11872,N_7544,N_8493);
and U11873 (N_11873,N_7907,N_7857);
nor U11874 (N_11874,N_8138,N_6923);
nor U11875 (N_11875,N_8711,N_8194);
and U11876 (N_11876,N_7115,N_6104);
xnor U11877 (N_11877,N_7415,N_7225);
nand U11878 (N_11878,N_7796,N_8207);
nand U11879 (N_11879,N_8177,N_7326);
and U11880 (N_11880,N_7665,N_6389);
xnor U11881 (N_11881,N_8573,N_6869);
xor U11882 (N_11882,N_6836,N_7651);
nor U11883 (N_11883,N_7619,N_8969);
nor U11884 (N_11884,N_8132,N_8951);
xor U11885 (N_11885,N_6478,N_7754);
nor U11886 (N_11886,N_8372,N_6905);
nor U11887 (N_11887,N_8256,N_7038);
nor U11888 (N_11888,N_8447,N_8550);
or U11889 (N_11889,N_7899,N_7708);
nand U11890 (N_11890,N_8057,N_7880);
xor U11891 (N_11891,N_7337,N_6840);
nand U11892 (N_11892,N_8356,N_8669);
or U11893 (N_11893,N_8362,N_6988);
and U11894 (N_11894,N_7338,N_6184);
nor U11895 (N_11895,N_6994,N_7231);
or U11896 (N_11896,N_7195,N_8713);
xor U11897 (N_11897,N_7024,N_6915);
and U11898 (N_11898,N_6757,N_8450);
and U11899 (N_11899,N_7635,N_6821);
nand U11900 (N_11900,N_8288,N_6584);
nand U11901 (N_11901,N_8990,N_6380);
xnor U11902 (N_11902,N_7428,N_8114);
xor U11903 (N_11903,N_7734,N_7892);
nand U11904 (N_11904,N_8373,N_8798);
or U11905 (N_11905,N_6719,N_6068);
or U11906 (N_11906,N_8040,N_6269);
xnor U11907 (N_11907,N_7028,N_8358);
nor U11908 (N_11908,N_6663,N_6337);
xor U11909 (N_11909,N_8096,N_7008);
or U11910 (N_11910,N_8574,N_6731);
xor U11911 (N_11911,N_7779,N_8926);
nor U11912 (N_11912,N_6110,N_6890);
and U11913 (N_11913,N_7590,N_6378);
and U11914 (N_11914,N_8210,N_7379);
nor U11915 (N_11915,N_6409,N_8792);
nand U11916 (N_11916,N_8589,N_7176);
or U11917 (N_11917,N_7835,N_7382);
nand U11918 (N_11918,N_6157,N_6631);
nand U11919 (N_11919,N_8208,N_7024);
or U11920 (N_11920,N_6286,N_8695);
or U11921 (N_11921,N_6692,N_7251);
xor U11922 (N_11922,N_7716,N_6875);
and U11923 (N_11923,N_6938,N_8632);
and U11924 (N_11924,N_8192,N_8884);
xnor U11925 (N_11925,N_6708,N_8770);
nor U11926 (N_11926,N_6827,N_7815);
nand U11927 (N_11927,N_8623,N_8776);
xnor U11928 (N_11928,N_8063,N_7246);
xnor U11929 (N_11929,N_7535,N_8053);
nor U11930 (N_11930,N_6775,N_8454);
or U11931 (N_11931,N_7069,N_6764);
xnor U11932 (N_11932,N_8433,N_8654);
nor U11933 (N_11933,N_8592,N_8040);
nor U11934 (N_11934,N_7761,N_6626);
nand U11935 (N_11935,N_6681,N_6016);
and U11936 (N_11936,N_6838,N_6638);
and U11937 (N_11937,N_7867,N_8386);
or U11938 (N_11938,N_6750,N_8813);
nand U11939 (N_11939,N_6083,N_8916);
xnor U11940 (N_11940,N_6547,N_7566);
and U11941 (N_11941,N_7796,N_8557);
nor U11942 (N_11942,N_6172,N_7791);
or U11943 (N_11943,N_7462,N_7042);
or U11944 (N_11944,N_7543,N_6105);
and U11945 (N_11945,N_7857,N_7625);
nand U11946 (N_11946,N_7431,N_8566);
nor U11947 (N_11947,N_6988,N_7108);
xor U11948 (N_11948,N_7699,N_7703);
nand U11949 (N_11949,N_7187,N_7074);
nand U11950 (N_11950,N_7243,N_7100);
nand U11951 (N_11951,N_6595,N_8266);
nand U11952 (N_11952,N_7946,N_7772);
and U11953 (N_11953,N_8986,N_6854);
nor U11954 (N_11954,N_8032,N_7805);
and U11955 (N_11955,N_8662,N_7122);
or U11956 (N_11956,N_6670,N_6904);
nand U11957 (N_11957,N_8171,N_7437);
nand U11958 (N_11958,N_8962,N_7768);
and U11959 (N_11959,N_6120,N_7973);
and U11960 (N_11960,N_6344,N_8277);
nand U11961 (N_11961,N_8499,N_7312);
nor U11962 (N_11962,N_6988,N_8996);
nand U11963 (N_11963,N_8410,N_6155);
or U11964 (N_11964,N_6302,N_7748);
and U11965 (N_11965,N_7129,N_8962);
or U11966 (N_11966,N_6274,N_8205);
or U11967 (N_11967,N_6279,N_6798);
or U11968 (N_11968,N_8194,N_7609);
nor U11969 (N_11969,N_6879,N_7241);
nand U11970 (N_11970,N_6801,N_6747);
or U11971 (N_11971,N_7526,N_6091);
and U11972 (N_11972,N_7202,N_6436);
nor U11973 (N_11973,N_7825,N_8516);
nor U11974 (N_11974,N_6426,N_8538);
and U11975 (N_11975,N_6606,N_7911);
and U11976 (N_11976,N_7896,N_6726);
nor U11977 (N_11977,N_8280,N_7643);
nor U11978 (N_11978,N_6829,N_6497);
nand U11979 (N_11979,N_7984,N_8462);
nor U11980 (N_11980,N_8850,N_8904);
and U11981 (N_11981,N_8430,N_7866);
nand U11982 (N_11982,N_6155,N_8041);
and U11983 (N_11983,N_6451,N_6953);
nor U11984 (N_11984,N_7514,N_7557);
and U11985 (N_11985,N_6288,N_7209);
and U11986 (N_11986,N_6733,N_7250);
and U11987 (N_11987,N_7476,N_7020);
and U11988 (N_11988,N_8672,N_6582);
or U11989 (N_11989,N_7581,N_8009);
nor U11990 (N_11990,N_8897,N_7803);
nor U11991 (N_11991,N_8927,N_6870);
or U11992 (N_11992,N_7532,N_6773);
nand U11993 (N_11993,N_8092,N_6706);
and U11994 (N_11994,N_6200,N_7131);
or U11995 (N_11995,N_6445,N_6243);
nor U11996 (N_11996,N_6224,N_8737);
nor U11997 (N_11997,N_8413,N_7017);
or U11998 (N_11998,N_8789,N_8119);
nand U11999 (N_11999,N_8111,N_6977);
nor U12000 (N_12000,N_11249,N_9709);
nor U12001 (N_12001,N_11586,N_9918);
nand U12002 (N_12002,N_9271,N_9064);
nand U12003 (N_12003,N_9603,N_11217);
or U12004 (N_12004,N_9058,N_11908);
xor U12005 (N_12005,N_10919,N_10504);
and U12006 (N_12006,N_10732,N_10337);
and U12007 (N_12007,N_11871,N_10891);
and U12008 (N_12008,N_10438,N_11110);
or U12009 (N_12009,N_9996,N_9289);
and U12010 (N_12010,N_9193,N_10882);
nand U12011 (N_12011,N_10635,N_11456);
nand U12012 (N_12012,N_9383,N_11530);
and U12013 (N_12013,N_11402,N_10658);
and U12014 (N_12014,N_10350,N_9067);
nor U12015 (N_12015,N_9148,N_11481);
or U12016 (N_12016,N_11968,N_10075);
nor U12017 (N_12017,N_10111,N_11044);
or U12018 (N_12018,N_9890,N_10482);
or U12019 (N_12019,N_10580,N_11882);
nand U12020 (N_12020,N_11264,N_9290);
nor U12021 (N_12021,N_10016,N_10720);
nand U12022 (N_12022,N_9763,N_9524);
xor U12023 (N_12023,N_9873,N_11146);
nor U12024 (N_12024,N_10553,N_10103);
nand U12025 (N_12025,N_10941,N_11250);
or U12026 (N_12026,N_10446,N_9886);
nor U12027 (N_12027,N_11702,N_10511);
and U12028 (N_12028,N_11141,N_9306);
nand U12029 (N_12029,N_11698,N_11738);
nor U12030 (N_12030,N_9874,N_10273);
nor U12031 (N_12031,N_9136,N_11444);
xnor U12032 (N_12032,N_11502,N_9002);
nor U12033 (N_12033,N_10462,N_10765);
or U12034 (N_12034,N_10122,N_9831);
or U12035 (N_12035,N_10409,N_10233);
nor U12036 (N_12036,N_9680,N_10678);
nor U12037 (N_12037,N_9182,N_11842);
nand U12038 (N_12038,N_11732,N_11520);
nand U12039 (N_12039,N_11446,N_9662);
or U12040 (N_12040,N_11621,N_10017);
xnor U12041 (N_12041,N_9055,N_11457);
nand U12042 (N_12042,N_11346,N_10519);
nor U12043 (N_12043,N_9702,N_10386);
nand U12044 (N_12044,N_11636,N_9165);
nor U12045 (N_12045,N_11877,N_10486);
or U12046 (N_12046,N_11454,N_11432);
xnor U12047 (N_12047,N_10844,N_10742);
nand U12048 (N_12048,N_10674,N_9957);
or U12049 (N_12049,N_11978,N_9794);
nand U12050 (N_12050,N_9034,N_11800);
nand U12051 (N_12051,N_10625,N_11229);
xor U12052 (N_12052,N_9587,N_9492);
xor U12053 (N_12053,N_11209,N_9677);
nand U12054 (N_12054,N_10505,N_10025);
xor U12055 (N_12055,N_9618,N_9628);
or U12056 (N_12056,N_10594,N_9589);
and U12057 (N_12057,N_10402,N_11259);
or U12058 (N_12058,N_9829,N_9561);
xor U12059 (N_12059,N_10334,N_9334);
nand U12060 (N_12060,N_10634,N_10556);
nor U12061 (N_12061,N_11508,N_11135);
or U12062 (N_12062,N_9443,N_11964);
nand U12063 (N_12063,N_9040,N_9620);
nand U12064 (N_12064,N_9440,N_9775);
nand U12065 (N_12065,N_9951,N_9705);
nand U12066 (N_12066,N_9954,N_11742);
or U12067 (N_12067,N_11565,N_10176);
or U12068 (N_12068,N_10593,N_9904);
nor U12069 (N_12069,N_9204,N_11900);
xnor U12070 (N_12070,N_10125,N_9211);
xnor U12071 (N_12071,N_9177,N_10567);
and U12072 (N_12072,N_9922,N_9739);
or U12073 (N_12073,N_9173,N_9156);
or U12074 (N_12074,N_11707,N_9310);
xnor U12075 (N_12075,N_11946,N_10682);
or U12076 (N_12076,N_10857,N_10066);
nor U12077 (N_12077,N_10053,N_11218);
or U12078 (N_12078,N_11181,N_10885);
and U12079 (N_12079,N_10824,N_9188);
and U12080 (N_12080,N_9862,N_9968);
nand U12081 (N_12081,N_10947,N_10317);
nor U12082 (N_12082,N_11306,N_11696);
xnor U12083 (N_12083,N_10225,N_9244);
or U12084 (N_12084,N_10179,N_10121);
and U12085 (N_12085,N_10734,N_9694);
and U12086 (N_12086,N_11921,N_11932);
xnor U12087 (N_12087,N_10725,N_9641);
xnor U12088 (N_12088,N_11241,N_11781);
or U12089 (N_12089,N_11518,N_9949);
nand U12090 (N_12090,N_10785,N_10791);
and U12091 (N_12091,N_11342,N_10305);
xnor U12092 (N_12092,N_9964,N_10663);
nand U12093 (N_12093,N_10360,N_11896);
and U12094 (N_12094,N_10114,N_11130);
xnor U12095 (N_12095,N_11156,N_10089);
nor U12096 (N_12096,N_10326,N_10733);
nor U12097 (N_12097,N_9434,N_11279);
nor U12098 (N_12098,N_10236,N_9593);
and U12099 (N_12099,N_11246,N_11780);
or U12100 (N_12100,N_9656,N_11776);
nand U12101 (N_12101,N_10840,N_10227);
nand U12102 (N_12102,N_9378,N_10633);
or U12103 (N_12103,N_11950,N_9909);
xor U12104 (N_12104,N_11855,N_11026);
nand U12105 (N_12105,N_10019,N_10557);
or U12106 (N_12106,N_10000,N_11100);
or U12107 (N_12107,N_9444,N_11362);
xor U12108 (N_12108,N_9780,N_11202);
or U12109 (N_12109,N_9217,N_10145);
or U12110 (N_12110,N_10893,N_11195);
nor U12111 (N_12111,N_10601,N_9130);
or U12112 (N_12112,N_10563,N_11323);
and U12113 (N_12113,N_10714,N_11343);
and U12114 (N_12114,N_11622,N_10414);
or U12115 (N_12115,N_11392,N_9133);
and U12116 (N_12116,N_9572,N_11017);
and U12117 (N_12117,N_11359,N_10549);
nor U12118 (N_12118,N_9191,N_11336);
or U12119 (N_12119,N_9733,N_11715);
nand U12120 (N_12120,N_10578,N_10669);
nand U12121 (N_12121,N_11262,N_11277);
or U12122 (N_12122,N_11869,N_9888);
nand U12123 (N_12123,N_10993,N_11762);
nand U12124 (N_12124,N_10029,N_11626);
nor U12125 (N_12125,N_11765,N_11079);
and U12126 (N_12126,N_9205,N_9273);
xnor U12127 (N_12127,N_10907,N_9554);
nor U12128 (N_12128,N_11095,N_9270);
or U12129 (N_12129,N_11210,N_11351);
nand U12130 (N_12130,N_9458,N_10131);
nor U12131 (N_12131,N_10464,N_9030);
or U12132 (N_12132,N_11007,N_11575);
and U12133 (N_12133,N_10716,N_10629);
or U12134 (N_12134,N_10271,N_9973);
nor U12135 (N_12135,N_11741,N_10169);
nand U12136 (N_12136,N_10499,N_9465);
xnor U12137 (N_12137,N_9144,N_11648);
xnor U12138 (N_12138,N_11623,N_11013);
or U12139 (N_12139,N_9539,N_10289);
nand U12140 (N_12140,N_11745,N_10985);
nor U12141 (N_12141,N_9377,N_10748);
and U12142 (N_12142,N_9274,N_10073);
nand U12143 (N_12143,N_11730,N_10659);
nand U12144 (N_12144,N_10437,N_10344);
or U12145 (N_12145,N_11397,N_10055);
and U12146 (N_12146,N_10672,N_10755);
and U12147 (N_12147,N_10341,N_11535);
and U12148 (N_12148,N_9102,N_11970);
nor U12149 (N_12149,N_10932,N_9602);
or U12150 (N_12150,N_9720,N_10666);
nand U12151 (N_12151,N_11977,N_9337);
xnor U12152 (N_12152,N_11638,N_10304);
or U12153 (N_12153,N_10485,N_9189);
xnor U12154 (N_12154,N_11695,N_10704);
nor U12155 (N_12155,N_11317,N_10280);
and U12156 (N_12156,N_11038,N_11265);
xor U12157 (N_12157,N_11806,N_9734);
xnor U12158 (N_12158,N_11352,N_11451);
and U12159 (N_12159,N_9810,N_9540);
or U12160 (N_12160,N_10298,N_10895);
nor U12161 (N_12161,N_11930,N_11369);
xnor U12162 (N_12162,N_11546,N_10761);
or U12163 (N_12163,N_9974,N_10497);
or U12164 (N_12164,N_11687,N_9152);
and U12165 (N_12165,N_9422,N_10194);
nand U12166 (N_12166,N_11204,N_11650);
and U12167 (N_12167,N_9318,N_9575);
nor U12168 (N_12168,N_10347,N_9804);
nor U12169 (N_12169,N_9562,N_9476);
xor U12170 (N_12170,N_9786,N_10590);
nor U12171 (N_12171,N_10309,N_9057);
and U12172 (N_12172,N_11054,N_10065);
xnor U12173 (N_12173,N_10364,N_9342);
and U12174 (N_12174,N_9495,N_11180);
and U12175 (N_12175,N_11627,N_10938);
or U12176 (N_12176,N_9781,N_9472);
and U12177 (N_12177,N_11425,N_10810);
nor U12178 (N_12178,N_9293,N_9517);
xor U12179 (N_12179,N_10996,N_10458);
or U12180 (N_12180,N_11881,N_11541);
and U12181 (N_12181,N_11281,N_9945);
or U12182 (N_12182,N_9218,N_11398);
nand U12183 (N_12183,N_9544,N_10604);
and U12184 (N_12184,N_9162,N_11886);
or U12185 (N_12185,N_9045,N_11302);
nor U12186 (N_12186,N_10232,N_11992);
nor U12187 (N_12187,N_11669,N_9570);
nor U12188 (N_12188,N_10400,N_9410);
xnor U12189 (N_12189,N_9256,N_10788);
or U12190 (N_12190,N_11588,N_11803);
xnor U12191 (N_12191,N_10287,N_9283);
and U12192 (N_12192,N_10603,N_11072);
and U12193 (N_12193,N_10877,N_9339);
nor U12194 (N_12194,N_9860,N_11314);
xnor U12195 (N_12195,N_10118,N_10838);
and U12196 (N_12196,N_9678,N_10512);
or U12197 (N_12197,N_9326,N_10849);
and U12198 (N_12198,N_10258,N_9092);
nor U12199 (N_12199,N_9948,N_10835);
nor U12200 (N_12200,N_10863,N_9843);
and U12201 (N_12201,N_9574,N_10676);
or U12202 (N_12202,N_11163,N_11274);
or U12203 (N_12203,N_9632,N_10268);
xnor U12204 (N_12204,N_10170,N_9013);
nand U12205 (N_12205,N_11601,N_9275);
and U12206 (N_12206,N_9473,N_9880);
nor U12207 (N_12207,N_9297,N_9559);
and U12208 (N_12208,N_9053,N_9239);
nand U12209 (N_12209,N_11419,N_10244);
and U12210 (N_12210,N_9496,N_11985);
and U12211 (N_12211,N_10128,N_11216);
nand U12212 (N_12212,N_11923,N_10712);
or U12213 (N_12213,N_9898,N_11207);
nor U12214 (N_12214,N_11168,N_9891);
nor U12215 (N_12215,N_11562,N_11147);
nand U12216 (N_12216,N_10048,N_10101);
xor U12217 (N_12217,N_10952,N_10319);
xor U12218 (N_12218,N_9069,N_10508);
xnor U12219 (N_12219,N_9851,N_11828);
or U12220 (N_12220,N_9346,N_9199);
xor U12221 (N_12221,N_9819,N_9418);
nand U12222 (N_12222,N_10410,N_10311);
or U12223 (N_12223,N_11603,N_11925);
nor U12224 (N_12224,N_11850,N_9697);
or U12225 (N_12225,N_9625,N_10834);
and U12226 (N_12226,N_11248,N_10096);
nor U12227 (N_12227,N_9645,N_9363);
and U12228 (N_12228,N_10132,N_11651);
nand U12229 (N_12229,N_9097,N_9784);
nor U12230 (N_12230,N_10760,N_10677);
and U12231 (N_12231,N_10861,N_11372);
or U12232 (N_12232,N_11475,N_10622);
nand U12233 (N_12233,N_11152,N_10694);
nor U12234 (N_12234,N_11555,N_10027);
xnor U12235 (N_12235,N_11827,N_9646);
xnor U12236 (N_12236,N_9348,N_10046);
and U12237 (N_12237,N_11931,N_11361);
nor U12238 (N_12238,N_11866,N_9266);
nand U12239 (N_12239,N_11185,N_9160);
and U12240 (N_12240,N_11324,N_9281);
nor U12241 (N_12241,N_11734,N_10898);
and U12242 (N_12242,N_11678,N_10193);
xnor U12243 (N_12243,N_11176,N_9050);
or U12244 (N_12244,N_11581,N_11247);
nand U12245 (N_12245,N_9450,N_9416);
nand U12246 (N_12246,N_11461,N_10463);
nand U12247 (N_12247,N_11383,N_11727);
nand U12248 (N_12248,N_10671,N_10422);
and U12249 (N_12249,N_10968,N_9036);
and U12250 (N_12250,N_11006,N_9665);
nand U12251 (N_12251,N_10889,N_9600);
nor U12252 (N_12252,N_9436,N_11106);
nor U12253 (N_12253,N_11655,N_10159);
and U12254 (N_12254,N_11551,N_9965);
nor U12255 (N_12255,N_10291,N_10809);
or U12256 (N_12256,N_10220,N_9877);
nor U12257 (N_12257,N_9247,N_10180);
nand U12258 (N_12258,N_10967,N_11466);
nand U12259 (N_12259,N_10026,N_11310);
or U12260 (N_12260,N_9820,N_11945);
xnor U12261 (N_12261,N_9866,N_10452);
or U12262 (N_12262,N_10476,N_10215);
and U12263 (N_12263,N_10272,N_11459);
xnor U12264 (N_12264,N_10007,N_9333);
and U12265 (N_12265,N_11979,N_11613);
nor U12266 (N_12266,N_10130,N_9487);
and U12267 (N_12267,N_10398,N_9532);
xnor U12268 (N_12268,N_11971,N_11020);
or U12269 (N_12269,N_11365,N_10698);
nor U12270 (N_12270,N_11848,N_9608);
and U12271 (N_12271,N_9300,N_10701);
nor U12272 (N_12272,N_11086,N_10149);
and U12273 (N_12273,N_11775,N_11339);
nor U12274 (N_12274,N_9841,N_9456);
nand U12275 (N_12275,N_9549,N_9717);
xor U12276 (N_12276,N_11831,N_10082);
or U12277 (N_12277,N_9533,N_9176);
nand U12278 (N_12278,N_9746,N_10987);
nor U12279 (N_12279,N_10752,N_9966);
xnor U12280 (N_12280,N_11068,N_10837);
and U12281 (N_12281,N_10173,N_11774);
xor U12282 (N_12282,N_11538,N_10379);
or U12283 (N_12283,N_11462,N_9061);
xor U12284 (N_12284,N_10113,N_9718);
or U12285 (N_12285,N_9923,N_9028);
nand U12286 (N_12286,N_11426,N_9134);
nand U12287 (N_12287,N_11667,N_11993);
and U12288 (N_12288,N_11942,N_10296);
nand U12289 (N_12289,N_10391,N_10241);
or U12290 (N_12290,N_9338,N_11969);
or U12291 (N_12291,N_10481,N_11286);
and U12292 (N_12292,N_11566,N_10831);
and U12293 (N_12293,N_11818,N_11153);
or U12294 (N_12294,N_11944,N_11697);
nor U12295 (N_12295,N_10406,N_9399);
nor U12296 (N_12296,N_10421,N_9384);
and U12297 (N_12297,N_10306,N_11884);
nor U12298 (N_12298,N_10295,N_10697);
and U12299 (N_12299,N_11252,N_11620);
nand U12300 (N_12300,N_9634,N_9785);
xor U12301 (N_12301,N_11256,N_11761);
or U12302 (N_12302,N_11037,N_9833);
nor U12303 (N_12303,N_10252,N_9824);
and U12304 (N_12304,N_11858,N_9301);
and U12305 (N_12305,N_10670,N_11770);
xnor U12306 (N_12306,N_10913,N_11901);
xnor U12307 (N_12307,N_10571,N_9195);
and U12308 (N_12308,N_10617,N_10267);
nor U12309 (N_12309,N_10349,N_11878);
or U12310 (N_12310,N_10804,N_10407);
and U12311 (N_12311,N_9741,N_9499);
and U12312 (N_12312,N_9027,N_10690);
and U12313 (N_12313,N_9683,N_11064);
nand U12314 (N_12314,N_10702,N_9375);
nor U12315 (N_12315,N_11568,N_11201);
nand U12316 (N_12316,N_9942,N_10195);
and U12317 (N_12317,N_11769,N_10535);
xnor U12318 (N_12318,N_11673,N_9770);
and U12319 (N_12319,N_10023,N_11830);
nor U12320 (N_12320,N_10187,N_9609);
or U12321 (N_12321,N_11231,N_11238);
and U12322 (N_12322,N_11737,N_9558);
nand U12323 (N_12323,N_10956,N_9779);
or U12324 (N_12324,N_9196,N_9861);
or U12325 (N_12325,N_11554,N_9541);
nand U12326 (N_12326,N_9569,N_9868);
nor U12327 (N_12327,N_9743,N_11124);
and U12328 (N_12328,N_11128,N_9967);
nor U12329 (N_12329,N_10240,N_10492);
nand U12330 (N_12330,N_11609,N_9240);
xnor U12331 (N_12331,N_10847,N_10049);
and U12332 (N_12332,N_9463,N_10077);
xnor U12333 (N_12333,N_11799,N_11998);
xor U12334 (N_12334,N_10954,N_9395);
nand U12335 (N_12335,N_9415,N_10653);
or U12336 (N_12336,N_11718,N_9579);
nor U12337 (N_12337,N_9936,N_10906);
xor U12338 (N_12338,N_10598,N_11088);
nand U12339 (N_12339,N_10275,N_10152);
nand U12340 (N_12340,N_9721,N_10450);
or U12341 (N_12341,N_9917,N_11332);
xnor U12342 (N_12342,N_10052,N_9071);
nor U12343 (N_12343,N_10183,N_10028);
or U12344 (N_12344,N_11497,N_10106);
xnor U12345 (N_12345,N_10691,N_10070);
nand U12346 (N_12346,N_9538,N_9699);
nand U12347 (N_12347,N_9494,N_10502);
xnor U12348 (N_12348,N_10636,N_9844);
or U12349 (N_12349,N_10314,N_11364);
or U12350 (N_12350,N_10420,N_10825);
or U12351 (N_12351,N_11236,N_10681);
and U12352 (N_12352,N_11504,N_11463);
nor U12353 (N_12353,N_9818,N_10856);
or U12354 (N_12354,N_11579,N_9285);
nor U12355 (N_12355,N_11490,N_10966);
nand U12356 (N_12356,N_11187,N_9186);
nand U12357 (N_12357,N_11990,N_11863);
or U12358 (N_12358,N_10310,N_11164);
xor U12359 (N_12359,N_10044,N_9754);
nor U12360 (N_12360,N_10978,N_9952);
nor U12361 (N_12361,N_10336,N_10591);
or U12362 (N_12362,N_10894,N_11967);
nand U12363 (N_12363,N_11282,N_9567);
nand U12364 (N_12364,N_11870,N_10221);
nand U12365 (N_12365,N_10097,N_11237);
and U12366 (N_12366,N_10444,N_10262);
nor U12367 (N_12367,N_10403,N_9714);
or U12368 (N_12368,N_11529,N_9518);
nor U12369 (N_12369,N_11213,N_11108);
xor U12370 (N_12370,N_9481,N_11689);
nor U12371 (N_12371,N_9352,N_9666);
nand U12372 (N_12372,N_10724,N_10875);
and U12373 (N_12373,N_11292,N_11948);
xnor U12374 (N_12374,N_11919,N_11471);
nand U12375 (N_12375,N_9316,N_11654);
nand U12376 (N_12376,N_10864,N_11391);
and U12377 (N_12377,N_9219,N_10214);
nor U12378 (N_12378,N_10265,N_10014);
nand U12379 (N_12379,N_9582,N_10270);
nand U12380 (N_12380,N_9612,N_9099);
or U12381 (N_12381,N_11356,N_11078);
xnor U12382 (N_12382,N_11101,N_11251);
or U12383 (N_12383,N_9519,N_11066);
xor U12384 (N_12384,N_9288,N_11127);
xnor U12385 (N_12385,N_10886,N_10279);
or U12386 (N_12386,N_10550,N_9286);
or U12387 (N_12387,N_10308,N_9046);
xnor U12388 (N_12388,N_10248,N_9469);
xor U12389 (N_12389,N_9427,N_9224);
nor U12390 (N_12390,N_9510,N_9525);
or U12391 (N_12391,N_9428,N_9054);
nand U12392 (N_12392,N_10608,N_10127);
and U12393 (N_12393,N_11709,N_9950);
xnor U12394 (N_12394,N_10828,N_10143);
nor U12395 (N_12395,N_10425,N_9413);
or U12396 (N_12396,N_10362,N_9406);
or U12397 (N_12397,N_11417,N_10107);
nand U12398 (N_12398,N_11658,N_10646);
xor U12399 (N_12399,N_11531,N_11771);
xnor U12400 (N_12400,N_11393,N_10708);
or U12401 (N_12401,N_9236,N_10884);
and U12402 (N_12402,N_10206,N_11008);
xnor U12403 (N_12403,N_10493,N_11812);
or U12404 (N_12404,N_9726,N_10772);
nor U12405 (N_12405,N_9358,N_9907);
and U12406 (N_12406,N_9096,N_10781);
and U12407 (N_12407,N_10439,N_10582);
or U12408 (N_12408,N_10538,N_9577);
nor U12409 (N_12409,N_11928,N_10491);
or U12410 (N_12410,N_9308,N_10892);
or U12411 (N_12411,N_10247,N_11533);
xnor U12412 (N_12412,N_9588,N_10527);
and U12413 (N_12413,N_10867,N_10948);
or U12414 (N_12414,N_10202,N_11728);
xnor U12415 (N_12415,N_9139,N_9477);
or U12416 (N_12416,N_11065,N_10728);
nand U12417 (N_12417,N_9123,N_11191);
and U12418 (N_12418,N_10056,N_9257);
or U12419 (N_12419,N_11384,N_11593);
nand U12420 (N_12420,N_11167,N_10754);
xor U12421 (N_12421,N_9263,N_10986);
nor U12422 (N_12422,N_11639,N_10461);
nand U12423 (N_12423,N_9586,N_11382);
nand U12424 (N_12424,N_10168,N_10256);
or U12425 (N_12425,N_10934,N_11032);
or U12426 (N_12426,N_9708,N_10239);
nor U12427 (N_12427,N_10933,N_10587);
nand U12428 (N_12428,N_10374,N_11660);
xnor U12429 (N_12429,N_10163,N_10184);
nand U12430 (N_12430,N_10243,N_11646);
xor U12431 (N_12431,N_9738,N_11489);
and U12432 (N_12432,N_11747,N_11094);
xor U12433 (N_12433,N_10078,N_10532);
nand U12434 (N_12434,N_11184,N_9488);
xnor U12435 (N_12435,N_10365,N_11080);
xor U12436 (N_12436,N_9124,N_9563);
nand U12437 (N_12437,N_11148,N_11486);
or U12438 (N_12438,N_9762,N_11345);
and U12439 (N_12439,N_9507,N_9424);
or U12440 (N_12440,N_11899,N_11194);
nor U12441 (N_12441,N_10696,N_9014);
and U12442 (N_12442,N_11482,N_11099);
xor U12443 (N_12443,N_9000,N_11027);
nand U12444 (N_12444,N_11485,N_11791);
and U12445 (N_12445,N_11073,N_11506);
or U12446 (N_12446,N_10290,N_9341);
or U12447 (N_12447,N_10573,N_11093);
or U12448 (N_12448,N_10261,N_10037);
nor U12449 (N_12449,N_9007,N_11939);
or U12450 (N_12450,N_11120,N_11906);
and U12451 (N_12451,N_11350,N_9085);
xor U12452 (N_12452,N_9613,N_11266);
nand U12453 (N_12453,N_10998,N_10651);
nor U12454 (N_12454,N_11595,N_9088);
nor U12455 (N_12455,N_10626,N_11991);
and U12456 (N_12456,N_9068,N_11898);
xnor U12457 (N_12457,N_10012,N_10230);
or U12458 (N_12458,N_11368,N_10134);
nor U12459 (N_12459,N_11675,N_11179);
xor U12460 (N_12460,N_10812,N_11516);
or U12461 (N_12461,N_11452,N_9800);
xor U12462 (N_12462,N_10162,N_9379);
or U12463 (N_12463,N_11172,N_10839);
xor U12464 (N_12464,N_9117,N_9938);
or U12465 (N_12465,N_9475,N_9806);
and U12466 (N_12466,N_9052,N_9089);
xor U12467 (N_12467,N_10484,N_10345);
nand U12468 (N_12468,N_10042,N_9687);
and U12469 (N_12469,N_11267,N_9548);
nor U12470 (N_12470,N_11140,N_11768);
or U12471 (N_12471,N_9788,N_11584);
and U12472 (N_12472,N_10841,N_11022);
nand U12473 (N_12473,N_9940,N_10808);
and U12474 (N_12474,N_11851,N_11354);
or U12475 (N_12475,N_11683,N_9190);
nor U12476 (N_12476,N_9899,N_10100);
nor U12477 (N_12477,N_9848,N_11597);
nor U12478 (N_12478,N_10005,N_9856);
xor U12479 (N_12479,N_11652,N_10854);
nor U12480 (N_12480,N_11599,N_10595);
or U12481 (N_12481,N_11860,N_10148);
or U12482 (N_12482,N_10147,N_11242);
nor U12483 (N_12483,N_11115,N_10076);
nor U12484 (N_12484,N_10548,N_9063);
xor U12485 (N_12485,N_9528,N_11772);
xor U12486 (N_12486,N_11790,N_9262);
nand U12487 (N_12487,N_11817,N_10514);
or U12488 (N_12488,N_10031,N_10822);
nor U12489 (N_12489,N_11744,N_10599);
nand U12490 (N_12490,N_9724,N_10441);
nand U12491 (N_12491,N_9466,N_9093);
nand U12492 (N_12492,N_10560,N_9303);
nand U12493 (N_12493,N_10084,N_9876);
xor U12494 (N_12494,N_10606,N_11750);
nand U12495 (N_12495,N_11496,N_11714);
nand U12496 (N_12496,N_9977,N_11606);
xnor U12497 (N_12497,N_11994,N_10596);
or U12498 (N_12498,N_9845,N_10253);
xnor U12499 (N_12499,N_9684,N_9910);
xnor U12500 (N_12500,N_10417,N_11577);
xnor U12501 (N_12501,N_10088,N_11890);
nand U12502 (N_12502,N_9181,N_11708);
or U12503 (N_12503,N_11903,N_9381);
xnor U12504 (N_12504,N_10235,N_11221);
nor U12505 (N_12505,N_11914,N_11003);
and U12506 (N_12506,N_9079,N_11922);
nor U12507 (N_12507,N_10513,N_11825);
nand U12508 (N_12508,N_9592,N_11234);
nand U12509 (N_12509,N_10480,N_9459);
and U12510 (N_12510,N_10286,N_10440);
or U12511 (N_12511,N_9278,N_9004);
or U12512 (N_12512,N_10085,N_10385);
or U12513 (N_12513,N_9241,N_11966);
nor U12514 (N_12514,N_10736,N_10940);
nand U12515 (N_12515,N_9047,N_10302);
xor U12516 (N_12516,N_9693,N_10917);
nand U12517 (N_12517,N_9005,N_10650);
and U12518 (N_12518,N_9471,N_11014);
xor U12519 (N_12519,N_9894,N_10842);
nand U12520 (N_12520,N_11227,N_10902);
or U12521 (N_12521,N_11082,N_9411);
nand U12522 (N_12522,N_9846,N_9043);
or U12523 (N_12523,N_11379,N_11902);
nand U12524 (N_12524,N_11494,N_11959);
or U12525 (N_12525,N_11074,N_9216);
or U12526 (N_12526,N_9566,N_9887);
nor U12527 (N_12527,N_9998,N_10722);
or U12528 (N_12528,N_11590,N_10866);
or U12529 (N_12529,N_11976,N_9268);
and U12530 (N_12530,N_11605,N_11987);
or U12531 (N_12531,N_11837,N_11713);
or U12532 (N_12532,N_9111,N_10301);
nand U12533 (N_12533,N_11570,N_10764);
and U12534 (N_12534,N_11677,N_10137);
xnor U12535 (N_12535,N_10786,N_9706);
or U12536 (N_12536,N_11413,N_11102);
nand U12537 (N_12537,N_10367,N_10359);
and U12538 (N_12538,N_11492,N_9878);
and U12539 (N_12539,N_9398,N_9276);
xor U12540 (N_12540,N_11142,N_10459);
nand U12541 (N_12541,N_11170,N_11411);
nand U12542 (N_12542,N_11285,N_10405);
and U12543 (N_12543,N_9202,N_11291);
and U12544 (N_12544,N_9143,N_10200);
nand U12545 (N_12545,N_10713,N_10520);
and U12546 (N_12546,N_9650,N_9606);
xor U12547 (N_12547,N_10777,N_10328);
and U12548 (N_12548,N_11938,N_10135);
and U12549 (N_12549,N_9637,N_9327);
and U12550 (N_12550,N_10165,N_9787);
and U12551 (N_12551,N_11671,N_10496);
nand U12552 (N_12552,N_11048,N_10637);
and U12553 (N_12553,N_11540,N_11134);
nor U12554 (N_12554,N_11924,N_9581);
nor U12555 (N_12555,N_10284,N_9686);
xnor U12556 (N_12556,N_9553,N_11637);
or U12557 (N_12557,N_9969,N_10638);
and U12558 (N_12558,N_11739,N_10102);
or U12559 (N_12559,N_9048,N_9201);
xor U12560 (N_12560,N_11060,N_10383);
or U12561 (N_12561,N_11331,N_10411);
xor U12562 (N_12562,N_11717,N_9223);
nor U12563 (N_12563,N_9639,N_10997);
or U12564 (N_12564,N_11469,N_11641);
nand U12565 (N_12565,N_9980,N_11909);
nand U12566 (N_12566,N_9703,N_9489);
nand U12567 (N_12567,N_10449,N_10832);
xnor U12568 (N_12568,N_10536,N_10353);
nand U12569 (N_12569,N_11125,N_10909);
nor U12570 (N_12570,N_11394,N_11557);
xnor U12571 (N_12571,N_9799,N_10980);
xor U12572 (N_12572,N_9530,N_11476);
xor U12573 (N_12573,N_9197,N_10992);
nor U12574 (N_12574,N_10186,N_11450);
and U12575 (N_12575,N_10282,N_10624);
xnor U12576 (N_12576,N_10443,N_9500);
or U12577 (N_12577,N_10836,N_10451);
or U12578 (N_12578,N_10123,N_10630);
xor U12579 (N_12579,N_10177,N_9238);
nand U12580 (N_12580,N_10018,N_9961);
xnor U12581 (N_12581,N_11049,N_10881);
and U12582 (N_12582,N_11634,N_9429);
or U12583 (N_12583,N_11527,N_10339);
and U12584 (N_12584,N_10494,N_10381);
or U12585 (N_12585,N_9020,N_11521);
nand U12586 (N_12586,N_10155,N_11619);
and U12587 (N_12587,N_9246,N_10191);
nand U12588 (N_12588,N_10960,N_11400);
nor U12589 (N_12589,N_10830,N_10801);
and U12590 (N_12590,N_11534,N_11387);
xnor U12591 (N_12591,N_9016,N_10994);
or U12592 (N_12592,N_9598,N_9091);
nor U12593 (N_12593,N_11573,N_10815);
nor U12594 (N_12594,N_10488,N_11004);
or U12595 (N_12595,N_10307,N_11759);
and U12596 (N_12596,N_11625,N_10559);
nand U12597 (N_12597,N_11642,N_9937);
or U12598 (N_12598,N_9758,N_9944);
xnor U12599 (N_12599,N_10746,N_9445);
or U12600 (N_12600,N_9943,N_9146);
nand U12601 (N_12601,N_10963,N_10710);
nand U12602 (N_12602,N_11308,N_9412);
nor U12603 (N_12603,N_10723,N_11563);
xnor U12604 (N_12604,N_9215,N_11666);
nor U12605 (N_12605,N_11933,N_9448);
nor U12606 (N_12606,N_10680,N_10616);
or U12607 (N_12607,N_11370,N_11113);
or U12608 (N_12608,N_10531,N_11786);
or U12609 (N_12609,N_9675,N_9735);
or U12610 (N_12610,N_9601,N_10942);
nand U12611 (N_12611,N_10013,N_9222);
nand U12612 (N_12612,N_9023,N_9371);
or U12613 (N_12613,N_9921,N_10949);
and U12614 (N_12614,N_10858,N_9812);
xnor U12615 (N_12615,N_10098,N_11723);
and U12616 (N_12616,N_9155,N_10212);
nor U12617 (N_12617,N_10904,N_9402);
nor U12618 (N_12618,N_11297,N_11289);
nor U12619 (N_12619,N_11253,N_10756);
xnor U12620 (N_12620,N_9287,N_11340);
and U12621 (N_12621,N_9081,N_10370);
and U12622 (N_12622,N_11320,N_9883);
nand U12623 (N_12623,N_10292,N_9685);
nor U12624 (N_12624,N_10259,N_10945);
or U12625 (N_12625,N_10615,N_10845);
xor U12626 (N_12626,N_9347,N_9772);
and U12627 (N_12627,N_9660,N_10126);
nor U12628 (N_12628,N_9362,N_9396);
nand U12629 (N_12629,N_11169,N_10529);
xnor U12630 (N_12630,N_11334,N_11644);
xor U12631 (N_12631,N_11046,N_9547);
nor U12632 (N_12632,N_11879,N_9971);
and U12633 (N_12633,N_11012,N_10355);
nand U12634 (N_12634,N_9988,N_11686);
xnor U12635 (N_12635,N_9291,N_9748);
and U12636 (N_12636,N_9031,N_11178);
and U12637 (N_12637,N_11057,N_10340);
nor U12638 (N_12638,N_10015,N_9546);
nor U12639 (N_12639,N_9832,N_10047);
and U12640 (N_12640,N_10793,N_11270);
and U12641 (N_12641,N_10879,N_10813);
or U12642 (N_12642,N_11423,N_10878);
nor U12643 (N_12643,N_9209,N_9329);
or U12644 (N_12644,N_9512,N_9503);
nor U12645 (N_12645,N_9590,N_9521);
or U12646 (N_12646,N_10823,N_10377);
nand U12647 (N_12647,N_10982,N_10719);
and U12648 (N_12648,N_10922,N_10888);
xnor U12649 (N_12649,N_10293,N_10537);
xor U12650 (N_12650,N_9369,N_10961);
and U12651 (N_12651,N_10500,N_10530);
or U12652 (N_12652,N_10346,N_10679);
or U12653 (N_12653,N_9101,N_11061);
xnor U12654 (N_12654,N_10853,N_10652);
or U12655 (N_12655,N_10711,N_10552);
or U12656 (N_12656,N_11853,N_11975);
and U12657 (N_12657,N_9389,N_10060);
and U12658 (N_12658,N_11963,N_11208);
or U12659 (N_12659,N_11755,N_11894);
nand U12660 (N_12660,N_11920,N_9312);
nand U12661 (N_12661,N_10642,N_9038);
nand U12662 (N_12662,N_9745,N_9857);
nand U12663 (N_12663,N_11659,N_10970);
and U12664 (N_12664,N_11300,N_9529);
and U12665 (N_12665,N_11158,N_9336);
xor U12666 (N_12666,N_9033,N_11787);
or U12667 (N_12667,N_10718,N_11684);
nand U12668 (N_12668,N_11883,N_10802);
nor U12669 (N_12669,N_11907,N_10780);
and U12670 (N_12670,N_9987,N_11547);
or U12671 (N_12671,N_11616,N_11558);
or U12672 (N_12672,N_10178,N_10447);
xor U12673 (N_12673,N_11797,N_9803);
nor U12674 (N_12674,N_11353,N_9253);
nand U12675 (N_12675,N_10700,N_9690);
and U12676 (N_12676,N_9435,N_10255);
or U12677 (N_12677,N_11941,N_9084);
or U12678 (N_12678,N_9929,N_10977);
xor U12679 (N_12679,N_11031,N_9610);
xnor U12680 (N_12680,N_9716,N_11729);
nor U12681 (N_12681,N_9296,N_10787);
and U12682 (N_12682,N_10445,N_9478);
xnor U12683 (N_12683,N_10196,N_10953);
or U12684 (N_12684,N_9365,N_11983);
nor U12685 (N_12685,N_9017,N_11859);
nor U12686 (N_12686,N_9118,N_9364);
and U12687 (N_12687,N_11955,N_11981);
nand U12688 (N_12688,N_9821,N_10995);
and U12689 (N_12689,N_11421,N_10971);
nand U12690 (N_12690,N_9490,N_11445);
xnor U12691 (N_12691,N_10572,N_9032);
nor U12692 (N_12692,N_9884,N_9565);
nor U12693 (N_12693,N_11422,N_11674);
xor U12694 (N_12694,N_9631,N_11510);
xnor U12695 (N_12695,N_9930,N_10453);
nor U12696 (N_12696,N_11974,N_10975);
xor U12697 (N_12697,N_11550,N_10080);
nor U12698 (N_12698,N_11553,N_11442);
nand U12699 (N_12699,N_9095,N_9461);
or U12700 (N_12700,N_10846,N_10285);
nor U12701 (N_12701,N_10104,N_9928);
and U12702 (N_12702,N_11258,N_10380);
xnor U12703 (N_12703,N_9372,N_10773);
nand U12704 (N_12704,N_10589,N_11439);
nand U12705 (N_12705,N_9915,N_9467);
nor U12706 (N_12706,N_10001,N_9353);
nor U12707 (N_12707,N_10627,N_9169);
nand U12708 (N_12708,N_11254,N_9376);
xnor U12709 (N_12709,N_9982,N_10164);
xor U12710 (N_12710,N_11186,N_9019);
xnor U12711 (N_12711,N_9853,N_11151);
and U12712 (N_12712,N_9235,N_9919);
nand U12713 (N_12713,N_10375,N_9447);
xnor U12714 (N_12714,N_10526,N_11823);
nor U12715 (N_12715,N_10868,N_10498);
nand U12716 (N_12716,N_11341,N_10715);
xor U12717 (N_12717,N_9849,N_11583);
nor U12718 (N_12718,N_11433,N_10351);
nor U12719 (N_12719,N_11615,N_9151);
nand U12720 (N_12720,N_9707,N_10192);
nor U12721 (N_12721,N_10661,N_11681);
and U12722 (N_12722,N_9895,N_11029);
and U12723 (N_12723,N_10641,N_9464);
xor U12724 (N_12724,N_11499,N_11617);
and U12725 (N_12725,N_11160,N_11552);
nor U12726 (N_12726,N_11532,N_9506);
or U12727 (N_12727,N_10092,N_9985);
nor U12728 (N_12728,N_10914,N_9897);
nor U12729 (N_12729,N_9171,N_9037);
xor U12730 (N_12730,N_11255,N_11980);
nand U12731 (N_12731,N_9098,N_9652);
nor U12732 (N_12732,N_10393,N_10401);
nor U12733 (N_12733,N_9958,N_9557);
xnor U12734 (N_12734,N_9438,N_9227);
nor U12735 (N_12735,N_11731,N_9747);
nor U12736 (N_12736,N_10782,N_10779);
nand U12737 (N_12737,N_10245,N_9523);
nor U12738 (N_12738,N_9692,N_10352);
nor U12739 (N_12739,N_11814,N_9903);
nor U12740 (N_12740,N_9505,N_9863);
nor U12741 (N_12741,N_10376,N_11834);
and U12742 (N_12742,N_10657,N_10099);
nand U12743 (N_12743,N_10392,N_10965);
nand U12744 (N_12744,N_10964,N_10607);
nor U12745 (N_12745,N_9168,N_9902);
and U12746 (N_12746,N_11107,N_11298);
nor U12747 (N_12747,N_9425,N_9768);
nand U12748 (N_12748,N_11699,N_11329);
nor U12749 (N_12749,N_10141,N_11913);
xor U12750 (N_12750,N_9147,N_11395);
nor U12751 (N_12751,N_9100,N_11611);
xnor U12752 (N_12752,N_10382,N_10086);
nor U12753 (N_12753,N_10454,N_11098);
or U12754 (N_12754,N_10269,N_9368);
or U12755 (N_12755,N_11607,N_9736);
or U12756 (N_12756,N_9042,N_9319);
xnor U12757 (N_12757,N_11749,N_9103);
nor U12758 (N_12758,N_11630,N_11680);
or U12759 (N_12759,N_10506,N_10095);
and U12760 (N_12760,N_9827,N_9356);
or U12761 (N_12761,N_9433,N_10745);
nand U12762 (N_12762,N_11647,N_11736);
nand U12763 (N_12763,N_9370,N_11240);
or U12764 (N_12764,N_10632,N_9715);
nand U12765 (N_12765,N_10683,N_11631);
or U12766 (N_12766,N_9731,N_10051);
xnor U12767 (N_12767,N_11288,N_9330);
and U12768 (N_12768,N_9127,N_10503);
xor U12769 (N_12769,N_11260,N_10487);
or U12770 (N_12770,N_11373,N_11269);
nand U12771 (N_12771,N_10418,N_10331);
and U12772 (N_12772,N_10859,N_10387);
or U12773 (N_12773,N_10705,N_9676);
and U12774 (N_12774,N_9914,N_9649);
or U12775 (N_12775,N_11335,N_9995);
xnor U12776 (N_12776,N_10460,N_9916);
and U12777 (N_12777,N_11710,N_10766);
xor U12778 (N_12778,N_10806,N_9298);
xor U12779 (N_12779,N_10816,N_10278);
nand U12780 (N_12780,N_10923,N_10620);
xor U12781 (N_12781,N_9669,N_11155);
nor U12782 (N_12782,N_11668,N_10726);
or U12783 (N_12783,N_9388,N_9110);
nor U12784 (N_12784,N_11893,N_11171);
nand U12785 (N_12785,N_11716,N_11083);
and U12786 (N_12786,N_10943,N_11321);
and U12787 (N_12787,N_11561,N_10743);
xor U12788 (N_12788,N_10011,N_9206);
or U12789 (N_12789,N_9056,N_11333);
and U12790 (N_12790,N_9867,N_11067);
xor U12791 (N_12791,N_9742,N_9324);
or U12792 (N_12792,N_11556,N_9021);
xor U12793 (N_12793,N_11760,N_10564);
or U12794 (N_12794,N_10057,N_10045);
and U12795 (N_12795,N_9926,N_11819);
nand U12796 (N_12796,N_11166,N_9822);
nor U12797 (N_12797,N_9657,N_9183);
nand U12798 (N_12798,N_10883,N_11706);
nand U12799 (N_12799,N_11918,N_11542);
or U12800 (N_12800,N_11794,N_9638);
nand U12801 (N_12801,N_10767,N_9924);
and U12802 (N_12802,N_11777,N_11338);
or U12803 (N_12803,N_9194,N_11327);
nor U12804 (N_12804,N_10727,N_9614);
xor U12805 (N_12805,N_11543,N_11512);
nand U12806 (N_12806,N_10432,N_9366);
xnor U12807 (N_12807,N_11596,N_9259);
nand U12808 (N_12808,N_11629,N_9029);
nand U12809 (N_12809,N_11690,N_11071);
nand U12810 (N_12810,N_11157,N_9830);
or U12811 (N_12811,N_10431,N_9167);
nand U12812 (N_12812,N_11437,N_10471);
xor U12813 (N_12813,N_10565,N_11096);
and U12814 (N_12814,N_9322,N_11844);
nand U12815 (N_12815,N_11911,N_11287);
xnor U12816 (N_12816,N_11560,N_9307);
or U12817 (N_12817,N_11821,N_9653);
xor U12818 (N_12818,N_11785,N_9695);
or U12819 (N_12819,N_10213,N_10062);
nand U12820 (N_12820,N_9164,N_9723);
nand U12821 (N_12821,N_10783,N_11144);
and U12822 (N_12822,N_11005,N_10792);
xor U12823 (N_12823,N_9451,N_11443);
nor U12824 (N_12824,N_11813,N_11230);
nand U12825 (N_12825,N_10955,N_11640);
or U12826 (N_12826,N_11464,N_10899);
or U12827 (N_12827,N_9701,N_9470);
and U12828 (N_12828,N_11885,N_11618);
nor U12829 (N_12829,N_11491,N_9513);
or U12830 (N_12830,N_10264,N_11449);
xor U12831 (N_12831,N_9254,N_11028);
nor U12832 (N_12832,N_9970,N_9430);
xor U12833 (N_12833,N_9931,N_9309);
xnor U12834 (N_12834,N_9145,N_10551);
xnor U12835 (N_12835,N_11740,N_10033);
xnor U12836 (N_12836,N_11011,N_9220);
and U12837 (N_12837,N_9386,N_11847);
nor U12838 (N_12838,N_10611,N_11703);
nand U12839 (N_12839,N_11722,N_9390);
nor U12840 (N_12840,N_10605,N_10246);
nand U12841 (N_12841,N_10950,N_10721);
xor U12842 (N_12842,N_10602,N_9109);
or U12843 (N_12843,N_10667,N_9550);
and U12844 (N_12844,N_9725,N_11197);
nand U12845 (N_12845,N_11801,N_10897);
or U12846 (N_12846,N_9783,N_11757);
or U12847 (N_12847,N_10869,N_10928);
nor U12848 (N_12848,N_10160,N_9142);
nand U12849 (N_12849,N_9039,N_11838);
xor U12850 (N_12850,N_11081,N_11934);
and U12851 (N_12851,N_9452,N_11525);
nand U12852 (N_12852,N_9229,N_11414);
and U12853 (N_12853,N_10554,N_9864);
or U12854 (N_12854,N_11091,N_9192);
or U12855 (N_12855,N_10799,N_11058);
xnor U12856 (N_12856,N_10662,N_9847);
or U12857 (N_12857,N_11097,N_11578);
or U12858 (N_12858,N_10687,N_10217);
or U12859 (N_12859,N_10778,N_10277);
or U12860 (N_12860,N_10378,N_9159);
nand U12861 (N_12861,N_10218,N_11424);
and U12862 (N_12862,N_10926,N_10577);
nand U12863 (N_12863,N_11493,N_9534);
or U12864 (N_12864,N_9981,N_11539);
xnor U12865 (N_12865,N_9421,N_9597);
or U12866 (N_12866,N_10588,N_10474);
nand U12867 (N_12867,N_9682,N_11435);
xor U12868 (N_12868,N_10584,N_9132);
nand U12869 (N_12869,N_11733,N_10518);
or U12870 (N_12870,N_11753,N_9543);
xor U12871 (N_12871,N_10373,N_9617);
nand U12872 (N_12872,N_10618,N_11656);
or U12873 (N_12873,N_9520,N_9939);
and U12874 (N_12874,N_9568,N_10930);
or U12875 (N_12875,N_9761,N_10807);
or U12876 (N_12876,N_11488,N_11874);
nand U12877 (N_12877,N_11211,N_10912);
xor U12878 (N_12878,N_9320,N_11290);
xnor U12879 (N_12879,N_10931,N_10254);
xor U12880 (N_12880,N_9972,N_10154);
and U12881 (N_12881,N_10108,N_9892);
nand U12882 (N_12882,N_10796,N_9823);
and U12883 (N_12883,N_10988,N_10656);
and U12884 (N_12884,N_10614,N_10534);
xor U12885 (N_12885,N_11121,N_9753);
xnor U12886 (N_12886,N_9423,N_10231);
or U12887 (N_12887,N_10091,N_11779);
nor U12888 (N_12888,N_10161,N_11763);
and U12889 (N_12889,N_9552,N_9825);
or U12890 (N_12890,N_11910,N_10872);
xor U12891 (N_12891,N_11138,N_11371);
or U12892 (N_12892,N_10717,N_11478);
nor U12893 (N_12893,N_9462,N_10609);
xnor U12894 (N_12894,N_10413,N_9323);
or U12895 (N_12895,N_9927,N_9766);
nor U12896 (N_12896,N_10600,N_11111);
nor U12897 (N_12897,N_11326,N_10814);
xor U12898 (N_12898,N_10219,N_11965);
nor U12899 (N_12899,N_11131,N_10545);
and U12900 (N_12900,N_11219,N_9571);
or U12901 (N_12901,N_11245,N_9374);
or U12902 (N_12902,N_10142,N_9912);
nand U12903 (N_12903,N_10643,N_9710);
and U12904 (N_12904,N_9576,N_11069);
nor U12905 (N_12905,N_11628,N_11337);
and U12906 (N_12906,N_10731,N_11087);
or U12907 (N_12907,N_10041,N_10855);
nor U12908 (N_12908,N_9485,N_11700);
nand U12909 (N_12909,N_10043,N_11052);
or U12910 (N_12910,N_9811,N_9984);
xnor U12911 (N_12911,N_11165,N_11474);
or U12912 (N_12912,N_10079,N_11429);
nand U12913 (N_12913,N_9207,N_10320);
or U12914 (N_12914,N_11685,N_10981);
nand U12915 (N_12915,N_10083,N_11085);
or U12916 (N_12916,N_11077,N_10918);
nor U12917 (N_12917,N_11347,N_11957);
nand U12918 (N_12918,N_10706,N_11926);
and U12919 (N_12919,N_11212,N_10361);
nand U12920 (N_12920,N_11023,N_9267);
and U12921 (N_12921,N_10821,N_9870);
or U12922 (N_12922,N_9062,N_11325);
nor U12923 (N_12923,N_9114,N_11839);
nor U12924 (N_12924,N_9882,N_9355);
nor U12925 (N_12925,N_11024,N_9508);
and U12926 (N_12926,N_10660,N_10115);
nand U12927 (N_12927,N_9635,N_10871);
xor U12928 (N_12928,N_10876,N_9722);
xor U12929 (N_12929,N_10138,N_11243);
or U12930 (N_12930,N_10260,N_11889);
nor U12931 (N_12931,N_10035,N_10639);
and U12932 (N_12932,N_11935,N_10759);
and U12933 (N_12933,N_10771,N_11608);
and U12934 (N_12934,N_9826,N_11261);
nand U12935 (N_12935,N_11294,N_9203);
and U12936 (N_12936,N_11042,N_11143);
and U12937 (N_12937,N_11386,N_10490);
nand U12938 (N_12938,N_9394,N_10002);
nor U12939 (N_12939,N_11764,N_10795);
nor U12940 (N_12940,N_9774,N_10762);
nor U12941 (N_12941,N_11296,N_10229);
nand U12942 (N_12942,N_11927,N_11272);
nor U12943 (N_12943,N_9872,N_10575);
nand U12944 (N_12944,N_9491,N_9125);
nor U12945 (N_12945,N_11301,N_11810);
nor U12946 (N_12946,N_11175,N_10798);
nor U12947 (N_12947,N_9556,N_10020);
and U12948 (N_12948,N_10833,N_10818);
or U12949 (N_12949,N_11472,N_11917);
nor U12950 (N_12950,N_10465,N_10004);
nor U12951 (N_12951,N_9185,N_10312);
or U12952 (N_12952,N_9728,N_9258);
nor U12953 (N_12953,N_11041,N_11805);
or U12954 (N_12954,N_11030,N_10058);
or U12955 (N_12955,N_11664,N_10501);
nand U12956 (N_12956,N_10299,N_11852);
or U12957 (N_12957,N_11206,N_9161);
or U12958 (N_12958,N_10182,N_11598);
nor U12959 (N_12959,N_9397,N_9807);
nor U12960 (N_12960,N_11358,N_9049);
xnor U12961 (N_12961,N_10937,N_10216);
nand U12962 (N_12962,N_10133,N_10740);
nand U12963 (N_12963,N_10144,N_11430);
and U12964 (N_12964,N_9282,N_9018);
xnor U12965 (N_12965,N_10522,N_10250);
or U12966 (N_12966,N_11633,N_9442);
or U12967 (N_12967,N_9730,N_11388);
nand U12968 (N_12968,N_11385,N_9403);
or U12969 (N_12969,N_11665,N_9642);
and U12970 (N_12970,N_11145,N_11198);
nand U12971 (N_12971,N_11002,N_9956);
nor U12972 (N_12972,N_9986,N_9230);
nor U12973 (N_12973,N_11154,N_9066);
nor U12974 (N_12974,N_11773,N_10921);
nor U12975 (N_12975,N_9796,N_9689);
or U12976 (N_12976,N_9591,N_10695);
and U12977 (N_12977,N_11409,N_10315);
xor U12978 (N_12978,N_9305,N_10613);
or U12979 (N_12979,N_10294,N_10581);
xnor U12980 (N_12980,N_11724,N_11278);
or U12981 (N_12981,N_9504,N_11025);
xnor U12982 (N_12982,N_10890,N_10873);
xor U12983 (N_12983,N_11312,N_11162);
nand U12984 (N_12984,N_10034,N_10038);
nor U12985 (N_12985,N_10935,N_11876);
xnor U12986 (N_12986,N_10870,N_9141);
or U12987 (N_12987,N_11316,N_10120);
and U12988 (N_12988,N_11524,N_11712);
or U12989 (N_12989,N_11123,N_10848);
nor U12990 (N_12990,N_10430,N_11726);
nor U12991 (N_12991,N_11767,N_11600);
or U12992 (N_12992,N_11305,N_9001);
and U12993 (N_12993,N_9304,N_10860);
xor U12994 (N_12994,N_11233,N_10208);
nor U12995 (N_12995,N_11783,N_11136);
xor U12996 (N_12996,N_10770,N_11010);
xor U12997 (N_12997,N_10054,N_9901);
nor U12998 (N_12998,N_10744,N_11594);
xor U12999 (N_12999,N_10862,N_10249);
nor U13000 (N_13000,N_10558,N_9387);
xnor U13001 (N_13001,N_9889,N_9250);
xor U13002 (N_13002,N_10851,N_10916);
nand U13003 (N_13003,N_9727,N_9498);
nand U13004 (N_13004,N_11205,N_9776);
nor U13005 (N_13005,N_10357,N_11357);
nor U13006 (N_13006,N_10612,N_9838);
and U13007 (N_13007,N_10263,N_11268);
nor U13008 (N_13008,N_9385,N_9137);
or U13009 (N_13009,N_11549,N_9140);
nand U13010 (N_13010,N_11311,N_9083);
nand U13011 (N_13011,N_11416,N_11193);
or U13012 (N_13012,N_9679,N_9840);
xor U13013 (N_13013,N_10507,N_9208);
and U13014 (N_13014,N_9426,N_9808);
or U13015 (N_13015,N_9393,N_11988);
nor U13016 (N_13016,N_10242,N_10579);
nor U13017 (N_13017,N_10547,N_9647);
and U13018 (N_13018,N_10368,N_9691);
xor U13019 (N_13019,N_11816,N_10415);
or U13020 (N_13020,N_9749,N_11410);
or U13021 (N_13021,N_10524,N_10189);
nor U13022 (N_13022,N_11056,N_9060);
nand U13023 (N_13023,N_9869,N_11480);
or U13024 (N_13024,N_11089,N_9214);
or U13025 (N_13025,N_9509,N_11215);
and U13026 (N_13026,N_11440,N_11501);
or U13027 (N_13027,N_9264,N_10167);
xor U13028 (N_13028,N_11192,N_11840);
or U13029 (N_13029,N_9627,N_11470);
or U13030 (N_13030,N_9537,N_9228);
or U13031 (N_13031,N_9480,N_11244);
nor U13032 (N_13032,N_10063,N_9226);
xor U13033 (N_13033,N_11427,N_10116);
or U13034 (N_13034,N_9391,N_11704);
and U13035 (N_13035,N_11505,N_11214);
xnor U13036 (N_13036,N_9769,N_11720);
and U13037 (N_13037,N_11864,N_9953);
or U13038 (N_13038,N_11513,N_9015);
and U13039 (N_13039,N_9663,N_10737);
and U13040 (N_13040,N_10850,N_10039);
and U13041 (N_13041,N_11947,N_9180);
or U13042 (N_13042,N_11754,N_11062);
xor U13043 (N_13043,N_9187,N_10201);
xor U13044 (N_13044,N_10283,N_9771);
and U13045 (N_13045,N_11415,N_9367);
nand U13046 (N_13046,N_9975,N_11009);
nor U13047 (N_13047,N_11035,N_10583);
and U13048 (N_13048,N_10150,N_9409);
or U13049 (N_13049,N_9704,N_9345);
xnor U13050 (N_13050,N_11751,N_10396);
and U13051 (N_13051,N_11571,N_9673);
or U13052 (N_13052,N_9809,N_10156);
or U13053 (N_13053,N_11313,N_11614);
and U13054 (N_13054,N_9595,N_9668);
and U13055 (N_13055,N_10251,N_9493);
and U13056 (N_13056,N_11405,N_9925);
and U13057 (N_13057,N_10050,N_10297);
xor U13058 (N_13058,N_9759,N_9484);
or U13059 (N_13059,N_10467,N_10852);
or U13060 (N_13060,N_9502,N_10388);
and U13061 (N_13061,N_10924,N_10354);
nand U13062 (N_13062,N_11348,N_11122);
xnor U13063 (N_13063,N_10969,N_11982);
nand U13064 (N_13064,N_10332,N_10435);
nand U13065 (N_13065,N_10198,N_10171);
xor U13066 (N_13066,N_11304,N_10419);
or U13067 (N_13067,N_9315,N_11447);
xor U13068 (N_13068,N_9022,N_10688);
xor U13069 (N_13069,N_9828,N_9343);
nand U13070 (N_13070,N_10790,N_10316);
and U13071 (N_13071,N_9332,N_9026);
and U13072 (N_13072,N_9357,N_10699);
nand U13073 (N_13073,N_9698,N_11453);
and U13074 (N_13074,N_10910,N_11076);
or U13075 (N_13075,N_9076,N_10006);
nand U13076 (N_13076,N_9871,N_9640);
nor U13077 (N_13077,N_11428,N_9420);
nand U13078 (N_13078,N_9482,N_9314);
xor U13079 (N_13079,N_9255,N_10566);
or U13080 (N_13080,N_10008,N_10157);
nand U13081 (N_13081,N_11868,N_9793);
nand U13082 (N_13082,N_10372,N_11150);
or U13083 (N_13083,N_9989,N_9175);
and U13084 (N_13084,N_11129,N_9059);
or U13085 (N_13085,N_11711,N_10692);
or U13086 (N_13086,N_9453,N_11958);
nand U13087 (N_13087,N_9955,N_10946);
nor U13088 (N_13088,N_9911,N_11183);
nor U13089 (N_13089,N_11511,N_9407);
and U13090 (N_13090,N_9834,N_10466);
or U13091 (N_13091,N_10390,N_10384);
nor U13092 (N_13092,N_11784,N_9331);
or U13093 (N_13093,N_9536,N_9149);
and U13094 (N_13094,N_9755,N_11672);
nand U13095 (N_13095,N_10072,N_9767);
xor U13096 (N_13096,N_11569,N_10030);
nand U13097 (N_13097,N_10473,N_9760);
nor U13098 (N_13098,N_9113,N_9350);
or U13099 (N_13099,N_10069,N_9457);
xnor U13100 (N_13100,N_10619,N_9431);
nand U13101 (N_13101,N_10119,N_9087);
or U13102 (N_13102,N_9626,N_9752);
and U13103 (N_13103,N_10769,N_10820);
nand U13104 (N_13104,N_10472,N_11483);
xnor U13105 (N_13105,N_11363,N_10592);
nor U13106 (N_13106,N_10896,N_9655);
or U13107 (N_13107,N_10404,N_9221);
nand U13108 (N_13108,N_9622,N_10561);
and U13109 (N_13109,N_11051,N_9086);
or U13110 (N_13110,N_10224,N_9112);
and U13111 (N_13111,N_9497,N_9906);
nand U13112 (N_13112,N_10190,N_10238);
and U13113 (N_13113,N_11572,N_10517);
and U13114 (N_13114,N_10758,N_11330);
nand U13115 (N_13115,N_11782,N_9802);
nor U13116 (N_13116,N_11815,N_11841);
xor U13117 (N_13117,N_9801,N_10521);
xor U13118 (N_13118,N_9859,N_10665);
xnor U13119 (N_13119,N_11473,N_9119);
or U13120 (N_13120,N_9245,N_10205);
nor U13121 (N_13121,N_9392,N_10689);
nor U13122 (N_13122,N_11159,N_10811);
xnor U13123 (N_13123,N_10234,N_11574);
nand U13124 (N_13124,N_9035,N_10911);
nand U13125 (N_13125,N_9659,N_9732);
and U13126 (N_13126,N_9439,N_10009);
xor U13127 (N_13127,N_11200,N_11986);
nor U13128 (N_13128,N_11748,N_9583);
nand U13129 (N_13129,N_11792,N_10789);
nand U13130 (N_13130,N_11399,N_11455);
or U13131 (N_13131,N_11746,N_10457);
nand U13132 (N_13132,N_10228,N_9080);
nor U13133 (N_13133,N_10369,N_11293);
nor U13134 (N_13134,N_11824,N_9933);
and U13135 (N_13135,N_9252,N_9963);
xor U13136 (N_13136,N_11811,N_10515);
and U13137 (N_13137,N_11043,N_10819);
and U13138 (N_13138,N_9596,N_9474);
xnor U13139 (N_13139,N_11624,N_9128);
nor U13140 (N_13140,N_10211,N_9941);
and U13141 (N_13141,N_9605,N_9321);
nor U13142 (N_13142,N_11448,N_11404);
nand U13143 (N_13143,N_10303,N_9789);
nand U13144 (N_13144,N_11996,N_10542);
and U13145 (N_13145,N_9280,N_9837);
or U13146 (N_13146,N_11161,N_11826);
nand U13147 (N_13147,N_10434,N_9248);
xnor U13148 (N_13148,N_9115,N_11039);
nand U13149 (N_13149,N_10040,N_10094);
xnor U13150 (N_13150,N_11271,N_10516);
and U13151 (N_13151,N_10470,N_11952);
xor U13152 (N_13152,N_9349,N_9179);
nand U13153 (N_13153,N_9814,N_10389);
xor U13154 (N_13154,N_9545,N_11795);
and U13155 (N_13155,N_9074,N_11315);
and U13156 (N_13156,N_11544,N_9879);
xnor U13157 (N_13157,N_11514,N_10645);
or U13158 (N_13158,N_10003,N_10972);
xor U13159 (N_13159,N_10775,N_10348);
and U13160 (N_13160,N_11322,N_9090);
xnor U13161 (N_13161,N_10412,N_11344);
xnor U13162 (N_13162,N_11487,N_11721);
nand U13163 (N_13163,N_11103,N_11585);
or U13164 (N_13164,N_11055,N_11796);
and U13165 (N_13165,N_11807,N_9279);
nor U13166 (N_13166,N_10059,N_11888);
or U13167 (N_13167,N_9401,N_11349);
nor U13168 (N_13168,N_9242,N_11591);
xor U13169 (N_13169,N_11915,N_10800);
nor U13170 (N_13170,N_11756,N_10210);
and U13171 (N_13171,N_11854,N_10322);
or U13172 (N_13172,N_11059,N_10032);
nor U13173 (N_13173,N_10730,N_11632);
nor U13174 (N_13174,N_11653,N_11196);
and U13175 (N_13175,N_11376,N_11670);
and U13176 (N_13176,N_10090,N_9865);
xor U13177 (N_13177,N_11587,N_9405);
or U13178 (N_13178,N_9999,N_11188);
and U13179 (N_13179,N_11075,N_10223);
or U13180 (N_13180,N_9414,N_11537);
or U13181 (N_13181,N_9455,N_9792);
or U13182 (N_13182,N_10158,N_10649);
xor U13183 (N_13183,N_11116,N_10684);
xnor U13184 (N_13184,N_9875,N_11936);
nor U13185 (N_13185,N_9077,N_10338);
nor U13186 (N_13186,N_10568,N_11705);
and U13187 (N_13187,N_9711,N_11693);
nor U13188 (N_13188,N_9990,N_11182);
nand U13189 (N_13189,N_11880,N_10703);
xor U13190 (N_13190,N_11793,N_10081);
or U13191 (N_13191,N_11001,N_11283);
xnor U13192 (N_13192,N_10363,N_11845);
nor U13193 (N_13193,N_10794,N_10528);
and U13194 (N_13194,N_10327,N_9277);
or U13195 (N_13195,N_10525,N_9382);
nand U13196 (N_13196,N_9585,N_10757);
nor U13197 (N_13197,N_10631,N_10523);
or U13198 (N_13198,N_11053,N_10197);
and U13199 (N_13199,N_9858,N_10539);
xor U13200 (N_13200,N_10477,N_10673);
nor U13201 (N_13201,N_9009,N_9243);
or U13202 (N_13202,N_9373,N_11940);
nand U13203 (N_13203,N_11190,N_9531);
xnor U13204 (N_13204,N_9905,N_11408);
and U13205 (N_13205,N_11843,N_11401);
and U13206 (N_13206,N_11832,N_9850);
xor U13207 (N_13207,N_11835,N_11407);
nand U13208 (N_13208,N_11610,N_11517);
or U13209 (N_13209,N_9797,N_11460);
and U13210 (N_13210,N_11360,N_11701);
nor U13211 (N_13211,N_9460,N_9302);
nor U13212 (N_13212,N_11036,N_9135);
and U13213 (N_13213,N_10610,N_11284);
and U13214 (N_13214,N_11303,N_9893);
nand U13215 (N_13215,N_9798,N_11118);
or U13216 (N_13216,N_11232,N_9630);
or U13217 (N_13217,N_11589,N_9325);
xnor U13218 (N_13218,N_11015,N_10843);
nand U13219 (N_13219,N_10874,N_10397);
nor U13220 (N_13220,N_9842,N_9479);
nor U13221 (N_13221,N_10540,N_9126);
and U13222 (N_13222,N_10333,N_10675);
nand U13223 (N_13223,N_10763,N_9404);
xor U13224 (N_13224,N_9008,N_9516);
and U13225 (N_13225,N_11559,N_10064);
nand U13226 (N_13226,N_11548,N_11033);
and U13227 (N_13227,N_9852,N_11222);
nand U13228 (N_13228,N_9154,N_10654);
nand U13229 (N_13229,N_10281,N_11090);
nor U13230 (N_13230,N_11431,N_11420);
xnor U13231 (N_13231,N_11367,N_10021);
nor U13232 (N_13232,N_11692,N_9231);
and U13233 (N_13233,N_11808,N_10395);
xnor U13234 (N_13234,N_9313,N_9791);
and U13235 (N_13235,N_11802,N_11412);
xnor U13236 (N_13236,N_10544,N_9178);
and U13237 (N_13237,N_10900,N_9082);
and U13238 (N_13238,N_11523,N_11467);
nand U13239 (N_13239,N_10648,N_11114);
or U13240 (N_13240,N_11836,N_9051);
nor U13241 (N_13241,N_11396,N_11275);
nand U13242 (N_13242,N_9361,N_10753);
nor U13243 (N_13243,N_10483,N_10074);
nand U13244 (N_13244,N_10424,N_9335);
or U13245 (N_13245,N_11117,N_9900);
xor U13246 (N_13246,N_9265,N_9764);
nand U13247 (N_13247,N_9959,N_9483);
or U13248 (N_13248,N_9773,N_10335);
xor U13249 (N_13249,N_10399,N_11034);
nand U13250 (N_13250,N_10709,N_9648);
and U13251 (N_13251,N_10105,N_11109);
xnor U13252 (N_13252,N_11567,N_9170);
nor U13253 (N_13253,N_9611,N_10110);
nand U13254 (N_13254,N_11526,N_11228);
nand U13255 (N_13255,N_9454,N_11235);
nand U13256 (N_13256,N_10944,N_9551);
xnor U13257 (N_13257,N_10936,N_11528);
nand U13258 (N_13258,N_9729,N_9643);
nor U13259 (N_13259,N_9672,N_11895);
and U13260 (N_13260,N_9782,N_10693);
or U13261 (N_13261,N_10433,N_9813);
and U13262 (N_13262,N_9651,N_10067);
xnor U13263 (N_13263,N_11380,N_11522);
and U13264 (N_13264,N_9232,N_10325);
xnor U13265 (N_13265,N_11691,N_11822);
nor U13266 (N_13266,N_10510,N_10735);
and U13267 (N_13267,N_11951,N_10408);
or U13268 (N_13268,N_11112,N_10533);
nand U13269 (N_13269,N_10416,N_11133);
nand U13270 (N_13270,N_10989,N_11375);
or U13271 (N_13271,N_9578,N_9184);
and U13272 (N_13272,N_11126,N_11418);
and U13273 (N_13273,N_11500,N_10623);
xnor U13274 (N_13274,N_11458,N_10991);
or U13275 (N_13275,N_10151,N_9163);
nor U13276 (N_13276,N_10469,N_10071);
or U13277 (N_13277,N_10427,N_11257);
xor U13278 (N_13278,N_11891,N_11973);
or U13279 (N_13279,N_9932,N_9751);
xnor U13280 (N_13280,N_11820,N_9960);
or U13281 (N_13281,N_11441,N_11477);
xnor U13282 (N_13282,N_11905,N_11649);
xor U13283 (N_13283,N_9962,N_11954);
or U13284 (N_13284,N_10751,N_11189);
xnor U13285 (N_13285,N_11203,N_11949);
or U13286 (N_13286,N_11225,N_11063);
nand U13287 (N_13287,N_9979,N_10750);
nor U13288 (N_13288,N_11084,N_10468);
nor U13289 (N_13289,N_9213,N_9555);
or U13290 (N_13290,N_9157,N_11295);
and U13291 (N_13291,N_9511,N_9012);
and U13292 (N_13292,N_11897,N_9599);
and U13293 (N_13293,N_10174,N_10951);
nor U13294 (N_13294,N_9644,N_10826);
and U13295 (N_13295,N_10803,N_9817);
nor U13296 (N_13296,N_10686,N_10456);
and U13297 (N_13297,N_11961,N_9486);
and U13298 (N_13298,N_9075,N_10973);
or U13299 (N_13299,N_10323,N_10175);
or U13300 (N_13300,N_10655,N_9934);
xor U13301 (N_13301,N_9311,N_11045);
nand U13302 (N_13302,N_9580,N_9976);
nor U13303 (N_13303,N_9615,N_10366);
xor U13304 (N_13304,N_10093,N_10429);
xnor U13305 (N_13305,N_9667,N_10570);
nand U13306 (N_13306,N_10300,N_10185);
or U13307 (N_13307,N_11798,N_11105);
nand U13308 (N_13308,N_10768,N_11468);
or U13309 (N_13309,N_10329,N_11580);
nand U13310 (N_13310,N_9351,N_10124);
or U13311 (N_13311,N_10562,N_9636);
nor U13312 (N_13312,N_10668,N_11643);
and U13313 (N_13313,N_9441,N_9200);
xnor U13314 (N_13314,N_10685,N_10647);
xor U13315 (N_13315,N_10747,N_9855);
nor U13316 (N_13316,N_10576,N_9006);
or U13317 (N_13317,N_11273,N_10983);
or U13318 (N_13318,N_9713,N_9072);
and U13319 (N_13319,N_9604,N_9419);
nand U13320 (N_13320,N_11092,N_10423);
and U13321 (N_13321,N_10226,N_11378);
or U13322 (N_13322,N_10109,N_10644);
xor U13323 (N_13323,N_11676,N_9120);
and U13324 (N_13324,N_9522,N_9514);
xor U13325 (N_13325,N_10574,N_11018);
nand U13326 (N_13326,N_9992,N_11997);
nor U13327 (N_13327,N_11545,N_11602);
and U13328 (N_13328,N_11495,N_11119);
nor U13329 (N_13329,N_9947,N_11406);
nand U13330 (N_13330,N_10426,N_10455);
and U13331 (N_13331,N_11515,N_9836);
and U13332 (N_13332,N_11132,N_9994);
xor U13333 (N_13333,N_10990,N_10999);
nor U13334 (N_13334,N_10749,N_10478);
nand U13335 (N_13335,N_11016,N_11220);
nor U13336 (N_13336,N_11989,N_9560);
nor U13337 (N_13337,N_9284,N_10024);
nand U13338 (N_13338,N_11995,N_11892);
nand U13339 (N_13339,N_9107,N_10962);
and U13340 (N_13340,N_11682,N_9674);
and U13341 (N_13341,N_10203,N_10707);
xor U13342 (N_13342,N_9619,N_11174);
nor U13343 (N_13343,N_11309,N_11688);
nand U13344 (N_13344,N_10640,N_10984);
xor U13345 (N_13345,N_9664,N_9138);
and U13346 (N_13346,N_10905,N_10901);
nand U13347 (N_13347,N_10865,N_9712);
nand U13348 (N_13348,N_11735,N_9041);
xnor U13349 (N_13349,N_10237,N_11743);
and U13350 (N_13350,N_10664,N_10010);
nand U13351 (N_13351,N_11137,N_11752);
or U13352 (N_13352,N_9756,N_10199);
nand U13353 (N_13353,N_11503,N_9681);
nor U13354 (N_13354,N_9106,N_9295);
or U13355 (N_13355,N_11662,N_9737);
or U13356 (N_13356,N_11536,N_11846);
and U13357 (N_13357,N_9158,N_11766);
nor U13358 (N_13358,N_11645,N_11381);
xnor U13359 (N_13359,N_9688,N_11436);
or U13360 (N_13360,N_10739,N_9225);
xor U13361 (N_13361,N_10805,N_11226);
or U13362 (N_13362,N_9234,N_9750);
nand U13363 (N_13363,N_9233,N_11872);
xnor U13364 (N_13364,N_9629,N_9354);
nand U13365 (N_13365,N_11833,N_9896);
or U13366 (N_13366,N_10586,N_10209);
or U13367 (N_13367,N_10939,N_9654);
or U13368 (N_13368,N_11374,N_9432);
or U13369 (N_13369,N_11953,N_10257);
and U13370 (N_13370,N_10022,N_10774);
xnor U13371 (N_13371,N_10776,N_11778);
xor U13372 (N_13372,N_11679,N_10358);
or U13373 (N_13373,N_10741,N_10129);
or U13374 (N_13374,N_10330,N_11592);
and U13375 (N_13375,N_11177,N_9408);
nand U13376 (N_13376,N_11299,N_10543);
nand U13377 (N_13377,N_10448,N_10222);
xor U13378 (N_13378,N_11849,N_11263);
nor U13379 (N_13379,N_11912,N_9360);
and U13380 (N_13380,N_9359,N_11403);
nand U13381 (N_13381,N_10266,N_9122);
or U13382 (N_13382,N_9526,N_9108);
or U13383 (N_13383,N_9908,N_11788);
nor U13384 (N_13384,N_11307,N_9065);
nand U13385 (N_13385,N_10541,N_11434);
and U13386 (N_13386,N_9449,N_10061);
nor U13387 (N_13387,N_11829,N_11438);
or U13388 (N_13388,N_9121,N_11519);
nor U13389 (N_13389,N_11657,N_10628);
and U13390 (N_13390,N_10957,N_9340);
nand U13391 (N_13391,N_9129,N_10903);
nor U13392 (N_13392,N_10181,N_9344);
nand U13393 (N_13393,N_10321,N_11663);
nand U13394 (N_13394,N_10827,N_9328);
and U13395 (N_13395,N_9261,N_9237);
xor U13396 (N_13396,N_9299,N_11019);
nor U13397 (N_13397,N_9380,N_11465);
nand U13398 (N_13398,N_9573,N_9997);
nand U13399 (N_13399,N_9795,N_11377);
nor U13400 (N_13400,N_9778,N_10146);
or U13401 (N_13401,N_11149,N_9437);
xor U13402 (N_13402,N_9671,N_9272);
nor U13403 (N_13403,N_9116,N_9885);
xnor U13404 (N_13404,N_9607,N_10569);
nand U13405 (N_13405,N_10738,N_9757);
and U13406 (N_13406,N_11962,N_10342);
and U13407 (N_13407,N_11809,N_10394);
and U13408 (N_13408,N_10489,N_10920);
or U13409 (N_13409,N_10318,N_9446);
or U13410 (N_13410,N_9515,N_10729);
nor U13411 (N_13411,N_9011,N_11479);
nand U13412 (N_13412,N_9913,N_9527);
or U13413 (N_13413,N_11862,N_11789);
and U13414 (N_13414,N_11021,N_11484);
or U13415 (N_13415,N_11984,N_10475);
and U13416 (N_13416,N_11498,N_9935);
nor U13417 (N_13417,N_10274,N_9584);
xnor U13418 (N_13418,N_11875,N_11355);
nand U13419 (N_13419,N_11223,N_9501);
nand U13420 (N_13420,N_10139,N_10343);
xnor U13421 (N_13421,N_10797,N_10204);
or U13422 (N_13422,N_11725,N_9417);
nand U13423 (N_13423,N_9658,N_10959);
nand U13424 (N_13424,N_11604,N_11366);
nor U13425 (N_13425,N_11576,N_9696);
nor U13426 (N_13426,N_9564,N_11873);
xnor U13427 (N_13427,N_11960,N_11509);
nor U13428 (N_13428,N_9881,N_9150);
and U13429 (N_13429,N_11661,N_10313);
or U13430 (N_13430,N_9198,N_9740);
nand U13431 (N_13431,N_9542,N_11929);
or U13432 (N_13432,N_9210,N_11564);
nand U13433 (N_13433,N_10509,N_10958);
xor U13434 (N_13434,N_11104,N_9003);
and U13435 (N_13435,N_10436,N_11173);
and U13436 (N_13436,N_9805,N_9765);
and U13437 (N_13437,N_9010,N_9624);
nor U13438 (N_13438,N_11635,N_10172);
xnor U13439 (N_13439,N_10324,N_11224);
nor U13440 (N_13440,N_9104,N_11050);
xor U13441 (N_13441,N_9044,N_9174);
nor U13442 (N_13442,N_9983,N_10880);
xnor U13443 (N_13443,N_9260,N_10356);
nor U13444 (N_13444,N_11887,N_9633);
nand U13445 (N_13445,N_9153,N_11390);
or U13446 (N_13446,N_11865,N_9854);
or U13447 (N_13447,N_10555,N_10829);
nand U13448 (N_13448,N_10276,N_9070);
or U13449 (N_13449,N_9594,N_9535);
nand U13450 (N_13450,N_11070,N_10207);
and U13451 (N_13451,N_10117,N_10974);
or U13452 (N_13452,N_11276,N_11582);
nor U13453 (N_13453,N_9816,N_10976);
nor U13454 (N_13454,N_9078,N_11972);
nand U13455 (N_13455,N_9790,N_11719);
xnor U13456 (N_13456,N_11694,N_9400);
or U13457 (N_13457,N_9294,N_9839);
and U13458 (N_13458,N_10495,N_11857);
nand U13459 (N_13459,N_9024,N_9835);
xor U13460 (N_13460,N_11239,N_10585);
nor U13461 (N_13461,N_10925,N_11139);
xor U13462 (N_13462,N_11861,N_11804);
or U13463 (N_13463,N_10288,N_9920);
xor U13464 (N_13464,N_10153,N_9670);
nor U13465 (N_13465,N_10136,N_9317);
nor U13466 (N_13466,N_9212,N_11856);
nand U13467 (N_13467,N_10166,N_9025);
xor U13468 (N_13468,N_10621,N_10784);
or U13469 (N_13469,N_9623,N_11956);
xnor U13470 (N_13470,N_9993,N_11943);
or U13471 (N_13471,N_10908,N_10929);
or U13472 (N_13472,N_11758,N_11000);
and U13473 (N_13473,N_9249,N_9251);
and U13474 (N_13474,N_9719,N_11319);
xnor U13475 (N_13475,N_9621,N_10979);
xnor U13476 (N_13476,N_10087,N_9468);
and U13477 (N_13477,N_9166,N_9172);
or U13478 (N_13478,N_11999,N_11867);
or U13479 (N_13479,N_10428,N_10442);
or U13480 (N_13480,N_11507,N_10817);
nand U13481 (N_13481,N_11047,N_11389);
nor U13482 (N_13482,N_10036,N_9616);
xnor U13483 (N_13483,N_9105,N_9661);
nor U13484 (N_13484,N_9991,N_11280);
or U13485 (N_13485,N_10140,N_10546);
nor U13486 (N_13486,N_10887,N_9744);
nor U13487 (N_13487,N_10371,N_9700);
nand U13488 (N_13488,N_11199,N_10479);
and U13489 (N_13489,N_9815,N_9269);
xnor U13490 (N_13490,N_11904,N_10915);
nor U13491 (N_13491,N_9292,N_10188);
or U13492 (N_13492,N_11040,N_10112);
or U13493 (N_13493,N_11328,N_10597);
nor U13494 (N_13494,N_11612,N_11916);
nor U13495 (N_13495,N_11937,N_9073);
nand U13496 (N_13496,N_10068,N_9946);
xnor U13497 (N_13497,N_9978,N_9094);
xnor U13498 (N_13498,N_11318,N_9777);
nor U13499 (N_13499,N_9131,N_10927);
xnor U13500 (N_13500,N_11376,N_11320);
and U13501 (N_13501,N_10696,N_11813);
nand U13502 (N_13502,N_9789,N_10428);
xor U13503 (N_13503,N_10619,N_11663);
nand U13504 (N_13504,N_11992,N_11635);
nor U13505 (N_13505,N_11012,N_11178);
or U13506 (N_13506,N_9179,N_10926);
nand U13507 (N_13507,N_9009,N_9029);
or U13508 (N_13508,N_9326,N_9095);
nand U13509 (N_13509,N_9915,N_9937);
and U13510 (N_13510,N_11720,N_9977);
xnor U13511 (N_13511,N_10564,N_11511);
nor U13512 (N_13512,N_10473,N_11311);
xnor U13513 (N_13513,N_10805,N_10266);
xnor U13514 (N_13514,N_9945,N_9212);
nand U13515 (N_13515,N_10040,N_11442);
and U13516 (N_13516,N_10871,N_10719);
nor U13517 (N_13517,N_11314,N_9245);
nand U13518 (N_13518,N_10750,N_9382);
nor U13519 (N_13519,N_11815,N_10987);
nand U13520 (N_13520,N_11906,N_9969);
xnor U13521 (N_13521,N_9729,N_9975);
nand U13522 (N_13522,N_10629,N_11864);
nand U13523 (N_13523,N_9306,N_10188);
or U13524 (N_13524,N_9282,N_10876);
and U13525 (N_13525,N_9303,N_10183);
xor U13526 (N_13526,N_10674,N_11430);
xnor U13527 (N_13527,N_11229,N_11136);
nor U13528 (N_13528,N_10973,N_9590);
or U13529 (N_13529,N_11331,N_9796);
xor U13530 (N_13530,N_9207,N_10169);
or U13531 (N_13531,N_10414,N_9641);
and U13532 (N_13532,N_10770,N_9797);
or U13533 (N_13533,N_10567,N_10864);
or U13534 (N_13534,N_10886,N_10665);
nand U13535 (N_13535,N_10125,N_9898);
or U13536 (N_13536,N_11556,N_11681);
nor U13537 (N_13537,N_10340,N_11901);
nor U13538 (N_13538,N_9358,N_10720);
or U13539 (N_13539,N_10109,N_11422);
and U13540 (N_13540,N_10225,N_9238);
xnor U13541 (N_13541,N_9844,N_10149);
or U13542 (N_13542,N_10850,N_11295);
or U13543 (N_13543,N_10624,N_10271);
nor U13544 (N_13544,N_10117,N_9424);
and U13545 (N_13545,N_10241,N_11758);
or U13546 (N_13546,N_9072,N_9390);
xor U13547 (N_13547,N_11160,N_10187);
and U13548 (N_13548,N_9098,N_9749);
nor U13549 (N_13549,N_9685,N_10621);
nand U13550 (N_13550,N_11659,N_11802);
xor U13551 (N_13551,N_11091,N_10445);
and U13552 (N_13552,N_11792,N_10905);
or U13553 (N_13553,N_9097,N_10695);
and U13554 (N_13554,N_9532,N_10756);
and U13555 (N_13555,N_9039,N_10020);
xor U13556 (N_13556,N_10280,N_10252);
nand U13557 (N_13557,N_11799,N_11365);
nand U13558 (N_13558,N_11414,N_10875);
or U13559 (N_13559,N_9339,N_9181);
or U13560 (N_13560,N_11212,N_10282);
nand U13561 (N_13561,N_10385,N_9567);
and U13562 (N_13562,N_10380,N_11174);
xor U13563 (N_13563,N_11229,N_11005);
or U13564 (N_13564,N_9820,N_9671);
xnor U13565 (N_13565,N_10371,N_9742);
nor U13566 (N_13566,N_10765,N_9134);
xor U13567 (N_13567,N_11042,N_9490);
and U13568 (N_13568,N_9299,N_11142);
and U13569 (N_13569,N_10394,N_9022);
nand U13570 (N_13570,N_11385,N_10815);
and U13571 (N_13571,N_10031,N_11216);
or U13572 (N_13572,N_10748,N_9646);
xnor U13573 (N_13573,N_10599,N_9192);
or U13574 (N_13574,N_11320,N_11375);
nor U13575 (N_13575,N_11820,N_11283);
or U13576 (N_13576,N_11347,N_9369);
nand U13577 (N_13577,N_11600,N_11634);
nor U13578 (N_13578,N_9547,N_11580);
nand U13579 (N_13579,N_10203,N_9443);
or U13580 (N_13580,N_11598,N_11144);
or U13581 (N_13581,N_11235,N_11002);
nand U13582 (N_13582,N_11961,N_10653);
and U13583 (N_13583,N_10837,N_9677);
and U13584 (N_13584,N_10299,N_9058);
nand U13585 (N_13585,N_10150,N_11017);
nand U13586 (N_13586,N_10940,N_10691);
and U13587 (N_13587,N_10648,N_9097);
xnor U13588 (N_13588,N_11553,N_9652);
nand U13589 (N_13589,N_11405,N_11369);
nor U13590 (N_13590,N_10712,N_9448);
nor U13591 (N_13591,N_11634,N_9338);
and U13592 (N_13592,N_10946,N_9535);
nor U13593 (N_13593,N_9064,N_9048);
xnor U13594 (N_13594,N_9226,N_10962);
nand U13595 (N_13595,N_10923,N_11816);
xor U13596 (N_13596,N_9860,N_10019);
and U13597 (N_13597,N_11481,N_10402);
nor U13598 (N_13598,N_10075,N_9379);
nand U13599 (N_13599,N_11480,N_9130);
or U13600 (N_13600,N_9378,N_11251);
nand U13601 (N_13601,N_9960,N_10600);
or U13602 (N_13602,N_10435,N_11756);
xor U13603 (N_13603,N_9514,N_11069);
nor U13604 (N_13604,N_11382,N_10133);
or U13605 (N_13605,N_11213,N_10914);
and U13606 (N_13606,N_9793,N_11674);
nand U13607 (N_13607,N_11435,N_10607);
and U13608 (N_13608,N_10605,N_10209);
nor U13609 (N_13609,N_9808,N_9749);
xnor U13610 (N_13610,N_10776,N_9623);
or U13611 (N_13611,N_9500,N_10069);
nor U13612 (N_13612,N_11491,N_9569);
xor U13613 (N_13613,N_11884,N_11704);
or U13614 (N_13614,N_10289,N_9814);
nand U13615 (N_13615,N_10469,N_11555);
nand U13616 (N_13616,N_10812,N_11168);
xnor U13617 (N_13617,N_9765,N_10141);
nor U13618 (N_13618,N_9260,N_9853);
xor U13619 (N_13619,N_11135,N_9976);
nand U13620 (N_13620,N_9333,N_11440);
xor U13621 (N_13621,N_11142,N_11731);
nor U13622 (N_13622,N_11473,N_11142);
xnor U13623 (N_13623,N_11584,N_11395);
or U13624 (N_13624,N_10862,N_10389);
or U13625 (N_13625,N_9059,N_11744);
nand U13626 (N_13626,N_11870,N_9510);
nand U13627 (N_13627,N_11215,N_11648);
xnor U13628 (N_13628,N_9671,N_11082);
nor U13629 (N_13629,N_9139,N_9865);
nand U13630 (N_13630,N_10628,N_9784);
or U13631 (N_13631,N_9917,N_11446);
or U13632 (N_13632,N_11378,N_11747);
nor U13633 (N_13633,N_10709,N_9974);
nand U13634 (N_13634,N_10712,N_10640);
nor U13635 (N_13635,N_11535,N_11491);
nand U13636 (N_13636,N_10564,N_11409);
or U13637 (N_13637,N_10592,N_10643);
nor U13638 (N_13638,N_10159,N_11712);
or U13639 (N_13639,N_10180,N_9372);
xnor U13640 (N_13640,N_9121,N_11194);
or U13641 (N_13641,N_11323,N_9496);
nand U13642 (N_13642,N_9981,N_10875);
nand U13643 (N_13643,N_11264,N_10958);
xor U13644 (N_13644,N_10750,N_9671);
and U13645 (N_13645,N_9367,N_10126);
nor U13646 (N_13646,N_11878,N_10373);
xor U13647 (N_13647,N_10420,N_11684);
nor U13648 (N_13648,N_9591,N_11308);
nor U13649 (N_13649,N_9498,N_9712);
nor U13650 (N_13650,N_9670,N_11552);
nand U13651 (N_13651,N_10006,N_9256);
and U13652 (N_13652,N_11747,N_10732);
nand U13653 (N_13653,N_11807,N_9685);
nand U13654 (N_13654,N_10722,N_11775);
xor U13655 (N_13655,N_10535,N_10819);
and U13656 (N_13656,N_11468,N_9456);
nor U13657 (N_13657,N_10564,N_9847);
nand U13658 (N_13658,N_11110,N_11766);
and U13659 (N_13659,N_9056,N_9070);
and U13660 (N_13660,N_9543,N_10062);
xor U13661 (N_13661,N_10689,N_11783);
and U13662 (N_13662,N_11032,N_10360);
nand U13663 (N_13663,N_10433,N_10860);
nor U13664 (N_13664,N_10885,N_11123);
or U13665 (N_13665,N_10484,N_10207);
nor U13666 (N_13666,N_9420,N_10539);
or U13667 (N_13667,N_10816,N_10849);
xnor U13668 (N_13668,N_9551,N_11984);
or U13669 (N_13669,N_9908,N_10585);
xnor U13670 (N_13670,N_10451,N_11400);
nand U13671 (N_13671,N_10329,N_10228);
nor U13672 (N_13672,N_10542,N_10825);
nand U13673 (N_13673,N_11455,N_10351);
xor U13674 (N_13674,N_10367,N_11033);
and U13675 (N_13675,N_10216,N_11226);
nor U13676 (N_13676,N_10826,N_9410);
xnor U13677 (N_13677,N_9531,N_10841);
nor U13678 (N_13678,N_10420,N_9148);
or U13679 (N_13679,N_9356,N_10151);
nand U13680 (N_13680,N_9189,N_10150);
and U13681 (N_13681,N_11195,N_10886);
and U13682 (N_13682,N_9002,N_9455);
nor U13683 (N_13683,N_11865,N_11663);
nand U13684 (N_13684,N_10079,N_9098);
xnor U13685 (N_13685,N_9352,N_11612);
nor U13686 (N_13686,N_9124,N_11620);
or U13687 (N_13687,N_11672,N_10761);
nand U13688 (N_13688,N_11052,N_9873);
nand U13689 (N_13689,N_11109,N_11895);
xor U13690 (N_13690,N_11177,N_11411);
nor U13691 (N_13691,N_11475,N_10144);
and U13692 (N_13692,N_11169,N_10064);
xnor U13693 (N_13693,N_10742,N_9695);
and U13694 (N_13694,N_9845,N_9195);
and U13695 (N_13695,N_10596,N_10249);
and U13696 (N_13696,N_11177,N_9685);
and U13697 (N_13697,N_11786,N_10233);
and U13698 (N_13698,N_9630,N_9189);
and U13699 (N_13699,N_11187,N_9574);
xnor U13700 (N_13700,N_9227,N_9898);
nand U13701 (N_13701,N_11423,N_11395);
nor U13702 (N_13702,N_11724,N_9374);
nor U13703 (N_13703,N_11219,N_11113);
nand U13704 (N_13704,N_10993,N_11498);
or U13705 (N_13705,N_11558,N_9238);
xor U13706 (N_13706,N_11558,N_9525);
xnor U13707 (N_13707,N_11819,N_9787);
or U13708 (N_13708,N_11264,N_11865);
and U13709 (N_13709,N_11845,N_10776);
or U13710 (N_13710,N_11241,N_11783);
nand U13711 (N_13711,N_9378,N_10259);
nor U13712 (N_13712,N_9072,N_9426);
or U13713 (N_13713,N_11654,N_10157);
nand U13714 (N_13714,N_11718,N_9135);
xor U13715 (N_13715,N_11802,N_10740);
xor U13716 (N_13716,N_10015,N_10125);
nand U13717 (N_13717,N_9444,N_11080);
xnor U13718 (N_13718,N_11230,N_9835);
nor U13719 (N_13719,N_10544,N_9429);
nand U13720 (N_13720,N_11192,N_9333);
or U13721 (N_13721,N_11954,N_9322);
or U13722 (N_13722,N_10351,N_9590);
nand U13723 (N_13723,N_9844,N_9767);
or U13724 (N_13724,N_9138,N_9102);
xnor U13725 (N_13725,N_11608,N_11174);
and U13726 (N_13726,N_11797,N_11075);
nand U13727 (N_13727,N_11217,N_10691);
xnor U13728 (N_13728,N_10587,N_10846);
xor U13729 (N_13729,N_10256,N_9385);
xor U13730 (N_13730,N_10871,N_11056);
xnor U13731 (N_13731,N_11799,N_9701);
nand U13732 (N_13732,N_11655,N_11307);
nand U13733 (N_13733,N_10318,N_9954);
nand U13734 (N_13734,N_11716,N_11976);
xor U13735 (N_13735,N_10597,N_11813);
nor U13736 (N_13736,N_9482,N_11304);
nor U13737 (N_13737,N_10193,N_11830);
nand U13738 (N_13738,N_11559,N_11959);
xor U13739 (N_13739,N_9424,N_9401);
and U13740 (N_13740,N_9075,N_11187);
nand U13741 (N_13741,N_11019,N_10836);
and U13742 (N_13742,N_11492,N_11041);
nand U13743 (N_13743,N_11923,N_11456);
nor U13744 (N_13744,N_11512,N_11027);
xor U13745 (N_13745,N_10860,N_9402);
and U13746 (N_13746,N_10709,N_10627);
nand U13747 (N_13747,N_11032,N_10008);
nor U13748 (N_13748,N_10352,N_11552);
and U13749 (N_13749,N_9166,N_10194);
nand U13750 (N_13750,N_10616,N_11057);
xnor U13751 (N_13751,N_11153,N_10739);
nor U13752 (N_13752,N_10945,N_10855);
and U13753 (N_13753,N_11853,N_9097);
or U13754 (N_13754,N_10423,N_9811);
nand U13755 (N_13755,N_10721,N_9203);
nand U13756 (N_13756,N_11868,N_10361);
and U13757 (N_13757,N_11632,N_10703);
or U13758 (N_13758,N_11179,N_11422);
or U13759 (N_13759,N_11556,N_10459);
xnor U13760 (N_13760,N_10905,N_9842);
nor U13761 (N_13761,N_10281,N_11552);
or U13762 (N_13762,N_9199,N_9434);
nand U13763 (N_13763,N_9878,N_11870);
and U13764 (N_13764,N_9136,N_10439);
or U13765 (N_13765,N_9564,N_10458);
xnor U13766 (N_13766,N_11913,N_10155);
or U13767 (N_13767,N_11713,N_11625);
and U13768 (N_13768,N_10204,N_9620);
nand U13769 (N_13769,N_10314,N_10636);
and U13770 (N_13770,N_10361,N_9128);
nand U13771 (N_13771,N_10230,N_9663);
or U13772 (N_13772,N_9561,N_10613);
and U13773 (N_13773,N_10666,N_11145);
and U13774 (N_13774,N_11821,N_10807);
nand U13775 (N_13775,N_11513,N_10508);
xnor U13776 (N_13776,N_10827,N_11013);
or U13777 (N_13777,N_9252,N_9004);
xor U13778 (N_13778,N_9388,N_11665);
or U13779 (N_13779,N_11558,N_10761);
xnor U13780 (N_13780,N_9159,N_9757);
and U13781 (N_13781,N_11812,N_11775);
nand U13782 (N_13782,N_11663,N_9486);
xor U13783 (N_13783,N_11567,N_9292);
and U13784 (N_13784,N_11423,N_9697);
and U13785 (N_13785,N_9376,N_10724);
and U13786 (N_13786,N_11350,N_9513);
nand U13787 (N_13787,N_10021,N_10232);
nand U13788 (N_13788,N_10566,N_10942);
xor U13789 (N_13789,N_9747,N_9859);
or U13790 (N_13790,N_11931,N_9539);
or U13791 (N_13791,N_10141,N_11075);
and U13792 (N_13792,N_11392,N_10923);
nand U13793 (N_13793,N_9450,N_10946);
xnor U13794 (N_13794,N_10543,N_10559);
and U13795 (N_13795,N_10813,N_9063);
and U13796 (N_13796,N_9411,N_9935);
nand U13797 (N_13797,N_9239,N_11852);
xor U13798 (N_13798,N_10664,N_11524);
nor U13799 (N_13799,N_11891,N_9769);
nor U13800 (N_13800,N_11899,N_9700);
nand U13801 (N_13801,N_9366,N_9950);
and U13802 (N_13802,N_11049,N_9943);
xor U13803 (N_13803,N_10950,N_10648);
nor U13804 (N_13804,N_11170,N_9655);
nand U13805 (N_13805,N_11791,N_11272);
or U13806 (N_13806,N_10492,N_11472);
xor U13807 (N_13807,N_10972,N_9265);
and U13808 (N_13808,N_9979,N_11287);
nor U13809 (N_13809,N_11797,N_10453);
nor U13810 (N_13810,N_11418,N_9667);
nor U13811 (N_13811,N_10626,N_10230);
or U13812 (N_13812,N_11946,N_11168);
or U13813 (N_13813,N_11292,N_10969);
and U13814 (N_13814,N_10600,N_9674);
or U13815 (N_13815,N_9623,N_9320);
xnor U13816 (N_13816,N_11649,N_10913);
or U13817 (N_13817,N_9864,N_11399);
or U13818 (N_13818,N_9302,N_10527);
nand U13819 (N_13819,N_11643,N_9118);
nor U13820 (N_13820,N_10585,N_11966);
or U13821 (N_13821,N_10273,N_9079);
or U13822 (N_13822,N_10135,N_11669);
nor U13823 (N_13823,N_9055,N_9982);
nand U13824 (N_13824,N_9820,N_9654);
xnor U13825 (N_13825,N_9723,N_9471);
xor U13826 (N_13826,N_9499,N_9994);
nor U13827 (N_13827,N_10780,N_10616);
or U13828 (N_13828,N_9554,N_11672);
or U13829 (N_13829,N_11586,N_10735);
xnor U13830 (N_13830,N_11541,N_11575);
nand U13831 (N_13831,N_9995,N_9735);
xor U13832 (N_13832,N_9949,N_11011);
and U13833 (N_13833,N_10442,N_10914);
nand U13834 (N_13834,N_11161,N_10531);
nor U13835 (N_13835,N_10277,N_10259);
and U13836 (N_13836,N_10095,N_10957);
and U13837 (N_13837,N_10365,N_10462);
nand U13838 (N_13838,N_9322,N_10188);
xor U13839 (N_13839,N_9302,N_10800);
nor U13840 (N_13840,N_9415,N_11310);
and U13841 (N_13841,N_11605,N_11236);
and U13842 (N_13842,N_11874,N_10351);
and U13843 (N_13843,N_9687,N_10508);
or U13844 (N_13844,N_11580,N_10516);
xnor U13845 (N_13845,N_11375,N_10900);
nand U13846 (N_13846,N_9393,N_11934);
nor U13847 (N_13847,N_11284,N_11639);
and U13848 (N_13848,N_10770,N_10016);
nand U13849 (N_13849,N_11765,N_11134);
and U13850 (N_13850,N_11475,N_10854);
and U13851 (N_13851,N_10757,N_10466);
or U13852 (N_13852,N_9124,N_11597);
or U13853 (N_13853,N_10311,N_11294);
and U13854 (N_13854,N_9707,N_10544);
nand U13855 (N_13855,N_11306,N_10147);
xor U13856 (N_13856,N_11771,N_9112);
nor U13857 (N_13857,N_10027,N_10830);
nor U13858 (N_13858,N_10982,N_10318);
and U13859 (N_13859,N_11053,N_9598);
nand U13860 (N_13860,N_10266,N_9935);
nor U13861 (N_13861,N_10888,N_11362);
nand U13862 (N_13862,N_9298,N_11960);
nor U13863 (N_13863,N_11512,N_10466);
nor U13864 (N_13864,N_11323,N_10885);
xor U13865 (N_13865,N_10963,N_9816);
or U13866 (N_13866,N_9509,N_9254);
and U13867 (N_13867,N_11083,N_11516);
xor U13868 (N_13868,N_9551,N_11439);
nor U13869 (N_13869,N_10788,N_9364);
nand U13870 (N_13870,N_9166,N_10985);
nand U13871 (N_13871,N_9328,N_11900);
nor U13872 (N_13872,N_11414,N_10227);
and U13873 (N_13873,N_9641,N_10079);
xnor U13874 (N_13874,N_11613,N_9093);
nor U13875 (N_13875,N_11535,N_10756);
or U13876 (N_13876,N_11222,N_9067);
or U13877 (N_13877,N_9765,N_10259);
nor U13878 (N_13878,N_11169,N_10417);
xnor U13879 (N_13879,N_11556,N_10088);
nand U13880 (N_13880,N_11952,N_10162);
nand U13881 (N_13881,N_9550,N_11301);
nand U13882 (N_13882,N_10961,N_11377);
nor U13883 (N_13883,N_10971,N_10707);
or U13884 (N_13884,N_10085,N_9160);
or U13885 (N_13885,N_9630,N_10486);
or U13886 (N_13886,N_11722,N_9901);
xnor U13887 (N_13887,N_10401,N_9585);
and U13888 (N_13888,N_10428,N_11838);
nor U13889 (N_13889,N_10881,N_11057);
nand U13890 (N_13890,N_9313,N_9825);
nand U13891 (N_13891,N_10264,N_10282);
xnor U13892 (N_13892,N_10284,N_9871);
xor U13893 (N_13893,N_9976,N_9998);
nor U13894 (N_13894,N_11919,N_9864);
xnor U13895 (N_13895,N_10584,N_9791);
xor U13896 (N_13896,N_10905,N_11469);
xnor U13897 (N_13897,N_10738,N_11932);
and U13898 (N_13898,N_11649,N_10656);
or U13899 (N_13899,N_10467,N_10312);
nor U13900 (N_13900,N_9543,N_10714);
nand U13901 (N_13901,N_9781,N_10326);
and U13902 (N_13902,N_11629,N_11139);
nand U13903 (N_13903,N_11144,N_11121);
nand U13904 (N_13904,N_9384,N_9203);
and U13905 (N_13905,N_9988,N_11870);
xor U13906 (N_13906,N_10685,N_9804);
nor U13907 (N_13907,N_9831,N_11838);
nand U13908 (N_13908,N_9685,N_11492);
xnor U13909 (N_13909,N_11827,N_10838);
nand U13910 (N_13910,N_9184,N_11185);
xnor U13911 (N_13911,N_10184,N_10337);
or U13912 (N_13912,N_11075,N_10475);
nor U13913 (N_13913,N_11560,N_10244);
and U13914 (N_13914,N_10910,N_11478);
or U13915 (N_13915,N_9067,N_10651);
nor U13916 (N_13916,N_9800,N_10289);
and U13917 (N_13917,N_11222,N_10635);
and U13918 (N_13918,N_10427,N_11656);
nor U13919 (N_13919,N_9974,N_11890);
and U13920 (N_13920,N_11189,N_9559);
nor U13921 (N_13921,N_10471,N_9044);
nor U13922 (N_13922,N_10332,N_10640);
or U13923 (N_13923,N_11474,N_10591);
or U13924 (N_13924,N_11377,N_9461);
xor U13925 (N_13925,N_9208,N_11731);
and U13926 (N_13926,N_11178,N_10291);
nand U13927 (N_13927,N_11678,N_9297);
nor U13928 (N_13928,N_10131,N_10811);
or U13929 (N_13929,N_9776,N_11887);
nor U13930 (N_13930,N_11950,N_9841);
nor U13931 (N_13931,N_11200,N_9048);
or U13932 (N_13932,N_11470,N_11307);
and U13933 (N_13933,N_11988,N_11727);
nor U13934 (N_13934,N_9314,N_11102);
nand U13935 (N_13935,N_11385,N_9758);
nand U13936 (N_13936,N_11343,N_9531);
nor U13937 (N_13937,N_9919,N_9756);
nor U13938 (N_13938,N_9974,N_10114);
nor U13939 (N_13939,N_9076,N_11803);
xor U13940 (N_13940,N_9825,N_10229);
xnor U13941 (N_13941,N_9597,N_11288);
and U13942 (N_13942,N_9594,N_10219);
nor U13943 (N_13943,N_9122,N_10301);
or U13944 (N_13944,N_10789,N_9040);
nand U13945 (N_13945,N_9232,N_9683);
nand U13946 (N_13946,N_10950,N_11480);
nor U13947 (N_13947,N_9120,N_10786);
or U13948 (N_13948,N_9100,N_9557);
and U13949 (N_13949,N_9621,N_9321);
nand U13950 (N_13950,N_10286,N_10853);
nand U13951 (N_13951,N_9863,N_9710);
nor U13952 (N_13952,N_11488,N_9585);
and U13953 (N_13953,N_10446,N_9204);
nor U13954 (N_13954,N_9731,N_11103);
nand U13955 (N_13955,N_9481,N_10792);
nand U13956 (N_13956,N_10146,N_9025);
nand U13957 (N_13957,N_9734,N_9195);
xor U13958 (N_13958,N_10521,N_9132);
or U13959 (N_13959,N_10185,N_10629);
nor U13960 (N_13960,N_11322,N_10149);
xor U13961 (N_13961,N_11523,N_9130);
and U13962 (N_13962,N_10386,N_11701);
nand U13963 (N_13963,N_11264,N_9152);
xnor U13964 (N_13964,N_9269,N_10425);
nor U13965 (N_13965,N_10347,N_10430);
and U13966 (N_13966,N_11638,N_9625);
xor U13967 (N_13967,N_11515,N_9356);
nand U13968 (N_13968,N_9536,N_10738);
or U13969 (N_13969,N_9411,N_9427);
and U13970 (N_13970,N_9792,N_11883);
xor U13971 (N_13971,N_9688,N_11508);
xnor U13972 (N_13972,N_10802,N_9836);
xor U13973 (N_13973,N_9478,N_10558);
nor U13974 (N_13974,N_9460,N_11228);
and U13975 (N_13975,N_10641,N_9578);
and U13976 (N_13976,N_11167,N_11420);
nand U13977 (N_13977,N_11478,N_10315);
nand U13978 (N_13978,N_9200,N_11878);
and U13979 (N_13979,N_11432,N_9480);
xor U13980 (N_13980,N_9173,N_11714);
nor U13981 (N_13981,N_11365,N_10869);
xor U13982 (N_13982,N_9815,N_11909);
nor U13983 (N_13983,N_9743,N_9197);
or U13984 (N_13984,N_9977,N_11106);
and U13985 (N_13985,N_11188,N_9642);
nand U13986 (N_13986,N_11162,N_9666);
or U13987 (N_13987,N_9233,N_11660);
nor U13988 (N_13988,N_9906,N_11260);
and U13989 (N_13989,N_10392,N_11737);
and U13990 (N_13990,N_10953,N_11374);
xnor U13991 (N_13991,N_11788,N_9363);
and U13992 (N_13992,N_10059,N_9672);
and U13993 (N_13993,N_11469,N_10706);
nand U13994 (N_13994,N_9814,N_11338);
nand U13995 (N_13995,N_11553,N_9189);
or U13996 (N_13996,N_11034,N_11232);
or U13997 (N_13997,N_9736,N_10371);
or U13998 (N_13998,N_10032,N_10461);
or U13999 (N_13999,N_11334,N_11739);
xnor U14000 (N_14000,N_9267,N_11807);
nor U14001 (N_14001,N_11374,N_10555);
and U14002 (N_14002,N_9283,N_11205);
nor U14003 (N_14003,N_11181,N_9159);
and U14004 (N_14004,N_10685,N_11372);
xor U14005 (N_14005,N_11328,N_9529);
or U14006 (N_14006,N_11684,N_10529);
nand U14007 (N_14007,N_11322,N_9471);
xor U14008 (N_14008,N_11544,N_11804);
nor U14009 (N_14009,N_10031,N_10907);
nor U14010 (N_14010,N_10637,N_9735);
nor U14011 (N_14011,N_9627,N_11506);
xnor U14012 (N_14012,N_9308,N_11003);
nor U14013 (N_14013,N_10082,N_10213);
nand U14014 (N_14014,N_11897,N_10157);
and U14015 (N_14015,N_10399,N_11536);
and U14016 (N_14016,N_10831,N_11553);
or U14017 (N_14017,N_11703,N_9112);
and U14018 (N_14018,N_9091,N_10075);
or U14019 (N_14019,N_9300,N_11860);
nor U14020 (N_14020,N_10146,N_9739);
nand U14021 (N_14021,N_9534,N_9488);
and U14022 (N_14022,N_11523,N_11210);
nand U14023 (N_14023,N_9347,N_11823);
xnor U14024 (N_14024,N_10164,N_9343);
nand U14025 (N_14025,N_9464,N_9438);
nand U14026 (N_14026,N_11333,N_11925);
or U14027 (N_14027,N_9155,N_10442);
nor U14028 (N_14028,N_9077,N_11017);
xor U14029 (N_14029,N_10043,N_10204);
xnor U14030 (N_14030,N_11619,N_9505);
nand U14031 (N_14031,N_9287,N_11384);
xnor U14032 (N_14032,N_10544,N_11392);
xnor U14033 (N_14033,N_10079,N_11206);
xor U14034 (N_14034,N_10918,N_10897);
nor U14035 (N_14035,N_9243,N_10976);
nor U14036 (N_14036,N_11758,N_10925);
xnor U14037 (N_14037,N_9010,N_9050);
and U14038 (N_14038,N_11033,N_10096);
and U14039 (N_14039,N_10706,N_9361);
and U14040 (N_14040,N_9762,N_11642);
nor U14041 (N_14041,N_11409,N_9261);
xnor U14042 (N_14042,N_9691,N_9626);
xnor U14043 (N_14043,N_10660,N_9204);
and U14044 (N_14044,N_11987,N_9899);
or U14045 (N_14045,N_10269,N_10000);
nand U14046 (N_14046,N_11379,N_11716);
nand U14047 (N_14047,N_11681,N_9985);
and U14048 (N_14048,N_10360,N_11257);
nand U14049 (N_14049,N_10610,N_11154);
or U14050 (N_14050,N_10500,N_11816);
or U14051 (N_14051,N_9632,N_10113);
xnor U14052 (N_14052,N_10977,N_10162);
and U14053 (N_14053,N_11980,N_9268);
or U14054 (N_14054,N_9861,N_9032);
nor U14055 (N_14055,N_10513,N_9955);
nand U14056 (N_14056,N_11773,N_10720);
nand U14057 (N_14057,N_10160,N_11102);
and U14058 (N_14058,N_11378,N_10400);
xnor U14059 (N_14059,N_9316,N_11626);
nand U14060 (N_14060,N_11967,N_10861);
nand U14061 (N_14061,N_11796,N_10750);
and U14062 (N_14062,N_10398,N_9512);
xnor U14063 (N_14063,N_9203,N_9353);
nor U14064 (N_14064,N_9051,N_11783);
or U14065 (N_14065,N_9793,N_11475);
nand U14066 (N_14066,N_9457,N_11670);
and U14067 (N_14067,N_11841,N_10733);
nand U14068 (N_14068,N_11457,N_10326);
xnor U14069 (N_14069,N_10597,N_10171);
nand U14070 (N_14070,N_9411,N_11396);
nor U14071 (N_14071,N_9893,N_11766);
nor U14072 (N_14072,N_10386,N_9194);
nand U14073 (N_14073,N_10982,N_9815);
xor U14074 (N_14074,N_9101,N_9963);
nand U14075 (N_14075,N_10912,N_10858);
nor U14076 (N_14076,N_10748,N_9591);
or U14077 (N_14077,N_10214,N_10301);
and U14078 (N_14078,N_11553,N_9965);
xor U14079 (N_14079,N_9812,N_10537);
xnor U14080 (N_14080,N_11751,N_9438);
xor U14081 (N_14081,N_10893,N_10584);
nor U14082 (N_14082,N_11712,N_11209);
and U14083 (N_14083,N_11610,N_11964);
or U14084 (N_14084,N_11743,N_11175);
xor U14085 (N_14085,N_9578,N_9781);
xor U14086 (N_14086,N_10416,N_9201);
nand U14087 (N_14087,N_11983,N_10126);
nand U14088 (N_14088,N_10538,N_9642);
or U14089 (N_14089,N_11967,N_9288);
nand U14090 (N_14090,N_10025,N_10150);
xor U14091 (N_14091,N_10671,N_9672);
or U14092 (N_14092,N_11983,N_9243);
nand U14093 (N_14093,N_10208,N_10271);
nand U14094 (N_14094,N_9358,N_10027);
xnor U14095 (N_14095,N_9455,N_9199);
nor U14096 (N_14096,N_10369,N_10966);
nand U14097 (N_14097,N_10980,N_11905);
or U14098 (N_14098,N_9493,N_9678);
and U14099 (N_14099,N_10553,N_10233);
nor U14100 (N_14100,N_10706,N_9715);
nand U14101 (N_14101,N_9908,N_9853);
nor U14102 (N_14102,N_11117,N_10885);
xor U14103 (N_14103,N_11583,N_9239);
xnor U14104 (N_14104,N_10668,N_11806);
nand U14105 (N_14105,N_11437,N_10902);
nand U14106 (N_14106,N_9587,N_11252);
and U14107 (N_14107,N_10037,N_10358);
xor U14108 (N_14108,N_11550,N_10193);
and U14109 (N_14109,N_10961,N_10557);
xnor U14110 (N_14110,N_11958,N_11023);
and U14111 (N_14111,N_11355,N_9093);
xnor U14112 (N_14112,N_10345,N_10461);
and U14113 (N_14113,N_10770,N_11458);
and U14114 (N_14114,N_10878,N_11920);
and U14115 (N_14115,N_9856,N_11491);
and U14116 (N_14116,N_10155,N_9100);
and U14117 (N_14117,N_9907,N_10174);
nor U14118 (N_14118,N_9317,N_11042);
nor U14119 (N_14119,N_10819,N_11681);
xnor U14120 (N_14120,N_11423,N_11219);
or U14121 (N_14121,N_11432,N_9400);
nand U14122 (N_14122,N_11949,N_10945);
nor U14123 (N_14123,N_11575,N_9870);
nor U14124 (N_14124,N_11690,N_10166);
nand U14125 (N_14125,N_9374,N_9593);
nor U14126 (N_14126,N_11795,N_10081);
and U14127 (N_14127,N_11794,N_11281);
and U14128 (N_14128,N_11689,N_11407);
and U14129 (N_14129,N_9935,N_9799);
nor U14130 (N_14130,N_9489,N_10344);
and U14131 (N_14131,N_11256,N_11862);
nand U14132 (N_14132,N_11757,N_11714);
and U14133 (N_14133,N_9211,N_10656);
or U14134 (N_14134,N_10848,N_11150);
nor U14135 (N_14135,N_11976,N_9158);
xor U14136 (N_14136,N_10358,N_10860);
nor U14137 (N_14137,N_11064,N_10615);
nand U14138 (N_14138,N_11579,N_11637);
or U14139 (N_14139,N_10729,N_10752);
and U14140 (N_14140,N_11300,N_10497);
xnor U14141 (N_14141,N_11234,N_11481);
nor U14142 (N_14142,N_9696,N_9543);
nand U14143 (N_14143,N_11472,N_10248);
nor U14144 (N_14144,N_11983,N_11762);
nand U14145 (N_14145,N_9672,N_11420);
and U14146 (N_14146,N_9682,N_9809);
and U14147 (N_14147,N_11710,N_10539);
nor U14148 (N_14148,N_9079,N_10327);
xnor U14149 (N_14149,N_11468,N_11704);
and U14150 (N_14150,N_10010,N_10304);
xnor U14151 (N_14151,N_9826,N_11803);
and U14152 (N_14152,N_9625,N_9286);
and U14153 (N_14153,N_11339,N_10930);
or U14154 (N_14154,N_9877,N_11856);
and U14155 (N_14155,N_10321,N_9858);
and U14156 (N_14156,N_9352,N_10489);
nor U14157 (N_14157,N_9890,N_10316);
nor U14158 (N_14158,N_9062,N_9885);
nor U14159 (N_14159,N_10633,N_9857);
and U14160 (N_14160,N_11238,N_9141);
nand U14161 (N_14161,N_11128,N_11487);
or U14162 (N_14162,N_9079,N_11439);
nand U14163 (N_14163,N_10803,N_10835);
nor U14164 (N_14164,N_10863,N_9849);
and U14165 (N_14165,N_10679,N_9406);
and U14166 (N_14166,N_10438,N_9922);
nand U14167 (N_14167,N_10927,N_11694);
or U14168 (N_14168,N_10635,N_11200);
nand U14169 (N_14169,N_9010,N_9665);
nor U14170 (N_14170,N_11486,N_11427);
and U14171 (N_14171,N_11761,N_11417);
nor U14172 (N_14172,N_10965,N_9322);
nor U14173 (N_14173,N_9186,N_9910);
or U14174 (N_14174,N_11782,N_9034);
nand U14175 (N_14175,N_11730,N_10580);
or U14176 (N_14176,N_9968,N_9194);
nand U14177 (N_14177,N_10751,N_10964);
nor U14178 (N_14178,N_11881,N_10762);
and U14179 (N_14179,N_10592,N_10242);
or U14180 (N_14180,N_10003,N_10774);
nand U14181 (N_14181,N_10733,N_9153);
nand U14182 (N_14182,N_9198,N_11887);
or U14183 (N_14183,N_11265,N_10863);
or U14184 (N_14184,N_11551,N_9837);
and U14185 (N_14185,N_10354,N_9608);
xor U14186 (N_14186,N_11507,N_11259);
nor U14187 (N_14187,N_11928,N_9626);
nor U14188 (N_14188,N_11385,N_9648);
xor U14189 (N_14189,N_11792,N_11455);
nor U14190 (N_14190,N_9326,N_11492);
or U14191 (N_14191,N_9599,N_10103);
nand U14192 (N_14192,N_11070,N_11705);
nor U14193 (N_14193,N_9405,N_11789);
nor U14194 (N_14194,N_10868,N_9804);
xnor U14195 (N_14195,N_11672,N_10757);
nor U14196 (N_14196,N_9889,N_11313);
xor U14197 (N_14197,N_10092,N_9532);
or U14198 (N_14198,N_9830,N_10746);
and U14199 (N_14199,N_11710,N_11274);
nor U14200 (N_14200,N_11502,N_11692);
and U14201 (N_14201,N_9011,N_9996);
xor U14202 (N_14202,N_9884,N_11482);
nor U14203 (N_14203,N_10357,N_9895);
or U14204 (N_14204,N_10414,N_11959);
and U14205 (N_14205,N_10828,N_9209);
and U14206 (N_14206,N_9702,N_10822);
nor U14207 (N_14207,N_9610,N_9051);
nand U14208 (N_14208,N_11019,N_11952);
and U14209 (N_14209,N_11350,N_9265);
nand U14210 (N_14210,N_10287,N_10352);
nor U14211 (N_14211,N_9159,N_9295);
or U14212 (N_14212,N_9710,N_10370);
nor U14213 (N_14213,N_9135,N_11426);
and U14214 (N_14214,N_10215,N_9635);
and U14215 (N_14215,N_9067,N_11500);
or U14216 (N_14216,N_9577,N_9985);
or U14217 (N_14217,N_10663,N_11815);
nor U14218 (N_14218,N_11206,N_11575);
xnor U14219 (N_14219,N_10942,N_11879);
nand U14220 (N_14220,N_10003,N_10054);
and U14221 (N_14221,N_11583,N_10783);
xor U14222 (N_14222,N_11721,N_10139);
nor U14223 (N_14223,N_11479,N_11990);
or U14224 (N_14224,N_10561,N_9334);
nor U14225 (N_14225,N_9391,N_9655);
nand U14226 (N_14226,N_9142,N_11801);
nand U14227 (N_14227,N_9836,N_9904);
and U14228 (N_14228,N_11619,N_10431);
or U14229 (N_14229,N_10275,N_11505);
and U14230 (N_14230,N_11075,N_10516);
nand U14231 (N_14231,N_10755,N_9989);
nand U14232 (N_14232,N_10120,N_9001);
nor U14233 (N_14233,N_10852,N_10463);
and U14234 (N_14234,N_9764,N_11294);
xnor U14235 (N_14235,N_9508,N_11450);
or U14236 (N_14236,N_10334,N_10489);
nand U14237 (N_14237,N_9239,N_10971);
nor U14238 (N_14238,N_10364,N_11825);
nor U14239 (N_14239,N_10692,N_10864);
nor U14240 (N_14240,N_10861,N_10705);
nand U14241 (N_14241,N_9012,N_9423);
nand U14242 (N_14242,N_11230,N_11143);
and U14243 (N_14243,N_11683,N_11178);
xor U14244 (N_14244,N_9177,N_9326);
nor U14245 (N_14245,N_10085,N_11980);
and U14246 (N_14246,N_10670,N_10633);
nor U14247 (N_14247,N_11746,N_11605);
xor U14248 (N_14248,N_9059,N_11375);
xnor U14249 (N_14249,N_9719,N_9325);
and U14250 (N_14250,N_11972,N_11952);
or U14251 (N_14251,N_9354,N_9164);
or U14252 (N_14252,N_9244,N_9289);
nand U14253 (N_14253,N_11948,N_11607);
or U14254 (N_14254,N_10202,N_11980);
and U14255 (N_14255,N_9658,N_10594);
nor U14256 (N_14256,N_10770,N_9770);
and U14257 (N_14257,N_10790,N_9136);
xnor U14258 (N_14258,N_11802,N_10860);
or U14259 (N_14259,N_9351,N_11045);
nor U14260 (N_14260,N_10951,N_11619);
nand U14261 (N_14261,N_9993,N_11127);
nor U14262 (N_14262,N_9840,N_10522);
xnor U14263 (N_14263,N_11445,N_11287);
xor U14264 (N_14264,N_11899,N_9424);
or U14265 (N_14265,N_10066,N_9061);
nor U14266 (N_14266,N_10401,N_11876);
and U14267 (N_14267,N_10659,N_11521);
or U14268 (N_14268,N_9742,N_11985);
nand U14269 (N_14269,N_11264,N_11785);
nor U14270 (N_14270,N_10637,N_11195);
and U14271 (N_14271,N_9672,N_11030);
xnor U14272 (N_14272,N_10658,N_9929);
nand U14273 (N_14273,N_10275,N_9624);
xnor U14274 (N_14274,N_11657,N_10150);
and U14275 (N_14275,N_10544,N_9091);
and U14276 (N_14276,N_11786,N_9406);
nor U14277 (N_14277,N_10864,N_11062);
and U14278 (N_14278,N_10767,N_11013);
and U14279 (N_14279,N_11825,N_9097);
xnor U14280 (N_14280,N_9912,N_9209);
or U14281 (N_14281,N_11024,N_9189);
nand U14282 (N_14282,N_10597,N_11318);
nor U14283 (N_14283,N_9544,N_10283);
nor U14284 (N_14284,N_9953,N_10966);
or U14285 (N_14285,N_10475,N_9630);
xor U14286 (N_14286,N_10786,N_9260);
xor U14287 (N_14287,N_11674,N_11987);
or U14288 (N_14288,N_10397,N_11453);
and U14289 (N_14289,N_9488,N_11230);
nand U14290 (N_14290,N_10870,N_9486);
nand U14291 (N_14291,N_11974,N_11200);
and U14292 (N_14292,N_10953,N_11914);
xor U14293 (N_14293,N_10370,N_11534);
nand U14294 (N_14294,N_9929,N_11994);
nand U14295 (N_14295,N_10737,N_10805);
nor U14296 (N_14296,N_10043,N_10001);
or U14297 (N_14297,N_10910,N_10533);
nand U14298 (N_14298,N_10151,N_9968);
or U14299 (N_14299,N_9221,N_11326);
and U14300 (N_14300,N_10776,N_11083);
nor U14301 (N_14301,N_10564,N_11304);
nand U14302 (N_14302,N_10260,N_11880);
xor U14303 (N_14303,N_11813,N_9789);
and U14304 (N_14304,N_9871,N_11298);
xnor U14305 (N_14305,N_10363,N_9000);
xnor U14306 (N_14306,N_11816,N_10547);
xor U14307 (N_14307,N_11738,N_9376);
nor U14308 (N_14308,N_10329,N_11116);
and U14309 (N_14309,N_9660,N_10648);
and U14310 (N_14310,N_10051,N_11345);
and U14311 (N_14311,N_9841,N_11478);
nand U14312 (N_14312,N_9921,N_9125);
nand U14313 (N_14313,N_11754,N_10584);
nor U14314 (N_14314,N_11507,N_9549);
and U14315 (N_14315,N_9490,N_9600);
xor U14316 (N_14316,N_10759,N_9485);
and U14317 (N_14317,N_11045,N_9319);
nand U14318 (N_14318,N_10001,N_9996);
nor U14319 (N_14319,N_11489,N_10695);
nand U14320 (N_14320,N_10716,N_11068);
and U14321 (N_14321,N_9245,N_11564);
xor U14322 (N_14322,N_10826,N_11500);
xor U14323 (N_14323,N_9603,N_10867);
and U14324 (N_14324,N_11956,N_10965);
or U14325 (N_14325,N_9361,N_11391);
or U14326 (N_14326,N_11567,N_11296);
xor U14327 (N_14327,N_10169,N_9512);
and U14328 (N_14328,N_11882,N_9412);
xor U14329 (N_14329,N_10542,N_10975);
or U14330 (N_14330,N_9337,N_11741);
xor U14331 (N_14331,N_9031,N_9775);
nand U14332 (N_14332,N_10115,N_10391);
and U14333 (N_14333,N_11408,N_9712);
nand U14334 (N_14334,N_9541,N_9386);
and U14335 (N_14335,N_10403,N_11863);
nor U14336 (N_14336,N_11399,N_10305);
or U14337 (N_14337,N_9874,N_9610);
or U14338 (N_14338,N_11880,N_11086);
and U14339 (N_14339,N_11910,N_10332);
and U14340 (N_14340,N_9896,N_10780);
nor U14341 (N_14341,N_9332,N_10526);
nor U14342 (N_14342,N_10275,N_9822);
xor U14343 (N_14343,N_9636,N_10789);
nor U14344 (N_14344,N_10692,N_9592);
nand U14345 (N_14345,N_9465,N_9483);
xnor U14346 (N_14346,N_9183,N_10967);
xnor U14347 (N_14347,N_9326,N_11041);
nand U14348 (N_14348,N_11839,N_10887);
and U14349 (N_14349,N_9248,N_9093);
xnor U14350 (N_14350,N_9458,N_9372);
or U14351 (N_14351,N_11536,N_9023);
or U14352 (N_14352,N_9795,N_9592);
or U14353 (N_14353,N_9189,N_11638);
nand U14354 (N_14354,N_10739,N_10431);
xnor U14355 (N_14355,N_11208,N_10019);
and U14356 (N_14356,N_11973,N_10512);
nand U14357 (N_14357,N_9439,N_9576);
xor U14358 (N_14358,N_11790,N_11815);
nand U14359 (N_14359,N_9254,N_11101);
nand U14360 (N_14360,N_9264,N_9631);
xnor U14361 (N_14361,N_9002,N_10238);
and U14362 (N_14362,N_11332,N_9811);
or U14363 (N_14363,N_10284,N_9959);
xor U14364 (N_14364,N_11870,N_9959);
and U14365 (N_14365,N_10930,N_10615);
or U14366 (N_14366,N_10805,N_11086);
nand U14367 (N_14367,N_11296,N_11255);
and U14368 (N_14368,N_11015,N_9666);
nor U14369 (N_14369,N_10240,N_10415);
nor U14370 (N_14370,N_11732,N_11005);
nor U14371 (N_14371,N_11057,N_10167);
nor U14372 (N_14372,N_11521,N_11490);
nor U14373 (N_14373,N_10192,N_11787);
and U14374 (N_14374,N_9592,N_10942);
and U14375 (N_14375,N_10603,N_10630);
xor U14376 (N_14376,N_9938,N_11481);
nor U14377 (N_14377,N_11190,N_11064);
xor U14378 (N_14378,N_9120,N_9136);
xor U14379 (N_14379,N_10130,N_11320);
xnor U14380 (N_14380,N_10751,N_9302);
nand U14381 (N_14381,N_11697,N_9984);
and U14382 (N_14382,N_11027,N_11034);
nand U14383 (N_14383,N_11936,N_9239);
xor U14384 (N_14384,N_10735,N_11281);
and U14385 (N_14385,N_10593,N_9616);
nand U14386 (N_14386,N_11838,N_10409);
or U14387 (N_14387,N_11925,N_9157);
and U14388 (N_14388,N_9449,N_10672);
xnor U14389 (N_14389,N_11517,N_9218);
or U14390 (N_14390,N_9542,N_11709);
nand U14391 (N_14391,N_11567,N_11764);
or U14392 (N_14392,N_10053,N_10406);
and U14393 (N_14393,N_9139,N_9004);
or U14394 (N_14394,N_10012,N_9843);
nor U14395 (N_14395,N_9896,N_11967);
xnor U14396 (N_14396,N_9358,N_11251);
nor U14397 (N_14397,N_11941,N_11580);
or U14398 (N_14398,N_9045,N_10219);
xnor U14399 (N_14399,N_11722,N_10677);
nand U14400 (N_14400,N_9486,N_10084);
and U14401 (N_14401,N_11237,N_11658);
or U14402 (N_14402,N_10315,N_11518);
nand U14403 (N_14403,N_10566,N_11759);
nand U14404 (N_14404,N_9988,N_10393);
or U14405 (N_14405,N_11109,N_11771);
xnor U14406 (N_14406,N_10341,N_11938);
or U14407 (N_14407,N_9521,N_11984);
nand U14408 (N_14408,N_9661,N_9969);
or U14409 (N_14409,N_10019,N_10231);
nand U14410 (N_14410,N_9041,N_10811);
nand U14411 (N_14411,N_10978,N_11329);
or U14412 (N_14412,N_10498,N_10017);
nand U14413 (N_14413,N_10397,N_10439);
or U14414 (N_14414,N_10081,N_11466);
nand U14415 (N_14415,N_9199,N_11156);
nor U14416 (N_14416,N_10112,N_11196);
and U14417 (N_14417,N_11688,N_11631);
xor U14418 (N_14418,N_9902,N_10193);
nor U14419 (N_14419,N_10804,N_9145);
and U14420 (N_14420,N_11497,N_9891);
nand U14421 (N_14421,N_11461,N_11803);
and U14422 (N_14422,N_11025,N_9542);
nor U14423 (N_14423,N_11135,N_11026);
and U14424 (N_14424,N_11198,N_11603);
or U14425 (N_14425,N_9636,N_10337);
nand U14426 (N_14426,N_10918,N_9021);
xnor U14427 (N_14427,N_10881,N_10411);
nand U14428 (N_14428,N_10099,N_11161);
and U14429 (N_14429,N_11931,N_10524);
nor U14430 (N_14430,N_11974,N_11404);
and U14431 (N_14431,N_10171,N_10411);
nor U14432 (N_14432,N_9069,N_10960);
nor U14433 (N_14433,N_11082,N_10786);
or U14434 (N_14434,N_11819,N_10444);
nor U14435 (N_14435,N_10626,N_11597);
or U14436 (N_14436,N_9378,N_10738);
nand U14437 (N_14437,N_11274,N_10478);
and U14438 (N_14438,N_11344,N_11267);
nor U14439 (N_14439,N_10427,N_11337);
or U14440 (N_14440,N_10664,N_9998);
nor U14441 (N_14441,N_9411,N_9321);
and U14442 (N_14442,N_10498,N_10251);
and U14443 (N_14443,N_10251,N_11797);
or U14444 (N_14444,N_11575,N_9543);
nor U14445 (N_14445,N_10137,N_9899);
and U14446 (N_14446,N_9262,N_10959);
nor U14447 (N_14447,N_9288,N_9957);
nor U14448 (N_14448,N_10465,N_10767);
nor U14449 (N_14449,N_9471,N_9618);
or U14450 (N_14450,N_9505,N_10447);
nor U14451 (N_14451,N_11129,N_10314);
xor U14452 (N_14452,N_11700,N_9369);
or U14453 (N_14453,N_10419,N_11334);
or U14454 (N_14454,N_10804,N_9341);
and U14455 (N_14455,N_9485,N_11377);
and U14456 (N_14456,N_10204,N_9565);
nor U14457 (N_14457,N_10006,N_10574);
and U14458 (N_14458,N_9531,N_10216);
nand U14459 (N_14459,N_11266,N_10111);
or U14460 (N_14460,N_10125,N_10357);
nor U14461 (N_14461,N_11531,N_11787);
xnor U14462 (N_14462,N_10913,N_10103);
nand U14463 (N_14463,N_10868,N_9000);
xnor U14464 (N_14464,N_10913,N_11737);
nor U14465 (N_14465,N_11007,N_10995);
nor U14466 (N_14466,N_10059,N_11102);
and U14467 (N_14467,N_10429,N_10786);
nor U14468 (N_14468,N_10609,N_10252);
xor U14469 (N_14469,N_11175,N_11647);
nand U14470 (N_14470,N_11790,N_9207);
nand U14471 (N_14471,N_10453,N_9038);
nand U14472 (N_14472,N_11539,N_10631);
nand U14473 (N_14473,N_9307,N_10819);
nand U14474 (N_14474,N_11321,N_10821);
nand U14475 (N_14475,N_9205,N_11214);
and U14476 (N_14476,N_9607,N_10070);
and U14477 (N_14477,N_9540,N_9427);
or U14478 (N_14478,N_9785,N_10561);
nand U14479 (N_14479,N_11960,N_9568);
nand U14480 (N_14480,N_10972,N_9273);
and U14481 (N_14481,N_10099,N_10076);
nand U14482 (N_14482,N_9302,N_9145);
nand U14483 (N_14483,N_10490,N_10709);
or U14484 (N_14484,N_10963,N_10662);
nor U14485 (N_14485,N_9914,N_10733);
and U14486 (N_14486,N_11214,N_9316);
or U14487 (N_14487,N_11290,N_11025);
and U14488 (N_14488,N_11555,N_9829);
nor U14489 (N_14489,N_9900,N_9502);
xnor U14490 (N_14490,N_10349,N_10697);
or U14491 (N_14491,N_9782,N_10170);
and U14492 (N_14492,N_11428,N_9275);
or U14493 (N_14493,N_9072,N_10483);
and U14494 (N_14494,N_11344,N_11770);
or U14495 (N_14495,N_11877,N_11467);
xnor U14496 (N_14496,N_11962,N_11024);
xor U14497 (N_14497,N_9736,N_10027);
xnor U14498 (N_14498,N_11443,N_10384);
or U14499 (N_14499,N_9241,N_10597);
or U14500 (N_14500,N_11203,N_10213);
or U14501 (N_14501,N_11327,N_9938);
nor U14502 (N_14502,N_10432,N_9202);
xnor U14503 (N_14503,N_11629,N_11640);
nand U14504 (N_14504,N_9357,N_9771);
xor U14505 (N_14505,N_10551,N_10726);
nand U14506 (N_14506,N_11764,N_11164);
and U14507 (N_14507,N_10403,N_11056);
nor U14508 (N_14508,N_9535,N_10786);
nand U14509 (N_14509,N_9920,N_11657);
and U14510 (N_14510,N_9541,N_11115);
xor U14511 (N_14511,N_10389,N_11394);
nand U14512 (N_14512,N_11540,N_10521);
nand U14513 (N_14513,N_10577,N_10726);
nor U14514 (N_14514,N_11323,N_9682);
or U14515 (N_14515,N_10911,N_10264);
nor U14516 (N_14516,N_11125,N_11316);
nand U14517 (N_14517,N_9305,N_9956);
or U14518 (N_14518,N_11009,N_9718);
nand U14519 (N_14519,N_11354,N_10337);
and U14520 (N_14520,N_9012,N_11213);
or U14521 (N_14521,N_10812,N_11281);
nand U14522 (N_14522,N_11266,N_10952);
and U14523 (N_14523,N_9292,N_11443);
nand U14524 (N_14524,N_9064,N_9676);
and U14525 (N_14525,N_10051,N_10324);
nor U14526 (N_14526,N_11952,N_9834);
xnor U14527 (N_14527,N_9574,N_9057);
xnor U14528 (N_14528,N_11815,N_11792);
or U14529 (N_14529,N_9721,N_11326);
and U14530 (N_14530,N_9561,N_9030);
or U14531 (N_14531,N_9652,N_11843);
or U14532 (N_14532,N_11020,N_11503);
or U14533 (N_14533,N_11730,N_11071);
xnor U14534 (N_14534,N_11198,N_9517);
and U14535 (N_14535,N_11706,N_9617);
or U14536 (N_14536,N_9310,N_10651);
or U14537 (N_14537,N_10526,N_10557);
xor U14538 (N_14538,N_11770,N_11346);
nor U14539 (N_14539,N_11840,N_11225);
and U14540 (N_14540,N_11863,N_10741);
or U14541 (N_14541,N_11662,N_10793);
xor U14542 (N_14542,N_9872,N_11988);
and U14543 (N_14543,N_9554,N_9379);
or U14544 (N_14544,N_9639,N_9913);
xor U14545 (N_14545,N_10841,N_9235);
and U14546 (N_14546,N_9658,N_9166);
nor U14547 (N_14547,N_9140,N_11678);
or U14548 (N_14548,N_10048,N_11447);
nand U14549 (N_14549,N_11086,N_11362);
or U14550 (N_14550,N_10889,N_9614);
or U14551 (N_14551,N_9335,N_11760);
or U14552 (N_14552,N_11110,N_9333);
or U14553 (N_14553,N_11196,N_9280);
xor U14554 (N_14554,N_9765,N_10473);
xnor U14555 (N_14555,N_9626,N_9531);
or U14556 (N_14556,N_9674,N_10284);
and U14557 (N_14557,N_11209,N_10545);
nand U14558 (N_14558,N_9344,N_11591);
and U14559 (N_14559,N_9171,N_9983);
nand U14560 (N_14560,N_10922,N_10359);
nor U14561 (N_14561,N_10747,N_9621);
xor U14562 (N_14562,N_9858,N_11247);
xor U14563 (N_14563,N_10972,N_11183);
xnor U14564 (N_14564,N_9881,N_11620);
nor U14565 (N_14565,N_10842,N_9193);
and U14566 (N_14566,N_11585,N_11260);
and U14567 (N_14567,N_9817,N_11748);
nor U14568 (N_14568,N_11937,N_11685);
nor U14569 (N_14569,N_9509,N_9351);
and U14570 (N_14570,N_9780,N_11012);
xor U14571 (N_14571,N_10246,N_9757);
or U14572 (N_14572,N_9495,N_9939);
and U14573 (N_14573,N_11668,N_10811);
or U14574 (N_14574,N_9321,N_11463);
and U14575 (N_14575,N_11341,N_11678);
nand U14576 (N_14576,N_10989,N_9508);
or U14577 (N_14577,N_11938,N_9760);
xnor U14578 (N_14578,N_11408,N_9535);
and U14579 (N_14579,N_9085,N_10156);
nor U14580 (N_14580,N_9991,N_11607);
xnor U14581 (N_14581,N_9091,N_9375);
and U14582 (N_14582,N_9052,N_9233);
xor U14583 (N_14583,N_10325,N_9747);
nor U14584 (N_14584,N_9322,N_10217);
or U14585 (N_14585,N_11544,N_10061);
or U14586 (N_14586,N_9101,N_11642);
and U14587 (N_14587,N_10765,N_9613);
nand U14588 (N_14588,N_9771,N_10757);
nand U14589 (N_14589,N_11935,N_9326);
nor U14590 (N_14590,N_11005,N_11416);
nor U14591 (N_14591,N_11779,N_9980);
xnor U14592 (N_14592,N_9310,N_10528);
and U14593 (N_14593,N_9268,N_9827);
or U14594 (N_14594,N_9631,N_9598);
and U14595 (N_14595,N_9654,N_11766);
and U14596 (N_14596,N_10874,N_11086);
or U14597 (N_14597,N_9007,N_11301);
xor U14598 (N_14598,N_11246,N_10823);
xnor U14599 (N_14599,N_11078,N_11113);
nor U14600 (N_14600,N_11666,N_11516);
nand U14601 (N_14601,N_11531,N_11848);
nor U14602 (N_14602,N_9724,N_11159);
xnor U14603 (N_14603,N_11170,N_10942);
or U14604 (N_14604,N_9041,N_11386);
nand U14605 (N_14605,N_11791,N_9390);
nand U14606 (N_14606,N_9785,N_11788);
and U14607 (N_14607,N_10304,N_9253);
and U14608 (N_14608,N_10627,N_9532);
or U14609 (N_14609,N_11301,N_9912);
nor U14610 (N_14610,N_9260,N_10389);
and U14611 (N_14611,N_10890,N_10367);
xnor U14612 (N_14612,N_9118,N_11694);
or U14613 (N_14613,N_11714,N_9845);
xor U14614 (N_14614,N_9440,N_10536);
or U14615 (N_14615,N_9218,N_10604);
nand U14616 (N_14616,N_10984,N_10002);
nand U14617 (N_14617,N_9506,N_10527);
or U14618 (N_14618,N_11699,N_9792);
and U14619 (N_14619,N_11497,N_11047);
and U14620 (N_14620,N_11117,N_11087);
xor U14621 (N_14621,N_9926,N_9382);
nand U14622 (N_14622,N_10581,N_9905);
or U14623 (N_14623,N_10937,N_10512);
and U14624 (N_14624,N_10806,N_9647);
and U14625 (N_14625,N_9189,N_10610);
or U14626 (N_14626,N_11558,N_11093);
nor U14627 (N_14627,N_10418,N_9426);
and U14628 (N_14628,N_10361,N_10005);
or U14629 (N_14629,N_10850,N_11273);
and U14630 (N_14630,N_11690,N_10498);
xor U14631 (N_14631,N_10260,N_9654);
and U14632 (N_14632,N_11078,N_10576);
nor U14633 (N_14633,N_10862,N_11899);
nor U14634 (N_14634,N_9119,N_9979);
nor U14635 (N_14635,N_9390,N_11119);
xnor U14636 (N_14636,N_9935,N_11250);
nor U14637 (N_14637,N_9646,N_10505);
nor U14638 (N_14638,N_11200,N_10185);
nand U14639 (N_14639,N_9056,N_10714);
and U14640 (N_14640,N_9642,N_10928);
nor U14641 (N_14641,N_9325,N_9404);
or U14642 (N_14642,N_10119,N_10974);
xnor U14643 (N_14643,N_11452,N_10507);
or U14644 (N_14644,N_9945,N_10943);
nand U14645 (N_14645,N_11470,N_11950);
nor U14646 (N_14646,N_9843,N_11038);
or U14647 (N_14647,N_11122,N_10941);
or U14648 (N_14648,N_11935,N_10660);
nor U14649 (N_14649,N_9460,N_10695);
nand U14650 (N_14650,N_11472,N_9883);
and U14651 (N_14651,N_9220,N_10634);
or U14652 (N_14652,N_11413,N_10647);
and U14653 (N_14653,N_9071,N_11191);
nor U14654 (N_14654,N_11736,N_11237);
xnor U14655 (N_14655,N_11858,N_11291);
and U14656 (N_14656,N_11785,N_10274);
and U14657 (N_14657,N_9567,N_11583);
nor U14658 (N_14658,N_9731,N_11661);
and U14659 (N_14659,N_9339,N_9021);
or U14660 (N_14660,N_9497,N_10624);
nor U14661 (N_14661,N_10850,N_9370);
nor U14662 (N_14662,N_11815,N_11668);
or U14663 (N_14663,N_11356,N_11583);
nor U14664 (N_14664,N_9470,N_9537);
and U14665 (N_14665,N_9754,N_10001);
nand U14666 (N_14666,N_10096,N_11378);
nand U14667 (N_14667,N_10986,N_10763);
xor U14668 (N_14668,N_9203,N_10000);
xor U14669 (N_14669,N_10622,N_10924);
or U14670 (N_14670,N_9581,N_11268);
nand U14671 (N_14671,N_11669,N_10504);
nand U14672 (N_14672,N_11013,N_11892);
xnor U14673 (N_14673,N_11844,N_10124);
or U14674 (N_14674,N_11600,N_10830);
nand U14675 (N_14675,N_10477,N_9947);
and U14676 (N_14676,N_10004,N_9532);
or U14677 (N_14677,N_10701,N_11412);
and U14678 (N_14678,N_10398,N_10092);
nor U14679 (N_14679,N_10125,N_11156);
and U14680 (N_14680,N_9168,N_9928);
xnor U14681 (N_14681,N_9379,N_10145);
xor U14682 (N_14682,N_10136,N_9645);
nand U14683 (N_14683,N_9001,N_9354);
nand U14684 (N_14684,N_11763,N_11190);
xor U14685 (N_14685,N_9060,N_11965);
or U14686 (N_14686,N_9731,N_11269);
or U14687 (N_14687,N_9545,N_10594);
nor U14688 (N_14688,N_9444,N_9561);
and U14689 (N_14689,N_11676,N_10702);
and U14690 (N_14690,N_11041,N_10142);
nand U14691 (N_14691,N_9565,N_9070);
or U14692 (N_14692,N_11065,N_11026);
xnor U14693 (N_14693,N_9884,N_11918);
nor U14694 (N_14694,N_9432,N_11622);
or U14695 (N_14695,N_9992,N_11962);
nor U14696 (N_14696,N_10031,N_11209);
xnor U14697 (N_14697,N_10433,N_11612);
xnor U14698 (N_14698,N_10497,N_11947);
or U14699 (N_14699,N_10301,N_10804);
nand U14700 (N_14700,N_10586,N_11334);
nor U14701 (N_14701,N_9674,N_10680);
nor U14702 (N_14702,N_11399,N_10213);
nor U14703 (N_14703,N_11731,N_10819);
and U14704 (N_14704,N_10064,N_10798);
nor U14705 (N_14705,N_11743,N_9713);
xor U14706 (N_14706,N_10452,N_10049);
xnor U14707 (N_14707,N_9884,N_10164);
xor U14708 (N_14708,N_10949,N_11740);
xor U14709 (N_14709,N_11080,N_9267);
nor U14710 (N_14710,N_9917,N_11024);
and U14711 (N_14711,N_9345,N_9675);
nand U14712 (N_14712,N_11191,N_11659);
xor U14713 (N_14713,N_11670,N_9009);
or U14714 (N_14714,N_10157,N_10958);
xor U14715 (N_14715,N_9296,N_9083);
and U14716 (N_14716,N_9760,N_11989);
nor U14717 (N_14717,N_10254,N_10347);
and U14718 (N_14718,N_10120,N_11516);
nor U14719 (N_14719,N_9763,N_11295);
nor U14720 (N_14720,N_11865,N_9697);
or U14721 (N_14721,N_9486,N_9234);
nor U14722 (N_14722,N_10061,N_10754);
nand U14723 (N_14723,N_10883,N_9355);
and U14724 (N_14724,N_11419,N_10786);
and U14725 (N_14725,N_10183,N_10182);
nand U14726 (N_14726,N_11267,N_9195);
or U14727 (N_14727,N_9380,N_9299);
xnor U14728 (N_14728,N_10223,N_11173);
xor U14729 (N_14729,N_11578,N_10470);
nand U14730 (N_14730,N_9329,N_11468);
nand U14731 (N_14731,N_9633,N_11835);
or U14732 (N_14732,N_10895,N_10811);
xnor U14733 (N_14733,N_10094,N_9435);
xnor U14734 (N_14734,N_11588,N_10999);
xor U14735 (N_14735,N_11329,N_9615);
nand U14736 (N_14736,N_9183,N_11914);
nand U14737 (N_14737,N_9458,N_10658);
or U14738 (N_14738,N_11314,N_10692);
and U14739 (N_14739,N_11845,N_10234);
or U14740 (N_14740,N_9435,N_10710);
xnor U14741 (N_14741,N_11015,N_11071);
nor U14742 (N_14742,N_9388,N_11446);
or U14743 (N_14743,N_11958,N_9059);
or U14744 (N_14744,N_9571,N_9704);
or U14745 (N_14745,N_11535,N_10140);
nand U14746 (N_14746,N_9428,N_9735);
nor U14747 (N_14747,N_11849,N_9759);
or U14748 (N_14748,N_10434,N_9055);
nor U14749 (N_14749,N_10934,N_10420);
or U14750 (N_14750,N_11439,N_11675);
nor U14751 (N_14751,N_9496,N_11612);
or U14752 (N_14752,N_9011,N_9534);
and U14753 (N_14753,N_9118,N_9066);
or U14754 (N_14754,N_9892,N_9459);
and U14755 (N_14755,N_10990,N_9933);
and U14756 (N_14756,N_10376,N_10973);
nor U14757 (N_14757,N_11717,N_9476);
and U14758 (N_14758,N_11498,N_11488);
or U14759 (N_14759,N_10907,N_9153);
and U14760 (N_14760,N_11695,N_9692);
nand U14761 (N_14761,N_11025,N_10135);
nand U14762 (N_14762,N_10064,N_9460);
xnor U14763 (N_14763,N_9267,N_10132);
and U14764 (N_14764,N_11160,N_10814);
or U14765 (N_14765,N_10670,N_9311);
nand U14766 (N_14766,N_10208,N_10326);
nor U14767 (N_14767,N_10033,N_11718);
xnor U14768 (N_14768,N_9485,N_9723);
or U14769 (N_14769,N_10802,N_10034);
nand U14770 (N_14770,N_11303,N_10804);
xor U14771 (N_14771,N_9494,N_9401);
or U14772 (N_14772,N_9837,N_11477);
or U14773 (N_14773,N_9868,N_11714);
or U14774 (N_14774,N_11735,N_9492);
or U14775 (N_14775,N_9867,N_11726);
or U14776 (N_14776,N_10342,N_9475);
nor U14777 (N_14777,N_11418,N_10008);
nand U14778 (N_14778,N_10277,N_9073);
xor U14779 (N_14779,N_10712,N_11826);
nand U14780 (N_14780,N_9584,N_9335);
or U14781 (N_14781,N_10529,N_11560);
or U14782 (N_14782,N_10437,N_9685);
and U14783 (N_14783,N_11547,N_11961);
nand U14784 (N_14784,N_10686,N_9242);
nand U14785 (N_14785,N_10168,N_10625);
or U14786 (N_14786,N_9530,N_11725);
nor U14787 (N_14787,N_10346,N_9481);
nand U14788 (N_14788,N_9305,N_10543);
nor U14789 (N_14789,N_10367,N_9109);
and U14790 (N_14790,N_10132,N_9537);
or U14791 (N_14791,N_11563,N_10505);
nand U14792 (N_14792,N_10378,N_9154);
nand U14793 (N_14793,N_10438,N_10566);
xnor U14794 (N_14794,N_9817,N_9972);
xor U14795 (N_14795,N_9531,N_10188);
or U14796 (N_14796,N_9195,N_11814);
nor U14797 (N_14797,N_10807,N_11358);
or U14798 (N_14798,N_10553,N_9125);
xnor U14799 (N_14799,N_10470,N_10722);
or U14800 (N_14800,N_9924,N_11023);
and U14801 (N_14801,N_9291,N_11340);
or U14802 (N_14802,N_10319,N_9419);
nor U14803 (N_14803,N_9929,N_9748);
xor U14804 (N_14804,N_10915,N_11248);
nor U14805 (N_14805,N_11181,N_9689);
nor U14806 (N_14806,N_11521,N_10376);
or U14807 (N_14807,N_10383,N_11416);
nand U14808 (N_14808,N_11333,N_11145);
xnor U14809 (N_14809,N_11783,N_10475);
xnor U14810 (N_14810,N_11256,N_10885);
xor U14811 (N_14811,N_9971,N_9243);
nor U14812 (N_14812,N_10365,N_9730);
and U14813 (N_14813,N_11990,N_9228);
nor U14814 (N_14814,N_9920,N_9368);
nand U14815 (N_14815,N_10201,N_10885);
xor U14816 (N_14816,N_9785,N_11579);
or U14817 (N_14817,N_10735,N_11823);
xor U14818 (N_14818,N_10755,N_11426);
and U14819 (N_14819,N_11287,N_10851);
nand U14820 (N_14820,N_9958,N_10217);
and U14821 (N_14821,N_9367,N_10563);
xnor U14822 (N_14822,N_11492,N_11835);
xnor U14823 (N_14823,N_10263,N_11421);
nand U14824 (N_14824,N_9709,N_11283);
xor U14825 (N_14825,N_10178,N_9997);
xnor U14826 (N_14826,N_10835,N_11036);
xor U14827 (N_14827,N_9284,N_10489);
or U14828 (N_14828,N_9325,N_10164);
or U14829 (N_14829,N_10990,N_11351);
nand U14830 (N_14830,N_9328,N_10774);
and U14831 (N_14831,N_10111,N_11318);
or U14832 (N_14832,N_10219,N_11846);
or U14833 (N_14833,N_11423,N_10018);
nand U14834 (N_14834,N_10991,N_11083);
or U14835 (N_14835,N_9909,N_11474);
xnor U14836 (N_14836,N_11553,N_11683);
nor U14837 (N_14837,N_11931,N_10964);
and U14838 (N_14838,N_11929,N_10653);
and U14839 (N_14839,N_10334,N_10299);
or U14840 (N_14840,N_11464,N_11001);
nand U14841 (N_14841,N_11587,N_9701);
xor U14842 (N_14842,N_11031,N_9243);
nand U14843 (N_14843,N_9735,N_10728);
xnor U14844 (N_14844,N_11155,N_11366);
nor U14845 (N_14845,N_11161,N_9223);
or U14846 (N_14846,N_11439,N_11129);
nor U14847 (N_14847,N_10745,N_9893);
nand U14848 (N_14848,N_11802,N_9974);
nor U14849 (N_14849,N_11951,N_11953);
nand U14850 (N_14850,N_10874,N_11815);
nand U14851 (N_14851,N_9278,N_9128);
nand U14852 (N_14852,N_10695,N_10289);
nand U14853 (N_14853,N_11335,N_10121);
and U14854 (N_14854,N_10247,N_11841);
and U14855 (N_14855,N_10806,N_10184);
and U14856 (N_14856,N_11952,N_9000);
and U14857 (N_14857,N_11492,N_10271);
or U14858 (N_14858,N_11178,N_10321);
nor U14859 (N_14859,N_11108,N_11471);
nor U14860 (N_14860,N_9385,N_10204);
nor U14861 (N_14861,N_10095,N_11381);
and U14862 (N_14862,N_10499,N_9767);
nand U14863 (N_14863,N_9878,N_10547);
nor U14864 (N_14864,N_9192,N_11585);
xor U14865 (N_14865,N_10429,N_11885);
nand U14866 (N_14866,N_10943,N_11785);
or U14867 (N_14867,N_10514,N_10115);
or U14868 (N_14868,N_9508,N_10790);
or U14869 (N_14869,N_10936,N_9225);
xnor U14870 (N_14870,N_11392,N_10313);
or U14871 (N_14871,N_9464,N_10308);
or U14872 (N_14872,N_11830,N_9360);
nand U14873 (N_14873,N_10576,N_9881);
nor U14874 (N_14874,N_11109,N_11017);
nor U14875 (N_14875,N_10331,N_10464);
nor U14876 (N_14876,N_10774,N_10659);
nand U14877 (N_14877,N_11056,N_9907);
or U14878 (N_14878,N_11791,N_10928);
and U14879 (N_14879,N_11243,N_9539);
xor U14880 (N_14880,N_10549,N_11391);
and U14881 (N_14881,N_10183,N_9422);
or U14882 (N_14882,N_9295,N_9130);
and U14883 (N_14883,N_11920,N_11814);
and U14884 (N_14884,N_10745,N_10292);
nor U14885 (N_14885,N_10954,N_10480);
nor U14886 (N_14886,N_10109,N_10657);
nor U14887 (N_14887,N_9827,N_11473);
nand U14888 (N_14888,N_9374,N_11284);
xnor U14889 (N_14889,N_11017,N_10700);
nand U14890 (N_14890,N_10633,N_10269);
and U14891 (N_14891,N_11011,N_11798);
or U14892 (N_14892,N_11037,N_10735);
and U14893 (N_14893,N_9562,N_9699);
and U14894 (N_14894,N_9716,N_11369);
xor U14895 (N_14895,N_10338,N_9125);
and U14896 (N_14896,N_10697,N_9926);
nor U14897 (N_14897,N_10600,N_11534);
xnor U14898 (N_14898,N_9121,N_9734);
xor U14899 (N_14899,N_11025,N_10976);
or U14900 (N_14900,N_10859,N_11428);
xnor U14901 (N_14901,N_10843,N_9111);
and U14902 (N_14902,N_9005,N_10940);
nand U14903 (N_14903,N_11235,N_11623);
or U14904 (N_14904,N_10945,N_11888);
nand U14905 (N_14905,N_9216,N_10944);
or U14906 (N_14906,N_9420,N_9797);
nand U14907 (N_14907,N_11227,N_11083);
nor U14908 (N_14908,N_10015,N_11348);
and U14909 (N_14909,N_10997,N_10642);
or U14910 (N_14910,N_9551,N_9658);
nor U14911 (N_14911,N_10037,N_11048);
or U14912 (N_14912,N_11598,N_10472);
nor U14913 (N_14913,N_10118,N_11255);
xor U14914 (N_14914,N_10410,N_11481);
nand U14915 (N_14915,N_10714,N_11052);
nor U14916 (N_14916,N_11483,N_10318);
nand U14917 (N_14917,N_9385,N_9889);
xnor U14918 (N_14918,N_10319,N_9983);
nand U14919 (N_14919,N_10439,N_11128);
nand U14920 (N_14920,N_11397,N_9147);
nand U14921 (N_14921,N_9383,N_9419);
xor U14922 (N_14922,N_10428,N_9705);
xor U14923 (N_14923,N_9827,N_11408);
nand U14924 (N_14924,N_11290,N_9512);
nand U14925 (N_14925,N_9033,N_11373);
or U14926 (N_14926,N_11261,N_11279);
or U14927 (N_14927,N_10104,N_10159);
or U14928 (N_14928,N_10328,N_10912);
xor U14929 (N_14929,N_10826,N_10899);
nand U14930 (N_14930,N_9861,N_9046);
nor U14931 (N_14931,N_10912,N_11945);
and U14932 (N_14932,N_11403,N_10937);
and U14933 (N_14933,N_9220,N_11483);
nor U14934 (N_14934,N_10039,N_10800);
and U14935 (N_14935,N_9881,N_10243);
nor U14936 (N_14936,N_10957,N_9982);
xor U14937 (N_14937,N_9460,N_10620);
and U14938 (N_14938,N_9216,N_11721);
xnor U14939 (N_14939,N_10133,N_9934);
nor U14940 (N_14940,N_11123,N_9302);
or U14941 (N_14941,N_9588,N_11512);
and U14942 (N_14942,N_11999,N_10567);
nand U14943 (N_14943,N_10519,N_11329);
xor U14944 (N_14944,N_9448,N_10155);
nand U14945 (N_14945,N_9227,N_10760);
xnor U14946 (N_14946,N_11063,N_10547);
xnor U14947 (N_14947,N_9009,N_9207);
nand U14948 (N_14948,N_9890,N_10419);
nand U14949 (N_14949,N_9695,N_10532);
xnor U14950 (N_14950,N_11604,N_9752);
nor U14951 (N_14951,N_9551,N_11495);
xor U14952 (N_14952,N_11237,N_10183);
and U14953 (N_14953,N_9471,N_10717);
xor U14954 (N_14954,N_10261,N_9874);
nand U14955 (N_14955,N_10045,N_11989);
nand U14956 (N_14956,N_11686,N_10537);
nand U14957 (N_14957,N_11713,N_10529);
nand U14958 (N_14958,N_9931,N_10183);
nand U14959 (N_14959,N_9392,N_10213);
nor U14960 (N_14960,N_9740,N_10532);
nor U14961 (N_14961,N_10812,N_11150);
and U14962 (N_14962,N_11532,N_9123);
nand U14963 (N_14963,N_9621,N_9191);
xnor U14964 (N_14964,N_11916,N_11651);
and U14965 (N_14965,N_11758,N_9627);
nor U14966 (N_14966,N_11700,N_10489);
and U14967 (N_14967,N_10541,N_10980);
and U14968 (N_14968,N_11375,N_11532);
or U14969 (N_14969,N_10852,N_9764);
nand U14970 (N_14970,N_9661,N_9431);
nand U14971 (N_14971,N_9179,N_9082);
xor U14972 (N_14972,N_11240,N_10976);
nor U14973 (N_14973,N_11139,N_10328);
or U14974 (N_14974,N_9243,N_9695);
or U14975 (N_14975,N_10972,N_9341);
nor U14976 (N_14976,N_9639,N_9778);
nand U14977 (N_14977,N_11145,N_9955);
nor U14978 (N_14978,N_9620,N_9432);
xor U14979 (N_14979,N_10849,N_9344);
nor U14980 (N_14980,N_10233,N_11455);
and U14981 (N_14981,N_10886,N_9249);
xor U14982 (N_14982,N_10255,N_11651);
or U14983 (N_14983,N_9496,N_11366);
nand U14984 (N_14984,N_9359,N_10435);
nor U14985 (N_14985,N_9389,N_9653);
nor U14986 (N_14986,N_9085,N_11242);
xor U14987 (N_14987,N_11551,N_10162);
and U14988 (N_14988,N_10541,N_11184);
or U14989 (N_14989,N_9832,N_9906);
or U14990 (N_14990,N_10932,N_10115);
nand U14991 (N_14991,N_10592,N_11526);
nor U14992 (N_14992,N_11659,N_10315);
nor U14993 (N_14993,N_9042,N_9063);
nand U14994 (N_14994,N_9734,N_10578);
and U14995 (N_14995,N_9576,N_9302);
xor U14996 (N_14996,N_9536,N_11337);
or U14997 (N_14997,N_10794,N_11134);
nand U14998 (N_14998,N_11654,N_10690);
nand U14999 (N_14999,N_11842,N_9664);
nor U15000 (N_15000,N_13465,N_14966);
xor U15001 (N_15001,N_13315,N_12026);
xnor U15002 (N_15002,N_13349,N_12000);
and U15003 (N_15003,N_13331,N_12400);
and U15004 (N_15004,N_12747,N_12037);
nor U15005 (N_15005,N_14435,N_14479);
nor U15006 (N_15006,N_13788,N_14950);
or U15007 (N_15007,N_12124,N_14862);
or U15008 (N_15008,N_12750,N_12092);
nor U15009 (N_15009,N_12500,N_12880);
xnor U15010 (N_15010,N_14442,N_14212);
or U15011 (N_15011,N_14684,N_12133);
and U15012 (N_15012,N_14523,N_12835);
or U15013 (N_15013,N_14674,N_12686);
and U15014 (N_15014,N_13474,N_14353);
xnor U15015 (N_15015,N_13037,N_14658);
xor U15016 (N_15016,N_13908,N_14404);
nand U15017 (N_15017,N_14813,N_13204);
nor U15018 (N_15018,N_12371,N_12962);
xor U15019 (N_15019,N_14800,N_14176);
nand U15020 (N_15020,N_13257,N_13581);
or U15021 (N_15021,N_13499,N_12227);
or U15022 (N_15022,N_14791,N_12040);
and U15023 (N_15023,N_13605,N_12061);
nand U15024 (N_15024,N_13805,N_13309);
or U15025 (N_15025,N_14043,N_13435);
nor U15026 (N_15026,N_12292,N_12640);
or U15027 (N_15027,N_14417,N_12138);
nand U15028 (N_15028,N_12873,N_14771);
xnor U15029 (N_15029,N_13119,N_14588);
or U15030 (N_15030,N_13999,N_14906);
or U15031 (N_15031,N_13348,N_13302);
and U15032 (N_15032,N_12552,N_12452);
and U15033 (N_15033,N_12267,N_13490);
and U15034 (N_15034,N_14820,N_14829);
xor U15035 (N_15035,N_13537,N_12679);
xor U15036 (N_15036,N_13114,N_14466);
nand U15037 (N_15037,N_13065,N_14833);
nand U15038 (N_15038,N_12905,N_13481);
xnor U15039 (N_15039,N_14840,N_14857);
nand U15040 (N_15040,N_13216,N_13663);
xor U15041 (N_15041,N_12929,N_13542);
or U15042 (N_15042,N_13325,N_12957);
or U15043 (N_15043,N_13638,N_12297);
nor U15044 (N_15044,N_13368,N_14320);
or U15045 (N_15045,N_13755,N_14072);
nor U15046 (N_15046,N_13797,N_12847);
xnor U15047 (N_15047,N_14991,N_13219);
nor U15048 (N_15048,N_14868,N_13764);
nor U15049 (N_15049,N_12579,N_12570);
nor U15050 (N_15050,N_12763,N_14084);
nand U15051 (N_15051,N_13033,N_13190);
and U15052 (N_15052,N_14690,N_12421);
nand U15053 (N_15053,N_14807,N_14068);
or U15054 (N_15054,N_14896,N_12461);
xnor U15055 (N_15055,N_12869,N_13191);
xor U15056 (N_15056,N_13978,N_14784);
or U15057 (N_15057,N_12906,N_13273);
or U15058 (N_15058,N_14639,N_12872);
nor U15059 (N_15059,N_12364,N_12740);
nor U15060 (N_15060,N_12648,N_13765);
and U15061 (N_15061,N_12870,N_12256);
and U15062 (N_15062,N_13824,N_13710);
nor U15063 (N_15063,N_12814,N_12715);
nor U15064 (N_15064,N_13704,N_12973);
or U15065 (N_15065,N_13342,N_14629);
and U15066 (N_15066,N_13462,N_14729);
and U15067 (N_15067,N_14631,N_12088);
and U15068 (N_15068,N_13120,N_12871);
xnor U15069 (N_15069,N_12219,N_14923);
nand U15070 (N_15070,N_13672,N_12649);
xnor U15071 (N_15071,N_12882,N_14201);
nor U15072 (N_15072,N_13473,N_13926);
or U15073 (N_15073,N_14134,N_12622);
and U15074 (N_15074,N_14766,N_12819);
or U15075 (N_15075,N_13711,N_14108);
and U15076 (N_15076,N_13981,N_12471);
nor U15077 (N_15077,N_14902,N_12165);
and U15078 (N_15078,N_13528,N_12466);
or U15079 (N_15079,N_12111,N_12140);
and U15080 (N_15080,N_12619,N_14093);
nand U15081 (N_15081,N_12337,N_14814);
nand U15082 (N_15082,N_12894,N_14749);
xnor U15083 (N_15083,N_14037,N_14760);
xnor U15084 (N_15084,N_13073,N_14924);
nand U15085 (N_15085,N_12407,N_13720);
and U15086 (N_15086,N_14617,N_13971);
and U15087 (N_15087,N_13066,N_14495);
and U15088 (N_15088,N_13579,N_13627);
nor U15089 (N_15089,N_13398,N_14436);
and U15090 (N_15090,N_14712,N_12776);
xnor U15091 (N_15091,N_12463,N_13659);
xor U15092 (N_15092,N_13090,N_14438);
nor U15093 (N_15093,N_12368,N_12222);
nand U15094 (N_15094,N_12303,N_14052);
xnor U15095 (N_15095,N_12498,N_13799);
nand U15096 (N_15096,N_14850,N_13818);
xor U15097 (N_15097,N_14010,N_12098);
xor U15098 (N_15098,N_13957,N_12330);
nand U15099 (N_15099,N_13222,N_13654);
xor U15100 (N_15100,N_14682,N_12845);
nor U15101 (N_15101,N_12947,N_13186);
nand U15102 (N_15102,N_13743,N_12029);
nor U15103 (N_15103,N_13646,N_13378);
nand U15104 (N_15104,N_12356,N_14194);
nor U15105 (N_15105,N_13941,N_12258);
and U15106 (N_15106,N_12423,N_12441);
or U15107 (N_15107,N_13841,N_13949);
nand U15108 (N_15108,N_14211,N_12735);
or U15109 (N_15109,N_12109,N_12879);
nor U15110 (N_15110,N_13652,N_12172);
or U15111 (N_15111,N_12090,N_13123);
or U15112 (N_15112,N_13624,N_13265);
nor U15113 (N_15113,N_12002,N_14964);
nor U15114 (N_15114,N_12593,N_13723);
nand U15115 (N_15115,N_12709,N_12033);
nor U15116 (N_15116,N_14382,N_14024);
nor U15117 (N_15117,N_13236,N_12313);
nor U15118 (N_15118,N_13148,N_12772);
xor U15119 (N_15119,N_14488,N_14511);
nor U15120 (N_15120,N_13272,N_12044);
nor U15121 (N_15121,N_14501,N_12557);
nand U15122 (N_15122,N_12866,N_12827);
and U15123 (N_15123,N_14255,N_13596);
nor U15124 (N_15124,N_13238,N_14313);
nand U15125 (N_15125,N_12157,N_14516);
xor U15126 (N_15126,N_13958,N_12083);
nor U15127 (N_15127,N_12363,N_13449);
nor U15128 (N_15128,N_12399,N_14431);
nand U15129 (N_15129,N_13112,N_13443);
or U15130 (N_15130,N_12568,N_13850);
nor U15131 (N_15131,N_12308,N_14195);
nand U15132 (N_15132,N_13021,N_12526);
xor U15133 (N_15133,N_12417,N_14196);
xnor U15134 (N_15134,N_14224,N_14292);
nand U15135 (N_15135,N_13403,N_14260);
nor U15136 (N_15136,N_14803,N_13223);
xnor U15137 (N_15137,N_12006,N_13567);
xor U15138 (N_15138,N_12253,N_12147);
nand U15139 (N_15139,N_13504,N_14133);
nand U15140 (N_15140,N_12966,N_12774);
xnor U15141 (N_15141,N_13385,N_13514);
and U15142 (N_15142,N_14032,N_14337);
nand U15143 (N_15143,N_14143,N_13811);
nor U15144 (N_15144,N_14054,N_13893);
or U15145 (N_15145,N_13386,N_12606);
nand U15146 (N_15146,N_12202,N_14519);
nor U15147 (N_15147,N_14701,N_14200);
nand U15148 (N_15148,N_12344,N_13096);
and U15149 (N_15149,N_14244,N_13545);
or U15150 (N_15150,N_14508,N_14344);
and U15151 (N_15151,N_14559,N_12112);
nor U15152 (N_15152,N_12554,N_13880);
xor U15153 (N_15153,N_13457,N_14379);
nor U15154 (N_15154,N_13943,N_14048);
or U15155 (N_15155,N_12838,N_12720);
or U15156 (N_15156,N_12346,N_14047);
or U15157 (N_15157,N_13661,N_12608);
and U15158 (N_15158,N_14920,N_14467);
nor U15159 (N_15159,N_14533,N_12472);
or U15160 (N_15160,N_14461,N_13715);
xnor U15161 (N_15161,N_13305,N_14447);
nor U15162 (N_15162,N_13275,N_14492);
or U15163 (N_15163,N_12639,N_13778);
and U15164 (N_15164,N_13869,N_13217);
nor U15165 (N_15165,N_12700,N_13707);
and U15166 (N_15166,N_14755,N_14737);
nand U15167 (N_15167,N_13936,N_14969);
xnor U15168 (N_15168,N_14262,N_14103);
or U15169 (N_15169,N_12723,N_14149);
and U15170 (N_15170,N_12315,N_14022);
nor U15171 (N_15171,N_14377,N_13396);
and U15172 (N_15172,N_12183,N_13050);
and U15173 (N_15173,N_13290,N_13166);
nand U15174 (N_15174,N_13431,N_13780);
nor U15175 (N_15175,N_13650,N_12110);
xnor U15176 (N_15176,N_12285,N_13301);
nand U15177 (N_15177,N_13790,N_12385);
or U15178 (N_15178,N_12612,N_14997);
or U15179 (N_15179,N_14939,N_14387);
nor U15180 (N_15180,N_13669,N_12078);
xor U15181 (N_15181,N_13994,N_14935);
and U15182 (N_15182,N_12493,N_13702);
or U15183 (N_15183,N_12232,N_13570);
or U15184 (N_15184,N_12668,N_13133);
nor U15185 (N_15185,N_12372,N_13234);
or U15186 (N_15186,N_12597,N_14153);
nand U15187 (N_15187,N_12724,N_13218);
nand U15188 (N_15188,N_14240,N_13067);
and U15189 (N_15189,N_14276,N_14191);
and U15190 (N_15190,N_13501,N_13135);
and U15191 (N_15191,N_13782,N_12024);
nor U15192 (N_15192,N_12178,N_13251);
or U15193 (N_15193,N_12596,N_12139);
nor U15194 (N_15194,N_14113,N_13529);
and U15195 (N_15195,N_12143,N_13823);
and U15196 (N_15196,N_14651,N_13170);
or U15197 (N_15197,N_12938,N_13752);
and U15198 (N_15198,N_13513,N_14897);
nand U15199 (N_15199,N_14376,N_14159);
nor U15200 (N_15200,N_13634,N_13747);
or U15201 (N_15201,N_14815,N_14750);
or U15202 (N_15202,N_13837,N_13987);
or U15203 (N_15203,N_13288,N_12121);
or U15204 (N_15204,N_13608,N_12120);
and U15205 (N_15205,N_13918,N_12376);
nor U15206 (N_15206,N_12004,N_12361);
and U15207 (N_15207,N_12924,N_12064);
xor U15208 (N_15208,N_14926,N_14463);
nor U15209 (N_15209,N_14056,N_13919);
or U15210 (N_15210,N_12142,N_12296);
nand U15211 (N_15211,N_12739,N_13871);
nor U15212 (N_15212,N_12341,N_12997);
xor U15213 (N_15213,N_12177,N_14356);
nand U15214 (N_15214,N_14128,N_13613);
and U15215 (N_15215,N_13963,N_12413);
nor U15216 (N_15216,N_13068,N_13184);
xnor U15217 (N_15217,N_12795,N_12940);
nand U15218 (N_15218,N_14555,N_14077);
nor U15219 (N_15219,N_14940,N_14537);
nand U15220 (N_15220,N_13952,N_14531);
and U15221 (N_15221,N_13072,N_14172);
nand U15222 (N_15222,N_13269,N_13716);
and U15223 (N_15223,N_14206,N_14328);
nand U15224 (N_15224,N_13134,N_13617);
nand U15225 (N_15225,N_13489,N_12751);
and U15226 (N_15226,N_13069,N_14947);
and U15227 (N_15227,N_14319,N_14247);
nand U15228 (N_15228,N_13372,N_14780);
nand U15229 (N_15229,N_14876,N_12843);
nand U15230 (N_15230,N_13682,N_14756);
nor U15231 (N_15231,N_13569,N_13556);
nor U15232 (N_15232,N_13879,N_12789);
nand U15233 (N_15233,N_12848,N_12107);
xor U15234 (N_15234,N_14859,N_14861);
or U15235 (N_15235,N_12416,N_14647);
xor U15236 (N_15236,N_13897,N_14823);
and U15237 (N_15237,N_12479,N_13580);
and U15238 (N_15238,N_14065,N_14021);
nor U15239 (N_15239,N_14066,N_14480);
or U15240 (N_15240,N_14595,N_13891);
or U15241 (N_15241,N_14165,N_12213);
or U15242 (N_15242,N_12660,N_12068);
and U15243 (N_15243,N_14996,N_13945);
nand U15244 (N_15244,N_12710,N_13175);
and U15245 (N_15245,N_13576,N_13227);
nor U15246 (N_15246,N_14816,N_13420);
xor U15247 (N_15247,N_13336,N_12742);
and U15248 (N_15248,N_14992,N_12212);
nand U15249 (N_15249,N_13200,N_13611);
nand U15250 (N_15250,N_12013,N_14100);
nor U15251 (N_15251,N_14144,N_14767);
nand U15252 (N_15252,N_14029,N_12974);
nor U15253 (N_15253,N_13598,N_13022);
or U15254 (N_15254,N_12066,N_13754);
nand U15255 (N_15255,N_13180,N_12022);
nor U15256 (N_15256,N_13258,N_13464);
nand U15257 (N_15257,N_12295,N_13008);
xnor U15258 (N_15258,N_14246,N_12489);
and U15259 (N_15259,N_13430,N_13688);
xor U15260 (N_15260,N_12225,N_13507);
nand U15261 (N_15261,N_14624,N_14359);
nand U15262 (N_15262,N_12440,N_13736);
nor U15263 (N_15263,N_12338,N_14653);
or U15264 (N_15264,N_14424,N_14297);
nor U15265 (N_15265,N_13318,N_14887);
nor U15266 (N_15266,N_14142,N_12290);
nor U15267 (N_15267,N_14703,N_14728);
or U15268 (N_15268,N_13140,N_12696);
and U15269 (N_15269,N_12888,N_14156);
xor U15270 (N_15270,N_14104,N_14409);
or U15271 (N_15271,N_14931,N_12490);
nand U15272 (N_15272,N_12837,N_13359);
nand U15273 (N_15273,N_13966,N_14787);
or U15274 (N_15274,N_13027,N_14584);
xnor U15275 (N_15275,N_12398,N_12070);
or U15276 (N_15276,N_13758,N_13341);
nand U15277 (N_15277,N_14087,N_14311);
nand U15278 (N_15278,N_13517,N_13121);
and U15279 (N_15279,N_13032,N_13375);
nand U15280 (N_15280,N_12584,N_13480);
xor U15281 (N_15281,N_14918,N_12706);
or U15282 (N_15282,N_12983,N_13195);
xnor U15283 (N_15283,N_13012,N_14395);
nand U15284 (N_15284,N_12049,N_12126);
nor U15285 (N_15285,N_12573,N_12443);
nor U15286 (N_15286,N_14761,N_13374);
or U15287 (N_15287,N_14589,N_14943);
xor U15288 (N_15288,N_13577,N_14822);
nor U15289 (N_15289,N_13831,N_14788);
or U15290 (N_15290,N_14838,N_12023);
nor U15291 (N_15291,N_14839,N_14139);
and U15292 (N_15292,N_13434,N_12555);
or U15293 (N_15293,N_13300,N_12692);
nand U15294 (N_15294,N_12652,N_13593);
nor U15295 (N_15295,N_12893,N_14632);
and U15296 (N_15296,N_12482,N_14659);
nor U15297 (N_15297,N_13395,N_12276);
nand U15298 (N_15298,N_13802,N_14683);
and U15299 (N_15299,N_14942,N_12424);
and U15300 (N_15300,N_12305,N_13011);
xor U15301 (N_15301,N_14117,N_12512);
nand U15302 (N_15302,N_14827,N_14455);
or U15303 (N_15303,N_12569,N_12743);
xnor U15304 (N_15304,N_13165,N_14673);
and U15305 (N_15305,N_14535,N_14173);
or U15306 (N_15306,N_14768,N_14323);
nor U15307 (N_15307,N_14972,N_12603);
nor U15308 (N_15308,N_13295,N_12239);
and U15309 (N_15309,N_12190,N_12056);
and U15310 (N_15310,N_13651,N_13345);
and U15311 (N_15311,N_13083,N_14114);
or U15312 (N_15312,N_14953,N_14871);
nor U15313 (N_15313,N_14470,N_14818);
or U15314 (N_15314,N_14486,N_13533);
and U15315 (N_15315,N_12846,N_12200);
nand U15316 (N_15316,N_12884,N_14672);
or U15317 (N_15317,N_12647,N_14708);
nor U15318 (N_15318,N_13137,N_12809);
and U15319 (N_15319,N_12684,N_12547);
nand U15320 (N_15320,N_12455,N_13129);
nand U15321 (N_15321,N_13583,N_14059);
nand U15322 (N_15322,N_12299,N_13245);
or U15323 (N_15323,N_14085,N_14169);
xor U15324 (N_15324,N_12486,N_13587);
nor U15325 (N_15325,N_14355,N_12430);
nand U15326 (N_15326,N_12558,N_12127);
xnor U15327 (N_15327,N_12345,N_13687);
nor U15328 (N_15328,N_12535,N_12448);
or U15329 (N_15329,N_13093,N_12229);
nand U15330 (N_15330,N_13351,N_12651);
xnor U15331 (N_15331,N_12524,N_14221);
and U15332 (N_15332,N_14762,N_14154);
nor U15333 (N_15333,N_14882,N_13019);
nor U15334 (N_15334,N_14158,N_14977);
nor U15335 (N_15335,N_12021,N_14464);
nor U15336 (N_15336,N_12528,N_13920);
xnor U15337 (N_15337,N_14229,N_13559);
or U15338 (N_15338,N_14805,N_12807);
nand U15339 (N_15339,N_12980,N_12970);
or U15340 (N_15340,N_13494,N_13762);
or U15341 (N_15341,N_14704,N_13785);
or U15342 (N_15342,N_14569,N_12084);
nor U15343 (N_15343,N_14975,N_12699);
nor U15344 (N_15344,N_14284,N_13154);
xnor U15345 (N_15345,N_12708,N_13772);
and U15346 (N_15346,N_13080,N_13940);
and U15347 (N_15347,N_14676,N_13684);
nor U15348 (N_15348,N_12758,N_14643);
xor U15349 (N_15349,N_14853,N_14619);
xor U15350 (N_15350,N_13621,N_13260);
and U15351 (N_15351,N_12867,N_13010);
and U15352 (N_15352,N_14951,N_14952);
nand U15353 (N_15353,N_14558,N_13967);
or U15354 (N_15354,N_12682,N_12946);
and U15355 (N_15355,N_13822,N_13064);
nor U15356 (N_15356,N_12504,N_12265);
or U15357 (N_15357,N_14548,N_14257);
or U15358 (N_15358,N_13052,N_13402);
xnor U15359 (N_15359,N_13894,N_13673);
or U15360 (N_15360,N_12101,N_13319);
and U15361 (N_15361,N_12250,N_14922);
xnor U15362 (N_15362,N_12826,N_12839);
and U15363 (N_15363,N_13700,N_12615);
nand U15364 (N_15364,N_14001,N_13146);
xor U15365 (N_15365,N_14270,N_13000);
nor U15366 (N_15366,N_13708,N_14763);
nand U15367 (N_15367,N_13872,N_14097);
nor U15368 (N_15368,N_12760,N_12063);
or U15369 (N_15369,N_13411,N_14462);
xor U15370 (N_15370,N_14306,N_14864);
and U15371 (N_15371,N_13699,N_13429);
nand U15372 (N_15372,N_13025,N_12234);
or U15373 (N_15373,N_13535,N_13326);
nor U15374 (N_15374,N_12678,N_14581);
nand U15375 (N_15375,N_12041,N_12191);
xnor U15376 (N_15376,N_13070,N_13224);
or U15377 (N_15377,N_13992,N_14654);
nand U15378 (N_15378,N_13857,N_13902);
nand U15379 (N_15379,N_12716,N_13968);
nor U15380 (N_15380,N_12333,N_12354);
or U15381 (N_15381,N_13697,N_12560);
nand U15382 (N_15382,N_14677,N_12707);
nand U15383 (N_15383,N_12633,N_12726);
nand U15384 (N_15384,N_14667,N_14491);
nor U15385 (N_15385,N_12446,N_13844);
nor U15386 (N_15386,N_12670,N_14811);
nor U15387 (N_15387,N_13082,N_14266);
nand U15388 (N_15388,N_14640,N_14405);
and U15389 (N_15389,N_13107,N_13448);
or U15390 (N_15390,N_13206,N_12192);
nor U15391 (N_15391,N_12806,N_13158);
nor U15392 (N_15392,N_12144,N_12808);
or U15393 (N_15393,N_12397,N_13192);
and U15394 (N_15394,N_13212,N_12357);
nor U15395 (N_15395,N_14529,N_14331);
xor U15396 (N_15396,N_12018,N_13575);
and U15397 (N_15397,N_12168,N_13827);
or U15398 (N_15398,N_12347,N_12264);
xor U15399 (N_15399,N_14759,N_13680);
and U15400 (N_15400,N_13405,N_12895);
or U15401 (N_15401,N_14810,N_13671);
nand U15402 (N_15402,N_14723,N_13532);
nor U15403 (N_15403,N_14626,N_14053);
and U15404 (N_15404,N_14202,N_13739);
or U15405 (N_15405,N_13503,N_14913);
xor U15406 (N_15406,N_13267,N_13103);
and U15407 (N_15407,N_13769,N_14120);
and U15408 (N_15408,N_13214,N_12517);
and U15409 (N_15409,N_14241,N_13479);
xor U15410 (N_15410,N_14388,N_12851);
and U15411 (N_15411,N_13925,N_13383);
or U15412 (N_15412,N_12152,N_12289);
nand U15413 (N_15413,N_14801,N_14493);
nand U15414 (N_15414,N_14646,N_12465);
xor U15415 (N_15415,N_14129,N_14506);
nand U15416 (N_15416,N_12223,N_12175);
nor U15417 (N_15417,N_14809,N_12811);
nand U15418 (N_15418,N_14457,N_14573);
and U15419 (N_15419,N_13692,N_14845);
or U15420 (N_15420,N_14606,N_12734);
xnor U15421 (N_15421,N_12487,N_14718);
nor U15422 (N_15422,N_12729,N_13807);
nand U15423 (N_15423,N_12282,N_14986);
or U15424 (N_15424,N_12307,N_12171);
nand U15425 (N_15425,N_12450,N_12391);
nand U15426 (N_15426,N_12829,N_12920);
or U15427 (N_15427,N_14426,N_14099);
nor U15428 (N_15428,N_13510,N_13746);
and U15429 (N_15429,N_12717,N_13796);
and U15430 (N_15430,N_12667,N_14530);
nand U15431 (N_15431,N_12702,N_14795);
xnor U15432 (N_15432,N_14773,N_13491);
xor U15433 (N_15433,N_13938,N_13923);
nand U15434 (N_15434,N_12325,N_12431);
xnor U15435 (N_15435,N_13757,N_12833);
nor U15436 (N_15436,N_13156,N_14502);
and U15437 (N_15437,N_14781,N_14638);
xor U15438 (N_15438,N_14711,N_12977);
xnor U15439 (N_15439,N_12328,N_14118);
nor U15440 (N_15440,N_13777,N_14338);
and U15441 (N_15441,N_13609,N_13492);
or U15442 (N_15442,N_12242,N_12787);
nand U15443 (N_15443,N_13328,N_12062);
nand U15444 (N_15444,N_12320,N_12409);
nor U15445 (N_15445,N_12134,N_13105);
and U15446 (N_15446,N_14391,N_12852);
or U15447 (N_15447,N_14049,N_13896);
and U15448 (N_15448,N_12351,N_13571);
nand U15449 (N_15449,N_12211,N_12657);
xnor U15450 (N_15450,N_12671,N_14296);
or U15451 (N_15451,N_14254,N_12360);
xnor U15452 (N_15452,N_12336,N_14786);
or U15453 (N_15453,N_12105,N_14278);
nand U15454 (N_15454,N_12079,N_13995);
xor U15455 (N_15455,N_12331,N_14515);
or U15456 (N_15456,N_12759,N_13338);
and U15457 (N_15457,N_12616,N_12269);
or U15458 (N_15458,N_12859,N_14277);
xnor U15459 (N_15459,N_13839,N_12950);
xor U15460 (N_15460,N_14340,N_13885);
or U15461 (N_15461,N_14259,N_13693);
or U15462 (N_15462,N_13237,N_14577);
xor U15463 (N_15463,N_14448,N_13679);
nor U15464 (N_15464,N_12773,N_13884);
and U15465 (N_15465,N_13459,N_14329);
xnor U15466 (N_15466,N_13155,N_12036);
and U15467 (N_15467,N_14967,N_13582);
or U15468 (N_15468,N_14305,N_14288);
xor U15469 (N_15469,N_12028,N_14532);
nand U15470 (N_15470,N_13486,N_14834);
nor U15471 (N_15471,N_12402,N_12031);
nand U15472 (N_15472,N_12404,N_12992);
and U15473 (N_15473,N_14738,N_14851);
or U15474 (N_15474,N_12677,N_13870);
nand U15475 (N_15475,N_14450,N_14751);
xnor U15476 (N_15476,N_14858,N_13097);
or U15477 (N_15477,N_13589,N_13565);
nand U15478 (N_15478,N_13944,N_12664);
nand U15479 (N_15479,N_12949,N_13914);
or U15480 (N_15480,N_13293,N_12745);
or U15481 (N_15481,N_13882,N_13607);
nand U15482 (N_15482,N_12598,N_14790);
nor U15483 (N_15483,N_12681,N_13889);
and U15484 (N_15484,N_13418,N_14747);
or U15485 (N_15485,N_13117,N_12892);
nand U15486 (N_15486,N_13197,N_12802);
nand U15487 (N_15487,N_13544,N_13899);
nor U15488 (N_15488,N_14067,N_12624);
nor U15489 (N_15489,N_13637,N_12459);
xor U15490 (N_15490,N_13628,N_14303);
or U15491 (N_15491,N_14189,N_12050);
or U15492 (N_15492,N_13436,N_13380);
nand U15493 (N_15493,N_13770,N_13546);
nand U15494 (N_15494,N_12816,N_14497);
nand U15495 (N_15495,N_13643,N_12069);
and U15496 (N_15496,N_12245,N_14383);
or U15497 (N_15497,N_14399,N_12812);
nand U15498 (N_15498,N_13040,N_14524);
or U15499 (N_15499,N_14783,N_13803);
or U15500 (N_15500,N_12327,N_12505);
or U15501 (N_15501,N_13719,N_13915);
or U15502 (N_15502,N_14177,N_13183);
nor U15503 (N_15503,N_14141,N_14429);
and U15504 (N_15504,N_13228,N_14289);
or U15505 (N_15505,N_14451,N_13210);
nor U15506 (N_15506,N_13043,N_14956);
and U15507 (N_15507,N_12959,N_13002);
or U15508 (N_15508,N_13401,N_13006);
nand U15509 (N_15509,N_14549,N_14927);
nand U15510 (N_15510,N_12387,N_14469);
and U15511 (N_15511,N_13079,N_13965);
xnor U15512 (N_15512,N_13705,N_14880);
nor U15513 (N_15513,N_14199,N_14027);
and U15514 (N_15514,N_14908,N_14112);
and U15515 (N_15515,N_13960,N_14441);
nand U15516 (N_15516,N_14959,N_13522);
or U15517 (N_15517,N_13306,N_12883);
nand U15518 (N_15518,N_13560,N_12689);
or U15519 (N_15519,N_12060,N_12737);
or U15520 (N_15520,N_14550,N_12551);
xnor U15521 (N_15521,N_13690,N_12255);
nand U15522 (N_15522,N_13815,N_12104);
or U15523 (N_15523,N_12468,N_12928);
or U15524 (N_15524,N_13525,N_14089);
xnor U15525 (N_15525,N_12359,N_14557);
xor U15526 (N_15526,N_14343,N_12697);
nor U15527 (N_15527,N_13698,N_12458);
or U15528 (N_15528,N_14420,N_13487);
nand U15529 (N_15529,N_13060,N_12790);
nand U15530 (N_15530,N_12011,N_12844);
nand U15531 (N_15531,N_14026,N_12767);
nor U15532 (N_15532,N_12599,N_14637);
xnor U15533 (N_15533,N_12984,N_14752);
nand U15534 (N_15534,N_14476,N_13005);
nand U15535 (N_15535,N_13922,N_14609);
nor U15536 (N_15536,N_14733,N_13722);
nand U15537 (N_15537,N_12577,N_13390);
nand U15538 (N_15538,N_13427,N_13883);
and U15539 (N_15539,N_14375,N_13685);
nor U15540 (N_15540,N_14452,N_14765);
nand U15541 (N_15541,N_14105,N_14490);
and U15542 (N_15542,N_12861,N_13864);
nor U15543 (N_15543,N_12817,N_14109);
or U15544 (N_15544,N_13982,N_13614);
nor U15545 (N_15545,N_14916,N_13404);
nand U15546 (N_15546,N_14693,N_14999);
xnor U15547 (N_15547,N_14870,N_13364);
and U15548 (N_15548,N_13703,N_13534);
nand U15549 (N_15549,N_13139,N_13733);
or U15550 (N_15550,N_14846,N_14171);
xor U15551 (N_15551,N_14365,N_12301);
and U15552 (N_15552,N_12159,N_13619);
or U15553 (N_15553,N_13388,N_14957);
nor U15554 (N_15554,N_12964,N_13773);
xor U15555 (N_15555,N_13907,N_12293);
and U15556 (N_15556,N_12923,N_12730);
or U15557 (N_15557,N_13713,N_13730);
xnor U15558 (N_15558,N_13604,N_12335);
nand U15559 (N_15559,N_14691,N_12864);
or U15560 (N_15560,N_12663,N_14362);
or U15561 (N_15561,N_14033,N_12785);
nor U15562 (N_15562,N_13298,N_12771);
nor U15563 (N_15563,N_14419,N_13104);
nand U15564 (N_15564,N_13160,N_14251);
xor U15565 (N_15565,N_14970,N_13985);
and U15566 (N_15566,N_12214,N_12945);
and U15567 (N_15567,N_12875,N_12972);
nor U15568 (N_15568,N_13094,N_14782);
and U15569 (N_15569,N_14526,N_14094);
xor U15570 (N_15570,N_13816,N_14610);
or U15571 (N_15571,N_14422,N_12621);
nor U15572 (N_15572,N_13821,N_13303);
nand U15573 (N_15573,N_13658,N_14095);
nand U15574 (N_15574,N_14290,N_12353);
nor U15575 (N_15575,N_14613,N_13728);
nor U15576 (N_15576,N_12511,N_14603);
xor U15577 (N_15577,N_14096,N_14697);
xnor U15578 (N_15578,N_13519,N_12187);
and U15579 (N_15579,N_14849,N_12752);
xor U15580 (N_15580,N_12382,N_14612);
or U15581 (N_15581,N_13555,N_14321);
nand U15582 (N_15582,N_14116,N_13458);
xnor U15583 (N_15583,N_14778,N_12799);
or U15584 (N_15584,N_14279,N_12095);
or U15585 (N_15585,N_14025,N_14265);
xnor U15586 (N_15586,N_12329,N_12129);
or U15587 (N_15587,N_12655,N_12447);
and U15588 (N_15588,N_12097,N_13676);
nand U15589 (N_15589,N_14650,N_14011);
nand U15590 (N_15590,N_12993,N_12913);
nand U15591 (N_15591,N_13826,N_13353);
or U15592 (N_15592,N_12174,N_14869);
or U15593 (N_15593,N_13741,N_14070);
xnor U15594 (N_15594,N_14473,N_13861);
xor U15595 (N_15595,N_12266,N_14601);
nor U15596 (N_15596,N_13497,N_12015);
nand U15597 (N_15597,N_14228,N_12437);
nor U15598 (N_15598,N_13447,N_13947);
or U15599 (N_15599,N_13159,N_13877);
xnor U15600 (N_15600,N_12220,N_13738);
nand U15601 (N_15601,N_14806,N_12525);
xnor U15602 (N_15602,N_12496,N_14465);
xnor U15603 (N_15603,N_12273,N_12196);
and U15604 (N_15604,N_14520,N_12150);
or U15605 (N_15605,N_13724,N_14794);
nand U15606 (N_15606,N_13182,N_12470);
nand U15607 (N_15607,N_14204,N_14400);
nor U15608 (N_15608,N_14724,N_12830);
xnor U15609 (N_15609,N_13508,N_12204);
nor U15610 (N_15610,N_13167,N_14147);
nand U15611 (N_15611,N_13421,N_12247);
nand U15612 (N_15612,N_14243,N_14798);
or U15613 (N_15613,N_12203,N_14168);
or U15614 (N_15614,N_12567,N_12953);
xnor U15615 (N_15615,N_13794,N_12287);
and U15616 (N_15616,N_13574,N_13437);
nand U15617 (N_15617,N_14742,N_13440);
nor U15618 (N_15618,N_12367,N_14645);
nand U15619 (N_15619,N_13207,N_14962);
nor U15620 (N_15620,N_13742,N_13886);
or U15621 (N_15621,N_13863,N_12932);
nand U15622 (N_15622,N_13511,N_12236);
nor U15623 (N_15623,N_12925,N_14406);
nor U15624 (N_15624,N_12971,N_12676);
and U15625 (N_15625,N_13578,N_13048);
xnor U15626 (N_15626,N_14592,N_13161);
nor U15627 (N_15627,N_12286,N_14272);
nand U15628 (N_15628,N_12757,N_14616);
or U15629 (N_15629,N_14151,N_14883);
xor U15630 (N_15630,N_13644,N_12252);
xnor U15631 (N_15631,N_12549,N_13394);
or U15632 (N_15632,N_12768,N_13745);
xnor U15633 (N_15633,N_14456,N_13426);
and U15634 (N_15634,N_12012,N_14552);
nor U15635 (N_15635,N_12057,N_14514);
nand U15636 (N_15636,N_14536,N_14625);
xor U15637 (N_15637,N_13558,N_12659);
or U15638 (N_15638,N_12491,N_12017);
xnor U15639 (N_15639,N_12444,N_13928);
nand U15640 (N_15640,N_14299,N_13789);
and U15641 (N_15641,N_13162,N_12502);
xor U15642 (N_15642,N_12927,N_12374);
nand U15643 (N_15643,N_13313,N_13128);
or U15644 (N_15644,N_12155,N_12712);
and U15645 (N_15645,N_12395,N_12027);
and U15646 (N_15646,N_14847,N_13756);
or U15647 (N_15647,N_13087,N_12581);
nor U15648 (N_15648,N_13732,N_14102);
or U15649 (N_15649,N_12281,N_14135);
nand U15650 (N_15650,N_14895,N_13176);
nor U15651 (N_15651,N_13470,N_12607);
xor U15652 (N_15652,N_13475,N_13538);
and U15653 (N_15653,N_14046,N_14258);
xnor U15654 (N_15654,N_12449,N_12460);
or U15655 (N_15655,N_13523,N_12432);
nand U15656 (N_15656,N_14933,N_13376);
or U15657 (N_15657,N_13285,N_13042);
or U15658 (N_15658,N_14336,N_14444);
or U15659 (N_15659,N_14357,N_14454);
or U15660 (N_15660,N_14418,N_14339);
or U15661 (N_15661,N_14837,N_14035);
nand U15662 (N_15662,N_14275,N_12497);
or U15663 (N_15663,N_14496,N_14013);
and U15664 (N_15664,N_12563,N_14891);
nor U15665 (N_15665,N_13976,N_13681);
xnor U15666 (N_15666,N_13075,N_13817);
and U15667 (N_15667,N_12904,N_13996);
xnor U15668 (N_15668,N_14627,N_14274);
or U15669 (N_15669,N_13955,N_12778);
xor U15670 (N_15670,N_12506,N_14681);
nor U15671 (N_15671,N_12467,N_12545);
xor U15672 (N_15672,N_12588,N_14666);
nor U15673 (N_15673,N_12154,N_12189);
xor U15674 (N_15674,N_13231,N_14757);
nor U15675 (N_15675,N_12262,N_13187);
xor U15676 (N_15676,N_12480,N_14754);
nand U15677 (N_15677,N_13324,N_12304);
and U15678 (N_15678,N_14350,N_13686);
xnor U15679 (N_15679,N_13526,N_12071);
nor U15680 (N_15680,N_13800,N_14985);
nand U15681 (N_15681,N_14715,N_14079);
and U15682 (N_15682,N_14655,N_14263);
and U15683 (N_15683,N_12373,N_13412);
nor U15684 (N_15684,N_12484,N_14984);
nor U15685 (N_15685,N_14332,N_12166);
nand U15686 (N_15686,N_12003,N_12494);
nand U15687 (N_15687,N_12197,N_12248);
nand U15688 (N_15688,N_14425,N_12319);
xor U15689 (N_15689,N_14408,N_14374);
and U15690 (N_15690,N_12221,N_14250);
nor U15691 (N_15691,N_12316,N_12961);
xor U15692 (N_15692,N_14322,N_13361);
nor U15693 (N_15693,N_13890,N_12379);
nand U15694 (N_15694,N_14505,N_12912);
nor U15695 (N_15695,N_12691,N_14354);
and U15696 (N_15696,N_12451,N_14190);
xnor U15697 (N_15697,N_14416,N_14449);
nand U15698 (N_15698,N_14744,N_13744);
nand U15699 (N_15699,N_12001,N_14346);
and U15700 (N_15700,N_13865,N_12508);
nor U15701 (N_15701,N_13906,N_12130);
and U15702 (N_15702,N_14286,N_13601);
or U15703 (N_15703,N_12080,N_12326);
or U15704 (N_15704,N_12592,N_12137);
xnor U15705 (N_15705,N_12765,N_14217);
nor U15706 (N_15706,N_12094,N_12690);
or U15707 (N_15707,N_12085,N_14434);
nand U15708 (N_15708,N_14227,N_12823);
xnor U15709 (N_15709,N_14091,N_14423);
and U15710 (N_15710,N_14092,N_13633);
and U15711 (N_15711,N_13640,N_12156);
and U15712 (N_15712,N_12548,N_12401);
nor U15713 (N_15713,N_12237,N_14914);
and U15714 (N_15714,N_14062,N_13354);
xor U15715 (N_15715,N_12251,N_14468);
or U15716 (N_15716,N_14083,N_14656);
or U15717 (N_15717,N_14620,N_13235);
nor U15718 (N_15718,N_13951,N_12048);
nand U15719 (N_15719,N_12828,N_13721);
or U15720 (N_15720,N_12342,N_13356);
nor U15721 (N_15721,N_12499,N_13062);
and U15722 (N_15722,N_14309,N_14894);
or U15723 (N_15723,N_13691,N_13456);
nor U15724 (N_15724,N_12117,N_12714);
xor U15725 (N_15725,N_13111,N_12673);
nor U15726 (N_15726,N_14877,N_13471);
and U15727 (N_15727,N_12510,N_14386);
nand U15728 (N_15728,N_13820,N_14993);
nor U15729 (N_15729,N_14061,N_13292);
and U15730 (N_15730,N_12995,N_12944);
nor U15731 (N_15731,N_12666,N_14660);
xor U15732 (N_15732,N_13502,N_12918);
nand U15733 (N_15733,N_12406,N_14622);
xor U15734 (N_15734,N_12410,N_12182);
nor U15735 (N_15735,N_13626,N_13874);
nand U15736 (N_15736,N_14960,N_13106);
nand U15737 (N_15737,N_14596,N_14184);
nand U15738 (N_15738,N_12428,N_14662);
nand U15739 (N_15739,N_14649,N_14598);
nor U15740 (N_15740,N_12038,N_12917);
nor U15741 (N_15741,N_13866,N_14563);
or U15742 (N_15742,N_14004,N_13076);
and U15743 (N_15743,N_14576,N_12915);
and U15744 (N_15744,N_14358,N_14007);
and U15745 (N_15745,N_14776,N_14963);
xnor U15746 (N_15746,N_12891,N_13895);
nor U15747 (N_15747,N_13130,N_12609);
and U15748 (N_15748,N_13108,N_13875);
xor U15749 (N_15749,N_12414,N_14157);
and U15750 (N_15750,N_14973,N_14714);
or U15751 (N_15751,N_14855,N_14844);
xnor U15752 (N_15752,N_13280,N_14236);
nand U15753 (N_15753,N_12352,N_14875);
nand U15754 (N_15754,N_14432,N_13563);
and U15755 (N_15755,N_14580,N_13786);
xor U15756 (N_15756,N_12877,N_13808);
nor U15757 (N_15757,N_12518,N_12705);
and U15758 (N_15758,N_12065,N_12375);
xor U15759 (N_15759,N_13612,N_13858);
nand U15760 (N_15760,N_13683,N_14064);
and U15761 (N_15761,N_13392,N_12199);
and U15762 (N_15762,N_12749,N_12638);
nand U15763 (N_15763,N_12791,N_13198);
or U15764 (N_15764,N_12243,N_14140);
or U15765 (N_15765,N_13828,N_12514);
or U15766 (N_15766,N_14594,N_14216);
nor U15767 (N_15767,N_13615,N_14398);
or U15768 (N_15768,N_13979,N_14904);
xor U15769 (N_15769,N_13442,N_13282);
nor U15770 (N_15770,N_12941,N_14335);
nor U15771 (N_15771,N_13098,N_13389);
or U15772 (N_15772,N_13586,N_13330);
nand U15773 (N_15773,N_13842,N_12100);
xor U15774 (N_15774,N_12711,N_12858);
nand U15775 (N_15775,N_14621,N_13438);
xnor U15776 (N_15776,N_12149,N_12756);
nor U15777 (N_15777,N_13515,N_13393);
or U15778 (N_15778,N_14209,N_12170);
nand U15779 (N_15779,N_14641,N_14611);
or U15780 (N_15780,N_13028,N_12796);
or U15781 (N_15781,N_12793,N_13053);
nor U15782 (N_15782,N_14411,N_14812);
or U15783 (N_15783,N_13618,N_13370);
xnor U15784 (N_15784,N_13379,N_13026);
and U15785 (N_15785,N_13734,N_13964);
xnor U15786 (N_15786,N_14802,N_14590);
xnor U15787 (N_15787,N_12762,N_12614);
xnor U15788 (N_15788,N_12310,N_14239);
nor U15789 (N_15789,N_14345,N_12865);
nand U15790 (N_15790,N_14186,N_12803);
nor U15791 (N_15791,N_14553,N_12741);
nand U15792 (N_15792,N_12481,N_13856);
and U15793 (N_15793,N_14050,N_14045);
nand U15794 (N_15794,N_13332,N_14223);
or U15795 (N_15795,N_14831,N_13548);
nand U15796 (N_15796,N_14132,N_14758);
or U15797 (N_15797,N_12118,N_13813);
or U15798 (N_15798,N_12334,N_13568);
nand U15799 (N_15799,N_12908,N_12218);
nand U15800 (N_15800,N_14585,N_13798);
xnor U15801 (N_15801,N_12850,N_14389);
and U15802 (N_15802,N_13727,N_14785);
and U15803 (N_15803,N_13848,N_13916);
or U15804 (N_15804,N_13215,N_12988);
xor U15805 (N_15805,N_13903,N_13149);
nor U15806 (N_15806,N_12698,N_14214);
nand U15807 (N_15807,N_12145,N_14808);
xnor U15808 (N_15808,N_12268,N_14793);
and U15809 (N_15809,N_12426,N_12754);
and U15810 (N_15810,N_14019,N_12476);
or U15811 (N_15811,N_13014,N_14568);
and U15812 (N_15812,N_13482,N_14041);
nor U15813 (N_15813,N_14872,N_14657);
and U15814 (N_15814,N_12902,N_13735);
nor U15815 (N_15815,N_13202,N_13179);
or U15816 (N_15816,N_13784,N_13468);
or U15817 (N_15817,N_12636,N_12805);
nor U15818 (N_15818,N_13573,N_14976);
nand U15819 (N_15819,N_13461,N_13446);
nand U15820 (N_15820,N_12862,N_13329);
or U15821 (N_15821,N_13675,N_14825);
nor U15822 (N_15822,N_12798,N_12283);
nor U15823 (N_15823,N_12571,N_13414);
nor U15824 (N_15824,N_14098,N_13591);
xnor U15825 (N_15825,N_12332,N_12205);
nand U15826 (N_15826,N_12257,N_14561);
xnor U15827 (N_15827,N_13761,N_13622);
xnor U15828 (N_15828,N_13317,N_12931);
nand U15829 (N_15829,N_13749,N_13049);
or U15830 (N_15830,N_14688,N_14324);
nand U15831 (N_15831,N_14775,N_12792);
and U15832 (N_15832,N_13441,N_12625);
and U15833 (N_15833,N_13795,N_14893);
or U15834 (N_15834,N_14122,N_12576);
and U15835 (N_15835,N_13543,N_12005);
nand U15836 (N_15836,N_14138,N_12122);
or U15837 (N_15837,N_14018,N_14088);
nand U15838 (N_15838,N_12116,N_14057);
xor U15839 (N_15839,N_13152,N_12719);
nor U15840 (N_15840,N_14965,N_12921);
xnor U15841 (N_15841,N_12939,N_12611);
nand U15842 (N_15842,N_13561,N_12010);
xor U15843 (N_15843,N_12911,N_13974);
nand U15844 (N_15844,N_13181,N_13382);
and U15845 (N_15845,N_13363,N_13725);
xor U15846 (N_15846,N_13900,N_14944);
and U15847 (N_15847,N_13086,N_13150);
xnor U15848 (N_15848,N_14937,N_14604);
nand U15849 (N_15849,N_12181,N_13592);
or U15850 (N_15850,N_14696,N_13603);
nand U15851 (N_15851,N_12975,N_14979);
xnor U15852 (N_15852,N_14739,N_13051);
nor U15853 (N_15853,N_12162,N_13059);
nor U15854 (N_15854,N_14009,N_12886);
and U15855 (N_15855,N_13812,N_13901);
or U15856 (N_15856,N_14233,N_13384);
nor U15857 (N_15857,N_12322,N_12539);
or U15858 (N_15858,N_12076,N_12215);
xnor U15859 (N_15859,N_13041,N_12561);
xnor U15860 (N_15860,N_12148,N_14310);
nand U15861 (N_15861,N_14402,N_13986);
and U15862 (N_15862,N_12602,N_13793);
nor U15863 (N_15863,N_12631,N_12840);
and U15864 (N_15864,N_14614,N_13606);
nand U15865 (N_15865,N_12656,N_14544);
nor U15866 (N_15866,N_12389,N_14599);
nand U15867 (N_15867,N_13254,N_14234);
nor U15868 (N_15868,N_12909,N_12797);
and U15869 (N_15869,N_14038,N_14628);
and U15870 (N_15870,N_14136,N_12016);
xor U15871 (N_15871,N_12259,N_14316);
nor U15872 (N_15872,N_14522,N_12488);
xnor U15873 (N_15873,N_14797,N_14334);
xnor U15874 (N_15874,N_13023,N_13810);
or U15875 (N_15875,N_14472,N_12685);
nand U15876 (N_15876,N_14770,N_13851);
nand U15877 (N_15877,N_13588,N_13641);
or U15878 (N_15878,N_12842,N_14540);
xnor U15879 (N_15879,N_13779,N_14571);
nand U15880 (N_15880,N_13024,N_13413);
nand U15881 (N_15881,N_14925,N_14318);
nor U15882 (N_15882,N_14817,N_13759);
xor U15883 (N_15883,N_14556,N_14225);
nor U15884 (N_15884,N_13714,N_14668);
nand U15885 (N_15885,N_14689,N_14663);
xor U15886 (N_15886,N_14326,N_14124);
nand U15887 (N_15887,N_13029,N_12641);
nor U15888 (N_15888,N_13248,N_14071);
xor U15889 (N_15889,N_14570,N_13932);
nor U15890 (N_15890,N_13334,N_13495);
or U15891 (N_15891,N_12478,N_13695);
and U15892 (N_15892,N_12986,N_13632);
or U15893 (N_15893,N_14005,N_12849);
and U15894 (N_15894,N_12587,N_13670);
nand U15895 (N_15895,N_12935,N_13962);
xnor U15896 (N_15896,N_12693,N_13163);
nand U15897 (N_15897,N_12209,N_13444);
or U15898 (N_15898,N_13991,N_14185);
nor U15899 (N_15899,N_12030,N_12300);
or U15900 (N_15900,N_12454,N_12989);
xor U15901 (N_15901,N_12683,N_14081);
nor U15902 (N_15902,N_13268,N_14692);
or U15903 (N_15903,N_14921,N_12574);
nand U15904 (N_15904,N_14146,N_13616);
xor U15905 (N_15905,N_13845,N_13547);
nor U15906 (N_15906,N_14403,N_13381);
nand U15907 (N_15907,N_12291,N_13367);
and U15908 (N_15908,N_14458,N_14727);
nor U15909 (N_15909,N_14101,N_14575);
or U15910 (N_15910,N_13339,N_12348);
nand U15911 (N_15911,N_13058,N_13226);
or U15912 (N_15912,N_13623,N_12046);
nor U15913 (N_15913,N_12473,N_13343);
or U15914 (N_15914,N_12522,N_14076);
nand U15915 (N_15915,N_13445,N_12362);
xor U15916 (N_15916,N_14006,N_12513);
xor U15917 (N_15917,N_14178,N_12728);
xor U15918 (N_15918,N_12736,N_12727);
and U15919 (N_15919,N_12788,N_13057);
xnor U15920 (N_15920,N_12270,N_13400);
or U15921 (N_15921,N_12261,N_13500);
or U15922 (N_15922,N_13539,N_12136);
nor U15923 (N_15923,N_13088,N_13760);
nor U15924 (N_15924,N_14608,N_14899);
or U15925 (N_15925,N_14804,N_14955);
nor U15926 (N_15926,N_14974,N_13781);
or U15927 (N_15927,N_12532,N_13264);
nand U15928 (N_15928,N_14572,N_14518);
and U15929 (N_15929,N_12161,N_13116);
or U15930 (N_15930,N_13371,N_13599);
xnor U15931 (N_15931,N_13091,N_14769);
nand U15932 (N_15932,N_12868,N_12073);
or U15933 (N_15933,N_13977,N_12578);
nor U15934 (N_15934,N_13173,N_14205);
and U15935 (N_15935,N_13518,N_13061);
nor U15936 (N_15936,N_12721,N_13157);
or U15937 (N_15937,N_12780,N_13791);
nor U15938 (N_15938,N_13241,N_14301);
nand U15939 (N_15939,N_13610,N_13595);
and U15940 (N_15940,N_14208,N_13819);
or U15941 (N_15941,N_13927,N_13131);
nor U15942 (N_15942,N_12052,N_12167);
nor U15943 (N_15943,N_14008,N_13524);
and U15944 (N_15944,N_12403,N_13997);
nand U15945 (N_15945,N_14193,N_13278);
nand U15946 (N_15946,N_13020,N_12613);
nand U15947 (N_15947,N_12960,N_14369);
xor U15948 (N_15948,N_14664,N_14119);
nand U15949 (N_15949,N_12541,N_13552);
and U15950 (N_15950,N_12249,N_12412);
nand U15951 (N_15951,N_13294,N_13972);
nor U15952 (N_15952,N_12515,N_14866);
nand U15953 (N_15953,N_12766,N_12132);
or U15954 (N_15954,N_13550,N_13993);
nor U15955 (N_15955,N_13410,N_14248);
xor U15956 (N_15956,N_12195,N_12978);
nand U15957 (N_15957,N_14160,N_13366);
or U15958 (N_15958,N_14125,N_13849);
and U15959 (N_15959,N_13199,N_12629);
nor U15960 (N_15960,N_12669,N_14312);
nand U15961 (N_15961,N_13047,N_12919);
xnor U15962 (N_15962,N_12810,N_13256);
nand U15963 (N_15963,N_14245,N_12477);
nand U15964 (N_15964,N_14936,N_13855);
nand U15965 (N_15965,N_13242,N_13327);
nor U15966 (N_15966,N_14039,N_12885);
and U15967 (N_15967,N_14830,N_14314);
xnor U15968 (N_15968,N_14748,N_14459);
nand U15969 (N_15969,N_12857,N_14014);
nor U15970 (N_15970,N_12821,N_14415);
nand U15971 (N_15971,N_12106,N_12546);
and U15972 (N_15972,N_13834,N_12617);
nor U15973 (N_15973,N_12644,N_13585);
and U15974 (N_15974,N_14670,N_13249);
and U15975 (N_15975,N_13774,N_14888);
nand U15976 (N_15976,N_12047,N_13910);
nor U15977 (N_15977,N_14300,N_14706);
or U15978 (N_15978,N_14500,N_14487);
or U15979 (N_15979,N_14600,N_13562);
xor U15980 (N_15980,N_13536,N_13862);
nor U15981 (N_15981,N_12077,N_13039);
xnor U15982 (N_15982,N_12151,N_14554);
xor U15983 (N_15983,N_14835,N_14695);
or U15984 (N_15984,N_13003,N_12583);
nor U15985 (N_15985,N_13953,N_14384);
and U15986 (N_15986,N_13696,N_13171);
nor U15987 (N_15987,N_13868,N_12527);
xor U15988 (N_15988,N_12585,N_12096);
nand U15989 (N_15989,N_14110,N_12058);
xnor U15990 (N_15990,N_14987,N_13304);
nand U15991 (N_15991,N_14361,N_13873);
xnor U15992 (N_15992,N_14155,N_13631);
and U15993 (N_15993,N_13973,N_13998);
nand U15994 (N_15994,N_14702,N_13847);
and U15995 (N_15995,N_13840,N_13594);
or U15996 (N_15996,N_14210,N_14036);
or U15997 (N_15997,N_13665,N_13255);
or U15998 (N_15998,N_12284,N_12822);
xor U15999 (N_15999,N_13825,N_14602);
nor U16000 (N_16000,N_12764,N_14341);
nor U16001 (N_16001,N_14726,N_14885);
nand U16002 (N_16002,N_13100,N_14652);
xor U16003 (N_16003,N_13017,N_13929);
xor U16004 (N_16004,N_14799,N_12435);
and U16005 (N_16005,N_13483,N_13196);
or U16006 (N_16006,N_13666,N_13004);
and U16007 (N_16007,N_12240,N_12910);
or U16008 (N_16008,N_13144,N_14261);
xor U16009 (N_16009,N_13478,N_12244);
nor U16010 (N_16010,N_14741,N_12722);
and U16011 (N_16011,N_12637,N_13942);
and U16012 (N_16012,N_13809,N_12503);
and U16013 (N_16013,N_12102,N_13647);
and U16014 (N_16014,N_13001,N_14367);
nor U16015 (N_16015,N_13946,N_12339);
and U16016 (N_16016,N_14680,N_13211);
nand U16017 (N_16017,N_13505,N_12985);
or U16018 (N_16018,N_14539,N_13668);
xor U16019 (N_16019,N_14271,N_14485);
nand U16020 (N_16020,N_13887,N_14633);
xnor U16021 (N_16021,N_12725,N_12160);
nand U16022 (N_16022,N_13509,N_14994);
nand U16023 (N_16023,N_13279,N_13881);
nor U16024 (N_16024,N_12572,N_14285);
xor U16025 (N_16025,N_13333,N_13630);
or U16026 (N_16026,N_12039,N_14044);
or U16027 (N_16027,N_14000,N_13846);
nand U16028 (N_16028,N_12930,N_12856);
or U16029 (N_16029,N_13335,N_13209);
or U16030 (N_16030,N_12369,N_13220);
nand U16031 (N_16031,N_12818,N_14327);
or U16032 (N_16032,N_12650,N_13933);
nor U16033 (N_16033,N_12815,N_13753);
and U16034 (N_16034,N_14280,N_14481);
nor U16035 (N_16035,N_12020,N_14364);
or U16036 (N_16036,N_12556,N_12474);
nand U16037 (N_16037,N_14078,N_14489);
nand U16038 (N_16038,N_12318,N_12903);
and U16039 (N_16039,N_14503,N_13729);
nor U16040 (N_16040,N_13261,N_14740);
nor U16041 (N_16041,N_14293,N_12210);
nor U16042 (N_16042,N_14174,N_12321);
and U16043 (N_16043,N_12081,N_13046);
xor U16044 (N_16044,N_13554,N_14003);
or U16045 (N_16045,N_12958,N_12411);
or U16046 (N_16046,N_12365,N_14198);
nor U16047 (N_16047,N_12067,N_13045);
xnor U16048 (N_16048,N_12294,N_12694);
nand U16049 (N_16049,N_13127,N_13620);
nor U16050 (N_16050,N_13244,N_12942);
and U16051 (N_16051,N_14126,N_12565);
xor U16052 (N_16052,N_12008,N_12201);
and U16053 (N_16053,N_13541,N_12713);
nor U16054 (N_16054,N_13917,N_12834);
xnor U16055 (N_16055,N_14325,N_14836);
nand U16056 (N_16056,N_13783,N_14401);
nand U16057 (N_16057,N_13648,N_14330);
or U16058 (N_16058,N_14512,N_14698);
nor U16059 (N_16059,N_14308,N_13629);
and U16060 (N_16060,N_14483,N_13316);
nor U16061 (N_16061,N_12086,N_14063);
and U16062 (N_16062,N_14903,N_13904);
xor U16063 (N_16063,N_12180,N_12863);
xnor U16064 (N_16064,N_12425,N_12475);
nor U16065 (N_16065,N_12582,N_13584);
nor U16066 (N_16066,N_13147,N_12543);
or U16067 (N_16067,N_13600,N_13151);
or U16068 (N_16068,N_14579,N_13153);
nor U16069 (N_16069,N_14819,N_12439);
and U16070 (N_16070,N_13939,N_14232);
or U16071 (N_16071,N_13074,N_14253);
nand U16072 (N_16072,N_13801,N_13689);
nor U16073 (N_16073,N_12272,N_12956);
xor U16074 (N_16074,N_14700,N_13323);
or U16075 (N_16075,N_13299,N_14978);
xnor U16076 (N_16076,N_14460,N_13346);
or U16077 (N_16077,N_13013,N_12456);
xnor U16078 (N_16078,N_12775,N_13645);
nor U16079 (N_16079,N_12916,N_12377);
or U16080 (N_16080,N_14230,N_12429);
and U16081 (N_16081,N_14256,N_13031);
xor U16082 (N_16082,N_13677,N_13063);
and U16083 (N_16083,N_13422,N_12324);
nand U16084 (N_16084,N_14226,N_12955);
or U16085 (N_16085,N_13597,N_14792);
nor U16086 (N_16086,N_12836,N_12954);
or U16087 (N_16087,N_13193,N_12860);
nand U16088 (N_16088,N_12529,N_13307);
nor U16089 (N_16089,N_13843,N_13590);
and U16090 (N_16090,N_13286,N_12043);
and U16091 (N_16091,N_13387,N_13776);
or U16092 (N_16092,N_12531,N_13113);
xnor U16093 (N_16093,N_13230,N_13488);
xnor U16094 (N_16094,N_12595,N_12131);
nor U16095 (N_16095,N_12179,N_14796);
xnor U16096 (N_16096,N_14543,N_13036);
or U16097 (N_16097,N_12658,N_14106);
nand U16098 (N_16098,N_12559,N_13726);
or U16099 (N_16099,N_12216,N_12628);
and U16100 (N_16100,N_13731,N_12855);
or U16101 (N_16101,N_14315,N_14042);
or U16102 (N_16102,N_13101,N_14705);
nor U16103 (N_16103,N_12224,N_14982);
and U16104 (N_16104,N_13472,N_12813);
and U16105 (N_16105,N_13355,N_12976);
xnor U16106 (N_16106,N_14881,N_14772);
nand U16107 (N_16107,N_14686,N_12298);
nand U16108 (N_16108,N_12575,N_14453);
xnor U16109 (N_16109,N_13678,N_13233);
nand U16110 (N_16110,N_14878,N_14273);
and U16111 (N_16111,N_13296,N_14901);
nand U16112 (N_16112,N_13975,N_14499);
and U16113 (N_16113,N_12119,N_12254);
nor U16114 (N_16114,N_13089,N_13205);
nand U16115 (N_16115,N_13970,N_14989);
xnor U16116 (N_16116,N_14058,N_13109);
xnor U16117 (N_16117,N_14504,N_13564);
or U16118 (N_16118,N_13425,N_14988);
and U16119 (N_16119,N_14678,N_14779);
and U16120 (N_16120,N_13867,N_14605);
nor U16121 (N_16121,N_13984,N_12779);
nor U16122 (N_16122,N_13913,N_14743);
xor U16123 (N_16123,N_12761,N_14352);
xor U16124 (N_16124,N_13935,N_14069);
nand U16125 (N_16125,N_13287,N_12832);
nor U16126 (N_16126,N_12553,N_14366);
or U16127 (N_16127,N_12350,N_14123);
xnor U16128 (N_16128,N_13792,N_12876);
and U16129 (N_16129,N_13911,N_14707);
or U16130 (N_16130,N_13365,N_13391);
nand U16131 (N_16131,N_12922,N_13188);
xor U16132 (N_16132,N_14886,N_12128);
nand U16133 (N_16133,N_14865,N_14710);
or U16134 (N_16134,N_12804,N_14721);
nand U16135 (N_16135,N_12653,N_13439);
nor U16136 (N_16136,N_12343,N_12623);
and U16137 (N_16137,N_12824,N_12777);
or U16138 (N_16138,N_14694,N_13467);
and U16139 (N_16139,N_14826,N_14593);
nor U16140 (N_16140,N_13284,N_14439);
and U16141 (N_16141,N_14302,N_14051);
and U16142 (N_16142,N_14934,N_14521);
and U16143 (N_16143,N_12646,N_12226);
or U16144 (N_16144,N_13143,N_14207);
and U16145 (N_16145,N_13078,N_12507);
xnor U16146 (N_16146,N_13553,N_12701);
nand U16147 (N_16147,N_14644,N_14231);
or U16148 (N_16148,N_14397,N_14002);
or U16149 (N_16149,N_14242,N_13602);
or U16150 (N_16150,N_13912,N_14909);
nor U16151 (N_16151,N_13990,N_14832);
xor U16152 (N_16152,N_13340,N_13961);
and U16153 (N_16153,N_12396,N_12279);
nand U16154 (N_16154,N_12099,N_12394);
nor U16155 (N_16155,N_13243,N_12469);
xor U16156 (N_16156,N_12271,N_12087);
or U16157 (N_16157,N_13009,N_12453);
nand U16158 (N_16158,N_13095,N_13635);
nand U16159 (N_16159,N_12542,N_14218);
xor U16160 (N_16160,N_14445,N_12054);
nand U16161 (N_16161,N_14854,N_13110);
and U16162 (N_16162,N_13455,N_13289);
or U16163 (N_16163,N_12994,N_12943);
or U16164 (N_16164,N_13948,N_13347);
and U16165 (N_16165,N_14777,N_14368);
nand U16166 (N_16166,N_13717,N_13653);
xnor U16167 (N_16167,N_13450,N_14736);
or U16168 (N_16168,N_12380,N_14564);
and U16169 (N_16169,N_13969,N_12238);
xnor U16170 (N_16170,N_13806,N_12704);
xnor U16171 (N_16171,N_14824,N_14115);
and U16172 (N_16172,N_12042,N_14735);
or U16173 (N_16173,N_12185,N_12278);
xnor U16174 (N_16174,N_14669,N_14012);
nand U16175 (N_16175,N_13836,N_14040);
or U16176 (N_16176,N_14015,N_12630);
nor U16177 (N_16177,N_14932,N_14220);
nand U16178 (N_16178,N_12275,N_14390);
or U16179 (N_16179,N_12643,N_14949);
nand U16180 (N_16180,N_13878,N_12314);
nand U16181 (N_16181,N_13551,N_14541);
nand U16182 (N_16182,N_12604,N_13406);
xnor U16183 (N_16183,N_14130,N_14222);
nor U16184 (N_16184,N_14587,N_14482);
xor U16185 (N_16185,N_13835,N_13126);
or U16186 (N_16186,N_14583,N_14030);
nand U16187 (N_16187,N_14671,N_13639);
nor U16188 (N_16188,N_14889,N_12184);
xnor U16189 (N_16189,N_12672,N_14349);
xnor U16190 (N_16190,N_12241,N_14034);
nand U16191 (N_16191,N_12233,N_12384);
nor U16192 (N_16192,N_14510,N_12035);
nand U16193 (N_16193,N_13321,N_13674);
nand U16194 (N_16194,N_14545,N_14392);
or U16195 (N_16195,N_13373,N_14547);
or U16196 (N_16196,N_14717,N_14578);
nand U16197 (N_16197,N_12786,N_14874);
nor U16198 (N_16198,N_12260,N_13768);
xor U16199 (N_16199,N_13898,N_14121);
or U16200 (N_16200,N_14591,N_14342);
nand U16201 (N_16201,N_13859,N_14080);
nand U16202 (N_16202,N_13454,N_12055);
nor U16203 (N_16203,N_12590,N_12340);
nor U16204 (N_16204,N_12485,N_12627);
nand U16205 (N_16205,N_12405,N_12309);
xnor U16206 (N_16206,N_14269,N_13451);
nand U16207 (N_16207,N_12530,N_14699);
nand U16208 (N_16208,N_12951,N_12889);
xor U16209 (N_16209,N_14215,N_13208);
nand U16210 (N_16210,N_13521,N_14363);
nor U16211 (N_16211,N_13466,N_14219);
or U16212 (N_16212,N_13397,N_12153);
nor U16213 (N_16213,N_14167,N_12703);
xnor U16214 (N_16214,N_13876,N_14348);
nand U16215 (N_16215,N_12538,N_13477);
xnor U16216 (N_16216,N_14910,N_13221);
nor U16217 (N_16217,N_14360,N_13664);
nand U16218 (N_16218,N_14282,N_12695);
xnor U16219 (N_16219,N_13118,N_12748);
or U16220 (N_16220,N_14351,N_14086);
xor U16221 (N_16221,N_13084,N_14873);
xnor U16222 (N_16222,N_13102,N_13415);
and U16223 (N_16223,N_13660,N_13709);
nor U16224 (N_16224,N_13262,N_12665);
nand U16225 (N_16225,N_13718,N_12948);
nor U16226 (N_16226,N_13852,N_12914);
or U16227 (N_16227,N_12164,N_12901);
nor U16228 (N_16228,N_14028,N_12952);
nand U16229 (N_16229,N_12277,N_13460);
or U16230 (N_16230,N_13246,N_13174);
xnor U16231 (N_16231,N_14525,N_14370);
and U16232 (N_16232,N_12163,N_12998);
xor U16233 (N_16233,N_14437,N_12620);
nand U16234 (N_16234,N_12230,N_12586);
and U16235 (N_16235,N_13838,N_13737);
nor U16236 (N_16236,N_13369,N_12438);
and U16237 (N_16237,N_13229,N_12523);
nand U16238 (N_16238,N_12520,N_14730);
and U16239 (N_16239,N_12349,N_14413);
or U16240 (N_16240,N_14433,N_12123);
xor U16241 (N_16241,N_12509,N_12378);
or U16242 (N_16242,N_13194,N_14421);
nor U16243 (N_16243,N_13934,N_13030);
and U16244 (N_16244,N_12492,N_14745);
and U16245 (N_16245,N_13748,N_12853);
xnor U16246 (N_16246,N_14148,N_12173);
and U16247 (N_16247,N_14990,N_12781);
or U16248 (N_16248,N_12217,N_14848);
and U16249 (N_16249,N_13667,N_13239);
and U16250 (N_16250,N_14980,N_12544);
nand U16251 (N_16251,N_13297,N_12146);
nand U16252 (N_16252,N_12135,N_14917);
nor U16253 (N_16253,N_14298,N_12045);
and U16254 (N_16254,N_14430,N_14446);
or U16255 (N_16255,N_12355,N_12208);
nor U16256 (N_16256,N_14407,N_14378);
xnor U16257 (N_16257,N_13099,N_14513);
nor U16258 (N_16258,N_14634,N_12537);
or U16259 (N_16259,N_12887,N_12235);
nor U16260 (N_16260,N_13138,N_13276);
and U16261 (N_16261,N_12115,N_12207);
or U16262 (N_16262,N_12462,N_14618);
and U16263 (N_16263,N_13931,N_12419);
nor U16264 (N_16264,N_14879,N_14679);
and U16265 (N_16265,N_12907,N_12025);
nand U16266 (N_16266,N_12897,N_12246);
and U16267 (N_16267,N_13905,N_12738);
xor U16268 (N_16268,N_14720,N_13775);
and U16269 (N_16269,N_14175,N_12687);
nand U16270 (N_16270,N_14180,N_14687);
nand U16271 (N_16271,N_13956,N_13814);
and U16272 (N_16272,N_14732,N_12442);
xnor U16273 (N_16273,N_14958,N_12415);
nor U16274 (N_16274,N_13655,N_14031);
or U16275 (N_16275,N_13520,N_12589);
or U16276 (N_16276,N_14725,N_14661);
nor U16277 (N_16277,N_13310,N_13185);
nor U16278 (N_16278,N_14414,N_14183);
or U16279 (N_16279,N_14131,N_12288);
and U16280 (N_16280,N_14635,N_12536);
and U16281 (N_16281,N_13337,N_14841);
xnor U16282 (N_16282,N_14427,N_13177);
or U16283 (N_16283,N_13125,N_12566);
or U16284 (N_16284,N_13496,N_14474);
nand U16285 (N_16285,N_14317,N_14281);
or U16286 (N_16286,N_13311,N_14722);
nand U16287 (N_16287,N_14675,N_12141);
and U16288 (N_16288,N_12753,N_14494);
and U16289 (N_16289,N_14648,N_12436);
nor U16290 (N_16290,N_12987,N_13132);
and U16291 (N_16291,N_12675,N_14197);
nand U16292 (N_16292,N_13751,N_12733);
xnor U16293 (N_16293,N_12445,N_14020);
nor U16294 (N_16294,N_13512,N_12306);
or U16295 (N_16295,N_13527,N_12007);
nor U16296 (N_16296,N_14716,N_14546);
nand U16297 (N_16297,N_12896,N_12642);
or U16298 (N_16298,N_14252,N_14517);
xor U16299 (N_16299,N_14188,N_13549);
xor U16300 (N_16300,N_12386,N_12169);
or U16301 (N_16301,N_13203,N_13250);
or U16302 (N_16302,N_13740,N_12188);
nor U16303 (N_16303,N_12075,N_13115);
or U16304 (N_16304,N_12422,N_14294);
nor U16305 (N_16305,N_12464,N_14478);
and U16306 (N_16306,N_14333,N_13516);
nor U16307 (N_16307,N_14981,N_14394);
nand U16308 (N_16308,N_12433,N_13038);
xor U16309 (N_16309,N_12516,N_13493);
or U16310 (N_16310,N_13476,N_12533);
and U16311 (N_16311,N_12420,N_14179);
or U16312 (N_16312,N_14860,N_14630);
xor U16313 (N_16313,N_14074,N_12228);
nor U16314 (N_16314,N_14385,N_12661);
nand U16315 (N_16315,N_14075,N_13266);
nand U16316 (N_16316,N_14295,N_14954);
and U16317 (N_16317,N_14565,N_12457);
nand U16318 (N_16318,N_12501,N_13959);
nand U16319 (N_16319,N_14498,N_12051);
nor U16320 (N_16320,N_14182,N_14764);
and U16321 (N_16321,N_12206,N_13054);
nand U16322 (N_16322,N_12263,N_13832);
nor U16323 (N_16323,N_13463,N_13416);
and U16324 (N_16324,N_12519,N_14082);
xor U16325 (N_16325,N_13453,N_13830);
xor U16326 (N_16326,N_14164,N_12933);
or U16327 (N_16327,N_13274,N_14393);
nand U16328 (N_16328,N_14192,N_14852);
xor U16329 (N_16329,N_12965,N_14203);
nor U16330 (N_16330,N_12967,N_14161);
nor U16331 (N_16331,N_12312,N_14238);
xor U16332 (N_16332,N_14307,N_12564);
nor U16333 (N_16333,N_14821,N_12550);
nor U16334 (N_16334,N_14235,N_13015);
nor U16335 (N_16335,N_13201,N_12898);
xor U16336 (N_16336,N_12890,N_14471);
nand U16337 (N_16337,N_12662,N_13016);
and U16338 (N_16338,N_14928,N_13350);
and U16339 (N_16339,N_13071,N_14560);
nand U16340 (N_16340,N_13950,N_13804);
nor U16341 (N_16341,N_13352,N_12082);
xor U16342 (N_16342,N_14163,N_13983);
and U16343 (N_16343,N_14900,N_14919);
or U16344 (N_16344,N_14842,N_13833);
or U16345 (N_16345,N_14443,N_14867);
and U16346 (N_16346,N_14347,N_14534);
nand U16347 (N_16347,N_14213,N_13909);
or U16348 (N_16348,N_14150,N_12674);
nor U16349 (N_16349,N_12926,N_12610);
nor U16350 (N_16350,N_14380,N_14428);
xor U16351 (N_16351,N_14642,N_13281);
nor U16352 (N_16352,N_12937,N_13168);
and U16353 (N_16353,N_14685,N_13892);
nor U16354 (N_16354,N_12635,N_13360);
nor U16355 (N_16355,N_13056,N_13485);
nor U16356 (N_16356,N_13854,N_12618);
or U16357 (N_16357,N_12534,N_13145);
or U16358 (N_16358,N_14789,N_12059);
nor U16359 (N_16359,N_12999,N_12074);
or U16360 (N_16360,N_13283,N_13136);
and U16361 (N_16361,N_13314,N_13232);
nor U16362 (N_16362,N_12769,N_13253);
nand U16363 (N_16363,N_12194,N_14372);
nand U16364 (N_16364,N_13937,N_14930);
xor U16365 (N_16365,N_12731,N_12495);
nor U16366 (N_16366,N_14137,N_12645);
nor U16367 (N_16367,N_12176,N_12591);
or U16368 (N_16368,N_13649,N_12982);
or U16369 (N_16369,N_13124,N_14863);
nand U16370 (N_16370,N_12841,N_14586);
or U16371 (N_16371,N_14527,N_12418);
nor U16372 (N_16372,N_14016,N_14946);
nand U16373 (N_16373,N_14538,N_13989);
nor U16374 (N_16374,N_12634,N_12594);
xnor U16375 (N_16375,N_13263,N_13247);
nor U16376 (N_16376,N_12103,N_14746);
nor U16377 (N_16377,N_14509,N_14884);
nor U16378 (N_16378,N_12770,N_14304);
xor U16379 (N_16379,N_12383,N_13172);
xnor U16380 (N_16380,N_14929,N_13706);
nor U16381 (N_16381,N_13712,N_14828);
nand U16382 (N_16382,N_12434,N_13409);
xnor U16383 (N_16383,N_14507,N_13358);
nand U16384 (N_16384,N_13498,N_13213);
xnor U16385 (N_16385,N_14477,N_13921);
nand U16386 (N_16386,N_13540,N_13225);
and U16387 (N_16387,N_12034,N_12991);
and U16388 (N_16388,N_13417,N_14373);
and U16389 (N_16389,N_13763,N_13164);
and U16390 (N_16390,N_13767,N_13357);
nand U16391 (N_16391,N_13860,N_13531);
or U16392 (N_16392,N_12521,N_12600);
and U16393 (N_16393,N_14484,N_12794);
nand U16394 (N_16394,N_13035,N_12825);
nand U16395 (N_16395,N_12198,N_14055);
xnor U16396 (N_16396,N_14551,N_14774);
nand U16397 (N_16397,N_12562,N_12108);
nor U16398 (N_16398,N_14107,N_14574);
or U16399 (N_16399,N_13259,N_13018);
xnor U16400 (N_16400,N_12979,N_14998);
and U16401 (N_16401,N_12483,N_12366);
xnor U16402 (N_16402,N_12014,N_14597);
or U16403 (N_16403,N_12381,N_12800);
nor U16404 (N_16404,N_12540,N_12158);
nand U16405 (N_16405,N_14023,N_14890);
xor U16406 (N_16406,N_12019,N_12370);
or U16407 (N_16407,N_12580,N_14961);
nor U16408 (N_16408,N_13988,N_12874);
nor U16409 (N_16409,N_14090,N_14719);
and U16410 (N_16410,N_13377,N_12601);
xor U16411 (N_16411,N_13787,N_13271);
and U16412 (N_16412,N_14145,N_14187);
nor U16413 (N_16413,N_13322,N_14731);
and U16414 (N_16414,N_12782,N_14170);
or U16415 (N_16415,N_14995,N_14948);
nor U16416 (N_16416,N_13980,N_14542);
xor U16417 (N_16417,N_13452,N_14111);
nand U16418 (N_16418,N_12231,N_13657);
xnor U16419 (N_16419,N_13853,N_14665);
nor U16420 (N_16420,N_13930,N_13240);
nand U16421 (N_16421,N_14475,N_13424);
nor U16422 (N_16422,N_12969,N_14412);
xnor U16423 (N_16423,N_12032,N_14941);
nor U16424 (N_16424,N_13750,N_13432);
and U16425 (N_16425,N_14892,N_13270);
nor U16426 (N_16426,N_14567,N_14713);
nor U16427 (N_16427,N_13662,N_14267);
and U16428 (N_16428,N_12746,N_13771);
nor U16429 (N_16429,N_13924,N_14017);
nor U16430 (N_16430,N_14060,N_12783);
nand U16431 (N_16431,N_12654,N_12388);
or U16432 (N_16432,N_12899,N_12317);
nor U16433 (N_16433,N_13169,N_14636);
nor U16434 (N_16434,N_14566,N_13484);
and U16435 (N_16435,N_13277,N_14905);
and U16436 (N_16436,N_12311,N_14968);
and U16437 (N_16437,N_12632,N_13433);
or U16438 (N_16438,N_12881,N_13034);
and U16439 (N_16439,N_12392,N_14410);
nand U16440 (N_16440,N_12408,N_13252);
xnor U16441 (N_16441,N_14371,N_14166);
nor U16442 (N_16442,N_12831,N_14381);
xor U16443 (N_16443,N_13557,N_12605);
and U16444 (N_16444,N_14582,N_14268);
and U16445 (N_16445,N_13766,N_12784);
or U16446 (N_16446,N_12744,N_12427);
xor U16447 (N_16447,N_13642,N_14291);
and U16448 (N_16448,N_14237,N_13081);
nand U16449 (N_16449,N_14615,N_14856);
or U16450 (N_16450,N_13308,N_14440);
nor U16451 (N_16451,N_12114,N_12968);
and U16452 (N_16452,N_14912,N_13469);
or U16453 (N_16453,N_13142,N_13506);
xor U16454 (N_16454,N_14753,N_14911);
xor U16455 (N_16455,N_12801,N_12390);
and U16456 (N_16456,N_12091,N_12936);
and U16457 (N_16457,N_14983,N_13656);
nand U16458 (N_16458,N_14938,N_13077);
xor U16459 (N_16459,N_12393,N_13085);
and U16460 (N_16460,N_13044,N_14181);
and U16461 (N_16461,N_13122,N_12626);
xor U16462 (N_16462,N_13407,N_12186);
nor U16463 (N_16463,N_14528,N_12125);
xnor U16464 (N_16464,N_12323,N_12302);
nor U16465 (N_16465,N_13625,N_13007);
xnor U16466 (N_16466,N_14734,N_12280);
or U16467 (N_16467,N_12274,N_12688);
xor U16468 (N_16468,N_14907,N_14249);
and U16469 (N_16469,N_14623,N_13428);
or U16470 (N_16470,N_13530,N_13312);
nor U16471 (N_16471,N_12820,N_12358);
and U16472 (N_16472,N_12089,N_12680);
nand U16473 (N_16473,N_14396,N_12093);
nor U16474 (N_16474,N_13141,N_12113);
or U16475 (N_16475,N_14152,N_14127);
and U16476 (N_16476,N_12072,N_13291);
nor U16477 (N_16477,N_14898,N_13829);
or U16478 (N_16478,N_14283,N_12732);
xor U16479 (N_16479,N_14607,N_14287);
nand U16480 (N_16480,N_13636,N_13888);
and U16481 (N_16481,N_12990,N_12996);
nor U16482 (N_16482,N_13344,N_13419);
or U16483 (N_16483,N_12981,N_13408);
xor U16484 (N_16484,N_13362,N_12053);
and U16485 (N_16485,N_13954,N_12193);
xor U16486 (N_16486,N_12854,N_14915);
nor U16487 (N_16487,N_13178,N_13092);
and U16488 (N_16488,N_12963,N_14264);
xor U16489 (N_16489,N_12900,N_14971);
nand U16490 (N_16490,N_13055,N_13423);
and U16491 (N_16491,N_13566,N_12934);
nor U16492 (N_16492,N_12878,N_14843);
nor U16493 (N_16493,N_14562,N_14709);
xnor U16494 (N_16494,N_12718,N_14073);
and U16495 (N_16495,N_12009,N_13701);
and U16496 (N_16496,N_13694,N_13189);
or U16497 (N_16497,N_14162,N_13320);
and U16498 (N_16498,N_12755,N_14945);
xnor U16499 (N_16499,N_13399,N_13572);
nand U16500 (N_16500,N_13362,N_12041);
and U16501 (N_16501,N_14243,N_13845);
and U16502 (N_16502,N_14887,N_13947);
and U16503 (N_16503,N_13515,N_13145);
nand U16504 (N_16504,N_14097,N_12771);
xnor U16505 (N_16505,N_14870,N_12928);
nand U16506 (N_16506,N_12670,N_12027);
nor U16507 (N_16507,N_13788,N_13174);
nor U16508 (N_16508,N_12010,N_14330);
and U16509 (N_16509,N_14448,N_13837);
or U16510 (N_16510,N_13726,N_13919);
or U16511 (N_16511,N_12487,N_14224);
xor U16512 (N_16512,N_12904,N_14414);
and U16513 (N_16513,N_13208,N_13449);
or U16514 (N_16514,N_12796,N_12043);
nor U16515 (N_16515,N_13563,N_14104);
and U16516 (N_16516,N_12529,N_12931);
xor U16517 (N_16517,N_13252,N_14443);
xor U16518 (N_16518,N_12106,N_13584);
xnor U16519 (N_16519,N_14744,N_14674);
nor U16520 (N_16520,N_12808,N_13061);
and U16521 (N_16521,N_12296,N_13808);
or U16522 (N_16522,N_14184,N_14573);
or U16523 (N_16523,N_14743,N_12629);
xor U16524 (N_16524,N_12600,N_14945);
xor U16525 (N_16525,N_14068,N_14256);
and U16526 (N_16526,N_14796,N_14034);
xnor U16527 (N_16527,N_12970,N_12414);
nor U16528 (N_16528,N_14519,N_12704);
or U16529 (N_16529,N_12472,N_14212);
and U16530 (N_16530,N_12389,N_12868);
or U16531 (N_16531,N_12975,N_12580);
nor U16532 (N_16532,N_14833,N_13776);
or U16533 (N_16533,N_14461,N_14935);
and U16534 (N_16534,N_14911,N_13209);
and U16535 (N_16535,N_13351,N_13201);
nor U16536 (N_16536,N_12708,N_12521);
xnor U16537 (N_16537,N_14168,N_13624);
and U16538 (N_16538,N_14774,N_14779);
xor U16539 (N_16539,N_12253,N_14327);
or U16540 (N_16540,N_14497,N_14390);
or U16541 (N_16541,N_12824,N_14190);
nand U16542 (N_16542,N_13548,N_12688);
xnor U16543 (N_16543,N_14585,N_14095);
xor U16544 (N_16544,N_13840,N_14707);
nand U16545 (N_16545,N_14354,N_14660);
and U16546 (N_16546,N_14580,N_13860);
xnor U16547 (N_16547,N_13808,N_13904);
nand U16548 (N_16548,N_12243,N_12770);
nand U16549 (N_16549,N_14008,N_12266);
and U16550 (N_16550,N_14718,N_14703);
or U16551 (N_16551,N_13131,N_13426);
xor U16552 (N_16552,N_14411,N_12957);
and U16553 (N_16553,N_14208,N_12605);
or U16554 (N_16554,N_12008,N_13823);
or U16555 (N_16555,N_14409,N_12448);
nand U16556 (N_16556,N_14482,N_14914);
nand U16557 (N_16557,N_14961,N_12022);
and U16558 (N_16558,N_12770,N_13424);
nor U16559 (N_16559,N_12034,N_13965);
nand U16560 (N_16560,N_14299,N_13635);
and U16561 (N_16561,N_12114,N_14396);
nor U16562 (N_16562,N_13273,N_12971);
and U16563 (N_16563,N_14868,N_14057);
nand U16564 (N_16564,N_14862,N_12359);
and U16565 (N_16565,N_13030,N_13267);
nand U16566 (N_16566,N_13020,N_13241);
nand U16567 (N_16567,N_14090,N_13116);
nor U16568 (N_16568,N_12104,N_13812);
nand U16569 (N_16569,N_12080,N_14917);
nor U16570 (N_16570,N_14649,N_12029);
nor U16571 (N_16571,N_14227,N_12373);
and U16572 (N_16572,N_14429,N_14188);
xor U16573 (N_16573,N_14624,N_14626);
nor U16574 (N_16574,N_14468,N_12026);
nor U16575 (N_16575,N_12742,N_13723);
and U16576 (N_16576,N_13442,N_14099);
or U16577 (N_16577,N_14634,N_14942);
and U16578 (N_16578,N_12715,N_14283);
nor U16579 (N_16579,N_14593,N_14539);
nor U16580 (N_16580,N_13692,N_13068);
or U16581 (N_16581,N_14929,N_14620);
nor U16582 (N_16582,N_14195,N_14271);
xnor U16583 (N_16583,N_12497,N_13333);
nor U16584 (N_16584,N_12582,N_12998);
and U16585 (N_16585,N_14576,N_14326);
xor U16586 (N_16586,N_12885,N_12124);
nor U16587 (N_16587,N_13472,N_13612);
and U16588 (N_16588,N_12227,N_14216);
nand U16589 (N_16589,N_12213,N_14724);
and U16590 (N_16590,N_12081,N_13076);
nand U16591 (N_16591,N_13950,N_12368);
or U16592 (N_16592,N_13526,N_12384);
nand U16593 (N_16593,N_14846,N_14243);
nand U16594 (N_16594,N_14881,N_14731);
or U16595 (N_16595,N_14120,N_12231);
and U16596 (N_16596,N_14972,N_13234);
or U16597 (N_16597,N_13812,N_12249);
or U16598 (N_16598,N_12853,N_14873);
nor U16599 (N_16599,N_13219,N_13096);
xor U16600 (N_16600,N_14089,N_14090);
xnor U16601 (N_16601,N_14992,N_14659);
or U16602 (N_16602,N_14825,N_12673);
and U16603 (N_16603,N_14617,N_12115);
and U16604 (N_16604,N_13767,N_13137);
nor U16605 (N_16605,N_14710,N_14115);
or U16606 (N_16606,N_12364,N_12181);
nand U16607 (N_16607,N_14406,N_14701);
xnor U16608 (N_16608,N_14905,N_13871);
and U16609 (N_16609,N_12453,N_12352);
and U16610 (N_16610,N_13586,N_13034);
nand U16611 (N_16611,N_13806,N_13655);
xor U16612 (N_16612,N_13379,N_12823);
or U16613 (N_16613,N_14376,N_14193);
or U16614 (N_16614,N_14470,N_12809);
nand U16615 (N_16615,N_12790,N_13546);
xor U16616 (N_16616,N_12785,N_13746);
nand U16617 (N_16617,N_14730,N_13032);
xor U16618 (N_16618,N_14943,N_12663);
and U16619 (N_16619,N_13399,N_14982);
xnor U16620 (N_16620,N_12701,N_12050);
and U16621 (N_16621,N_14874,N_12759);
nor U16622 (N_16622,N_12535,N_12787);
nand U16623 (N_16623,N_12372,N_14762);
xnor U16624 (N_16624,N_12097,N_13191);
nand U16625 (N_16625,N_12552,N_12212);
or U16626 (N_16626,N_13188,N_13740);
or U16627 (N_16627,N_13301,N_12861);
nand U16628 (N_16628,N_14034,N_12542);
nand U16629 (N_16629,N_12982,N_13407);
nand U16630 (N_16630,N_12359,N_14589);
xor U16631 (N_16631,N_12714,N_13183);
xor U16632 (N_16632,N_12998,N_13869);
nand U16633 (N_16633,N_14880,N_14483);
nand U16634 (N_16634,N_14505,N_12921);
xnor U16635 (N_16635,N_12372,N_14942);
nand U16636 (N_16636,N_13039,N_12029);
nor U16637 (N_16637,N_14680,N_12388);
nand U16638 (N_16638,N_13591,N_12763);
xnor U16639 (N_16639,N_14547,N_13468);
nor U16640 (N_16640,N_14844,N_14203);
nor U16641 (N_16641,N_13236,N_12856);
nand U16642 (N_16642,N_12812,N_13677);
and U16643 (N_16643,N_13930,N_14166);
and U16644 (N_16644,N_13193,N_13710);
nand U16645 (N_16645,N_12275,N_12668);
or U16646 (N_16646,N_12953,N_13365);
xor U16647 (N_16647,N_14820,N_12976);
nor U16648 (N_16648,N_12531,N_14329);
or U16649 (N_16649,N_12858,N_13600);
nor U16650 (N_16650,N_12876,N_12958);
or U16651 (N_16651,N_14400,N_12209);
nand U16652 (N_16652,N_12411,N_13343);
nand U16653 (N_16653,N_12971,N_12388);
and U16654 (N_16654,N_14424,N_12957);
and U16655 (N_16655,N_12014,N_13716);
or U16656 (N_16656,N_13210,N_13258);
or U16657 (N_16657,N_12785,N_13870);
nand U16658 (N_16658,N_12742,N_14218);
nand U16659 (N_16659,N_12181,N_12506);
nand U16660 (N_16660,N_13473,N_13869);
or U16661 (N_16661,N_12901,N_12447);
and U16662 (N_16662,N_13449,N_12272);
and U16663 (N_16663,N_14572,N_12102);
nor U16664 (N_16664,N_12787,N_13072);
xor U16665 (N_16665,N_13094,N_13629);
nand U16666 (N_16666,N_12344,N_14492);
and U16667 (N_16667,N_14599,N_13636);
or U16668 (N_16668,N_14895,N_14391);
and U16669 (N_16669,N_14469,N_14971);
xor U16670 (N_16670,N_14467,N_12159);
or U16671 (N_16671,N_12068,N_14622);
xnor U16672 (N_16672,N_14977,N_12113);
xor U16673 (N_16673,N_14566,N_12664);
nor U16674 (N_16674,N_14881,N_12942);
nor U16675 (N_16675,N_14385,N_12589);
xor U16676 (N_16676,N_13974,N_13049);
and U16677 (N_16677,N_14419,N_12375);
nor U16678 (N_16678,N_12317,N_13097);
nand U16679 (N_16679,N_14327,N_12712);
and U16680 (N_16680,N_12963,N_13726);
nand U16681 (N_16681,N_14872,N_14154);
or U16682 (N_16682,N_13807,N_12793);
nand U16683 (N_16683,N_13718,N_14336);
nand U16684 (N_16684,N_13159,N_12427);
and U16685 (N_16685,N_14626,N_13472);
xnor U16686 (N_16686,N_14203,N_13854);
xor U16687 (N_16687,N_13510,N_13341);
nor U16688 (N_16688,N_12531,N_12698);
and U16689 (N_16689,N_13744,N_12125);
nand U16690 (N_16690,N_12667,N_14602);
and U16691 (N_16691,N_14496,N_14066);
nand U16692 (N_16692,N_13984,N_14544);
xor U16693 (N_16693,N_12553,N_13329);
and U16694 (N_16694,N_13028,N_13965);
and U16695 (N_16695,N_12527,N_13128);
and U16696 (N_16696,N_12368,N_12092);
and U16697 (N_16697,N_13030,N_13410);
and U16698 (N_16698,N_13940,N_14014);
or U16699 (N_16699,N_12431,N_12010);
or U16700 (N_16700,N_13992,N_14102);
xnor U16701 (N_16701,N_13848,N_13492);
xor U16702 (N_16702,N_12646,N_14008);
nand U16703 (N_16703,N_13252,N_12828);
nand U16704 (N_16704,N_12053,N_12072);
xnor U16705 (N_16705,N_13505,N_12710);
xor U16706 (N_16706,N_14505,N_12691);
and U16707 (N_16707,N_14818,N_14842);
nor U16708 (N_16708,N_13965,N_12262);
xnor U16709 (N_16709,N_14473,N_13290);
xor U16710 (N_16710,N_12053,N_14705);
nand U16711 (N_16711,N_14785,N_14134);
nand U16712 (N_16712,N_13951,N_12368);
nand U16713 (N_16713,N_14237,N_13034);
nand U16714 (N_16714,N_14649,N_14505);
xnor U16715 (N_16715,N_14544,N_12708);
xnor U16716 (N_16716,N_14393,N_12294);
or U16717 (N_16717,N_12987,N_13547);
nand U16718 (N_16718,N_12076,N_12512);
nor U16719 (N_16719,N_13068,N_14526);
nand U16720 (N_16720,N_13218,N_13954);
nand U16721 (N_16721,N_14986,N_12999);
nor U16722 (N_16722,N_12646,N_12395);
or U16723 (N_16723,N_12682,N_12172);
xor U16724 (N_16724,N_13027,N_13750);
or U16725 (N_16725,N_13602,N_12467);
nor U16726 (N_16726,N_12719,N_13921);
or U16727 (N_16727,N_13199,N_14610);
and U16728 (N_16728,N_12847,N_14198);
nor U16729 (N_16729,N_14731,N_13474);
and U16730 (N_16730,N_14047,N_12459);
or U16731 (N_16731,N_12022,N_14670);
nand U16732 (N_16732,N_13180,N_13853);
or U16733 (N_16733,N_12813,N_13320);
nor U16734 (N_16734,N_13113,N_12825);
nor U16735 (N_16735,N_13442,N_13674);
nand U16736 (N_16736,N_14956,N_14548);
or U16737 (N_16737,N_14076,N_12114);
nor U16738 (N_16738,N_13138,N_14674);
nand U16739 (N_16739,N_13376,N_12800);
nor U16740 (N_16740,N_12854,N_12726);
or U16741 (N_16741,N_13793,N_12377);
xnor U16742 (N_16742,N_12793,N_13706);
or U16743 (N_16743,N_13477,N_14628);
nand U16744 (N_16744,N_13275,N_13378);
nand U16745 (N_16745,N_13598,N_14742);
or U16746 (N_16746,N_12977,N_12630);
and U16747 (N_16747,N_14923,N_13177);
nor U16748 (N_16748,N_14945,N_12378);
nor U16749 (N_16749,N_12272,N_12371);
nor U16750 (N_16750,N_14501,N_14391);
nor U16751 (N_16751,N_14371,N_13893);
and U16752 (N_16752,N_13886,N_13624);
or U16753 (N_16753,N_13598,N_14094);
or U16754 (N_16754,N_13253,N_13917);
nand U16755 (N_16755,N_13047,N_14542);
or U16756 (N_16756,N_12627,N_14625);
nor U16757 (N_16757,N_12405,N_13733);
and U16758 (N_16758,N_12485,N_14763);
and U16759 (N_16759,N_12823,N_14811);
xnor U16760 (N_16760,N_14879,N_12346);
and U16761 (N_16761,N_14740,N_13345);
or U16762 (N_16762,N_13071,N_12473);
nand U16763 (N_16763,N_14674,N_13905);
or U16764 (N_16764,N_12765,N_14440);
nand U16765 (N_16765,N_12821,N_14500);
and U16766 (N_16766,N_13862,N_14445);
xnor U16767 (N_16767,N_13662,N_13139);
xor U16768 (N_16768,N_13975,N_14647);
and U16769 (N_16769,N_13387,N_14146);
and U16770 (N_16770,N_13434,N_14901);
nand U16771 (N_16771,N_14075,N_14386);
xnor U16772 (N_16772,N_12442,N_13636);
nor U16773 (N_16773,N_14645,N_12886);
nor U16774 (N_16774,N_14612,N_13350);
and U16775 (N_16775,N_14778,N_12841);
xnor U16776 (N_16776,N_14870,N_13739);
or U16777 (N_16777,N_13016,N_13206);
or U16778 (N_16778,N_12167,N_14669);
or U16779 (N_16779,N_14365,N_12491);
xor U16780 (N_16780,N_12160,N_14487);
nand U16781 (N_16781,N_14815,N_12657);
nand U16782 (N_16782,N_12321,N_12985);
xnor U16783 (N_16783,N_12160,N_13022);
or U16784 (N_16784,N_12737,N_13142);
xnor U16785 (N_16785,N_14215,N_12650);
xnor U16786 (N_16786,N_13687,N_14734);
nand U16787 (N_16787,N_13182,N_13052);
nand U16788 (N_16788,N_14524,N_13855);
and U16789 (N_16789,N_13746,N_12610);
or U16790 (N_16790,N_13140,N_12483);
and U16791 (N_16791,N_14156,N_12176);
or U16792 (N_16792,N_14884,N_12218);
nor U16793 (N_16793,N_13465,N_12909);
xnor U16794 (N_16794,N_14122,N_14518);
or U16795 (N_16795,N_12994,N_14285);
xor U16796 (N_16796,N_13918,N_12001);
nand U16797 (N_16797,N_13557,N_14566);
and U16798 (N_16798,N_14280,N_13278);
nor U16799 (N_16799,N_12524,N_14928);
and U16800 (N_16800,N_12734,N_13065);
nand U16801 (N_16801,N_12928,N_13098);
xor U16802 (N_16802,N_12078,N_14580);
and U16803 (N_16803,N_13746,N_12130);
xnor U16804 (N_16804,N_14061,N_13320);
or U16805 (N_16805,N_12962,N_14757);
nor U16806 (N_16806,N_14651,N_12394);
xor U16807 (N_16807,N_12511,N_13372);
and U16808 (N_16808,N_13451,N_12222);
or U16809 (N_16809,N_12666,N_12287);
nor U16810 (N_16810,N_12635,N_12214);
xor U16811 (N_16811,N_14147,N_13819);
nand U16812 (N_16812,N_12914,N_13519);
xor U16813 (N_16813,N_12171,N_13251);
xnor U16814 (N_16814,N_14635,N_12679);
or U16815 (N_16815,N_14036,N_13889);
and U16816 (N_16816,N_12240,N_13823);
or U16817 (N_16817,N_12615,N_12345);
nor U16818 (N_16818,N_13118,N_12818);
or U16819 (N_16819,N_12341,N_14013);
xor U16820 (N_16820,N_13454,N_13529);
nand U16821 (N_16821,N_12925,N_14648);
nand U16822 (N_16822,N_14231,N_13346);
or U16823 (N_16823,N_14629,N_14098);
nor U16824 (N_16824,N_13549,N_13098);
xor U16825 (N_16825,N_12499,N_13565);
nand U16826 (N_16826,N_14709,N_13225);
xnor U16827 (N_16827,N_13516,N_14365);
nand U16828 (N_16828,N_14218,N_13848);
nand U16829 (N_16829,N_14676,N_14141);
xor U16830 (N_16830,N_13533,N_12216);
nor U16831 (N_16831,N_14304,N_12335);
xor U16832 (N_16832,N_12427,N_12993);
nand U16833 (N_16833,N_12434,N_13675);
nand U16834 (N_16834,N_14794,N_13767);
nor U16835 (N_16835,N_13210,N_14051);
and U16836 (N_16836,N_12836,N_12911);
or U16837 (N_16837,N_13020,N_12854);
xnor U16838 (N_16838,N_13717,N_13786);
or U16839 (N_16839,N_13640,N_12599);
or U16840 (N_16840,N_13131,N_13361);
xnor U16841 (N_16841,N_13457,N_14185);
nand U16842 (N_16842,N_13452,N_14524);
nand U16843 (N_16843,N_14216,N_14609);
xor U16844 (N_16844,N_13009,N_14995);
and U16845 (N_16845,N_13135,N_12572);
xnor U16846 (N_16846,N_14369,N_14569);
nor U16847 (N_16847,N_13417,N_14474);
xor U16848 (N_16848,N_13093,N_13938);
xor U16849 (N_16849,N_12433,N_12778);
xor U16850 (N_16850,N_14084,N_14328);
and U16851 (N_16851,N_14710,N_14926);
nand U16852 (N_16852,N_14409,N_12148);
and U16853 (N_16853,N_14072,N_13566);
nand U16854 (N_16854,N_14055,N_13113);
and U16855 (N_16855,N_13707,N_12575);
or U16856 (N_16856,N_12373,N_12952);
nand U16857 (N_16857,N_12920,N_13359);
xnor U16858 (N_16858,N_14601,N_13732);
and U16859 (N_16859,N_13095,N_14537);
nand U16860 (N_16860,N_12924,N_13169);
and U16861 (N_16861,N_12627,N_13726);
xnor U16862 (N_16862,N_13469,N_14244);
nand U16863 (N_16863,N_14381,N_13679);
nand U16864 (N_16864,N_14026,N_12602);
xor U16865 (N_16865,N_12878,N_14680);
nand U16866 (N_16866,N_13693,N_12758);
or U16867 (N_16867,N_13386,N_14211);
and U16868 (N_16868,N_13656,N_14037);
xnor U16869 (N_16869,N_13990,N_14403);
xnor U16870 (N_16870,N_12132,N_13827);
nor U16871 (N_16871,N_12923,N_13121);
nand U16872 (N_16872,N_12837,N_13800);
nor U16873 (N_16873,N_14232,N_12180);
and U16874 (N_16874,N_13120,N_12593);
or U16875 (N_16875,N_12217,N_13698);
xor U16876 (N_16876,N_12183,N_12241);
xnor U16877 (N_16877,N_12461,N_14894);
or U16878 (N_16878,N_12157,N_14618);
nor U16879 (N_16879,N_13838,N_13278);
or U16880 (N_16880,N_14022,N_13816);
nand U16881 (N_16881,N_13526,N_12309);
nor U16882 (N_16882,N_12658,N_12987);
nand U16883 (N_16883,N_14223,N_13375);
xnor U16884 (N_16884,N_14439,N_14361);
nor U16885 (N_16885,N_13476,N_14864);
or U16886 (N_16886,N_13954,N_12662);
xor U16887 (N_16887,N_12081,N_14671);
xor U16888 (N_16888,N_14338,N_12328);
and U16889 (N_16889,N_13761,N_12477);
or U16890 (N_16890,N_14822,N_13740);
or U16891 (N_16891,N_13732,N_14757);
xor U16892 (N_16892,N_14963,N_14406);
nand U16893 (N_16893,N_14241,N_14079);
or U16894 (N_16894,N_14592,N_13151);
nand U16895 (N_16895,N_12621,N_14865);
or U16896 (N_16896,N_12592,N_12085);
or U16897 (N_16897,N_14259,N_14963);
and U16898 (N_16898,N_12329,N_14287);
nand U16899 (N_16899,N_13133,N_14442);
xor U16900 (N_16900,N_14269,N_12744);
nand U16901 (N_16901,N_13638,N_12534);
or U16902 (N_16902,N_12103,N_14177);
xnor U16903 (N_16903,N_12441,N_13108);
nor U16904 (N_16904,N_14284,N_12086);
xor U16905 (N_16905,N_14707,N_14894);
nand U16906 (N_16906,N_14718,N_12318);
xnor U16907 (N_16907,N_13033,N_12396);
and U16908 (N_16908,N_12199,N_13437);
and U16909 (N_16909,N_12610,N_13134);
nand U16910 (N_16910,N_14816,N_13546);
or U16911 (N_16911,N_13907,N_13334);
and U16912 (N_16912,N_14488,N_12535);
nor U16913 (N_16913,N_12069,N_12693);
xnor U16914 (N_16914,N_13440,N_14450);
and U16915 (N_16915,N_12668,N_14726);
nand U16916 (N_16916,N_14053,N_14355);
nand U16917 (N_16917,N_14642,N_13454);
xnor U16918 (N_16918,N_13615,N_14183);
or U16919 (N_16919,N_13146,N_14965);
nor U16920 (N_16920,N_12704,N_13731);
nor U16921 (N_16921,N_12195,N_12547);
nand U16922 (N_16922,N_14548,N_12989);
xnor U16923 (N_16923,N_12437,N_12512);
xor U16924 (N_16924,N_14399,N_12708);
or U16925 (N_16925,N_12910,N_14614);
nand U16926 (N_16926,N_13842,N_14051);
xor U16927 (N_16927,N_13732,N_12171);
and U16928 (N_16928,N_12406,N_12355);
nand U16929 (N_16929,N_12757,N_14928);
and U16930 (N_16930,N_14751,N_12645);
xor U16931 (N_16931,N_12921,N_12347);
xnor U16932 (N_16932,N_14849,N_13834);
nand U16933 (N_16933,N_13956,N_12011);
or U16934 (N_16934,N_13457,N_14970);
nand U16935 (N_16935,N_14402,N_12342);
xor U16936 (N_16936,N_13041,N_14754);
xnor U16937 (N_16937,N_12903,N_14022);
nand U16938 (N_16938,N_13489,N_14927);
nor U16939 (N_16939,N_13650,N_13280);
xnor U16940 (N_16940,N_14951,N_13771);
nor U16941 (N_16941,N_13716,N_12543);
and U16942 (N_16942,N_13231,N_12164);
xnor U16943 (N_16943,N_14929,N_14334);
xnor U16944 (N_16944,N_12958,N_13779);
nand U16945 (N_16945,N_13872,N_13311);
xnor U16946 (N_16946,N_14220,N_12021);
or U16947 (N_16947,N_13437,N_13301);
and U16948 (N_16948,N_12454,N_14662);
or U16949 (N_16949,N_13777,N_12653);
nand U16950 (N_16950,N_14236,N_14890);
nor U16951 (N_16951,N_12869,N_13733);
xor U16952 (N_16952,N_14955,N_14960);
xor U16953 (N_16953,N_14362,N_14088);
nand U16954 (N_16954,N_12615,N_14040);
nand U16955 (N_16955,N_13971,N_14003);
xnor U16956 (N_16956,N_12135,N_12616);
nand U16957 (N_16957,N_12753,N_13178);
or U16958 (N_16958,N_13496,N_12756);
xnor U16959 (N_16959,N_13399,N_14806);
or U16960 (N_16960,N_13414,N_12230);
nand U16961 (N_16961,N_14124,N_13660);
nor U16962 (N_16962,N_14086,N_14312);
xor U16963 (N_16963,N_14080,N_12175);
and U16964 (N_16964,N_14664,N_13147);
and U16965 (N_16965,N_13720,N_14805);
xor U16966 (N_16966,N_14993,N_13857);
nor U16967 (N_16967,N_14798,N_12971);
xor U16968 (N_16968,N_12537,N_13193);
xnor U16969 (N_16969,N_14876,N_13563);
nand U16970 (N_16970,N_13999,N_13310);
or U16971 (N_16971,N_14845,N_13046);
nand U16972 (N_16972,N_12223,N_14900);
xnor U16973 (N_16973,N_13919,N_13183);
and U16974 (N_16974,N_13548,N_14614);
xnor U16975 (N_16975,N_12999,N_14208);
and U16976 (N_16976,N_13853,N_12350);
nor U16977 (N_16977,N_12959,N_13669);
or U16978 (N_16978,N_14198,N_14242);
nand U16979 (N_16979,N_12573,N_14745);
xor U16980 (N_16980,N_13919,N_13548);
nand U16981 (N_16981,N_13014,N_14929);
xor U16982 (N_16982,N_13835,N_13196);
nor U16983 (N_16983,N_12022,N_14845);
nand U16984 (N_16984,N_12421,N_12214);
xnor U16985 (N_16985,N_12678,N_14946);
and U16986 (N_16986,N_12422,N_14867);
or U16987 (N_16987,N_13012,N_13709);
nor U16988 (N_16988,N_13125,N_14728);
nor U16989 (N_16989,N_12103,N_12497);
or U16990 (N_16990,N_12984,N_14691);
and U16991 (N_16991,N_13042,N_14798);
or U16992 (N_16992,N_13201,N_13232);
nand U16993 (N_16993,N_12139,N_14844);
nor U16994 (N_16994,N_13273,N_12004);
and U16995 (N_16995,N_13967,N_12684);
xor U16996 (N_16996,N_13579,N_13260);
xnor U16997 (N_16997,N_12984,N_14260);
or U16998 (N_16998,N_12531,N_14348);
nor U16999 (N_16999,N_13479,N_13179);
nor U17000 (N_17000,N_12745,N_12080);
nand U17001 (N_17001,N_14835,N_12327);
nor U17002 (N_17002,N_13348,N_12213);
and U17003 (N_17003,N_12580,N_14481);
nand U17004 (N_17004,N_14009,N_12167);
or U17005 (N_17005,N_12216,N_12090);
xnor U17006 (N_17006,N_13563,N_14535);
xor U17007 (N_17007,N_13328,N_14667);
xnor U17008 (N_17008,N_12480,N_14389);
and U17009 (N_17009,N_13072,N_12909);
or U17010 (N_17010,N_12288,N_12019);
xnor U17011 (N_17011,N_13890,N_13910);
nand U17012 (N_17012,N_12948,N_14088);
and U17013 (N_17013,N_12358,N_13345);
xnor U17014 (N_17014,N_13039,N_12398);
xor U17015 (N_17015,N_12558,N_12018);
and U17016 (N_17016,N_12896,N_13533);
and U17017 (N_17017,N_13212,N_12935);
nor U17018 (N_17018,N_13505,N_12425);
nor U17019 (N_17019,N_14719,N_14829);
nand U17020 (N_17020,N_14932,N_12891);
or U17021 (N_17021,N_13510,N_12215);
or U17022 (N_17022,N_13321,N_13493);
xor U17023 (N_17023,N_12626,N_13997);
nand U17024 (N_17024,N_13459,N_12931);
nor U17025 (N_17025,N_13778,N_13602);
xor U17026 (N_17026,N_12075,N_14448);
nand U17027 (N_17027,N_12779,N_14658);
xor U17028 (N_17028,N_14298,N_13375);
nand U17029 (N_17029,N_13832,N_13796);
and U17030 (N_17030,N_13667,N_13003);
nand U17031 (N_17031,N_14911,N_12480);
nand U17032 (N_17032,N_12325,N_14396);
nand U17033 (N_17033,N_13809,N_12992);
or U17034 (N_17034,N_14954,N_12569);
and U17035 (N_17035,N_12140,N_14628);
or U17036 (N_17036,N_14290,N_14520);
and U17037 (N_17037,N_14645,N_14180);
nand U17038 (N_17038,N_13378,N_14295);
nor U17039 (N_17039,N_14704,N_13567);
xnor U17040 (N_17040,N_14405,N_14490);
or U17041 (N_17041,N_13121,N_14575);
and U17042 (N_17042,N_14149,N_14304);
or U17043 (N_17043,N_12785,N_12079);
or U17044 (N_17044,N_14495,N_14863);
or U17045 (N_17045,N_13282,N_13633);
and U17046 (N_17046,N_13934,N_12184);
and U17047 (N_17047,N_13525,N_12450);
nor U17048 (N_17048,N_12417,N_14533);
and U17049 (N_17049,N_12895,N_14241);
or U17050 (N_17050,N_14083,N_13010);
or U17051 (N_17051,N_13641,N_12925);
nand U17052 (N_17052,N_12353,N_13731);
nor U17053 (N_17053,N_12413,N_14714);
xnor U17054 (N_17054,N_14047,N_14236);
and U17055 (N_17055,N_14923,N_13809);
and U17056 (N_17056,N_12832,N_12774);
nor U17057 (N_17057,N_14589,N_13228);
nor U17058 (N_17058,N_14415,N_12105);
nand U17059 (N_17059,N_14500,N_14582);
nor U17060 (N_17060,N_14275,N_12294);
or U17061 (N_17061,N_12199,N_12834);
or U17062 (N_17062,N_14171,N_14149);
or U17063 (N_17063,N_13916,N_14960);
or U17064 (N_17064,N_13984,N_14221);
or U17065 (N_17065,N_13869,N_12418);
or U17066 (N_17066,N_12838,N_12483);
nor U17067 (N_17067,N_12657,N_12989);
or U17068 (N_17068,N_12643,N_13113);
xor U17069 (N_17069,N_12489,N_12793);
and U17070 (N_17070,N_12016,N_14468);
nand U17071 (N_17071,N_13836,N_14391);
nand U17072 (N_17072,N_13435,N_14426);
or U17073 (N_17073,N_14900,N_14813);
and U17074 (N_17074,N_12273,N_13369);
nor U17075 (N_17075,N_13949,N_13301);
nor U17076 (N_17076,N_14889,N_14838);
nor U17077 (N_17077,N_13056,N_13294);
nor U17078 (N_17078,N_13381,N_13593);
nor U17079 (N_17079,N_13042,N_14359);
and U17080 (N_17080,N_13132,N_13450);
nand U17081 (N_17081,N_13047,N_12204);
xor U17082 (N_17082,N_12356,N_14677);
nand U17083 (N_17083,N_13453,N_12157);
and U17084 (N_17084,N_12871,N_12249);
nand U17085 (N_17085,N_12527,N_14352);
xor U17086 (N_17086,N_14597,N_13155);
and U17087 (N_17087,N_12710,N_12787);
nor U17088 (N_17088,N_12978,N_12504);
and U17089 (N_17089,N_12233,N_13454);
or U17090 (N_17090,N_12722,N_12791);
xor U17091 (N_17091,N_13608,N_13784);
or U17092 (N_17092,N_12733,N_13105);
nor U17093 (N_17093,N_12993,N_14912);
or U17094 (N_17094,N_14338,N_12491);
nand U17095 (N_17095,N_12147,N_12734);
nand U17096 (N_17096,N_13484,N_13597);
nor U17097 (N_17097,N_13413,N_12907);
xor U17098 (N_17098,N_12394,N_13112);
xor U17099 (N_17099,N_13540,N_12123);
xor U17100 (N_17100,N_14317,N_12107);
or U17101 (N_17101,N_14868,N_13890);
nor U17102 (N_17102,N_12885,N_12961);
nand U17103 (N_17103,N_13200,N_12530);
and U17104 (N_17104,N_12643,N_12162);
and U17105 (N_17105,N_13238,N_14706);
nand U17106 (N_17106,N_14545,N_12336);
and U17107 (N_17107,N_13720,N_12311);
and U17108 (N_17108,N_14278,N_13654);
xor U17109 (N_17109,N_12776,N_12125);
xor U17110 (N_17110,N_12227,N_13536);
and U17111 (N_17111,N_13747,N_14474);
or U17112 (N_17112,N_12461,N_12569);
nand U17113 (N_17113,N_14121,N_14160);
or U17114 (N_17114,N_14664,N_13311);
nor U17115 (N_17115,N_14017,N_12546);
nand U17116 (N_17116,N_12622,N_12709);
xnor U17117 (N_17117,N_12119,N_13899);
and U17118 (N_17118,N_14104,N_13666);
nand U17119 (N_17119,N_13261,N_12174);
nand U17120 (N_17120,N_12910,N_12772);
or U17121 (N_17121,N_14245,N_14621);
nor U17122 (N_17122,N_14087,N_14679);
xnor U17123 (N_17123,N_14693,N_13134);
xnor U17124 (N_17124,N_14501,N_13945);
or U17125 (N_17125,N_12639,N_13436);
and U17126 (N_17126,N_13488,N_14967);
or U17127 (N_17127,N_13617,N_13362);
nor U17128 (N_17128,N_13496,N_13791);
and U17129 (N_17129,N_14553,N_14333);
or U17130 (N_17130,N_14780,N_14177);
nor U17131 (N_17131,N_14461,N_12736);
nor U17132 (N_17132,N_12766,N_12089);
xor U17133 (N_17133,N_13497,N_13522);
nand U17134 (N_17134,N_14155,N_14578);
nor U17135 (N_17135,N_13592,N_14685);
xor U17136 (N_17136,N_13764,N_14252);
xnor U17137 (N_17137,N_12830,N_13471);
nor U17138 (N_17138,N_13437,N_12750);
or U17139 (N_17139,N_14294,N_14331);
nor U17140 (N_17140,N_12269,N_12377);
nor U17141 (N_17141,N_12558,N_12478);
xor U17142 (N_17142,N_13671,N_12765);
and U17143 (N_17143,N_14425,N_13364);
and U17144 (N_17144,N_14973,N_12841);
nand U17145 (N_17145,N_14916,N_12499);
xor U17146 (N_17146,N_12894,N_12325);
and U17147 (N_17147,N_14203,N_14799);
nor U17148 (N_17148,N_12632,N_13167);
or U17149 (N_17149,N_14818,N_14059);
nand U17150 (N_17150,N_13887,N_12216);
and U17151 (N_17151,N_14506,N_14335);
or U17152 (N_17152,N_12029,N_13780);
or U17153 (N_17153,N_14338,N_12352);
or U17154 (N_17154,N_12230,N_13079);
xnor U17155 (N_17155,N_14289,N_12093);
xor U17156 (N_17156,N_13857,N_13654);
xnor U17157 (N_17157,N_13130,N_12042);
nand U17158 (N_17158,N_13880,N_13856);
or U17159 (N_17159,N_12372,N_12902);
or U17160 (N_17160,N_12751,N_13666);
nor U17161 (N_17161,N_14903,N_14249);
nor U17162 (N_17162,N_13278,N_12006);
xor U17163 (N_17163,N_14743,N_13855);
and U17164 (N_17164,N_14238,N_13371);
xor U17165 (N_17165,N_13695,N_13839);
and U17166 (N_17166,N_13294,N_12993);
or U17167 (N_17167,N_14134,N_13615);
nor U17168 (N_17168,N_14352,N_12017);
xnor U17169 (N_17169,N_14372,N_13955);
nand U17170 (N_17170,N_12496,N_14949);
or U17171 (N_17171,N_12728,N_13163);
xnor U17172 (N_17172,N_12020,N_13861);
or U17173 (N_17173,N_13710,N_14944);
nand U17174 (N_17174,N_14137,N_12124);
or U17175 (N_17175,N_12273,N_13849);
or U17176 (N_17176,N_14953,N_13042);
xnor U17177 (N_17177,N_12486,N_13500);
nand U17178 (N_17178,N_13833,N_14960);
xor U17179 (N_17179,N_13127,N_12574);
nor U17180 (N_17180,N_14206,N_12589);
or U17181 (N_17181,N_13881,N_12972);
or U17182 (N_17182,N_13251,N_14105);
xnor U17183 (N_17183,N_12320,N_14209);
xnor U17184 (N_17184,N_14774,N_14002);
xor U17185 (N_17185,N_13129,N_13733);
xor U17186 (N_17186,N_13317,N_12253);
nor U17187 (N_17187,N_14425,N_14137);
and U17188 (N_17188,N_14666,N_13899);
nor U17189 (N_17189,N_13189,N_12058);
or U17190 (N_17190,N_13134,N_12060);
nand U17191 (N_17191,N_14722,N_13734);
nand U17192 (N_17192,N_12307,N_14463);
xor U17193 (N_17193,N_12834,N_14389);
nor U17194 (N_17194,N_14144,N_13486);
nor U17195 (N_17195,N_14600,N_14663);
nand U17196 (N_17196,N_13180,N_14253);
nand U17197 (N_17197,N_13678,N_14793);
and U17198 (N_17198,N_14973,N_13857);
nor U17199 (N_17199,N_14384,N_12008);
nand U17200 (N_17200,N_12974,N_13805);
nor U17201 (N_17201,N_14307,N_14350);
and U17202 (N_17202,N_14145,N_14877);
xor U17203 (N_17203,N_13691,N_13888);
or U17204 (N_17204,N_12371,N_14594);
and U17205 (N_17205,N_13965,N_13203);
xnor U17206 (N_17206,N_14338,N_13366);
or U17207 (N_17207,N_13890,N_12443);
nand U17208 (N_17208,N_12116,N_14090);
or U17209 (N_17209,N_13193,N_12280);
xnor U17210 (N_17210,N_13876,N_14465);
and U17211 (N_17211,N_14657,N_14672);
nor U17212 (N_17212,N_14336,N_12402);
xnor U17213 (N_17213,N_13677,N_14503);
and U17214 (N_17214,N_12559,N_12447);
xnor U17215 (N_17215,N_12538,N_13849);
xnor U17216 (N_17216,N_12858,N_14033);
nor U17217 (N_17217,N_13719,N_13458);
nor U17218 (N_17218,N_13070,N_14934);
nor U17219 (N_17219,N_14646,N_12430);
nand U17220 (N_17220,N_13432,N_12113);
xor U17221 (N_17221,N_13017,N_14492);
nor U17222 (N_17222,N_13347,N_12153);
or U17223 (N_17223,N_14151,N_14126);
nand U17224 (N_17224,N_14379,N_13078);
and U17225 (N_17225,N_14040,N_12303);
nand U17226 (N_17226,N_13973,N_12548);
or U17227 (N_17227,N_14350,N_12506);
nor U17228 (N_17228,N_14894,N_14437);
xnor U17229 (N_17229,N_14560,N_13656);
nor U17230 (N_17230,N_13248,N_13500);
and U17231 (N_17231,N_14555,N_12625);
and U17232 (N_17232,N_13538,N_12025);
nand U17233 (N_17233,N_13329,N_12777);
nand U17234 (N_17234,N_13335,N_14783);
nor U17235 (N_17235,N_12721,N_12759);
or U17236 (N_17236,N_14512,N_14558);
or U17237 (N_17237,N_12597,N_13372);
or U17238 (N_17238,N_14187,N_13708);
nand U17239 (N_17239,N_13014,N_13549);
xor U17240 (N_17240,N_13099,N_14420);
and U17241 (N_17241,N_12295,N_14536);
nand U17242 (N_17242,N_13194,N_14846);
nand U17243 (N_17243,N_12645,N_14975);
nand U17244 (N_17244,N_13175,N_13220);
and U17245 (N_17245,N_13571,N_13888);
nor U17246 (N_17246,N_12607,N_14153);
or U17247 (N_17247,N_13383,N_13760);
or U17248 (N_17248,N_13332,N_13481);
nor U17249 (N_17249,N_13938,N_13560);
or U17250 (N_17250,N_12155,N_13798);
xnor U17251 (N_17251,N_14477,N_14465);
nand U17252 (N_17252,N_14387,N_14892);
xnor U17253 (N_17253,N_13611,N_14665);
and U17254 (N_17254,N_13548,N_14866);
xnor U17255 (N_17255,N_14350,N_13399);
and U17256 (N_17256,N_13978,N_13184);
nor U17257 (N_17257,N_14734,N_13190);
or U17258 (N_17258,N_14657,N_13404);
or U17259 (N_17259,N_14945,N_12468);
nor U17260 (N_17260,N_12972,N_13339);
nand U17261 (N_17261,N_14130,N_13185);
nand U17262 (N_17262,N_13561,N_12743);
or U17263 (N_17263,N_12007,N_14240);
or U17264 (N_17264,N_13155,N_12927);
or U17265 (N_17265,N_13375,N_14620);
and U17266 (N_17266,N_13748,N_13646);
xor U17267 (N_17267,N_13101,N_12081);
nor U17268 (N_17268,N_12621,N_14204);
or U17269 (N_17269,N_13447,N_13258);
nand U17270 (N_17270,N_12033,N_14312);
xor U17271 (N_17271,N_12003,N_13459);
and U17272 (N_17272,N_14696,N_13819);
nor U17273 (N_17273,N_13493,N_13573);
nor U17274 (N_17274,N_12516,N_12007);
nand U17275 (N_17275,N_14248,N_12595);
nand U17276 (N_17276,N_14060,N_14745);
nor U17277 (N_17277,N_14580,N_13237);
nand U17278 (N_17278,N_12506,N_12798);
and U17279 (N_17279,N_14454,N_13420);
nor U17280 (N_17280,N_14881,N_14221);
or U17281 (N_17281,N_13060,N_12014);
nand U17282 (N_17282,N_14059,N_14291);
xnor U17283 (N_17283,N_13742,N_14437);
and U17284 (N_17284,N_12426,N_13739);
xor U17285 (N_17285,N_12854,N_14898);
nor U17286 (N_17286,N_14583,N_14660);
nor U17287 (N_17287,N_14450,N_14901);
or U17288 (N_17288,N_13474,N_12742);
and U17289 (N_17289,N_14889,N_12447);
nand U17290 (N_17290,N_14761,N_13219);
nor U17291 (N_17291,N_13595,N_13352);
nor U17292 (N_17292,N_14588,N_12412);
nor U17293 (N_17293,N_13997,N_13427);
nand U17294 (N_17294,N_14668,N_13504);
xnor U17295 (N_17295,N_13232,N_12823);
and U17296 (N_17296,N_12736,N_12193);
xor U17297 (N_17297,N_14730,N_13669);
and U17298 (N_17298,N_12590,N_13918);
nand U17299 (N_17299,N_13330,N_13000);
and U17300 (N_17300,N_14281,N_14981);
and U17301 (N_17301,N_12086,N_14697);
or U17302 (N_17302,N_14338,N_12825);
nor U17303 (N_17303,N_13067,N_13189);
nor U17304 (N_17304,N_13507,N_14574);
nand U17305 (N_17305,N_12028,N_14614);
and U17306 (N_17306,N_14455,N_12016);
or U17307 (N_17307,N_12246,N_13111);
or U17308 (N_17308,N_14833,N_13064);
xor U17309 (N_17309,N_13260,N_14733);
nor U17310 (N_17310,N_14197,N_14107);
and U17311 (N_17311,N_12365,N_12570);
and U17312 (N_17312,N_14023,N_14103);
xnor U17313 (N_17313,N_13891,N_12954);
and U17314 (N_17314,N_14115,N_14374);
nor U17315 (N_17315,N_13788,N_13614);
nand U17316 (N_17316,N_14928,N_13367);
nand U17317 (N_17317,N_13817,N_14115);
xnor U17318 (N_17318,N_14515,N_13205);
nand U17319 (N_17319,N_12013,N_14002);
xnor U17320 (N_17320,N_14410,N_12664);
nand U17321 (N_17321,N_12427,N_13958);
nor U17322 (N_17322,N_14995,N_13754);
nand U17323 (N_17323,N_12889,N_12569);
or U17324 (N_17324,N_14217,N_12214);
and U17325 (N_17325,N_13154,N_12867);
or U17326 (N_17326,N_12353,N_12383);
nor U17327 (N_17327,N_13354,N_12537);
nand U17328 (N_17328,N_13037,N_13826);
or U17329 (N_17329,N_12005,N_12868);
and U17330 (N_17330,N_14991,N_14701);
nand U17331 (N_17331,N_12965,N_12757);
xor U17332 (N_17332,N_13570,N_13849);
nand U17333 (N_17333,N_13434,N_12228);
and U17334 (N_17334,N_14688,N_13969);
or U17335 (N_17335,N_13596,N_14647);
nor U17336 (N_17336,N_14893,N_14938);
xor U17337 (N_17337,N_13352,N_14430);
nand U17338 (N_17338,N_12424,N_13922);
nor U17339 (N_17339,N_13346,N_12802);
or U17340 (N_17340,N_14318,N_14003);
nand U17341 (N_17341,N_13204,N_14384);
nor U17342 (N_17342,N_14015,N_12430);
nor U17343 (N_17343,N_14045,N_12750);
xnor U17344 (N_17344,N_13827,N_12143);
and U17345 (N_17345,N_13140,N_13244);
nand U17346 (N_17346,N_14414,N_13316);
nand U17347 (N_17347,N_13753,N_12085);
xor U17348 (N_17348,N_14003,N_13033);
and U17349 (N_17349,N_13472,N_13796);
or U17350 (N_17350,N_14116,N_13445);
nor U17351 (N_17351,N_13085,N_13681);
xor U17352 (N_17352,N_13773,N_13462);
nand U17353 (N_17353,N_13032,N_14081);
or U17354 (N_17354,N_13673,N_13843);
or U17355 (N_17355,N_12673,N_14659);
or U17356 (N_17356,N_12820,N_13939);
nand U17357 (N_17357,N_14085,N_12749);
xor U17358 (N_17358,N_14716,N_13629);
nand U17359 (N_17359,N_13161,N_14353);
nand U17360 (N_17360,N_12827,N_13681);
xor U17361 (N_17361,N_12366,N_13140);
xnor U17362 (N_17362,N_13064,N_12991);
xnor U17363 (N_17363,N_12193,N_13314);
or U17364 (N_17364,N_12015,N_13550);
xor U17365 (N_17365,N_13094,N_13658);
and U17366 (N_17366,N_13761,N_12828);
and U17367 (N_17367,N_12017,N_12079);
nor U17368 (N_17368,N_13871,N_12973);
and U17369 (N_17369,N_12180,N_12387);
nor U17370 (N_17370,N_13422,N_12166);
xor U17371 (N_17371,N_12163,N_14436);
nand U17372 (N_17372,N_12501,N_14253);
nand U17373 (N_17373,N_13427,N_13670);
or U17374 (N_17374,N_13302,N_13709);
xnor U17375 (N_17375,N_12201,N_12708);
or U17376 (N_17376,N_12344,N_14362);
and U17377 (N_17377,N_14504,N_14292);
and U17378 (N_17378,N_13212,N_14864);
xor U17379 (N_17379,N_13402,N_14347);
and U17380 (N_17380,N_12948,N_14214);
nor U17381 (N_17381,N_12232,N_13230);
or U17382 (N_17382,N_12929,N_12580);
nand U17383 (N_17383,N_12820,N_13953);
nor U17384 (N_17384,N_12582,N_14824);
or U17385 (N_17385,N_14503,N_13250);
nor U17386 (N_17386,N_14878,N_13952);
xnor U17387 (N_17387,N_14291,N_12962);
xnor U17388 (N_17388,N_14456,N_14873);
and U17389 (N_17389,N_12246,N_14836);
and U17390 (N_17390,N_14784,N_12427);
nor U17391 (N_17391,N_13197,N_12197);
nor U17392 (N_17392,N_14677,N_13491);
xnor U17393 (N_17393,N_13917,N_12631);
nor U17394 (N_17394,N_13369,N_13953);
or U17395 (N_17395,N_14188,N_14836);
nand U17396 (N_17396,N_14866,N_14850);
or U17397 (N_17397,N_13374,N_14247);
nor U17398 (N_17398,N_14130,N_13328);
and U17399 (N_17399,N_13396,N_14385);
nor U17400 (N_17400,N_12752,N_13311);
or U17401 (N_17401,N_12263,N_14121);
nor U17402 (N_17402,N_12352,N_13698);
xnor U17403 (N_17403,N_14005,N_12409);
nor U17404 (N_17404,N_14203,N_14766);
nor U17405 (N_17405,N_13775,N_12648);
nor U17406 (N_17406,N_13242,N_12604);
nor U17407 (N_17407,N_14087,N_12559);
or U17408 (N_17408,N_13244,N_14796);
nor U17409 (N_17409,N_12844,N_14584);
nor U17410 (N_17410,N_12726,N_12012);
nor U17411 (N_17411,N_12026,N_12336);
xor U17412 (N_17412,N_14741,N_12922);
nor U17413 (N_17413,N_12972,N_14560);
nor U17414 (N_17414,N_12595,N_14317);
or U17415 (N_17415,N_13909,N_12585);
or U17416 (N_17416,N_13589,N_13908);
nor U17417 (N_17417,N_13453,N_13898);
or U17418 (N_17418,N_13746,N_13681);
nand U17419 (N_17419,N_14107,N_12542);
xnor U17420 (N_17420,N_12814,N_13881);
or U17421 (N_17421,N_12019,N_14691);
and U17422 (N_17422,N_13641,N_14784);
nand U17423 (N_17423,N_12327,N_12609);
and U17424 (N_17424,N_14209,N_14099);
nand U17425 (N_17425,N_14711,N_13367);
nand U17426 (N_17426,N_14024,N_13500);
xor U17427 (N_17427,N_13715,N_13289);
and U17428 (N_17428,N_14837,N_12148);
or U17429 (N_17429,N_13272,N_14159);
nor U17430 (N_17430,N_13096,N_13480);
or U17431 (N_17431,N_14185,N_12983);
xor U17432 (N_17432,N_14271,N_13737);
and U17433 (N_17433,N_13172,N_12626);
or U17434 (N_17434,N_13848,N_12307);
nor U17435 (N_17435,N_12008,N_12337);
nor U17436 (N_17436,N_14338,N_14285);
or U17437 (N_17437,N_14183,N_13075);
or U17438 (N_17438,N_14319,N_13224);
xnor U17439 (N_17439,N_13397,N_13726);
xnor U17440 (N_17440,N_13169,N_12268);
or U17441 (N_17441,N_12748,N_13056);
or U17442 (N_17442,N_14504,N_12677);
and U17443 (N_17443,N_14569,N_12918);
or U17444 (N_17444,N_14498,N_12006);
nand U17445 (N_17445,N_12637,N_14541);
xor U17446 (N_17446,N_14312,N_14503);
xnor U17447 (N_17447,N_13746,N_13991);
and U17448 (N_17448,N_13020,N_12383);
or U17449 (N_17449,N_12616,N_13200);
xor U17450 (N_17450,N_12202,N_14695);
xnor U17451 (N_17451,N_13266,N_12146);
or U17452 (N_17452,N_13334,N_14323);
xnor U17453 (N_17453,N_12391,N_14109);
or U17454 (N_17454,N_13777,N_14861);
nor U17455 (N_17455,N_13009,N_12893);
xnor U17456 (N_17456,N_13604,N_12302);
or U17457 (N_17457,N_13548,N_12847);
and U17458 (N_17458,N_13545,N_13276);
nand U17459 (N_17459,N_14343,N_13586);
nand U17460 (N_17460,N_14941,N_14549);
nor U17461 (N_17461,N_12277,N_13967);
xnor U17462 (N_17462,N_13618,N_14576);
and U17463 (N_17463,N_13538,N_12488);
xor U17464 (N_17464,N_14355,N_13615);
xor U17465 (N_17465,N_13122,N_12328);
xnor U17466 (N_17466,N_13971,N_13927);
nor U17467 (N_17467,N_12832,N_13726);
and U17468 (N_17468,N_13837,N_14049);
nor U17469 (N_17469,N_14550,N_14095);
xor U17470 (N_17470,N_12619,N_12368);
and U17471 (N_17471,N_14847,N_13031);
xor U17472 (N_17472,N_12956,N_14205);
nor U17473 (N_17473,N_13262,N_12250);
or U17474 (N_17474,N_14245,N_12935);
xnor U17475 (N_17475,N_12115,N_14303);
or U17476 (N_17476,N_12832,N_12926);
xnor U17477 (N_17477,N_14756,N_14113);
xnor U17478 (N_17478,N_12758,N_14562);
and U17479 (N_17479,N_14516,N_14284);
xor U17480 (N_17480,N_12161,N_13272);
or U17481 (N_17481,N_14286,N_13890);
or U17482 (N_17482,N_12261,N_14960);
or U17483 (N_17483,N_12656,N_12851);
nor U17484 (N_17484,N_14194,N_12346);
nand U17485 (N_17485,N_13614,N_12342);
nand U17486 (N_17486,N_14693,N_13771);
or U17487 (N_17487,N_13607,N_13808);
nor U17488 (N_17488,N_14363,N_14681);
xnor U17489 (N_17489,N_13308,N_13248);
nand U17490 (N_17490,N_13360,N_13464);
xor U17491 (N_17491,N_14626,N_13706);
xor U17492 (N_17492,N_13088,N_12454);
xor U17493 (N_17493,N_13154,N_13844);
or U17494 (N_17494,N_13612,N_14252);
or U17495 (N_17495,N_14805,N_14299);
nor U17496 (N_17496,N_13001,N_13534);
nor U17497 (N_17497,N_14603,N_14184);
or U17498 (N_17498,N_14329,N_12148);
or U17499 (N_17499,N_13369,N_13419);
or U17500 (N_17500,N_12937,N_12034);
nand U17501 (N_17501,N_13720,N_13294);
or U17502 (N_17502,N_13348,N_13525);
or U17503 (N_17503,N_14363,N_13386);
nor U17504 (N_17504,N_13355,N_13925);
or U17505 (N_17505,N_12940,N_12720);
or U17506 (N_17506,N_12136,N_14077);
nor U17507 (N_17507,N_13889,N_14294);
xor U17508 (N_17508,N_13221,N_13778);
or U17509 (N_17509,N_13324,N_14386);
and U17510 (N_17510,N_14100,N_12421);
xnor U17511 (N_17511,N_12583,N_12603);
nand U17512 (N_17512,N_14350,N_13764);
or U17513 (N_17513,N_12473,N_12555);
nand U17514 (N_17514,N_14122,N_12111);
nand U17515 (N_17515,N_12471,N_13945);
xor U17516 (N_17516,N_13859,N_13216);
nand U17517 (N_17517,N_12182,N_13148);
and U17518 (N_17518,N_12654,N_13595);
and U17519 (N_17519,N_14472,N_13881);
nor U17520 (N_17520,N_12496,N_12041);
and U17521 (N_17521,N_13552,N_14345);
nand U17522 (N_17522,N_13999,N_14683);
and U17523 (N_17523,N_14146,N_12031);
and U17524 (N_17524,N_12046,N_13364);
and U17525 (N_17525,N_12461,N_13003);
or U17526 (N_17526,N_14818,N_14448);
nand U17527 (N_17527,N_13425,N_12157);
nand U17528 (N_17528,N_14116,N_12818);
xnor U17529 (N_17529,N_13774,N_12295);
and U17530 (N_17530,N_14790,N_13594);
nor U17531 (N_17531,N_13427,N_12905);
or U17532 (N_17532,N_12844,N_13107);
and U17533 (N_17533,N_12150,N_14102);
nand U17534 (N_17534,N_12013,N_12656);
nand U17535 (N_17535,N_13368,N_14651);
xnor U17536 (N_17536,N_12735,N_13974);
xor U17537 (N_17537,N_13785,N_14348);
nand U17538 (N_17538,N_14565,N_12937);
xor U17539 (N_17539,N_14045,N_12792);
nor U17540 (N_17540,N_13194,N_13390);
nor U17541 (N_17541,N_12296,N_12466);
or U17542 (N_17542,N_14325,N_12181);
and U17543 (N_17543,N_14595,N_13321);
nand U17544 (N_17544,N_12726,N_13274);
or U17545 (N_17545,N_13216,N_12219);
nor U17546 (N_17546,N_14157,N_12269);
or U17547 (N_17547,N_13185,N_14562);
nor U17548 (N_17548,N_13776,N_12552);
nor U17549 (N_17549,N_12053,N_12088);
and U17550 (N_17550,N_13558,N_12795);
nor U17551 (N_17551,N_13035,N_13667);
nor U17552 (N_17552,N_14511,N_14869);
and U17553 (N_17553,N_12385,N_14426);
and U17554 (N_17554,N_12474,N_13890);
xnor U17555 (N_17555,N_14236,N_13716);
and U17556 (N_17556,N_14888,N_13294);
xor U17557 (N_17557,N_14618,N_14514);
xor U17558 (N_17558,N_14556,N_12445);
nor U17559 (N_17559,N_14479,N_13685);
nand U17560 (N_17560,N_13224,N_13434);
nor U17561 (N_17561,N_12109,N_12374);
nand U17562 (N_17562,N_14017,N_14593);
nor U17563 (N_17563,N_13818,N_14672);
and U17564 (N_17564,N_12588,N_12906);
nand U17565 (N_17565,N_12419,N_14903);
nor U17566 (N_17566,N_13520,N_12633);
nand U17567 (N_17567,N_13279,N_14777);
nor U17568 (N_17568,N_14022,N_12042);
nand U17569 (N_17569,N_12764,N_13707);
nand U17570 (N_17570,N_14046,N_13009);
xor U17571 (N_17571,N_13730,N_12061);
xor U17572 (N_17572,N_13495,N_12075);
or U17573 (N_17573,N_13537,N_12225);
or U17574 (N_17574,N_14746,N_12013);
xor U17575 (N_17575,N_12419,N_13793);
xnor U17576 (N_17576,N_13245,N_12604);
and U17577 (N_17577,N_13837,N_14550);
or U17578 (N_17578,N_13601,N_12792);
nand U17579 (N_17579,N_12024,N_12394);
nand U17580 (N_17580,N_14367,N_14891);
nand U17581 (N_17581,N_13647,N_13526);
nand U17582 (N_17582,N_12342,N_13213);
xor U17583 (N_17583,N_12254,N_13273);
nor U17584 (N_17584,N_12160,N_14902);
and U17585 (N_17585,N_14574,N_12288);
nand U17586 (N_17586,N_13121,N_13187);
and U17587 (N_17587,N_12714,N_12594);
nand U17588 (N_17588,N_13719,N_13859);
nand U17589 (N_17589,N_12911,N_13528);
xor U17590 (N_17590,N_14107,N_14693);
xnor U17591 (N_17591,N_13376,N_13248);
or U17592 (N_17592,N_14732,N_13440);
nand U17593 (N_17593,N_14889,N_12187);
or U17594 (N_17594,N_13860,N_13937);
or U17595 (N_17595,N_12392,N_12276);
and U17596 (N_17596,N_13703,N_12395);
or U17597 (N_17597,N_14696,N_14959);
xnor U17598 (N_17598,N_14452,N_13937);
nor U17599 (N_17599,N_14178,N_14796);
and U17600 (N_17600,N_12510,N_14931);
nand U17601 (N_17601,N_14011,N_12177);
or U17602 (N_17602,N_13006,N_14312);
nor U17603 (N_17603,N_13473,N_13991);
nor U17604 (N_17604,N_14461,N_14647);
or U17605 (N_17605,N_12011,N_13934);
and U17606 (N_17606,N_14036,N_12433);
xor U17607 (N_17607,N_14898,N_13213);
and U17608 (N_17608,N_13174,N_14150);
xnor U17609 (N_17609,N_13018,N_12019);
and U17610 (N_17610,N_12785,N_12892);
nand U17611 (N_17611,N_14517,N_13412);
and U17612 (N_17612,N_12447,N_14156);
xnor U17613 (N_17613,N_13532,N_12115);
and U17614 (N_17614,N_13767,N_13780);
and U17615 (N_17615,N_14331,N_14995);
and U17616 (N_17616,N_13577,N_14016);
and U17617 (N_17617,N_14605,N_12550);
or U17618 (N_17618,N_14613,N_14462);
and U17619 (N_17619,N_14989,N_13756);
and U17620 (N_17620,N_12330,N_12548);
xnor U17621 (N_17621,N_14370,N_12179);
xor U17622 (N_17622,N_12306,N_14850);
nand U17623 (N_17623,N_13384,N_13827);
nand U17624 (N_17624,N_13049,N_13748);
or U17625 (N_17625,N_12772,N_13346);
or U17626 (N_17626,N_14217,N_14317);
xor U17627 (N_17627,N_14769,N_13393);
nor U17628 (N_17628,N_13888,N_14238);
nand U17629 (N_17629,N_14129,N_13038);
nor U17630 (N_17630,N_13019,N_13989);
or U17631 (N_17631,N_14532,N_13035);
and U17632 (N_17632,N_12598,N_12008);
nor U17633 (N_17633,N_14281,N_12161);
nor U17634 (N_17634,N_14387,N_12836);
or U17635 (N_17635,N_12942,N_14954);
xor U17636 (N_17636,N_14041,N_14082);
nand U17637 (N_17637,N_12900,N_12205);
and U17638 (N_17638,N_12691,N_14443);
or U17639 (N_17639,N_14186,N_13756);
and U17640 (N_17640,N_14109,N_14993);
xnor U17641 (N_17641,N_12863,N_13788);
nand U17642 (N_17642,N_12586,N_12109);
and U17643 (N_17643,N_13255,N_14683);
or U17644 (N_17644,N_12023,N_13993);
and U17645 (N_17645,N_14154,N_14585);
xor U17646 (N_17646,N_13907,N_13260);
or U17647 (N_17647,N_14193,N_14093);
nand U17648 (N_17648,N_13242,N_13390);
nand U17649 (N_17649,N_12896,N_13660);
nor U17650 (N_17650,N_13799,N_13076);
nor U17651 (N_17651,N_12945,N_14829);
nand U17652 (N_17652,N_12837,N_12097);
nand U17653 (N_17653,N_13710,N_13636);
nor U17654 (N_17654,N_12439,N_13107);
xor U17655 (N_17655,N_12765,N_14639);
or U17656 (N_17656,N_12207,N_12147);
nor U17657 (N_17657,N_14586,N_14878);
nor U17658 (N_17658,N_13985,N_13970);
and U17659 (N_17659,N_14270,N_12617);
and U17660 (N_17660,N_13512,N_13966);
xor U17661 (N_17661,N_12224,N_13291);
or U17662 (N_17662,N_12511,N_13145);
and U17663 (N_17663,N_13405,N_14820);
or U17664 (N_17664,N_12266,N_12870);
or U17665 (N_17665,N_13282,N_14722);
nand U17666 (N_17666,N_13718,N_12037);
and U17667 (N_17667,N_14803,N_13766);
xor U17668 (N_17668,N_12557,N_13905);
xnor U17669 (N_17669,N_12171,N_13059);
nor U17670 (N_17670,N_14077,N_14414);
nand U17671 (N_17671,N_12476,N_13719);
and U17672 (N_17672,N_12217,N_14633);
xnor U17673 (N_17673,N_12873,N_14342);
xor U17674 (N_17674,N_12929,N_13796);
and U17675 (N_17675,N_13214,N_12142);
nand U17676 (N_17676,N_12116,N_14737);
and U17677 (N_17677,N_14794,N_13865);
nor U17678 (N_17678,N_13901,N_14856);
and U17679 (N_17679,N_14648,N_12690);
and U17680 (N_17680,N_14502,N_13960);
and U17681 (N_17681,N_14582,N_14401);
and U17682 (N_17682,N_13212,N_12857);
or U17683 (N_17683,N_14598,N_14711);
nor U17684 (N_17684,N_14816,N_13876);
and U17685 (N_17685,N_13645,N_14406);
or U17686 (N_17686,N_12143,N_14123);
xor U17687 (N_17687,N_12277,N_14132);
nor U17688 (N_17688,N_13685,N_12374);
or U17689 (N_17689,N_13647,N_14008);
nand U17690 (N_17690,N_13251,N_14186);
nand U17691 (N_17691,N_12071,N_13502);
xnor U17692 (N_17692,N_12644,N_13863);
xor U17693 (N_17693,N_13156,N_14097);
and U17694 (N_17694,N_13821,N_12035);
xnor U17695 (N_17695,N_14819,N_14879);
xnor U17696 (N_17696,N_13529,N_12629);
xor U17697 (N_17697,N_14738,N_14896);
or U17698 (N_17698,N_12929,N_13734);
or U17699 (N_17699,N_14341,N_14579);
nand U17700 (N_17700,N_12746,N_13215);
xnor U17701 (N_17701,N_12969,N_12335);
and U17702 (N_17702,N_12927,N_14010);
nor U17703 (N_17703,N_14039,N_14207);
nand U17704 (N_17704,N_12193,N_12536);
and U17705 (N_17705,N_14427,N_13922);
xnor U17706 (N_17706,N_12057,N_13508);
or U17707 (N_17707,N_13178,N_12818);
or U17708 (N_17708,N_13268,N_12162);
nand U17709 (N_17709,N_13154,N_12682);
and U17710 (N_17710,N_13150,N_12183);
and U17711 (N_17711,N_13955,N_13721);
and U17712 (N_17712,N_14335,N_12581);
xor U17713 (N_17713,N_13429,N_14630);
nand U17714 (N_17714,N_12280,N_12786);
or U17715 (N_17715,N_13678,N_13657);
xnor U17716 (N_17716,N_12161,N_14230);
nand U17717 (N_17717,N_13908,N_12264);
xor U17718 (N_17718,N_13971,N_14111);
xor U17719 (N_17719,N_13715,N_14245);
xnor U17720 (N_17720,N_14160,N_14472);
or U17721 (N_17721,N_14152,N_12466);
nand U17722 (N_17722,N_13057,N_13298);
or U17723 (N_17723,N_12327,N_14732);
xor U17724 (N_17724,N_13070,N_12514);
and U17725 (N_17725,N_13348,N_13962);
or U17726 (N_17726,N_12742,N_13203);
and U17727 (N_17727,N_12975,N_13219);
xnor U17728 (N_17728,N_13495,N_14656);
and U17729 (N_17729,N_14578,N_13621);
nand U17730 (N_17730,N_13004,N_13886);
or U17731 (N_17731,N_13491,N_13354);
nand U17732 (N_17732,N_14300,N_12425);
or U17733 (N_17733,N_13966,N_13742);
and U17734 (N_17734,N_12467,N_14290);
nor U17735 (N_17735,N_13300,N_13369);
nand U17736 (N_17736,N_14255,N_12378);
or U17737 (N_17737,N_13302,N_13085);
xnor U17738 (N_17738,N_12864,N_14003);
or U17739 (N_17739,N_12941,N_13069);
nor U17740 (N_17740,N_14404,N_13552);
nor U17741 (N_17741,N_12307,N_13000);
xor U17742 (N_17742,N_12939,N_14465);
or U17743 (N_17743,N_13146,N_12481);
nor U17744 (N_17744,N_14823,N_14014);
nor U17745 (N_17745,N_14651,N_12489);
and U17746 (N_17746,N_13299,N_14039);
or U17747 (N_17747,N_13800,N_12107);
nor U17748 (N_17748,N_14384,N_14540);
nand U17749 (N_17749,N_14831,N_13944);
xnor U17750 (N_17750,N_12630,N_14180);
or U17751 (N_17751,N_14982,N_14609);
nand U17752 (N_17752,N_13087,N_12572);
and U17753 (N_17753,N_13978,N_12379);
or U17754 (N_17754,N_13239,N_12317);
nand U17755 (N_17755,N_14639,N_12495);
xnor U17756 (N_17756,N_13176,N_13612);
nand U17757 (N_17757,N_12837,N_12617);
or U17758 (N_17758,N_13346,N_14627);
or U17759 (N_17759,N_13334,N_13021);
or U17760 (N_17760,N_12085,N_14002);
and U17761 (N_17761,N_13613,N_14083);
nand U17762 (N_17762,N_13809,N_12522);
or U17763 (N_17763,N_13629,N_13551);
or U17764 (N_17764,N_14462,N_14302);
xor U17765 (N_17765,N_12270,N_12328);
or U17766 (N_17766,N_14966,N_13287);
nand U17767 (N_17767,N_14390,N_13049);
and U17768 (N_17768,N_12523,N_13840);
xnor U17769 (N_17769,N_12005,N_13461);
nand U17770 (N_17770,N_13175,N_14262);
xor U17771 (N_17771,N_13438,N_13035);
nor U17772 (N_17772,N_13734,N_13444);
nor U17773 (N_17773,N_13883,N_12729);
or U17774 (N_17774,N_14045,N_14621);
or U17775 (N_17775,N_14310,N_12667);
or U17776 (N_17776,N_14131,N_12853);
and U17777 (N_17777,N_13157,N_12545);
nand U17778 (N_17778,N_12614,N_13861);
or U17779 (N_17779,N_13704,N_13788);
nand U17780 (N_17780,N_13505,N_12496);
or U17781 (N_17781,N_14182,N_14851);
nor U17782 (N_17782,N_13819,N_13081);
nand U17783 (N_17783,N_14683,N_13945);
xnor U17784 (N_17784,N_14980,N_12479);
nand U17785 (N_17785,N_12318,N_12224);
nor U17786 (N_17786,N_14183,N_13761);
nor U17787 (N_17787,N_14090,N_12194);
nor U17788 (N_17788,N_14667,N_14600);
nand U17789 (N_17789,N_14564,N_13828);
nand U17790 (N_17790,N_14874,N_14497);
and U17791 (N_17791,N_13247,N_13930);
or U17792 (N_17792,N_13433,N_12438);
nand U17793 (N_17793,N_14880,N_12094);
nor U17794 (N_17794,N_12287,N_14727);
or U17795 (N_17795,N_12721,N_14936);
and U17796 (N_17796,N_14760,N_12204);
nor U17797 (N_17797,N_13561,N_13898);
and U17798 (N_17798,N_12426,N_12385);
nor U17799 (N_17799,N_12635,N_13166);
nand U17800 (N_17800,N_13896,N_12138);
or U17801 (N_17801,N_14782,N_12174);
and U17802 (N_17802,N_12516,N_14573);
xnor U17803 (N_17803,N_14406,N_12530);
or U17804 (N_17804,N_13803,N_14022);
or U17805 (N_17805,N_13645,N_14132);
and U17806 (N_17806,N_12473,N_14482);
nor U17807 (N_17807,N_13042,N_14942);
nor U17808 (N_17808,N_14590,N_12470);
nand U17809 (N_17809,N_13883,N_14036);
nor U17810 (N_17810,N_13408,N_13082);
nor U17811 (N_17811,N_13514,N_12830);
nand U17812 (N_17812,N_14441,N_14876);
nand U17813 (N_17813,N_14277,N_12556);
nand U17814 (N_17814,N_14671,N_14074);
xor U17815 (N_17815,N_12194,N_12282);
and U17816 (N_17816,N_13174,N_14154);
nand U17817 (N_17817,N_12653,N_14697);
and U17818 (N_17818,N_14617,N_12397);
xnor U17819 (N_17819,N_14479,N_12639);
or U17820 (N_17820,N_13685,N_12412);
and U17821 (N_17821,N_13168,N_14861);
and U17822 (N_17822,N_14039,N_12386);
nand U17823 (N_17823,N_13630,N_12733);
and U17824 (N_17824,N_13068,N_12602);
and U17825 (N_17825,N_12084,N_12263);
nand U17826 (N_17826,N_14875,N_12123);
nor U17827 (N_17827,N_14586,N_14714);
and U17828 (N_17828,N_13127,N_14806);
nor U17829 (N_17829,N_12382,N_12283);
xnor U17830 (N_17830,N_12995,N_12981);
or U17831 (N_17831,N_12854,N_13084);
nand U17832 (N_17832,N_13032,N_12585);
xnor U17833 (N_17833,N_14044,N_14612);
or U17834 (N_17834,N_14153,N_13408);
nand U17835 (N_17835,N_12795,N_13464);
xnor U17836 (N_17836,N_12037,N_14112);
nand U17837 (N_17837,N_13035,N_12163);
nand U17838 (N_17838,N_14216,N_12811);
nand U17839 (N_17839,N_14304,N_14532);
nand U17840 (N_17840,N_12365,N_13103);
xnor U17841 (N_17841,N_12240,N_12258);
and U17842 (N_17842,N_13080,N_13983);
xnor U17843 (N_17843,N_13858,N_14280);
and U17844 (N_17844,N_14871,N_13228);
or U17845 (N_17845,N_14245,N_12427);
nand U17846 (N_17846,N_14280,N_14624);
xnor U17847 (N_17847,N_14468,N_13234);
xor U17848 (N_17848,N_13703,N_14231);
xor U17849 (N_17849,N_13118,N_14885);
xor U17850 (N_17850,N_12394,N_12047);
nor U17851 (N_17851,N_14844,N_13383);
or U17852 (N_17852,N_13976,N_14578);
and U17853 (N_17853,N_12837,N_14942);
nor U17854 (N_17854,N_14100,N_13762);
nor U17855 (N_17855,N_13728,N_12684);
nor U17856 (N_17856,N_13555,N_14769);
and U17857 (N_17857,N_14917,N_13877);
or U17858 (N_17858,N_13395,N_14380);
or U17859 (N_17859,N_14309,N_12406);
xnor U17860 (N_17860,N_14929,N_14162);
nor U17861 (N_17861,N_13118,N_12221);
and U17862 (N_17862,N_13674,N_12458);
or U17863 (N_17863,N_14540,N_13310);
xor U17864 (N_17864,N_13928,N_14305);
or U17865 (N_17865,N_13352,N_13917);
nand U17866 (N_17866,N_13134,N_12085);
nor U17867 (N_17867,N_14363,N_12824);
nand U17868 (N_17868,N_12505,N_13731);
or U17869 (N_17869,N_12765,N_13111);
xor U17870 (N_17870,N_13055,N_14112);
nand U17871 (N_17871,N_12715,N_14467);
or U17872 (N_17872,N_12409,N_14499);
and U17873 (N_17873,N_13356,N_13157);
nor U17874 (N_17874,N_14270,N_14685);
nor U17875 (N_17875,N_13309,N_12977);
nand U17876 (N_17876,N_13838,N_13450);
nand U17877 (N_17877,N_14030,N_12855);
nor U17878 (N_17878,N_14695,N_12990);
nand U17879 (N_17879,N_12154,N_14096);
or U17880 (N_17880,N_13054,N_13568);
xor U17881 (N_17881,N_12784,N_14309);
or U17882 (N_17882,N_14793,N_13334);
or U17883 (N_17883,N_12482,N_12576);
or U17884 (N_17884,N_12760,N_12830);
nand U17885 (N_17885,N_14971,N_12312);
or U17886 (N_17886,N_12169,N_12254);
and U17887 (N_17887,N_14186,N_13810);
nand U17888 (N_17888,N_12309,N_12793);
nor U17889 (N_17889,N_12732,N_13369);
or U17890 (N_17890,N_13968,N_13683);
nand U17891 (N_17891,N_13262,N_12410);
nor U17892 (N_17892,N_12282,N_12509);
nand U17893 (N_17893,N_13526,N_14178);
nand U17894 (N_17894,N_14335,N_14959);
xnor U17895 (N_17895,N_14732,N_13093);
xor U17896 (N_17896,N_14652,N_12658);
and U17897 (N_17897,N_13149,N_12731);
or U17898 (N_17898,N_12260,N_12653);
xnor U17899 (N_17899,N_12382,N_12939);
nor U17900 (N_17900,N_13636,N_12131);
nand U17901 (N_17901,N_14921,N_12458);
nand U17902 (N_17902,N_14583,N_12762);
or U17903 (N_17903,N_14707,N_14777);
nand U17904 (N_17904,N_13010,N_14621);
xor U17905 (N_17905,N_13352,N_12570);
xor U17906 (N_17906,N_14013,N_13870);
or U17907 (N_17907,N_14610,N_12451);
xnor U17908 (N_17908,N_12996,N_14647);
nor U17909 (N_17909,N_13031,N_12294);
or U17910 (N_17910,N_12178,N_13642);
xor U17911 (N_17911,N_12219,N_13058);
and U17912 (N_17912,N_13875,N_14527);
xnor U17913 (N_17913,N_14652,N_13184);
or U17914 (N_17914,N_12937,N_13929);
or U17915 (N_17915,N_12772,N_14070);
nor U17916 (N_17916,N_13852,N_12771);
xnor U17917 (N_17917,N_14046,N_13548);
or U17918 (N_17918,N_12554,N_14490);
nand U17919 (N_17919,N_13927,N_13391);
nor U17920 (N_17920,N_14658,N_14588);
or U17921 (N_17921,N_12434,N_14855);
nand U17922 (N_17922,N_12685,N_14438);
or U17923 (N_17923,N_14992,N_12331);
xor U17924 (N_17924,N_14707,N_14306);
or U17925 (N_17925,N_12467,N_12437);
xnor U17926 (N_17926,N_12490,N_14848);
and U17927 (N_17927,N_12983,N_14228);
and U17928 (N_17928,N_14899,N_14925);
or U17929 (N_17929,N_14011,N_14630);
and U17930 (N_17930,N_14696,N_14898);
or U17931 (N_17931,N_12105,N_12659);
nand U17932 (N_17932,N_12809,N_12126);
or U17933 (N_17933,N_12064,N_13567);
nand U17934 (N_17934,N_13498,N_13964);
or U17935 (N_17935,N_14386,N_13008);
nor U17936 (N_17936,N_12503,N_14441);
nand U17937 (N_17937,N_14350,N_14419);
and U17938 (N_17938,N_13751,N_13551);
nor U17939 (N_17939,N_14325,N_14062);
or U17940 (N_17940,N_12723,N_14870);
nor U17941 (N_17941,N_12035,N_13177);
or U17942 (N_17942,N_13224,N_13751);
nor U17943 (N_17943,N_14367,N_13832);
nand U17944 (N_17944,N_13498,N_12033);
nor U17945 (N_17945,N_14877,N_14747);
and U17946 (N_17946,N_13330,N_12485);
and U17947 (N_17947,N_12073,N_12279);
nor U17948 (N_17948,N_14596,N_12282);
xor U17949 (N_17949,N_13765,N_13227);
or U17950 (N_17950,N_13818,N_14237);
nand U17951 (N_17951,N_12166,N_14968);
nor U17952 (N_17952,N_13295,N_12607);
or U17953 (N_17953,N_12553,N_14580);
nor U17954 (N_17954,N_12622,N_12514);
nor U17955 (N_17955,N_14218,N_12464);
and U17956 (N_17956,N_14079,N_12197);
and U17957 (N_17957,N_12684,N_13324);
nor U17958 (N_17958,N_12601,N_12361);
and U17959 (N_17959,N_13752,N_14312);
or U17960 (N_17960,N_14137,N_12271);
or U17961 (N_17961,N_14357,N_14224);
or U17962 (N_17962,N_12202,N_12551);
nor U17963 (N_17963,N_12026,N_14976);
xor U17964 (N_17964,N_14800,N_12912);
or U17965 (N_17965,N_13371,N_13383);
and U17966 (N_17966,N_13133,N_13097);
xnor U17967 (N_17967,N_14344,N_12127);
xor U17968 (N_17968,N_12842,N_14985);
xor U17969 (N_17969,N_14403,N_14948);
nor U17970 (N_17970,N_14185,N_13165);
nor U17971 (N_17971,N_12616,N_12478);
xnor U17972 (N_17972,N_12478,N_13879);
xor U17973 (N_17973,N_13107,N_13473);
nand U17974 (N_17974,N_13911,N_14996);
and U17975 (N_17975,N_12371,N_13452);
and U17976 (N_17976,N_14414,N_14356);
nor U17977 (N_17977,N_12908,N_14499);
xor U17978 (N_17978,N_13825,N_13477);
nor U17979 (N_17979,N_14722,N_12508);
nor U17980 (N_17980,N_13086,N_12818);
xnor U17981 (N_17981,N_13604,N_14996);
nand U17982 (N_17982,N_12159,N_12967);
xor U17983 (N_17983,N_12784,N_12754);
and U17984 (N_17984,N_13461,N_12667);
or U17985 (N_17985,N_13495,N_12534);
nor U17986 (N_17986,N_14419,N_12167);
and U17987 (N_17987,N_13460,N_12965);
and U17988 (N_17988,N_13416,N_14830);
xnor U17989 (N_17989,N_14289,N_12515);
nor U17990 (N_17990,N_13843,N_14099);
nand U17991 (N_17991,N_14613,N_14815);
or U17992 (N_17992,N_14922,N_14558);
nand U17993 (N_17993,N_14396,N_14707);
and U17994 (N_17994,N_13931,N_13510);
nor U17995 (N_17995,N_13645,N_13229);
xnor U17996 (N_17996,N_13906,N_14998);
or U17997 (N_17997,N_13945,N_14666);
or U17998 (N_17998,N_12473,N_12519);
nand U17999 (N_17999,N_12006,N_12906);
xor U18000 (N_18000,N_15368,N_15567);
xor U18001 (N_18001,N_17936,N_16495);
nor U18002 (N_18002,N_16116,N_17365);
nor U18003 (N_18003,N_15172,N_15525);
and U18004 (N_18004,N_17712,N_16878);
and U18005 (N_18005,N_16625,N_15377);
xnor U18006 (N_18006,N_16520,N_15408);
and U18007 (N_18007,N_17143,N_16782);
or U18008 (N_18008,N_17681,N_17741);
nand U18009 (N_18009,N_16893,N_16390);
or U18010 (N_18010,N_17783,N_15969);
and U18011 (N_18011,N_16405,N_15034);
xor U18012 (N_18012,N_16820,N_17894);
xor U18013 (N_18013,N_16045,N_15621);
and U18014 (N_18014,N_17135,N_16688);
nand U18015 (N_18015,N_15836,N_17503);
nor U18016 (N_18016,N_15324,N_17256);
and U18017 (N_18017,N_16598,N_15346);
xnor U18018 (N_18018,N_15307,N_16616);
or U18019 (N_18019,N_16691,N_17015);
and U18020 (N_18020,N_17166,N_16169);
xor U18021 (N_18021,N_17163,N_15560);
nand U18022 (N_18022,N_15513,N_16106);
xnor U18023 (N_18023,N_16133,N_16997);
and U18024 (N_18024,N_15711,N_16319);
nand U18025 (N_18025,N_16504,N_17179);
nand U18026 (N_18026,N_15634,N_15350);
xnor U18027 (N_18027,N_16898,N_15618);
and U18028 (N_18028,N_17927,N_16995);
and U18029 (N_18029,N_16561,N_15680);
and U18030 (N_18030,N_17651,N_16917);
or U18031 (N_18031,N_15600,N_15370);
or U18032 (N_18032,N_16541,N_16177);
and U18033 (N_18033,N_15274,N_16971);
xor U18034 (N_18034,N_17563,N_15250);
nor U18035 (N_18035,N_17102,N_16939);
nor U18036 (N_18036,N_16124,N_15824);
xor U18037 (N_18037,N_16394,N_15966);
nor U18038 (N_18038,N_17835,N_16718);
nand U18039 (N_18039,N_15866,N_16784);
nand U18040 (N_18040,N_17603,N_15331);
nor U18041 (N_18041,N_17930,N_17650);
nor U18042 (N_18042,N_16547,N_16510);
or U18043 (N_18043,N_16373,N_17085);
nand U18044 (N_18044,N_17117,N_16522);
nor U18045 (N_18045,N_16258,N_15801);
or U18046 (N_18046,N_15890,N_15737);
and U18047 (N_18047,N_15811,N_16223);
nor U18048 (N_18048,N_16796,N_16257);
xor U18049 (N_18049,N_17730,N_15631);
or U18050 (N_18050,N_17279,N_16415);
xor U18051 (N_18051,N_17542,N_16368);
or U18052 (N_18052,N_17181,N_17668);
and U18053 (N_18053,N_16247,N_17373);
or U18054 (N_18054,N_17352,N_17857);
nand U18055 (N_18055,N_16723,N_17165);
and U18056 (N_18056,N_16352,N_17825);
nand U18057 (N_18057,N_17295,N_16243);
or U18058 (N_18058,N_17381,N_15336);
nand U18059 (N_18059,N_17514,N_17899);
or U18060 (N_18060,N_15017,N_15626);
nor U18061 (N_18061,N_17327,N_16089);
nor U18062 (N_18062,N_15786,N_16340);
or U18063 (N_18063,N_16629,N_15715);
xor U18064 (N_18064,N_16470,N_15552);
xnor U18065 (N_18065,N_17187,N_17746);
and U18066 (N_18066,N_15654,N_16166);
and U18067 (N_18067,N_17601,N_17891);
nor U18068 (N_18068,N_16052,N_16608);
or U18069 (N_18069,N_15135,N_17257);
and U18070 (N_18070,N_17366,N_15572);
nor U18071 (N_18071,N_17995,N_15716);
nor U18072 (N_18072,N_16865,N_17066);
nand U18073 (N_18073,N_16269,N_17680);
nand U18074 (N_18074,N_16010,N_15101);
nand U18075 (N_18075,N_17223,N_16099);
xor U18076 (N_18076,N_17579,N_15920);
and U18077 (N_18077,N_17199,N_17308);
nand U18078 (N_18078,N_17008,N_17644);
nor U18079 (N_18079,N_16392,N_17214);
nand U18080 (N_18080,N_15465,N_16699);
nand U18081 (N_18081,N_16197,N_16521);
nor U18082 (N_18082,N_15073,N_16739);
nand U18083 (N_18083,N_16426,N_16827);
nor U18084 (N_18084,N_15089,N_16492);
nand U18085 (N_18085,N_15774,N_15007);
xnor U18086 (N_18086,N_15526,N_15819);
or U18087 (N_18087,N_16057,N_15130);
and U18088 (N_18088,N_16696,N_16343);
nand U18089 (N_18089,N_16850,N_16653);
nor U18090 (N_18090,N_17659,N_16261);
nor U18091 (N_18091,N_15458,N_15499);
and U18092 (N_18092,N_15795,N_16551);
nor U18093 (N_18093,N_17531,N_17701);
nand U18094 (N_18094,N_15823,N_15293);
or U18095 (N_18095,N_15473,N_15476);
nand U18096 (N_18096,N_17148,N_17304);
nand U18097 (N_18097,N_17326,N_17598);
nor U18098 (N_18098,N_15975,N_15205);
nor U18099 (N_18099,N_15435,N_16256);
nor U18100 (N_18100,N_15687,N_15883);
and U18101 (N_18101,N_15486,N_17594);
and U18102 (N_18102,N_17753,N_16336);
or U18103 (N_18103,N_15178,N_16412);
or U18104 (N_18104,N_16557,N_15676);
nand U18105 (N_18105,N_15049,N_16966);
or U18106 (N_18106,N_15629,N_15867);
and U18107 (N_18107,N_17617,N_17404);
or U18108 (N_18108,N_16081,N_17149);
or U18109 (N_18109,N_15599,N_17255);
and U18110 (N_18110,N_15538,N_16095);
and U18111 (N_18111,N_15997,N_17299);
xnor U18112 (N_18112,N_15053,N_17465);
nor U18113 (N_18113,N_15899,N_16981);
nor U18114 (N_18114,N_15507,N_17582);
and U18115 (N_18115,N_16437,N_17915);
or U18116 (N_18116,N_15218,N_17971);
nor U18117 (N_18117,N_15758,N_16952);
nor U18118 (N_18118,N_15903,N_17168);
or U18119 (N_18119,N_16601,N_15134);
or U18120 (N_18120,N_16158,N_15059);
nand U18121 (N_18121,N_15886,N_15396);
or U18122 (N_18122,N_15672,N_17926);
xnor U18123 (N_18123,N_15229,N_15865);
xnor U18124 (N_18124,N_16769,N_15561);
nor U18125 (N_18125,N_16974,N_17072);
nand U18126 (N_18126,N_17131,N_15647);
nor U18127 (N_18127,N_15694,N_16906);
nor U18128 (N_18128,N_15490,N_16185);
nor U18129 (N_18129,N_15138,N_16051);
and U18130 (N_18130,N_17377,N_15746);
xor U18131 (N_18131,N_15963,N_15166);
nor U18132 (N_18132,N_17948,N_17739);
or U18133 (N_18133,N_15853,N_16056);
xnor U18134 (N_18134,N_17750,N_16485);
and U18135 (N_18135,N_15074,N_16559);
xnor U18136 (N_18136,N_15231,N_15553);
or U18137 (N_18137,N_15998,N_17482);
and U18138 (N_18138,N_15937,N_17436);
and U18139 (N_18139,N_17871,N_15832);
nor U18140 (N_18140,N_17541,N_16190);
nand U18141 (N_18141,N_15285,N_16369);
nand U18142 (N_18142,N_15203,N_17050);
nand U18143 (N_18143,N_17128,N_15400);
or U18144 (N_18144,N_17405,N_16728);
xnor U18145 (N_18145,N_17578,N_17538);
or U18146 (N_18146,N_17422,N_16867);
nor U18147 (N_18147,N_15539,N_16754);
nor U18148 (N_18148,N_17252,N_17283);
xor U18149 (N_18149,N_15273,N_17147);
xor U18150 (N_18150,N_15682,N_16722);
xor U18151 (N_18151,N_16466,N_15712);
or U18152 (N_18152,N_17061,N_15095);
or U18153 (N_18153,N_16672,N_16473);
and U18154 (N_18154,N_15121,N_17878);
nand U18155 (N_18155,N_17609,N_17637);
or U18156 (N_18156,N_16710,N_15357);
nand U18157 (N_18157,N_16249,N_16229);
or U18158 (N_18158,N_16170,N_15728);
xor U18159 (N_18159,N_17743,N_16685);
and U18160 (N_18160,N_17953,N_16174);
xnor U18161 (N_18161,N_16970,N_16076);
or U18162 (N_18162,N_16799,N_16950);
nand U18163 (N_18163,N_17307,N_15536);
and U18164 (N_18164,N_15642,N_15768);
nand U18165 (N_18165,N_15943,N_17216);
nor U18166 (N_18166,N_16125,N_16160);
nand U18167 (N_18167,N_16073,N_15117);
nor U18168 (N_18168,N_15126,N_17121);
or U18169 (N_18169,N_17488,N_15615);
or U18170 (N_18170,N_16749,N_15663);
nand U18171 (N_18171,N_16862,N_16586);
or U18172 (N_18172,N_15338,N_15511);
nor U18173 (N_18173,N_15762,N_16102);
xnor U18174 (N_18174,N_16254,N_16640);
nand U18175 (N_18175,N_15308,N_15448);
nor U18176 (N_18176,N_15748,N_15419);
xor U18177 (N_18177,N_15945,N_16695);
or U18178 (N_18178,N_17144,N_17711);
nor U18179 (N_18179,N_16425,N_16980);
nor U18180 (N_18180,N_16323,N_16617);
or U18181 (N_18181,N_17839,N_15732);
and U18182 (N_18182,N_17720,N_16539);
and U18183 (N_18183,N_17842,N_15988);
nand U18184 (N_18184,N_15453,N_17454);
or U18185 (N_18185,N_16015,N_16355);
xnor U18186 (N_18186,N_16128,N_16932);
nand U18187 (N_18187,N_16698,N_17966);
nor U18188 (N_18188,N_15718,N_16578);
xor U18189 (N_18189,N_15688,N_15147);
nor U18190 (N_18190,N_15692,N_17790);
xnor U18191 (N_18191,N_15857,N_17905);
or U18192 (N_18192,N_17397,N_15472);
nor U18193 (N_18193,N_15043,N_16849);
nor U18194 (N_18194,N_16940,N_17274);
or U18195 (N_18195,N_17303,N_15504);
and U18196 (N_18196,N_16476,N_17374);
nand U18197 (N_18197,N_16549,N_17254);
nand U18198 (N_18198,N_17133,N_17778);
and U18199 (N_18199,N_15420,N_15403);
and U18200 (N_18200,N_16484,N_17054);
nand U18201 (N_18201,N_17230,N_16419);
nand U18202 (N_18202,N_16227,N_15763);
and U18203 (N_18203,N_15780,N_17105);
nor U18204 (N_18204,N_16948,N_17607);
xnor U18205 (N_18205,N_17885,N_16575);
xnor U18206 (N_18206,N_16304,N_17799);
and U18207 (N_18207,N_16202,N_15120);
and U18208 (N_18208,N_17378,N_15882);
xnor U18209 (N_18209,N_17947,N_16915);
xor U18210 (N_18210,N_16988,N_17771);
or U18211 (N_18211,N_16292,N_15924);
or U18212 (N_18212,N_15141,N_16212);
nand U18213 (N_18213,N_17992,N_15702);
and U18214 (N_18214,N_15657,N_17747);
and U18215 (N_18215,N_16667,N_16609);
xor U18216 (N_18216,N_17840,N_16322);
or U18217 (N_18217,N_16705,N_16218);
xor U18218 (N_18218,N_17889,N_17698);
nor U18219 (N_18219,N_15411,N_16524);
nor U18220 (N_18220,N_16221,N_16448);
or U18221 (N_18221,N_16478,N_15311);
xor U18222 (N_18222,N_16398,N_17073);
or U18223 (N_18223,N_16280,N_16807);
nand U18224 (N_18224,N_15491,N_15829);
xnor U18225 (N_18225,N_16025,N_17587);
or U18226 (N_18226,N_17564,N_15952);
and U18227 (N_18227,N_15955,N_15393);
xor U18228 (N_18228,N_16897,N_15656);
nand U18229 (N_18229,N_15257,N_16758);
nand U18230 (N_18230,N_15651,N_15846);
nor U18231 (N_18231,N_16297,N_15689);
xor U18232 (N_18232,N_15805,N_16930);
and U18233 (N_18233,N_17850,N_15330);
nor U18234 (N_18234,N_17934,N_15830);
nor U18235 (N_18235,N_15481,N_15840);
xnor U18236 (N_18236,N_15785,N_15287);
nand U18237 (N_18237,N_15013,N_15183);
and U18238 (N_18238,N_17464,N_15484);
and U18239 (N_18239,N_17424,N_17445);
nand U18240 (N_18240,N_17142,N_17824);
or U18241 (N_18241,N_16555,N_15045);
xnor U18242 (N_18242,N_16509,N_16381);
nor U18243 (N_18243,N_15091,N_15399);
xor U18244 (N_18244,N_17776,N_16353);
nor U18245 (N_18245,N_15496,N_17211);
xnor U18246 (N_18246,N_17939,N_17146);
and U18247 (N_18247,N_16331,N_16922);
and U18248 (N_18248,N_17290,N_15301);
and U18249 (N_18249,N_16498,N_17826);
or U18250 (N_18250,N_15217,N_16721);
or U18251 (N_18251,N_16921,N_16645);
or U18252 (N_18252,N_17141,N_15046);
nor U18253 (N_18253,N_15123,N_16196);
xor U18254 (N_18254,N_17034,N_15317);
and U18255 (N_18255,N_15014,N_16211);
nand U18256 (N_18256,N_16112,N_17717);
or U18257 (N_18257,N_15508,N_15910);
nand U18258 (N_18258,N_15838,N_16761);
or U18259 (N_18259,N_15204,N_16067);
xor U18260 (N_18260,N_15442,N_15165);
nor U18261 (N_18261,N_15637,N_15220);
or U18262 (N_18262,N_15674,N_16277);
nor U18263 (N_18263,N_17942,N_15666);
or U18264 (N_18264,N_17756,N_17497);
or U18265 (N_18265,N_15582,N_16454);
nor U18266 (N_18266,N_16533,N_15421);
or U18267 (N_18267,N_16738,N_15455);
xor U18268 (N_18268,N_16287,N_16872);
xnor U18269 (N_18269,N_17537,N_15133);
or U18270 (N_18270,N_15885,N_17870);
xnor U18271 (N_18271,N_15518,N_17569);
or U18272 (N_18272,N_15608,N_17353);
nand U18273 (N_18273,N_15437,N_15497);
xnor U18274 (N_18274,N_15213,N_15787);
and U18275 (N_18275,N_15489,N_16386);
or U18276 (N_18276,N_17493,N_16725);
and U18277 (N_18277,N_16389,N_16194);
and U18278 (N_18278,N_16604,N_15392);
nor U18279 (N_18279,N_16975,N_15658);
or U18280 (N_18280,N_16902,N_16821);
nand U18281 (N_18281,N_17392,N_15793);
or U18282 (N_18282,N_15207,N_17626);
nor U18283 (N_18283,N_16456,N_17757);
and U18284 (N_18284,N_16765,N_16399);
and U18285 (N_18285,N_16181,N_17703);
or U18286 (N_18286,N_17184,N_17620);
and U18287 (N_18287,N_16032,N_15429);
or U18288 (N_18288,N_15054,N_17551);
nand U18289 (N_18289,N_15964,N_16508);
xor U18290 (N_18290,N_17173,N_16162);
or U18291 (N_18291,N_15784,N_17055);
nor U18292 (N_18292,N_17411,N_15241);
nor U18293 (N_18293,N_16395,N_15256);
or U18294 (N_18294,N_17190,N_15747);
and U18295 (N_18295,N_16204,N_15949);
or U18296 (N_18296,N_15659,N_16839);
or U18297 (N_18297,N_15816,N_16383);
or U18298 (N_18298,N_17232,N_16724);
and U18299 (N_18299,N_16517,N_17595);
or U18300 (N_18300,N_15551,N_16318);
or U18301 (N_18301,N_15083,N_15474);
nor U18302 (N_18302,N_15136,N_17820);
nor U18303 (N_18303,N_17629,N_16942);
or U18304 (N_18304,N_17244,N_15398);
nor U18305 (N_18305,N_15036,N_16733);
or U18306 (N_18306,N_17762,N_16363);
nor U18307 (N_18307,N_15590,N_15556);
or U18308 (N_18308,N_17566,N_16358);
or U18309 (N_18309,N_16016,N_16283);
or U18310 (N_18310,N_16063,N_17913);
nor U18311 (N_18311,N_15451,N_15105);
or U18312 (N_18312,N_16475,N_16251);
xnor U18313 (N_18313,N_16994,N_15833);
and U18314 (N_18314,N_15757,N_16438);
xor U18315 (N_18315,N_16944,N_17047);
nand U18316 (N_18316,N_16104,N_15641);
and U18317 (N_18317,N_16387,N_17911);
nand U18318 (N_18318,N_16396,N_15972);
and U18319 (N_18319,N_15628,N_15807);
xnor U18320 (N_18320,N_15669,N_17896);
and U18321 (N_18321,N_17805,N_15253);
nand U18322 (N_18322,N_16018,N_17386);
or U18323 (N_18323,N_16071,N_17170);
and U18324 (N_18324,N_17237,N_16896);
and U18325 (N_18325,N_15655,N_16823);
nand U18326 (N_18326,N_17127,N_15635);
nand U18327 (N_18327,N_15861,N_17113);
and U18328 (N_18328,N_16191,N_16468);
or U18329 (N_18329,N_16694,N_15144);
nand U18330 (N_18330,N_15334,N_17003);
nor U18331 (N_18331,N_16819,N_15827);
xor U18332 (N_18332,N_16459,N_17636);
nor U18333 (N_18333,N_17343,N_15340);
xnor U18334 (N_18334,N_17688,N_16631);
xor U18335 (N_18335,N_16615,N_15164);
nor U18336 (N_18336,N_17276,N_15322);
or U18337 (N_18337,N_16420,N_15443);
xnor U18338 (N_18338,N_16450,N_17337);
nand U18339 (N_18339,N_15825,N_15543);
xor U18340 (N_18340,N_16883,N_16963);
xor U18341 (N_18341,N_16458,N_15848);
and U18342 (N_18342,N_15516,N_15528);
and U18343 (N_18343,N_16841,N_15367);
and U18344 (N_18344,N_15261,N_16829);
or U18345 (N_18345,N_16690,N_17075);
or U18346 (N_18346,N_16856,N_17695);
xnor U18347 (N_18347,N_17263,N_17819);
nand U18348 (N_18348,N_17961,N_15452);
xor U18349 (N_18349,N_17027,N_15585);
xor U18350 (N_18350,N_16577,N_17038);
and U18351 (N_18351,N_16644,N_16416);
nor U18352 (N_18352,N_17413,N_16637);
xor U18353 (N_18353,N_16764,N_15173);
nand U18354 (N_18354,N_17818,N_15817);
and U18355 (N_18355,N_17065,N_17409);
or U18356 (N_18356,N_17388,N_16595);
or U18357 (N_18357,N_17322,N_15765);
nand U18358 (N_18358,N_15850,N_17094);
and U18359 (N_18359,N_15990,N_16082);
xnor U18360 (N_18360,N_16719,N_16585);
or U18361 (N_18361,N_15559,N_16656);
and U18362 (N_18362,N_17396,N_17811);
xnor U18363 (N_18363,N_17051,N_16147);
or U18364 (N_18364,N_15303,N_16424);
nor U18365 (N_18365,N_15100,N_17410);
and U18366 (N_18366,N_17647,N_16665);
or U18367 (N_18367,N_16193,N_15546);
nand U18368 (N_18368,N_15313,N_15610);
nand U18369 (N_18369,N_17286,N_16774);
nor U18370 (N_18370,N_15500,N_15877);
or U18371 (N_18371,N_16418,N_16511);
and U18372 (N_18372,N_15364,N_16252);
nand U18373 (N_18373,N_15245,N_17954);
or U18374 (N_18374,N_17605,N_17585);
or U18375 (N_18375,N_17432,N_16597);
nand U18376 (N_18376,N_15871,N_15035);
xor U18377 (N_18377,N_16792,N_17275);
nand U18378 (N_18378,N_15271,N_16427);
and U18379 (N_18379,N_15001,N_16977);
nor U18380 (N_18380,N_17555,N_16746);
nor U18381 (N_18381,N_17340,N_17952);
nand U18382 (N_18382,N_15015,N_16027);
nand U18383 (N_18383,N_15032,N_15810);
nor U18384 (N_18384,N_16003,N_17116);
nand U18385 (N_18385,N_16845,N_15971);
and U18386 (N_18386,N_16143,N_15932);
or U18387 (N_18387,N_17728,N_17266);
or U18388 (N_18388,N_17649,N_16235);
or U18389 (N_18389,N_17421,N_16033);
nor U18390 (N_18390,N_15480,N_16793);
and U18391 (N_18391,N_15695,N_17922);
nand U18392 (N_18392,N_17002,N_16264);
or U18393 (N_18393,N_15304,N_16668);
nand U18394 (N_18394,N_16164,N_17191);
xor U18395 (N_18395,N_17202,N_17914);
or U18396 (N_18396,N_16430,N_15510);
xor U18397 (N_18397,N_15412,N_15351);
nor U18398 (N_18398,N_15961,N_16567);
or U18399 (N_18399,N_15246,N_17964);
and U18400 (N_18400,N_17821,N_16186);
and U18401 (N_18401,N_17705,N_17780);
xnor U18402 (N_18402,N_16350,N_16781);
xnor U18403 (N_18403,N_16907,N_17990);
xor U18404 (N_18404,N_17260,N_17249);
nand U18405 (N_18405,N_17658,N_17986);
and U18406 (N_18406,N_17735,N_17156);
or U18407 (N_18407,N_17502,N_17732);
xor U18408 (N_18408,N_17796,N_17526);
xnor U18409 (N_18409,N_16836,N_15620);
xnor U18410 (N_18410,N_17597,N_15354);
nand U18411 (N_18411,N_15189,N_15265);
nand U18412 (N_18412,N_16298,N_16713);
and U18413 (N_18413,N_17134,N_16619);
and U18414 (N_18414,N_16863,N_15337);
nand U18415 (N_18415,N_17226,N_16624);
xor U18416 (N_18416,N_17250,N_17999);
and U18417 (N_18417,N_16926,N_15162);
nor U18418 (N_18418,N_17028,N_17646);
or U18419 (N_18419,N_15921,N_15995);
nand U18420 (N_18420,N_15630,N_16927);
nand U18421 (N_18421,N_16242,N_16382);
nand U18422 (N_18422,N_17364,N_15869);
nor U18423 (N_18423,N_16432,N_16550);
and U18424 (N_18424,N_15815,N_15740);
nor U18425 (N_18425,N_15065,N_16660);
and U18426 (N_18426,N_17440,N_17606);
xor U18427 (N_18427,N_16041,N_15167);
nand U18428 (N_18428,N_16832,N_15859);
and U18429 (N_18429,N_17074,N_17185);
nor U18430 (N_18430,N_16145,N_16880);
or U18431 (N_18431,N_15005,N_17760);
nor U18432 (N_18432,N_16013,N_15569);
nand U18433 (N_18433,N_17511,N_15422);
and U18434 (N_18434,N_17363,N_17315);
nand U18435 (N_18435,N_16982,N_15096);
and U18436 (N_18436,N_16462,N_17063);
or U18437 (N_18437,N_17692,N_15640);
xnor U18438 (N_18438,N_17469,N_17604);
nor U18439 (N_18439,N_15122,N_15532);
xor U18440 (N_18440,N_17689,N_17235);
nor U18441 (N_18441,N_17151,N_16881);
nor U18442 (N_18442,N_17349,N_17407);
xor U18443 (N_18443,N_16712,N_17662);
or U18444 (N_18444,N_16360,N_17985);
or U18445 (N_18445,N_15826,N_17096);
nand U18446 (N_18446,N_17434,N_15025);
nand U18447 (N_18447,N_15703,N_16736);
xnor U18448 (N_18448,N_15349,N_15845);
nor U18449 (N_18449,N_17838,N_15232);
and U18450 (N_18450,N_17809,N_16537);
nor U18451 (N_18451,N_17356,N_16161);
nor U18452 (N_18452,N_15382,N_15520);
nor U18453 (N_18453,N_16490,N_17849);
xor U18454 (N_18454,N_16080,N_15450);
xor U18455 (N_18455,N_16641,N_17175);
or U18456 (N_18456,N_15649,N_16599);
and U18457 (N_18457,N_17246,N_15228);
or U18458 (N_18458,N_15487,N_16487);
and U18459 (N_18459,N_17916,N_16934);
nand U18460 (N_18460,N_16078,N_17892);
or U18461 (N_18461,N_15872,N_15940);
nor U18462 (N_18462,N_17158,N_17494);
nand U18463 (N_18463,N_17860,N_17748);
or U18464 (N_18464,N_15206,N_17476);
xor U18465 (N_18465,N_16961,N_15870);
nand U18466 (N_18466,N_15644,N_17622);
xnor U18467 (N_18467,N_15233,N_16518);
and U18468 (N_18468,N_16515,N_15447);
nor U18469 (N_18469,N_16855,N_15544);
xnor U18470 (N_18470,N_16762,N_17420);
or U18471 (N_18471,N_15247,N_15925);
xor U18472 (N_18472,N_17517,N_15353);
xor U18473 (N_18473,N_16763,N_16851);
nand U18474 (N_18474,N_15851,N_15352);
nand U18475 (N_18475,N_16650,N_16936);
nor U18476 (N_18476,N_16742,N_15057);
nand U18477 (N_18477,N_17157,N_15316);
and U18478 (N_18478,N_16065,N_17361);
nor U18479 (N_18479,N_17103,N_17462);
or U18480 (N_18480,N_16532,N_16467);
and U18481 (N_18481,N_16516,N_17251);
or U18482 (N_18482,N_17040,N_15729);
and U18483 (N_18483,N_16060,N_16421);
or U18484 (N_18484,N_15031,N_15799);
and U18485 (N_18485,N_16132,N_17714);
and U18486 (N_18486,N_16852,N_16131);
nor U18487 (N_18487,N_16957,N_17877);
xnor U18488 (N_18488,N_16876,N_15426);
and U18489 (N_18489,N_16529,N_17160);
and U18490 (N_18490,N_16165,N_17836);
nand U18491 (N_18491,N_16805,N_15200);
or U18492 (N_18492,N_15591,N_15214);
xor U18493 (N_18493,N_16877,N_16964);
and U18494 (N_18494,N_17457,N_17793);
nor U18495 (N_18495,N_17794,N_15991);
xor U18496 (N_18496,N_15770,N_16565);
xor U18497 (N_18497,N_17600,N_17989);
and U18498 (N_18498,N_16324,N_16136);
and U18499 (N_18499,N_17044,N_17236);
nor U18500 (N_18500,N_15915,N_16813);
nand U18501 (N_18501,N_17929,N_15535);
nor U18502 (N_18502,N_17874,N_17602);
and U18503 (N_18503,N_15255,N_16810);
or U18504 (N_18504,N_16436,N_16357);
nor U18505 (N_18505,N_16693,N_16684);
xor U18506 (N_18506,N_16916,N_17568);
nand U18507 (N_18507,N_17625,N_16452);
nor U18508 (N_18508,N_17956,N_15668);
nor U18509 (N_18509,N_17431,N_15461);
or U18510 (N_18510,N_15363,N_16070);
xor U18511 (N_18511,N_17285,N_16226);
nor U18512 (N_18512,N_16613,N_17830);
xnor U18513 (N_18513,N_15194,N_16978);
xnor U18514 (N_18514,N_15583,N_17145);
nor U18515 (N_18515,N_15727,N_17248);
or U18516 (N_18516,N_15427,N_15153);
xor U18517 (N_18517,N_17522,N_16777);
xnor U18518 (N_18518,N_15822,N_16903);
nand U18519 (N_18519,N_16587,N_15471);
or U18520 (N_18520,N_15098,N_15140);
nor U18521 (N_18521,N_17227,N_16026);
nand U18522 (N_18522,N_16138,N_17509);
or U18523 (N_18523,N_15835,N_15433);
or U18524 (N_18524,N_17543,N_17451);
nor U18525 (N_18525,N_15752,N_15606);
nor U18526 (N_18526,N_16680,N_17708);
xnor U18527 (N_18527,N_17686,N_15283);
and U18528 (N_18528,N_15800,N_17459);
nor U18529 (N_18529,N_16449,N_16905);
xnor U18530 (N_18530,N_17499,N_15375);
xor U18531 (N_18531,N_17106,N_15298);
nand U18532 (N_18532,N_17376,N_15596);
and U18533 (N_18533,N_16726,N_15066);
nand U18534 (N_18534,N_15697,N_15965);
xor U18535 (N_18535,N_17855,N_17053);
or U18536 (N_18536,N_15062,N_15934);
or U18537 (N_18537,N_16985,N_17975);
nor U18538 (N_18538,N_15084,N_17866);
nor U18539 (N_18539,N_15388,N_15683);
xor U18540 (N_18540,N_16664,N_16176);
nor U18541 (N_18541,N_17501,N_15962);
and U18542 (N_18542,N_15266,N_17919);
and U18543 (N_18543,N_16711,N_15327);
xor U18544 (N_18544,N_16825,N_17725);
and U18545 (N_18545,N_16707,N_17507);
xor U18546 (N_18546,N_15477,N_16703);
xor U18547 (N_18547,N_16811,N_17946);
nor U18548 (N_18548,N_15956,N_17415);
nand U18549 (N_18549,N_16224,N_16795);
xnor U18550 (N_18550,N_15858,N_16992);
and U18551 (N_18551,N_16141,N_16914);
and U18552 (N_18552,N_15061,N_17492);
or U18553 (N_18553,N_16861,N_15554);
and U18554 (N_18554,N_17957,N_15542);
and U18555 (N_18555,N_17931,N_17908);
xor U18556 (N_18556,N_16195,N_15002);
xor U18557 (N_18557,N_15158,N_17974);
xnor U18558 (N_18558,N_15580,N_16417);
nor U18559 (N_18559,N_16759,N_17092);
xor U18560 (N_18560,N_15169,N_15482);
and U18561 (N_18561,N_16816,N_16442);
or U18562 (N_18562,N_15930,N_16822);
nand U18563 (N_18563,N_15063,N_17547);
nor U18564 (N_18564,N_16009,N_16499);
nor U18565 (N_18565,N_17675,N_16960);
nor U18566 (N_18566,N_17119,N_16666);
xor U18567 (N_18567,N_15996,N_17076);
xor U18568 (N_18568,N_15439,N_17172);
and U18569 (N_18569,N_15679,N_17525);
nor U18570 (N_18570,N_17897,N_15613);
xnor U18571 (N_18571,N_15685,N_15874);
or U18572 (N_18572,N_16377,N_15386);
nand U18573 (N_18573,N_16201,N_17864);
and U18574 (N_18574,N_16225,N_16072);
nand U18575 (N_18575,N_16238,N_17242);
or U18576 (N_18576,N_15821,N_17697);
and U18577 (N_18577,N_17486,N_15282);
nand U18578 (N_18578,N_15562,N_16361);
and U18579 (N_18579,N_17463,N_16607);
or U18580 (N_18580,N_15440,N_15633);
nor U18581 (N_18581,N_15696,N_15794);
nand U18582 (N_18582,N_15743,N_15754);
xor U18583 (N_18583,N_17473,N_17635);
nand U18584 (N_18584,N_15739,N_17408);
and U18585 (N_18585,N_15441,N_17539);
nor U18586 (N_18586,N_15994,N_15258);
and U18587 (N_18587,N_17311,N_15802);
xor U18588 (N_18588,N_17777,N_15478);
or U18589 (N_18589,N_15385,N_16828);
nor U18590 (N_18590,N_17847,N_15111);
xor U18591 (N_18591,N_17567,N_15589);
or U18592 (N_18592,N_17091,N_15201);
xnor U18593 (N_18593,N_15783,N_15960);
nand U18594 (N_18594,N_17903,N_17430);
xor U18595 (N_18595,N_17673,N_16801);
nand U18596 (N_18596,N_15109,N_16008);
nand U18597 (N_18597,N_16962,N_15366);
or U18598 (N_18598,N_16864,N_17443);
or U18599 (N_18599,N_15010,N_15725);
xor U18600 (N_18600,N_15395,N_16513);
nor U18601 (N_18601,N_16366,N_16127);
and U18602 (N_18602,N_15212,N_16919);
or U18603 (N_18603,N_17460,N_16757);
nor U18604 (N_18604,N_17480,N_16920);
nor U18605 (N_18605,N_17736,N_15907);
nand U18606 (N_18606,N_15113,N_15011);
nand U18607 (N_18607,N_16376,N_17297);
and U18608 (N_18608,N_17262,N_17982);
nor U18609 (N_18609,N_17487,N_16263);
xnor U18610 (N_18610,N_16255,N_16122);
nor U18611 (N_18611,N_15286,N_17576);
xor U18612 (N_18612,N_16312,N_16384);
xor U18613 (N_18613,N_15974,N_16843);
nand U18614 (N_18614,N_15855,N_17225);
or U18615 (N_18615,N_16649,N_16012);
nand U18616 (N_18616,N_17755,N_17391);
nor U18617 (N_18617,N_17767,N_17114);
xor U18618 (N_18618,N_16054,N_16958);
nand U18619 (N_18619,N_16407,N_16274);
and U18620 (N_18620,N_17446,N_15047);
nor U18621 (N_18621,N_17484,N_16286);
xor U18622 (N_18622,N_17412,N_16737);
xor U18623 (N_18623,N_16941,N_15008);
or U18624 (N_18624,N_15839,N_15678);
nand U18625 (N_18625,N_17983,N_17702);
xor U18626 (N_18626,N_15417,N_16623);
and U18627 (N_18627,N_16661,N_16313);
or U18628 (N_18628,N_15731,N_16605);
nand U18629 (N_18629,N_15502,N_15106);
xnor U18630 (N_18630,N_16972,N_15190);
and U18631 (N_18631,N_17150,N_15917);
nor U18632 (N_18632,N_16512,N_15104);
xnor U18633 (N_18633,N_17313,N_16891);
xnor U18634 (N_18634,N_17081,N_16446);
nand U18635 (N_18635,N_15180,N_15936);
and U18636 (N_18636,N_16523,N_17222);
nor U18637 (N_18637,N_15459,N_15533);
nand U18638 (N_18638,N_17331,N_17657);
nand U18639 (N_18639,N_16847,N_16835);
or U18640 (N_18640,N_16791,N_15645);
nand U18641 (N_18641,N_17271,N_15778);
nand U18642 (N_18642,N_15160,N_17310);
or U18643 (N_18643,N_16059,N_16479);
nand U18644 (N_18644,N_17631,N_16031);
nor U18645 (N_18645,N_17928,N_17959);
nor U18646 (N_18646,N_17853,N_17037);
nand U18647 (N_18647,N_17592,N_17155);
and U18648 (N_18648,N_16734,N_15044);
nor U18649 (N_18649,N_17513,N_17973);
nor U18650 (N_18650,N_16094,N_16134);
nand U18651 (N_18651,N_16976,N_15958);
nand U18652 (N_18652,N_16818,N_15812);
xor U18653 (N_18653,N_15849,N_15196);
xor U18654 (N_18654,N_17475,N_15977);
and U18655 (N_18655,N_17022,N_17344);
and U18656 (N_18656,N_16077,N_15197);
nor U18657 (N_18657,N_15248,N_16745);
or U18658 (N_18658,N_16594,N_17846);
nand U18659 (N_18659,N_16496,N_17880);
or U18660 (N_18660,N_17329,N_17898);
nor U18661 (N_18661,N_17231,N_16556);
xor U18662 (N_18662,N_16590,N_17640);
and U18663 (N_18663,N_16655,N_16538);
xnor U18664 (N_18664,N_17233,N_15856);
nor U18665 (N_18665,N_16182,N_17292);
nor U18666 (N_18666,N_15753,N_15627);
xnor U18667 (N_18667,N_15720,N_16047);
nor U18668 (N_18668,N_15012,N_17084);
nor U18669 (N_18669,N_15436,N_16760);
and U18670 (N_18670,N_17784,N_17371);
or U18671 (N_18671,N_17584,N_16403);
and U18672 (N_18672,N_17280,N_17951);
xnor U18673 (N_18673,N_17162,N_17791);
xnor U18674 (N_18674,N_16453,N_17192);
and U18675 (N_18675,N_16447,N_16780);
nand U18676 (N_18676,N_15092,N_17940);
or U18677 (N_18677,N_17367,N_17071);
xor U18678 (N_18678,N_17512,N_17282);
xor U18679 (N_18679,N_15760,N_17764);
xnor U18680 (N_18680,N_16114,N_15310);
and U18681 (N_18681,N_17571,N_15923);
nand U18682 (N_18682,N_17960,N_17766);
and U18683 (N_18683,N_16118,N_15094);
xnor U18684 (N_18684,N_16959,N_16494);
nand U18685 (N_18685,N_17140,N_15574);
and U18686 (N_18686,N_17333,N_16671);
and U18687 (N_18687,N_15380,N_16325);
or U18688 (N_18688,N_16678,N_15456);
and U18689 (N_18689,N_15792,N_17289);
and U18690 (N_18690,N_17997,N_17925);
or U18691 (N_18691,N_16612,N_16216);
xnor U18692 (N_18692,N_16560,N_16873);
or U18693 (N_18693,N_16282,N_15110);
xor U18694 (N_18694,N_17379,N_17580);
and U18695 (N_18695,N_17902,N_16004);
or U18696 (N_18696,N_17123,N_16267);
nand U18697 (N_18697,N_15129,N_17213);
nand U18698 (N_18698,N_15522,N_17895);
nand U18699 (N_18699,N_17833,N_17876);
nor U18700 (N_18700,N_15803,N_17048);
or U18701 (N_18701,N_15726,N_15643);
nand U18702 (N_18702,N_15404,N_16682);
nor U18703 (N_18703,N_16246,N_15305);
nand U18704 (N_18704,N_16569,N_15415);
nor U18705 (N_18705,N_16349,N_17057);
or U18706 (N_18706,N_17089,N_15254);
nand U18707 (N_18707,N_17270,N_16752);
nor U18708 (N_18708,N_16779,N_16083);
and U18709 (N_18709,N_17416,N_15900);
and U18710 (N_18710,N_15128,N_17769);
or U18711 (N_18711,N_15003,N_17706);
and U18712 (N_18712,N_15537,N_15594);
xor U18713 (N_18713,N_16574,N_15540);
nor U18714 (N_18714,N_17019,N_15880);
nor U18715 (N_18715,N_17924,N_16375);
and U18716 (N_18716,N_15413,N_17400);
or U18717 (N_18717,N_17490,N_17829);
and U18718 (N_18718,N_17212,N_17161);
nor U18719 (N_18719,N_17228,N_17761);
and U18720 (N_18720,N_16848,N_16111);
nand U18721 (N_18721,N_16911,N_15227);
xor U18722 (N_18722,N_15097,N_17558);
or U18723 (N_18723,N_16908,N_16697);
nor U18724 (N_18724,N_17535,N_16525);
or U18725 (N_18725,N_15378,N_16638);
nand U18726 (N_18726,N_17861,N_15660);
nor U18727 (N_18727,N_17079,N_15176);
xnor U18728 (N_18728,N_17518,N_15328);
or U18729 (N_18729,N_16570,N_15475);
nand U18730 (N_18730,N_16428,N_17229);
nand U18731 (N_18731,N_16986,N_17108);
nand U18732 (N_18732,N_17943,N_15577);
nor U18733 (N_18733,N_15345,N_16553);
and U18734 (N_18734,N_17095,N_16463);
nor U18735 (N_18735,N_16968,N_15521);
and U18736 (N_18736,N_17346,N_17086);
nand U18737 (N_18737,N_16773,N_15579);
nand U18738 (N_18738,N_17330,N_15115);
xnor U18739 (N_18739,N_17305,N_17078);
or U18740 (N_18740,N_17429,N_15722);
nor U18741 (N_18741,N_15506,N_17209);
xor U18742 (N_18742,N_15240,N_16755);
xor U18743 (N_18743,N_16727,N_16156);
nor U18744 (N_18744,N_16332,N_17029);
nor U18745 (N_18745,N_16788,N_15236);
nand U18746 (N_18746,N_17510,N_17345);
nor U18747 (N_18747,N_17426,N_15534);
nand U18748 (N_18748,N_15519,N_16639);
nand U18749 (N_18749,N_15766,N_15906);
nand U18750 (N_18750,N_17218,N_15992);
or U18751 (N_18751,N_15612,N_17302);
xor U18752 (N_18752,N_16953,N_15646);
nor U18753 (N_18753,N_16321,N_17557);
nor U18754 (N_18754,N_16302,N_17744);
xor U18755 (N_18755,N_17976,N_15318);
nand U18756 (N_18756,N_16101,N_17398);
nand U18757 (N_18757,N_17197,N_17742);
and U18758 (N_18758,N_16990,N_16562);
nor U18759 (N_18759,N_15425,N_15896);
xor U18760 (N_18760,N_15603,N_15431);
or U18761 (N_18761,N_15888,N_17309);
nor U18762 (N_18762,N_16281,N_17991);
or U18763 (N_18763,N_16391,N_16308);
or U18764 (N_18764,N_15587,N_15598);
and U18765 (N_18765,N_15192,N_17452);
nand U18766 (N_18766,N_16951,N_16097);
nand U18767 (N_18767,N_16148,N_15617);
nor U18768 (N_18768,N_15195,N_16787);
or U18769 (N_18769,N_16220,N_17196);
nor U18770 (N_18770,N_15919,N_16750);
and U18771 (N_18771,N_16393,N_15119);
nand U18772 (N_18772,N_15222,N_16770);
xnor U18773 (N_18773,N_16477,N_15373);
nand U18774 (N_18774,N_16732,N_17477);
nand U18775 (N_18775,N_17217,N_17506);
xor U18776 (N_18776,N_16885,N_16860);
nor U18777 (N_18777,N_17562,N_17610);
and U18778 (N_18778,N_17599,N_17298);
nor U18779 (N_18779,N_15675,N_15565);
and U18780 (N_18780,N_17194,N_16345);
or U18781 (N_18781,N_15950,N_15077);
or U18782 (N_18782,N_15979,N_17064);
and U18783 (N_18783,N_15745,N_15168);
and U18784 (N_18784,N_17152,N_17740);
nand U18785 (N_18785,N_16646,N_15681);
nor U18786 (N_18786,N_16947,N_15498);
or U18787 (N_18787,N_15323,N_16020);
or U18788 (N_18788,N_17077,N_15592);
nand U18789 (N_18789,N_16854,N_15650);
nor U18790 (N_18790,N_16279,N_17693);
or U18791 (N_18791,N_15755,N_16278);
nor U18792 (N_18792,N_16092,N_17005);
nand U18793 (N_18793,N_15854,N_16969);
nor U18794 (N_18794,N_17505,N_16730);
nor U18795 (N_18795,N_16785,N_15024);
nor U18796 (N_18796,N_17406,N_15299);
xor U18797 (N_18797,N_15623,N_17573);
or U18798 (N_18798,N_17201,N_15639);
or U18799 (N_18799,N_15051,N_16505);
or U18800 (N_18800,N_15706,N_17478);
nor U18801 (N_18801,N_16868,N_15834);
or U18802 (N_18802,N_15927,N_16157);
nor U18803 (N_18803,N_16214,N_15052);
nor U18804 (N_18804,N_17561,N_15987);
or U18805 (N_18805,N_17268,N_15369);
nor U18806 (N_18806,N_16751,N_17781);
or U18807 (N_18807,N_17968,N_17726);
and U18808 (N_18808,N_15276,N_16180);
and U18809 (N_18809,N_17724,N_17258);
nor U18810 (N_18810,N_15242,N_16767);
nor U18811 (N_18811,N_16021,N_17269);
xor U18812 (N_18812,N_17642,N_17383);
or U18813 (N_18813,N_16630,N_17634);
xor U18814 (N_18814,N_15578,N_15360);
or U18815 (N_18815,N_15912,N_15279);
xnor U18816 (N_18816,N_17977,N_16715);
nor U18817 (N_18817,N_15018,N_16055);
nand U18818 (N_18818,N_16205,N_16584);
xor U18819 (N_18819,N_16652,N_16149);
and U18820 (N_18820,N_17586,N_17798);
and U18821 (N_18821,N_16789,N_17614);
nor U18822 (N_18822,N_15913,N_16886);
xnor U18823 (N_18823,N_15881,N_16374);
or U18824 (N_18824,N_16402,N_17118);
nand U18825 (N_18825,N_15876,N_15769);
xor U18826 (N_18826,N_17471,N_17474);
nand U18827 (N_18827,N_16159,N_15494);
nand U18828 (N_18828,N_17923,N_16130);
and U18829 (N_18829,N_16931,N_15756);
nor U18830 (N_18830,N_15333,N_15549);
nor U18831 (N_18831,N_15664,N_16445);
and U18832 (N_18832,N_15079,N_16545);
or U18833 (N_18833,N_15277,N_15804);
or U18834 (N_18834,N_17938,N_16700);
nor U18835 (N_18835,N_17890,N_15488);
or U18836 (N_18836,N_17699,N_16596);
and U18837 (N_18837,N_17320,N_15423);
and U18838 (N_18838,N_15470,N_15151);
xnor U18839 (N_18839,N_17834,N_17540);
nor U18840 (N_18840,N_17354,N_15933);
or U18841 (N_18841,N_16979,N_15252);
xor U18842 (N_18842,N_15027,N_15914);
xnor U18843 (N_18843,N_15796,N_15193);
nor U18844 (N_18844,N_17122,N_17685);
or U18845 (N_18845,N_17823,N_17575);
nor U18846 (N_18846,N_15344,N_17641);
or U18847 (N_18847,N_16543,N_17667);
xnor U18848 (N_18848,N_15951,N_16315);
and U18849 (N_18849,N_16154,N_17210);
nand U18850 (N_18850,N_16507,N_15781);
and U18851 (N_18851,N_16858,N_16683);
or U18852 (N_18852,N_17020,N_15852);
xnor U18853 (N_18853,N_16248,N_17529);
xor U18854 (N_18854,N_15814,N_15321);
xor U18855 (N_18855,N_17439,N_17240);
and U18856 (N_18856,N_17611,N_16317);
and U18857 (N_18857,N_16657,N_17030);
xnor U18858 (N_18858,N_17498,N_15653);
or U18859 (N_18859,N_17731,N_15090);
nand U18860 (N_18860,N_15434,N_17504);
nand U18861 (N_18861,N_16334,N_15887);
nor U18862 (N_18862,N_15464,N_16044);
nand U18863 (N_18863,N_15263,N_15901);
nand U18864 (N_18864,N_15428,N_15391);
nor U18865 (N_18865,N_16483,N_16231);
xnor U18866 (N_18866,N_16434,N_16288);
nand U18867 (N_18867,N_16086,N_15555);
nor U18868 (N_18868,N_15315,N_17577);
nand U18869 (N_18869,N_17470,N_17536);
or U18870 (N_18870,N_16647,N_17300);
nor U18871 (N_18871,N_15260,N_16039);
nor U18872 (N_18872,N_16999,N_17713);
nand U18873 (N_18873,N_16344,N_16702);
and U18874 (N_18874,N_17453,N_16740);
nor U18875 (N_18875,N_17206,N_17009);
and U18876 (N_18876,N_16809,N_17182);
nor U18877 (N_18877,N_17241,N_15698);
nor U18878 (N_18878,N_15291,N_15208);
nand U18879 (N_18879,N_15161,N_15744);
nor U18880 (N_18880,N_17485,N_16563);
or U18881 (N_18881,N_16945,N_16330);
and U18882 (N_18882,N_15947,N_15791);
xnor U18883 (N_18883,N_15040,N_17013);
and U18884 (N_18884,N_16232,N_15430);
or U18885 (N_18885,N_16996,N_17450);
or U18886 (N_18886,N_16600,N_15581);
nor U18887 (N_18887,N_16576,N_16800);
nor U18888 (N_18888,N_17325,N_16895);
nor U18889 (N_18889,N_16984,N_17052);
and U18890 (N_18890,N_17671,N_17062);
nand U18891 (N_18891,N_17441,N_17590);
and U18892 (N_18892,N_15202,N_16423);
and U18893 (N_18893,N_15325,N_17572);
nor U18894 (N_18894,N_16748,N_17176);
nor U18895 (N_18895,N_16079,N_17679);
or U18896 (N_18896,N_16100,N_15347);
nor U18897 (N_18897,N_17120,N_17277);
xor U18898 (N_18898,N_16422,N_17362);
nor U18899 (N_18899,N_17852,N_17318);
or U18900 (N_18900,N_15788,N_17067);
and U18901 (N_18901,N_15717,N_17932);
and U18902 (N_18902,N_17979,N_17042);
nand U18903 (N_18903,N_17865,N_16689);
nor U18904 (N_18904,N_17316,N_17247);
xor U18905 (N_18905,N_16050,N_17253);
and U18906 (N_18906,N_15108,N_17278);
nor U18907 (N_18907,N_16464,N_16929);
xnor U18908 (N_18908,N_15563,N_17126);
and U18909 (N_18909,N_15967,N_15397);
or U18910 (N_18910,N_15777,N_15864);
or U18911 (N_18911,N_15982,N_15359);
xnor U18912 (N_18912,N_15070,N_17012);
or U18913 (N_18913,N_17710,N_17284);
nor U18914 (N_18914,N_16307,N_16236);
xnor U18915 (N_18915,N_17583,N_17788);
and U18916 (N_18916,N_17357,N_15733);
xnor U18917 (N_18917,N_15721,N_16245);
nor U18918 (N_18918,N_17854,N_17545);
nor U18919 (N_18919,N_15939,N_17980);
xor U18920 (N_18920,N_16935,N_16091);
nand U18921 (N_18921,N_16794,N_16946);
nor U18922 (N_18922,N_16709,N_17886);
nand U18923 (N_18923,N_17519,N_16662);
nand U18924 (N_18924,N_16167,N_15942);
nand U18925 (N_18925,N_15941,N_15916);
or U18926 (N_18926,N_17581,N_16564);
xor U18927 (N_18927,N_17967,N_17663);
or U18928 (N_18928,N_17917,N_15571);
nand U18929 (N_18929,N_17737,N_16093);
or U18930 (N_18930,N_17359,N_15019);
nand U18931 (N_18931,N_16579,N_16163);
xnor U18932 (N_18932,N_15406,N_16714);
or U18933 (N_18933,N_17859,N_17046);
and U18934 (N_18934,N_16444,N_15908);
or U18935 (N_18935,N_17417,N_16840);
or U18936 (N_18936,N_16005,N_15701);
or U18937 (N_18937,N_16552,N_17630);
and U18938 (N_18938,N_16912,N_15742);
nand U18939 (N_18939,N_17858,N_16614);
nand U18940 (N_18940,N_17665,N_16776);
nand U18941 (N_18941,N_15125,N_16837);
and U18942 (N_18942,N_16654,N_17570);
xnor U18943 (N_18943,N_15813,N_17083);
or U18944 (N_18944,N_17369,N_16069);
nor U18945 (N_18945,N_16756,N_16673);
or U18946 (N_18946,N_17935,N_16090);
or U18947 (N_18947,N_17347,N_17011);
nor U18948 (N_18948,N_15269,N_15708);
and U18949 (N_18949,N_16303,N_15329);
nand U18950 (N_18950,N_17204,N_16348);
nor U18951 (N_18951,N_15981,N_16435);
xnor U18952 (N_18952,N_15272,N_16019);
or U18953 (N_18953,N_16120,N_16489);
nand U18954 (N_18954,N_17723,N_15041);
or U18955 (N_18955,N_15843,N_15152);
nor U18956 (N_18956,N_16040,N_16199);
nand U18957 (N_18957,N_17851,N_15064);
or U18958 (N_18958,N_17674,N_17419);
nand U18959 (N_18959,N_16838,N_17645);
nor U18960 (N_18960,N_17907,N_17438);
and U18961 (N_18961,N_16342,N_17800);
xnor U18962 (N_18962,N_16831,N_15714);
nor U18963 (N_18963,N_17136,N_15102);
and U18964 (N_18964,N_15080,N_15004);
xnor U18965 (N_18965,N_16385,N_17822);
or U18966 (N_18966,N_16140,N_16546);
and U18967 (N_18967,N_15611,N_16046);
and U18968 (N_18968,N_17627,N_16200);
nor U18969 (N_18969,N_17869,N_15911);
xnor U18970 (N_18970,N_16766,N_17843);
nand U18971 (N_18971,N_17107,N_16798);
nor U18972 (N_18972,N_17380,N_17752);
or U18973 (N_18973,N_15905,N_17715);
or U18974 (N_18974,N_15186,N_16548);
nor U18975 (N_18975,N_15402,N_17393);
and U18976 (N_18976,N_15670,N_16611);
nand U18977 (N_18977,N_15042,N_17435);
or U18978 (N_18978,N_16028,N_17043);
nand U18979 (N_18979,N_16834,N_17845);
nor U18980 (N_18980,N_17690,N_16501);
or U18981 (N_18981,N_16451,N_16062);
xnor U18982 (N_18982,N_15414,N_17402);
or U18983 (N_18983,N_15595,N_15216);
and U18984 (N_18984,N_16237,N_15103);
or U18985 (N_18985,N_17893,N_17639);
or U18986 (N_18986,N_15225,N_16472);
nand U18987 (N_18987,N_17554,N_15381);
xor U18988 (N_18988,N_15223,N_17533);
or U18989 (N_18989,N_17664,N_17033);
and U18990 (N_18990,N_17998,N_16913);
and U18991 (N_18991,N_17941,N_16217);
nor U18992 (N_18992,N_15085,N_15394);
and U18993 (N_18993,N_16126,N_16284);
xor U18994 (N_18994,N_16554,N_17195);
xnor U18995 (N_18995,N_16610,N_15530);
xnor U18996 (N_18996,N_15922,N_15713);
nor U18997 (N_18997,N_15179,N_15638);
xnor U18998 (N_18998,N_15586,N_16493);
nand U18999 (N_18999,N_16139,N_15576);
and U19000 (N_19000,N_16320,N_16778);
and U19001 (N_19001,N_16949,N_16706);
or U19002 (N_19002,N_16503,N_17319);
xnor U19003 (N_19003,N_17041,N_15545);
nor U19004 (N_19004,N_16747,N_17653);
and U19005 (N_19005,N_17900,N_17729);
and U19006 (N_19006,N_15690,N_16273);
nor U19007 (N_19007,N_16064,N_17137);
nor U19008 (N_19008,N_16414,N_16651);
nor U19009 (N_19009,N_17016,N_17616);
nor U19010 (N_19010,N_16583,N_15973);
nand U19011 (N_19011,N_16899,N_16833);
nor U19012 (N_19012,N_15343,N_16643);
xnor U19013 (N_19013,N_15355,N_16593);
nor U19014 (N_19014,N_17321,N_16534);
nand U19015 (N_19015,N_16544,N_17920);
or U19016 (N_19016,N_16306,N_17969);
xnor U19017 (N_19017,N_16786,N_17888);
and U19018 (N_19018,N_16887,N_15099);
nand U19019 (N_19019,N_15069,N_16636);
and U19020 (N_19020,N_17444,N_15288);
or U19021 (N_19021,N_16606,N_17863);
nand U19022 (N_19022,N_15985,N_16676);
or U19023 (N_19023,N_16500,N_16804);
xor U19024 (N_19024,N_16270,N_17082);
or U19025 (N_19025,N_17036,N_17613);
and U19026 (N_19026,N_15661,N_17035);
and U19027 (N_19027,N_17205,N_16271);
nor U19028 (N_19028,N_15365,N_15072);
nand U19029 (N_19029,N_15636,N_17844);
or U19030 (N_19030,N_17615,N_15124);
nor U19031 (N_19031,N_17921,N_15029);
nand U19032 (N_19032,N_16378,N_17098);
nor U19033 (N_19033,N_17722,N_16144);
nand U19034 (N_19034,N_15021,N_16121);
or U19035 (N_19035,N_15314,N_17508);
xor U19036 (N_19036,N_16717,N_16735);
xnor U19037 (N_19037,N_15557,N_15665);
xnor U19038 (N_19038,N_16259,N_17912);
nor U19039 (N_19039,N_16354,N_15348);
or U19040 (N_19040,N_16155,N_16491);
nand U19041 (N_19041,N_15142,N_15148);
nand U19042 (N_19042,N_15515,N_16826);
xnor U19043 (N_19043,N_16299,N_15187);
or U19044 (N_19044,N_15060,N_16527);
nand U19045 (N_19045,N_16314,N_15632);
or U19046 (N_19046,N_15759,N_16888);
xnor U19047 (N_19047,N_17652,N_15198);
nand U19048 (N_19048,N_16153,N_15605);
or U19049 (N_19049,N_16842,N_16108);
xnor U19050 (N_19050,N_15405,N_17816);
nand U19051 (N_19051,N_15454,N_16103);
xnor U19052 (N_19052,N_17786,N_16311);
and U19053 (N_19053,N_17700,N_15970);
or U19054 (N_19054,N_17449,N_17709);
and U19055 (N_19055,N_16215,N_17623);
xnor U19056 (N_19056,N_17848,N_17101);
and U19057 (N_19057,N_17301,N_17970);
nand U19058 (N_19058,N_16998,N_17017);
nand U19059 (N_19059,N_16890,N_15219);
and U19060 (N_19060,N_17716,N_17324);
nor U19061 (N_19061,N_17782,N_15954);
nand U19062 (N_19062,N_17332,N_15093);
or U19063 (N_19063,N_17025,N_15289);
and U19064 (N_19064,N_16029,N_17294);
nor U19065 (N_19065,N_17049,N_15259);
and U19066 (N_19066,N_17334,N_17832);
or U19067 (N_19067,N_15891,N_16295);
nand U19068 (N_19068,N_17632,N_16460);
nor U19069 (N_19069,N_17243,N_15132);
xnor U19070 (N_19070,N_15199,N_17287);
and U19071 (N_19071,N_16925,N_15989);
nor U19072 (N_19072,N_16486,N_16889);
or U19073 (N_19073,N_15495,N_17024);
xor U19074 (N_19074,N_15667,N_17186);
nand U19075 (N_19075,N_17288,N_17328);
or U19076 (N_19076,N_16339,N_16171);
and U19077 (N_19077,N_15358,N_16329);
xnor U19078 (N_19078,N_17669,N_17129);
nand U19079 (N_19079,N_17552,N_16753);
or U19080 (N_19080,N_16002,N_16812);
nor U19081 (N_19081,N_17238,N_17428);
nor U19082 (N_19082,N_17950,N_17666);
and U19083 (N_19083,N_16203,N_16117);
xnor U19084 (N_19084,N_15137,N_15320);
or U19085 (N_19085,N_17801,N_16870);
nor U19086 (N_19086,N_15898,N_15597);
xor U19087 (N_19087,N_15860,N_16150);
nand U19088 (N_19088,N_15290,N_17589);
and U19089 (N_19089,N_16371,N_17088);
or U19090 (N_19090,N_16000,N_15771);
nand U19091 (N_19091,N_16129,N_15790);
and U19092 (N_19092,N_16882,N_16210);
nand U19093 (N_19093,N_16222,N_17338);
nand U19094 (N_19094,N_16879,N_17981);
and U19095 (N_19095,N_15039,N_17654);
nand U19096 (N_19096,N_15268,N_16123);
or U19097 (N_19097,N_16096,N_17987);
and U19098 (N_19098,N_15234,N_15339);
nor U19099 (N_19099,N_17621,N_16397);
nand U19100 (N_19100,N_15238,N_16955);
and U19101 (N_19101,N_15379,N_17109);
nand U19102 (N_19102,N_17707,N_15710);
or U19103 (N_19103,N_15847,N_16192);
and U19104 (N_19104,N_16558,N_15050);
or U19105 (N_19105,N_16316,N_15527);
nand U19106 (N_19106,N_15485,N_15893);
and U19107 (N_19107,N_16048,N_15895);
nor U19108 (N_19108,N_17612,N_15782);
xor U19109 (N_19109,N_16869,N_17045);
nand U19110 (N_19110,N_15022,N_17080);
nand U19111 (N_19111,N_16572,N_15118);
nor U19112 (N_19112,N_17591,N_17382);
nor U19113 (N_19113,N_17198,N_15009);
xnor U19114 (N_19114,N_15705,N_17177);
nor U19115 (N_19115,N_16954,N_15704);
nand U19116 (N_19116,N_17618,N_16146);
or U19117 (N_19117,N_16620,N_16300);
nand U19118 (N_19118,N_16289,N_16663);
xor U19119 (N_19119,N_17574,N_15112);
nor U19120 (N_19120,N_17189,N_15251);
nor U19121 (N_19121,N_15570,N_15684);
or U19122 (N_19122,N_16471,N_16310);
nand U19123 (N_19123,N_15319,N_17341);
or U19124 (N_19124,N_15030,N_17904);
and U19125 (N_19125,N_16061,N_16488);
xnor U19126 (N_19126,N_17032,N_16853);
nor U19127 (N_19127,N_16568,N_16198);
and U19128 (N_19128,N_16991,N_17906);
and U19129 (N_19129,N_17881,N_16168);
nor U19130 (N_19130,N_16034,N_17559);
and U19131 (N_19131,N_15693,N_17624);
xor U19132 (N_19132,N_15468,N_17773);
nand U19133 (N_19133,N_17556,N_15226);
xnor U19134 (N_19134,N_15270,N_15968);
nor U19135 (N_19135,N_16803,N_17104);
nor U19136 (N_19136,N_17468,N_17010);
nor U19137 (N_19137,N_16741,N_17368);
and U19138 (N_19138,N_16918,N_17996);
and U19139 (N_19139,N_15957,N_16075);
and U19140 (N_19140,N_17021,N_17831);
nand U19141 (N_19141,N_15648,N_16038);
nor U19142 (N_19142,N_17565,N_16589);
nand U19143 (N_19143,N_15483,N_17937);
or U19144 (N_19144,N_15547,N_15607);
nand U19145 (N_19145,N_17239,N_17550);
and U19146 (N_19146,N_15209,N_17608);
xor U19147 (N_19147,N_15243,N_15071);
and U19148 (N_19148,N_16540,N_16433);
or U19149 (N_19149,N_17972,N_17390);
nand U19150 (N_19150,N_15798,N_17944);
and U19151 (N_19151,N_17770,N_15466);
and U19152 (N_19152,N_15449,N_16049);
nand U19153 (N_19153,N_15764,N_16443);
nor U19154 (N_19154,N_16207,N_17458);
nor U19155 (N_19155,N_16874,N_16356);
and U19156 (N_19156,N_17909,N_16187);
xnor U19157 (N_19157,N_15938,N_15818);
nor U19158 (N_19158,N_15181,N_15550);
xnor U19159 (N_19159,N_15312,N_15390);
or U19160 (N_19160,N_17691,N_15081);
or U19161 (N_19161,N_17159,N_15772);
xor U19162 (N_19162,N_17125,N_16679);
nand U19163 (N_19163,N_17090,N_16455);
xor U19164 (N_19164,N_15779,N_16294);
xnor U19165 (N_19165,N_15150,N_16290);
nand U19166 (N_19166,N_16938,N_17070);
nand U19167 (N_19167,N_15407,N_15999);
nand U19168 (N_19168,N_15026,N_17058);
nor U19169 (N_19169,N_16783,N_16053);
xor U19170 (N_19170,N_17718,N_16172);
and U19171 (N_19171,N_17787,N_16372);
nor U19172 (N_19172,N_15332,N_16206);
nand U19173 (N_19173,N_17763,N_17530);
or U19174 (N_19174,N_17862,N_15127);
xor U19175 (N_19175,N_17803,N_16431);
or U19176 (N_19176,N_15409,N_16956);
or U19177 (N_19177,N_17596,N_15531);
and U19178 (N_19178,N_15902,N_17802);
nor U19179 (N_19179,N_15401,N_16859);
nor U19180 (N_19180,N_17466,N_15677);
or U19181 (N_19181,N_17765,N_15558);
or U19182 (N_19182,N_17384,N_16824);
nand U19183 (N_19183,N_17933,N_15418);
nor U19184 (N_19184,N_17719,N_16411);
xnor U19185 (N_19185,N_16581,N_16669);
or U19186 (N_19186,N_16142,N_16965);
and U19187 (N_19187,N_17549,N_15926);
and U19188 (N_19188,N_17389,N_15776);
and U19189 (N_19189,N_17455,N_17351);
nor U19190 (N_19190,N_15978,N_16692);
or U19191 (N_19191,N_17350,N_17772);
and U19192 (N_19192,N_17523,N_17461);
nor U19193 (N_19193,N_16265,N_15517);
nor U19194 (N_19194,N_15068,N_16571);
and U19195 (N_19195,N_16240,N_16173);
nand U19196 (N_19196,N_17984,N_16301);
xor U19197 (N_19197,N_15878,N_16309);
and U19198 (N_19198,N_16351,N_15935);
xnor U19199 (N_19199,N_15894,N_16894);
nand U19200 (N_19200,N_16175,N_16337);
nor U19201 (N_19201,N_17014,N_16772);
nor U19202 (N_19202,N_17483,N_17500);
xnor U19203 (N_19203,N_16704,N_17056);
nor U19204 (N_19204,N_15993,N_16268);
xor U19205 (N_19205,N_17215,N_17312);
nor U19206 (N_19206,N_16208,N_15215);
nor U19207 (N_19207,N_16474,N_16536);
xor U19208 (N_19208,N_15424,N_17178);
and U19209 (N_19209,N_16006,N_16635);
xor U19210 (N_19210,N_15928,N_15463);
nor U19211 (N_19211,N_15604,N_15267);
or U19212 (N_19212,N_15048,N_16482);
xnor U19213 (N_19213,N_17348,N_17174);
and U19214 (N_19214,N_15037,N_16973);
nand U19215 (N_19215,N_17945,N_16814);
and U19216 (N_19216,N_17068,N_16115);
nor U19217 (N_19217,N_17234,N_15067);
or U19218 (N_19218,N_16531,N_17360);
nor U19219 (N_19219,N_15541,N_15614);
and U19220 (N_19220,N_15376,N_15767);
and U19221 (N_19221,N_17442,N_15163);
or U19222 (N_19222,N_17918,N_15751);
nand U19223 (N_19223,N_17884,N_17115);
and U19224 (N_19224,N_16806,N_16528);
or U19225 (N_19225,N_15383,N_16213);
or U19226 (N_19226,N_15078,N_17775);
xor U19227 (N_19227,N_17527,N_16731);
or U19228 (N_19228,N_16272,N_16327);
nand U19229 (N_19229,N_17342,N_17395);
and U19230 (N_19230,N_17479,N_16815);
and U19231 (N_19231,N_16519,N_16335);
and U19232 (N_19232,N_16230,N_16184);
or U19233 (N_19233,N_17183,N_17774);
and U19234 (N_19234,N_16701,N_17259);
nor U19235 (N_19235,N_17656,N_17841);
xnor U19236 (N_19236,N_16253,N_16506);
nand U19237 (N_19237,N_16084,N_16659);
nand U19238 (N_19238,N_16634,N_15275);
or U19239 (N_19239,N_15953,N_17684);
nand U19240 (N_19240,N_17180,N_15087);
nand U19241 (N_19241,N_16266,N_17808);
xnor U19242 (N_19242,N_17910,N_16293);
or U19243 (N_19243,N_15262,N_16514);
and U19244 (N_19244,N_17648,N_17883);
or U19245 (N_19245,N_15038,N_16367);
xor U19246 (N_19246,N_17004,N_15188);
and U19247 (N_19247,N_16857,N_16441);
and U19248 (N_19248,N_17875,N_16410);
or U19249 (N_19249,N_16024,N_16007);
and U19250 (N_19250,N_15055,N_16790);
xnor U19251 (N_19251,N_17355,N_15976);
nand U19252 (N_19252,N_17560,N_17828);
xor U19253 (N_19253,N_16675,N_17031);
nor U19254 (N_19254,N_15862,N_17039);
or U19255 (N_19255,N_16677,N_16904);
nand U19256 (N_19256,N_15295,N_17687);
xor U19257 (N_19257,N_16729,N_17515);
nand U19258 (N_19258,N_15503,N_17491);
or U19259 (N_19259,N_15863,N_15493);
xor U19260 (N_19260,N_17856,N_15875);
nand U19261 (N_19261,N_16413,N_15879);
and U19262 (N_19262,N_15625,N_17759);
nor U19263 (N_19263,N_15139,N_16580);
xnor U19264 (N_19264,N_15306,N_15831);
or U19265 (N_19265,N_17678,N_17677);
nor U19266 (N_19266,N_16573,N_16135);
xor U19267 (N_19267,N_17272,N_16871);
xnor U19268 (N_19268,N_15750,N_17007);
nor U19269 (N_19269,N_15601,N_16291);
xor U19270 (N_19270,N_17403,N_16105);
nor U19271 (N_19271,N_17837,N_17779);
or U19272 (N_19272,N_16720,N_17001);
xnor U19273 (N_19273,N_16296,N_16967);
or U19274 (N_19274,N_16591,N_15082);
nand U19275 (N_19275,N_17683,N_15844);
and U19276 (N_19276,N_16439,N_17467);
nand U19277 (N_19277,N_15170,N_16137);
nand U19278 (N_19278,N_15145,N_17806);
or U19279 (N_19279,N_16884,N_15155);
and U19280 (N_19280,N_15146,N_15467);
and U19281 (N_19281,N_16406,N_16244);
or U19282 (N_19282,N_15568,N_15326);
and U19283 (N_19283,N_16042,N_17797);
nor U19284 (N_19284,N_15297,N_17219);
or U19285 (N_19285,N_15300,N_17955);
or U19286 (N_19286,N_17448,N_16582);
nand U19287 (N_19287,N_16909,N_17099);
and U19288 (N_19288,N_15619,N_15738);
and U19289 (N_19289,N_16328,N_17481);
or U19290 (N_19290,N_17661,N_16937);
nor U19291 (N_19291,N_16526,N_15868);
xor U19292 (N_19292,N_15761,N_15000);
nor U19293 (N_19293,N_17633,N_15280);
nand U19294 (N_19294,N_15058,N_17387);
nor U19295 (N_19295,N_16626,N_16989);
nand U19296 (N_19296,N_15410,N_15281);
nor U19297 (N_19297,N_16151,N_16001);
and U19298 (N_19298,N_17496,N_16036);
xnor U19299 (N_19299,N_17293,N_15086);
nor U19300 (N_19300,N_15512,N_17221);
or U19301 (N_19301,N_16542,N_15509);
nor U19302 (N_19302,N_17638,N_16910);
xnor U19303 (N_19303,N_15889,N_17643);
and U19304 (N_19304,N_16480,N_16603);
or U19305 (N_19305,N_16658,N_15548);
xor U19306 (N_19306,N_15897,N_16379);
or U19307 (N_19307,N_16189,N_16333);
nor U19308 (N_19308,N_17267,N_17745);
nor U19309 (N_19309,N_15699,N_17528);
xor U19310 (N_19310,N_15904,N_15789);
nor U19311 (N_19311,N_16183,N_17245);
xnor U19312 (N_19312,N_17296,N_15249);
xnor U19313 (N_19313,N_15884,N_15309);
or U19314 (N_19314,N_16933,N_15056);
and U19315 (N_19315,N_16901,N_15175);
nand U19316 (N_19316,N_16074,N_16943);
xnor U19317 (N_19317,N_17394,N_16457);
nand U19318 (N_19318,N_16775,N_15191);
nor U19319 (N_19319,N_16234,N_15341);
nand U19320 (N_19320,N_16400,N_17314);
nor U19321 (N_19321,N_15292,N_17000);
nor U19322 (N_19322,N_15741,N_17532);
nand U19323 (N_19323,N_16037,N_16642);
xnor U19324 (N_19324,N_17401,N_17887);
nand U19325 (N_19325,N_17167,N_16107);
xor U19326 (N_19326,N_15356,N_15624);
and U19327 (N_19327,N_17423,N_15588);
nor U19328 (N_19328,N_17827,N_17810);
nor U19329 (N_19329,N_15736,N_16928);
xnor U19330 (N_19330,N_16119,N_15239);
nor U19331 (N_19331,N_16113,N_15673);
xnor U19332 (N_19332,N_17812,N_15416);
xor U19333 (N_19333,N_16923,N_15211);
xnor U19334 (N_19334,N_15841,N_16588);
or U19335 (N_19335,N_16686,N_15114);
nor U19336 (N_19336,N_16983,N_15523);
nand U19337 (N_19337,N_16066,N_15235);
or U19338 (N_19338,N_17132,N_15182);
or U19339 (N_19339,N_15159,N_16716);
nand U19340 (N_19340,N_16275,N_16305);
xor U19341 (N_19341,N_17978,N_17619);
nor U19342 (N_19342,N_17817,N_15020);
nand U19343 (N_19343,N_16347,N_16844);
and U19344 (N_19344,N_15622,N_16346);
or U19345 (N_19345,N_17291,N_17281);
xor U19346 (N_19346,N_17060,N_17372);
xnor U19347 (N_19347,N_16228,N_16179);
nand U19348 (N_19348,N_15230,N_17670);
or U19349 (N_19349,N_17901,N_17306);
nor U19350 (N_19350,N_16058,N_16110);
xnor U19351 (N_19351,N_16817,N_15088);
xor U19352 (N_19352,N_17660,N_17704);
and U19353 (N_19353,N_17433,N_15116);
nand U19354 (N_19354,N_17339,N_16152);
and U19355 (N_19355,N_17548,N_17879);
nor U19356 (N_19356,N_17676,N_15023);
nor U19357 (N_19357,N_17749,N_17169);
nor U19358 (N_19358,N_16341,N_16440);
nand U19359 (N_19359,N_16627,N_15371);
or U19360 (N_19360,N_15662,N_15264);
nand U19361 (N_19361,N_15302,N_17544);
nand U19362 (N_19362,N_15828,N_17672);
nand U19363 (N_19363,N_16469,N_16465);
xnor U19364 (N_19364,N_17375,N_17358);
and U19365 (N_19365,N_17208,N_17385);
nand U19366 (N_19366,N_15892,N_16219);
nand U19367 (N_19367,N_15514,N_15983);
and U19368 (N_19368,N_16023,N_17873);
nand U19369 (N_19369,N_17988,N_15707);
and U19370 (N_19370,N_15149,N_17815);
xor U19371 (N_19371,N_16188,N_17447);
and U19372 (N_19372,N_17553,N_17261);
xnor U19373 (N_19373,N_15131,N_15446);
nor U19374 (N_19374,N_15929,N_17093);
nor U19375 (N_19375,N_15944,N_15387);
or U19376 (N_19376,N_16687,N_17593);
nor U19377 (N_19377,N_15362,N_15184);
xor U19378 (N_19378,N_15773,N_16892);
and U19379 (N_19379,N_15724,N_16481);
xnor U19380 (N_19380,N_16014,N_17437);
nand U19381 (N_19381,N_16461,N_17768);
nand U19382 (N_19382,N_17867,N_16622);
nor U19383 (N_19383,N_17963,N_16987);
and U19384 (N_19384,N_17273,N_15157);
nor U19385 (N_19385,N_17489,N_16900);
nor U19386 (N_19386,N_15244,N_15171);
or U19387 (N_19387,N_16743,N_15809);
nor U19388 (N_19388,N_16178,N_15457);
xnor U19389 (N_19389,N_16260,N_16621);
nor U19390 (N_19390,N_15156,N_15946);
nand U19391 (N_19391,N_15296,N_16408);
nor U19392 (N_19392,N_17427,N_15775);
nor U19393 (N_19393,N_16602,N_16404);
nor U19394 (N_19394,N_15185,N_17546);
nand U19395 (N_19395,N_16233,N_15909);
or U19396 (N_19396,N_17882,N_17124);
nand U19397 (N_19397,N_17006,N_16068);
xnor U19398 (N_19398,N_15033,N_17872);
or U19399 (N_19399,N_17804,N_15210);
and U19400 (N_19400,N_15984,N_15221);
xnor U19401 (N_19401,N_17993,N_15584);
or U19402 (N_19402,N_17111,N_17087);
nor U19403 (N_19403,N_16618,N_16085);
nand U19404 (N_19404,N_17200,N_17193);
nor U19405 (N_19405,N_15735,N_17795);
xor U19406 (N_19406,N_16362,N_16030);
nand U19407 (N_19407,N_15734,N_17323);
nor U19408 (N_19408,N_16109,N_17069);
nor U19409 (N_19409,N_16681,N_16364);
xor U19410 (N_19410,N_15224,N_15501);
nor U19411 (N_19411,N_17994,N_15700);
and U19412 (N_19412,N_15686,N_16530);
xnor U19413 (N_19413,N_15671,N_17758);
nand U19414 (N_19414,N_16262,N_17138);
nor U19415 (N_19415,N_17628,N_15564);
or U19416 (N_19416,N_15076,N_15016);
nor U19417 (N_19417,N_16592,N_17807);
and U19418 (N_19418,N_15154,N_15237);
or U19419 (N_19419,N_17335,N_17164);
xor U19420 (N_19420,N_16241,N_17418);
and U19421 (N_19421,N_15505,N_15107);
nand U19422 (N_19422,N_15372,N_15709);
and U19423 (N_19423,N_16802,N_17023);
nand U19424 (N_19424,N_15931,N_17962);
nand U19425 (N_19425,N_17813,N_15438);
nor U19426 (N_19426,N_17588,N_17097);
and U19427 (N_19427,N_17399,N_16768);
or U19428 (N_19428,N_15573,N_17792);
nor U19429 (N_19429,N_16674,N_15808);
xor U19430 (N_19430,N_15806,N_15143);
and U19431 (N_19431,N_17696,N_16797);
or U19432 (N_19432,N_16497,N_17370);
and U19433 (N_19433,N_16535,N_15460);
or U19434 (N_19434,N_15575,N_15723);
and U19435 (N_19435,N_15691,N_17965);
nand U19436 (N_19436,N_17655,N_15492);
nand U19437 (N_19437,N_15566,N_17694);
nand U19438 (N_19438,N_17754,N_15842);
or U19439 (N_19439,N_17524,N_16088);
xor U19440 (N_19440,N_16670,N_17534);
and U19441 (N_19441,N_17789,N_15462);
nor U19442 (N_19442,N_15284,N_16011);
and U19443 (N_19443,N_15797,N_16401);
nor U19444 (N_19444,N_15948,N_16239);
and U19445 (N_19445,N_17153,N_16209);
or U19446 (N_19446,N_16365,N_15294);
xnor U19447 (N_19447,N_16359,N_17949);
and U19448 (N_19448,N_17100,N_15609);
nor U19449 (N_19449,N_16098,N_16338);
and U19450 (N_19450,N_16633,N_17425);
nand U19451 (N_19451,N_17682,N_16409);
xnor U19452 (N_19452,N_17220,N_17727);
and U19453 (N_19453,N_17738,N_16502);
xnor U19454 (N_19454,N_15873,N_15006);
nand U19455 (N_19455,N_17264,N_17814);
nand U19456 (N_19456,N_15335,N_16087);
nand U19457 (N_19457,N_17203,N_15918);
or U19458 (N_19458,N_17018,N_17110);
or U19459 (N_19459,N_15524,N_17868);
xnor U19460 (N_19460,N_17472,N_17516);
or U19461 (N_19461,N_15278,N_16924);
xnor U19462 (N_19462,N_16035,N_16628);
and U19463 (N_19463,N_16744,N_16429);
or U19464 (N_19464,N_17059,N_15719);
xor U19465 (N_19465,N_15652,N_17733);
and U19466 (N_19466,N_15445,N_17207);
and U19467 (N_19467,N_16388,N_17414);
xnor U19468 (N_19468,N_15837,N_15389);
nor U19469 (N_19469,N_15980,N_17130);
xnor U19470 (N_19470,N_15749,N_15593);
or U19471 (N_19471,N_17224,N_15177);
or U19472 (N_19472,N_15529,N_17521);
xor U19473 (N_19473,N_16022,N_15616);
xor U19474 (N_19474,N_17317,N_16326);
or U19475 (N_19475,N_17139,N_17171);
nand U19476 (N_19476,N_17785,N_16866);
or U19477 (N_19477,N_16993,N_17188);
xnor U19478 (N_19478,N_16276,N_17265);
or U19479 (N_19479,N_17721,N_15469);
nor U19480 (N_19480,N_16285,N_17026);
and U19481 (N_19481,N_17336,N_17495);
nor U19482 (N_19482,N_15730,N_15959);
xnor U19483 (N_19483,N_15374,N_16632);
xor U19484 (N_19484,N_16250,N_16771);
xor U19485 (N_19485,N_17734,N_17958);
or U19486 (N_19486,N_16830,N_16566);
xnor U19487 (N_19487,N_15444,N_15384);
nor U19488 (N_19488,N_16017,N_15479);
xor U19489 (N_19489,N_15342,N_15820);
or U19490 (N_19490,N_16846,N_17154);
nor U19491 (N_19491,N_15986,N_16043);
nand U19492 (N_19492,N_16648,N_16708);
nand U19493 (N_19493,N_15361,N_16808);
nor U19494 (N_19494,N_16380,N_15602);
or U19495 (N_19495,N_15028,N_17520);
nand U19496 (N_19496,N_17751,N_15075);
nor U19497 (N_19497,N_16875,N_15432);
nor U19498 (N_19498,N_17112,N_17456);
nor U19499 (N_19499,N_15174,N_16370);
and U19500 (N_19500,N_17959,N_15448);
nand U19501 (N_19501,N_15329,N_16489);
nor U19502 (N_19502,N_17224,N_15644);
nand U19503 (N_19503,N_15962,N_17467);
or U19504 (N_19504,N_16704,N_16748);
or U19505 (N_19505,N_15096,N_17967);
or U19506 (N_19506,N_17261,N_17240);
or U19507 (N_19507,N_16350,N_17573);
nand U19508 (N_19508,N_15626,N_15921);
and U19509 (N_19509,N_16143,N_17325);
xor U19510 (N_19510,N_15487,N_16330);
and U19511 (N_19511,N_17807,N_17974);
or U19512 (N_19512,N_15947,N_15570);
nand U19513 (N_19513,N_16574,N_15150);
nand U19514 (N_19514,N_15636,N_17451);
nand U19515 (N_19515,N_16782,N_15629);
nand U19516 (N_19516,N_17254,N_17913);
or U19517 (N_19517,N_15345,N_17001);
or U19518 (N_19518,N_17352,N_16593);
or U19519 (N_19519,N_16283,N_15023);
nand U19520 (N_19520,N_17161,N_17172);
nor U19521 (N_19521,N_16220,N_15403);
nor U19522 (N_19522,N_16272,N_15674);
and U19523 (N_19523,N_15733,N_15160);
or U19524 (N_19524,N_16336,N_16770);
or U19525 (N_19525,N_15298,N_17505);
nand U19526 (N_19526,N_16340,N_17949);
or U19527 (N_19527,N_15979,N_16512);
xnor U19528 (N_19528,N_16035,N_17591);
nand U19529 (N_19529,N_16963,N_15315);
nand U19530 (N_19530,N_16446,N_17967);
or U19531 (N_19531,N_15601,N_16770);
or U19532 (N_19532,N_17289,N_16077);
xnor U19533 (N_19533,N_16507,N_15800);
or U19534 (N_19534,N_17512,N_16498);
and U19535 (N_19535,N_16364,N_17717);
nand U19536 (N_19536,N_17911,N_17563);
xnor U19537 (N_19537,N_15925,N_16502);
and U19538 (N_19538,N_17773,N_15607);
nand U19539 (N_19539,N_16071,N_15698);
nor U19540 (N_19540,N_17828,N_15947);
nor U19541 (N_19541,N_17359,N_15560);
nand U19542 (N_19542,N_17726,N_15014);
and U19543 (N_19543,N_17778,N_16924);
and U19544 (N_19544,N_17790,N_17316);
nor U19545 (N_19545,N_16406,N_16721);
or U19546 (N_19546,N_16661,N_17983);
or U19547 (N_19547,N_15251,N_17127);
xor U19548 (N_19548,N_17764,N_15296);
and U19549 (N_19549,N_17040,N_17948);
xor U19550 (N_19550,N_15338,N_16043);
nor U19551 (N_19551,N_16263,N_16686);
xor U19552 (N_19552,N_16312,N_15546);
nor U19553 (N_19553,N_15048,N_16975);
and U19554 (N_19554,N_16571,N_17325);
and U19555 (N_19555,N_17425,N_16543);
or U19556 (N_19556,N_16312,N_16511);
nand U19557 (N_19557,N_16367,N_15231);
or U19558 (N_19558,N_16983,N_15895);
nor U19559 (N_19559,N_16822,N_15175);
nor U19560 (N_19560,N_15897,N_16573);
nand U19561 (N_19561,N_15189,N_16570);
or U19562 (N_19562,N_15773,N_15700);
and U19563 (N_19563,N_17241,N_17788);
nor U19564 (N_19564,N_15067,N_17616);
nor U19565 (N_19565,N_15880,N_16649);
and U19566 (N_19566,N_17377,N_15657);
nand U19567 (N_19567,N_16793,N_16287);
nand U19568 (N_19568,N_17935,N_15115);
nand U19569 (N_19569,N_17461,N_15595);
nand U19570 (N_19570,N_15592,N_16841);
nand U19571 (N_19571,N_16589,N_17933);
nor U19572 (N_19572,N_17145,N_17085);
xor U19573 (N_19573,N_17036,N_16405);
and U19574 (N_19574,N_16687,N_15507);
nand U19575 (N_19575,N_17659,N_15121);
nand U19576 (N_19576,N_16889,N_16607);
nand U19577 (N_19577,N_17333,N_17601);
xor U19578 (N_19578,N_15115,N_16785);
nor U19579 (N_19579,N_17599,N_16114);
xor U19580 (N_19580,N_17151,N_17206);
nor U19581 (N_19581,N_17573,N_15522);
nor U19582 (N_19582,N_16164,N_17374);
nand U19583 (N_19583,N_15093,N_16572);
or U19584 (N_19584,N_16466,N_16518);
xor U19585 (N_19585,N_16711,N_16775);
xnor U19586 (N_19586,N_17646,N_15631);
xnor U19587 (N_19587,N_17828,N_15016);
and U19588 (N_19588,N_16327,N_15856);
or U19589 (N_19589,N_15479,N_17305);
xor U19590 (N_19590,N_16432,N_15164);
or U19591 (N_19591,N_16698,N_16830);
xor U19592 (N_19592,N_16484,N_16446);
xnor U19593 (N_19593,N_15306,N_15135);
or U19594 (N_19594,N_15400,N_17667);
nor U19595 (N_19595,N_16136,N_16713);
nor U19596 (N_19596,N_16785,N_15599);
nand U19597 (N_19597,N_16025,N_16885);
xnor U19598 (N_19598,N_17339,N_17658);
nor U19599 (N_19599,N_15671,N_15403);
or U19600 (N_19600,N_17912,N_17833);
and U19601 (N_19601,N_16584,N_15805);
nand U19602 (N_19602,N_15746,N_16688);
or U19603 (N_19603,N_17316,N_15510);
nor U19604 (N_19604,N_15894,N_15249);
and U19605 (N_19605,N_16674,N_16528);
xor U19606 (N_19606,N_16940,N_17133);
and U19607 (N_19607,N_17702,N_15159);
nand U19608 (N_19608,N_16906,N_17498);
nand U19609 (N_19609,N_15283,N_15617);
and U19610 (N_19610,N_15092,N_16561);
or U19611 (N_19611,N_15897,N_16632);
and U19612 (N_19612,N_16009,N_16811);
and U19613 (N_19613,N_15723,N_15540);
xor U19614 (N_19614,N_15749,N_16335);
xor U19615 (N_19615,N_15170,N_16067);
xor U19616 (N_19616,N_16111,N_16304);
nor U19617 (N_19617,N_16202,N_17760);
nor U19618 (N_19618,N_16911,N_15287);
or U19619 (N_19619,N_17429,N_16363);
or U19620 (N_19620,N_16429,N_16718);
nand U19621 (N_19621,N_15355,N_15919);
or U19622 (N_19622,N_16672,N_15167);
and U19623 (N_19623,N_15099,N_15811);
or U19624 (N_19624,N_16216,N_17720);
and U19625 (N_19625,N_15440,N_16562);
or U19626 (N_19626,N_17301,N_15300);
or U19627 (N_19627,N_16364,N_15288);
nor U19628 (N_19628,N_17862,N_16285);
and U19629 (N_19629,N_15816,N_17410);
and U19630 (N_19630,N_15129,N_16176);
and U19631 (N_19631,N_17799,N_17732);
nor U19632 (N_19632,N_15819,N_16227);
xor U19633 (N_19633,N_16246,N_16508);
xor U19634 (N_19634,N_16840,N_15950);
nand U19635 (N_19635,N_15061,N_15088);
and U19636 (N_19636,N_16563,N_17417);
nand U19637 (N_19637,N_16314,N_15523);
nor U19638 (N_19638,N_17573,N_15027);
or U19639 (N_19639,N_17583,N_17221);
xnor U19640 (N_19640,N_17273,N_15541);
xor U19641 (N_19641,N_15145,N_17765);
nand U19642 (N_19642,N_15552,N_16825);
xor U19643 (N_19643,N_17860,N_16312);
nand U19644 (N_19644,N_15926,N_17575);
nor U19645 (N_19645,N_17369,N_15879);
or U19646 (N_19646,N_16899,N_15503);
and U19647 (N_19647,N_15337,N_16576);
xnor U19648 (N_19648,N_16068,N_15516);
or U19649 (N_19649,N_17313,N_17569);
or U19650 (N_19650,N_15107,N_15904);
nor U19651 (N_19651,N_15596,N_16783);
nor U19652 (N_19652,N_17022,N_17181);
nand U19653 (N_19653,N_16458,N_17011);
nor U19654 (N_19654,N_15334,N_15885);
nor U19655 (N_19655,N_17911,N_17013);
nor U19656 (N_19656,N_16490,N_16122);
or U19657 (N_19657,N_16579,N_17411);
nor U19658 (N_19658,N_15021,N_16250);
or U19659 (N_19659,N_15374,N_17711);
or U19660 (N_19660,N_16593,N_16504);
or U19661 (N_19661,N_17548,N_16948);
or U19662 (N_19662,N_16099,N_16499);
xnor U19663 (N_19663,N_16293,N_16768);
or U19664 (N_19664,N_16812,N_16803);
xor U19665 (N_19665,N_16810,N_17905);
xnor U19666 (N_19666,N_16830,N_16258);
nand U19667 (N_19667,N_15866,N_16630);
nand U19668 (N_19668,N_17886,N_16693);
nor U19669 (N_19669,N_15511,N_17712);
nor U19670 (N_19670,N_17936,N_17599);
nor U19671 (N_19671,N_17485,N_16817);
nor U19672 (N_19672,N_17590,N_15289);
and U19673 (N_19673,N_15701,N_16274);
and U19674 (N_19674,N_17892,N_15208);
xor U19675 (N_19675,N_16603,N_17646);
nand U19676 (N_19676,N_15183,N_17993);
or U19677 (N_19677,N_16812,N_16994);
nand U19678 (N_19678,N_15943,N_16328);
nor U19679 (N_19679,N_15665,N_15051);
and U19680 (N_19680,N_16378,N_16279);
nor U19681 (N_19681,N_17932,N_15972);
or U19682 (N_19682,N_15278,N_17578);
or U19683 (N_19683,N_16833,N_17883);
and U19684 (N_19684,N_15679,N_16857);
xnor U19685 (N_19685,N_15247,N_15256);
nor U19686 (N_19686,N_17440,N_16043);
and U19687 (N_19687,N_15380,N_17196);
nand U19688 (N_19688,N_16871,N_15532);
nor U19689 (N_19689,N_17314,N_16797);
and U19690 (N_19690,N_17985,N_15914);
nor U19691 (N_19691,N_17456,N_16593);
xor U19692 (N_19692,N_15906,N_15557);
xor U19693 (N_19693,N_17059,N_15996);
nor U19694 (N_19694,N_16722,N_15179);
nand U19695 (N_19695,N_17523,N_15590);
nand U19696 (N_19696,N_16000,N_17116);
nand U19697 (N_19697,N_15354,N_15880);
and U19698 (N_19698,N_15987,N_16309);
xnor U19699 (N_19699,N_15221,N_15235);
nor U19700 (N_19700,N_16140,N_16190);
xnor U19701 (N_19701,N_17805,N_15610);
nor U19702 (N_19702,N_17702,N_15673);
xnor U19703 (N_19703,N_15202,N_17695);
xnor U19704 (N_19704,N_16707,N_15544);
and U19705 (N_19705,N_17991,N_16643);
or U19706 (N_19706,N_17175,N_17303);
and U19707 (N_19707,N_16568,N_15677);
xnor U19708 (N_19708,N_15441,N_15558);
xor U19709 (N_19709,N_15308,N_16083);
or U19710 (N_19710,N_16331,N_16864);
and U19711 (N_19711,N_16724,N_16501);
xnor U19712 (N_19712,N_16156,N_15289);
nor U19713 (N_19713,N_17979,N_16565);
or U19714 (N_19714,N_17352,N_16418);
or U19715 (N_19715,N_16903,N_15772);
and U19716 (N_19716,N_15272,N_15735);
nor U19717 (N_19717,N_17842,N_15506);
xnor U19718 (N_19718,N_17486,N_16716);
or U19719 (N_19719,N_15971,N_16739);
nor U19720 (N_19720,N_15781,N_15023);
and U19721 (N_19721,N_17759,N_17708);
nand U19722 (N_19722,N_17637,N_17906);
and U19723 (N_19723,N_15173,N_15230);
and U19724 (N_19724,N_16299,N_17292);
or U19725 (N_19725,N_15742,N_16636);
nor U19726 (N_19726,N_15597,N_15409);
xnor U19727 (N_19727,N_17425,N_17103);
nand U19728 (N_19728,N_16862,N_16940);
nand U19729 (N_19729,N_17678,N_16029);
and U19730 (N_19730,N_17608,N_15340);
nor U19731 (N_19731,N_17079,N_15124);
nor U19732 (N_19732,N_17848,N_17150);
or U19733 (N_19733,N_16963,N_16145);
or U19734 (N_19734,N_17538,N_17108);
and U19735 (N_19735,N_15176,N_16128);
or U19736 (N_19736,N_15368,N_17558);
xnor U19737 (N_19737,N_17260,N_15524);
nor U19738 (N_19738,N_15197,N_16788);
xor U19739 (N_19739,N_16590,N_17483);
xor U19740 (N_19740,N_15167,N_17591);
nand U19741 (N_19741,N_17629,N_16100);
nand U19742 (N_19742,N_16108,N_17244);
nor U19743 (N_19743,N_17062,N_17676);
xor U19744 (N_19744,N_16665,N_15631);
or U19745 (N_19745,N_17558,N_15969);
nor U19746 (N_19746,N_15571,N_16750);
and U19747 (N_19747,N_16942,N_17159);
or U19748 (N_19748,N_16303,N_15159);
nand U19749 (N_19749,N_17066,N_15047);
nor U19750 (N_19750,N_17940,N_17548);
nor U19751 (N_19751,N_16545,N_17282);
xnor U19752 (N_19752,N_17547,N_15868);
or U19753 (N_19753,N_17680,N_16810);
nor U19754 (N_19754,N_15917,N_15975);
nor U19755 (N_19755,N_15016,N_16999);
nand U19756 (N_19756,N_16943,N_15041);
xnor U19757 (N_19757,N_15787,N_15512);
and U19758 (N_19758,N_17432,N_15145);
or U19759 (N_19759,N_17180,N_15186);
or U19760 (N_19760,N_15909,N_15863);
nand U19761 (N_19761,N_16192,N_15377);
and U19762 (N_19762,N_15509,N_15848);
nand U19763 (N_19763,N_17529,N_17937);
nand U19764 (N_19764,N_15636,N_17745);
nand U19765 (N_19765,N_17577,N_16754);
and U19766 (N_19766,N_16896,N_16679);
or U19767 (N_19767,N_17519,N_17565);
xnor U19768 (N_19768,N_17489,N_17631);
or U19769 (N_19769,N_17019,N_17211);
xor U19770 (N_19770,N_16310,N_15904);
nor U19771 (N_19771,N_17996,N_17927);
nor U19772 (N_19772,N_16435,N_15018);
nor U19773 (N_19773,N_17626,N_15465);
xnor U19774 (N_19774,N_15492,N_17788);
or U19775 (N_19775,N_17847,N_15552);
and U19776 (N_19776,N_15998,N_15099);
or U19777 (N_19777,N_15191,N_15013);
or U19778 (N_19778,N_17243,N_17591);
or U19779 (N_19779,N_17106,N_15213);
nand U19780 (N_19780,N_16589,N_16596);
nand U19781 (N_19781,N_17103,N_15554);
nor U19782 (N_19782,N_16062,N_15359);
xnor U19783 (N_19783,N_16872,N_16044);
nor U19784 (N_19784,N_15322,N_17928);
and U19785 (N_19785,N_16711,N_16284);
nand U19786 (N_19786,N_17993,N_16766);
nor U19787 (N_19787,N_15773,N_16077);
nor U19788 (N_19788,N_16376,N_17270);
nand U19789 (N_19789,N_17821,N_15137);
or U19790 (N_19790,N_15176,N_16439);
nor U19791 (N_19791,N_17463,N_15407);
or U19792 (N_19792,N_16600,N_15562);
nand U19793 (N_19793,N_17228,N_15772);
or U19794 (N_19794,N_16281,N_17070);
nand U19795 (N_19795,N_16049,N_17425);
and U19796 (N_19796,N_16085,N_16737);
nor U19797 (N_19797,N_15954,N_17136);
nor U19798 (N_19798,N_17901,N_17853);
and U19799 (N_19799,N_15576,N_17550);
or U19800 (N_19800,N_15823,N_17445);
nand U19801 (N_19801,N_17955,N_15442);
xor U19802 (N_19802,N_15918,N_17670);
and U19803 (N_19803,N_16741,N_17481);
and U19804 (N_19804,N_16721,N_15282);
nor U19805 (N_19805,N_15299,N_15385);
nand U19806 (N_19806,N_17690,N_15653);
xor U19807 (N_19807,N_16995,N_15009);
xnor U19808 (N_19808,N_16368,N_17195);
nor U19809 (N_19809,N_15546,N_15385);
nor U19810 (N_19810,N_16846,N_17220);
or U19811 (N_19811,N_15434,N_15078);
nand U19812 (N_19812,N_15517,N_15920);
nor U19813 (N_19813,N_15911,N_16272);
and U19814 (N_19814,N_16687,N_17504);
or U19815 (N_19815,N_16268,N_15235);
nor U19816 (N_19816,N_16964,N_17601);
or U19817 (N_19817,N_17796,N_15865);
nor U19818 (N_19818,N_17298,N_15910);
nor U19819 (N_19819,N_16867,N_17002);
nor U19820 (N_19820,N_17466,N_17573);
and U19821 (N_19821,N_17472,N_16740);
nor U19822 (N_19822,N_15132,N_17118);
nand U19823 (N_19823,N_17514,N_16319);
nor U19824 (N_19824,N_16006,N_17190);
or U19825 (N_19825,N_15007,N_17032);
nand U19826 (N_19826,N_16836,N_15566);
or U19827 (N_19827,N_17186,N_16162);
or U19828 (N_19828,N_17477,N_15787);
xor U19829 (N_19829,N_16739,N_16292);
or U19830 (N_19830,N_15591,N_17237);
or U19831 (N_19831,N_16039,N_15245);
and U19832 (N_19832,N_16816,N_17713);
xnor U19833 (N_19833,N_15451,N_16305);
and U19834 (N_19834,N_17741,N_17241);
nand U19835 (N_19835,N_17467,N_17168);
and U19836 (N_19836,N_15305,N_17255);
nor U19837 (N_19837,N_15928,N_16411);
nand U19838 (N_19838,N_15394,N_15271);
or U19839 (N_19839,N_17167,N_16959);
or U19840 (N_19840,N_17332,N_17065);
and U19841 (N_19841,N_16571,N_16929);
and U19842 (N_19842,N_15479,N_17132);
and U19843 (N_19843,N_16753,N_16345);
or U19844 (N_19844,N_15513,N_15912);
or U19845 (N_19845,N_15131,N_16680);
or U19846 (N_19846,N_15273,N_16353);
or U19847 (N_19847,N_17179,N_15837);
or U19848 (N_19848,N_16243,N_17185);
nor U19849 (N_19849,N_16470,N_17410);
nand U19850 (N_19850,N_15463,N_17675);
xnor U19851 (N_19851,N_16175,N_15816);
nand U19852 (N_19852,N_17688,N_16621);
or U19853 (N_19853,N_16747,N_15032);
or U19854 (N_19854,N_15498,N_17061);
xor U19855 (N_19855,N_16460,N_17344);
or U19856 (N_19856,N_17786,N_16980);
and U19857 (N_19857,N_15355,N_16509);
xnor U19858 (N_19858,N_17578,N_16591);
nand U19859 (N_19859,N_17694,N_17725);
nor U19860 (N_19860,N_16472,N_16001);
and U19861 (N_19861,N_16460,N_15128);
and U19862 (N_19862,N_16913,N_15596);
and U19863 (N_19863,N_15303,N_17183);
xnor U19864 (N_19864,N_16809,N_16545);
and U19865 (N_19865,N_16611,N_16652);
nor U19866 (N_19866,N_15324,N_17229);
nand U19867 (N_19867,N_17337,N_15055);
xor U19868 (N_19868,N_15627,N_15629);
and U19869 (N_19869,N_17084,N_16579);
or U19870 (N_19870,N_16445,N_17996);
or U19871 (N_19871,N_16891,N_16413);
xnor U19872 (N_19872,N_15676,N_15366);
nand U19873 (N_19873,N_17760,N_17265);
nor U19874 (N_19874,N_15696,N_17888);
nor U19875 (N_19875,N_15435,N_17929);
xor U19876 (N_19876,N_17296,N_17167);
nand U19877 (N_19877,N_15399,N_15338);
and U19878 (N_19878,N_17839,N_17584);
xnor U19879 (N_19879,N_16311,N_15571);
nor U19880 (N_19880,N_15284,N_15725);
nand U19881 (N_19881,N_16134,N_16236);
or U19882 (N_19882,N_15131,N_16968);
xor U19883 (N_19883,N_15936,N_16207);
or U19884 (N_19884,N_16764,N_16224);
and U19885 (N_19885,N_16471,N_15033);
xor U19886 (N_19886,N_16455,N_17584);
or U19887 (N_19887,N_16686,N_17695);
nand U19888 (N_19888,N_15876,N_17607);
and U19889 (N_19889,N_15738,N_15570);
xnor U19890 (N_19890,N_17620,N_17603);
or U19891 (N_19891,N_17022,N_16403);
nor U19892 (N_19892,N_16824,N_17073);
or U19893 (N_19893,N_15491,N_17552);
nor U19894 (N_19894,N_15025,N_17706);
nor U19895 (N_19895,N_17453,N_17418);
and U19896 (N_19896,N_15486,N_15462);
nand U19897 (N_19897,N_16635,N_15189);
nor U19898 (N_19898,N_17687,N_16832);
nand U19899 (N_19899,N_15527,N_16858);
or U19900 (N_19900,N_16787,N_15075);
xor U19901 (N_19901,N_17922,N_15376);
and U19902 (N_19902,N_15424,N_15121);
nor U19903 (N_19903,N_15678,N_16144);
nand U19904 (N_19904,N_17219,N_15468);
nand U19905 (N_19905,N_17857,N_15469);
or U19906 (N_19906,N_17213,N_17326);
nand U19907 (N_19907,N_16021,N_16031);
nor U19908 (N_19908,N_15930,N_15745);
and U19909 (N_19909,N_16526,N_15937);
nand U19910 (N_19910,N_15579,N_16462);
nor U19911 (N_19911,N_16262,N_16996);
or U19912 (N_19912,N_17762,N_16392);
nor U19913 (N_19913,N_17767,N_17686);
or U19914 (N_19914,N_16578,N_15374);
and U19915 (N_19915,N_15492,N_15475);
or U19916 (N_19916,N_17242,N_16848);
xor U19917 (N_19917,N_17110,N_15173);
nand U19918 (N_19918,N_16224,N_15013);
and U19919 (N_19919,N_16611,N_17503);
or U19920 (N_19920,N_15382,N_16925);
and U19921 (N_19921,N_16793,N_15178);
nor U19922 (N_19922,N_17312,N_15216);
nor U19923 (N_19923,N_15022,N_16740);
nor U19924 (N_19924,N_15460,N_17746);
and U19925 (N_19925,N_16901,N_16462);
xnor U19926 (N_19926,N_16846,N_16218);
xor U19927 (N_19927,N_15784,N_16467);
nor U19928 (N_19928,N_16813,N_15949);
and U19929 (N_19929,N_17494,N_17710);
or U19930 (N_19930,N_17857,N_17213);
xnor U19931 (N_19931,N_15214,N_17309);
or U19932 (N_19932,N_17209,N_15520);
or U19933 (N_19933,N_15268,N_15708);
nor U19934 (N_19934,N_16740,N_17683);
nor U19935 (N_19935,N_17571,N_16767);
nor U19936 (N_19936,N_17145,N_15283);
xor U19937 (N_19937,N_17021,N_17057);
or U19938 (N_19938,N_16012,N_17330);
nand U19939 (N_19939,N_16797,N_17811);
or U19940 (N_19940,N_17516,N_16605);
nand U19941 (N_19941,N_17338,N_16049);
and U19942 (N_19942,N_15560,N_15558);
xnor U19943 (N_19943,N_17967,N_17915);
and U19944 (N_19944,N_16707,N_15981);
or U19945 (N_19945,N_15516,N_17565);
xor U19946 (N_19946,N_17127,N_16588);
nand U19947 (N_19947,N_16647,N_15330);
or U19948 (N_19948,N_16116,N_17051);
nand U19949 (N_19949,N_17136,N_15725);
nand U19950 (N_19950,N_17154,N_16086);
or U19951 (N_19951,N_15367,N_17569);
nand U19952 (N_19952,N_15380,N_15699);
xor U19953 (N_19953,N_16943,N_17070);
or U19954 (N_19954,N_17115,N_16569);
nor U19955 (N_19955,N_15938,N_16243);
xnor U19956 (N_19956,N_17152,N_15594);
nand U19957 (N_19957,N_17189,N_15565);
xor U19958 (N_19958,N_17840,N_17894);
nand U19959 (N_19959,N_16183,N_15322);
nor U19960 (N_19960,N_16774,N_17443);
xor U19961 (N_19961,N_17400,N_16695);
and U19962 (N_19962,N_15159,N_16052);
nand U19963 (N_19963,N_15051,N_15019);
and U19964 (N_19964,N_17653,N_16202);
nor U19965 (N_19965,N_17424,N_17214);
or U19966 (N_19966,N_15777,N_17039);
xnor U19967 (N_19967,N_17375,N_15269);
xor U19968 (N_19968,N_15426,N_16775);
nand U19969 (N_19969,N_16640,N_17491);
xnor U19970 (N_19970,N_15362,N_17274);
nand U19971 (N_19971,N_17796,N_17528);
and U19972 (N_19972,N_17871,N_15735);
and U19973 (N_19973,N_16463,N_17584);
xnor U19974 (N_19974,N_15275,N_16766);
and U19975 (N_19975,N_15169,N_15501);
nand U19976 (N_19976,N_17306,N_17096);
or U19977 (N_19977,N_15395,N_17730);
nor U19978 (N_19978,N_17323,N_16638);
xnor U19979 (N_19979,N_15679,N_17049);
and U19980 (N_19980,N_17348,N_16307);
nor U19981 (N_19981,N_16231,N_15324);
and U19982 (N_19982,N_17908,N_16524);
xnor U19983 (N_19983,N_16382,N_17204);
xor U19984 (N_19984,N_16814,N_17152);
xor U19985 (N_19985,N_17081,N_16726);
nor U19986 (N_19986,N_15256,N_17607);
and U19987 (N_19987,N_16383,N_16473);
xor U19988 (N_19988,N_17859,N_15846);
or U19989 (N_19989,N_17178,N_15464);
xnor U19990 (N_19990,N_17899,N_15813);
nand U19991 (N_19991,N_16370,N_16887);
and U19992 (N_19992,N_15100,N_16404);
nand U19993 (N_19993,N_17859,N_17192);
nor U19994 (N_19994,N_17037,N_16550);
nor U19995 (N_19995,N_17444,N_16979);
nand U19996 (N_19996,N_15368,N_15071);
xor U19997 (N_19997,N_17215,N_17767);
nor U19998 (N_19998,N_15405,N_16254);
nand U19999 (N_19999,N_17433,N_17335);
nor U20000 (N_20000,N_16785,N_15709);
nand U20001 (N_20001,N_16652,N_17665);
and U20002 (N_20002,N_16180,N_15769);
and U20003 (N_20003,N_15958,N_15069);
nand U20004 (N_20004,N_15462,N_16579);
nand U20005 (N_20005,N_15806,N_15768);
nor U20006 (N_20006,N_16601,N_15782);
xor U20007 (N_20007,N_16920,N_15969);
nand U20008 (N_20008,N_16156,N_17197);
and U20009 (N_20009,N_17386,N_15301);
nand U20010 (N_20010,N_15487,N_17435);
nor U20011 (N_20011,N_17651,N_15126);
nor U20012 (N_20012,N_16970,N_17531);
nor U20013 (N_20013,N_16885,N_15175);
nand U20014 (N_20014,N_16009,N_15954);
xnor U20015 (N_20015,N_15111,N_16132);
nand U20016 (N_20016,N_15465,N_15075);
or U20017 (N_20017,N_15441,N_17329);
or U20018 (N_20018,N_17554,N_17271);
and U20019 (N_20019,N_15067,N_17383);
xor U20020 (N_20020,N_17876,N_17948);
or U20021 (N_20021,N_15174,N_17875);
xor U20022 (N_20022,N_17040,N_17018);
or U20023 (N_20023,N_17449,N_17410);
and U20024 (N_20024,N_17261,N_15906);
nor U20025 (N_20025,N_15670,N_17515);
nor U20026 (N_20026,N_16321,N_16557);
nand U20027 (N_20027,N_16759,N_15850);
or U20028 (N_20028,N_17947,N_16769);
or U20029 (N_20029,N_15219,N_17980);
nor U20030 (N_20030,N_16222,N_17978);
xor U20031 (N_20031,N_17455,N_16003);
and U20032 (N_20032,N_17342,N_16579);
or U20033 (N_20033,N_16223,N_16308);
xnor U20034 (N_20034,N_17185,N_16424);
or U20035 (N_20035,N_17172,N_16889);
and U20036 (N_20036,N_16298,N_16999);
nand U20037 (N_20037,N_15825,N_15690);
or U20038 (N_20038,N_16213,N_17254);
xor U20039 (N_20039,N_17408,N_15104);
and U20040 (N_20040,N_17179,N_16010);
xnor U20041 (N_20041,N_17229,N_17960);
or U20042 (N_20042,N_15412,N_16243);
and U20043 (N_20043,N_17752,N_17173);
nor U20044 (N_20044,N_17229,N_15163);
and U20045 (N_20045,N_17249,N_17869);
nand U20046 (N_20046,N_16912,N_16719);
or U20047 (N_20047,N_15518,N_16198);
and U20048 (N_20048,N_17957,N_15908);
nand U20049 (N_20049,N_17697,N_15430);
or U20050 (N_20050,N_15801,N_16747);
xnor U20051 (N_20051,N_15412,N_16301);
and U20052 (N_20052,N_15692,N_15530);
nand U20053 (N_20053,N_16381,N_17701);
or U20054 (N_20054,N_17767,N_17152);
and U20055 (N_20055,N_16894,N_15265);
and U20056 (N_20056,N_16837,N_16576);
nand U20057 (N_20057,N_17061,N_17608);
nand U20058 (N_20058,N_15542,N_16303);
or U20059 (N_20059,N_17924,N_15435);
and U20060 (N_20060,N_17178,N_16822);
nand U20061 (N_20061,N_16748,N_17387);
and U20062 (N_20062,N_16300,N_15488);
nand U20063 (N_20063,N_16572,N_17878);
nand U20064 (N_20064,N_16022,N_16901);
nand U20065 (N_20065,N_17676,N_17840);
xnor U20066 (N_20066,N_16902,N_17309);
nor U20067 (N_20067,N_17006,N_16924);
nand U20068 (N_20068,N_16369,N_15636);
and U20069 (N_20069,N_17140,N_16978);
or U20070 (N_20070,N_17114,N_16187);
nand U20071 (N_20071,N_15014,N_16304);
or U20072 (N_20072,N_16874,N_17611);
or U20073 (N_20073,N_16057,N_16624);
xor U20074 (N_20074,N_17292,N_17021);
nand U20075 (N_20075,N_16658,N_16175);
nor U20076 (N_20076,N_15667,N_16012);
and U20077 (N_20077,N_15834,N_17926);
or U20078 (N_20078,N_17416,N_16141);
or U20079 (N_20079,N_16718,N_15312);
nand U20080 (N_20080,N_15515,N_17001);
xnor U20081 (N_20081,N_15365,N_15011);
and U20082 (N_20082,N_15289,N_17945);
or U20083 (N_20083,N_16349,N_17968);
nor U20084 (N_20084,N_17939,N_16236);
nand U20085 (N_20085,N_16849,N_15999);
xnor U20086 (N_20086,N_15483,N_15821);
or U20087 (N_20087,N_15463,N_15809);
nand U20088 (N_20088,N_16649,N_15585);
or U20089 (N_20089,N_17864,N_17396);
and U20090 (N_20090,N_17937,N_17213);
nor U20091 (N_20091,N_15784,N_15396);
and U20092 (N_20092,N_16803,N_15147);
nor U20093 (N_20093,N_15226,N_17637);
xor U20094 (N_20094,N_17266,N_15814);
xnor U20095 (N_20095,N_15158,N_15388);
or U20096 (N_20096,N_16492,N_17833);
nor U20097 (N_20097,N_15960,N_16441);
or U20098 (N_20098,N_16711,N_17857);
nor U20099 (N_20099,N_15955,N_17798);
and U20100 (N_20100,N_17061,N_17167);
nand U20101 (N_20101,N_17537,N_17803);
and U20102 (N_20102,N_16265,N_16972);
nor U20103 (N_20103,N_15783,N_15224);
xnor U20104 (N_20104,N_15234,N_16513);
nand U20105 (N_20105,N_16238,N_17630);
and U20106 (N_20106,N_15848,N_17336);
nand U20107 (N_20107,N_15167,N_17258);
nor U20108 (N_20108,N_17648,N_16244);
xor U20109 (N_20109,N_17270,N_15484);
nand U20110 (N_20110,N_15329,N_17623);
nand U20111 (N_20111,N_15557,N_16776);
or U20112 (N_20112,N_16617,N_15774);
xor U20113 (N_20113,N_17475,N_15581);
nor U20114 (N_20114,N_15819,N_17342);
and U20115 (N_20115,N_17849,N_15321);
nor U20116 (N_20116,N_15641,N_16302);
xnor U20117 (N_20117,N_15307,N_15139);
or U20118 (N_20118,N_16461,N_16798);
or U20119 (N_20119,N_16495,N_16592);
nand U20120 (N_20120,N_16136,N_16332);
xnor U20121 (N_20121,N_17706,N_17863);
xnor U20122 (N_20122,N_15393,N_17993);
or U20123 (N_20123,N_17731,N_16344);
or U20124 (N_20124,N_17657,N_15988);
nand U20125 (N_20125,N_16972,N_15267);
xnor U20126 (N_20126,N_15765,N_17755);
or U20127 (N_20127,N_16229,N_17659);
nor U20128 (N_20128,N_17462,N_15573);
and U20129 (N_20129,N_16912,N_15473);
nor U20130 (N_20130,N_16878,N_16791);
nand U20131 (N_20131,N_15352,N_16620);
and U20132 (N_20132,N_16741,N_17209);
nand U20133 (N_20133,N_15497,N_17498);
or U20134 (N_20134,N_17640,N_15386);
and U20135 (N_20135,N_17123,N_15844);
and U20136 (N_20136,N_17786,N_17166);
nand U20137 (N_20137,N_17948,N_15356);
xor U20138 (N_20138,N_16423,N_16701);
and U20139 (N_20139,N_17019,N_16854);
xor U20140 (N_20140,N_16698,N_16926);
xor U20141 (N_20141,N_16146,N_17899);
or U20142 (N_20142,N_17754,N_15078);
and U20143 (N_20143,N_17285,N_16164);
nor U20144 (N_20144,N_15894,N_15316);
nand U20145 (N_20145,N_17893,N_16208);
xor U20146 (N_20146,N_17504,N_17011);
and U20147 (N_20147,N_16544,N_16731);
and U20148 (N_20148,N_15824,N_17134);
nand U20149 (N_20149,N_16154,N_15041);
and U20150 (N_20150,N_17808,N_16120);
and U20151 (N_20151,N_17126,N_16837);
and U20152 (N_20152,N_16259,N_15315);
nor U20153 (N_20153,N_16076,N_17100);
nor U20154 (N_20154,N_17664,N_17899);
nand U20155 (N_20155,N_15104,N_17698);
and U20156 (N_20156,N_17594,N_17411);
or U20157 (N_20157,N_15032,N_17090);
nor U20158 (N_20158,N_16226,N_16037);
xnor U20159 (N_20159,N_15467,N_16269);
and U20160 (N_20160,N_16915,N_15446);
xor U20161 (N_20161,N_17521,N_15355);
or U20162 (N_20162,N_15445,N_16196);
xnor U20163 (N_20163,N_16780,N_15058);
and U20164 (N_20164,N_15266,N_16477);
and U20165 (N_20165,N_17737,N_17629);
and U20166 (N_20166,N_17242,N_16508);
nand U20167 (N_20167,N_17920,N_16673);
nand U20168 (N_20168,N_17189,N_15863);
nor U20169 (N_20169,N_16210,N_15221);
xnor U20170 (N_20170,N_15775,N_15848);
nor U20171 (N_20171,N_16972,N_16629);
xnor U20172 (N_20172,N_17249,N_15630);
or U20173 (N_20173,N_17619,N_16860);
xnor U20174 (N_20174,N_16771,N_16941);
xor U20175 (N_20175,N_16763,N_16964);
or U20176 (N_20176,N_15713,N_17936);
nor U20177 (N_20177,N_17514,N_15202);
nand U20178 (N_20178,N_17039,N_16634);
and U20179 (N_20179,N_16645,N_15484);
nand U20180 (N_20180,N_15158,N_15765);
and U20181 (N_20181,N_17372,N_16036);
nand U20182 (N_20182,N_17872,N_15046);
xor U20183 (N_20183,N_17692,N_17710);
nand U20184 (N_20184,N_16308,N_15012);
nand U20185 (N_20185,N_16349,N_16518);
or U20186 (N_20186,N_17063,N_15040);
nor U20187 (N_20187,N_16446,N_15213);
or U20188 (N_20188,N_17181,N_15395);
nand U20189 (N_20189,N_16701,N_17389);
nor U20190 (N_20190,N_16655,N_16282);
nand U20191 (N_20191,N_16226,N_16956);
nand U20192 (N_20192,N_16556,N_17187);
and U20193 (N_20193,N_15672,N_16034);
nor U20194 (N_20194,N_17318,N_17135);
or U20195 (N_20195,N_16970,N_15726);
nand U20196 (N_20196,N_15402,N_17504);
or U20197 (N_20197,N_16304,N_16086);
nor U20198 (N_20198,N_17986,N_15149);
nand U20199 (N_20199,N_16061,N_15491);
nor U20200 (N_20200,N_16950,N_16098);
or U20201 (N_20201,N_17498,N_15534);
nand U20202 (N_20202,N_16687,N_17141);
nor U20203 (N_20203,N_17017,N_16301);
or U20204 (N_20204,N_16115,N_17417);
and U20205 (N_20205,N_16846,N_15511);
xnor U20206 (N_20206,N_16198,N_16319);
and U20207 (N_20207,N_17152,N_16669);
xnor U20208 (N_20208,N_17546,N_16504);
xnor U20209 (N_20209,N_17898,N_15204);
xor U20210 (N_20210,N_15249,N_17230);
and U20211 (N_20211,N_17095,N_16134);
and U20212 (N_20212,N_16423,N_16735);
or U20213 (N_20213,N_16063,N_17624);
nand U20214 (N_20214,N_15840,N_15832);
xor U20215 (N_20215,N_16668,N_17377);
nor U20216 (N_20216,N_15133,N_17428);
nor U20217 (N_20217,N_16791,N_15012);
and U20218 (N_20218,N_16647,N_15783);
xnor U20219 (N_20219,N_17845,N_15636);
nor U20220 (N_20220,N_16544,N_16418);
or U20221 (N_20221,N_17731,N_15608);
xor U20222 (N_20222,N_17644,N_17801);
nand U20223 (N_20223,N_16508,N_15781);
xor U20224 (N_20224,N_15977,N_17551);
and U20225 (N_20225,N_15289,N_16398);
xnor U20226 (N_20226,N_17395,N_16086);
nor U20227 (N_20227,N_17656,N_16329);
xnor U20228 (N_20228,N_15244,N_17822);
nand U20229 (N_20229,N_15703,N_16808);
and U20230 (N_20230,N_17820,N_17278);
or U20231 (N_20231,N_15322,N_16587);
and U20232 (N_20232,N_16834,N_15534);
or U20233 (N_20233,N_17893,N_15201);
and U20234 (N_20234,N_15834,N_16665);
xor U20235 (N_20235,N_15010,N_17423);
or U20236 (N_20236,N_16209,N_17990);
nand U20237 (N_20237,N_15667,N_15858);
nand U20238 (N_20238,N_16320,N_17605);
and U20239 (N_20239,N_17341,N_17940);
nand U20240 (N_20240,N_16496,N_16587);
xor U20241 (N_20241,N_16403,N_16276);
nor U20242 (N_20242,N_17727,N_16737);
nand U20243 (N_20243,N_16155,N_17618);
or U20244 (N_20244,N_16398,N_17254);
or U20245 (N_20245,N_17199,N_17237);
and U20246 (N_20246,N_16778,N_17959);
nor U20247 (N_20247,N_15648,N_17110);
or U20248 (N_20248,N_17188,N_15073);
nor U20249 (N_20249,N_16419,N_15107);
nor U20250 (N_20250,N_15968,N_15083);
xnor U20251 (N_20251,N_17100,N_16829);
xnor U20252 (N_20252,N_17115,N_16975);
nand U20253 (N_20253,N_15823,N_16608);
nor U20254 (N_20254,N_15009,N_17631);
and U20255 (N_20255,N_15210,N_17583);
xnor U20256 (N_20256,N_17430,N_16935);
nor U20257 (N_20257,N_17364,N_17463);
or U20258 (N_20258,N_16305,N_15512);
and U20259 (N_20259,N_16182,N_15825);
nand U20260 (N_20260,N_16375,N_15373);
nor U20261 (N_20261,N_16559,N_15883);
nand U20262 (N_20262,N_16312,N_16020);
xor U20263 (N_20263,N_16977,N_17970);
nor U20264 (N_20264,N_15007,N_17465);
and U20265 (N_20265,N_15734,N_17984);
nor U20266 (N_20266,N_17834,N_17215);
and U20267 (N_20267,N_15036,N_15436);
or U20268 (N_20268,N_17376,N_16099);
nor U20269 (N_20269,N_17902,N_17799);
and U20270 (N_20270,N_15118,N_17196);
and U20271 (N_20271,N_17177,N_16648);
or U20272 (N_20272,N_17955,N_15101);
xnor U20273 (N_20273,N_17459,N_17398);
or U20274 (N_20274,N_15884,N_16403);
or U20275 (N_20275,N_15867,N_16374);
xnor U20276 (N_20276,N_16395,N_17404);
and U20277 (N_20277,N_16045,N_15988);
or U20278 (N_20278,N_17367,N_15125);
nand U20279 (N_20279,N_16392,N_16585);
nor U20280 (N_20280,N_16437,N_17538);
nor U20281 (N_20281,N_15551,N_17921);
xor U20282 (N_20282,N_17853,N_17557);
nand U20283 (N_20283,N_15806,N_16641);
xor U20284 (N_20284,N_15850,N_17532);
nand U20285 (N_20285,N_15295,N_17034);
xor U20286 (N_20286,N_17685,N_17072);
or U20287 (N_20287,N_15216,N_17184);
nor U20288 (N_20288,N_15828,N_17735);
xor U20289 (N_20289,N_17687,N_16336);
and U20290 (N_20290,N_16126,N_16754);
and U20291 (N_20291,N_16468,N_16407);
nand U20292 (N_20292,N_15446,N_17374);
and U20293 (N_20293,N_17722,N_17880);
nand U20294 (N_20294,N_16614,N_16617);
nor U20295 (N_20295,N_16330,N_17296);
and U20296 (N_20296,N_17843,N_17291);
or U20297 (N_20297,N_17073,N_15489);
and U20298 (N_20298,N_17688,N_17797);
or U20299 (N_20299,N_17068,N_17324);
nor U20300 (N_20300,N_15982,N_15479);
nand U20301 (N_20301,N_16518,N_17551);
xnor U20302 (N_20302,N_17020,N_16018);
and U20303 (N_20303,N_16779,N_15512);
xor U20304 (N_20304,N_16437,N_17198);
or U20305 (N_20305,N_16183,N_15039);
nor U20306 (N_20306,N_16702,N_17608);
or U20307 (N_20307,N_17085,N_17121);
nor U20308 (N_20308,N_16495,N_17466);
xor U20309 (N_20309,N_15845,N_16961);
or U20310 (N_20310,N_16407,N_16479);
nor U20311 (N_20311,N_17630,N_16785);
or U20312 (N_20312,N_16076,N_16428);
xnor U20313 (N_20313,N_15726,N_15881);
xor U20314 (N_20314,N_17668,N_16140);
or U20315 (N_20315,N_17818,N_17509);
xor U20316 (N_20316,N_17621,N_17981);
nor U20317 (N_20317,N_15766,N_15765);
nor U20318 (N_20318,N_15162,N_17923);
nor U20319 (N_20319,N_17962,N_17608);
nor U20320 (N_20320,N_16178,N_17210);
nand U20321 (N_20321,N_16865,N_17974);
or U20322 (N_20322,N_16114,N_15787);
nor U20323 (N_20323,N_17891,N_15219);
nor U20324 (N_20324,N_17607,N_16037);
or U20325 (N_20325,N_17712,N_15604);
or U20326 (N_20326,N_17657,N_15032);
nand U20327 (N_20327,N_15428,N_17963);
nor U20328 (N_20328,N_15188,N_17968);
nor U20329 (N_20329,N_15427,N_17947);
nor U20330 (N_20330,N_16934,N_17804);
nand U20331 (N_20331,N_15772,N_15746);
nand U20332 (N_20332,N_15135,N_15265);
and U20333 (N_20333,N_17724,N_16588);
nand U20334 (N_20334,N_16961,N_15663);
nand U20335 (N_20335,N_15860,N_16183);
xor U20336 (N_20336,N_16613,N_17035);
nor U20337 (N_20337,N_17817,N_16367);
xnor U20338 (N_20338,N_16698,N_15948);
and U20339 (N_20339,N_15139,N_17181);
or U20340 (N_20340,N_16021,N_16155);
or U20341 (N_20341,N_17725,N_15926);
xor U20342 (N_20342,N_17110,N_15971);
or U20343 (N_20343,N_15436,N_16549);
nand U20344 (N_20344,N_17452,N_15502);
nor U20345 (N_20345,N_15596,N_15497);
and U20346 (N_20346,N_17722,N_15145);
nand U20347 (N_20347,N_15916,N_17034);
nor U20348 (N_20348,N_17038,N_16671);
xnor U20349 (N_20349,N_16946,N_16872);
or U20350 (N_20350,N_16057,N_15040);
or U20351 (N_20351,N_16032,N_17117);
nand U20352 (N_20352,N_16745,N_15667);
xor U20353 (N_20353,N_16624,N_15087);
xnor U20354 (N_20354,N_16289,N_16598);
nor U20355 (N_20355,N_15766,N_15227);
xnor U20356 (N_20356,N_17518,N_15884);
xor U20357 (N_20357,N_15241,N_16871);
xnor U20358 (N_20358,N_15787,N_15777);
and U20359 (N_20359,N_15700,N_17290);
nor U20360 (N_20360,N_16881,N_16826);
and U20361 (N_20361,N_15093,N_15809);
nand U20362 (N_20362,N_15782,N_16943);
xnor U20363 (N_20363,N_15799,N_16502);
and U20364 (N_20364,N_17016,N_15350);
nand U20365 (N_20365,N_17444,N_17989);
and U20366 (N_20366,N_16038,N_15220);
or U20367 (N_20367,N_16597,N_15857);
nor U20368 (N_20368,N_16751,N_16061);
nor U20369 (N_20369,N_16608,N_16580);
and U20370 (N_20370,N_15562,N_15928);
nor U20371 (N_20371,N_15584,N_16745);
or U20372 (N_20372,N_15877,N_17481);
xor U20373 (N_20373,N_16993,N_17755);
xnor U20374 (N_20374,N_15806,N_16741);
nor U20375 (N_20375,N_16225,N_15791);
and U20376 (N_20376,N_15161,N_17587);
xnor U20377 (N_20377,N_15184,N_17350);
or U20378 (N_20378,N_15153,N_16859);
xor U20379 (N_20379,N_17766,N_15627);
or U20380 (N_20380,N_16627,N_15591);
or U20381 (N_20381,N_17929,N_17854);
xnor U20382 (N_20382,N_16933,N_17580);
xnor U20383 (N_20383,N_15198,N_16715);
nand U20384 (N_20384,N_15257,N_16666);
and U20385 (N_20385,N_15065,N_17601);
xor U20386 (N_20386,N_15398,N_16124);
and U20387 (N_20387,N_15018,N_17853);
nand U20388 (N_20388,N_15212,N_15788);
xor U20389 (N_20389,N_15646,N_17967);
and U20390 (N_20390,N_16024,N_15091);
or U20391 (N_20391,N_16298,N_17880);
xnor U20392 (N_20392,N_15904,N_16801);
nor U20393 (N_20393,N_17238,N_15354);
xnor U20394 (N_20394,N_16168,N_15314);
nor U20395 (N_20395,N_16952,N_17057);
and U20396 (N_20396,N_15738,N_17457);
nor U20397 (N_20397,N_17203,N_17560);
nand U20398 (N_20398,N_17385,N_17481);
or U20399 (N_20399,N_15416,N_16855);
and U20400 (N_20400,N_16791,N_17790);
nand U20401 (N_20401,N_16572,N_15475);
and U20402 (N_20402,N_16517,N_16056);
xnor U20403 (N_20403,N_15090,N_15858);
nor U20404 (N_20404,N_16098,N_17379);
nor U20405 (N_20405,N_17751,N_15188);
xnor U20406 (N_20406,N_16442,N_15506);
nor U20407 (N_20407,N_17203,N_17679);
xor U20408 (N_20408,N_16007,N_17323);
and U20409 (N_20409,N_15964,N_16036);
nand U20410 (N_20410,N_16781,N_15249);
or U20411 (N_20411,N_16606,N_16927);
nand U20412 (N_20412,N_15518,N_15275);
nand U20413 (N_20413,N_16164,N_17517);
and U20414 (N_20414,N_17302,N_16513);
nor U20415 (N_20415,N_15270,N_15070);
xor U20416 (N_20416,N_16634,N_15761);
nor U20417 (N_20417,N_15998,N_17430);
xor U20418 (N_20418,N_17452,N_17851);
nor U20419 (N_20419,N_15453,N_17405);
or U20420 (N_20420,N_17232,N_15855);
xnor U20421 (N_20421,N_16687,N_17533);
nor U20422 (N_20422,N_15065,N_15403);
nand U20423 (N_20423,N_16672,N_17176);
xor U20424 (N_20424,N_15446,N_16899);
and U20425 (N_20425,N_16759,N_17196);
nor U20426 (N_20426,N_16525,N_16935);
nand U20427 (N_20427,N_15452,N_17925);
nor U20428 (N_20428,N_15917,N_16917);
nand U20429 (N_20429,N_16143,N_16765);
or U20430 (N_20430,N_15125,N_15279);
or U20431 (N_20431,N_15090,N_15410);
xor U20432 (N_20432,N_16242,N_16029);
nor U20433 (N_20433,N_15640,N_17233);
nand U20434 (N_20434,N_15698,N_16345);
xor U20435 (N_20435,N_16512,N_16511);
nor U20436 (N_20436,N_16456,N_15270);
nand U20437 (N_20437,N_15465,N_15355);
and U20438 (N_20438,N_15671,N_15993);
or U20439 (N_20439,N_16746,N_16551);
nor U20440 (N_20440,N_15098,N_17090);
xnor U20441 (N_20441,N_17684,N_15531);
and U20442 (N_20442,N_17634,N_15659);
nand U20443 (N_20443,N_16267,N_16792);
or U20444 (N_20444,N_16796,N_17237);
nand U20445 (N_20445,N_16668,N_17675);
xnor U20446 (N_20446,N_16216,N_17989);
and U20447 (N_20447,N_17625,N_16494);
nand U20448 (N_20448,N_15922,N_16583);
and U20449 (N_20449,N_16916,N_17295);
nand U20450 (N_20450,N_17996,N_16954);
nand U20451 (N_20451,N_16453,N_16652);
xor U20452 (N_20452,N_16294,N_17564);
or U20453 (N_20453,N_15091,N_17016);
or U20454 (N_20454,N_15158,N_16274);
xor U20455 (N_20455,N_16778,N_17254);
xnor U20456 (N_20456,N_16412,N_16148);
or U20457 (N_20457,N_15106,N_15301);
xnor U20458 (N_20458,N_16500,N_15029);
xnor U20459 (N_20459,N_17604,N_16277);
xnor U20460 (N_20460,N_17720,N_17206);
and U20461 (N_20461,N_15032,N_17826);
and U20462 (N_20462,N_16701,N_16738);
nor U20463 (N_20463,N_17073,N_16027);
or U20464 (N_20464,N_15943,N_15793);
or U20465 (N_20465,N_17122,N_16299);
and U20466 (N_20466,N_15467,N_15259);
or U20467 (N_20467,N_17227,N_16462);
or U20468 (N_20468,N_16602,N_17435);
xor U20469 (N_20469,N_16040,N_16758);
or U20470 (N_20470,N_15922,N_15528);
xnor U20471 (N_20471,N_17448,N_16866);
xnor U20472 (N_20472,N_17230,N_16533);
nor U20473 (N_20473,N_15322,N_17585);
or U20474 (N_20474,N_17619,N_17069);
nand U20475 (N_20475,N_15751,N_15749);
xnor U20476 (N_20476,N_15666,N_15505);
xor U20477 (N_20477,N_15525,N_15841);
or U20478 (N_20478,N_15747,N_15470);
nor U20479 (N_20479,N_15106,N_17219);
nor U20480 (N_20480,N_15728,N_17605);
or U20481 (N_20481,N_16369,N_17149);
or U20482 (N_20482,N_16698,N_15460);
nor U20483 (N_20483,N_15127,N_16325);
or U20484 (N_20484,N_16326,N_17372);
and U20485 (N_20485,N_16616,N_16093);
or U20486 (N_20486,N_16569,N_15302);
xor U20487 (N_20487,N_17103,N_17752);
xor U20488 (N_20488,N_16399,N_16368);
and U20489 (N_20489,N_15811,N_16898);
nor U20490 (N_20490,N_16429,N_16295);
nand U20491 (N_20491,N_15205,N_16442);
xnor U20492 (N_20492,N_16904,N_16854);
nor U20493 (N_20493,N_15725,N_17482);
or U20494 (N_20494,N_17690,N_17447);
xor U20495 (N_20495,N_16882,N_17709);
xor U20496 (N_20496,N_15439,N_16221);
xnor U20497 (N_20497,N_17665,N_16760);
nor U20498 (N_20498,N_17318,N_16100);
nand U20499 (N_20499,N_16750,N_16987);
nand U20500 (N_20500,N_17073,N_17545);
and U20501 (N_20501,N_15057,N_16897);
and U20502 (N_20502,N_17049,N_17057);
nand U20503 (N_20503,N_15294,N_16054);
nor U20504 (N_20504,N_17905,N_15038);
and U20505 (N_20505,N_16999,N_16750);
and U20506 (N_20506,N_16038,N_16080);
nand U20507 (N_20507,N_15018,N_16531);
and U20508 (N_20508,N_15700,N_17420);
nand U20509 (N_20509,N_17150,N_17510);
nand U20510 (N_20510,N_15312,N_16209);
nor U20511 (N_20511,N_17151,N_16242);
nor U20512 (N_20512,N_15629,N_16833);
nand U20513 (N_20513,N_15473,N_17022);
and U20514 (N_20514,N_17012,N_15293);
xnor U20515 (N_20515,N_17604,N_15585);
xor U20516 (N_20516,N_17114,N_15183);
nor U20517 (N_20517,N_16390,N_17321);
or U20518 (N_20518,N_15327,N_16585);
nor U20519 (N_20519,N_16783,N_17605);
or U20520 (N_20520,N_16759,N_17425);
nor U20521 (N_20521,N_16050,N_16926);
nand U20522 (N_20522,N_15663,N_16172);
nor U20523 (N_20523,N_16244,N_15271);
and U20524 (N_20524,N_17922,N_16933);
or U20525 (N_20525,N_17687,N_15501);
nand U20526 (N_20526,N_16489,N_15992);
or U20527 (N_20527,N_17672,N_16272);
xnor U20528 (N_20528,N_16910,N_16006);
nor U20529 (N_20529,N_15611,N_16988);
nand U20530 (N_20530,N_16436,N_15275);
or U20531 (N_20531,N_15022,N_16474);
or U20532 (N_20532,N_16221,N_17890);
nand U20533 (N_20533,N_15552,N_17043);
and U20534 (N_20534,N_16582,N_16859);
nand U20535 (N_20535,N_17835,N_16262);
nand U20536 (N_20536,N_17419,N_15364);
nor U20537 (N_20537,N_17718,N_15831);
and U20538 (N_20538,N_16577,N_15005);
nand U20539 (N_20539,N_15782,N_16501);
xnor U20540 (N_20540,N_16638,N_15595);
nand U20541 (N_20541,N_15657,N_15313);
nor U20542 (N_20542,N_16494,N_15458);
xnor U20543 (N_20543,N_16845,N_17488);
and U20544 (N_20544,N_17165,N_15577);
nor U20545 (N_20545,N_16549,N_16404);
or U20546 (N_20546,N_15145,N_17075);
nor U20547 (N_20547,N_15339,N_16421);
nor U20548 (N_20548,N_15238,N_17571);
or U20549 (N_20549,N_17888,N_17612);
nand U20550 (N_20550,N_17706,N_16843);
xor U20551 (N_20551,N_16065,N_17478);
or U20552 (N_20552,N_17035,N_17417);
nor U20553 (N_20553,N_16988,N_15863);
or U20554 (N_20554,N_15973,N_17456);
xor U20555 (N_20555,N_17180,N_16779);
nor U20556 (N_20556,N_17126,N_16409);
nand U20557 (N_20557,N_17043,N_15408);
and U20558 (N_20558,N_15155,N_16304);
or U20559 (N_20559,N_17845,N_15087);
nand U20560 (N_20560,N_17012,N_17621);
nor U20561 (N_20561,N_16988,N_15164);
or U20562 (N_20562,N_15336,N_17575);
nor U20563 (N_20563,N_15201,N_15864);
or U20564 (N_20564,N_15791,N_16843);
nand U20565 (N_20565,N_15827,N_17232);
nand U20566 (N_20566,N_16903,N_16577);
nor U20567 (N_20567,N_17135,N_15635);
nor U20568 (N_20568,N_15034,N_17292);
nand U20569 (N_20569,N_17416,N_17962);
xnor U20570 (N_20570,N_15585,N_15687);
xor U20571 (N_20571,N_17963,N_15801);
or U20572 (N_20572,N_15955,N_16836);
or U20573 (N_20573,N_15889,N_16233);
xor U20574 (N_20574,N_17214,N_15843);
nand U20575 (N_20575,N_17331,N_16309);
nor U20576 (N_20576,N_16107,N_16317);
xnor U20577 (N_20577,N_17646,N_15962);
and U20578 (N_20578,N_17399,N_17773);
nor U20579 (N_20579,N_15466,N_17635);
nand U20580 (N_20580,N_17663,N_17905);
or U20581 (N_20581,N_17564,N_15412);
or U20582 (N_20582,N_15876,N_15067);
and U20583 (N_20583,N_17001,N_17484);
nand U20584 (N_20584,N_16271,N_15110);
and U20585 (N_20585,N_15380,N_16915);
nor U20586 (N_20586,N_16275,N_17607);
and U20587 (N_20587,N_16055,N_15000);
or U20588 (N_20588,N_17771,N_16481);
xor U20589 (N_20589,N_15422,N_15945);
nor U20590 (N_20590,N_17454,N_17908);
nor U20591 (N_20591,N_16954,N_17137);
nor U20592 (N_20592,N_17810,N_15462);
xnor U20593 (N_20593,N_16234,N_16862);
xnor U20594 (N_20594,N_16932,N_16766);
nor U20595 (N_20595,N_16627,N_15286);
nor U20596 (N_20596,N_17521,N_15109);
nor U20597 (N_20597,N_15414,N_15944);
nand U20598 (N_20598,N_17371,N_15569);
nor U20599 (N_20599,N_16333,N_16943);
nor U20600 (N_20600,N_17946,N_15009);
and U20601 (N_20601,N_16151,N_16564);
and U20602 (N_20602,N_17082,N_17742);
nand U20603 (N_20603,N_15392,N_15981);
xnor U20604 (N_20604,N_16097,N_17282);
xnor U20605 (N_20605,N_17063,N_17191);
xor U20606 (N_20606,N_17957,N_16459);
nor U20607 (N_20607,N_15592,N_17429);
xor U20608 (N_20608,N_15314,N_15971);
and U20609 (N_20609,N_17065,N_15457);
nor U20610 (N_20610,N_16556,N_15834);
and U20611 (N_20611,N_15608,N_15073);
nand U20612 (N_20612,N_15154,N_15630);
and U20613 (N_20613,N_17129,N_17754);
nor U20614 (N_20614,N_15259,N_16319);
or U20615 (N_20615,N_15363,N_17718);
xnor U20616 (N_20616,N_16548,N_17588);
nor U20617 (N_20617,N_15024,N_16161);
nor U20618 (N_20618,N_15921,N_15425);
nand U20619 (N_20619,N_15321,N_17640);
xnor U20620 (N_20620,N_17672,N_16199);
and U20621 (N_20621,N_17119,N_17965);
nor U20622 (N_20622,N_15451,N_16757);
or U20623 (N_20623,N_15639,N_15631);
nor U20624 (N_20624,N_16439,N_16080);
or U20625 (N_20625,N_15437,N_15768);
xnor U20626 (N_20626,N_15989,N_16803);
nor U20627 (N_20627,N_16655,N_15631);
xnor U20628 (N_20628,N_17579,N_15181);
nand U20629 (N_20629,N_17389,N_16258);
nand U20630 (N_20630,N_16678,N_17214);
and U20631 (N_20631,N_16604,N_16681);
nand U20632 (N_20632,N_15187,N_15758);
xor U20633 (N_20633,N_16168,N_15159);
xnor U20634 (N_20634,N_16570,N_15931);
and U20635 (N_20635,N_15736,N_16969);
or U20636 (N_20636,N_16171,N_16765);
and U20637 (N_20637,N_17399,N_15314);
xor U20638 (N_20638,N_16301,N_16792);
or U20639 (N_20639,N_15461,N_17233);
nor U20640 (N_20640,N_17031,N_15980);
xor U20641 (N_20641,N_17590,N_17939);
xnor U20642 (N_20642,N_17262,N_17217);
nor U20643 (N_20643,N_17525,N_16415);
or U20644 (N_20644,N_15243,N_16091);
nand U20645 (N_20645,N_17152,N_16680);
and U20646 (N_20646,N_15111,N_16040);
nor U20647 (N_20647,N_15580,N_15776);
or U20648 (N_20648,N_15034,N_16300);
nand U20649 (N_20649,N_17848,N_17648);
and U20650 (N_20650,N_17319,N_17789);
nor U20651 (N_20651,N_16855,N_15966);
nand U20652 (N_20652,N_17158,N_15308);
or U20653 (N_20653,N_17435,N_16348);
nor U20654 (N_20654,N_16694,N_17349);
and U20655 (N_20655,N_17893,N_17219);
xnor U20656 (N_20656,N_17608,N_15017);
nor U20657 (N_20657,N_15475,N_17868);
or U20658 (N_20658,N_17006,N_17226);
xor U20659 (N_20659,N_15646,N_17105);
xnor U20660 (N_20660,N_15852,N_17980);
and U20661 (N_20661,N_16495,N_15256);
xor U20662 (N_20662,N_15117,N_17458);
or U20663 (N_20663,N_17586,N_16526);
nor U20664 (N_20664,N_17518,N_15541);
xor U20665 (N_20665,N_15531,N_16373);
and U20666 (N_20666,N_17966,N_16125);
or U20667 (N_20667,N_15980,N_15729);
nand U20668 (N_20668,N_17903,N_15673);
nand U20669 (N_20669,N_17880,N_17685);
nand U20670 (N_20670,N_17376,N_16368);
nand U20671 (N_20671,N_17179,N_16497);
or U20672 (N_20672,N_15385,N_16090);
xor U20673 (N_20673,N_16969,N_15290);
nor U20674 (N_20674,N_16538,N_17760);
nor U20675 (N_20675,N_17195,N_15546);
and U20676 (N_20676,N_16068,N_16931);
nor U20677 (N_20677,N_15282,N_15064);
nand U20678 (N_20678,N_16190,N_16621);
nand U20679 (N_20679,N_15006,N_17879);
nor U20680 (N_20680,N_17143,N_16220);
or U20681 (N_20681,N_17208,N_15748);
or U20682 (N_20682,N_16567,N_17155);
nand U20683 (N_20683,N_15326,N_17028);
xor U20684 (N_20684,N_15982,N_15228);
nor U20685 (N_20685,N_17426,N_15865);
xor U20686 (N_20686,N_15549,N_15990);
or U20687 (N_20687,N_17886,N_16039);
nor U20688 (N_20688,N_16736,N_15800);
xnor U20689 (N_20689,N_17202,N_16391);
nor U20690 (N_20690,N_16029,N_17545);
nor U20691 (N_20691,N_17172,N_17460);
and U20692 (N_20692,N_16003,N_15154);
or U20693 (N_20693,N_17713,N_17119);
xnor U20694 (N_20694,N_16851,N_15043);
xor U20695 (N_20695,N_15762,N_15572);
nand U20696 (N_20696,N_15849,N_17777);
or U20697 (N_20697,N_17636,N_17472);
or U20698 (N_20698,N_15610,N_15016);
or U20699 (N_20699,N_17582,N_16599);
nor U20700 (N_20700,N_16069,N_17027);
nor U20701 (N_20701,N_15114,N_17155);
nor U20702 (N_20702,N_17610,N_17305);
nor U20703 (N_20703,N_15958,N_17202);
nand U20704 (N_20704,N_17159,N_15561);
nand U20705 (N_20705,N_16662,N_15731);
nand U20706 (N_20706,N_15796,N_17910);
and U20707 (N_20707,N_16590,N_15310);
xnor U20708 (N_20708,N_17839,N_15909);
nand U20709 (N_20709,N_15692,N_17838);
and U20710 (N_20710,N_15653,N_16629);
and U20711 (N_20711,N_17722,N_15743);
nor U20712 (N_20712,N_15150,N_16203);
nor U20713 (N_20713,N_15205,N_15179);
xor U20714 (N_20714,N_17892,N_16932);
and U20715 (N_20715,N_17271,N_15842);
nand U20716 (N_20716,N_15459,N_17700);
xor U20717 (N_20717,N_15146,N_16845);
or U20718 (N_20718,N_17583,N_15776);
nand U20719 (N_20719,N_16416,N_16501);
xnor U20720 (N_20720,N_15822,N_15385);
nand U20721 (N_20721,N_17589,N_15049);
nor U20722 (N_20722,N_15099,N_16287);
or U20723 (N_20723,N_16368,N_15810);
nand U20724 (N_20724,N_15541,N_17327);
and U20725 (N_20725,N_15650,N_17527);
nor U20726 (N_20726,N_16067,N_15169);
nand U20727 (N_20727,N_17257,N_17201);
nor U20728 (N_20728,N_15404,N_17064);
nor U20729 (N_20729,N_17867,N_16644);
xnor U20730 (N_20730,N_15389,N_15606);
xnor U20731 (N_20731,N_17720,N_17280);
nand U20732 (N_20732,N_16606,N_17414);
nor U20733 (N_20733,N_16493,N_16505);
nand U20734 (N_20734,N_15586,N_15171);
xor U20735 (N_20735,N_17488,N_16135);
or U20736 (N_20736,N_15314,N_17366);
xnor U20737 (N_20737,N_15141,N_17961);
nand U20738 (N_20738,N_17271,N_17044);
or U20739 (N_20739,N_15186,N_15882);
xnor U20740 (N_20740,N_15709,N_16577);
or U20741 (N_20741,N_16194,N_15425);
and U20742 (N_20742,N_17234,N_16534);
or U20743 (N_20743,N_15797,N_17119);
nor U20744 (N_20744,N_16847,N_17307);
nand U20745 (N_20745,N_16996,N_17733);
xor U20746 (N_20746,N_16820,N_15243);
nand U20747 (N_20747,N_17663,N_16338);
nand U20748 (N_20748,N_17584,N_15943);
nor U20749 (N_20749,N_15998,N_17669);
xnor U20750 (N_20750,N_15667,N_17529);
or U20751 (N_20751,N_15053,N_17527);
and U20752 (N_20752,N_16522,N_17603);
nor U20753 (N_20753,N_17748,N_16010);
xor U20754 (N_20754,N_17685,N_15280);
or U20755 (N_20755,N_17952,N_16801);
nand U20756 (N_20756,N_16440,N_15279);
xor U20757 (N_20757,N_17826,N_16024);
nand U20758 (N_20758,N_16293,N_15302);
xor U20759 (N_20759,N_17703,N_17802);
nor U20760 (N_20760,N_15333,N_15368);
xor U20761 (N_20761,N_16486,N_17753);
or U20762 (N_20762,N_16727,N_17498);
nor U20763 (N_20763,N_17805,N_15949);
and U20764 (N_20764,N_15575,N_15695);
nor U20765 (N_20765,N_16173,N_17578);
or U20766 (N_20766,N_15403,N_16972);
xnor U20767 (N_20767,N_16286,N_17488);
or U20768 (N_20768,N_15869,N_15236);
or U20769 (N_20769,N_17978,N_15829);
nand U20770 (N_20770,N_16655,N_15476);
xor U20771 (N_20771,N_17840,N_15081);
or U20772 (N_20772,N_17812,N_16172);
nand U20773 (N_20773,N_17763,N_17592);
or U20774 (N_20774,N_15213,N_16325);
nor U20775 (N_20775,N_15377,N_15429);
nor U20776 (N_20776,N_16130,N_16456);
nor U20777 (N_20777,N_17606,N_17389);
nand U20778 (N_20778,N_15492,N_16525);
xnor U20779 (N_20779,N_16044,N_16375);
and U20780 (N_20780,N_16748,N_15420);
or U20781 (N_20781,N_15410,N_15448);
xnor U20782 (N_20782,N_17387,N_15257);
nor U20783 (N_20783,N_15721,N_15922);
nand U20784 (N_20784,N_17725,N_16132);
xnor U20785 (N_20785,N_16614,N_17962);
nor U20786 (N_20786,N_15406,N_16920);
and U20787 (N_20787,N_15826,N_16185);
nand U20788 (N_20788,N_17653,N_16395);
nand U20789 (N_20789,N_16928,N_15581);
nand U20790 (N_20790,N_15077,N_17452);
xnor U20791 (N_20791,N_17856,N_15247);
nor U20792 (N_20792,N_17597,N_17142);
xnor U20793 (N_20793,N_15971,N_15761);
nand U20794 (N_20794,N_17960,N_16738);
nand U20795 (N_20795,N_17683,N_17178);
and U20796 (N_20796,N_17377,N_16816);
xnor U20797 (N_20797,N_15642,N_15439);
or U20798 (N_20798,N_15491,N_15873);
or U20799 (N_20799,N_17820,N_15911);
and U20800 (N_20800,N_17363,N_15012);
xor U20801 (N_20801,N_15541,N_16635);
nand U20802 (N_20802,N_16990,N_17837);
and U20803 (N_20803,N_16942,N_15236);
xor U20804 (N_20804,N_16671,N_15656);
and U20805 (N_20805,N_15622,N_17089);
and U20806 (N_20806,N_16013,N_17823);
and U20807 (N_20807,N_17875,N_17060);
nand U20808 (N_20808,N_15318,N_17353);
nor U20809 (N_20809,N_17389,N_16888);
xor U20810 (N_20810,N_15173,N_17594);
nor U20811 (N_20811,N_16594,N_16659);
nor U20812 (N_20812,N_16324,N_17220);
nand U20813 (N_20813,N_17477,N_16003);
xnor U20814 (N_20814,N_15397,N_17097);
and U20815 (N_20815,N_16972,N_17758);
nor U20816 (N_20816,N_15366,N_17787);
xnor U20817 (N_20817,N_17818,N_17020);
or U20818 (N_20818,N_15507,N_17746);
nor U20819 (N_20819,N_15290,N_16387);
or U20820 (N_20820,N_16264,N_17298);
nand U20821 (N_20821,N_17308,N_16778);
or U20822 (N_20822,N_16611,N_16497);
nand U20823 (N_20823,N_16271,N_17988);
or U20824 (N_20824,N_17975,N_17540);
nand U20825 (N_20825,N_15755,N_16571);
or U20826 (N_20826,N_15508,N_16868);
nand U20827 (N_20827,N_16846,N_16727);
and U20828 (N_20828,N_17461,N_16261);
and U20829 (N_20829,N_16658,N_17983);
or U20830 (N_20830,N_15405,N_17131);
nor U20831 (N_20831,N_16234,N_17935);
nand U20832 (N_20832,N_15264,N_17891);
and U20833 (N_20833,N_16360,N_15631);
xor U20834 (N_20834,N_16017,N_17928);
xor U20835 (N_20835,N_17169,N_15152);
nand U20836 (N_20836,N_15442,N_15369);
xor U20837 (N_20837,N_16369,N_16662);
and U20838 (N_20838,N_16438,N_15865);
xnor U20839 (N_20839,N_15264,N_16933);
nand U20840 (N_20840,N_15160,N_15384);
or U20841 (N_20841,N_16431,N_17915);
nor U20842 (N_20842,N_15950,N_16361);
xor U20843 (N_20843,N_16431,N_15171);
nand U20844 (N_20844,N_17976,N_17276);
xnor U20845 (N_20845,N_16533,N_15288);
nand U20846 (N_20846,N_17207,N_15035);
and U20847 (N_20847,N_15465,N_16885);
or U20848 (N_20848,N_16392,N_16522);
nand U20849 (N_20849,N_16102,N_16523);
and U20850 (N_20850,N_16033,N_17576);
xor U20851 (N_20851,N_16589,N_15979);
nor U20852 (N_20852,N_16390,N_16650);
or U20853 (N_20853,N_16943,N_17240);
nand U20854 (N_20854,N_17555,N_16896);
xnor U20855 (N_20855,N_16567,N_15259);
nand U20856 (N_20856,N_16535,N_16258);
or U20857 (N_20857,N_17355,N_17656);
or U20858 (N_20858,N_16515,N_17080);
nand U20859 (N_20859,N_15862,N_17645);
nand U20860 (N_20860,N_17739,N_16144);
nor U20861 (N_20861,N_17708,N_16714);
and U20862 (N_20862,N_15072,N_15067);
xor U20863 (N_20863,N_16971,N_16799);
and U20864 (N_20864,N_16283,N_15831);
and U20865 (N_20865,N_16677,N_15789);
xnor U20866 (N_20866,N_15320,N_16567);
or U20867 (N_20867,N_16648,N_16765);
xor U20868 (N_20868,N_17237,N_15404);
nand U20869 (N_20869,N_16560,N_15613);
or U20870 (N_20870,N_15679,N_16985);
or U20871 (N_20871,N_16150,N_16856);
nand U20872 (N_20872,N_17572,N_15167);
nand U20873 (N_20873,N_15077,N_15018);
and U20874 (N_20874,N_15557,N_17006);
xor U20875 (N_20875,N_17256,N_17466);
nand U20876 (N_20876,N_16723,N_17612);
and U20877 (N_20877,N_15698,N_15185);
nand U20878 (N_20878,N_16633,N_16950);
or U20879 (N_20879,N_17012,N_17849);
and U20880 (N_20880,N_15677,N_15291);
or U20881 (N_20881,N_16642,N_16994);
xor U20882 (N_20882,N_15865,N_15881);
nor U20883 (N_20883,N_16387,N_15998);
xor U20884 (N_20884,N_17282,N_17713);
xnor U20885 (N_20885,N_17493,N_17370);
nor U20886 (N_20886,N_16557,N_17829);
nand U20887 (N_20887,N_17824,N_15383);
or U20888 (N_20888,N_17544,N_17576);
or U20889 (N_20889,N_16521,N_16595);
xnor U20890 (N_20890,N_15135,N_15368);
or U20891 (N_20891,N_15926,N_15860);
and U20892 (N_20892,N_15701,N_15275);
nand U20893 (N_20893,N_15534,N_17563);
or U20894 (N_20894,N_17245,N_17042);
xor U20895 (N_20895,N_17397,N_16059);
nand U20896 (N_20896,N_17071,N_17053);
nor U20897 (N_20897,N_17441,N_16973);
and U20898 (N_20898,N_17347,N_15452);
and U20899 (N_20899,N_15609,N_16126);
nand U20900 (N_20900,N_15619,N_16414);
nor U20901 (N_20901,N_17334,N_16725);
nand U20902 (N_20902,N_15310,N_17730);
nor U20903 (N_20903,N_17515,N_15882);
and U20904 (N_20904,N_17637,N_16494);
nand U20905 (N_20905,N_15435,N_17104);
or U20906 (N_20906,N_15937,N_16407);
nand U20907 (N_20907,N_15777,N_16531);
nand U20908 (N_20908,N_16906,N_15008);
or U20909 (N_20909,N_17426,N_15904);
xnor U20910 (N_20910,N_15883,N_15674);
nand U20911 (N_20911,N_15809,N_15430);
xor U20912 (N_20912,N_17362,N_16337);
or U20913 (N_20913,N_15267,N_15655);
nand U20914 (N_20914,N_17848,N_17023);
or U20915 (N_20915,N_15626,N_17899);
or U20916 (N_20916,N_15864,N_17836);
or U20917 (N_20917,N_15252,N_16954);
xor U20918 (N_20918,N_17515,N_16714);
nand U20919 (N_20919,N_16998,N_17778);
and U20920 (N_20920,N_17989,N_16577);
xor U20921 (N_20921,N_16781,N_16590);
nor U20922 (N_20922,N_16053,N_16198);
nand U20923 (N_20923,N_17642,N_16668);
and U20924 (N_20924,N_15733,N_15291);
nor U20925 (N_20925,N_16062,N_16076);
nor U20926 (N_20926,N_17811,N_16990);
and U20927 (N_20927,N_16780,N_16743);
nand U20928 (N_20928,N_15908,N_15598);
nor U20929 (N_20929,N_15919,N_16564);
xor U20930 (N_20930,N_16365,N_17790);
and U20931 (N_20931,N_17482,N_17226);
or U20932 (N_20932,N_15939,N_17201);
xor U20933 (N_20933,N_15068,N_16785);
xnor U20934 (N_20934,N_16185,N_16451);
and U20935 (N_20935,N_17647,N_15906);
or U20936 (N_20936,N_15403,N_15733);
nand U20937 (N_20937,N_17722,N_15633);
xnor U20938 (N_20938,N_16771,N_17381);
nand U20939 (N_20939,N_16543,N_17190);
nor U20940 (N_20940,N_15278,N_16998);
xnor U20941 (N_20941,N_17197,N_16089);
nor U20942 (N_20942,N_15430,N_16753);
and U20943 (N_20943,N_16043,N_17177);
nor U20944 (N_20944,N_16000,N_15859);
xnor U20945 (N_20945,N_16470,N_15196);
and U20946 (N_20946,N_16942,N_15628);
nand U20947 (N_20947,N_15774,N_16911);
nand U20948 (N_20948,N_17078,N_16937);
nor U20949 (N_20949,N_16196,N_17020);
and U20950 (N_20950,N_15564,N_17807);
or U20951 (N_20951,N_15345,N_17949);
nor U20952 (N_20952,N_17744,N_15327);
nand U20953 (N_20953,N_15928,N_17897);
or U20954 (N_20954,N_15198,N_15793);
or U20955 (N_20955,N_17655,N_16924);
nand U20956 (N_20956,N_16730,N_17201);
nand U20957 (N_20957,N_17824,N_15232);
nand U20958 (N_20958,N_17380,N_15037);
or U20959 (N_20959,N_17284,N_15020);
and U20960 (N_20960,N_15941,N_16555);
nand U20961 (N_20961,N_16134,N_16276);
xor U20962 (N_20962,N_15139,N_16161);
nand U20963 (N_20963,N_17393,N_15509);
nand U20964 (N_20964,N_17517,N_15623);
xnor U20965 (N_20965,N_16110,N_17914);
and U20966 (N_20966,N_17989,N_17164);
nand U20967 (N_20967,N_15328,N_15258);
nor U20968 (N_20968,N_15971,N_15213);
and U20969 (N_20969,N_15470,N_15635);
xor U20970 (N_20970,N_15610,N_16242);
and U20971 (N_20971,N_16756,N_17485);
nand U20972 (N_20972,N_16162,N_16431);
nand U20973 (N_20973,N_15674,N_15061);
and U20974 (N_20974,N_15711,N_16355);
or U20975 (N_20975,N_16696,N_17059);
nor U20976 (N_20976,N_17071,N_16742);
nor U20977 (N_20977,N_15203,N_16759);
nand U20978 (N_20978,N_17592,N_16433);
nand U20979 (N_20979,N_15884,N_15310);
or U20980 (N_20980,N_16484,N_16201);
nand U20981 (N_20981,N_16739,N_15687);
xor U20982 (N_20982,N_16116,N_17006);
and U20983 (N_20983,N_15624,N_16806);
nand U20984 (N_20984,N_15103,N_17655);
xor U20985 (N_20985,N_15461,N_15426);
nor U20986 (N_20986,N_16310,N_16288);
and U20987 (N_20987,N_17477,N_17381);
or U20988 (N_20988,N_15018,N_17176);
xor U20989 (N_20989,N_15384,N_16770);
xnor U20990 (N_20990,N_16574,N_15984);
and U20991 (N_20991,N_17185,N_16569);
nand U20992 (N_20992,N_17012,N_15463);
nor U20993 (N_20993,N_15759,N_15592);
xor U20994 (N_20994,N_17202,N_16431);
xor U20995 (N_20995,N_17323,N_16281);
nand U20996 (N_20996,N_16438,N_15924);
nor U20997 (N_20997,N_15012,N_16893);
or U20998 (N_20998,N_16739,N_17779);
or U20999 (N_20999,N_16609,N_17993);
xor U21000 (N_21000,N_20041,N_20149);
nor U21001 (N_21001,N_18860,N_19268);
nor U21002 (N_21002,N_19617,N_20960);
or U21003 (N_21003,N_19272,N_20166);
nor U21004 (N_21004,N_19912,N_18850);
and U21005 (N_21005,N_19071,N_19868);
nand U21006 (N_21006,N_20984,N_20843);
nand U21007 (N_21007,N_20785,N_19765);
and U21008 (N_21008,N_19607,N_18011);
nand U21009 (N_21009,N_18483,N_19081);
nand U21010 (N_21010,N_20205,N_19914);
nor U21011 (N_21011,N_19286,N_18665);
nor U21012 (N_21012,N_18197,N_20179);
xor U21013 (N_21013,N_19861,N_20493);
nand U21014 (N_21014,N_20589,N_18061);
or U21015 (N_21015,N_19599,N_20020);
xnor U21016 (N_21016,N_19988,N_20007);
or U21017 (N_21017,N_18682,N_18005);
and U21018 (N_21018,N_18637,N_19485);
nor U21019 (N_21019,N_18644,N_19123);
nand U21020 (N_21020,N_19616,N_18864);
or U21021 (N_21021,N_18835,N_18287);
or U21022 (N_21022,N_19828,N_19696);
xor U21023 (N_21023,N_20518,N_19686);
nand U21024 (N_21024,N_20686,N_20378);
or U21025 (N_21025,N_18261,N_18757);
nand U21026 (N_21026,N_18063,N_20894);
xor U21027 (N_21027,N_18456,N_18609);
or U21028 (N_21028,N_19254,N_18723);
nand U21029 (N_21029,N_20082,N_19243);
nand U21030 (N_21030,N_19595,N_18398);
nand U21031 (N_21031,N_20510,N_19945);
nand U21032 (N_21032,N_18461,N_18085);
or U21033 (N_21033,N_18927,N_18848);
and U21034 (N_21034,N_18556,N_19074);
or U21035 (N_21035,N_20612,N_19288);
nand U21036 (N_21036,N_18250,N_19966);
nand U21037 (N_21037,N_19682,N_20327);
or U21038 (N_21038,N_20426,N_20946);
nor U21039 (N_21039,N_18341,N_18970);
and U21040 (N_21040,N_19421,N_19709);
nand U21041 (N_21041,N_19880,N_20341);
xnor U21042 (N_21042,N_20629,N_19721);
xnor U21043 (N_21043,N_18877,N_18078);
or U21044 (N_21044,N_18529,N_19805);
nand U21045 (N_21045,N_20116,N_18347);
and U21046 (N_21046,N_18954,N_19314);
xnor U21047 (N_21047,N_18965,N_20918);
nor U21048 (N_21048,N_19655,N_18696);
xor U21049 (N_21049,N_20316,N_20927);
and U21050 (N_21050,N_20942,N_19598);
or U21051 (N_21051,N_18445,N_18620);
nor U21052 (N_21052,N_20321,N_18365);
xnor U21053 (N_21053,N_19487,N_18091);
or U21054 (N_21054,N_19725,N_18630);
nand U21055 (N_21055,N_18361,N_20738);
xnor U21056 (N_21056,N_18929,N_18565);
and U21057 (N_21057,N_18714,N_19163);
and U21058 (N_21058,N_20030,N_19813);
and U21059 (N_21059,N_19859,N_18245);
or U21060 (N_21060,N_18298,N_18258);
nor U21061 (N_21061,N_20873,N_19028);
or U21062 (N_21062,N_18564,N_19716);
nor U21063 (N_21063,N_19482,N_20617);
or U21064 (N_21064,N_19306,N_20988);
and U21065 (N_21065,N_18832,N_18846);
nor U21066 (N_21066,N_18519,N_19582);
or U21067 (N_21067,N_18499,N_20161);
or U21068 (N_21068,N_20641,N_18136);
xnor U21069 (N_21069,N_20133,N_18616);
or U21070 (N_21070,N_18304,N_20837);
and U21071 (N_21071,N_20303,N_19559);
or U21072 (N_21072,N_18058,N_19791);
xor U21073 (N_21073,N_19405,N_20292);
or U21074 (N_21074,N_19006,N_19415);
or U21075 (N_21075,N_19430,N_20648);
or U21076 (N_21076,N_19501,N_19674);
and U21077 (N_21077,N_20394,N_20382);
nor U21078 (N_21078,N_18133,N_20753);
or U21079 (N_21079,N_19670,N_20369);
xnor U21080 (N_21080,N_19905,N_19741);
nor U21081 (N_21081,N_18415,N_19798);
nand U21082 (N_21082,N_20143,N_19414);
or U21083 (N_21083,N_19992,N_20035);
nand U21084 (N_21084,N_18703,N_19833);
nand U21085 (N_21085,N_20729,N_20485);
nor U21086 (N_21086,N_19503,N_19646);
nor U21087 (N_21087,N_19207,N_18704);
xor U21088 (N_21088,N_18976,N_18613);
xnor U21089 (N_21089,N_18962,N_18791);
nor U21090 (N_21090,N_19338,N_18656);
and U21091 (N_21091,N_20293,N_19358);
nand U21092 (N_21092,N_19838,N_18272);
nor U21093 (N_21093,N_20836,N_20553);
xor U21094 (N_21094,N_19809,N_18685);
nand U21095 (N_21095,N_19799,N_18301);
xor U21096 (N_21096,N_19139,N_19939);
and U21097 (N_21097,N_20416,N_18026);
nor U21098 (N_21098,N_18165,N_20377);
and U21099 (N_21099,N_19863,N_19279);
xnor U21100 (N_21100,N_18467,N_20905);
and U21101 (N_21101,N_20447,N_19916);
or U21102 (N_21102,N_18554,N_20379);
and U21103 (N_21103,N_20135,N_18025);
nand U21104 (N_21104,N_20242,N_19223);
nand U21105 (N_21105,N_18442,N_19715);
or U21106 (N_21106,N_18469,N_18568);
xor U21107 (N_21107,N_20492,N_20432);
and U21108 (N_21108,N_18225,N_19017);
xor U21109 (N_21109,N_18514,N_19151);
nor U21110 (N_21110,N_20311,N_20900);
nor U21111 (N_21111,N_20576,N_20345);
and U21112 (N_21112,N_20401,N_19416);
or U21113 (N_21113,N_20839,N_18366);
nand U21114 (N_21114,N_20326,N_19604);
or U21115 (N_21115,N_20801,N_19649);
nand U21116 (N_21116,N_19463,N_20779);
nand U21117 (N_21117,N_18115,N_19219);
nor U21118 (N_21118,N_18187,N_19312);
nand U21119 (N_21119,N_20031,N_18198);
xor U21120 (N_21120,N_19236,N_19862);
or U21121 (N_21121,N_18614,N_18646);
xnor U21122 (N_21122,N_20328,N_18649);
xor U21123 (N_21123,N_19736,N_18060);
nor U21124 (N_21124,N_18847,N_19909);
or U21125 (N_21125,N_18351,N_20909);
nor U21126 (N_21126,N_19450,N_19099);
xor U21127 (N_21127,N_20757,N_19057);
nor U21128 (N_21128,N_18434,N_20340);
nor U21129 (N_21129,N_19845,N_20430);
and U21130 (N_21130,N_19636,N_18840);
xor U21131 (N_21131,N_19987,N_20564);
nand U21132 (N_21132,N_19520,N_18804);
or U21133 (N_21133,N_20540,N_20986);
or U21134 (N_21134,N_20777,N_20809);
xor U21135 (N_21135,N_18371,N_20195);
nor U21136 (N_21136,N_18561,N_18511);
nand U21137 (N_21137,N_19156,N_19882);
nor U21138 (N_21138,N_18578,N_18606);
and U21139 (N_21139,N_20145,N_19082);
xor U21140 (N_21140,N_20971,N_18913);
xnor U21141 (N_21141,N_19129,N_20818);
nor U21142 (N_21142,N_18596,N_18159);
xnor U21143 (N_21143,N_19318,N_18701);
or U21144 (N_21144,N_19227,N_19049);
xor U21145 (N_21145,N_20176,N_19937);
nand U21146 (N_21146,N_18183,N_18244);
and U21147 (N_21147,N_18873,N_20749);
xor U21148 (N_21148,N_18503,N_20804);
and U21149 (N_21149,N_18688,N_18633);
nor U21150 (N_21150,N_19294,N_18032);
and U21151 (N_21151,N_18824,N_19737);
xor U21152 (N_21152,N_18935,N_19407);
nor U21153 (N_21153,N_20286,N_19111);
or U21154 (N_21154,N_19879,N_20395);
nor U21155 (N_21155,N_20998,N_20004);
nand U21156 (N_21156,N_19618,N_18849);
nand U21157 (N_21157,N_19730,N_20289);
and U21158 (N_21158,N_20167,N_18892);
nand U21159 (N_21159,N_20055,N_20719);
nand U21160 (N_21160,N_18755,N_20938);
and U21161 (N_21161,N_18132,N_18774);
and U21162 (N_21162,N_18908,N_18331);
or U21163 (N_21163,N_18404,N_18672);
or U21164 (N_21164,N_20137,N_20500);
nand U21165 (N_21165,N_18653,N_19775);
and U21166 (N_21166,N_18342,N_19735);
nand U21167 (N_21167,N_18584,N_20476);
and U21168 (N_21168,N_19353,N_20951);
nor U21169 (N_21169,N_19785,N_19275);
xor U21170 (N_21170,N_20561,N_19213);
nand U21171 (N_21171,N_20472,N_20989);
nand U21172 (N_21172,N_18603,N_19391);
and U21173 (N_21173,N_19989,N_18731);
and U21174 (N_21174,N_18277,N_19533);
xnor U21175 (N_21175,N_20634,N_19110);
nand U21176 (N_21176,N_18255,N_20644);
nand U21177 (N_21177,N_20953,N_19424);
nor U21178 (N_21178,N_20978,N_18880);
xnor U21179 (N_21179,N_19792,N_20064);
xor U21180 (N_21180,N_18080,N_18153);
nand U21181 (N_21181,N_18619,N_19509);
nor U21182 (N_21182,N_18195,N_18724);
and U21183 (N_21183,N_18409,N_19570);
nor U21184 (N_21184,N_20872,N_19027);
nand U21185 (N_21185,N_18113,N_19278);
nor U21186 (N_21186,N_20467,N_19085);
nand U21187 (N_21187,N_20233,N_18819);
nor U21188 (N_21188,N_19147,N_20755);
and U21189 (N_21189,N_18390,N_19297);
nor U21190 (N_21190,N_20353,N_20083);
xor U21191 (N_21191,N_18585,N_20615);
nor U21192 (N_21192,N_20936,N_19778);
nand U21193 (N_21193,N_20052,N_18911);
and U21194 (N_21194,N_19892,N_19619);
nand U21195 (N_21195,N_20387,N_20619);
or U21196 (N_21196,N_19355,N_19269);
nand U21197 (N_21197,N_19201,N_19708);
xnor U21198 (N_21198,N_19927,N_20402);
or U21199 (N_21199,N_18505,N_20040);
xor U21200 (N_21200,N_19155,N_20763);
and U21201 (N_21201,N_18781,N_20764);
nand U21202 (N_21202,N_19036,N_19853);
nor U21203 (N_21203,N_19105,N_18745);
nand U21204 (N_21204,N_18681,N_18312);
xor U21205 (N_21205,N_18344,N_18858);
xor U21206 (N_21206,N_18383,N_18663);
nor U21207 (N_21207,N_20603,N_18715);
and U21208 (N_21208,N_20527,N_18795);
nor U21209 (N_21209,N_18050,N_20390);
or U21210 (N_21210,N_20670,N_19499);
nor U21211 (N_21211,N_20868,N_18833);
nor U21212 (N_21212,N_19968,N_20660);
nor U21213 (N_21213,N_18702,N_20788);
nor U21214 (N_21214,N_20489,N_20637);
or U21215 (N_21215,N_19982,N_18157);
or U21216 (N_21216,N_20294,N_18140);
nor U21217 (N_21217,N_18161,N_18462);
nor U21218 (N_21218,N_20618,N_18203);
nor U21219 (N_21219,N_18654,N_18604);
and U21220 (N_21220,N_19724,N_18112);
xor U21221 (N_21221,N_19336,N_18303);
and U21222 (N_21222,N_20044,N_19621);
and U21223 (N_21223,N_20955,N_19376);
nor U21224 (N_21224,N_20972,N_20783);
or U21225 (N_21225,N_18362,N_18018);
and U21226 (N_21226,N_20663,N_19045);
and U21227 (N_21227,N_20696,N_18540);
and U21228 (N_21228,N_20762,N_19934);
nand U21229 (N_21229,N_18273,N_18088);
and U21230 (N_21230,N_19656,N_19876);
nor U21231 (N_21231,N_20099,N_18925);
nor U21232 (N_21232,N_19133,N_20970);
nor U21233 (N_21233,N_19034,N_18662);
xor U21234 (N_21234,N_18176,N_19844);
nor U21235 (N_21235,N_18575,N_18089);
nand U21236 (N_21236,N_18983,N_18215);
xnor U21237 (N_21237,N_18974,N_19854);
nand U21238 (N_21238,N_19544,N_18270);
xnor U21239 (N_21239,N_19667,N_18611);
nand U21240 (N_21240,N_20354,N_19335);
and U21241 (N_21241,N_18170,N_18697);
nor U21242 (N_21242,N_19320,N_18266);
and U21243 (N_21243,N_20053,N_18555);
and U21244 (N_21244,N_20620,N_18259);
nand U21245 (N_21245,N_20019,N_20943);
and U21246 (N_21246,N_18436,N_19368);
nor U21247 (N_21247,N_19552,N_20334);
xor U21248 (N_21248,N_20468,N_20844);
nor U21249 (N_21249,N_19007,N_19583);
xor U21250 (N_21250,N_19115,N_18571);
xnor U21251 (N_21251,N_18493,N_19168);
and U21252 (N_21252,N_19596,N_20814);
or U21253 (N_21253,N_19098,N_18508);
or U21254 (N_21254,N_19182,N_19812);
or U21255 (N_21255,N_19238,N_20123);
or U21256 (N_21256,N_20735,N_20203);
xor U21257 (N_21257,N_18979,N_20089);
nor U21258 (N_21258,N_20305,N_20084);
xnor U21259 (N_21259,N_20535,N_19193);
and U21260 (N_21260,N_19712,N_18049);
and U21261 (N_21261,N_18968,N_18098);
or U21262 (N_21262,N_18126,N_18453);
nand U21263 (N_21263,N_19210,N_20559);
xor U21264 (N_21264,N_20556,N_19829);
nor U21265 (N_21265,N_19114,N_20445);
nor U21266 (N_21266,N_18352,N_18816);
nor U21267 (N_21267,N_20924,N_18617);
nand U21268 (N_21268,N_20758,N_20086);
or U21269 (N_21269,N_18507,N_19050);
nor U21270 (N_21270,N_20833,N_20528);
xor U21271 (N_21271,N_19642,N_20995);
nor U21272 (N_21272,N_20318,N_20156);
nand U21273 (N_21273,N_19153,N_20743);
or U21274 (N_21274,N_19920,N_18125);
xnor U21275 (N_21275,N_20679,N_19032);
or U21276 (N_21276,N_18015,N_18713);
or U21277 (N_21277,N_19240,N_18057);
or U21278 (N_21278,N_20707,N_20555);
xor U21279 (N_21279,N_20144,N_18392);
nor U21280 (N_21280,N_18315,N_20636);
nand U21281 (N_21281,N_18317,N_20787);
nor U21282 (N_21282,N_20330,N_19169);
nor U21283 (N_21283,N_18275,N_19116);
and U21284 (N_21284,N_19466,N_20794);
xor U21285 (N_21285,N_20093,N_18865);
and U21286 (N_21286,N_20916,N_19823);
nand U21287 (N_21287,N_18587,N_19332);
and U21288 (N_21288,N_19756,N_20593);
nor U21289 (N_21289,N_19422,N_20079);
nor U21290 (N_21290,N_19867,N_19048);
and U21291 (N_21291,N_18921,N_19706);
xnor U21292 (N_21292,N_20880,N_19490);
xnor U21293 (N_21293,N_19979,N_18875);
nand U21294 (N_21294,N_20198,N_20652);
nor U21295 (N_21295,N_18010,N_19200);
or U21296 (N_21296,N_20874,N_19342);
nand U21297 (N_21297,N_18053,N_19692);
xor U21298 (N_21298,N_18978,N_20542);
nor U21299 (N_21299,N_19797,N_18894);
and U21300 (N_21300,N_20616,N_18280);
nor U21301 (N_21301,N_19299,N_18586);
xor U21302 (N_21302,N_18432,N_19751);
or U21303 (N_21303,N_20845,N_19013);
or U21304 (N_21304,N_20599,N_19963);
xor U21305 (N_21305,N_18999,N_18118);
xor U21306 (N_21306,N_20209,N_20152);
or U21307 (N_21307,N_18289,N_20550);
nand U21308 (N_21308,N_18830,N_19431);
nand U21309 (N_21309,N_19390,N_20388);
or U21310 (N_21310,N_18727,N_20338);
or U21311 (N_21311,N_18168,N_20012);
nand U21312 (N_21312,N_19203,N_18042);
or U21313 (N_21313,N_18355,N_19280);
xnor U21314 (N_21314,N_18471,N_18881);
nor U21315 (N_21315,N_18635,N_20892);
nand U21316 (N_21316,N_19516,N_20739);
xor U21317 (N_21317,N_20147,N_20858);
nand U21318 (N_21318,N_18815,N_19410);
and U21319 (N_21319,N_18583,N_19883);
or U21320 (N_21320,N_18156,N_20002);
xor U21321 (N_21321,N_18759,N_20677);
or U21322 (N_21322,N_20852,N_19825);
and U21323 (N_21323,N_18201,N_18147);
xor U21324 (N_21324,N_20813,N_19075);
or U21325 (N_21325,N_20054,N_19576);
nor U21326 (N_21326,N_18236,N_18484);
xnor U21327 (N_21327,N_20760,N_19317);
nor U21328 (N_21328,N_18749,N_19150);
nor U21329 (N_21329,N_19540,N_19580);
nand U21330 (N_21330,N_18207,N_19023);
and U21331 (N_21331,N_19371,N_18320);
or U21332 (N_21332,N_19525,N_18799);
and U21333 (N_21333,N_18354,N_20419);
or U21334 (N_21334,N_20239,N_20132);
nand U21335 (N_21335,N_18420,N_20141);
nor U21336 (N_21336,N_20462,N_19250);
xor U21337 (N_21337,N_20796,N_19707);
nand U21338 (N_21338,N_18878,N_20568);
and U21339 (N_21339,N_20992,N_20119);
or U21340 (N_21340,N_18631,N_19970);
nor U21341 (N_21341,N_18497,N_19330);
or U21342 (N_21342,N_20473,N_20185);
nor U21343 (N_21343,N_20904,N_19840);
nand U21344 (N_21344,N_20827,N_18845);
nand U21345 (N_21345,N_20952,N_18648);
or U21346 (N_21346,N_18706,N_19634);
or U21347 (N_21347,N_18326,N_20213);
xnor U21348 (N_21348,N_18691,N_18668);
or U21349 (N_21349,N_18732,N_18457);
or U21350 (N_21350,N_20422,N_19900);
xnor U21351 (N_21351,N_19820,N_19745);
xor U21352 (N_21352,N_19774,N_18933);
nand U21353 (N_21353,N_18944,N_18750);
or U21354 (N_21354,N_19185,N_19896);
nor U21355 (N_21355,N_19484,N_20165);
and U21356 (N_21356,N_20940,N_19690);
nand U21357 (N_21357,N_18693,N_19697);
nor U21358 (N_21358,N_18155,N_18044);
nor U21359 (N_21359,N_19729,N_19020);
nor U21360 (N_21360,N_20247,N_20966);
and U21361 (N_21361,N_19313,N_18523);
nor U21362 (N_21362,N_18076,N_20680);
or U21363 (N_21363,N_20668,N_20003);
nor U21364 (N_21364,N_20057,N_20291);
nand U21365 (N_21365,N_19538,N_19472);
or U21366 (N_21366,N_18389,N_20898);
xor U21367 (N_21367,N_18059,N_20786);
and U21368 (N_21368,N_20333,N_18370);
or U21369 (N_21369,N_20684,N_20182);
xor U21370 (N_21370,N_20375,N_18741);
xnor U21371 (N_21371,N_18676,N_18369);
nor U21372 (N_21372,N_18622,N_19392);
nor U21373 (N_21373,N_18671,N_20773);
or U21374 (N_21374,N_20106,N_18117);
nand U21375 (N_21375,N_18422,N_20346);
xnor U21376 (N_21376,N_18570,N_18910);
nand U21377 (N_21377,N_20253,N_18019);
or U21378 (N_21378,N_19753,N_18577);
xnor U21379 (N_21379,N_19009,N_18557);
and U21380 (N_21380,N_19884,N_20150);
nand U21381 (N_21381,N_20162,N_19467);
nand U21382 (N_21382,N_19901,N_19800);
and U21383 (N_21383,N_18281,N_20180);
nor U21384 (N_21384,N_18391,N_18516);
nand U21385 (N_21385,N_19964,N_18230);
nor U21386 (N_21386,N_18145,N_20921);
nor U21387 (N_21387,N_18437,N_19244);
nand U21388 (N_21388,N_20347,N_19594);
or U21389 (N_21389,N_19003,N_20626);
xor U21390 (N_21390,N_20526,N_18629);
and U21391 (N_21391,N_19388,N_20155);
or U21392 (N_21392,N_20479,N_18162);
or U21393 (N_21393,N_20315,N_18859);
and U21394 (N_21394,N_19241,N_20931);
nand U21395 (N_21395,N_20826,N_18380);
nand U21396 (N_21396,N_19569,N_19993);
or U21397 (N_21397,N_20163,N_18382);
and U21398 (N_21398,N_20077,N_18844);
or U21399 (N_21399,N_20627,N_18890);
xnor U21400 (N_21400,N_20391,N_18108);
and U21401 (N_21401,N_18101,N_19766);
nand U21402 (N_21402,N_19852,N_18756);
nor U21403 (N_21403,N_20359,N_18924);
nand U21404 (N_21404,N_18659,N_19929);
nor U21405 (N_21405,N_20120,N_20243);
and U21406 (N_21406,N_19031,N_18097);
xor U21407 (N_21407,N_19149,N_18995);
nand U21408 (N_21408,N_19319,N_20323);
or U21409 (N_21409,N_19700,N_19586);
and U21410 (N_21410,N_20234,N_18135);
or U21411 (N_21411,N_19597,N_19941);
and U21412 (N_21412,N_18051,N_18222);
or U21413 (N_21413,N_18348,N_19850);
and U21414 (N_21414,N_18610,N_20950);
and U21415 (N_21415,N_20797,N_20199);
nor U21416 (N_21416,N_20097,N_20699);
and U21417 (N_21417,N_18430,N_18683);
or U21418 (N_21418,N_18917,N_20562);
nand U21419 (N_21419,N_18022,N_18185);
and U21420 (N_21420,N_20870,N_19659);
nand U21421 (N_21421,N_20557,N_18034);
or U21422 (N_21422,N_18936,N_19780);
nand U21423 (N_21423,N_19531,N_20171);
xor U21424 (N_21424,N_18541,N_20320);
and U21425 (N_21425,N_18385,N_18651);
nor U21426 (N_21426,N_18975,N_18695);
or U21427 (N_21427,N_18504,N_20611);
or U21428 (N_21428,N_19784,N_19301);
or U21429 (N_21429,N_19274,N_18216);
nor U21430 (N_21430,N_20081,N_18188);
or U21431 (N_21431,N_18137,N_19625);
xor U21432 (N_21432,N_19441,N_18454);
nand U21433 (N_21433,N_19107,N_20486);
and U21434 (N_21434,N_20228,N_18127);
nand U21435 (N_21435,N_18014,N_20256);
nand U21436 (N_21436,N_19505,N_20575);
and U21437 (N_21437,N_18283,N_19305);
xnor U21438 (N_21438,N_19551,N_20733);
nand U21439 (N_21439,N_18253,N_20765);
or U21440 (N_21440,N_19906,N_19526);
xor U21441 (N_21441,N_20703,N_19806);
xor U21442 (N_21442,N_19258,N_19308);
nand U21443 (N_21443,N_20768,N_20574);
xnor U21444 (N_21444,N_18397,N_18803);
nand U21445 (N_21445,N_20584,N_18942);
nand U21446 (N_21446,N_20262,N_18861);
nor U21447 (N_21447,N_18334,N_19041);
nor U21448 (N_21448,N_20704,N_18670);
nor U21449 (N_21449,N_18086,N_19389);
or U21450 (N_21450,N_18521,N_19412);
nor U21451 (N_21451,N_20306,N_19518);
or U21452 (N_21452,N_18916,N_18870);
and U21453 (N_21453,N_19340,N_18090);
and U21454 (N_21454,N_20717,N_19030);
xnor U21455 (N_21455,N_19871,N_18869);
and U21456 (N_21456,N_19237,N_19652);
xor U21457 (N_21457,N_19787,N_18152);
or U21458 (N_21458,N_19865,N_20937);
xnor U21459 (N_21459,N_20360,N_20424);
or U21460 (N_21460,N_20811,N_18898);
nand U21461 (N_21461,N_20245,N_19606);
or U21462 (N_21462,N_20109,N_19470);
nor U21463 (N_21463,N_20543,N_19581);
nor U21464 (N_21464,N_20560,N_19816);
nand U21465 (N_21465,N_19125,N_20159);
xnor U21466 (N_21466,N_18186,N_19888);
or U21467 (N_21467,N_18307,N_19015);
or U21468 (N_21468,N_19413,N_18421);
nor U21469 (N_21469,N_19315,N_19411);
and U21470 (N_21470,N_19921,N_18003);
xnor U21471 (N_21471,N_19681,N_19984);
nand U21472 (N_21472,N_19016,N_19949);
or U21473 (N_21473,N_18311,N_19327);
or U21474 (N_21474,N_19091,N_20495);
nand U21475 (N_21475,N_20647,N_20533);
nor U21476 (N_21476,N_19356,N_19891);
nor U21477 (N_21477,N_19383,N_20314);
nor U21478 (N_21478,N_20525,N_18728);
nand U21479 (N_21479,N_20255,N_19699);
and U21480 (N_21480,N_18753,N_19624);
or U21481 (N_21481,N_18411,N_19764);
nor U21482 (N_21482,N_18364,N_20687);
xor U21483 (N_21483,N_18863,N_20349);
nand U21484 (N_21484,N_18031,N_20581);
or U21485 (N_21485,N_18533,N_20929);
and U21486 (N_21486,N_18444,N_19205);
nor U21487 (N_21487,N_19858,N_18600);
nor U21488 (N_21488,N_19191,N_19456);
and U21489 (N_21489,N_20269,N_19029);
or U21490 (N_21490,N_19423,N_19478);
and U21491 (N_21491,N_20941,N_20499);
or U21492 (N_21492,N_20189,N_20522);
xor U21493 (N_21493,N_19761,N_19046);
and U21494 (N_21494,N_19418,N_19396);
nand U21495 (N_21495,N_19384,N_19465);
and U21496 (N_21496,N_20958,N_19851);
nor U21497 (N_21497,N_18268,N_20018);
and U21498 (N_21498,N_20871,N_20795);
nand U21499 (N_21499,N_18820,N_20678);
and U21500 (N_21500,N_19821,N_20418);
nand U21501 (N_21501,N_20903,N_19469);
and U21502 (N_21502,N_19372,N_19255);
nor U21503 (N_21503,N_20780,N_19277);
nor U21504 (N_21504,N_19374,N_19924);
nor U21505 (N_21505,N_20830,N_20112);
xnor U21506 (N_21506,N_20945,N_19628);
nand U21507 (N_21507,N_20625,N_18257);
and U21508 (N_21508,N_19794,N_19047);
nand U21509 (N_21509,N_19839,N_18491);
xor U21510 (N_21510,N_18807,N_19186);
xor U21511 (N_21511,N_19287,N_19873);
or U21512 (N_21512,N_18329,N_19425);
nor U21513 (N_21513,N_18180,N_19452);
and U21514 (N_21514,N_20290,N_20480);
nor U21515 (N_21515,N_19662,N_18017);
nand U21516 (N_21516,N_20973,N_20477);
or U21517 (N_21517,N_20383,N_19980);
and U21518 (N_21518,N_20569,N_18544);
nand U21519 (N_21519,N_20734,N_19251);
or U21520 (N_21520,N_18582,N_20798);
xnor U21521 (N_21521,N_18416,N_18915);
and U21522 (N_21522,N_18747,N_20807);
or U21523 (N_21523,N_19698,N_19398);
xor U21524 (N_21524,N_19995,N_18477);
or U21525 (N_21525,N_20235,N_19807);
and U21526 (N_21526,N_19429,N_20708);
nor U21527 (N_21527,N_19627,N_20997);
nor U21528 (N_21528,N_19519,N_18641);
nor U21529 (N_21529,N_20170,N_20690);
nor U21530 (N_21530,N_18573,N_20565);
xnor U21531 (N_21531,N_20279,N_20329);
nor U21532 (N_21532,N_18752,N_20299);
nor U21533 (N_21533,N_20767,N_18906);
xor U21534 (N_21534,N_19510,N_19677);
and U21535 (N_21535,N_18350,N_20563);
or U21536 (N_21536,N_18427,N_20138);
nor U21537 (N_21537,N_19897,N_20014);
xor U21538 (N_21538,N_18036,N_20091);
and U21539 (N_21539,N_19119,N_20036);
xor U21540 (N_21540,N_19864,N_18475);
or U21541 (N_21541,N_19890,N_18530);
and U21542 (N_21542,N_20805,N_19898);
nand U21543 (N_21543,N_20348,N_20076);
nor U21544 (N_21544,N_20598,N_20016);
nor U21545 (N_21545,N_19904,N_19530);
and U21546 (N_21546,N_20990,N_20173);
nor U21547 (N_21547,N_19922,N_18426);
and U21548 (N_21548,N_20066,N_18992);
or U21549 (N_21549,N_20406,N_19361);
nand U21550 (N_21550,N_18551,N_18856);
xnor U21551 (N_21551,N_19399,N_19947);
nand U21552 (N_21552,N_18020,N_19348);
or U21553 (N_21553,N_19959,N_20539);
xor U21554 (N_21554,N_18282,N_19506);
xnor U21555 (N_21555,N_19008,N_19060);
and U21556 (N_21556,N_19121,N_20840);
nand U21557 (N_21557,N_18743,N_19488);
and U21558 (N_21558,N_19334,N_19063);
nor U21559 (N_21559,N_18590,N_19276);
and U21560 (N_21560,N_19592,N_18041);
nand U21561 (N_21561,N_19417,N_19351);
nand U21562 (N_21562,N_19843,N_19419);
nand U21563 (N_21563,N_20274,N_19403);
nand U21564 (N_21564,N_18615,N_19167);
nor U21565 (N_21565,N_18407,N_20781);
nand U21566 (N_21566,N_18621,N_19558);
nand U21567 (N_21567,N_19534,N_20448);
xor U21568 (N_21568,N_20771,N_19188);
nor U21569 (N_21569,N_18151,N_20580);
xor U21570 (N_21570,N_19940,N_19770);
or U21571 (N_21571,N_18123,N_18675);
and U21572 (N_21572,N_20108,N_20792);
nand U21573 (N_21573,N_19899,N_18934);
xnor U21574 (N_21574,N_19640,N_19130);
nand U21575 (N_21575,N_18306,N_19427);
or U21576 (N_21576,N_18106,N_19572);
nand U21577 (N_21577,N_20655,N_18879);
and U21578 (N_21578,N_20222,N_18340);
and U21579 (N_21579,N_20548,N_18852);
and U21580 (N_21580,N_20396,N_19647);
nor U21581 (N_21581,N_20922,N_20846);
nand U21582 (N_21582,N_18636,N_20039);
or U21583 (N_21583,N_20283,N_20175);
nand U21584 (N_21584,N_19090,N_18492);
or U21585 (N_21585,N_20643,N_20435);
nor U21586 (N_21586,N_20017,N_18038);
and U21587 (N_21587,N_18353,N_20683);
nand U21588 (N_21588,N_20015,N_18993);
or U21589 (N_21589,N_20164,N_20146);
or U21590 (N_21590,N_19380,N_18045);
xor U21591 (N_21591,N_18517,N_19284);
and U21592 (N_21592,N_18740,N_18829);
xor U21593 (N_21593,N_20246,N_19550);
nor U21594 (N_21594,N_20541,N_19171);
nand U21595 (N_21595,N_20398,N_20069);
xnor U21596 (N_21596,N_20888,N_18866);
nand U21597 (N_21597,N_20357,N_20633);
nor U21598 (N_21598,N_19629,N_18928);
xnor U21599 (N_21599,N_19072,N_19705);
xor U21600 (N_21600,N_19495,N_19720);
or U21601 (N_21601,N_20605,N_18932);
xor U21602 (N_21602,N_19143,N_20026);
or U21603 (N_21603,N_20128,N_19341);
nand U21604 (N_21604,N_18429,N_18733);
nand U21605 (N_21605,N_20364,N_20043);
nor U21606 (N_21606,N_20869,N_18680);
nand U21607 (N_21607,N_19704,N_20808);
or U21608 (N_21608,N_19885,N_18698);
xor U21609 (N_21609,N_19180,N_20883);
nand U21610 (N_21610,N_20608,N_18193);
nand U21611 (N_21611,N_18912,N_19608);
nand U21612 (N_21612,N_20371,N_20050);
nand U21613 (N_21613,N_18982,N_20741);
nor U21614 (N_21614,N_19349,N_20947);
or U21615 (N_21615,N_19202,N_19204);
and U21616 (N_21616,N_18376,N_20368);
nand U21617 (N_21617,N_20711,N_19915);
xor U21618 (N_21618,N_19365,N_20464);
nand U21619 (N_21619,N_20628,N_20221);
or U21620 (N_21620,N_19035,N_18149);
xor U21621 (N_21621,N_19869,N_20932);
nor U21622 (N_21622,N_19759,N_18322);
xor U21623 (N_21623,N_19100,N_20915);
xor U21624 (N_21624,N_19134,N_19172);
nor U21625 (N_21625,N_19164,N_18081);
nand U21626 (N_21626,N_20142,N_19170);
xnor U21627 (N_21627,N_19728,N_18534);
or U21628 (N_21628,N_20460,N_18827);
xor U21629 (N_21629,N_20688,N_20373);
nand U21630 (N_21630,N_18452,N_19458);
xnor U21631 (N_21631,N_18506,N_20466);
nor U21632 (N_21632,N_18040,N_20899);
xnor U21633 (N_21633,N_19841,N_18789);
or U21634 (N_21634,N_19962,N_19026);
nor U21635 (N_21635,N_19842,N_19094);
xnor U21636 (N_21636,N_20169,N_20723);
and U21637 (N_21637,N_18802,N_19108);
nand U21638 (N_21638,N_19449,N_19097);
xor U21639 (N_21639,N_18288,N_20632);
nor U21640 (N_21640,N_20621,N_20122);
or U21641 (N_21641,N_19270,N_20029);
xor U21642 (N_21642,N_20957,N_18160);
nand U21643 (N_21643,N_18037,N_19184);
xnor U21644 (N_21644,N_18196,N_18955);
nand U21645 (N_21645,N_18532,N_20886);
nand U21646 (N_21646,N_18213,N_20207);
nor U21647 (N_21647,N_18291,N_18961);
xor U21648 (N_21648,N_19126,N_20304);
and U21649 (N_21649,N_19262,N_19718);
nand U21650 (N_21650,N_18023,N_19507);
or U21651 (N_21651,N_20417,N_19943);
or U21652 (N_21652,N_19460,N_18838);
nor U21653 (N_21653,N_18100,N_19259);
and U21654 (N_21654,N_19215,N_18569);
xnor U21655 (N_21655,N_20134,N_19566);
nand U21656 (N_21656,N_20537,N_18110);
nor U21657 (N_21657,N_20939,N_19158);
nand U21658 (N_21658,N_19480,N_18052);
nand U21659 (N_21659,N_20350,N_19144);
nand U21660 (N_21660,N_18692,N_18930);
nand U21661 (N_21661,N_18264,N_20646);
and U21662 (N_21662,N_19093,N_19434);
and U21663 (N_21663,N_18773,N_19779);
nor U21664 (N_21664,N_19554,N_19435);
or U21665 (N_21665,N_20901,N_20158);
nand U21666 (N_21666,N_18817,N_19626);
nand U21667 (N_21667,N_18128,N_19782);
or U21668 (N_21668,N_18294,N_20236);
xnor U21669 (N_21669,N_19894,N_19228);
nor U21670 (N_21670,N_19154,N_20325);
or U21671 (N_21671,N_18262,N_18095);
and U21672 (N_21672,N_20730,N_18500);
and U21673 (N_21673,N_19610,N_19444);
xnor U21674 (N_21674,N_20981,N_18808);
and U21675 (N_21675,N_20102,N_18158);
nand U21676 (N_21676,N_18093,N_20669);
or U21677 (N_21677,N_19225,N_20671);
xor U21678 (N_21678,N_20456,N_18016);
xor U21679 (N_21679,N_20731,N_18798);
nor U21680 (N_21680,N_20168,N_18588);
nand U21681 (N_21681,N_20296,N_19192);
or U21682 (N_21682,N_19769,N_18684);
nor U21683 (N_21683,N_19038,N_18903);
nand U21684 (N_21684,N_19918,N_20115);
nand U21685 (N_21685,N_18678,N_18219);
nand U21686 (N_21686,N_19381,N_18528);
and U21687 (N_21687,N_18142,N_18559);
and U21688 (N_21688,N_20072,N_20265);
nor U21689 (N_21689,N_19161,N_20381);
or U21690 (N_21690,N_19731,N_20752);
and U21691 (N_21691,N_20212,N_18512);
nand U21692 (N_21692,N_18823,N_20399);
nand U21693 (N_21693,N_19326,N_19574);
nor U21694 (N_21694,N_20011,N_19808);
or U21695 (N_21695,N_20545,N_19693);
xor U21696 (N_21696,N_20497,N_19584);
and U21697 (N_21697,N_19776,N_18806);
nand U21698 (N_21698,N_19496,N_20639);
nand U21699 (N_21699,N_18977,N_19887);
or U21700 (N_21700,N_19522,N_18470);
and U21701 (N_21701,N_19974,N_20863);
nand U21702 (N_21702,N_18981,N_19504);
xor U21703 (N_21703,N_20121,N_19432);
xnor U21704 (N_21704,N_20470,N_20667);
or U21705 (N_21705,N_20691,N_20389);
xor U21706 (N_21706,N_18384,N_20068);
nand U21707 (N_21707,N_18284,N_20214);
and U21708 (N_21708,N_20547,N_20197);
nor U21709 (N_21709,N_19364,N_19292);
nand U21710 (N_21710,N_18338,N_20751);
nor U21711 (N_21711,N_18260,N_18996);
or U21712 (N_21712,N_20718,N_20407);
and U21713 (N_21713,N_19285,N_19395);
nand U21714 (N_21714,N_20544,N_18246);
xnor U21715 (N_21715,N_19950,N_18576);
nor U21716 (N_21716,N_18602,N_18460);
and U21717 (N_21717,N_20664,N_19638);
and U21718 (N_21718,N_18776,N_18046);
nand U21719 (N_21719,N_20604,N_20716);
nor U21720 (N_21720,N_18372,N_19406);
nand U21721 (N_21721,N_18634,N_20876);
or U21722 (N_21722,N_18226,N_19568);
nor U21723 (N_21723,N_18386,N_18842);
or U21724 (N_21724,N_20380,N_19021);
and U21725 (N_21725,N_20766,N_18305);
nor U21726 (N_21726,N_18794,N_19448);
or U21727 (N_21727,N_20538,N_20622);
nor U21728 (N_21728,N_18455,N_19935);
nor U21729 (N_21729,N_19291,N_19300);
xnor U21730 (N_21730,N_20051,N_20983);
xnor U21731 (N_21731,N_18984,N_19409);
nand U21732 (N_21732,N_18446,N_18997);
and U21733 (N_21733,N_20775,N_19302);
nor U21734 (N_21734,N_20906,N_19973);
nand U21735 (N_21735,N_18639,N_18096);
and U21736 (N_21736,N_18580,N_18231);
or U21737 (N_21737,N_20853,N_19577);
or U21738 (N_21738,N_19657,N_18689);
xnor U21739 (N_21739,N_18234,N_18987);
nor U21740 (N_21740,N_19933,N_18595);
and U21741 (N_21741,N_20889,N_18909);
and U21742 (N_21742,N_18030,N_18472);
xor U21743 (N_21743,N_19084,N_18336);
or U21744 (N_21744,N_20692,N_18969);
nand U21745 (N_21745,N_19178,N_20045);
nor U21746 (N_21746,N_19468,N_20444);
or U21747 (N_21747,N_19985,N_19831);
nor U21748 (N_21748,N_20129,N_19079);
xor U21749 (N_21749,N_18419,N_19726);
nor U21750 (N_21750,N_19878,N_20793);
xnor U21751 (N_21751,N_18940,N_20606);
nor U21752 (N_21752,N_20835,N_18501);
nand U21753 (N_21753,N_20782,N_20806);
nand U21754 (N_21754,N_18599,N_19231);
nor U21755 (N_21755,N_20088,N_19768);
nand U21756 (N_21756,N_19141,N_18267);
and U21757 (N_21757,N_20895,N_18632);
or U21758 (N_21758,N_19137,N_19738);
nor U21759 (N_21759,N_18498,N_18782);
and U21760 (N_21760,N_20126,N_19230);
nor U21761 (N_21761,N_18666,N_20546);
nor U21762 (N_21762,N_19714,N_18399);
nand U21763 (N_21763,N_18318,N_20920);
xor U21764 (N_21764,N_20095,N_19672);
xnor U21765 (N_21765,N_20851,N_18562);
xor U21766 (N_21766,N_20107,N_20096);
or U21767 (N_21767,N_18194,N_20591);
nor U21768 (N_21768,N_20850,N_20263);
xnor U21769 (N_21769,N_18739,N_18959);
nor U21770 (N_21770,N_19474,N_19454);
and U21771 (N_21771,N_20985,N_19165);
or U21772 (N_21772,N_19058,N_20085);
nand U21773 (N_21773,N_18831,N_20481);
and U21774 (N_21774,N_20962,N_19211);
or U21775 (N_21775,N_20218,N_19886);
nand U21776 (N_21776,N_18006,N_18146);
nor U21777 (N_21777,N_20160,N_19996);
and U21778 (N_21778,N_20307,N_20337);
nor U21779 (N_21779,N_20393,N_20558);
nor U21780 (N_21780,N_19311,N_19179);
or U21781 (N_21781,N_19723,N_18077);
or U21782 (N_21782,N_18094,N_20278);
nand U21783 (N_21783,N_20478,N_20504);
or U21784 (N_21784,N_20186,N_20740);
xor U21785 (N_21785,N_20210,N_20650);
and U21786 (N_21786,N_18204,N_18425);
or U21787 (N_21787,N_19960,N_18103);
nor U21788 (N_21788,N_18337,N_19663);
xor U21789 (N_21789,N_19246,N_19786);
xor U21790 (N_21790,N_18439,N_19109);
xor U21791 (N_21791,N_20261,N_19952);
nand U21792 (N_21792,N_19609,N_20975);
nor U21793 (N_21793,N_19561,N_19483);
or U21794 (N_21794,N_19679,N_20656);
xnor U21795 (N_21795,N_19245,N_19819);
and U21796 (N_21796,N_18661,N_18172);
nor U21797 (N_21797,N_19632,N_18024);
or U21798 (N_21798,N_19446,N_19666);
and U21799 (N_21799,N_18292,N_20384);
nand U21800 (N_21800,N_20725,N_20907);
and U21801 (N_21801,N_20659,N_18887);
nand U21802 (N_21802,N_20944,N_18647);
xor U21803 (N_21803,N_20867,N_19242);
nand U21804 (N_21804,N_19103,N_19124);
or U21805 (N_21805,N_18007,N_20352);
xnor U21806 (N_21806,N_19895,N_18111);
nand U21807 (N_21807,N_19162,N_20259);
xnor U21808 (N_21808,N_19557,N_19363);
nor U21809 (N_21809,N_19443,N_19535);
or U21810 (N_21810,N_18937,N_19695);
or U21811 (N_21811,N_18896,N_20370);
nand U21812 (N_21812,N_18527,N_20454);
nand U21813 (N_21813,N_18719,N_18405);
xor U21814 (N_21814,N_20817,N_20154);
nor U21815 (N_21815,N_20491,N_20842);
xor U21816 (N_21816,N_18593,N_20487);
xor U21817 (N_21817,N_19796,N_18413);
nor U21818 (N_21818,N_18343,N_19717);
xor U21819 (N_21819,N_18988,N_20819);
nand U21820 (N_21820,N_19986,N_18947);
nand U21821 (N_21821,N_19919,N_20759);
or U21822 (N_21822,N_18319,N_20721);
nor U21823 (N_21823,N_18169,N_20397);
and U21824 (N_21824,N_19969,N_18558);
xnor U21825 (N_21825,N_18949,N_19512);
or U21826 (N_21826,N_20551,N_20033);
xnor U21827 (N_21827,N_19740,N_19846);
nand U21828 (N_21828,N_20977,N_19438);
nor U21829 (N_21829,N_18116,N_18537);
or U21830 (N_21830,N_19590,N_18751);
nand U21831 (N_21831,N_19022,N_18761);
and U21832 (N_21832,N_19104,N_18594);
nand U21833 (N_21833,N_18513,N_20078);
nand U21834 (N_21834,N_18777,N_18235);
nor U21835 (N_21835,N_19054,N_20676);
xnor U21836 (N_21836,N_20187,N_18447);
and U21837 (N_21837,N_20993,N_20732);
nand U21838 (N_21838,N_18325,N_18082);
nand U21839 (N_21839,N_18396,N_18356);
xnor U21840 (N_21840,N_20048,N_18218);
nand U21841 (N_21841,N_20461,N_19077);
xor U21842 (N_21842,N_19752,N_20585);
nor U21843 (N_21843,N_18202,N_20114);
xor U21844 (N_21844,N_18251,N_18769);
nor U21845 (N_21845,N_18725,N_20410);
xnor U21846 (N_21846,N_20596,N_18550);
xor U21847 (N_21847,N_18851,N_20074);
and U21848 (N_21848,N_19059,N_18468);
or U21849 (N_21849,N_19080,N_19571);
and U21850 (N_21850,N_20912,N_20217);
nand U21851 (N_21851,N_18360,N_19260);
or U21852 (N_21852,N_20362,N_19575);
or U21853 (N_21853,N_20474,N_20594);
xnor U21854 (N_21854,N_20302,N_19673);
or U21855 (N_21855,N_20021,N_19781);
and U21856 (N_21856,N_18956,N_19189);
or U21857 (N_21857,N_18406,N_18718);
or U21858 (N_21858,N_18748,N_18837);
or U21859 (N_21859,N_19420,N_20282);
or U21860 (N_21860,N_20073,N_20194);
nand U21861 (N_21861,N_20503,N_20298);
nor U21862 (N_21862,N_20281,N_19529);
or U21863 (N_21863,N_20193,N_19127);
and U21864 (N_21864,N_19910,N_18418);
nor U21865 (N_21865,N_19394,N_19061);
nand U21866 (N_21866,N_20552,N_20737);
xnor U21867 (N_21867,N_18394,N_20061);
xnor U21868 (N_21868,N_20654,N_19486);
and U21869 (N_21869,N_20961,N_19322);
nand U21870 (N_21870,N_20319,N_20200);
or U21871 (N_21871,N_19343,N_20854);
xor U21872 (N_21872,N_19822,N_20251);
or U21873 (N_21873,N_20301,N_18891);
nor U21874 (N_21874,N_20963,N_19479);
nor U21875 (N_21875,N_20177,N_18991);
nand U21876 (N_21876,N_19589,N_20772);
nor U21877 (N_21877,N_18358,N_18346);
nor U21878 (N_21878,N_20532,N_18669);
nand U21879 (N_21879,N_18134,N_20712);
nor U21880 (N_21880,N_20490,N_18775);
nor U21881 (N_21881,N_19198,N_20184);
nor U21882 (N_21882,N_19152,N_20413);
xor U21883 (N_21883,N_18926,N_18067);
xor U21884 (N_21884,N_19553,N_18474);
xnor U21885 (N_21885,N_20080,N_19746);
nor U21886 (N_21886,N_20505,N_18843);
nand U21887 (N_21887,N_18951,N_18001);
xor U21888 (N_21888,N_19999,N_19613);
and U21889 (N_21889,N_20902,N_19903);
and U21890 (N_21890,N_20697,N_20070);
and U21891 (N_21891,N_19713,N_20288);
nor U21892 (N_21892,N_18945,N_18805);
nand U21893 (N_21893,N_18783,N_19536);
nand U21894 (N_21894,N_18479,N_19856);
xnor U21895 (N_21895,N_18013,N_20434);
nand U21896 (N_21896,N_18228,N_19062);
xnor U21897 (N_21897,N_18720,N_18953);
nor U21898 (N_21898,N_18099,N_20272);
or U21899 (N_21899,N_19146,N_19065);
xnor U21900 (N_21900,N_19096,N_19067);
or U21901 (N_21901,N_19762,N_18868);
and U21902 (N_21902,N_20969,N_18760);
nor U21903 (N_21903,N_18542,N_19857);
nor U21904 (N_21904,N_20227,N_20412);
nand U21905 (N_21905,N_20153,N_18008);
xnor U21906 (N_21906,N_20736,N_19683);
nand U21907 (N_21907,N_19175,N_18690);
or U21908 (N_21908,N_18252,N_20855);
nor U21909 (N_21909,N_18464,N_18000);
nor U21910 (N_21910,N_19199,N_18138);
nor U21911 (N_21911,N_19298,N_19234);
or U21912 (N_21912,N_20662,N_18834);
xnor U21913 (N_21913,N_20573,N_20372);
nor U21914 (N_21914,N_19281,N_20202);
and U21915 (N_21915,N_19370,N_18073);
nor U21916 (N_21916,N_19001,N_19815);
xnor U21917 (N_21917,N_19874,N_18515);
nor U21918 (N_21918,N_19033,N_19359);
nor U21919 (N_21919,N_18314,N_18638);
nor U21920 (N_21920,N_18531,N_18217);
or U21921 (N_21921,N_20063,N_20885);
nand U21922 (N_21922,N_20386,N_19177);
or U21923 (N_21923,N_20420,N_20645);
xor U21924 (N_21924,N_19282,N_20404);
nor U21925 (N_21925,N_20948,N_20705);
xor U21926 (N_21926,N_20810,N_19772);
xor U21927 (N_21927,N_20999,N_18387);
xor U21928 (N_21928,N_18191,N_19527);
nor U21929 (N_21929,N_19818,N_19451);
nand U21930 (N_21930,N_20925,N_20756);
or U21931 (N_21931,N_19832,N_20666);
nand U21932 (N_21932,N_18002,N_18302);
nand U21933 (N_21933,N_18102,N_19521);
nand U21934 (N_21934,N_19977,N_18581);
and U21935 (N_21935,N_18324,N_20226);
nand U21936 (N_21936,N_18950,N_18120);
nor U21937 (N_21937,N_20220,N_20877);
and U21938 (N_21938,N_20875,N_19493);
nand U21939 (N_21939,N_18627,N_19991);
or U21940 (N_21940,N_20715,N_20893);
and U21941 (N_21941,N_18828,N_18494);
or U21942 (N_21942,N_20570,N_19475);
or U21943 (N_21943,N_18884,N_20308);
nand U21944 (N_21944,N_20776,N_19965);
xnor U21945 (N_21945,N_19140,N_20881);
nand U21946 (N_21946,N_20964,N_19400);
or U21947 (N_21947,N_20784,N_20244);
xnor U21948 (N_21948,N_19978,N_19307);
or U21949 (N_21949,N_19051,N_20832);
and U21950 (N_21950,N_18489,N_19719);
xor U21951 (N_21951,N_19913,N_19684);
xnor U21952 (N_21952,N_19605,N_19795);
or U21953 (N_21953,N_20223,N_18605);
nand U21954 (N_21954,N_18286,N_18836);
nand U21955 (N_21955,N_20597,N_18064);
or U21956 (N_21956,N_18758,N_18211);
or U21957 (N_21957,N_19481,N_18657);
xnor U21958 (N_21958,N_19639,N_18109);
nor U21959 (N_21959,N_19086,N_20452);
nor U21960 (N_21960,N_18607,N_18687);
or U21961 (N_21961,N_18029,N_19687);
nor U21962 (N_21962,N_18994,N_19386);
and U21963 (N_21963,N_20421,N_20789);
nand U21964 (N_21964,N_19541,N_19265);
or U21965 (N_21965,N_20672,N_19357);
or U21966 (N_21966,N_20339,N_20742);
xnor U21967 (N_21967,N_18148,N_18335);
nor U21968 (N_21968,N_20822,N_19337);
nand U21969 (N_21969,N_19083,N_18821);
xor U21970 (N_21970,N_18899,N_20911);
xnor U21971 (N_21971,N_18368,N_19426);
or U21972 (N_21972,N_18674,N_20127);
nor U21973 (N_21973,N_19459,N_20600);
nor U21974 (N_21974,N_20367,N_18066);
or U21975 (N_21975,N_20693,N_19612);
nor U21976 (N_21976,N_18119,N_18762);
nand U21977 (N_21977,N_19102,N_18874);
nand U21978 (N_21978,N_19513,N_20215);
and U21979 (N_21979,N_18401,N_20847);
nand U21980 (N_21980,N_19593,N_18563);
and U21981 (N_21981,N_20774,N_18973);
or U21982 (N_21982,N_18787,N_19827);
and U21983 (N_21983,N_20140,N_18300);
xnor U21984 (N_21984,N_20954,N_18793);
nor U21985 (N_21985,N_18265,N_20219);
and U21986 (N_21986,N_19788,N_18876);
and U21987 (N_21987,N_20856,N_19848);
nor U21988 (N_21988,N_18239,N_18967);
nand U21989 (N_21989,N_18931,N_20117);
or U21990 (N_21990,N_18809,N_18074);
or U21991 (N_21991,N_19360,N_20438);
nor U21992 (N_21992,N_20475,N_20609);
nor U21993 (N_21993,N_20812,N_19176);
xnor U21994 (N_21994,N_20658,N_20829);
and U21995 (N_21995,N_18826,N_20374);
or U21996 (N_21996,N_18443,N_18520);
and U21997 (N_21997,N_19564,N_19076);
or U21998 (N_21998,N_19377,N_18673);
nor U21999 (N_21999,N_19393,N_19018);
nand U22000 (N_22000,N_20322,N_19042);
nor U22001 (N_22001,N_18033,N_20514);
or U22002 (N_22002,N_18248,N_18192);
nor U22003 (N_22003,N_20579,N_20453);
nor U22004 (N_22004,N_20427,N_18964);
xnor U22005 (N_22005,N_20882,N_18092);
and U22006 (N_22006,N_19329,N_18709);
nor U22007 (N_22007,N_20746,N_20509);
or U22008 (N_22008,N_18972,N_19267);
nor U22009 (N_22009,N_18367,N_19671);
xor U22010 (N_22010,N_20483,N_19217);
and U22011 (N_22011,N_18960,N_20770);
and U22012 (N_22012,N_19653,N_19428);
nor U22013 (N_22013,N_19971,N_19498);
or U22014 (N_22014,N_18359,N_18171);
or U22015 (N_22015,N_19688,N_20923);
xor U22016 (N_22016,N_20285,N_19946);
and U22017 (N_22017,N_20934,N_19194);
or U22018 (N_22018,N_20284,N_18509);
xor U22019 (N_22019,N_18279,N_19024);
nor U22020 (N_22020,N_18466,N_18901);
xor U22021 (N_22021,N_20196,N_19668);
nor U22022 (N_22022,N_20572,N_19658);
or U22023 (N_22023,N_19235,N_20273);
nand U22024 (N_22024,N_19710,N_18814);
and U22025 (N_22025,N_18224,N_19087);
nand U22026 (N_22026,N_18643,N_20825);
xor U22027 (N_22027,N_20034,N_20356);
xnor U22028 (N_22028,N_18502,N_18212);
and U22029 (N_22029,N_19754,N_19324);
or U22030 (N_22030,N_18608,N_18247);
or U22031 (N_22031,N_19711,N_18174);
and U22032 (N_22032,N_20726,N_19239);
or U22033 (N_22033,N_19689,N_19588);
xnor U22034 (N_22034,N_20358,N_18285);
or U22035 (N_22035,N_18548,N_19257);
nand U22036 (N_22036,N_18862,N_19548);
or U22037 (N_22037,N_19757,N_19611);
or U22038 (N_22038,N_20583,N_19722);
or U22039 (N_22039,N_18652,N_18485);
or U22040 (N_22040,N_19685,N_19404);
nand U22041 (N_22041,N_20249,N_19981);
nand U22042 (N_22042,N_20685,N_19680);
nand U22043 (N_22043,N_18624,N_19835);
nor U22044 (N_22044,N_19181,N_18181);
xor U22045 (N_22045,N_20536,N_20254);
nor U22046 (N_22046,N_20046,N_18768);
nor U22047 (N_22047,N_18451,N_19870);
and U22048 (N_22048,N_20361,N_20592);
and U22049 (N_22049,N_18567,N_19983);
xor U22050 (N_22050,N_19447,N_18946);
and U22051 (N_22051,N_20727,N_18107);
xnor U22052 (N_22052,N_20653,N_19002);
and U22053 (N_22053,N_20578,N_18321);
nor U22054 (N_22054,N_19802,N_18907);
or U22055 (N_22055,N_19369,N_19958);
xor U22056 (N_22056,N_20484,N_19068);
and U22057 (N_22057,N_20728,N_18237);
or U22058 (N_22058,N_19641,N_20860);
nor U22059 (N_22059,N_19889,N_18009);
and U22060 (N_22060,N_20204,N_20113);
and U22061 (N_22061,N_19044,N_18487);
nor U22062 (N_22062,N_19218,N_20250);
or U22063 (N_22063,N_19826,N_19755);
nor U22064 (N_22064,N_20816,N_20376);
or U22065 (N_22065,N_18478,N_19209);
nor U22066 (N_22066,N_19347,N_19489);
and U22067 (N_22067,N_18122,N_19064);
and U22068 (N_22068,N_20722,N_19539);
or U22069 (N_22069,N_18242,N_18012);
xnor U22070 (N_22070,N_20586,N_19206);
nor U22071 (N_22071,N_18431,N_20897);
nor U22072 (N_22072,N_20400,N_18952);
and U22073 (N_22073,N_19549,N_18241);
or U22074 (N_22074,N_20450,N_19148);
nand U22075 (N_22075,N_19092,N_20513);
nand U22076 (N_22076,N_18839,N_20682);
nor U22077 (N_22077,N_20192,N_19600);
nor U22078 (N_22078,N_19352,N_20482);
xnor U22079 (N_22079,N_19492,N_20000);
or U22080 (N_22080,N_20630,N_18070);
and U22081 (N_22081,N_18985,N_19073);
nor U22082 (N_22082,N_20206,N_18480);
and U22083 (N_22083,N_18373,N_18710);
nand U22084 (N_22084,N_18524,N_20267);
nand U22085 (N_22085,N_18711,N_19744);
nor U22086 (N_22086,N_18792,N_20042);
nand U22087 (N_22087,N_20190,N_19316);
nand U22088 (N_22088,N_19615,N_20511);
xnor U22089 (N_22089,N_19373,N_18746);
nand U22090 (N_22090,N_18872,N_20191);
or U22091 (N_22091,N_20130,N_20429);
xnor U22092 (N_22092,N_19956,N_18902);
and U22093 (N_22093,N_19650,N_20744);
xor U22094 (N_22094,N_18278,N_18296);
nand U22095 (N_22095,N_19602,N_19220);
and U22096 (N_22096,N_18966,N_18163);
xnor U22097 (N_22097,N_18395,N_20987);
nand U22098 (N_22098,N_20027,N_18154);
xnor U22099 (N_22099,N_19266,N_18175);
or U22100 (N_22100,N_20098,N_20065);
nand U22101 (N_22101,N_18779,N_19367);
xnor U22102 (N_22102,N_18227,N_19560);
nor U22103 (N_22103,N_19767,N_19543);
or U22104 (N_22104,N_20980,N_19039);
or U22105 (N_22105,N_20949,N_20312);
and U22106 (N_22106,N_20188,N_20517);
nor U22107 (N_22107,N_19346,N_18249);
and U22108 (N_22108,N_18589,N_20136);
or U22109 (N_22109,N_18035,N_20529);
or U22110 (N_22110,N_19532,N_18786);
nand U22111 (N_22111,N_18883,N_20295);
or U22112 (N_22112,N_19037,N_19734);
nand U22113 (N_22113,N_20878,N_19132);
xor U22114 (N_22114,N_20791,N_19453);
and U22115 (N_22115,N_20125,N_20459);
or U22116 (N_22116,N_19052,N_18543);
and U22117 (N_22117,N_18545,N_19789);
nor U22118 (N_22118,N_20661,N_18922);
nor U22119 (N_22119,N_19310,N_20101);
nand U22120 (N_22120,N_18818,N_20343);
or U22121 (N_22121,N_20965,N_20103);
xnor U22122 (N_22122,N_20100,N_18141);
xnor U22123 (N_22123,N_20455,N_18131);
nor U22124 (N_22124,N_19654,N_18841);
nor U22125 (N_22125,N_20910,N_19145);
and U22126 (N_22126,N_19811,N_18700);
or U22127 (N_22127,N_19221,N_20216);
nor U22128 (N_22128,N_19273,N_20778);
xnor U22129 (N_22129,N_19040,N_20139);
xor U22130 (N_22130,N_20446,N_18737);
or U22131 (N_22131,N_18433,N_20521);
xnor U22132 (N_22132,N_20428,N_18295);
and U22133 (N_22133,N_19676,N_18525);
nor U22134 (N_22134,N_19066,N_19004);
and U22135 (N_22135,N_20238,N_20651);
or U22136 (N_22136,N_19801,N_18375);
nor U22137 (N_22137,N_19354,N_19005);
xor U22138 (N_22138,N_20994,N_19990);
and U22139 (N_22139,N_18601,N_20022);
xnor U22140 (N_22140,N_19742,N_19494);
and U22141 (N_22141,N_18233,N_19847);
and U22142 (N_22142,N_20815,N_19855);
xnor U22143 (N_22143,N_19166,N_19758);
and U22144 (N_22144,N_18349,N_18205);
and U22145 (N_22145,N_18299,N_20549);
and U22146 (N_22146,N_18735,N_20392);
or U22147 (N_22147,N_19556,N_18223);
or U22148 (N_22148,N_19635,N_19817);
nand U22149 (N_22149,N_19440,N_20313);
xnor U22150 (N_22150,N_18167,N_19542);
and U22151 (N_22151,N_20803,N_18721);
and U22152 (N_22152,N_18626,N_20124);
nor U22153 (N_22153,N_20224,N_20635);
xnor U22154 (N_22154,N_18297,N_18200);
or U22155 (N_22155,N_19069,N_19252);
or U22156 (N_22156,N_19442,N_19290);
and U22157 (N_22157,N_19436,N_19953);
and U22158 (N_22158,N_19837,N_20508);
nor U22159 (N_22159,N_19321,N_18667);
nand U22160 (N_22160,N_20933,N_19309);
or U22161 (N_22161,N_20232,N_19401);
or U22162 (N_22162,N_19019,N_20891);
and U22163 (N_22163,N_19579,N_19877);
and U22164 (N_22164,N_19614,N_18199);
xnor U22165 (N_22165,N_18707,N_20761);
nor U22166 (N_22166,N_18206,N_20512);
or U22167 (N_22167,N_18220,N_18612);
and U22168 (N_22168,N_18269,N_18178);
xor U22169 (N_22169,N_18941,N_19911);
and U22170 (N_22170,N_18764,N_19830);
nand U22171 (N_22171,N_18423,N_18597);
nor U22172 (N_22172,N_18822,N_19954);
or U22173 (N_22173,N_18271,N_20610);
xnor U22174 (N_22174,N_20624,N_20363);
or U22175 (N_22175,N_18812,N_20657);
or U22176 (N_22176,N_20336,N_20440);
nand U22177 (N_22177,N_19727,N_19623);
nand U22178 (N_22178,N_20056,N_18778);
xor U22179 (N_22179,N_20974,N_18381);
xnor U22180 (N_22180,N_18263,N_19160);
xnor U22181 (N_22181,N_20060,N_20037);
nor U22182 (N_22182,N_20087,N_19120);
nand U22183 (N_22183,N_18021,N_18726);
nor U22184 (N_22184,N_20001,N_20038);
xor U22185 (N_22185,N_20431,N_20275);
and U22186 (N_22186,N_18989,N_18904);
xnor U22187 (N_22187,N_18027,N_20110);
xor U22188 (N_22188,N_20820,N_20673);
xor U22189 (N_22189,N_18958,N_19375);
or U22190 (N_22190,N_18905,N_19461);
nand U22191 (N_22191,N_19917,N_18290);
nor U22192 (N_22192,N_19620,N_18150);
xnor U22193 (N_22193,N_20092,N_19733);
and U22194 (N_22194,N_19248,N_18459);
and U22195 (N_22195,N_20351,N_19328);
or U22196 (N_22196,N_19502,N_19630);
nor U22197 (N_22197,N_18694,N_18441);
and U22198 (N_22198,N_20623,N_19256);
nor U22199 (N_22199,N_19222,N_19208);
nor U22200 (N_22200,N_19247,N_19224);
or U22201 (N_22201,N_19402,N_18328);
nand U22202 (N_22202,N_20841,N_18071);
and U22203 (N_22203,N_20488,N_20229);
nand U22204 (N_22204,N_19537,N_20859);
xor U22205 (N_22205,N_20857,N_20342);
xnor U22206 (N_22206,N_18510,N_18414);
xor U22207 (N_22207,N_18623,N_18784);
nor U22208 (N_22208,N_18871,N_20607);
and U22209 (N_22209,N_18450,N_18068);
nor U22210 (N_22210,N_19000,N_18867);
xor U22211 (N_22211,N_20248,N_18449);
or U22212 (N_22212,N_20178,N_20523);
nand U22213 (N_22213,N_19197,N_20104);
nand U22214 (N_22214,N_18716,N_18209);
or U22215 (N_22215,N_20366,N_18190);
and U22216 (N_22216,N_18853,N_18579);
and U22217 (N_22217,N_20058,N_20449);
or U22218 (N_22218,N_19793,N_19187);
xor U22219 (N_22219,N_19562,N_20075);
nand U22220 (N_22220,N_19477,N_20747);
and U22221 (N_22221,N_20928,N_18770);
or U22222 (N_22222,N_18963,N_19464);
and U22223 (N_22223,N_18079,N_18744);
xor U22224 (N_22224,N_18885,N_18813);
xnor U22225 (N_22225,N_19128,N_20297);
and U22226 (N_22226,N_20148,N_18403);
nor U22227 (N_22227,N_18428,N_18412);
xnor U22228 (N_22228,N_20968,N_18062);
nor U22229 (N_22229,N_19702,N_18722);
or U22230 (N_22230,N_19691,N_18143);
xnor U22231 (N_22231,N_20496,N_19295);
or U22232 (N_22232,N_19631,N_19088);
or U22233 (N_22233,N_20890,N_18345);
nand U22234 (N_22234,N_18189,N_20441);
xnor U22235 (N_22235,N_19345,N_20613);
nor U22236 (N_22236,N_19439,N_18895);
or U22237 (N_22237,N_19387,N_19118);
or U22238 (N_22238,N_18566,N_18893);
and U22239 (N_22239,N_20047,N_18378);
nor U22240 (N_22240,N_20111,N_18084);
nor U22241 (N_22241,N_19951,N_19159);
and U22242 (N_22242,N_18650,N_20317);
xnor U22243 (N_22243,N_19664,N_20706);
xor U22244 (N_22244,N_19053,N_18495);
xor U22245 (N_22245,N_18232,N_19195);
xnor U22246 (N_22246,N_20516,N_18075);
nand U22247 (N_22247,N_20094,N_20059);
nand U22248 (N_22248,N_20268,N_20131);
or U22249 (N_22249,N_19138,N_19976);
and U22250 (N_22250,N_19382,N_20405);
xnor U22251 (N_22251,N_19339,N_20264);
nand U22252 (N_22252,N_20834,N_20515);
and U22253 (N_22253,N_18943,N_18208);
xnor U22254 (N_22254,N_19437,N_19379);
nand U22255 (N_22255,N_19948,N_18882);
and U22256 (N_22256,N_18811,N_19573);
nand U22257 (N_22257,N_19476,N_20277);
xor U22258 (N_22258,N_18363,N_19814);
and U22259 (N_22259,N_18309,N_18801);
nand U22260 (N_22260,N_19926,N_20365);
xnor U22261 (N_22261,N_20465,N_20595);
and U22262 (N_22262,N_20908,N_18918);
nand U22263 (N_22263,N_19881,N_19078);
or U22264 (N_22264,N_18028,N_19810);
or U22265 (N_22265,N_20331,N_18072);
and U22266 (N_22266,N_18047,N_18900);
xor U22267 (N_22267,N_19936,N_20520);
or U22268 (N_22268,N_20865,N_18276);
or U22269 (N_22269,N_20005,N_18857);
xor U22270 (N_22270,N_19747,N_19122);
xnor U22271 (N_22271,N_18214,N_19669);
nor U22272 (N_22272,N_20385,N_20831);
and U22273 (N_22273,N_18476,N_18645);
and U22274 (N_22274,N_19385,N_18310);
nand U22275 (N_22275,N_18546,N_20403);
nand U22276 (N_22276,N_18986,N_18655);
nor U22277 (N_22277,N_20790,N_19660);
nor U22278 (N_22278,N_19633,N_20062);
nand U22279 (N_22279,N_20010,N_18488);
or U22280 (N_22280,N_18243,N_18800);
nor U22281 (N_22281,N_19665,N_18182);
nand U22282 (N_22282,N_20266,N_19925);
nor U22283 (N_22283,N_18465,N_19212);
and U22284 (N_22284,N_19760,N_18177);
xnor U22285 (N_22285,N_18560,N_20506);
nand U22286 (N_22286,N_18699,N_18166);
and U22287 (N_22287,N_19739,N_19232);
xor U22288 (N_22288,N_19455,N_18574);
nor U22289 (N_22289,N_18121,N_19457);
nand U22290 (N_22290,N_19834,N_20524);
or U22291 (N_22291,N_20642,N_19113);
nor U22292 (N_22292,N_20260,N_19875);
or U22293 (N_22293,N_20919,N_18069);
nand U22294 (N_22294,N_20799,N_20694);
nand U22295 (N_22295,N_19293,N_19261);
and U22296 (N_22296,N_19043,N_20917);
nor U22297 (N_22297,N_20714,N_18139);
and U22298 (N_22298,N_18729,N_18734);
or U22299 (N_22299,N_19567,N_20309);
or U22300 (N_22300,N_19743,N_19216);
or U22301 (N_22301,N_19025,N_18327);
or U22302 (N_22302,N_20310,N_20501);
nor U22303 (N_22303,N_18736,N_18408);
nand U22304 (N_22304,N_18129,N_20930);
xnor U22305 (N_22305,N_18591,N_18417);
xor U22306 (N_22306,N_20745,N_18914);
nand U22307 (N_22307,N_20601,N_19528);
xor U22308 (N_22308,N_19836,N_19748);
and U22309 (N_22309,N_18854,N_20280);
and U22310 (N_22310,N_19462,N_20067);
nand U22311 (N_22311,N_19183,N_20151);
nand U22312 (N_22312,N_19555,N_19771);
nor U22313 (N_22313,N_20225,N_19271);
or U22314 (N_22314,N_19975,N_18766);
xor U22315 (N_22315,N_20577,N_19233);
nand U22316 (N_22316,N_20498,N_20502);
or U22317 (N_22317,N_20849,N_18539);
nor U22318 (N_22318,N_18535,N_18658);
nor U22319 (N_22319,N_20530,N_19643);
and U22320 (N_22320,N_20959,N_20174);
and U22321 (N_22321,N_18377,N_20344);
and U22322 (N_22322,N_18660,N_20821);
xnor U22323 (N_22323,N_18810,N_20240);
nor U22324 (N_22324,N_19344,N_18889);
and U22325 (N_22325,N_18308,N_19289);
nor U22326 (N_22326,N_20439,N_19106);
and U22327 (N_22327,N_18164,N_20006);
or U22328 (N_22328,N_20408,N_18496);
xnor U22329 (N_22329,N_18424,N_20698);
nor U22330 (N_22330,N_19362,N_19433);
xor U22331 (N_22331,N_19014,N_18481);
and U22332 (N_22332,N_19932,N_19773);
nand U22333 (N_22333,N_19471,N_20471);
nor U22334 (N_22334,N_18686,N_18482);
or U22335 (N_22335,N_18771,N_19893);
nor U22336 (N_22336,N_18229,N_20769);
nor U22337 (N_22337,N_19678,N_19955);
or U22338 (N_22338,N_20862,N_20436);
or U22339 (N_22339,N_18938,N_18897);
nand U22340 (N_22340,N_20602,N_20415);
nor U22341 (N_22341,N_20913,N_19196);
and U22342 (N_22342,N_18254,N_19497);
nor U22343 (N_22343,N_19942,N_20049);
nand U22344 (N_22344,N_19944,N_19961);
and U22345 (N_22345,N_18705,N_18104);
xnor U22346 (N_22346,N_20674,N_19585);
nand U22347 (N_22347,N_19296,N_19010);
nand U22348 (N_22348,N_20425,N_18919);
and U22349 (N_22349,N_19249,N_18054);
nor U22350 (N_22350,N_19651,N_18393);
nor U22351 (N_22351,N_20355,N_18458);
and U22352 (N_22352,N_20848,N_19563);
xor U22353 (N_22353,N_18313,N_20554);
or U22354 (N_22354,N_20828,N_19902);
nand U22355 (N_22355,N_20024,N_19514);
nor U22356 (N_22356,N_19303,N_18547);
xnor U22357 (N_22357,N_18357,N_18526);
or U22358 (N_22358,N_18238,N_19997);
or U22359 (N_22359,N_20258,N_18625);
nand U22360 (N_22360,N_20914,N_18780);
nand U22361 (N_22361,N_20996,N_18592);
xor U22362 (N_22362,N_19283,N_18788);
nor U22363 (N_22363,N_18438,N_18980);
nand U22364 (N_22364,N_20709,N_20838);
or U22365 (N_22365,N_20442,N_20800);
and U22366 (N_22366,N_18004,N_20701);
nand U22367 (N_22367,N_19253,N_19783);
and U22368 (N_22368,N_19694,N_18553);
xor U22369 (N_22369,N_18448,N_18754);
xnor U22370 (N_22370,N_19591,N_19675);
and U22371 (N_22371,N_19644,N_19491);
or U22372 (N_22372,N_19804,N_19136);
nand U22373 (N_22373,N_19055,N_19408);
nor U22374 (N_22374,N_19547,N_18640);
nor U22375 (N_22375,N_20935,N_20009);
xor U22376 (N_22376,N_20823,N_19523);
xor U22377 (N_22377,N_19264,N_18173);
and U22378 (N_22378,N_18048,N_18388);
nor U22379 (N_22379,N_20754,N_20681);
nor U22380 (N_22380,N_20013,N_20531);
or U22381 (N_22381,N_18772,N_18990);
nor U22382 (N_22382,N_20534,N_20237);
and U22383 (N_22383,N_18463,N_20720);
and U22384 (N_22384,N_20896,N_20183);
or U22385 (N_22385,N_18486,N_19994);
nand U22386 (N_22386,N_19957,N_18888);
or U22387 (N_22387,N_20590,N_18742);
xnor U22388 (N_22388,N_18998,N_19603);
xnor U22389 (N_22389,N_19648,N_20587);
nand U22390 (N_22390,N_18522,N_19500);
or U22391 (N_22391,N_20926,N_20231);
nand U22392 (N_22392,N_19777,N_20451);
or U22393 (N_22393,N_18400,N_19263);
xnor U22394 (N_22394,N_19173,N_19117);
and U22395 (N_22395,N_20324,N_18402);
xor U22396 (N_22396,N_19190,N_19601);
or U22397 (N_22397,N_19587,N_20409);
xnor U22398 (N_22398,N_19229,N_19515);
and U22399 (N_22399,N_20443,N_18763);
xor U22400 (N_22400,N_19089,N_18221);
nor U22401 (N_22401,N_20276,N_18679);
xor U22402 (N_22402,N_19931,N_20710);
or U22403 (N_22403,N_19763,N_19012);
and U22404 (N_22404,N_18293,N_19849);
nor U22405 (N_22405,N_19214,N_19545);
and U22406 (N_22406,N_20976,N_18790);
nand U22407 (N_22407,N_20105,N_19095);
nor U22408 (N_22408,N_20494,N_20241);
nor U22409 (N_22409,N_20335,N_20208);
and U22410 (N_22410,N_20649,N_18274);
nor U22411 (N_22411,N_19112,N_19622);
nand U22412 (N_22412,N_19803,N_20519);
or U22413 (N_22413,N_18572,N_19325);
nand U22414 (N_22414,N_20507,N_20025);
nand U22415 (N_22415,N_20713,N_20695);
and U22416 (N_22416,N_18549,N_20702);
nor U22417 (N_22417,N_18379,N_20967);
and U22418 (N_22418,N_20571,N_20469);
or U22419 (N_22419,N_20287,N_20689);
nand U22420 (N_22420,N_18124,N_19972);
and U22421 (N_22421,N_19907,N_20631);
nand U22422 (N_22422,N_18765,N_18738);
or U22423 (N_22423,N_20861,N_18440);
nand U22424 (N_22424,N_18339,N_18708);
nor U22425 (N_22425,N_18552,N_18323);
nand U22426 (N_22426,N_19928,N_20457);
and U22427 (N_22427,N_20257,N_18333);
xor U22428 (N_22428,N_18796,N_18039);
nor U22429 (N_22429,N_20458,N_20748);
or U22430 (N_22430,N_19331,N_19860);
nor U22431 (N_22431,N_20071,N_20750);
xor U22432 (N_22432,N_18939,N_18923);
and U22433 (N_22433,N_19565,N_20879);
and U22434 (N_22434,N_20582,N_19508);
nor U22435 (N_22435,N_18628,N_18435);
xnor U22436 (N_22436,N_19157,N_18642);
nor U22437 (N_22437,N_18374,N_18043);
nor U22438 (N_22438,N_19908,N_20181);
or U22439 (N_22439,N_18957,N_19323);
nor U22440 (N_22440,N_20665,N_19938);
and U22441 (N_22441,N_20023,N_19750);
or U22442 (N_22442,N_20638,N_18855);
or U22443 (N_22443,N_20614,N_18518);
nand U22444 (N_22444,N_18712,N_20979);
and U22445 (N_22445,N_20700,N_20433);
xnor U22446 (N_22446,N_19661,N_19923);
or U22447 (N_22447,N_18677,N_20802);
and U22448 (N_22448,N_19824,N_18087);
xnor U22449 (N_22449,N_19226,N_19101);
and U22450 (N_22450,N_18240,N_20090);
nand U22451 (N_22451,N_19790,N_18971);
xnor U22452 (N_22452,N_18717,N_20956);
and U22453 (N_22453,N_18538,N_18785);
nor U22454 (N_22454,N_19998,N_18055);
or U22455 (N_22455,N_18184,N_20211);
or U22456 (N_22456,N_19397,N_20463);
and U22457 (N_22457,N_19546,N_19511);
nand U22458 (N_22458,N_20567,N_18536);
or U22459 (N_22459,N_19701,N_20884);
or U22460 (N_22460,N_20271,N_18210);
and U22461 (N_22461,N_20640,N_19645);
nand U22462 (N_22462,N_18410,N_19749);
nand U22463 (N_22463,N_18664,N_18473);
or U22464 (N_22464,N_20887,N_20566);
xnor U22465 (N_22465,N_19174,N_20270);
nand U22466 (N_22466,N_18114,N_20118);
nand U22467 (N_22467,N_18330,N_18144);
and U22468 (N_22468,N_19637,N_20201);
and U22469 (N_22469,N_19135,N_20411);
nor U22470 (N_22470,N_19473,N_18332);
or U22471 (N_22471,N_19011,N_20008);
or U22472 (N_22472,N_20982,N_18730);
nor U22473 (N_22473,N_18618,N_19866);
xnor U22474 (N_22474,N_19378,N_20332);
xor U22475 (N_22475,N_20866,N_19070);
and U22476 (N_22476,N_18316,N_18256);
nor U22477 (N_22477,N_20252,N_18825);
xor U22478 (N_22478,N_20414,N_19056);
nand U22479 (N_22479,N_20028,N_20675);
nand U22480 (N_22480,N_20588,N_18797);
nand U22481 (N_22481,N_19524,N_20157);
xnor U22482 (N_22482,N_18130,N_18065);
xor U22483 (N_22483,N_19703,N_18490);
or U22484 (N_22484,N_19304,N_19872);
and U22485 (N_22485,N_20724,N_19366);
nor U22486 (N_22486,N_20172,N_18179);
nor U22487 (N_22487,N_18920,N_19578);
xnor U22488 (N_22488,N_20423,N_19142);
nor U22489 (N_22489,N_19732,N_19350);
and U22490 (N_22490,N_18056,N_19445);
xnor U22491 (N_22491,N_20864,N_18767);
and U22492 (N_22492,N_18083,N_19333);
xnor U22493 (N_22493,N_20300,N_19967);
and U22494 (N_22494,N_19930,N_20824);
nand U22495 (N_22495,N_19517,N_19131);
nor U22496 (N_22496,N_20230,N_20032);
and U22497 (N_22497,N_20991,N_18948);
xnor U22498 (N_22498,N_20437,N_18886);
nand U22499 (N_22499,N_18598,N_18105);
nand U22500 (N_22500,N_19061,N_20023);
or U22501 (N_22501,N_19230,N_19833);
nand U22502 (N_22502,N_18877,N_18662);
and U22503 (N_22503,N_18548,N_18950);
and U22504 (N_22504,N_18997,N_19433);
nand U22505 (N_22505,N_20569,N_20084);
and U22506 (N_22506,N_19872,N_19886);
and U22507 (N_22507,N_19156,N_18295);
xor U22508 (N_22508,N_20995,N_19918);
nor U22509 (N_22509,N_18427,N_18989);
xor U22510 (N_22510,N_19477,N_20105);
nand U22511 (N_22511,N_20119,N_19792);
or U22512 (N_22512,N_18452,N_20952);
nand U22513 (N_22513,N_20617,N_19671);
or U22514 (N_22514,N_19042,N_19126);
or U22515 (N_22515,N_19147,N_19972);
or U22516 (N_22516,N_20853,N_19788);
xor U22517 (N_22517,N_18136,N_20558);
or U22518 (N_22518,N_19469,N_20496);
and U22519 (N_22519,N_20518,N_18188);
and U22520 (N_22520,N_20887,N_18524);
nor U22521 (N_22521,N_19888,N_18082);
xnor U22522 (N_22522,N_19683,N_18036);
or U22523 (N_22523,N_19583,N_19817);
and U22524 (N_22524,N_19228,N_19556);
and U22525 (N_22525,N_20544,N_20200);
nand U22526 (N_22526,N_18406,N_18328);
or U22527 (N_22527,N_19582,N_20129);
and U22528 (N_22528,N_19319,N_18194);
or U22529 (N_22529,N_20365,N_18935);
xnor U22530 (N_22530,N_20915,N_18321);
and U22531 (N_22531,N_18926,N_20138);
or U22532 (N_22532,N_18749,N_19591);
nor U22533 (N_22533,N_20871,N_19582);
nor U22534 (N_22534,N_20763,N_20066);
or U22535 (N_22535,N_18040,N_18338);
and U22536 (N_22536,N_19632,N_20271);
nor U22537 (N_22537,N_18423,N_20937);
and U22538 (N_22538,N_19492,N_19455);
or U22539 (N_22539,N_18992,N_20097);
and U22540 (N_22540,N_18684,N_18430);
nor U22541 (N_22541,N_19867,N_19712);
xnor U22542 (N_22542,N_19040,N_19663);
and U22543 (N_22543,N_18992,N_18977);
nand U22544 (N_22544,N_18425,N_20235);
xnor U22545 (N_22545,N_20953,N_18700);
nand U22546 (N_22546,N_18298,N_20416);
xor U22547 (N_22547,N_20374,N_19206);
nand U22548 (N_22548,N_18035,N_19648);
nand U22549 (N_22549,N_19049,N_19701);
nor U22550 (N_22550,N_19651,N_19290);
nor U22551 (N_22551,N_19912,N_19952);
nand U22552 (N_22552,N_20126,N_19237);
nand U22553 (N_22553,N_19324,N_18687);
xor U22554 (N_22554,N_18011,N_19094);
nor U22555 (N_22555,N_18414,N_20634);
nand U22556 (N_22556,N_20558,N_20561);
nand U22557 (N_22557,N_18593,N_18675);
or U22558 (N_22558,N_18991,N_20618);
xnor U22559 (N_22559,N_20675,N_18021);
xor U22560 (N_22560,N_20402,N_18061);
nand U22561 (N_22561,N_20020,N_18958);
nor U22562 (N_22562,N_19912,N_18727);
xor U22563 (N_22563,N_20064,N_19876);
nor U22564 (N_22564,N_19439,N_20689);
and U22565 (N_22565,N_18052,N_18838);
or U22566 (N_22566,N_19640,N_19010);
nand U22567 (N_22567,N_19123,N_20512);
nor U22568 (N_22568,N_20121,N_19744);
nand U22569 (N_22569,N_18431,N_20183);
and U22570 (N_22570,N_20066,N_18275);
and U22571 (N_22571,N_19112,N_20862);
nand U22572 (N_22572,N_18675,N_18253);
nor U22573 (N_22573,N_20089,N_20565);
or U22574 (N_22574,N_20570,N_20079);
and U22575 (N_22575,N_18920,N_18344);
xnor U22576 (N_22576,N_19674,N_19783);
nor U22577 (N_22577,N_20825,N_18603);
nand U22578 (N_22578,N_19934,N_20629);
or U22579 (N_22579,N_19264,N_20674);
or U22580 (N_22580,N_19761,N_20424);
or U22581 (N_22581,N_19170,N_20350);
and U22582 (N_22582,N_19575,N_19735);
and U22583 (N_22583,N_18644,N_19112);
nand U22584 (N_22584,N_18407,N_19843);
and U22585 (N_22585,N_18085,N_19191);
nand U22586 (N_22586,N_19512,N_20970);
and U22587 (N_22587,N_19633,N_20473);
nor U22588 (N_22588,N_19210,N_19856);
and U22589 (N_22589,N_20208,N_20822);
xor U22590 (N_22590,N_20017,N_18367);
xnor U22591 (N_22591,N_20566,N_20796);
or U22592 (N_22592,N_19209,N_20353);
nand U22593 (N_22593,N_19425,N_18405);
nor U22594 (N_22594,N_18976,N_18558);
and U22595 (N_22595,N_20467,N_19968);
nand U22596 (N_22596,N_20277,N_18110);
nor U22597 (N_22597,N_19716,N_19858);
nand U22598 (N_22598,N_18071,N_20461);
nor U22599 (N_22599,N_18296,N_19871);
nor U22600 (N_22600,N_20440,N_18000);
and U22601 (N_22601,N_20293,N_18485);
nor U22602 (N_22602,N_19791,N_18117);
and U22603 (N_22603,N_18761,N_18990);
xor U22604 (N_22604,N_19992,N_19835);
and U22605 (N_22605,N_19440,N_18002);
and U22606 (N_22606,N_19339,N_19514);
or U22607 (N_22607,N_19386,N_20956);
xnor U22608 (N_22608,N_20078,N_19890);
xnor U22609 (N_22609,N_20877,N_20532);
or U22610 (N_22610,N_18845,N_18794);
and U22611 (N_22611,N_20421,N_18214);
nor U22612 (N_22612,N_20811,N_20829);
or U22613 (N_22613,N_20508,N_20869);
and U22614 (N_22614,N_20471,N_18358);
nor U22615 (N_22615,N_19524,N_20905);
or U22616 (N_22616,N_18077,N_19783);
nand U22617 (N_22617,N_18580,N_20458);
nor U22618 (N_22618,N_19665,N_19214);
nand U22619 (N_22619,N_19710,N_20049);
nand U22620 (N_22620,N_20079,N_19327);
xor U22621 (N_22621,N_20225,N_19789);
nor U22622 (N_22622,N_20463,N_18196);
nand U22623 (N_22623,N_20683,N_20425);
nor U22624 (N_22624,N_18555,N_20292);
and U22625 (N_22625,N_18445,N_18573);
xor U22626 (N_22626,N_19006,N_18391);
or U22627 (N_22627,N_20525,N_18334);
xnor U22628 (N_22628,N_18975,N_20903);
or U22629 (N_22629,N_20829,N_20941);
nor U22630 (N_22630,N_19157,N_20476);
and U22631 (N_22631,N_18897,N_18491);
and U22632 (N_22632,N_18484,N_20465);
and U22633 (N_22633,N_20123,N_18730);
nand U22634 (N_22634,N_18893,N_19290);
xor U22635 (N_22635,N_20985,N_18938);
xor U22636 (N_22636,N_18193,N_19683);
nor U22637 (N_22637,N_19278,N_19296);
xor U22638 (N_22638,N_19797,N_18153);
nand U22639 (N_22639,N_20745,N_19975);
nor U22640 (N_22640,N_20530,N_20230);
or U22641 (N_22641,N_18798,N_19862);
and U22642 (N_22642,N_19107,N_20325);
xnor U22643 (N_22643,N_19085,N_20016);
nand U22644 (N_22644,N_20550,N_19541);
and U22645 (N_22645,N_20912,N_19635);
xnor U22646 (N_22646,N_20380,N_20609);
and U22647 (N_22647,N_20400,N_19568);
xnor U22648 (N_22648,N_20424,N_18878);
and U22649 (N_22649,N_19546,N_20132);
xnor U22650 (N_22650,N_18598,N_18080);
and U22651 (N_22651,N_18113,N_18333);
and U22652 (N_22652,N_19478,N_18095);
nand U22653 (N_22653,N_19211,N_20913);
xor U22654 (N_22654,N_20659,N_19802);
and U22655 (N_22655,N_18029,N_18147);
xor U22656 (N_22656,N_18984,N_18334);
xnor U22657 (N_22657,N_18902,N_19135);
or U22658 (N_22658,N_18779,N_20168);
xnor U22659 (N_22659,N_19677,N_20226);
xor U22660 (N_22660,N_18372,N_20733);
xnor U22661 (N_22661,N_18148,N_18289);
nand U22662 (N_22662,N_19393,N_19202);
nor U22663 (N_22663,N_20463,N_20423);
or U22664 (N_22664,N_19088,N_19875);
nand U22665 (N_22665,N_18339,N_19557);
xor U22666 (N_22666,N_19605,N_20905);
nand U22667 (N_22667,N_19869,N_19257);
and U22668 (N_22668,N_20342,N_18559);
xor U22669 (N_22669,N_18336,N_20030);
and U22670 (N_22670,N_18597,N_19206);
xor U22671 (N_22671,N_20854,N_19789);
or U22672 (N_22672,N_20320,N_18865);
nor U22673 (N_22673,N_20992,N_20941);
xnor U22674 (N_22674,N_20619,N_18955);
nor U22675 (N_22675,N_19628,N_20145);
or U22676 (N_22676,N_20133,N_20362);
xnor U22677 (N_22677,N_19896,N_19655);
or U22678 (N_22678,N_19471,N_18007);
and U22679 (N_22679,N_18445,N_20961);
xor U22680 (N_22680,N_18404,N_19957);
nor U22681 (N_22681,N_18150,N_18849);
xor U22682 (N_22682,N_18066,N_19212);
nor U22683 (N_22683,N_18373,N_19640);
nor U22684 (N_22684,N_19175,N_19660);
or U22685 (N_22685,N_18874,N_18064);
or U22686 (N_22686,N_20439,N_19320);
xor U22687 (N_22687,N_18149,N_18304);
nand U22688 (N_22688,N_19088,N_18197);
xnor U22689 (N_22689,N_19394,N_20350);
nor U22690 (N_22690,N_19389,N_20443);
and U22691 (N_22691,N_19990,N_19906);
xnor U22692 (N_22692,N_20772,N_19131);
xnor U22693 (N_22693,N_19110,N_20201);
nor U22694 (N_22694,N_18169,N_20959);
nor U22695 (N_22695,N_19290,N_20155);
xor U22696 (N_22696,N_19434,N_18318);
or U22697 (N_22697,N_18637,N_18067);
and U22698 (N_22698,N_19563,N_19575);
and U22699 (N_22699,N_20741,N_19440);
and U22700 (N_22700,N_19301,N_19928);
nor U22701 (N_22701,N_19368,N_20454);
xnor U22702 (N_22702,N_18496,N_18267);
or U22703 (N_22703,N_19269,N_18722);
nor U22704 (N_22704,N_20836,N_18242);
nand U22705 (N_22705,N_20054,N_18043);
and U22706 (N_22706,N_19041,N_18951);
xor U22707 (N_22707,N_20143,N_20490);
or U22708 (N_22708,N_18318,N_18925);
nor U22709 (N_22709,N_19593,N_18140);
or U22710 (N_22710,N_19912,N_18342);
and U22711 (N_22711,N_18582,N_20621);
nand U22712 (N_22712,N_18907,N_18852);
xnor U22713 (N_22713,N_18922,N_20347);
nand U22714 (N_22714,N_20941,N_19505);
and U22715 (N_22715,N_18452,N_19944);
nand U22716 (N_22716,N_20053,N_20394);
and U22717 (N_22717,N_20101,N_19940);
xor U22718 (N_22718,N_20884,N_20750);
nand U22719 (N_22719,N_18796,N_18497);
nand U22720 (N_22720,N_19606,N_19730);
and U22721 (N_22721,N_19305,N_19410);
xor U22722 (N_22722,N_18356,N_18181);
nand U22723 (N_22723,N_18318,N_20242);
or U22724 (N_22724,N_18288,N_19068);
nor U22725 (N_22725,N_19844,N_19188);
or U22726 (N_22726,N_18281,N_18864);
nor U22727 (N_22727,N_18546,N_18796);
xor U22728 (N_22728,N_18716,N_19332);
xnor U22729 (N_22729,N_19560,N_20024);
or U22730 (N_22730,N_18424,N_18931);
or U22731 (N_22731,N_19155,N_18203);
nor U22732 (N_22732,N_20233,N_19575);
nand U22733 (N_22733,N_20329,N_18179);
and U22734 (N_22734,N_20009,N_19479);
and U22735 (N_22735,N_19456,N_20224);
and U22736 (N_22736,N_18390,N_19038);
nor U22737 (N_22737,N_18627,N_18543);
or U22738 (N_22738,N_19642,N_20233);
nand U22739 (N_22739,N_18649,N_19207);
nor U22740 (N_22740,N_18568,N_18138);
xor U22741 (N_22741,N_18880,N_18856);
or U22742 (N_22742,N_18007,N_19909);
xor U22743 (N_22743,N_20227,N_18442);
and U22744 (N_22744,N_20009,N_20615);
nor U22745 (N_22745,N_20733,N_19872);
or U22746 (N_22746,N_18009,N_19518);
and U22747 (N_22747,N_18497,N_19268);
nand U22748 (N_22748,N_18458,N_18426);
nor U22749 (N_22749,N_18371,N_19555);
nand U22750 (N_22750,N_18693,N_19956);
or U22751 (N_22751,N_20475,N_20593);
nor U22752 (N_22752,N_20098,N_18138);
or U22753 (N_22753,N_20323,N_18510);
nor U22754 (N_22754,N_20556,N_18164);
nor U22755 (N_22755,N_19269,N_18303);
and U22756 (N_22756,N_18463,N_20962);
xnor U22757 (N_22757,N_19617,N_19352);
or U22758 (N_22758,N_20438,N_18289);
xnor U22759 (N_22759,N_20006,N_20576);
nor U22760 (N_22760,N_20749,N_19572);
or U22761 (N_22761,N_20696,N_19673);
and U22762 (N_22762,N_18471,N_20317);
xor U22763 (N_22763,N_20207,N_19465);
xnor U22764 (N_22764,N_20350,N_19630);
xor U22765 (N_22765,N_19647,N_18262);
or U22766 (N_22766,N_19264,N_19912);
or U22767 (N_22767,N_19731,N_20731);
xnor U22768 (N_22768,N_18403,N_20517);
xor U22769 (N_22769,N_20054,N_18928);
xor U22770 (N_22770,N_18782,N_20052);
xor U22771 (N_22771,N_19008,N_19767);
or U22772 (N_22772,N_20471,N_20455);
nand U22773 (N_22773,N_19843,N_20567);
nand U22774 (N_22774,N_19185,N_18755);
or U22775 (N_22775,N_20166,N_19226);
or U22776 (N_22776,N_18737,N_18859);
nand U22777 (N_22777,N_20857,N_18707);
nor U22778 (N_22778,N_19547,N_19079);
nand U22779 (N_22779,N_20600,N_20360);
and U22780 (N_22780,N_20277,N_19789);
nor U22781 (N_22781,N_19972,N_18261);
nor U22782 (N_22782,N_18845,N_18926);
xor U22783 (N_22783,N_19299,N_20586);
nor U22784 (N_22784,N_20605,N_18389);
or U22785 (N_22785,N_18126,N_18042);
and U22786 (N_22786,N_19388,N_18449);
nor U22787 (N_22787,N_19194,N_19453);
nor U22788 (N_22788,N_19020,N_19473);
nor U22789 (N_22789,N_20307,N_20908);
xnor U22790 (N_22790,N_19483,N_20371);
xnor U22791 (N_22791,N_20525,N_19922);
and U22792 (N_22792,N_20734,N_19510);
nand U22793 (N_22793,N_18679,N_19420);
nand U22794 (N_22794,N_18079,N_20965);
or U22795 (N_22795,N_20288,N_18309);
nand U22796 (N_22796,N_18434,N_19808);
nand U22797 (N_22797,N_19353,N_18327);
or U22798 (N_22798,N_20229,N_20567);
xnor U22799 (N_22799,N_19298,N_18696);
nand U22800 (N_22800,N_19875,N_18386);
or U22801 (N_22801,N_18932,N_20047);
xnor U22802 (N_22802,N_18596,N_20295);
or U22803 (N_22803,N_20937,N_19427);
xor U22804 (N_22804,N_18674,N_18582);
or U22805 (N_22805,N_19226,N_18527);
xnor U22806 (N_22806,N_19279,N_18736);
nor U22807 (N_22807,N_20745,N_18197);
nor U22808 (N_22808,N_19041,N_20871);
nor U22809 (N_22809,N_20839,N_20771);
and U22810 (N_22810,N_18701,N_18471);
and U22811 (N_22811,N_19042,N_19567);
nor U22812 (N_22812,N_20558,N_18534);
nor U22813 (N_22813,N_19384,N_20738);
nand U22814 (N_22814,N_18383,N_19111);
and U22815 (N_22815,N_20034,N_20666);
and U22816 (N_22816,N_19143,N_19246);
or U22817 (N_22817,N_20004,N_20503);
nand U22818 (N_22818,N_19915,N_18672);
nor U22819 (N_22819,N_18732,N_20350);
or U22820 (N_22820,N_20833,N_18195);
and U22821 (N_22821,N_18096,N_19983);
xor U22822 (N_22822,N_19326,N_19358);
and U22823 (N_22823,N_19570,N_18153);
xor U22824 (N_22824,N_20447,N_18143);
or U22825 (N_22825,N_19385,N_19344);
nor U22826 (N_22826,N_20475,N_19847);
and U22827 (N_22827,N_19761,N_18131);
and U22828 (N_22828,N_19580,N_20861);
and U22829 (N_22829,N_18200,N_19274);
or U22830 (N_22830,N_20084,N_19574);
and U22831 (N_22831,N_20726,N_18260);
and U22832 (N_22832,N_20664,N_20812);
xor U22833 (N_22833,N_20327,N_18751);
xnor U22834 (N_22834,N_18308,N_20386);
nor U22835 (N_22835,N_20676,N_20782);
xor U22836 (N_22836,N_20735,N_20626);
or U22837 (N_22837,N_19070,N_18722);
xnor U22838 (N_22838,N_19122,N_19666);
or U22839 (N_22839,N_18036,N_19627);
nand U22840 (N_22840,N_18646,N_19787);
or U22841 (N_22841,N_20674,N_20828);
nand U22842 (N_22842,N_20422,N_18702);
nor U22843 (N_22843,N_20345,N_18815);
xnor U22844 (N_22844,N_18360,N_18177);
or U22845 (N_22845,N_18763,N_18447);
xnor U22846 (N_22846,N_19613,N_19079);
nand U22847 (N_22847,N_19510,N_20916);
xnor U22848 (N_22848,N_18360,N_18318);
xnor U22849 (N_22849,N_20318,N_20483);
nand U22850 (N_22850,N_20039,N_18664);
nor U22851 (N_22851,N_20705,N_19995);
and U22852 (N_22852,N_19201,N_19124);
xor U22853 (N_22853,N_18899,N_18360);
nand U22854 (N_22854,N_18816,N_18967);
or U22855 (N_22855,N_18093,N_18314);
nand U22856 (N_22856,N_19992,N_20244);
xnor U22857 (N_22857,N_19594,N_18791);
nand U22858 (N_22858,N_18303,N_18412);
or U22859 (N_22859,N_18185,N_20430);
xor U22860 (N_22860,N_20100,N_19740);
nor U22861 (N_22861,N_19909,N_19897);
and U22862 (N_22862,N_19141,N_20223);
nor U22863 (N_22863,N_20212,N_20103);
and U22864 (N_22864,N_18375,N_18530);
or U22865 (N_22865,N_18858,N_19246);
xnor U22866 (N_22866,N_20655,N_18224);
nand U22867 (N_22867,N_18448,N_20017);
or U22868 (N_22868,N_18052,N_18140);
and U22869 (N_22869,N_18834,N_20902);
nand U22870 (N_22870,N_20708,N_20688);
or U22871 (N_22871,N_19225,N_19338);
nor U22872 (N_22872,N_18548,N_19496);
nand U22873 (N_22873,N_18378,N_19763);
xnor U22874 (N_22874,N_20507,N_20408);
and U22875 (N_22875,N_18196,N_19512);
and U22876 (N_22876,N_20222,N_18542);
and U22877 (N_22877,N_19062,N_19536);
nor U22878 (N_22878,N_18752,N_19448);
or U22879 (N_22879,N_18016,N_19042);
xnor U22880 (N_22880,N_19396,N_18539);
and U22881 (N_22881,N_19766,N_20784);
nor U22882 (N_22882,N_19219,N_20791);
nand U22883 (N_22883,N_20482,N_19798);
xor U22884 (N_22884,N_20074,N_19681);
nor U22885 (N_22885,N_20328,N_20877);
nand U22886 (N_22886,N_20184,N_18205);
nand U22887 (N_22887,N_18951,N_18997);
and U22888 (N_22888,N_18975,N_20397);
xnor U22889 (N_22889,N_19698,N_19748);
nand U22890 (N_22890,N_19056,N_18533);
and U22891 (N_22891,N_20162,N_18896);
nand U22892 (N_22892,N_19235,N_19427);
nor U22893 (N_22893,N_18531,N_18869);
and U22894 (N_22894,N_18599,N_20298);
and U22895 (N_22895,N_18161,N_18032);
or U22896 (N_22896,N_18012,N_19133);
or U22897 (N_22897,N_19995,N_18902);
nor U22898 (N_22898,N_20692,N_20895);
nand U22899 (N_22899,N_18070,N_20639);
xnor U22900 (N_22900,N_18961,N_18795);
nor U22901 (N_22901,N_19711,N_18587);
nand U22902 (N_22902,N_19062,N_18172);
and U22903 (N_22903,N_20790,N_18952);
xnor U22904 (N_22904,N_19449,N_19345);
xnor U22905 (N_22905,N_18938,N_20779);
xnor U22906 (N_22906,N_20983,N_18958);
nor U22907 (N_22907,N_19516,N_18067);
xor U22908 (N_22908,N_18844,N_19517);
nand U22909 (N_22909,N_18210,N_18300);
xnor U22910 (N_22910,N_20330,N_20544);
or U22911 (N_22911,N_18853,N_20864);
nor U22912 (N_22912,N_19673,N_18886);
nand U22913 (N_22913,N_19483,N_20608);
and U22914 (N_22914,N_20114,N_20015);
nand U22915 (N_22915,N_19120,N_18824);
or U22916 (N_22916,N_20093,N_18695);
or U22917 (N_22917,N_20709,N_20680);
nand U22918 (N_22918,N_19482,N_19051);
or U22919 (N_22919,N_19943,N_18487);
and U22920 (N_22920,N_18758,N_18249);
and U22921 (N_22921,N_18510,N_20022);
nand U22922 (N_22922,N_18050,N_19389);
nor U22923 (N_22923,N_20844,N_20211);
nand U22924 (N_22924,N_20541,N_18803);
xor U22925 (N_22925,N_19185,N_18608);
nand U22926 (N_22926,N_18551,N_18170);
nand U22927 (N_22927,N_18576,N_18043);
nor U22928 (N_22928,N_20992,N_20490);
nor U22929 (N_22929,N_18918,N_18281);
and U22930 (N_22930,N_18740,N_18410);
or U22931 (N_22931,N_19934,N_18748);
xnor U22932 (N_22932,N_18447,N_20158);
or U22933 (N_22933,N_19007,N_19867);
or U22934 (N_22934,N_19264,N_19674);
nand U22935 (N_22935,N_20999,N_18091);
nand U22936 (N_22936,N_19573,N_20985);
nor U22937 (N_22937,N_20828,N_18541);
and U22938 (N_22938,N_19253,N_19432);
xor U22939 (N_22939,N_20814,N_18437);
and U22940 (N_22940,N_18451,N_20136);
or U22941 (N_22941,N_20590,N_18166);
and U22942 (N_22942,N_18693,N_19919);
or U22943 (N_22943,N_20233,N_18320);
or U22944 (N_22944,N_18174,N_19705);
nand U22945 (N_22945,N_18520,N_18797);
and U22946 (N_22946,N_19560,N_20824);
and U22947 (N_22947,N_20143,N_20012);
nor U22948 (N_22948,N_20337,N_19637);
nor U22949 (N_22949,N_20435,N_18211);
nand U22950 (N_22950,N_19348,N_18557);
or U22951 (N_22951,N_20275,N_19121);
nand U22952 (N_22952,N_19743,N_19778);
nor U22953 (N_22953,N_18871,N_20955);
nand U22954 (N_22954,N_20214,N_19968);
or U22955 (N_22955,N_18263,N_20202);
or U22956 (N_22956,N_20314,N_19351);
or U22957 (N_22957,N_19910,N_20097);
and U22958 (N_22958,N_19366,N_20811);
xnor U22959 (N_22959,N_20332,N_20295);
and U22960 (N_22960,N_20695,N_18493);
nor U22961 (N_22961,N_20033,N_20640);
nand U22962 (N_22962,N_20517,N_20358);
xnor U22963 (N_22963,N_18185,N_20475);
and U22964 (N_22964,N_20989,N_20997);
or U22965 (N_22965,N_20975,N_19584);
nand U22966 (N_22966,N_19411,N_18024);
nor U22967 (N_22967,N_18391,N_18875);
nor U22968 (N_22968,N_20246,N_18241);
and U22969 (N_22969,N_18208,N_18247);
xor U22970 (N_22970,N_20386,N_19105);
nand U22971 (N_22971,N_19220,N_18073);
nor U22972 (N_22972,N_19713,N_20872);
nor U22973 (N_22973,N_19426,N_19024);
nand U22974 (N_22974,N_18384,N_18079);
nand U22975 (N_22975,N_18762,N_20136);
xnor U22976 (N_22976,N_19534,N_18197);
and U22977 (N_22977,N_20758,N_19869);
xnor U22978 (N_22978,N_18000,N_19791);
nor U22979 (N_22979,N_20940,N_19023);
or U22980 (N_22980,N_20475,N_20134);
and U22981 (N_22981,N_20954,N_19241);
nand U22982 (N_22982,N_19014,N_19930);
or U22983 (N_22983,N_19931,N_20519);
nor U22984 (N_22984,N_19262,N_18366);
xor U22985 (N_22985,N_18772,N_18830);
or U22986 (N_22986,N_18467,N_20406);
nor U22987 (N_22987,N_20031,N_19403);
nor U22988 (N_22988,N_20800,N_18933);
xor U22989 (N_22989,N_20636,N_20838);
xnor U22990 (N_22990,N_18388,N_19060);
and U22991 (N_22991,N_19493,N_20472);
nand U22992 (N_22992,N_19708,N_19066);
or U22993 (N_22993,N_20553,N_18093);
nor U22994 (N_22994,N_20467,N_20848);
or U22995 (N_22995,N_18374,N_18939);
xnor U22996 (N_22996,N_19820,N_18788);
or U22997 (N_22997,N_18714,N_19385);
and U22998 (N_22998,N_19406,N_18869);
and U22999 (N_22999,N_18763,N_20960);
or U23000 (N_23000,N_18414,N_18151);
or U23001 (N_23001,N_19678,N_19861);
xnor U23002 (N_23002,N_18018,N_20064);
xor U23003 (N_23003,N_18078,N_20066);
nor U23004 (N_23004,N_19275,N_18490);
nand U23005 (N_23005,N_19406,N_19204);
nor U23006 (N_23006,N_20778,N_20706);
nor U23007 (N_23007,N_19282,N_18589);
or U23008 (N_23008,N_19893,N_18041);
and U23009 (N_23009,N_20730,N_19382);
nand U23010 (N_23010,N_20463,N_18601);
nor U23011 (N_23011,N_20730,N_19604);
xor U23012 (N_23012,N_19288,N_19289);
and U23013 (N_23013,N_18803,N_18498);
and U23014 (N_23014,N_19726,N_19363);
xor U23015 (N_23015,N_19007,N_19271);
xor U23016 (N_23016,N_20550,N_18814);
and U23017 (N_23017,N_19552,N_20048);
xnor U23018 (N_23018,N_20401,N_19130);
nand U23019 (N_23019,N_19331,N_20496);
or U23020 (N_23020,N_18967,N_19410);
xnor U23021 (N_23021,N_19652,N_18536);
nor U23022 (N_23022,N_20145,N_19033);
nor U23023 (N_23023,N_18548,N_18152);
xor U23024 (N_23024,N_18112,N_20938);
xor U23025 (N_23025,N_19088,N_20660);
and U23026 (N_23026,N_18356,N_18459);
or U23027 (N_23027,N_19194,N_20164);
and U23028 (N_23028,N_19124,N_19827);
nor U23029 (N_23029,N_20038,N_19835);
nor U23030 (N_23030,N_18941,N_18002);
nand U23031 (N_23031,N_18181,N_18345);
or U23032 (N_23032,N_19771,N_20330);
xor U23033 (N_23033,N_19772,N_20051);
and U23034 (N_23034,N_18531,N_19803);
or U23035 (N_23035,N_19062,N_20481);
nand U23036 (N_23036,N_18421,N_19289);
and U23037 (N_23037,N_18428,N_20583);
or U23038 (N_23038,N_19066,N_19080);
and U23039 (N_23039,N_18896,N_19567);
nand U23040 (N_23040,N_20518,N_19948);
nor U23041 (N_23041,N_20611,N_20995);
xor U23042 (N_23042,N_20422,N_20633);
or U23043 (N_23043,N_20963,N_20723);
xnor U23044 (N_23044,N_18586,N_20247);
or U23045 (N_23045,N_20947,N_18996);
xor U23046 (N_23046,N_20039,N_20704);
or U23047 (N_23047,N_18362,N_20501);
xnor U23048 (N_23048,N_20962,N_20123);
and U23049 (N_23049,N_20147,N_18079);
nand U23050 (N_23050,N_18388,N_20115);
nor U23051 (N_23051,N_20062,N_19987);
or U23052 (N_23052,N_20895,N_18232);
xnor U23053 (N_23053,N_18203,N_20577);
and U23054 (N_23054,N_18040,N_19338);
nand U23055 (N_23055,N_18809,N_20350);
nand U23056 (N_23056,N_18158,N_18898);
nor U23057 (N_23057,N_20757,N_20765);
nor U23058 (N_23058,N_19990,N_19178);
or U23059 (N_23059,N_20847,N_18521);
xor U23060 (N_23060,N_19713,N_19379);
nor U23061 (N_23061,N_18759,N_19241);
nor U23062 (N_23062,N_18251,N_19810);
nor U23063 (N_23063,N_20957,N_18324);
xnor U23064 (N_23064,N_18250,N_18081);
xnor U23065 (N_23065,N_20964,N_20032);
or U23066 (N_23066,N_18186,N_18669);
xor U23067 (N_23067,N_19805,N_18449);
and U23068 (N_23068,N_18479,N_20326);
or U23069 (N_23069,N_19865,N_19973);
or U23070 (N_23070,N_18085,N_18550);
or U23071 (N_23071,N_20757,N_19194);
xnor U23072 (N_23072,N_19388,N_20275);
nor U23073 (N_23073,N_20803,N_20939);
or U23074 (N_23074,N_18270,N_19166);
nand U23075 (N_23075,N_20184,N_20975);
nor U23076 (N_23076,N_20007,N_19834);
nor U23077 (N_23077,N_20877,N_18738);
xnor U23078 (N_23078,N_20339,N_18091);
nor U23079 (N_23079,N_18108,N_19578);
and U23080 (N_23080,N_18996,N_19046);
nor U23081 (N_23081,N_19875,N_20055);
nor U23082 (N_23082,N_19220,N_20586);
xnor U23083 (N_23083,N_18497,N_20551);
and U23084 (N_23084,N_20292,N_18982);
and U23085 (N_23085,N_20568,N_20718);
xor U23086 (N_23086,N_19291,N_18944);
nand U23087 (N_23087,N_20274,N_20037);
nor U23088 (N_23088,N_20656,N_18363);
or U23089 (N_23089,N_18745,N_18513);
nand U23090 (N_23090,N_18164,N_20715);
nor U23091 (N_23091,N_18588,N_18868);
nand U23092 (N_23092,N_18263,N_19316);
xor U23093 (N_23093,N_20749,N_19071);
xnor U23094 (N_23094,N_18967,N_19896);
xor U23095 (N_23095,N_18629,N_18938);
and U23096 (N_23096,N_19280,N_20020);
and U23097 (N_23097,N_18669,N_20587);
xor U23098 (N_23098,N_18092,N_19284);
xor U23099 (N_23099,N_19443,N_18525);
and U23100 (N_23100,N_18728,N_18910);
xnor U23101 (N_23101,N_20024,N_20148);
nand U23102 (N_23102,N_19238,N_20327);
or U23103 (N_23103,N_20019,N_20093);
and U23104 (N_23104,N_19976,N_19020);
and U23105 (N_23105,N_18942,N_18331);
xor U23106 (N_23106,N_20045,N_20849);
xnor U23107 (N_23107,N_19221,N_19551);
xor U23108 (N_23108,N_18164,N_19800);
xor U23109 (N_23109,N_19374,N_19635);
nor U23110 (N_23110,N_19602,N_19625);
nand U23111 (N_23111,N_18601,N_18289);
nand U23112 (N_23112,N_19068,N_20303);
nand U23113 (N_23113,N_20748,N_19440);
xor U23114 (N_23114,N_19456,N_20187);
nand U23115 (N_23115,N_18646,N_20402);
and U23116 (N_23116,N_19152,N_19478);
nand U23117 (N_23117,N_19289,N_19404);
nand U23118 (N_23118,N_18032,N_19043);
and U23119 (N_23119,N_19964,N_19645);
nand U23120 (N_23120,N_20711,N_19005);
nor U23121 (N_23121,N_19341,N_18196);
and U23122 (N_23122,N_19047,N_19490);
nand U23123 (N_23123,N_20594,N_18730);
xor U23124 (N_23124,N_20648,N_19581);
xnor U23125 (N_23125,N_18714,N_18631);
xnor U23126 (N_23126,N_18451,N_18322);
xor U23127 (N_23127,N_18291,N_18084);
and U23128 (N_23128,N_18186,N_18762);
nand U23129 (N_23129,N_19387,N_20029);
and U23130 (N_23130,N_19529,N_20119);
xor U23131 (N_23131,N_19921,N_19766);
nor U23132 (N_23132,N_20921,N_20868);
nor U23133 (N_23133,N_19624,N_18499);
nand U23134 (N_23134,N_18621,N_18932);
and U23135 (N_23135,N_18384,N_20158);
and U23136 (N_23136,N_19107,N_19131);
or U23137 (N_23137,N_19353,N_20075);
nand U23138 (N_23138,N_20841,N_18279);
nor U23139 (N_23139,N_20034,N_18638);
xnor U23140 (N_23140,N_20633,N_18604);
nor U23141 (N_23141,N_19956,N_19050);
nor U23142 (N_23142,N_18914,N_19852);
and U23143 (N_23143,N_18832,N_18822);
nand U23144 (N_23144,N_18974,N_20317);
xor U23145 (N_23145,N_19745,N_20044);
or U23146 (N_23146,N_19072,N_19562);
xor U23147 (N_23147,N_20279,N_18851);
xnor U23148 (N_23148,N_19269,N_18128);
xor U23149 (N_23149,N_20616,N_20864);
nor U23150 (N_23150,N_18375,N_19562);
and U23151 (N_23151,N_19813,N_20514);
xor U23152 (N_23152,N_19890,N_20524);
or U23153 (N_23153,N_18215,N_20567);
and U23154 (N_23154,N_19964,N_19068);
nor U23155 (N_23155,N_20664,N_18644);
nor U23156 (N_23156,N_18267,N_20633);
xnor U23157 (N_23157,N_19545,N_19967);
nor U23158 (N_23158,N_19862,N_19602);
xnor U23159 (N_23159,N_18115,N_18133);
or U23160 (N_23160,N_20955,N_19180);
and U23161 (N_23161,N_18509,N_19090);
xor U23162 (N_23162,N_19069,N_19173);
xnor U23163 (N_23163,N_18430,N_19823);
and U23164 (N_23164,N_19631,N_20983);
and U23165 (N_23165,N_18479,N_20607);
nor U23166 (N_23166,N_20402,N_20051);
xor U23167 (N_23167,N_18633,N_18183);
nand U23168 (N_23168,N_18137,N_19740);
or U23169 (N_23169,N_19817,N_19533);
or U23170 (N_23170,N_18668,N_19266);
and U23171 (N_23171,N_20310,N_18973);
and U23172 (N_23172,N_18074,N_18524);
nand U23173 (N_23173,N_19349,N_19277);
and U23174 (N_23174,N_20320,N_19612);
or U23175 (N_23175,N_20675,N_18006);
nand U23176 (N_23176,N_19525,N_20791);
or U23177 (N_23177,N_18358,N_20623);
nor U23178 (N_23178,N_18536,N_19208);
nor U23179 (N_23179,N_18415,N_20855);
nand U23180 (N_23180,N_20004,N_19145);
nor U23181 (N_23181,N_20019,N_19994);
nor U23182 (N_23182,N_18838,N_19734);
xnor U23183 (N_23183,N_18223,N_20718);
xor U23184 (N_23184,N_18863,N_20862);
xnor U23185 (N_23185,N_19205,N_20968);
xor U23186 (N_23186,N_18140,N_20675);
nand U23187 (N_23187,N_20190,N_20830);
nor U23188 (N_23188,N_19087,N_19043);
or U23189 (N_23189,N_19873,N_20120);
and U23190 (N_23190,N_20581,N_20092);
nor U23191 (N_23191,N_18664,N_20949);
xnor U23192 (N_23192,N_18426,N_20217);
or U23193 (N_23193,N_20233,N_20323);
and U23194 (N_23194,N_20419,N_18211);
nand U23195 (N_23195,N_18748,N_18784);
and U23196 (N_23196,N_20562,N_18610);
nor U23197 (N_23197,N_19869,N_18924);
nor U23198 (N_23198,N_20146,N_20606);
nor U23199 (N_23199,N_19187,N_20147);
nor U23200 (N_23200,N_18696,N_18374);
and U23201 (N_23201,N_18097,N_19258);
or U23202 (N_23202,N_20970,N_19020);
xor U23203 (N_23203,N_19570,N_20412);
nor U23204 (N_23204,N_18203,N_20998);
nand U23205 (N_23205,N_18062,N_18337);
and U23206 (N_23206,N_19401,N_19001);
nor U23207 (N_23207,N_19857,N_19651);
nand U23208 (N_23208,N_20679,N_19261);
or U23209 (N_23209,N_19251,N_18761);
and U23210 (N_23210,N_19458,N_19221);
nand U23211 (N_23211,N_20808,N_19263);
and U23212 (N_23212,N_18312,N_20765);
nand U23213 (N_23213,N_18340,N_20090);
or U23214 (N_23214,N_20200,N_19458);
nand U23215 (N_23215,N_18427,N_19367);
or U23216 (N_23216,N_19972,N_19428);
nand U23217 (N_23217,N_19929,N_20999);
xnor U23218 (N_23218,N_18219,N_18786);
or U23219 (N_23219,N_18129,N_20580);
nand U23220 (N_23220,N_20540,N_19851);
nand U23221 (N_23221,N_19159,N_19758);
and U23222 (N_23222,N_19685,N_20866);
and U23223 (N_23223,N_19268,N_18308);
xor U23224 (N_23224,N_19920,N_18485);
nand U23225 (N_23225,N_20222,N_20313);
and U23226 (N_23226,N_19598,N_20378);
nor U23227 (N_23227,N_18819,N_20903);
nand U23228 (N_23228,N_20282,N_20338);
or U23229 (N_23229,N_19189,N_19216);
or U23230 (N_23230,N_19344,N_19484);
and U23231 (N_23231,N_18092,N_19448);
xnor U23232 (N_23232,N_20089,N_18054);
nand U23233 (N_23233,N_20660,N_19779);
xor U23234 (N_23234,N_20342,N_18338);
or U23235 (N_23235,N_18533,N_20960);
nand U23236 (N_23236,N_18373,N_19814);
nand U23237 (N_23237,N_19714,N_19394);
nand U23238 (N_23238,N_20662,N_18994);
and U23239 (N_23239,N_18409,N_20372);
nand U23240 (N_23240,N_19528,N_20290);
xor U23241 (N_23241,N_19850,N_18325);
and U23242 (N_23242,N_20291,N_20739);
xnor U23243 (N_23243,N_19959,N_19647);
xor U23244 (N_23244,N_18390,N_18144);
nor U23245 (N_23245,N_20848,N_18920);
nor U23246 (N_23246,N_19223,N_18488);
nor U23247 (N_23247,N_20303,N_19556);
nor U23248 (N_23248,N_20324,N_20813);
xnor U23249 (N_23249,N_19196,N_19583);
and U23250 (N_23250,N_20460,N_20430);
nand U23251 (N_23251,N_20365,N_19671);
xnor U23252 (N_23252,N_20175,N_19143);
nor U23253 (N_23253,N_20839,N_18646);
nand U23254 (N_23254,N_19800,N_19726);
xnor U23255 (N_23255,N_18617,N_19241);
or U23256 (N_23256,N_18939,N_20657);
nor U23257 (N_23257,N_18659,N_20487);
or U23258 (N_23258,N_19450,N_18008);
xnor U23259 (N_23259,N_19032,N_18329);
and U23260 (N_23260,N_19608,N_20559);
and U23261 (N_23261,N_20024,N_19771);
nand U23262 (N_23262,N_19178,N_20582);
or U23263 (N_23263,N_18733,N_18239);
xor U23264 (N_23264,N_20609,N_19986);
nor U23265 (N_23265,N_18553,N_18154);
nor U23266 (N_23266,N_18489,N_20049);
or U23267 (N_23267,N_19403,N_20926);
or U23268 (N_23268,N_18228,N_19994);
or U23269 (N_23269,N_19929,N_19737);
nor U23270 (N_23270,N_18182,N_20487);
nor U23271 (N_23271,N_19432,N_20625);
nor U23272 (N_23272,N_20405,N_19070);
and U23273 (N_23273,N_19062,N_18721);
and U23274 (N_23274,N_19666,N_20408);
nor U23275 (N_23275,N_20812,N_18838);
and U23276 (N_23276,N_19311,N_19899);
xnor U23277 (N_23277,N_19736,N_19903);
nor U23278 (N_23278,N_18951,N_18109);
xnor U23279 (N_23279,N_19316,N_20509);
nand U23280 (N_23280,N_19413,N_20553);
and U23281 (N_23281,N_18897,N_20526);
or U23282 (N_23282,N_19010,N_19941);
nor U23283 (N_23283,N_19128,N_18751);
xor U23284 (N_23284,N_19753,N_19456);
nand U23285 (N_23285,N_18776,N_18680);
xor U23286 (N_23286,N_19040,N_19671);
nor U23287 (N_23287,N_18298,N_19822);
or U23288 (N_23288,N_20089,N_18070);
xnor U23289 (N_23289,N_19428,N_19961);
xnor U23290 (N_23290,N_18800,N_19233);
nor U23291 (N_23291,N_19459,N_18531);
nand U23292 (N_23292,N_20318,N_18483);
or U23293 (N_23293,N_19233,N_20416);
and U23294 (N_23294,N_19388,N_20739);
or U23295 (N_23295,N_18943,N_19905);
nand U23296 (N_23296,N_20382,N_20882);
or U23297 (N_23297,N_19230,N_18381);
nand U23298 (N_23298,N_19405,N_18344);
or U23299 (N_23299,N_18407,N_18191);
xor U23300 (N_23300,N_18192,N_19346);
nor U23301 (N_23301,N_19180,N_20197);
or U23302 (N_23302,N_18795,N_19757);
or U23303 (N_23303,N_19069,N_19505);
xor U23304 (N_23304,N_20645,N_18134);
and U23305 (N_23305,N_20218,N_20766);
and U23306 (N_23306,N_19166,N_18943);
nand U23307 (N_23307,N_19381,N_18077);
nor U23308 (N_23308,N_20321,N_20890);
and U23309 (N_23309,N_20348,N_20390);
xor U23310 (N_23310,N_20045,N_20281);
nor U23311 (N_23311,N_18731,N_19188);
nand U23312 (N_23312,N_19554,N_18709);
xnor U23313 (N_23313,N_19271,N_19198);
and U23314 (N_23314,N_20615,N_18774);
or U23315 (N_23315,N_19224,N_18072);
nor U23316 (N_23316,N_20055,N_19763);
nand U23317 (N_23317,N_20801,N_18921);
nor U23318 (N_23318,N_20497,N_19901);
and U23319 (N_23319,N_20383,N_20555);
and U23320 (N_23320,N_18184,N_18539);
xnor U23321 (N_23321,N_20831,N_19887);
or U23322 (N_23322,N_19029,N_18714);
nand U23323 (N_23323,N_18998,N_19223);
and U23324 (N_23324,N_19902,N_19552);
nand U23325 (N_23325,N_20054,N_19955);
and U23326 (N_23326,N_20371,N_19057);
nand U23327 (N_23327,N_19573,N_18562);
xor U23328 (N_23328,N_20587,N_18799);
and U23329 (N_23329,N_18362,N_19241);
nand U23330 (N_23330,N_18290,N_19947);
xnor U23331 (N_23331,N_19481,N_18362);
or U23332 (N_23332,N_18259,N_19887);
or U23333 (N_23333,N_20881,N_20392);
nand U23334 (N_23334,N_18674,N_19976);
nand U23335 (N_23335,N_18510,N_18939);
or U23336 (N_23336,N_19228,N_20463);
nand U23337 (N_23337,N_19769,N_18883);
nor U23338 (N_23338,N_20105,N_19546);
xor U23339 (N_23339,N_18949,N_18101);
and U23340 (N_23340,N_18603,N_18740);
nor U23341 (N_23341,N_18242,N_20128);
nor U23342 (N_23342,N_20972,N_20421);
nand U23343 (N_23343,N_18296,N_19261);
nand U23344 (N_23344,N_19837,N_20013);
nand U23345 (N_23345,N_18846,N_19800);
nor U23346 (N_23346,N_20552,N_18682);
nand U23347 (N_23347,N_19007,N_18353);
nor U23348 (N_23348,N_19187,N_19498);
and U23349 (N_23349,N_19733,N_19930);
nand U23350 (N_23350,N_18898,N_18306);
and U23351 (N_23351,N_20088,N_18228);
or U23352 (N_23352,N_19962,N_20392);
xor U23353 (N_23353,N_19441,N_18075);
xnor U23354 (N_23354,N_19140,N_19225);
or U23355 (N_23355,N_18935,N_19479);
and U23356 (N_23356,N_19326,N_20062);
or U23357 (N_23357,N_19848,N_18020);
nand U23358 (N_23358,N_19004,N_19392);
nand U23359 (N_23359,N_20280,N_18310);
nor U23360 (N_23360,N_19769,N_18648);
nand U23361 (N_23361,N_18127,N_19913);
and U23362 (N_23362,N_18193,N_19419);
and U23363 (N_23363,N_18433,N_20767);
xnor U23364 (N_23364,N_20902,N_18346);
and U23365 (N_23365,N_18119,N_20750);
nor U23366 (N_23366,N_19028,N_18556);
and U23367 (N_23367,N_20771,N_18661);
and U23368 (N_23368,N_18411,N_20825);
nand U23369 (N_23369,N_19462,N_19948);
or U23370 (N_23370,N_18017,N_18873);
nand U23371 (N_23371,N_20301,N_19777);
nor U23372 (N_23372,N_18907,N_19979);
nor U23373 (N_23373,N_18470,N_20116);
or U23374 (N_23374,N_18904,N_18458);
nand U23375 (N_23375,N_19580,N_18816);
nor U23376 (N_23376,N_19130,N_20260);
nor U23377 (N_23377,N_20875,N_18384);
xor U23378 (N_23378,N_20871,N_18441);
and U23379 (N_23379,N_19421,N_19770);
and U23380 (N_23380,N_19707,N_20742);
or U23381 (N_23381,N_20306,N_19920);
or U23382 (N_23382,N_19928,N_18263);
and U23383 (N_23383,N_20228,N_19472);
xor U23384 (N_23384,N_19037,N_20619);
xnor U23385 (N_23385,N_19085,N_19929);
and U23386 (N_23386,N_18841,N_18734);
xor U23387 (N_23387,N_18973,N_18847);
nor U23388 (N_23388,N_19173,N_19608);
nor U23389 (N_23389,N_20966,N_18834);
xor U23390 (N_23390,N_19496,N_19767);
and U23391 (N_23391,N_18285,N_18861);
nand U23392 (N_23392,N_20085,N_20341);
or U23393 (N_23393,N_18529,N_20897);
nand U23394 (N_23394,N_19908,N_18627);
and U23395 (N_23395,N_19266,N_20887);
or U23396 (N_23396,N_18621,N_19768);
xor U23397 (N_23397,N_19555,N_18620);
or U23398 (N_23398,N_18062,N_19546);
nand U23399 (N_23399,N_18050,N_19847);
or U23400 (N_23400,N_18686,N_19315);
or U23401 (N_23401,N_20389,N_20217);
and U23402 (N_23402,N_18802,N_18104);
nor U23403 (N_23403,N_20635,N_19876);
nand U23404 (N_23404,N_20171,N_18985);
and U23405 (N_23405,N_19279,N_20882);
or U23406 (N_23406,N_20683,N_19748);
or U23407 (N_23407,N_20421,N_18935);
and U23408 (N_23408,N_18983,N_18687);
xor U23409 (N_23409,N_18676,N_18035);
nor U23410 (N_23410,N_19901,N_18637);
nor U23411 (N_23411,N_19431,N_18125);
or U23412 (N_23412,N_20743,N_20582);
xnor U23413 (N_23413,N_18029,N_19441);
nand U23414 (N_23414,N_20637,N_18556);
or U23415 (N_23415,N_20484,N_19422);
nand U23416 (N_23416,N_19218,N_18742);
or U23417 (N_23417,N_19215,N_19487);
xor U23418 (N_23418,N_18404,N_18570);
and U23419 (N_23419,N_20810,N_19347);
xor U23420 (N_23420,N_18170,N_19477);
and U23421 (N_23421,N_20860,N_20942);
and U23422 (N_23422,N_19756,N_20181);
xnor U23423 (N_23423,N_19893,N_20167);
and U23424 (N_23424,N_18148,N_18967);
or U23425 (N_23425,N_19157,N_20542);
xor U23426 (N_23426,N_19535,N_20445);
xor U23427 (N_23427,N_20717,N_18556);
xnor U23428 (N_23428,N_20122,N_18771);
or U23429 (N_23429,N_19436,N_18812);
nor U23430 (N_23430,N_18128,N_19466);
xnor U23431 (N_23431,N_19384,N_19922);
and U23432 (N_23432,N_20794,N_20832);
nand U23433 (N_23433,N_19145,N_19049);
nor U23434 (N_23434,N_20708,N_18654);
nor U23435 (N_23435,N_18515,N_19222);
nand U23436 (N_23436,N_19872,N_19778);
nor U23437 (N_23437,N_20340,N_19039);
nor U23438 (N_23438,N_19703,N_19020);
or U23439 (N_23439,N_19445,N_19644);
or U23440 (N_23440,N_19636,N_20591);
and U23441 (N_23441,N_20661,N_20642);
and U23442 (N_23442,N_19319,N_19129);
nor U23443 (N_23443,N_19319,N_18276);
xor U23444 (N_23444,N_19191,N_20476);
or U23445 (N_23445,N_20807,N_19272);
nand U23446 (N_23446,N_18935,N_20684);
nor U23447 (N_23447,N_18112,N_20954);
nand U23448 (N_23448,N_18385,N_19517);
xor U23449 (N_23449,N_20414,N_18165);
nand U23450 (N_23450,N_18397,N_18589);
nand U23451 (N_23451,N_18600,N_18033);
or U23452 (N_23452,N_20931,N_18184);
nor U23453 (N_23453,N_19036,N_18156);
or U23454 (N_23454,N_18955,N_18362);
nor U23455 (N_23455,N_19751,N_19546);
nand U23456 (N_23456,N_20953,N_18304);
xnor U23457 (N_23457,N_19955,N_19177);
nand U23458 (N_23458,N_18724,N_20237);
nor U23459 (N_23459,N_19533,N_20742);
and U23460 (N_23460,N_20619,N_20474);
nor U23461 (N_23461,N_18224,N_20884);
or U23462 (N_23462,N_18097,N_18188);
and U23463 (N_23463,N_20674,N_20350);
nor U23464 (N_23464,N_18794,N_19385);
or U23465 (N_23465,N_20930,N_20210);
nor U23466 (N_23466,N_19142,N_19188);
and U23467 (N_23467,N_18918,N_20154);
nor U23468 (N_23468,N_20631,N_20840);
nor U23469 (N_23469,N_20078,N_18489);
nand U23470 (N_23470,N_18374,N_19828);
nor U23471 (N_23471,N_19843,N_19606);
xor U23472 (N_23472,N_19650,N_19211);
and U23473 (N_23473,N_20908,N_19112);
nor U23474 (N_23474,N_19803,N_20220);
xor U23475 (N_23475,N_18312,N_20152);
and U23476 (N_23476,N_19199,N_19590);
and U23477 (N_23477,N_19011,N_18906);
nor U23478 (N_23478,N_20678,N_19852);
xnor U23479 (N_23479,N_19176,N_19540);
or U23480 (N_23480,N_18023,N_18337);
nor U23481 (N_23481,N_19692,N_20543);
or U23482 (N_23482,N_18948,N_19375);
and U23483 (N_23483,N_19442,N_19791);
and U23484 (N_23484,N_19167,N_18526);
and U23485 (N_23485,N_19450,N_19827);
nand U23486 (N_23486,N_18722,N_20118);
xnor U23487 (N_23487,N_18974,N_20047);
xnor U23488 (N_23488,N_19705,N_20206);
and U23489 (N_23489,N_18747,N_19769);
nor U23490 (N_23490,N_19825,N_18324);
and U23491 (N_23491,N_19034,N_18921);
xnor U23492 (N_23492,N_19065,N_19142);
nor U23493 (N_23493,N_20811,N_18594);
or U23494 (N_23494,N_19727,N_20311);
and U23495 (N_23495,N_18469,N_20223);
nand U23496 (N_23496,N_18583,N_18391);
xor U23497 (N_23497,N_19103,N_20741);
xor U23498 (N_23498,N_19398,N_19122);
and U23499 (N_23499,N_19611,N_19005);
and U23500 (N_23500,N_19962,N_20606);
nand U23501 (N_23501,N_20031,N_18822);
nor U23502 (N_23502,N_19203,N_18371);
or U23503 (N_23503,N_20905,N_19363);
nand U23504 (N_23504,N_19385,N_19560);
and U23505 (N_23505,N_20617,N_20536);
nor U23506 (N_23506,N_19087,N_20934);
or U23507 (N_23507,N_19523,N_20162);
nand U23508 (N_23508,N_18971,N_18702);
xor U23509 (N_23509,N_19127,N_19517);
and U23510 (N_23510,N_20504,N_20809);
and U23511 (N_23511,N_20799,N_20352);
and U23512 (N_23512,N_20489,N_18213);
nand U23513 (N_23513,N_20480,N_20967);
nand U23514 (N_23514,N_18590,N_20713);
nand U23515 (N_23515,N_18590,N_19817);
and U23516 (N_23516,N_18740,N_19602);
nand U23517 (N_23517,N_20338,N_18643);
and U23518 (N_23518,N_20394,N_20313);
nand U23519 (N_23519,N_20333,N_20082);
nand U23520 (N_23520,N_20207,N_20479);
xor U23521 (N_23521,N_20112,N_19626);
or U23522 (N_23522,N_20575,N_18652);
and U23523 (N_23523,N_19717,N_19964);
nand U23524 (N_23524,N_18481,N_20784);
xnor U23525 (N_23525,N_18772,N_19613);
nor U23526 (N_23526,N_19981,N_19770);
and U23527 (N_23527,N_18648,N_20710);
and U23528 (N_23528,N_20430,N_18077);
nor U23529 (N_23529,N_19512,N_18319);
xnor U23530 (N_23530,N_18959,N_18681);
or U23531 (N_23531,N_18347,N_18858);
nand U23532 (N_23532,N_19924,N_20271);
and U23533 (N_23533,N_19577,N_20450);
xnor U23534 (N_23534,N_19997,N_18181);
nand U23535 (N_23535,N_18295,N_20164);
nor U23536 (N_23536,N_19924,N_18584);
and U23537 (N_23537,N_19936,N_18485);
nand U23538 (N_23538,N_19934,N_18762);
and U23539 (N_23539,N_20834,N_18404);
nand U23540 (N_23540,N_18811,N_19215);
or U23541 (N_23541,N_19257,N_18933);
or U23542 (N_23542,N_19340,N_19076);
and U23543 (N_23543,N_20024,N_20691);
or U23544 (N_23544,N_18694,N_20120);
or U23545 (N_23545,N_18851,N_20645);
or U23546 (N_23546,N_18410,N_19789);
nand U23547 (N_23547,N_20086,N_19127);
or U23548 (N_23548,N_18730,N_20931);
xnor U23549 (N_23549,N_20086,N_18933);
nand U23550 (N_23550,N_18494,N_19626);
or U23551 (N_23551,N_19669,N_19597);
nand U23552 (N_23552,N_20908,N_20598);
and U23553 (N_23553,N_18655,N_18798);
xnor U23554 (N_23554,N_18801,N_18438);
and U23555 (N_23555,N_19704,N_19972);
and U23556 (N_23556,N_18439,N_19350);
nand U23557 (N_23557,N_20886,N_20172);
nand U23558 (N_23558,N_20909,N_20554);
xor U23559 (N_23559,N_20232,N_18829);
xor U23560 (N_23560,N_19491,N_18687);
xor U23561 (N_23561,N_20748,N_18561);
or U23562 (N_23562,N_18741,N_18299);
or U23563 (N_23563,N_19150,N_19409);
nor U23564 (N_23564,N_18865,N_20177);
or U23565 (N_23565,N_19556,N_20821);
xnor U23566 (N_23566,N_20664,N_19360);
or U23567 (N_23567,N_20906,N_18294);
and U23568 (N_23568,N_20470,N_18923);
or U23569 (N_23569,N_20289,N_20274);
nor U23570 (N_23570,N_18781,N_20223);
xnor U23571 (N_23571,N_19295,N_18281);
nand U23572 (N_23572,N_20152,N_18099);
xnor U23573 (N_23573,N_19115,N_18118);
nor U23574 (N_23574,N_20878,N_18596);
nor U23575 (N_23575,N_20742,N_19218);
and U23576 (N_23576,N_20731,N_18467);
nor U23577 (N_23577,N_18306,N_20724);
and U23578 (N_23578,N_19541,N_18219);
nand U23579 (N_23579,N_18893,N_18971);
nor U23580 (N_23580,N_19111,N_18910);
nor U23581 (N_23581,N_18256,N_19671);
xor U23582 (N_23582,N_20947,N_20880);
nor U23583 (N_23583,N_19023,N_20342);
nor U23584 (N_23584,N_20488,N_19564);
nor U23585 (N_23585,N_18663,N_18806);
nand U23586 (N_23586,N_19631,N_20198);
or U23587 (N_23587,N_20196,N_20544);
and U23588 (N_23588,N_20355,N_19288);
nor U23589 (N_23589,N_20986,N_20116);
nor U23590 (N_23590,N_19298,N_19799);
xnor U23591 (N_23591,N_18213,N_20972);
nand U23592 (N_23592,N_19210,N_19462);
nand U23593 (N_23593,N_19690,N_18839);
nand U23594 (N_23594,N_18960,N_18755);
nand U23595 (N_23595,N_20893,N_19620);
or U23596 (N_23596,N_20437,N_19356);
xnor U23597 (N_23597,N_18095,N_19131);
and U23598 (N_23598,N_19900,N_19770);
nor U23599 (N_23599,N_18661,N_18797);
xor U23600 (N_23600,N_20503,N_18884);
or U23601 (N_23601,N_19334,N_19451);
xor U23602 (N_23602,N_19071,N_18518);
or U23603 (N_23603,N_19293,N_19548);
xor U23604 (N_23604,N_20281,N_20378);
and U23605 (N_23605,N_19798,N_20145);
xor U23606 (N_23606,N_20149,N_18545);
xnor U23607 (N_23607,N_20649,N_19961);
nor U23608 (N_23608,N_19881,N_19491);
nand U23609 (N_23609,N_18004,N_19820);
nor U23610 (N_23610,N_19032,N_18881);
nor U23611 (N_23611,N_18070,N_20403);
xnor U23612 (N_23612,N_20830,N_19413);
xor U23613 (N_23613,N_20027,N_18308);
nand U23614 (N_23614,N_18964,N_19388);
and U23615 (N_23615,N_20647,N_19661);
and U23616 (N_23616,N_19382,N_18041);
xor U23617 (N_23617,N_20707,N_18827);
and U23618 (N_23618,N_19724,N_20539);
and U23619 (N_23619,N_19892,N_20045);
nand U23620 (N_23620,N_18385,N_19305);
xor U23621 (N_23621,N_19604,N_20698);
and U23622 (N_23622,N_19599,N_19480);
and U23623 (N_23623,N_18134,N_19192);
or U23624 (N_23624,N_20083,N_20720);
nand U23625 (N_23625,N_20611,N_18805);
nor U23626 (N_23626,N_20863,N_18495);
nor U23627 (N_23627,N_19359,N_20280);
nor U23628 (N_23628,N_19627,N_18835);
and U23629 (N_23629,N_19533,N_18440);
xnor U23630 (N_23630,N_19381,N_20173);
or U23631 (N_23631,N_19770,N_20320);
xor U23632 (N_23632,N_20597,N_20576);
nor U23633 (N_23633,N_18664,N_20979);
nand U23634 (N_23634,N_20782,N_18693);
xnor U23635 (N_23635,N_19619,N_18633);
nand U23636 (N_23636,N_18266,N_20225);
nor U23637 (N_23637,N_20333,N_19436);
xnor U23638 (N_23638,N_18873,N_18289);
and U23639 (N_23639,N_20425,N_20356);
or U23640 (N_23640,N_18175,N_18026);
and U23641 (N_23641,N_18292,N_19883);
and U23642 (N_23642,N_18171,N_18250);
nand U23643 (N_23643,N_18007,N_18986);
and U23644 (N_23644,N_19787,N_18030);
nand U23645 (N_23645,N_19346,N_18091);
and U23646 (N_23646,N_19012,N_20652);
and U23647 (N_23647,N_18182,N_19101);
xor U23648 (N_23648,N_18518,N_20232);
xnor U23649 (N_23649,N_20404,N_19336);
and U23650 (N_23650,N_19112,N_18661);
or U23651 (N_23651,N_18365,N_19241);
nand U23652 (N_23652,N_18936,N_18635);
xnor U23653 (N_23653,N_19731,N_18819);
nand U23654 (N_23654,N_20707,N_19860);
xor U23655 (N_23655,N_19980,N_19918);
or U23656 (N_23656,N_20936,N_20747);
nor U23657 (N_23657,N_18538,N_19131);
xor U23658 (N_23658,N_18246,N_20669);
and U23659 (N_23659,N_19200,N_18744);
or U23660 (N_23660,N_19617,N_18492);
and U23661 (N_23661,N_19417,N_18664);
or U23662 (N_23662,N_18058,N_19136);
nand U23663 (N_23663,N_20265,N_20261);
nor U23664 (N_23664,N_20619,N_19782);
or U23665 (N_23665,N_18551,N_18120);
xnor U23666 (N_23666,N_20109,N_20491);
nor U23667 (N_23667,N_20889,N_19489);
or U23668 (N_23668,N_19822,N_18738);
nand U23669 (N_23669,N_20534,N_19510);
xnor U23670 (N_23670,N_20962,N_19191);
nor U23671 (N_23671,N_20134,N_18818);
xnor U23672 (N_23672,N_20380,N_18201);
or U23673 (N_23673,N_19728,N_20444);
and U23674 (N_23674,N_20036,N_20734);
nand U23675 (N_23675,N_18032,N_18772);
xor U23676 (N_23676,N_18412,N_19048);
and U23677 (N_23677,N_20663,N_19830);
nand U23678 (N_23678,N_19228,N_20157);
nor U23679 (N_23679,N_19449,N_19959);
nor U23680 (N_23680,N_18792,N_18800);
and U23681 (N_23681,N_18805,N_20531);
xnor U23682 (N_23682,N_20809,N_18315);
or U23683 (N_23683,N_20942,N_19785);
or U23684 (N_23684,N_18182,N_20434);
nor U23685 (N_23685,N_18406,N_19501);
xor U23686 (N_23686,N_18529,N_18056);
or U23687 (N_23687,N_20403,N_20364);
nor U23688 (N_23688,N_18904,N_20399);
nand U23689 (N_23689,N_19355,N_19516);
nand U23690 (N_23690,N_18698,N_18469);
and U23691 (N_23691,N_20391,N_19637);
or U23692 (N_23692,N_20026,N_20361);
nor U23693 (N_23693,N_18569,N_19721);
nand U23694 (N_23694,N_20969,N_20884);
nand U23695 (N_23695,N_19935,N_19444);
and U23696 (N_23696,N_20633,N_18790);
xnor U23697 (N_23697,N_19069,N_18200);
xnor U23698 (N_23698,N_19911,N_18109);
nor U23699 (N_23699,N_18356,N_18499);
nand U23700 (N_23700,N_20584,N_19752);
nand U23701 (N_23701,N_20108,N_19573);
and U23702 (N_23702,N_19507,N_19937);
xor U23703 (N_23703,N_20487,N_18118);
or U23704 (N_23704,N_20098,N_20540);
xor U23705 (N_23705,N_18233,N_18837);
and U23706 (N_23706,N_18090,N_18536);
xor U23707 (N_23707,N_18114,N_19394);
xor U23708 (N_23708,N_19678,N_18302);
or U23709 (N_23709,N_20310,N_18188);
and U23710 (N_23710,N_20015,N_20231);
and U23711 (N_23711,N_18011,N_19395);
nand U23712 (N_23712,N_19618,N_20196);
nand U23713 (N_23713,N_18690,N_20298);
and U23714 (N_23714,N_18090,N_18419);
nor U23715 (N_23715,N_18649,N_20334);
nor U23716 (N_23716,N_20884,N_19480);
nand U23717 (N_23717,N_18459,N_18156);
xnor U23718 (N_23718,N_18310,N_20388);
xnor U23719 (N_23719,N_19062,N_20052);
nand U23720 (N_23720,N_20909,N_18215);
nor U23721 (N_23721,N_18867,N_18427);
xnor U23722 (N_23722,N_18110,N_19626);
xnor U23723 (N_23723,N_20036,N_19232);
and U23724 (N_23724,N_18257,N_19782);
nor U23725 (N_23725,N_18618,N_18267);
nor U23726 (N_23726,N_20650,N_19815);
and U23727 (N_23727,N_18808,N_19954);
xor U23728 (N_23728,N_19756,N_19257);
xnor U23729 (N_23729,N_18919,N_20119);
nand U23730 (N_23730,N_20064,N_19497);
nand U23731 (N_23731,N_18481,N_19952);
or U23732 (N_23732,N_20182,N_18990);
or U23733 (N_23733,N_19666,N_18026);
nand U23734 (N_23734,N_20331,N_18348);
xnor U23735 (N_23735,N_18582,N_20248);
xor U23736 (N_23736,N_20917,N_18985);
and U23737 (N_23737,N_20310,N_18372);
nand U23738 (N_23738,N_19427,N_18011);
or U23739 (N_23739,N_20586,N_20548);
xnor U23740 (N_23740,N_19125,N_20938);
xor U23741 (N_23741,N_20414,N_20357);
xor U23742 (N_23742,N_18306,N_19471);
or U23743 (N_23743,N_19910,N_19559);
nand U23744 (N_23744,N_19787,N_20492);
xor U23745 (N_23745,N_19266,N_19586);
nand U23746 (N_23746,N_18257,N_20165);
xor U23747 (N_23747,N_19010,N_19711);
and U23748 (N_23748,N_18155,N_18151);
xnor U23749 (N_23749,N_20951,N_19209);
nand U23750 (N_23750,N_19414,N_19848);
or U23751 (N_23751,N_20738,N_20677);
and U23752 (N_23752,N_19648,N_20265);
and U23753 (N_23753,N_18250,N_20309);
or U23754 (N_23754,N_19290,N_20898);
nand U23755 (N_23755,N_19273,N_18603);
nand U23756 (N_23756,N_18397,N_18674);
nor U23757 (N_23757,N_18176,N_19501);
nor U23758 (N_23758,N_20368,N_19261);
nand U23759 (N_23759,N_20621,N_18786);
and U23760 (N_23760,N_19221,N_20802);
nor U23761 (N_23761,N_18330,N_18343);
nor U23762 (N_23762,N_19098,N_20432);
xor U23763 (N_23763,N_19230,N_19074);
xnor U23764 (N_23764,N_20334,N_18342);
and U23765 (N_23765,N_20336,N_20750);
and U23766 (N_23766,N_20609,N_20370);
xnor U23767 (N_23767,N_18299,N_18303);
xor U23768 (N_23768,N_20201,N_18177);
nand U23769 (N_23769,N_20874,N_18687);
and U23770 (N_23770,N_19184,N_18266);
nor U23771 (N_23771,N_20494,N_19114);
or U23772 (N_23772,N_19787,N_18682);
and U23773 (N_23773,N_19240,N_20172);
xnor U23774 (N_23774,N_20527,N_19402);
and U23775 (N_23775,N_19446,N_19148);
nand U23776 (N_23776,N_18286,N_18216);
xor U23777 (N_23777,N_19858,N_18003);
xor U23778 (N_23778,N_18817,N_18545);
nor U23779 (N_23779,N_19383,N_18477);
or U23780 (N_23780,N_19887,N_19624);
or U23781 (N_23781,N_18931,N_20684);
and U23782 (N_23782,N_19206,N_19246);
and U23783 (N_23783,N_19231,N_20334);
nand U23784 (N_23784,N_18217,N_20079);
nor U23785 (N_23785,N_19464,N_20388);
nand U23786 (N_23786,N_18839,N_18937);
nor U23787 (N_23787,N_18215,N_20553);
and U23788 (N_23788,N_20843,N_19616);
nand U23789 (N_23789,N_18340,N_19181);
or U23790 (N_23790,N_20523,N_18756);
and U23791 (N_23791,N_18961,N_18910);
and U23792 (N_23792,N_20737,N_20962);
xor U23793 (N_23793,N_18943,N_19193);
or U23794 (N_23794,N_19704,N_20460);
or U23795 (N_23795,N_20245,N_19784);
xnor U23796 (N_23796,N_19772,N_19108);
nand U23797 (N_23797,N_18964,N_20645);
and U23798 (N_23798,N_18882,N_18742);
nor U23799 (N_23799,N_19631,N_20757);
and U23800 (N_23800,N_20613,N_18601);
nand U23801 (N_23801,N_20502,N_20250);
xnor U23802 (N_23802,N_18836,N_18955);
xnor U23803 (N_23803,N_20622,N_20165);
and U23804 (N_23804,N_20950,N_20173);
xnor U23805 (N_23805,N_20874,N_20193);
and U23806 (N_23806,N_18956,N_19026);
nor U23807 (N_23807,N_18452,N_18115);
or U23808 (N_23808,N_18223,N_20730);
nor U23809 (N_23809,N_19431,N_20880);
nand U23810 (N_23810,N_18137,N_18450);
nor U23811 (N_23811,N_19522,N_19541);
or U23812 (N_23812,N_20693,N_20633);
and U23813 (N_23813,N_20085,N_19089);
nor U23814 (N_23814,N_20376,N_18714);
xor U23815 (N_23815,N_19562,N_19892);
and U23816 (N_23816,N_19884,N_20163);
and U23817 (N_23817,N_20570,N_18088);
and U23818 (N_23818,N_19339,N_18738);
and U23819 (N_23819,N_19849,N_18209);
and U23820 (N_23820,N_19623,N_20021);
nor U23821 (N_23821,N_20674,N_18536);
nor U23822 (N_23822,N_19785,N_18223);
and U23823 (N_23823,N_19193,N_18413);
xnor U23824 (N_23824,N_19728,N_20454);
xor U23825 (N_23825,N_19500,N_18827);
and U23826 (N_23826,N_19858,N_19475);
and U23827 (N_23827,N_18530,N_18039);
and U23828 (N_23828,N_19635,N_20971);
or U23829 (N_23829,N_19439,N_19429);
nand U23830 (N_23830,N_18825,N_18635);
nand U23831 (N_23831,N_20943,N_20458);
nor U23832 (N_23832,N_20579,N_18960);
or U23833 (N_23833,N_20964,N_18242);
nor U23834 (N_23834,N_20734,N_19577);
or U23835 (N_23835,N_18497,N_19316);
nand U23836 (N_23836,N_19351,N_18304);
nor U23837 (N_23837,N_20259,N_20949);
nand U23838 (N_23838,N_18444,N_19815);
xor U23839 (N_23839,N_19453,N_19920);
nor U23840 (N_23840,N_19650,N_20538);
and U23841 (N_23841,N_19007,N_19789);
or U23842 (N_23842,N_18048,N_20614);
nand U23843 (N_23843,N_19135,N_20257);
nor U23844 (N_23844,N_20471,N_19877);
nand U23845 (N_23845,N_18642,N_18103);
nand U23846 (N_23846,N_19138,N_20437);
and U23847 (N_23847,N_18293,N_19999);
xnor U23848 (N_23848,N_20534,N_19301);
xor U23849 (N_23849,N_19145,N_18610);
xnor U23850 (N_23850,N_19566,N_19159);
nand U23851 (N_23851,N_19652,N_19642);
nor U23852 (N_23852,N_20089,N_19967);
and U23853 (N_23853,N_20151,N_20650);
nor U23854 (N_23854,N_19799,N_19374);
nor U23855 (N_23855,N_20007,N_18279);
and U23856 (N_23856,N_20282,N_20768);
or U23857 (N_23857,N_20282,N_19418);
xnor U23858 (N_23858,N_19486,N_19503);
xor U23859 (N_23859,N_20967,N_18853);
xor U23860 (N_23860,N_20476,N_20886);
xor U23861 (N_23861,N_18648,N_20648);
and U23862 (N_23862,N_20013,N_19448);
nor U23863 (N_23863,N_18493,N_20455);
and U23864 (N_23864,N_18947,N_19232);
and U23865 (N_23865,N_20444,N_20221);
and U23866 (N_23866,N_18631,N_18464);
xnor U23867 (N_23867,N_20286,N_18425);
nor U23868 (N_23868,N_18895,N_20751);
nand U23869 (N_23869,N_20039,N_19310);
or U23870 (N_23870,N_20799,N_20896);
or U23871 (N_23871,N_18290,N_20990);
or U23872 (N_23872,N_20538,N_20390);
and U23873 (N_23873,N_19043,N_20338);
and U23874 (N_23874,N_19997,N_18797);
and U23875 (N_23875,N_19201,N_18451);
and U23876 (N_23876,N_18248,N_18304);
or U23877 (N_23877,N_20773,N_19720);
nor U23878 (N_23878,N_19811,N_18604);
and U23879 (N_23879,N_19406,N_19296);
or U23880 (N_23880,N_19640,N_18509);
or U23881 (N_23881,N_19173,N_20690);
xor U23882 (N_23882,N_19599,N_18062);
nor U23883 (N_23883,N_20980,N_19834);
nor U23884 (N_23884,N_19572,N_18816);
nand U23885 (N_23885,N_18000,N_18446);
xor U23886 (N_23886,N_18226,N_20051);
or U23887 (N_23887,N_20226,N_19823);
and U23888 (N_23888,N_19901,N_20413);
or U23889 (N_23889,N_20088,N_20037);
nand U23890 (N_23890,N_18407,N_18984);
and U23891 (N_23891,N_20392,N_20955);
and U23892 (N_23892,N_20287,N_18340);
nand U23893 (N_23893,N_19195,N_18883);
or U23894 (N_23894,N_20544,N_20798);
nor U23895 (N_23895,N_19515,N_18446);
nor U23896 (N_23896,N_18805,N_19414);
nor U23897 (N_23897,N_18562,N_18071);
nand U23898 (N_23898,N_19176,N_20886);
xnor U23899 (N_23899,N_19399,N_18845);
and U23900 (N_23900,N_19058,N_19110);
nand U23901 (N_23901,N_19790,N_20028);
nand U23902 (N_23902,N_20629,N_19579);
and U23903 (N_23903,N_19355,N_20134);
nand U23904 (N_23904,N_18209,N_20734);
nand U23905 (N_23905,N_19820,N_19301);
xnor U23906 (N_23906,N_19420,N_18402);
nand U23907 (N_23907,N_19005,N_20578);
nand U23908 (N_23908,N_20777,N_18685);
xor U23909 (N_23909,N_18076,N_19781);
or U23910 (N_23910,N_20298,N_19876);
nand U23911 (N_23911,N_18139,N_18589);
nand U23912 (N_23912,N_19808,N_20386);
and U23913 (N_23913,N_19015,N_20490);
or U23914 (N_23914,N_18768,N_19765);
nor U23915 (N_23915,N_18343,N_20936);
or U23916 (N_23916,N_19592,N_18649);
nand U23917 (N_23917,N_19899,N_20059);
xnor U23918 (N_23918,N_18126,N_18156);
nand U23919 (N_23919,N_20158,N_18804);
xor U23920 (N_23920,N_19685,N_20085);
nor U23921 (N_23921,N_20046,N_19604);
and U23922 (N_23922,N_20702,N_20241);
xor U23923 (N_23923,N_19572,N_19457);
nor U23924 (N_23924,N_18615,N_19796);
and U23925 (N_23925,N_19902,N_19576);
and U23926 (N_23926,N_19547,N_18597);
and U23927 (N_23927,N_18441,N_20562);
nand U23928 (N_23928,N_20459,N_20549);
and U23929 (N_23929,N_18099,N_18880);
nand U23930 (N_23930,N_19825,N_19069);
and U23931 (N_23931,N_20409,N_20457);
or U23932 (N_23932,N_20715,N_20467);
nand U23933 (N_23933,N_19405,N_18763);
and U23934 (N_23934,N_20946,N_20850);
nand U23935 (N_23935,N_18143,N_19580);
nor U23936 (N_23936,N_20287,N_20927);
xor U23937 (N_23937,N_19698,N_20024);
nor U23938 (N_23938,N_20154,N_19282);
or U23939 (N_23939,N_19259,N_20866);
nand U23940 (N_23940,N_19768,N_18813);
and U23941 (N_23941,N_19989,N_18342);
nand U23942 (N_23942,N_19211,N_18317);
xnor U23943 (N_23943,N_18696,N_18440);
nor U23944 (N_23944,N_19047,N_18376);
nand U23945 (N_23945,N_19441,N_18330);
and U23946 (N_23946,N_18374,N_20533);
xor U23947 (N_23947,N_20332,N_18161);
nand U23948 (N_23948,N_20960,N_20280);
xor U23949 (N_23949,N_20561,N_18152);
and U23950 (N_23950,N_19599,N_20115);
or U23951 (N_23951,N_19731,N_20118);
and U23952 (N_23952,N_18679,N_18849);
nor U23953 (N_23953,N_19652,N_19173);
xor U23954 (N_23954,N_19583,N_20896);
and U23955 (N_23955,N_20953,N_19387);
nand U23956 (N_23956,N_19773,N_19763);
and U23957 (N_23957,N_20196,N_20219);
nor U23958 (N_23958,N_18262,N_18766);
nor U23959 (N_23959,N_18137,N_20076);
nand U23960 (N_23960,N_19996,N_20247);
or U23961 (N_23961,N_20910,N_19140);
and U23962 (N_23962,N_19147,N_19154);
xnor U23963 (N_23963,N_18590,N_20481);
nand U23964 (N_23964,N_18957,N_18596);
nor U23965 (N_23965,N_18575,N_18323);
or U23966 (N_23966,N_19920,N_18703);
or U23967 (N_23967,N_19631,N_19336);
or U23968 (N_23968,N_19787,N_20191);
nor U23969 (N_23969,N_19438,N_20337);
xnor U23970 (N_23970,N_18314,N_18363);
xnor U23971 (N_23971,N_20144,N_18954);
nand U23972 (N_23972,N_20574,N_20669);
or U23973 (N_23973,N_20839,N_18200);
or U23974 (N_23974,N_19867,N_18675);
nor U23975 (N_23975,N_18872,N_20504);
nor U23976 (N_23976,N_20957,N_20053);
xnor U23977 (N_23977,N_19019,N_18945);
nand U23978 (N_23978,N_20632,N_18144);
xor U23979 (N_23979,N_19696,N_19737);
nand U23980 (N_23980,N_19477,N_20352);
or U23981 (N_23981,N_20383,N_18564);
or U23982 (N_23982,N_19078,N_20025);
xor U23983 (N_23983,N_19434,N_18993);
nand U23984 (N_23984,N_18448,N_18554);
nand U23985 (N_23985,N_19871,N_20555);
nor U23986 (N_23986,N_18341,N_20151);
nor U23987 (N_23987,N_20738,N_19590);
or U23988 (N_23988,N_20937,N_19272);
nor U23989 (N_23989,N_19287,N_19720);
nand U23990 (N_23990,N_20059,N_18876);
and U23991 (N_23991,N_19793,N_19480);
xnor U23992 (N_23992,N_18043,N_19951);
or U23993 (N_23993,N_20401,N_18727);
nand U23994 (N_23994,N_20036,N_18176);
and U23995 (N_23995,N_19784,N_19315);
nand U23996 (N_23996,N_19783,N_19178);
xnor U23997 (N_23997,N_18829,N_18807);
nand U23998 (N_23998,N_19859,N_20490);
and U23999 (N_23999,N_18771,N_18754);
xnor U24000 (N_24000,N_23696,N_23918);
nand U24001 (N_24001,N_21832,N_23639);
nor U24002 (N_24002,N_21535,N_21584);
nor U24003 (N_24003,N_22254,N_21516);
and U24004 (N_24004,N_23675,N_21747);
and U24005 (N_24005,N_23564,N_21794);
xnor U24006 (N_24006,N_23504,N_23016);
nand U24007 (N_24007,N_21543,N_23673);
xnor U24008 (N_24008,N_22148,N_22162);
nor U24009 (N_24009,N_22319,N_22851);
or U24010 (N_24010,N_21190,N_21672);
nor U24011 (N_24011,N_21382,N_21362);
nor U24012 (N_24012,N_21618,N_23969);
and U24013 (N_24013,N_23135,N_21941);
nand U24014 (N_24014,N_21592,N_22527);
nand U24015 (N_24015,N_22607,N_21448);
nor U24016 (N_24016,N_23864,N_21748);
nor U24017 (N_24017,N_22272,N_21069);
and U24018 (N_24018,N_21761,N_23351);
nor U24019 (N_24019,N_21716,N_22292);
nor U24020 (N_24020,N_21368,N_23129);
nor U24021 (N_24021,N_21329,N_22082);
or U24022 (N_24022,N_23746,N_23621);
or U24023 (N_24023,N_23807,N_22230);
xnor U24024 (N_24024,N_22391,N_21176);
nand U24025 (N_24025,N_22641,N_22328);
nor U24026 (N_24026,N_22260,N_22504);
or U24027 (N_24027,N_22951,N_21731);
or U24028 (N_24028,N_21287,N_23837);
xor U24029 (N_24029,N_23790,N_21180);
nor U24030 (N_24030,N_23556,N_21870);
nor U24031 (N_24031,N_23769,N_23430);
and U24032 (N_24032,N_23501,N_21299);
xnor U24033 (N_24033,N_22117,N_23578);
and U24034 (N_24034,N_22021,N_23065);
or U24035 (N_24035,N_22635,N_22928);
or U24036 (N_24036,N_23882,N_23455);
xor U24037 (N_24037,N_21943,N_23829);
nand U24038 (N_24038,N_21578,N_23147);
nand U24039 (N_24039,N_21415,N_23684);
xnor U24040 (N_24040,N_23298,N_22445);
or U24041 (N_24041,N_23678,N_21637);
and U24042 (N_24042,N_22190,N_21890);
nor U24043 (N_24043,N_22070,N_21946);
nor U24044 (N_24044,N_21239,N_23938);
and U24045 (N_24045,N_22772,N_23984);
xnor U24046 (N_24046,N_21458,N_21040);
nor U24047 (N_24047,N_21151,N_21929);
and U24048 (N_24048,N_23432,N_21325);
nor U24049 (N_24049,N_23749,N_22521);
nand U24050 (N_24050,N_23560,N_21529);
nand U24051 (N_24051,N_23895,N_23723);
xnor U24052 (N_24052,N_21878,N_23617);
and U24053 (N_24053,N_23354,N_23728);
and U24054 (N_24054,N_21928,N_21704);
xnor U24055 (N_24055,N_22047,N_23857);
xnor U24056 (N_24056,N_21266,N_21787);
or U24057 (N_24057,N_23263,N_22582);
nor U24058 (N_24058,N_22662,N_22933);
nand U24059 (N_24059,N_21046,N_21285);
nand U24060 (N_24060,N_23277,N_21322);
or U24061 (N_24061,N_21392,N_23220);
nand U24062 (N_24062,N_23656,N_22197);
nand U24063 (N_24063,N_22247,N_22996);
or U24064 (N_24064,N_22845,N_21348);
xor U24065 (N_24065,N_23862,N_21453);
or U24066 (N_24066,N_21948,N_22303);
nand U24067 (N_24067,N_23246,N_23706);
and U24068 (N_24068,N_23628,N_22330);
or U24069 (N_24069,N_21791,N_23497);
nor U24070 (N_24070,N_21260,N_22136);
and U24071 (N_24071,N_23954,N_23572);
xor U24072 (N_24072,N_21998,N_22693);
nand U24073 (N_24073,N_21923,N_22010);
or U24074 (N_24074,N_22747,N_21682);
nand U24075 (N_24075,N_21616,N_23204);
nor U24076 (N_24076,N_22156,N_21188);
xor U24077 (N_24077,N_23633,N_23577);
nand U24078 (N_24078,N_23883,N_21739);
and U24079 (N_24079,N_23152,N_21455);
nand U24080 (N_24080,N_23308,N_22433);
or U24081 (N_24081,N_21252,N_22726);
nor U24082 (N_24082,N_21214,N_22222);
nor U24083 (N_24083,N_22114,N_21119);
nor U24084 (N_24084,N_21251,N_21953);
nand U24085 (N_24085,N_22627,N_22837);
xor U24086 (N_24086,N_21875,N_23653);
nor U24087 (N_24087,N_23665,N_23717);
nand U24088 (N_24088,N_22874,N_23978);
nor U24089 (N_24089,N_22231,N_23319);
nor U24090 (N_24090,N_21595,N_23571);
nor U24091 (N_24091,N_21658,N_23553);
nand U24092 (N_24092,N_23171,N_22967);
nand U24093 (N_24093,N_23608,N_23921);
nand U24094 (N_24094,N_22903,N_23975);
or U24095 (N_24095,N_22728,N_23485);
nor U24096 (N_24096,N_22606,N_22334);
or U24097 (N_24097,N_23652,N_21416);
nor U24098 (N_24098,N_23048,N_23218);
xnor U24099 (N_24099,N_21961,N_22949);
and U24100 (N_24100,N_23264,N_23378);
nor U24101 (N_24101,N_22408,N_21937);
nor U24102 (N_24102,N_21861,N_21924);
or U24103 (N_24103,N_22137,N_21717);
nand U24104 (N_24104,N_23757,N_23916);
and U24105 (N_24105,N_21031,N_22895);
xnor U24106 (N_24106,N_21017,N_23278);
or U24107 (N_24107,N_22807,N_23899);
nand U24108 (N_24108,N_22357,N_21311);
nand U24109 (N_24109,N_23813,N_23067);
and U24110 (N_24110,N_22628,N_23262);
nand U24111 (N_24111,N_23116,N_23035);
and U24112 (N_24112,N_23959,N_23090);
and U24113 (N_24113,N_22192,N_22171);
or U24114 (N_24114,N_21141,N_23976);
or U24115 (N_24115,N_21697,N_21819);
xor U24116 (N_24116,N_23960,N_22346);
nor U24117 (N_24117,N_22769,N_23846);
and U24118 (N_24118,N_21118,N_23335);
xnor U24119 (N_24119,N_22699,N_23407);
nand U24120 (N_24120,N_23655,N_23691);
or U24121 (N_24121,N_23915,N_23603);
xnor U24122 (N_24122,N_23986,N_23231);
nand U24123 (N_24123,N_23327,N_21737);
xor U24124 (N_24124,N_23042,N_23050);
and U24125 (N_24125,N_21891,N_21625);
nor U24126 (N_24126,N_22109,N_21706);
nor U24127 (N_24127,N_21511,N_23440);
xor U24128 (N_24128,N_23227,N_21892);
nand U24129 (N_24129,N_21075,N_23239);
nand U24130 (N_24130,N_22487,N_23206);
or U24131 (N_24131,N_23436,N_21883);
xor U24132 (N_24132,N_22207,N_22760);
and U24133 (N_24133,N_23352,N_23459);
nor U24134 (N_24134,N_22108,N_22266);
xor U24135 (N_24135,N_22348,N_21154);
nor U24136 (N_24136,N_23654,N_21234);
and U24137 (N_24137,N_22615,N_23437);
and U24138 (N_24138,N_23318,N_21184);
and U24139 (N_24139,N_22263,N_21855);
or U24140 (N_24140,N_22539,N_23242);
xor U24141 (N_24141,N_23020,N_22926);
nor U24142 (N_24142,N_21408,N_22520);
or U24143 (N_24143,N_22923,N_22495);
nor U24144 (N_24144,N_21806,N_23953);
or U24145 (N_24145,N_21396,N_22738);
and U24146 (N_24146,N_23950,N_23531);
or U24147 (N_24147,N_21499,N_22857);
nor U24148 (N_24148,N_22887,N_21241);
or U24149 (N_24149,N_21312,N_23592);
or U24150 (N_24150,N_22469,N_23506);
xnor U24151 (N_24151,N_22096,N_23126);
nor U24152 (N_24152,N_23333,N_21104);
and U24153 (N_24153,N_23397,N_22869);
nor U24154 (N_24154,N_22203,N_23060);
xnor U24155 (N_24155,N_21345,N_23205);
nand U24156 (N_24156,N_21050,N_23366);
nand U24157 (N_24157,N_23568,N_23527);
xnor U24158 (N_24158,N_22396,N_22358);
or U24159 (N_24159,N_21060,N_21821);
and U24160 (N_24160,N_22649,N_21420);
nor U24161 (N_24161,N_22675,N_21997);
or U24162 (N_24162,N_21082,N_22161);
nor U24163 (N_24163,N_21236,N_22172);
xnor U24164 (N_24164,N_22663,N_23386);
or U24165 (N_24165,N_23533,N_21403);
xor U24166 (N_24166,N_22033,N_21183);
and U24167 (N_24167,N_21170,N_21983);
or U24168 (N_24168,N_22905,N_23207);
nor U24169 (N_24169,N_21874,N_22743);
and U24170 (N_24170,N_22473,N_22121);
or U24171 (N_24171,N_23461,N_21011);
or U24172 (N_24172,N_21033,N_21256);
and U24173 (N_24173,N_21440,N_23269);
or U24174 (N_24174,N_22523,N_23481);
nand U24175 (N_24175,N_23783,N_23258);
nor U24176 (N_24176,N_23086,N_21800);
nand U24177 (N_24177,N_22604,N_21581);
nand U24178 (N_24178,N_23845,N_22555);
xor U24179 (N_24179,N_23478,N_21845);
and U24180 (N_24180,N_22689,N_23620);
xnor U24181 (N_24181,N_22101,N_22638);
and U24182 (N_24182,N_23186,N_21942);
nand U24183 (N_24183,N_23694,N_23519);
nand U24184 (N_24184,N_23767,N_22794);
or U24185 (N_24185,N_21365,N_22339);
or U24186 (N_24186,N_21156,N_21675);
or U24187 (N_24187,N_21776,N_21958);
nor U24188 (N_24188,N_22127,N_23816);
xnor U24189 (N_24189,N_21985,N_23663);
nand U24190 (N_24190,N_21566,N_22763);
nor U24191 (N_24191,N_22583,N_21292);
nand U24192 (N_24192,N_23237,N_21038);
nand U24193 (N_24193,N_23994,N_21539);
and U24194 (N_24194,N_22703,N_21277);
and U24195 (N_24195,N_23989,N_23228);
and U24196 (N_24196,N_23838,N_23192);
xor U24197 (N_24197,N_23772,N_23569);
and U24198 (N_24198,N_21555,N_23713);
nand U24199 (N_24199,N_22786,N_23700);
xnor U24200 (N_24200,N_22016,N_23834);
nand U24201 (N_24201,N_23629,N_21494);
nand U24202 (N_24202,N_23662,N_22170);
nand U24203 (N_24203,N_22911,N_21579);
nand U24204 (N_24204,N_23342,N_21444);
or U24205 (N_24205,N_23222,N_23765);
xnor U24206 (N_24206,N_23013,N_23064);
nor U24207 (N_24207,N_21871,N_23551);
and U24208 (N_24208,N_21117,N_23869);
xnor U24209 (N_24209,N_21564,N_21102);
and U24210 (N_24210,N_22361,N_23529);
or U24211 (N_24211,N_23474,N_23898);
or U24212 (N_24212,N_23505,N_22425);
xnor U24213 (N_24213,N_21810,N_23539);
and U24214 (N_24214,N_21058,N_22100);
nor U24215 (N_24215,N_23089,N_21201);
and U24216 (N_24216,N_22018,N_21351);
and U24217 (N_24217,N_22955,N_23260);
nand U24218 (N_24218,N_23049,N_22378);
nand U24219 (N_24219,N_23840,N_23203);
nor U24220 (N_24220,N_22655,N_21096);
and U24221 (N_24221,N_22516,N_23646);
nand U24222 (N_24222,N_22574,N_23842);
nor U24223 (N_24223,N_22512,N_21041);
nand U24224 (N_24224,N_21346,N_22347);
nor U24225 (N_24225,N_22145,N_21081);
xor U24226 (N_24226,N_21160,N_23518);
nor U24227 (N_24227,N_22572,N_22372);
nor U24228 (N_24228,N_21729,N_22936);
or U24229 (N_24229,N_23624,N_22983);
or U24230 (N_24230,N_22065,N_21386);
nand U24231 (N_24231,N_23712,N_21931);
nor U24232 (N_24232,N_23347,N_23359);
xnor U24233 (N_24233,N_22915,N_23151);
and U24234 (N_24234,N_21247,N_22733);
or U24235 (N_24235,N_21418,N_21614);
or U24236 (N_24236,N_21713,N_21417);
and U24237 (N_24237,N_23053,N_22988);
or U24238 (N_24238,N_23515,N_23516);
nand U24239 (N_24239,N_22669,N_21908);
nor U24240 (N_24240,N_22106,N_21061);
nand U24241 (N_24241,N_21037,N_22842);
and U24242 (N_24242,N_22797,N_21628);
xor U24243 (N_24243,N_23725,N_22024);
and U24244 (N_24244,N_21509,N_23146);
xor U24245 (N_24245,N_22731,N_22467);
or U24246 (N_24246,N_23120,N_23810);
xnor U24247 (N_24247,N_22723,N_23784);
nand U24248 (N_24248,N_22300,N_21865);
nand U24249 (N_24249,N_21710,N_22614);
or U24250 (N_24250,N_23174,N_21823);
nor U24251 (N_24251,N_21064,N_22213);
nand U24252 (N_24252,N_22630,N_23693);
and U24253 (N_24253,N_23949,N_23737);
xnor U24254 (N_24254,N_22317,N_23296);
or U24255 (N_24255,N_21841,N_22461);
xnor U24256 (N_24256,N_23348,N_23877);
nand U24257 (N_24257,N_21390,N_22793);
nor U24258 (N_24258,N_21824,N_21836);
nor U24259 (N_24259,N_21079,N_22687);
or U24260 (N_24260,N_21634,N_21626);
xnor U24261 (N_24261,N_23026,N_22563);
and U24262 (N_24262,N_22633,N_21816);
xor U24263 (N_24263,N_22414,N_23900);
xnor U24264 (N_24264,N_23072,N_22449);
nor U24265 (N_24265,N_23598,N_22506);
or U24266 (N_24266,N_22700,N_23188);
xor U24267 (N_24267,N_21438,N_21853);
nor U24268 (N_24268,N_22363,N_23362);
or U24269 (N_24269,N_22907,N_22560);
xor U24270 (N_24270,N_22287,N_22830);
or U24271 (N_24271,N_22864,N_22778);
xnor U24272 (N_24272,N_21080,N_21827);
nor U24273 (N_24273,N_22128,N_23685);
xnor U24274 (N_24274,N_22402,N_22636);
nor U24275 (N_24275,N_23894,N_22052);
and U24276 (N_24276,N_21629,N_21758);
nor U24277 (N_24277,N_22881,N_22997);
or U24278 (N_24278,N_21089,N_22817);
nand U24279 (N_24279,N_21221,N_23099);
or U24280 (N_24280,N_22113,N_22546);
or U24281 (N_24281,N_22569,N_23763);
nand U24282 (N_24282,N_22011,N_23910);
or U24283 (N_24283,N_21261,N_23558);
or U24284 (N_24284,N_21240,N_22694);
xnor U24285 (N_24285,N_23643,N_23486);
or U24286 (N_24286,N_22316,N_23615);
xor U24287 (N_24287,N_23881,N_22087);
or U24288 (N_24288,N_21431,N_21215);
or U24289 (N_24289,N_21515,N_23219);
or U24290 (N_24290,N_23261,N_23555);
nand U24291 (N_24291,N_21849,N_21763);
nand U24292 (N_24292,N_22773,N_21206);
and U24293 (N_24293,N_23626,N_23044);
or U24294 (N_24294,N_23526,N_22532);
nor U24295 (N_24295,N_22775,N_21217);
xor U24296 (N_24296,N_21934,N_23704);
and U24297 (N_24297,N_22494,N_22825);
or U24298 (N_24298,N_21182,N_23886);
or U24299 (N_24299,N_23401,N_21767);
xor U24300 (N_24300,N_22322,N_23136);
and U24301 (N_24301,N_23159,N_22354);
nand U24302 (N_24302,N_21968,N_23730);
xor U24303 (N_24303,N_21964,N_22152);
nand U24304 (N_24304,N_23051,N_21361);
nand U24305 (N_24305,N_22344,N_22884);
nor U24306 (N_24306,N_21447,N_23332);
xnor U24307 (N_24307,N_21088,N_23311);
or U24308 (N_24308,N_21880,N_23280);
xnor U24309 (N_24309,N_21620,N_21213);
and U24310 (N_24310,N_21210,N_23415);
and U24311 (N_24311,N_22729,N_22716);
or U24312 (N_24312,N_23443,N_22673);
xor U24313 (N_24313,N_22525,N_22882);
nor U24314 (N_24314,N_22169,N_22939);
xor U24315 (N_24315,N_22745,N_22737);
nand U24316 (N_24316,N_23304,N_21834);
or U24317 (N_24317,N_23500,N_22455);
or U24318 (N_24318,N_22919,N_21817);
or U24319 (N_24319,N_21355,N_23750);
xnor U24320 (N_24320,N_23538,N_21043);
xor U24321 (N_24321,N_22540,N_21332);
nor U24322 (N_24322,N_23449,N_22659);
nor U24323 (N_24323,N_22125,N_22086);
xor U24324 (N_24324,N_21021,N_22522);
and U24325 (N_24325,N_21254,N_23111);
nor U24326 (N_24326,N_21839,N_22019);
nand U24327 (N_24327,N_21072,N_22576);
and U24328 (N_24328,N_23144,N_21436);
or U24329 (N_24329,N_21779,N_21813);
xnor U24330 (N_24330,N_21619,N_22844);
nand U24331 (N_24331,N_23047,N_21569);
or U24332 (N_24332,N_23101,N_23075);
nand U24333 (N_24333,N_21967,N_21280);
and U24334 (N_24334,N_23305,N_22877);
xor U24335 (N_24335,N_21424,N_21410);
nand U24336 (N_24336,N_21385,N_23389);
or U24337 (N_24337,N_21955,N_23779);
nor U24338 (N_24338,N_22674,N_22995);
nand U24339 (N_24339,N_21301,N_23887);
or U24340 (N_24340,N_23683,N_21973);
or U24341 (N_24341,N_21657,N_23912);
or U24342 (N_24342,N_22173,N_23388);
xor U24343 (N_24343,N_22083,N_23173);
nor U24344 (N_24344,N_22430,N_21684);
xnor U24345 (N_24345,N_22686,N_21570);
xnor U24346 (N_24346,N_23891,N_21427);
or U24347 (N_24347,N_23282,N_22243);
nand U24348 (N_24348,N_22284,N_22032);
nor U24349 (N_24349,N_21127,N_22258);
nand U24350 (N_24350,N_23524,N_23306);
nand U24351 (N_24351,N_22329,N_21318);
and U24352 (N_24352,N_23991,N_23917);
nor U24353 (N_24353,N_22643,N_23800);
nand U24354 (N_24354,N_21111,N_22538);
xnor U24355 (N_24355,N_22820,N_21762);
or U24356 (N_24356,N_23119,N_22601);
nor U24357 (N_24357,N_21901,N_23480);
and U24358 (N_24358,N_22376,N_21723);
or U24359 (N_24359,N_22557,N_23574);
nor U24360 (N_24360,N_22337,N_22352);
nand U24361 (N_24361,N_21186,N_23454);
nor U24362 (N_24362,N_23863,N_22095);
or U24363 (N_24363,N_21708,N_23931);
nor U24364 (N_24364,N_22834,N_23365);
nand U24365 (N_24365,N_22298,N_21143);
xor U24366 (N_24366,N_22634,N_22696);
xor U24367 (N_24367,N_22921,N_22041);
xor U24368 (N_24368,N_21015,N_21822);
and U24369 (N_24369,N_23326,N_21700);
and U24370 (N_24370,N_21464,N_23372);
and U24371 (N_24371,N_22447,N_23233);
xor U24372 (N_24372,N_23300,N_23934);
xor U24373 (N_24373,N_21411,N_21711);
and U24374 (N_24374,N_21594,N_21425);
or U24375 (N_24375,N_23802,N_21087);
xnor U24376 (N_24376,N_21587,N_21722);
nor U24377 (N_24377,N_22476,N_23128);
nor U24378 (N_24378,N_22832,N_21608);
xor U24379 (N_24379,N_21725,N_22474);
nor U24380 (N_24380,N_21652,N_23856);
or U24381 (N_24381,N_22885,N_22039);
nand U24382 (N_24382,N_22484,N_21485);
and U24383 (N_24383,N_23382,N_22226);
nor U24384 (N_24384,N_22577,N_21381);
xor U24385 (N_24385,N_21323,N_22974);
nor U24386 (N_24386,N_21357,N_23627);
xnor U24387 (N_24387,N_23631,N_22390);
nor U24388 (N_24388,N_21617,N_21679);
and U24389 (N_24389,N_23092,N_22288);
nand U24390 (N_24390,N_23105,N_22701);
nand U24391 (N_24391,N_22736,N_22411);
xor U24392 (N_24392,N_22573,N_22306);
and U24393 (N_24393,N_21778,N_22448);
or U24394 (N_24394,N_22237,N_21740);
or U24395 (N_24395,N_22973,N_21898);
and U24396 (N_24396,N_22478,N_21507);
nand U24397 (N_24397,N_21641,N_23535);
xor U24398 (N_24398,N_22341,N_22558);
and U24399 (N_24399,N_22592,N_22074);
and U24400 (N_24400,N_22088,N_23434);
and U24401 (N_24401,N_23199,N_23732);
or U24402 (N_24402,N_22941,N_21030);
or U24403 (N_24403,N_23573,N_21987);
and U24404 (N_24404,N_22417,N_21622);
or U24405 (N_24405,N_23880,N_21733);
nor U24406 (N_24406,N_23266,N_22790);
nand U24407 (N_24407,N_21523,N_23875);
xnor U24408 (N_24408,N_23114,N_22900);
and U24409 (N_24409,N_23272,N_23177);
or U24410 (N_24410,N_23328,N_21772);
and U24411 (N_24411,N_21765,N_21712);
or U24412 (N_24412,N_22286,N_22454);
and U24413 (N_24413,N_23602,N_23477);
xnor U24414 (N_24414,N_22970,N_23906);
and U24415 (N_24415,N_21294,N_22945);
or U24416 (N_24416,N_22862,N_21388);
xnor U24417 (N_24417,N_23036,N_21720);
or U24418 (N_24418,N_23447,N_22924);
xnor U24419 (N_24419,N_21687,N_22925);
nand U24420 (N_24420,N_21460,N_22922);
or U24421 (N_24421,N_23141,N_22684);
or U24422 (N_24422,N_22759,N_22228);
nor U24423 (N_24423,N_23212,N_21225);
nand U24424 (N_24424,N_22429,N_21468);
and U24425 (N_24425,N_23927,N_23541);
xor U24426 (N_24426,N_21429,N_21273);
xnor U24427 (N_24427,N_21475,N_23786);
nand U24428 (N_24428,N_23438,N_22964);
nor U24429 (N_24429,N_22890,N_23285);
or U24430 (N_24430,N_22751,N_23343);
xor U24431 (N_24431,N_21175,N_23017);
nor U24432 (N_24432,N_23510,N_23364);
or U24433 (N_24433,N_21423,N_23297);
and U24434 (N_24434,N_21848,N_23517);
nand U24435 (N_24435,N_23429,N_23698);
nor U24436 (N_24436,N_21873,N_22822);
nand U24437 (N_24437,N_22710,N_23812);
xnor U24438 (N_24438,N_22727,N_22394);
and U24439 (N_24439,N_21812,N_21177);
and U24440 (N_24440,N_22665,N_23672);
nor U24441 (N_24441,N_22761,N_22840);
or U24442 (N_24442,N_21231,N_23736);
nor U24443 (N_24443,N_21915,N_21913);
nor U24444 (N_24444,N_23873,N_23705);
and U24445 (N_24445,N_21520,N_22119);
xnor U24446 (N_24446,N_22513,N_22819);
or U24447 (N_24447,N_23399,N_21734);
nand U24448 (N_24448,N_22456,N_21588);
or U24449 (N_24449,N_21056,N_22764);
nand U24450 (N_24450,N_23563,N_22301);
or U24451 (N_24451,N_23210,N_21450);
and U24452 (N_24452,N_22508,N_21042);
xor U24453 (N_24453,N_21583,N_23391);
and U24454 (N_24454,N_22014,N_22757);
or U24455 (N_24455,N_22690,N_23855);
or U24456 (N_24456,N_23033,N_22276);
or U24457 (N_24457,N_21370,N_23012);
and U24458 (N_24458,N_22575,N_22957);
nor U24459 (N_24459,N_22481,N_23742);
xnor U24460 (N_24460,N_22815,N_23940);
nor U24461 (N_24461,N_23970,N_23121);
nor U24462 (N_24462,N_23901,N_21589);
xor U24463 (N_24463,N_23396,N_23793);
and U24464 (N_24464,N_21728,N_22003);
xnor U24465 (N_24465,N_21971,N_23641);
or U24466 (N_24466,N_21905,N_23274);
nand U24467 (N_24467,N_23544,N_23371);
nor U24468 (N_24468,N_23988,N_22556);
nor U24469 (N_24469,N_22979,N_21798);
nand U24470 (N_24470,N_22360,N_23079);
xnor U24471 (N_24471,N_23238,N_21991);
xnor U24472 (N_24472,N_21642,N_22533);
xnor U24473 (N_24473,N_21130,N_23083);
or U24474 (N_24474,N_22383,N_23489);
or U24475 (N_24475,N_23309,N_21216);
nand U24476 (N_24476,N_22368,N_22289);
nand U24477 (N_24477,N_23279,N_23502);
xor U24478 (N_24478,N_23252,N_22424);
and U24479 (N_24479,N_21926,N_21498);
or U24480 (N_24480,N_22215,N_21391);
and U24481 (N_24481,N_21744,N_22158);
xnor U24482 (N_24482,N_23747,N_23611);
nand U24483 (N_24483,N_21894,N_21367);
and U24484 (N_24484,N_22917,N_22415);
or U24485 (N_24485,N_21877,N_21736);
and U24486 (N_24486,N_22722,N_21495);
and U24487 (N_24487,N_21092,N_21203);
nor U24488 (N_24488,N_21412,N_23464);
or U24489 (N_24489,N_21532,N_23346);
nor U24490 (N_24490,N_21406,N_21164);
and U24491 (N_24491,N_23292,N_22236);
and U24492 (N_24492,N_21648,N_21063);
nor U24493 (N_24493,N_21567,N_21545);
nor U24494 (N_24494,N_21128,N_21785);
xnor U24495 (N_24495,N_22587,N_23699);
nor U24496 (N_24496,N_23741,N_22992);
or U24497 (N_24497,N_21990,N_22972);
or U24498 (N_24498,N_22501,N_22962);
or U24499 (N_24499,N_21666,N_23613);
nor U24500 (N_24500,N_22327,N_23878);
nor U24501 (N_24501,N_23589,N_21477);
or U24502 (N_24502,N_21497,N_21524);
nor U24503 (N_24503,N_21268,N_22404);
xor U24504 (N_24504,N_22401,N_22488);
xnor U24505 (N_24505,N_23166,N_23968);
or U24506 (N_24506,N_23010,N_22631);
and U24507 (N_24507,N_22123,N_22971);
xnor U24508 (N_24508,N_22518,N_21680);
nor U24509 (N_24509,N_22045,N_22261);
nand U24510 (N_24510,N_21223,N_23007);
and U24511 (N_24511,N_21482,N_21930);
and U24512 (N_24512,N_21344,N_22253);
nor U24513 (N_24513,N_21897,N_22167);
nand U24514 (N_24514,N_21544,N_22739);
and U24515 (N_24515,N_22406,N_23738);
nor U24516 (N_24516,N_22283,N_23567);
nand U24517 (N_24517,N_21047,N_22749);
nor U24518 (N_24518,N_23462,N_23134);
nor U24519 (N_24519,N_22201,N_23761);
nand U24520 (N_24520,N_21333,N_21850);
xnor U24521 (N_24521,N_21109,N_23295);
and U24522 (N_24522,N_21781,N_21550);
nand U24523 (N_24523,N_21920,N_21709);
nand U24524 (N_24524,N_21646,N_21083);
xor U24525 (N_24525,N_22589,N_22613);
xor U24526 (N_24526,N_23123,N_21777);
nand U24527 (N_24527,N_22318,N_22485);
nor U24528 (N_24528,N_21965,N_21756);
nand U24529 (N_24529,N_21363,N_23139);
xor U24530 (N_24530,N_23680,N_23823);
nor U24531 (N_24531,N_22680,N_21445);
or U24532 (N_24532,N_23154,N_22661);
or U24533 (N_24533,N_23648,N_23708);
and U24534 (N_24534,N_21463,N_21159);
and U24535 (N_24535,N_23835,N_23385);
nand U24536 (N_24536,N_23193,N_21910);
nand U24537 (N_24537,N_21327,N_21243);
nor U24538 (N_24538,N_21563,N_22715);
and U24539 (N_24539,N_22085,N_21107);
or U24540 (N_24540,N_21889,N_21378);
and U24541 (N_24541,N_23302,N_23850);
or U24542 (N_24542,N_23339,N_23250);
xnor U24543 (N_24543,N_22821,N_21054);
nor U24544 (N_24544,N_22332,N_22600);
xnor U24545 (N_24545,N_21144,N_23425);
nand U24546 (N_24546,N_22529,N_22122);
and U24547 (N_24547,N_23795,N_22709);
or U24548 (N_24548,N_23496,N_23257);
nor U24549 (N_24549,N_21242,N_22938);
and U24550 (N_24550,N_23605,N_22846);
xor U24551 (N_24551,N_21685,N_23005);
nor U24552 (N_24552,N_23027,N_21707);
nand U24553 (N_24553,N_21289,N_21694);
xnor U24554 (N_24554,N_23865,N_21724);
nor U24555 (N_24555,N_21496,N_21461);
and U24556 (N_24556,N_23316,N_23132);
nand U24557 (N_24557,N_23637,N_23094);
and U24558 (N_24558,N_22718,N_21631);
nor U24559 (N_24559,N_23791,N_22989);
and U24560 (N_24560,N_22075,N_21833);
xor U24561 (N_24561,N_22492,N_22077);
or U24562 (N_24562,N_22452,N_22954);
or U24563 (N_24563,N_22963,N_21784);
nand U24564 (N_24564,N_23587,N_23373);
xor U24565 (N_24565,N_21501,N_21258);
nand U24566 (N_24566,N_21828,N_23866);
nand U24567 (N_24567,N_22894,N_21246);
nand U24568 (N_24568,N_22622,N_21632);
nor U24569 (N_24569,N_23068,N_21212);
xnor U24570 (N_24570,N_23720,N_21966);
xnor U24571 (N_24571,N_21574,N_22420);
or U24572 (N_24572,N_22566,N_22421);
nor U24573 (N_24573,N_22505,N_22326);
and U24574 (N_24574,N_21229,N_21936);
and U24575 (N_24575,N_23775,N_23087);
and U24576 (N_24576,N_21293,N_21989);
or U24577 (N_24577,N_22343,N_21753);
xor U24578 (N_24578,N_22199,N_21743);
nand U24579 (N_24579,N_21112,N_21996);
nor U24580 (N_24580,N_23039,N_21962);
nand U24581 (N_24581,N_22398,N_23201);
nand U24582 (N_24582,N_23057,N_22705);
and U24583 (N_24583,N_23902,N_23043);
nor U24584 (N_24584,N_21195,N_23697);
nor U24585 (N_24585,N_23175,N_23923);
xor U24586 (N_24586,N_23453,N_22629);
or U24587 (N_24587,N_23284,N_23457);
or U24588 (N_24588,N_22860,N_23759);
nor U24589 (N_24589,N_23456,N_22181);
and U24590 (N_24590,N_23286,N_22697);
xnor U24591 (N_24591,N_21992,N_22302);
or U24592 (N_24592,N_22581,N_23532);
or U24593 (N_24593,N_22564,N_22632);
xor U24594 (N_24594,N_21283,N_23659);
nand U24595 (N_24595,N_22027,N_23619);
nand U24596 (N_24596,N_23998,N_22942);
and U24597 (N_24597,N_23289,N_21066);
nand U24598 (N_24598,N_21586,N_23642);
nor U24599 (N_24599,N_23125,N_21149);
or U24600 (N_24600,N_21027,N_22943);
and U24601 (N_24601,N_21308,N_22852);
nand U24602 (N_24602,N_21237,N_22355);
and U24603 (N_24603,N_22839,N_23408);
and U24604 (N_24604,N_21670,N_23191);
or U24605 (N_24605,N_22756,N_21558);
xor U24606 (N_24606,N_23625,N_22782);
xor U24607 (N_24607,N_23872,N_21196);
or U24608 (N_24608,N_23824,N_23215);
nand U24609 (N_24609,N_23833,N_21275);
nand U24610 (N_24610,N_21590,N_22559);
xnor U24611 (N_24611,N_23780,N_23341);
nor U24612 (N_24612,N_23782,N_23113);
nand U24613 (N_24613,N_21886,N_22285);
nor U24614 (N_24614,N_22545,N_22711);
nand U24615 (N_24615,N_23904,N_21207);
or U24616 (N_24616,N_22366,N_21405);
nand U24617 (N_24617,N_23848,N_21265);
or U24618 (N_24618,N_22889,N_22090);
and U24619 (N_24619,N_22618,N_21178);
nor U24620 (N_24620,N_23666,N_21353);
or U24621 (N_24621,N_23350,N_22295);
nand U24622 (N_24622,N_23200,N_22080);
nor U24623 (N_24623,N_23547,N_21338);
or U24624 (N_24624,N_21259,N_22160);
nor U24625 (N_24625,N_21531,N_21655);
or U24626 (N_24626,N_23417,N_21944);
xor U24627 (N_24627,N_21219,N_22177);
nor U24628 (N_24628,N_21899,N_21960);
and U24629 (N_24629,N_23690,N_21826);
nor U24630 (N_24630,N_22281,N_21337);
nand U24631 (N_24631,N_22342,N_22994);
nor U24632 (N_24632,N_21358,N_23187);
nand U24633 (N_24633,N_21483,N_21023);
or U24634 (N_24634,N_21059,N_21211);
nand U24635 (N_24635,N_21123,N_22071);
and U24636 (N_24636,N_21389,N_22471);
or U24637 (N_24637,N_23511,N_22653);
and U24638 (N_24638,N_21305,N_23888);
xor U24639 (N_24639,N_22112,N_22946);
nor U24640 (N_24640,N_21419,N_23828);
xor U24641 (N_24641,N_21097,N_21609);
or U24642 (N_24642,N_21858,N_23240);
and U24643 (N_24643,N_21270,N_21471);
nand U24644 (N_24644,N_21683,N_23821);
nor U24645 (N_24645,N_22110,N_22683);
and U24646 (N_24646,N_21250,N_23768);
xnor U24647 (N_24647,N_21014,N_23392);
nor U24648 (N_24648,N_23576,N_22565);
and U24649 (N_24649,N_22528,N_23349);
nand U24650 (N_24650,N_23463,N_23424);
or U24651 (N_24651,N_21380,N_22969);
nand U24652 (N_24652,N_21788,N_22423);
nor U24653 (N_24653,N_21844,N_22927);
nand U24654 (N_24654,N_22233,N_21451);
or U24655 (N_24655,N_23788,N_21169);
or U24656 (N_24656,N_21220,N_21792);
xor U24657 (N_24657,N_21918,N_21230);
and U24658 (N_24658,N_21939,N_21094);
or U24659 (N_24659,N_21639,N_22791);
and U24660 (N_24660,N_23826,N_23508);
xnor U24661 (N_24661,N_23383,N_22947);
nand U24662 (N_24662,N_21528,N_21384);
xnor U24663 (N_24663,N_22278,N_23623);
xnor U24664 (N_24664,N_21029,N_22744);
or U24665 (N_24665,N_21959,N_22990);
xnor U24666 (N_24666,N_23145,N_21024);
and U24667 (N_24667,N_23607,N_23964);
or U24668 (N_24668,N_21982,N_23330);
xor U24669 (N_24669,N_22800,N_23892);
and U24670 (N_24670,N_23830,N_21470);
and U24671 (N_24671,N_23164,N_23980);
nor U24672 (N_24672,N_21101,N_21661);
or U24673 (N_24673,N_23046,N_23593);
and U24674 (N_24674,N_22060,N_21479);
nand U24675 (N_24675,N_23411,N_21802);
xor U24676 (N_24676,N_23803,N_21248);
and U24677 (N_24677,N_21076,N_21818);
nor U24678 (N_24678,N_23374,N_23808);
nor U24679 (N_24679,N_23729,N_21155);
xor U24680 (N_24680,N_23423,N_22888);
nand U24681 (N_24681,N_22380,N_22026);
nor U24682 (N_24682,N_21902,N_21291);
and U24683 (N_24683,N_21297,N_21738);
and U24684 (N_24684,N_22325,N_23676);
nand U24685 (N_24685,N_21932,N_23952);
nand U24686 (N_24686,N_23112,N_21122);
nor U24687 (N_24687,N_21703,N_22395);
xnor U24688 (N_24688,N_22274,N_23925);
or U24689 (N_24689,N_21377,N_22652);
nand U24690 (N_24690,N_22486,N_21115);
nor U24691 (N_24691,N_22142,N_21264);
or U24692 (N_24692,N_22509,N_21830);
nand U24693 (N_24693,N_22812,N_22388);
or U24694 (N_24694,N_21533,N_22400);
or U24695 (N_24695,N_23321,N_21397);
and U24696 (N_24696,N_21341,N_22297);
xor U24697 (N_24697,N_21842,N_22296);
and U24698 (N_24698,N_21466,N_22164);
and U24699 (N_24699,N_23479,N_22067);
and U24700 (N_24700,N_21715,N_21020);
nand U24701 (N_24701,N_22210,N_21852);
or U24702 (N_24702,N_22766,N_21263);
or U24703 (N_24703,N_21198,N_22410);
or U24704 (N_24704,N_22216,N_21073);
xor U24705 (N_24705,N_22536,N_23874);
and U24706 (N_24706,N_23475,N_23194);
xnor U24707 (N_24707,N_23983,N_22913);
nor U24708 (N_24708,N_22367,N_22179);
or U24709 (N_24709,N_22554,N_22847);
or U24710 (N_24710,N_22000,N_23731);
nor U24711 (N_24711,N_22124,N_22440);
nor U24712 (N_24712,N_21591,N_22184);
nand U24713 (N_24713,N_23011,N_22748);
nor U24714 (N_24714,N_23522,N_22843);
xnor U24715 (N_24715,N_22750,N_22658);
nor U24716 (N_24716,N_22498,N_22755);
nor U24717 (N_24717,N_23003,N_23841);
xnor U24718 (N_24718,N_21002,N_21662);
xnor U24719 (N_24719,N_21957,N_23937);
nor U24720 (N_24720,N_21185,N_21068);
nand U24721 (N_24721,N_22816,N_21754);
or U24722 (N_24722,N_23929,N_23601);
or U24723 (N_24723,N_22570,N_21200);
nor U24724 (N_24724,N_22975,N_21009);
or U24725 (N_24725,N_22138,N_23426);
nor U24726 (N_24726,N_22431,N_22140);
nor U24727 (N_24727,N_22350,N_21437);
and U24728 (N_24728,N_22340,N_23649);
nor U24729 (N_24729,N_22891,N_22012);
xor U24730 (N_24730,N_23368,N_23009);
xor U24731 (N_24731,N_23727,N_22929);
or U24732 (N_24732,N_21244,N_21452);
nor U24733 (N_24733,N_22829,N_22858);
or U24734 (N_24734,N_23419,N_21395);
nand U24735 (N_24735,N_21552,N_22541);
and U24736 (N_24736,N_22165,N_23836);
nand U24737 (N_24737,N_21859,N_22054);
nand U24738 (N_24738,N_21369,N_22702);
or U24739 (N_24739,N_21347,N_22553);
and U24740 (N_24740,N_21222,N_23973);
nor U24741 (N_24741,N_21150,N_21487);
nand U24742 (N_24742,N_22666,N_21008);
and U24743 (N_24743,N_21493,N_23861);
or U24744 (N_24744,N_22578,N_21310);
nand U24745 (N_24745,N_21433,N_22706);
and U24746 (N_24746,N_21189,N_23255);
nand U24747 (N_24747,N_21522,N_21663);
nand U24748 (N_24748,N_21227,N_22868);
or U24749 (N_24749,N_21490,N_22439);
nor U24750 (N_24750,N_21677,N_21714);
nor U24751 (N_24751,N_22444,N_22084);
nor U24752 (N_24752,N_21199,N_21257);
or U24753 (N_24753,N_21665,N_22044);
nand U24754 (N_24754,N_21300,N_22186);
xnor U24755 (N_24755,N_22500,N_23446);
nand U24756 (N_24756,N_23418,N_21862);
xnor U24757 (N_24757,N_22902,N_21596);
xor U24758 (N_24758,N_22517,N_21746);
xnor U24759 (N_24759,N_22803,N_23760);
nor U24760 (N_24760,N_22904,N_22379);
nor U24761 (N_24761,N_22005,N_23582);
xor U24762 (N_24762,N_22602,N_21922);
xor U24763 (N_24763,N_23491,N_23271);
and U24764 (N_24764,N_23163,N_22450);
nand U24765 (N_24765,N_23584,N_23202);
and U24766 (N_24766,N_21521,N_22503);
nor U24767 (N_24767,N_23528,N_22092);
nor U24768 (N_24768,N_22893,N_22310);
or U24769 (N_24769,N_22212,N_21925);
nor U24770 (N_24770,N_23165,N_23103);
and U24771 (N_24771,N_23847,N_21400);
or U24772 (N_24772,N_21409,N_22912);
or U24773 (N_24773,N_22001,N_23692);
or U24774 (N_24774,N_21012,N_23428);
nand U24775 (N_24775,N_22382,N_21055);
nor U24776 (N_24776,N_22813,N_23667);
xor U24777 (N_24777,N_21640,N_21272);
or U24778 (N_24778,N_23811,N_23562);
nor U24779 (N_24779,N_21636,N_21110);
or U24780 (N_24780,N_22134,N_23338);
xnor U24781 (N_24781,N_23859,N_23689);
nand U24782 (N_24782,N_21091,N_23579);
nand U24783 (N_24783,N_22648,N_23657);
xnor U24784 (N_24784,N_21449,N_23038);
nand U24785 (N_24785,N_23358,N_23061);
or U24786 (N_24786,N_23379,N_23465);
and U24787 (N_24787,N_23082,N_23645);
xor U24788 (N_24788,N_21978,N_23403);
nand U24789 (N_24789,N_21768,N_21446);
or U24790 (N_24790,N_21638,N_23548);
and U24791 (N_24791,N_21808,N_23507);
or U24792 (N_24792,N_22784,N_22034);
nor U24793 (N_24793,N_23041,N_22025);
xor U24794 (N_24794,N_22460,N_21360);
or U24795 (N_24795,N_21457,N_22187);
xnor U24796 (N_24796,N_22626,N_21313);
or U24797 (N_24797,N_23924,N_21194);
xor U24798 (N_24798,N_22029,N_22753);
nand U24799 (N_24799,N_23018,N_23357);
or U24800 (N_24800,N_21402,N_22654);
xor U24801 (N_24801,N_21651,N_23198);
nand U24802 (N_24802,N_21090,N_22056);
nor U24803 (N_24803,N_23226,N_23922);
and U24804 (N_24804,N_23074,N_21296);
nor U24805 (N_24805,N_21557,N_21290);
or U24806 (N_24806,N_22599,N_22959);
xor U24807 (N_24807,N_23008,N_21721);
xnor U24808 (N_24808,N_21245,N_21465);
nor U24809 (N_24809,N_23452,N_22419);
and U24810 (N_24810,N_22055,N_22767);
nor U24811 (N_24811,N_21695,N_22543);
nor U24812 (N_24812,N_21443,N_21321);
and U24813 (N_24813,N_21334,N_21693);
or U24814 (N_24814,N_21303,N_23503);
nand U24815 (N_24815,N_23804,N_23635);
nand U24816 (N_24816,N_21025,N_23208);
and U24817 (N_24817,N_23939,N_23247);
xnor U24818 (N_24818,N_23472,N_21374);
xnor U24819 (N_24819,N_23942,N_22811);
and U24820 (N_24820,N_23214,N_21049);
xor U24821 (N_24821,N_23996,N_22305);
nor U24822 (N_24822,N_22854,N_22413);
nand U24823 (N_24823,N_21205,N_21006);
or U24824 (N_24824,N_23974,N_21790);
nor U24825 (N_24825,N_22017,N_22804);
and U24826 (N_24826,N_21525,N_22605);
nand U24827 (N_24827,N_22878,N_21975);
nor U24828 (N_24828,N_22961,N_22031);
xor U24829 (N_24829,N_21484,N_21621);
and U24830 (N_24830,N_23320,N_22264);
xnor U24831 (N_24831,N_22861,N_21114);
or U24832 (N_24832,N_21224,N_22107);
or U24833 (N_24833,N_21903,N_22876);
and U24834 (N_24834,N_22267,N_22403);
nor U24835 (N_24835,N_22191,N_22679);
or U24836 (N_24836,N_21900,N_21032);
xor U24837 (N_24837,N_22144,N_22313);
nor U24838 (N_24838,N_23421,N_22956);
xnor U24839 (N_24839,N_21439,N_23552);
or U24840 (N_24840,N_21831,N_22625);
nand U24841 (N_24841,N_22965,N_21773);
nor U24842 (N_24842,N_22293,N_23066);
nor U24843 (N_24843,N_22477,N_22479);
xnor U24844 (N_24844,N_21492,N_23473);
nand U24845 (N_24845,N_21603,N_22046);
or U24846 (N_24846,N_22682,N_23367);
and U24847 (N_24847,N_21755,N_22976);
nand U24848 (N_24848,N_23458,N_22163);
nand U24849 (N_24849,N_21571,N_22735);
xnor U24850 (N_24850,N_22497,N_21500);
and U24851 (N_24851,N_22198,N_22856);
xor U24852 (N_24852,N_22309,N_23045);
nand U24853 (N_24853,N_21718,N_22051);
nor U24854 (N_24854,N_23604,N_23130);
xnor U24855 (N_24855,N_22091,N_23966);
and U24856 (N_24856,N_21512,N_22040);
nand U24857 (N_24857,N_21135,N_22180);
and U24858 (N_24858,N_22338,N_21172);
xor U24859 (N_24859,N_22814,N_21085);
xor U24860 (N_24860,N_21766,N_21304);
or U24861 (N_24861,N_21354,N_23679);
or U24862 (N_24862,N_21476,N_23907);
xor U24863 (N_24863,N_23844,N_21488);
or U24864 (N_24864,N_21686,N_22664);
nor U24865 (N_24865,N_23229,N_21888);
xor U24866 (N_24866,N_23570,N_21376);
and U24867 (N_24867,N_23565,N_23651);
and U24868 (N_24868,N_23785,N_22294);
xor U24869 (N_24869,N_23054,N_22561);
nor U24870 (N_24870,N_22028,N_22232);
nor U24871 (N_24871,N_23520,N_21598);
and U24872 (N_24872,N_21668,N_21343);
nor U24873 (N_24873,N_23052,N_23495);
or U24874 (N_24874,N_22270,N_23244);
xor U24875 (N_24875,N_22304,N_21124);
and U24876 (N_24876,N_21884,N_23876);
or U24877 (N_24877,N_22886,N_21869);
and U24878 (N_24878,N_21062,N_22780);
and U24879 (N_24879,N_21854,N_22621);
xnor U24880 (N_24880,N_22681,N_23993);
nand U24881 (N_24881,N_21399,N_22934);
or U24882 (N_24882,N_21867,N_23972);
nor U24883 (N_24883,N_21909,N_21801);
xnor U24884 (N_24884,N_21599,N_21847);
and U24885 (N_24885,N_21407,N_21956);
nor U24886 (N_24886,N_22126,N_22741);
nand U24887 (N_24887,N_21393,N_22779);
nor U24888 (N_24888,N_23137,N_21814);
xor U24889 (N_24889,N_22758,N_21404);
and U24890 (N_24890,N_23344,N_22859);
nand U24891 (N_24891,N_21627,N_22218);
nand U24892 (N_24892,N_21699,N_22848);
or U24893 (N_24893,N_23427,N_23248);
nor U24894 (N_24894,N_22809,N_22427);
xnor U24895 (N_24895,N_21052,N_23484);
nand U24896 (N_24896,N_21835,N_23070);
or U24897 (N_24897,N_21005,N_21147);
or U24898 (N_24898,N_21635,N_21838);
and U24899 (N_24899,N_23224,N_22416);
nor U24900 (N_24900,N_21681,N_22580);
xor U24901 (N_24901,N_21540,N_23957);
or U24902 (N_24902,N_23787,N_22154);
and U24903 (N_24903,N_21314,N_23671);
and U24904 (N_24904,N_22369,N_22549);
nand U24905 (N_24905,N_23451,N_22385);
nor U24906 (N_24906,N_21702,N_23029);
xor U24907 (N_24907,N_23268,N_21262);
and U24908 (N_24908,N_21504,N_22515);
or U24909 (N_24909,N_21752,N_23168);
xor U24910 (N_24910,N_23752,N_23167);
nand U24911 (N_24911,N_23638,N_22909);
and U24912 (N_24912,N_21513,N_22324);
xnor U24913 (N_24913,N_23537,N_23185);
xnor U24914 (N_24914,N_21454,N_21988);
xnor U24915 (N_24915,N_23234,N_21519);
xnor U24916 (N_24916,N_21757,N_22850);
and U24917 (N_24917,N_23071,N_21138);
or U24918 (N_24918,N_22612,N_22426);
nor U24919 (N_24919,N_23235,N_22371);
xnor U24920 (N_24920,N_23771,N_22932);
nand U24921 (N_24921,N_21286,N_22491);
xnor U24922 (N_24922,N_21204,N_23015);
nor U24923 (N_24923,N_23843,N_22132);
nand U24924 (N_24924,N_23726,N_22451);
nor U24925 (N_24925,N_21786,N_23380);
nor U24926 (N_24926,N_22240,N_21921);
xor U24927 (N_24927,N_21732,N_22930);
nand U24928 (N_24928,N_23256,N_22175);
xor U24929 (N_24929,N_21582,N_22015);
nor U24930 (N_24930,N_22853,N_21126);
and U24931 (N_24931,N_23591,N_22315);
or U24932 (N_24932,N_21336,N_23935);
nor U24933 (N_24933,N_23792,N_23142);
or U24934 (N_24934,N_23762,N_22174);
xnor U24935 (N_24935,N_22788,N_22880);
xor U24936 (N_24936,N_21770,N_23444);
nor U24937 (N_24937,N_22537,N_21366);
nor U24938 (N_24938,N_23023,N_23913);
xnor U24939 (N_24939,N_21659,N_23796);
and U24940 (N_24940,N_22585,N_22475);
xnor U24941 (N_24941,N_22002,N_21459);
xnor U24942 (N_24942,N_22805,N_22935);
nor U24943 (N_24943,N_23644,N_22079);
nor U24944 (N_24944,N_22239,N_23441);
and U24945 (N_24945,N_22713,N_23037);
nor U24946 (N_24946,N_21984,N_21035);
or U24947 (N_24947,N_23336,N_21803);
xor U24948 (N_24948,N_23832,N_21173);
and U24949 (N_24949,N_23143,N_21541);
and U24950 (N_24950,N_23356,N_21671);
xnor U24951 (N_24951,N_23195,N_22097);
nand U24952 (N_24952,N_21373,N_23905);
nor U24953 (N_24953,N_23160,N_21193);
nor U24954 (N_24954,N_23310,N_22437);
xnor U24955 (N_24955,N_21735,N_21726);
nor U24956 (N_24956,N_23040,N_23482);
xor U24957 (N_24957,N_21238,N_23404);
xnor U24958 (N_24958,N_22089,N_23716);
and U24959 (N_24959,N_21624,N_23585);
and U24960 (N_24960,N_22242,N_23622);
nor U24961 (N_24961,N_21108,N_23860);
and U24962 (N_24962,N_21698,N_22940);
and U24963 (N_24963,N_22464,N_22597);
nor U24964 (N_24964,N_23936,N_23445);
nand U24965 (N_24965,N_23971,N_22098);
nand U24966 (N_24966,N_23999,N_21916);
xnor U24967 (N_24967,N_23711,N_23109);
nor U24968 (N_24968,N_22624,N_23148);
nor U24969 (N_24969,N_22734,N_22496);
nor U24970 (N_24970,N_21105,N_21815);
nand U24971 (N_24971,N_22183,N_23521);
and U24972 (N_24972,N_23217,N_23557);
nand U24973 (N_24973,N_22009,N_22776);
nand U24974 (N_24974,N_22787,N_21469);
or U24975 (N_24975,N_21860,N_22234);
or U24976 (N_24976,N_22130,N_22194);
or U24977 (N_24977,N_21093,N_23944);
xor U24978 (N_24978,N_22982,N_23241);
xor U24979 (N_24979,N_23581,N_21168);
xor U24980 (N_24980,N_21769,N_22262);
nor U24981 (N_24981,N_23781,N_23839);
nor U24982 (N_24982,N_22640,N_22550);
nor U24983 (N_24983,N_22552,N_23930);
nand U24984 (N_24984,N_22149,N_21947);
nand U24985 (N_24985,N_21954,N_22241);
and U24986 (N_24986,N_23303,N_21969);
xnor U24987 (N_24987,N_21837,N_22249);
nand U24988 (N_24988,N_23745,N_21538);
and U24989 (N_24989,N_22235,N_21549);
xnor U24990 (N_24990,N_21480,N_22526);
and U24991 (N_24991,N_22831,N_23714);
xnor U24992 (N_24992,N_23634,N_22129);
or U24993 (N_24993,N_21807,N_22373);
or U24994 (N_24994,N_22252,N_21084);
nand U24995 (N_24995,N_23001,N_21142);
nor U24996 (N_24996,N_21187,N_23363);
xor U24997 (N_24997,N_23946,N_21799);
xnor U24998 (N_24998,N_21435,N_22579);
and U24999 (N_24999,N_21796,N_21537);
or U25000 (N_25000,N_21970,N_22268);
nand U25001 (N_25001,N_23766,N_21751);
nand U25002 (N_25002,N_22656,N_22993);
or U25003 (N_25003,N_23097,N_22950);
or U25004 (N_25004,N_21051,N_22275);
xor U25005 (N_25005,N_21904,N_22364);
nand U25006 (N_25006,N_23740,N_22676);
nand U25007 (N_25007,N_23301,N_21701);
nand U25008 (N_25008,N_23559,N_21401);
and U25009 (N_25009,N_23818,N_23182);
and U25010 (N_25010,N_21398,N_21745);
and U25011 (N_25011,N_22135,N_21106);
nor U25012 (N_25012,N_21218,N_23509);
xor U25013 (N_25013,N_23435,N_21057);
xnor U25014 (N_25014,N_22435,N_22072);
or U25015 (N_25015,N_23709,N_23719);
xor U25016 (N_25016,N_21705,N_22308);
and U25017 (N_25017,N_21505,N_22958);
or U25018 (N_25018,N_22977,N_21749);
nand U25019 (N_25019,N_21394,N_23355);
nor U25020 (N_25020,N_22567,N_21972);
nand U25021 (N_25021,N_23650,N_22131);
or U25022 (N_25022,N_23076,N_22438);
or U25023 (N_25023,N_23992,N_21623);
nand U25024 (N_25024,N_23743,N_23313);
and U25025 (N_25025,N_21284,N_22637);
nand U25026 (N_25026,N_23108,N_21099);
xnor U25027 (N_25027,N_22695,N_21045);
xor U25028 (N_25028,N_21288,N_22642);
and U25029 (N_25029,N_23854,N_21945);
xor U25030 (N_25030,N_21197,N_21153);
nor U25031 (N_25031,N_21919,N_22104);
nor U25032 (N_25032,N_23967,N_23660);
xnor U25033 (N_25033,N_22762,N_23947);
or U25034 (N_25034,N_21383,N_22660);
nand U25035 (N_25035,N_21432,N_23062);
xor U25036 (N_25036,N_22670,N_23809);
or U25037 (N_25037,N_23000,N_22155);
and U25038 (N_25038,N_21478,N_23077);
or U25039 (N_25039,N_23254,N_22200);
or U25040 (N_25040,N_23245,N_22265);
nor U25041 (N_25041,N_22193,N_23955);
nor U25042 (N_25042,N_22810,N_23981);
nand U25043 (N_25043,N_23941,N_23024);
xor U25044 (N_25044,N_22059,N_21789);
or U25045 (N_25045,N_23190,N_21977);
nand U25046 (N_25046,N_21610,N_22397);
nand U25047 (N_25047,N_21279,N_23739);
nor U25048 (N_25048,N_22568,N_22672);
and U25049 (N_25049,N_23794,N_22102);
nor U25050 (N_25050,N_23409,N_23293);
nand U25051 (N_25051,N_23588,N_22204);
or U25052 (N_25052,N_23322,N_23414);
or U25053 (N_25053,N_21857,N_21053);
and U25054 (N_25054,N_22006,N_21660);
or U25055 (N_25055,N_23098,N_23180);
or U25056 (N_25056,N_22841,N_21895);
or U25057 (N_25057,N_22133,N_23536);
nor U25058 (N_25058,N_21999,N_22007);
or U25059 (N_25059,N_23312,N_23006);
or U25060 (N_25060,N_22823,N_21750);
nand U25061 (N_25061,N_21502,N_22185);
or U25062 (N_25062,N_22048,N_21568);
and U25063 (N_25063,N_22732,N_22219);
and U25064 (N_25064,N_21034,N_23487);
nor U25065 (N_25065,N_23369,N_23979);
nand U25066 (N_25066,N_22802,N_23948);
and U25067 (N_25067,N_21414,N_21503);
and U25068 (N_25068,N_23133,N_21317);
or U25069 (N_25069,N_23381,N_22502);
or U25070 (N_25070,N_23030,N_22651);
nand U25071 (N_25071,N_22916,N_22937);
or U25072 (N_25072,N_21481,N_23963);
nand U25073 (N_25073,N_22514,N_21278);
nand U25074 (N_25074,N_21856,N_21534);
or U25075 (N_25075,N_23439,N_21601);
nor U25076 (N_25076,N_21226,N_21181);
or U25077 (N_25077,N_23172,N_22244);
or U25078 (N_25078,N_21233,N_22551);
and U25079 (N_25079,N_22591,N_23158);
nor U25080 (N_25080,N_23370,N_22432);
xnor U25081 (N_25081,N_23820,N_22387);
nand U25082 (N_25082,N_23004,N_23157);
nor U25083 (N_25083,N_23590,N_23687);
or U25084 (N_25084,N_21010,N_22465);
and U25085 (N_25085,N_21307,N_21098);
and U25086 (N_25086,N_23288,N_21774);
nor U25087 (N_25087,N_21597,N_22647);
nor U25088 (N_25088,N_22765,N_22507);
or U25089 (N_25089,N_23115,N_23753);
nand U25090 (N_25090,N_22205,N_21863);
xnor U25091 (N_25091,N_23721,N_21851);
nand U25092 (N_25092,N_22057,N_21678);
nand U25093 (N_25093,N_22849,N_23184);
xor U25094 (N_25094,N_23943,N_23118);
nand U25095 (N_25095,N_21486,N_23849);
nor U25096 (N_25096,N_21896,N_23664);
or U25097 (N_25097,N_22783,N_23259);
or U25098 (N_25098,N_21764,N_23243);
nor U25099 (N_25099,N_23686,N_21319);
nor U25100 (N_25100,N_21951,N_22867);
nand U25101 (N_25101,N_21580,N_22103);
and U25102 (N_25102,N_22049,N_22168);
nand U25103 (N_25103,N_23294,N_22146);
xor U25104 (N_25104,N_23566,N_22875);
or U25105 (N_25105,N_21315,N_21148);
nand U25106 (N_25106,N_23153,N_23958);
nand U25107 (N_25107,N_23817,N_23669);
xor U25108 (N_25108,N_22547,N_22742);
nor U25109 (N_25109,N_23647,N_23751);
nor U25110 (N_25110,N_21518,N_21950);
or U25111 (N_25111,N_23909,N_23450);
or U25112 (N_25112,N_22866,N_22022);
nand U25113 (N_25113,N_23748,N_21071);
nor U25114 (N_25114,N_23896,N_22774);
nor U25115 (N_25115,N_22066,N_22434);
xor U25116 (N_25116,N_23400,N_21940);
nand U25117 (N_25117,N_22151,N_21428);
nand U25118 (N_25118,N_21462,N_22225);
or U25119 (N_25119,N_21980,N_23390);
and U25120 (N_25120,N_22073,N_22838);
nand U25121 (N_25121,N_21235,N_22409);
nor U25122 (N_25122,N_22069,N_21018);
nor U25123 (N_25123,N_23058,N_22777);
nor U25124 (N_25124,N_21882,N_21805);
nand U25125 (N_25125,N_23025,N_23997);
nor U25126 (N_25126,N_22892,N_22312);
nor U25127 (N_25127,N_21330,N_21139);
and U25128 (N_25128,N_21730,N_22968);
or U25129 (N_25129,N_21517,N_22004);
xor U25130 (N_25130,N_21165,N_23334);
and U25131 (N_25131,N_23283,N_22824);
and U25132 (N_25132,N_22064,N_21783);
and U25133 (N_25133,N_23329,N_23095);
and U25134 (N_25134,N_23183,N_23494);
nand U25135 (N_25135,N_22899,N_22290);
xnor U25136 (N_25136,N_22229,N_23230);
or U25137 (N_25137,N_21202,N_23063);
nor U25138 (N_25138,N_21161,N_21116);
and U25139 (N_25139,N_22987,N_21167);
xnor U25140 (N_25140,N_21510,N_23908);
and U25141 (N_25141,N_22897,N_22872);
nand U25142 (N_25142,N_23806,N_23055);
and U25143 (N_25143,N_23682,N_21039);
xor U25144 (N_25144,N_23069,N_22480);
nand U25145 (N_25145,N_21536,N_23161);
and U25146 (N_25146,N_23530,N_23561);
or U25147 (N_25147,N_22948,N_22042);
xnor U25148 (N_25148,N_22960,N_23410);
nor U25149 (N_25149,N_23019,N_22678);
and U25150 (N_25150,N_23117,N_22359);
nand U25151 (N_25151,N_22299,N_22221);
xnor U25152 (N_25152,N_21893,N_21696);
nor U25153 (N_25153,N_22094,N_22209);
and U25154 (N_25154,N_23867,N_22443);
nor U25155 (N_25155,N_23695,N_22377);
or U25156 (N_25156,N_23345,N_21120);
xnor U25157 (N_25157,N_22436,N_22542);
and U25158 (N_25158,N_23080,N_23287);
nand U25159 (N_25159,N_22999,N_22770);
xnor U25160 (N_25160,N_21554,N_22441);
or U25161 (N_25161,N_21546,N_21633);
nor U25162 (N_25162,N_22349,N_21673);
or U25163 (N_25163,N_21825,N_23778);
xor U25164 (N_25164,N_22115,N_22384);
or U25165 (N_25165,N_21434,N_21506);
nor U25166 (N_25166,N_23149,N_23596);
and U25167 (N_25167,N_23710,N_22291);
nor U25168 (N_25168,N_22691,N_23032);
nand U25169 (N_25169,N_23744,N_22353);
and U25170 (N_25170,N_23618,N_21065);
nor U25171 (N_25171,N_22418,N_22206);
nand U25172 (N_25172,N_22901,N_22099);
and U25173 (N_25173,N_23550,N_21630);
nor U25174 (N_25174,N_23253,N_21797);
and U25175 (N_25175,N_21228,N_21912);
or U25176 (N_25176,N_23701,N_21335);
nor U25177 (N_25177,N_21077,N_23540);
nor U25178 (N_25178,N_21208,N_21604);
nor U25179 (N_25179,N_22510,N_22331);
nand U25180 (N_25180,N_22389,N_21364);
or U25181 (N_25181,N_23331,N_22898);
or U25182 (N_25182,N_21328,N_21140);
and U25183 (N_25183,N_21526,N_23932);
nor U25184 (N_25184,N_23606,N_22078);
or U25185 (N_25185,N_22781,N_23674);
or U25186 (N_25186,N_23387,N_21356);
xor U25187 (N_25187,N_23384,N_21232);
and U25188 (N_25188,N_21007,N_21136);
or U25189 (N_25189,N_23707,N_22118);
xor U25190 (N_25190,N_22798,N_23933);
and U25191 (N_25191,N_22251,N_23879);
and U25192 (N_25192,N_22399,N_21019);
xnor U25193 (N_25193,N_23636,N_21949);
nor U25194 (N_25194,N_21653,N_23770);
nor U25195 (N_25195,N_21927,N_21371);
or U25196 (N_25196,N_22620,N_23124);
nor U25197 (N_25197,N_22667,N_23393);
xnor U25198 (N_25198,N_23209,N_22826);
and U25199 (N_25199,N_21906,N_23911);
or U25200 (N_25200,N_23545,N_23091);
xnor U25201 (N_25201,N_21133,N_23977);
and U25202 (N_25202,N_21413,N_21067);
nand U25203 (N_25203,N_22796,N_23965);
xnor U25204 (N_25204,N_22259,N_22466);
xor U25205 (N_25205,N_23512,N_23249);
and U25206 (N_25206,N_21542,N_21209);
xor U25207 (N_25207,N_21001,N_21556);
and U25208 (N_25208,N_22795,N_21914);
or U25209 (N_25209,N_22282,N_23546);
and U25210 (N_25210,N_22483,N_22068);
xnor U25211 (N_25211,N_21163,N_23431);
nor U25212 (N_25212,N_23858,N_23084);
nand U25213 (N_25213,N_22446,N_21995);
nand U25214 (N_25214,N_22792,N_21044);
xor U25215 (N_25215,N_21422,N_22827);
and U25216 (N_25216,N_22692,N_23640);
nand U25217 (N_25217,N_23034,N_22143);
nor U25218 (N_25218,N_23575,N_23735);
nor U25219 (N_25219,N_23093,N_22023);
xnor U25220 (N_25220,N_22544,N_21145);
nor U25221 (N_25221,N_23127,N_22855);
nand U25222 (N_25222,N_22116,N_23758);
or U25223 (N_25223,N_23488,N_23987);
nor U25224 (N_25224,N_22178,N_23073);
nand U25225 (N_25225,N_22908,N_23777);
xor U25226 (N_25226,N_22375,N_22688);
and U25227 (N_25227,N_21281,N_21917);
xor U25228 (N_25228,N_23677,N_22269);
xnor U25229 (N_25229,N_23442,N_22428);
or U25230 (N_25230,N_21078,N_21298);
nand U25231 (N_25231,N_21171,N_21267);
nor U25232 (N_25232,N_22490,N_22978);
and U25233 (N_25233,N_23853,N_23549);
or U25234 (N_25234,N_21000,N_22714);
nand U25235 (N_25235,N_21611,N_22588);
or U25236 (N_25236,N_23920,N_22246);
nor U25237 (N_25237,N_22535,N_21689);
nand U25238 (N_25238,N_22828,N_21775);
xor U25239 (N_25239,N_23586,N_21573);
nand U25240 (N_25240,N_23889,N_22356);
nor U25241 (N_25241,N_21121,N_23534);
nor U25242 (N_25242,N_22593,N_23104);
xor U25243 (N_25243,N_22724,N_22196);
nand U25244 (N_25244,N_21340,N_21472);
xor U25245 (N_25245,N_22595,N_23176);
nor U25246 (N_25246,N_21473,N_22147);
nor U25247 (N_25247,N_21804,N_23773);
or U25248 (N_25248,N_21253,N_21820);
or U25249 (N_25249,N_21527,N_22562);
xnor U25250 (N_25250,N_22980,N_23490);
or U25251 (N_25251,N_23138,N_23323);
nand U25252 (N_25252,N_22730,N_21690);
or U25253 (N_25253,N_22808,N_23798);
xor U25254 (N_25254,N_22020,N_22063);
xnor U25255 (N_25255,N_21887,N_23827);
nor U25256 (N_25256,N_22217,N_23022);
xnor U25257 (N_25257,N_23460,N_21036);
xnor U25258 (N_25258,N_23469,N_21442);
nor U25259 (N_25259,N_23360,N_23756);
or U25260 (N_25260,N_22386,N_22610);
and U25261 (N_25261,N_23102,N_22320);
xnor U25262 (N_25262,N_21551,N_23554);
xnor U25263 (N_25263,N_21881,N_22381);
nand U25264 (N_25264,N_22277,N_22590);
or U25265 (N_25265,N_22224,N_22280);
nor U25266 (N_25266,N_23599,N_23542);
nor U25267 (N_25267,N_23513,N_21349);
nor U25268 (N_25268,N_22799,N_22981);
xor U25269 (N_25269,N_23755,N_23951);
xnor U25270 (N_25270,N_23085,N_23377);
or U25271 (N_25271,N_21491,N_21274);
xnor U25272 (N_25272,N_22470,N_23275);
xnor U25273 (N_25273,N_22314,N_22768);
xor U25274 (N_25274,N_21320,N_22609);
and U25275 (N_25275,N_22818,N_23236);
and U25276 (N_25276,N_23122,N_21938);
or U25277 (N_25277,N_21131,N_22801);
and U25278 (N_25278,N_21339,N_23616);
xor U25279 (N_25279,N_23221,N_22966);
nand U25280 (N_25280,N_21572,N_22952);
nor U25281 (N_25281,N_21645,N_23982);
nor U25282 (N_25282,N_22472,N_23600);
and U25283 (N_25283,N_22986,N_21795);
nor U25284 (N_25284,N_23110,N_21331);
nor U25285 (N_25285,N_23276,N_23990);
nor U25286 (N_25286,N_22931,N_22865);
nand U25287 (N_25287,N_22412,N_21013);
nor U25288 (N_25288,N_23995,N_21048);
nor U25289 (N_25289,N_23754,N_22453);
nor U25290 (N_25290,N_23307,N_22584);
nor U25291 (N_25291,N_21868,N_21316);
nand U25292 (N_25292,N_21372,N_22273);
xor U25293 (N_25293,N_21979,N_22058);
or U25294 (N_25294,N_22785,N_21644);
nor U25295 (N_25295,N_21615,N_23002);
nand U25296 (N_25296,N_21113,N_21719);
nor U25297 (N_25297,N_21137,N_21166);
nor U25298 (N_25298,N_21935,N_21192);
xnor U25299 (N_25299,N_22704,N_22462);
and U25300 (N_25300,N_23162,N_21375);
xor U25301 (N_25301,N_22030,N_23413);
and U25302 (N_25302,N_23189,N_21152);
or U25303 (N_25303,N_22093,N_22984);
and U25304 (N_25304,N_22719,N_23801);
nand U25305 (N_25305,N_23661,N_21811);
or U25306 (N_25306,N_22220,N_23232);
nor U25307 (N_25307,N_23776,N_21352);
or U25308 (N_25308,N_23251,N_23870);
nor U25309 (N_25309,N_22307,N_22910);
xnor U25310 (N_25310,N_21100,N_22141);
or U25311 (N_25311,N_22407,N_21174);
nor U25312 (N_25312,N_21741,N_23021);
nor U25313 (N_25313,N_21605,N_23852);
xor U25314 (N_25314,N_22646,N_21553);
or U25315 (N_25315,N_21306,N_23416);
or U25316 (N_25316,N_21885,N_21872);
or U25317 (N_25317,N_23514,N_21606);
nand U25318 (N_25318,N_22879,N_23774);
nor U25319 (N_25319,N_23499,N_21474);
xnor U25320 (N_25320,N_23281,N_22650);
nor U25321 (N_25321,N_23100,N_23493);
or U25322 (N_25322,N_21771,N_21759);
nand U25323 (N_25323,N_22836,N_22571);
or U25324 (N_25324,N_21669,N_23314);
nand U25325 (N_25325,N_23702,N_21162);
xor U25326 (N_25326,N_21688,N_22725);
and U25327 (N_25327,N_22351,N_23155);
xnor U25328 (N_25328,N_22362,N_23956);
xor U25329 (N_25329,N_23337,N_21295);
xor U25330 (N_25330,N_22603,N_22873);
xnor U25331 (N_25331,N_23078,N_23299);
and U25332 (N_25332,N_21994,N_22370);
nor U25333 (N_25333,N_23961,N_23169);
or U25334 (N_25334,N_21986,N_22985);
nand U25335 (N_25335,N_22257,N_21026);
nor U25336 (N_25336,N_22608,N_21613);
xor U25337 (N_25337,N_23805,N_23688);
xor U25338 (N_25338,N_21692,N_22458);
nand U25339 (N_25339,N_23985,N_21282);
nand U25340 (N_25340,N_22256,N_21760);
xor U25341 (N_25341,N_21974,N_21191);
and U25342 (N_25342,N_23213,N_23031);
and U25343 (N_25343,N_22365,N_22863);
or U25344 (N_25344,N_22534,N_22914);
nor U25345 (N_25345,N_22598,N_22920);
and U25346 (N_25346,N_22752,N_23483);
xor U25347 (N_25347,N_23926,N_21879);
xor U25348 (N_25348,N_23612,N_23014);
nand U25349 (N_25349,N_23028,N_22442);
nor U25350 (N_25350,N_22616,N_22771);
nor U25351 (N_25351,N_22335,N_23814);
nand U25352 (N_25352,N_21342,N_21421);
nand U25353 (N_25353,N_22105,N_22159);
xor U25354 (N_25354,N_23395,N_21649);
or U25355 (N_25355,N_21022,N_23170);
or U25356 (N_25356,N_21650,N_22740);
xnor U25357 (N_25357,N_21547,N_23394);
or U25358 (N_25358,N_21016,N_22998);
or U25359 (N_25359,N_23525,N_23724);
xnor U25360 (N_25360,N_21129,N_22321);
nand U25361 (N_25361,N_21602,N_22671);
or U25362 (N_25362,N_22530,N_23353);
nand U25363 (N_25363,N_21933,N_23405);
nor U25364 (N_25364,N_21095,N_22548);
or U25365 (N_25365,N_21691,N_23799);
xnor U25366 (N_25366,N_22188,N_21866);
nand U25367 (N_25367,N_22053,N_22482);
or U25368 (N_25368,N_23223,N_23081);
nor U25369 (N_25369,N_22596,N_23815);
nor U25370 (N_25370,N_22202,N_21576);
or U25371 (N_25371,N_21158,N_21309);
nand U25372 (N_25372,N_21561,N_21607);
xor U25373 (N_25373,N_21575,N_21441);
nor U25374 (N_25374,N_23420,N_22208);
nand U25375 (N_25375,N_22279,N_21829);
nor U25376 (N_25376,N_23523,N_23595);
nand U25377 (N_25377,N_21387,N_21793);
and U25378 (N_25378,N_22238,N_23851);
nor U25379 (N_25379,N_23914,N_22806);
or U25380 (N_25380,N_23764,N_22245);
xor U25381 (N_25381,N_22008,N_21430);
nand U25382 (N_25382,N_22707,N_22392);
or U25383 (N_25383,N_22038,N_22248);
and U25384 (N_25384,N_23325,N_22519);
nor U25385 (N_25385,N_22223,N_22586);
xnor U25386 (N_25386,N_22789,N_22139);
nor U25387 (N_25387,N_21907,N_21585);
or U25388 (N_25388,N_22668,N_23594);
nor U25389 (N_25389,N_22499,N_22944);
or U25390 (N_25390,N_21782,N_23703);
nor U25391 (N_25391,N_23156,N_22037);
or U25392 (N_25392,N_21249,N_21809);
nor U25393 (N_25393,N_21612,N_23267);
xor U25394 (N_25394,N_23179,N_22211);
and U25395 (N_25395,N_23107,N_23733);
nor U25396 (N_25396,N_22036,N_21004);
nand U25397 (N_25397,N_21134,N_21269);
xor U25398 (N_25398,N_23196,N_23583);
xnor U25399 (N_25399,N_22468,N_22061);
xnor U25400 (N_25400,N_21780,N_23884);
nand U25401 (N_25401,N_23630,N_23903);
and U25402 (N_25402,N_22214,N_23825);
xnor U25403 (N_25403,N_23789,N_23718);
xor U25404 (N_25404,N_23681,N_22182);
xnor U25405 (N_25405,N_22953,N_23265);
and U25406 (N_25406,N_23150,N_22712);
and U25407 (N_25407,N_23376,N_21911);
nand U25408 (N_25408,N_22323,N_21530);
xor U25409 (N_25409,N_21359,N_21508);
nor U25410 (N_25410,N_23470,N_21981);
nand U25411 (N_25411,N_22717,N_22489);
and U25412 (N_25412,N_23315,N_22459);
nand U25413 (N_25413,N_23131,N_23722);
and U25414 (N_25414,N_23375,N_22336);
or U25415 (N_25415,N_21302,N_23291);
xnor U25416 (N_25416,N_22013,N_22157);
and U25417 (N_25417,N_23945,N_22524);
xnor U25418 (N_25418,N_22035,N_23610);
nand U25419 (N_25419,N_23715,N_23897);
nor U25420 (N_25420,N_22150,N_23471);
nand U25421 (N_25421,N_22076,N_22720);
nand U25422 (N_25422,N_23893,N_22189);
nor U25423 (N_25423,N_23140,N_23632);
xor U25424 (N_25424,N_22657,N_23609);
nand U25425 (N_25425,N_22918,N_22883);
nand U25426 (N_25426,N_21742,N_22871);
nor U25427 (N_25427,N_21647,N_22457);
or U25428 (N_25428,N_22644,N_23402);
xor U25429 (N_25429,N_22050,N_23597);
xnor U25430 (N_25430,N_21132,N_22645);
xnor U25431 (N_25431,N_22677,N_23498);
nor U25432 (N_25432,N_21146,N_22043);
xnor U25433 (N_25433,N_22623,N_23433);
nand U25434 (N_25434,N_21271,N_22611);
and U25435 (N_25435,N_23962,N_23476);
and U25436 (N_25436,N_21350,N_22617);
or U25437 (N_25437,N_21489,N_22374);
nand U25438 (N_25438,N_22511,N_22250);
xnor U25439 (N_25439,N_23822,N_21577);
nand U25440 (N_25440,N_22195,N_21565);
xnor U25441 (N_25441,N_22493,N_21276);
or U25442 (N_25442,N_21560,N_22870);
and U25443 (N_25443,N_23797,N_22685);
or U25444 (N_25444,N_21676,N_23317);
nand U25445 (N_25445,N_22463,N_21548);
and U25446 (N_25446,N_23885,N_23468);
or U25447 (N_25447,N_22619,N_21600);
and U25448 (N_25448,N_22271,N_23658);
nand U25449 (N_25449,N_21456,N_22698);
xnor U25450 (N_25450,N_23580,N_23324);
or U25451 (N_25451,N_21643,N_22896);
xor U25452 (N_25452,N_23734,N_22176);
nand U25453 (N_25453,N_23668,N_22153);
xnor U25454 (N_25454,N_21562,N_21086);
xor U25455 (N_25455,N_22333,N_21426);
nor U25456 (N_25456,N_23197,N_21003);
and U25457 (N_25457,N_23466,N_22393);
nand U25458 (N_25458,N_22833,N_23181);
nand U25459 (N_25459,N_22255,N_23467);
xor U25460 (N_25460,N_23290,N_23340);
or U25461 (N_25461,N_23273,N_21993);
nand U25462 (N_25462,N_22746,N_21674);
xor U25463 (N_25463,N_21664,N_23831);
nor U25464 (N_25464,N_23543,N_21656);
nor U25465 (N_25465,N_21379,N_23096);
nand U25466 (N_25466,N_21840,N_21103);
nor U25467 (N_25467,N_21843,N_23890);
nand U25468 (N_25468,N_23088,N_22311);
nor U25469 (N_25469,N_23270,N_23614);
nand U25470 (N_25470,N_22531,N_21559);
xor U25471 (N_25471,N_22111,N_22639);
nor U25472 (N_25472,N_22991,N_23406);
xor U25473 (N_25473,N_23422,N_21255);
and U25474 (N_25474,N_22721,N_21727);
xor U25475 (N_25475,N_23059,N_21846);
xnor U25476 (N_25476,N_23819,N_21467);
and U25477 (N_25477,N_21125,N_22062);
nor U25478 (N_25478,N_23398,N_21667);
or U25479 (N_25479,N_21324,N_23361);
xor U25480 (N_25480,N_22227,N_22906);
and U25481 (N_25481,N_22594,N_22754);
and U25482 (N_25482,N_23919,N_23871);
nor U25483 (N_25483,N_21864,N_23492);
nor U25484 (N_25484,N_23448,N_22835);
xnor U25485 (N_25485,N_21070,N_21326);
xor U25486 (N_25486,N_21593,N_21028);
nand U25487 (N_25487,N_23868,N_21514);
nand U25488 (N_25488,N_22166,N_23056);
xor U25489 (N_25489,N_23216,N_22708);
xnor U25490 (N_25490,N_21952,N_21963);
or U25491 (N_25491,N_23928,N_21654);
nand U25492 (N_25492,N_23670,N_23412);
nand U25493 (N_25493,N_23178,N_23106);
xor U25494 (N_25494,N_22422,N_21179);
or U25495 (N_25495,N_22081,N_21876);
or U25496 (N_25496,N_21074,N_22120);
nor U25497 (N_25497,N_22345,N_23211);
nor U25498 (N_25498,N_22405,N_21157);
and U25499 (N_25499,N_21976,N_23225);
and U25500 (N_25500,N_23779,N_22135);
xnor U25501 (N_25501,N_21457,N_23557);
and U25502 (N_25502,N_21656,N_21533);
or U25503 (N_25503,N_22135,N_21579);
xor U25504 (N_25504,N_21936,N_23654);
and U25505 (N_25505,N_21086,N_22624);
nor U25506 (N_25506,N_23738,N_22903);
or U25507 (N_25507,N_22758,N_22227);
or U25508 (N_25508,N_23891,N_21460);
and U25509 (N_25509,N_22422,N_21515);
xor U25510 (N_25510,N_23302,N_23752);
nor U25511 (N_25511,N_22330,N_23713);
or U25512 (N_25512,N_23499,N_21929);
xnor U25513 (N_25513,N_22684,N_22117);
nor U25514 (N_25514,N_22432,N_23689);
or U25515 (N_25515,N_22018,N_21672);
nand U25516 (N_25516,N_22643,N_21692);
or U25517 (N_25517,N_22755,N_22387);
or U25518 (N_25518,N_22162,N_23310);
xor U25519 (N_25519,N_23529,N_22281);
nor U25520 (N_25520,N_21525,N_21576);
and U25521 (N_25521,N_22271,N_21688);
xor U25522 (N_25522,N_21538,N_21399);
and U25523 (N_25523,N_22222,N_22133);
and U25524 (N_25524,N_21126,N_23542);
and U25525 (N_25525,N_22567,N_22302);
nand U25526 (N_25526,N_21430,N_21568);
xnor U25527 (N_25527,N_23278,N_21460);
xnor U25528 (N_25528,N_21382,N_21172);
xor U25529 (N_25529,N_23692,N_21620);
nor U25530 (N_25530,N_21871,N_21677);
nand U25531 (N_25531,N_23851,N_23545);
nor U25532 (N_25532,N_21625,N_21056);
nand U25533 (N_25533,N_23043,N_21340);
xnor U25534 (N_25534,N_21890,N_21784);
nand U25535 (N_25535,N_23309,N_23313);
nand U25536 (N_25536,N_22300,N_23301);
nand U25537 (N_25537,N_23603,N_21126);
nand U25538 (N_25538,N_22703,N_22052);
nand U25539 (N_25539,N_22039,N_23134);
and U25540 (N_25540,N_22668,N_21332);
nor U25541 (N_25541,N_22677,N_21065);
nand U25542 (N_25542,N_23746,N_22746);
xnor U25543 (N_25543,N_21757,N_21001);
nor U25544 (N_25544,N_23911,N_22441);
nand U25545 (N_25545,N_22293,N_22111);
nand U25546 (N_25546,N_21844,N_21424);
xor U25547 (N_25547,N_21098,N_21429);
xnor U25548 (N_25548,N_22056,N_23974);
nor U25549 (N_25549,N_21864,N_23896);
nor U25550 (N_25550,N_21071,N_21674);
or U25551 (N_25551,N_22507,N_23831);
nor U25552 (N_25552,N_21179,N_21092);
xor U25553 (N_25553,N_23722,N_23453);
nand U25554 (N_25554,N_21685,N_21875);
and U25555 (N_25555,N_23973,N_23627);
nand U25556 (N_25556,N_22613,N_21817);
and U25557 (N_25557,N_22610,N_21178);
nor U25558 (N_25558,N_23110,N_22559);
xnor U25559 (N_25559,N_21013,N_23518);
nor U25560 (N_25560,N_21171,N_23899);
or U25561 (N_25561,N_22834,N_23219);
or U25562 (N_25562,N_23795,N_23299);
nor U25563 (N_25563,N_21489,N_21240);
xnor U25564 (N_25564,N_21142,N_22782);
nor U25565 (N_25565,N_22408,N_23371);
nand U25566 (N_25566,N_21017,N_23625);
nor U25567 (N_25567,N_21967,N_22723);
and U25568 (N_25568,N_23789,N_23823);
and U25569 (N_25569,N_23725,N_21765);
and U25570 (N_25570,N_22013,N_23839);
and U25571 (N_25571,N_23405,N_23768);
nor U25572 (N_25572,N_23776,N_21824);
nor U25573 (N_25573,N_23074,N_23258);
or U25574 (N_25574,N_21137,N_23220);
and U25575 (N_25575,N_21573,N_23308);
nor U25576 (N_25576,N_23297,N_22705);
nor U25577 (N_25577,N_23366,N_22115);
nand U25578 (N_25578,N_23065,N_21414);
nand U25579 (N_25579,N_23659,N_23417);
or U25580 (N_25580,N_23526,N_23596);
nand U25581 (N_25581,N_21559,N_22749);
nor U25582 (N_25582,N_23435,N_22651);
nand U25583 (N_25583,N_22347,N_22773);
or U25584 (N_25584,N_21713,N_23562);
xor U25585 (N_25585,N_23851,N_21590);
xor U25586 (N_25586,N_21245,N_22375);
and U25587 (N_25587,N_23903,N_22407);
nand U25588 (N_25588,N_22796,N_23679);
nand U25589 (N_25589,N_21142,N_21576);
or U25590 (N_25590,N_21786,N_22711);
or U25591 (N_25591,N_21569,N_21556);
and U25592 (N_25592,N_22689,N_23379);
nand U25593 (N_25593,N_21129,N_21477);
or U25594 (N_25594,N_23628,N_21832);
nor U25595 (N_25595,N_23965,N_22947);
or U25596 (N_25596,N_22933,N_22368);
and U25597 (N_25597,N_23158,N_23389);
or U25598 (N_25598,N_21298,N_23943);
nand U25599 (N_25599,N_22815,N_22082);
or U25600 (N_25600,N_23191,N_22911);
and U25601 (N_25601,N_21955,N_23313);
and U25602 (N_25602,N_21408,N_23340);
and U25603 (N_25603,N_23439,N_22660);
nand U25604 (N_25604,N_22277,N_23035);
and U25605 (N_25605,N_22980,N_23877);
nand U25606 (N_25606,N_23153,N_22722);
xor U25607 (N_25607,N_23834,N_21581);
or U25608 (N_25608,N_23270,N_21256);
or U25609 (N_25609,N_21778,N_22527);
nand U25610 (N_25610,N_22162,N_21186);
nand U25611 (N_25611,N_21599,N_22497);
nand U25612 (N_25612,N_22935,N_21379);
or U25613 (N_25613,N_21364,N_23432);
xnor U25614 (N_25614,N_23962,N_23506);
nor U25615 (N_25615,N_22137,N_23467);
and U25616 (N_25616,N_21802,N_21092);
nor U25617 (N_25617,N_22295,N_22704);
or U25618 (N_25618,N_21500,N_22610);
nor U25619 (N_25619,N_22080,N_21217);
nor U25620 (N_25620,N_21663,N_21908);
xnor U25621 (N_25621,N_21132,N_22323);
nor U25622 (N_25622,N_21463,N_21519);
nor U25623 (N_25623,N_23806,N_21259);
or U25624 (N_25624,N_23426,N_23142);
or U25625 (N_25625,N_23321,N_23219);
nand U25626 (N_25626,N_23896,N_23111);
or U25627 (N_25627,N_23594,N_22298);
or U25628 (N_25628,N_21787,N_22915);
and U25629 (N_25629,N_21387,N_21796);
and U25630 (N_25630,N_21031,N_21158);
nor U25631 (N_25631,N_21246,N_22937);
xnor U25632 (N_25632,N_22965,N_22138);
xnor U25633 (N_25633,N_23025,N_22435);
or U25634 (N_25634,N_22579,N_22506);
or U25635 (N_25635,N_21407,N_23240);
or U25636 (N_25636,N_23202,N_22225);
xor U25637 (N_25637,N_21367,N_21671);
xnor U25638 (N_25638,N_22929,N_21766);
or U25639 (N_25639,N_21602,N_21400);
or U25640 (N_25640,N_23918,N_21355);
xor U25641 (N_25641,N_21602,N_23131);
xor U25642 (N_25642,N_23695,N_23389);
nor U25643 (N_25643,N_23980,N_22717);
xor U25644 (N_25644,N_21944,N_21945);
or U25645 (N_25645,N_23806,N_23667);
and U25646 (N_25646,N_22668,N_22284);
nand U25647 (N_25647,N_21012,N_22058);
nand U25648 (N_25648,N_22862,N_21396);
nand U25649 (N_25649,N_21389,N_21975);
xnor U25650 (N_25650,N_22821,N_21923);
nor U25651 (N_25651,N_22018,N_22721);
xor U25652 (N_25652,N_22904,N_22568);
xnor U25653 (N_25653,N_22812,N_23053);
xnor U25654 (N_25654,N_23191,N_22809);
xor U25655 (N_25655,N_22889,N_21203);
xnor U25656 (N_25656,N_23261,N_22949);
and U25657 (N_25657,N_21169,N_21765);
nor U25658 (N_25658,N_23091,N_21558);
nand U25659 (N_25659,N_21405,N_23128);
nor U25660 (N_25660,N_22580,N_23580);
nor U25661 (N_25661,N_22338,N_21433);
nand U25662 (N_25662,N_23338,N_23089);
xnor U25663 (N_25663,N_21933,N_23765);
nand U25664 (N_25664,N_21550,N_21018);
xnor U25665 (N_25665,N_21532,N_22613);
nand U25666 (N_25666,N_21278,N_23802);
xor U25667 (N_25667,N_22782,N_22558);
and U25668 (N_25668,N_23490,N_23243);
nor U25669 (N_25669,N_23100,N_21650);
or U25670 (N_25670,N_22961,N_22009);
nor U25671 (N_25671,N_23058,N_23145);
nand U25672 (N_25672,N_22872,N_21907);
or U25673 (N_25673,N_21252,N_23018);
or U25674 (N_25674,N_22511,N_22939);
nand U25675 (N_25675,N_23985,N_21625);
and U25676 (N_25676,N_22741,N_23734);
xnor U25677 (N_25677,N_21362,N_23695);
nand U25678 (N_25678,N_21671,N_23584);
or U25679 (N_25679,N_21826,N_22334);
and U25680 (N_25680,N_21857,N_22690);
nand U25681 (N_25681,N_21651,N_21104);
nor U25682 (N_25682,N_21973,N_22333);
and U25683 (N_25683,N_22989,N_21518);
nand U25684 (N_25684,N_21781,N_23562);
nand U25685 (N_25685,N_22519,N_22336);
or U25686 (N_25686,N_21688,N_23118);
and U25687 (N_25687,N_22808,N_22404);
xnor U25688 (N_25688,N_23538,N_22576);
and U25689 (N_25689,N_21105,N_21551);
and U25690 (N_25690,N_21078,N_22318);
nand U25691 (N_25691,N_22953,N_21473);
xnor U25692 (N_25692,N_21838,N_21231);
nor U25693 (N_25693,N_22893,N_23574);
nand U25694 (N_25694,N_21912,N_21370);
or U25695 (N_25695,N_21800,N_23579);
nand U25696 (N_25696,N_21348,N_21146);
or U25697 (N_25697,N_22334,N_21889);
and U25698 (N_25698,N_22758,N_21668);
and U25699 (N_25699,N_21382,N_22937);
or U25700 (N_25700,N_23758,N_22812);
or U25701 (N_25701,N_21903,N_22689);
and U25702 (N_25702,N_23087,N_22718);
nand U25703 (N_25703,N_21523,N_23204);
and U25704 (N_25704,N_21306,N_21504);
and U25705 (N_25705,N_23785,N_22577);
nor U25706 (N_25706,N_23488,N_21841);
nor U25707 (N_25707,N_21447,N_22048);
or U25708 (N_25708,N_23377,N_21868);
nand U25709 (N_25709,N_21978,N_23915);
nor U25710 (N_25710,N_23638,N_22231);
and U25711 (N_25711,N_22121,N_23332);
xnor U25712 (N_25712,N_21946,N_22685);
nor U25713 (N_25713,N_22638,N_22740);
xnor U25714 (N_25714,N_21913,N_21388);
nor U25715 (N_25715,N_23454,N_23183);
xor U25716 (N_25716,N_22543,N_23774);
or U25717 (N_25717,N_21123,N_21739);
nor U25718 (N_25718,N_23653,N_21538);
nor U25719 (N_25719,N_23471,N_23109);
xnor U25720 (N_25720,N_22326,N_23074);
nand U25721 (N_25721,N_22782,N_23738);
xnor U25722 (N_25722,N_23199,N_21602);
nor U25723 (N_25723,N_23289,N_21727);
xnor U25724 (N_25724,N_23769,N_22956);
xor U25725 (N_25725,N_21409,N_21026);
nor U25726 (N_25726,N_23229,N_23948);
and U25727 (N_25727,N_23882,N_21552);
and U25728 (N_25728,N_21010,N_23720);
xor U25729 (N_25729,N_22934,N_23824);
nor U25730 (N_25730,N_21553,N_21361);
nand U25731 (N_25731,N_22739,N_23655);
nor U25732 (N_25732,N_22768,N_22385);
and U25733 (N_25733,N_21817,N_23656);
xor U25734 (N_25734,N_22513,N_23325);
nand U25735 (N_25735,N_21119,N_23984);
nand U25736 (N_25736,N_22328,N_22583);
nand U25737 (N_25737,N_23837,N_23818);
nand U25738 (N_25738,N_23029,N_22664);
or U25739 (N_25739,N_23716,N_22164);
nand U25740 (N_25740,N_22850,N_22202);
or U25741 (N_25741,N_22992,N_22679);
nand U25742 (N_25742,N_23778,N_22684);
nor U25743 (N_25743,N_23905,N_23435);
and U25744 (N_25744,N_23852,N_23047);
or U25745 (N_25745,N_22580,N_22026);
or U25746 (N_25746,N_21965,N_23910);
and U25747 (N_25747,N_23146,N_22022);
nor U25748 (N_25748,N_22923,N_23210);
and U25749 (N_25749,N_21480,N_23459);
and U25750 (N_25750,N_23699,N_22866);
nand U25751 (N_25751,N_21729,N_21018);
nor U25752 (N_25752,N_23566,N_22826);
or U25753 (N_25753,N_21222,N_21394);
nor U25754 (N_25754,N_22233,N_21059);
nor U25755 (N_25755,N_21873,N_21376);
nor U25756 (N_25756,N_23099,N_21213);
and U25757 (N_25757,N_21865,N_22894);
nand U25758 (N_25758,N_21834,N_23394);
xnor U25759 (N_25759,N_22748,N_21471);
and U25760 (N_25760,N_21098,N_21285);
or U25761 (N_25761,N_21588,N_23611);
xnor U25762 (N_25762,N_21540,N_23946);
xor U25763 (N_25763,N_21461,N_22241);
or U25764 (N_25764,N_21027,N_23710);
nand U25765 (N_25765,N_23330,N_22274);
xnor U25766 (N_25766,N_22282,N_21547);
xnor U25767 (N_25767,N_22198,N_21783);
and U25768 (N_25768,N_23770,N_23483);
nand U25769 (N_25769,N_21006,N_22711);
xnor U25770 (N_25770,N_21582,N_23640);
and U25771 (N_25771,N_21025,N_22537);
nand U25772 (N_25772,N_21303,N_21539);
nand U25773 (N_25773,N_23671,N_23739);
nor U25774 (N_25774,N_21087,N_23474);
and U25775 (N_25775,N_23321,N_23951);
and U25776 (N_25776,N_22250,N_23206);
nor U25777 (N_25777,N_22477,N_23881);
or U25778 (N_25778,N_22558,N_21885);
nor U25779 (N_25779,N_22470,N_21242);
or U25780 (N_25780,N_21896,N_23432);
and U25781 (N_25781,N_23097,N_21643);
nand U25782 (N_25782,N_21138,N_23629);
and U25783 (N_25783,N_23480,N_23343);
nand U25784 (N_25784,N_22063,N_21367);
nor U25785 (N_25785,N_22436,N_23983);
nand U25786 (N_25786,N_22897,N_23237);
xnor U25787 (N_25787,N_21855,N_22768);
nand U25788 (N_25788,N_21496,N_23423);
xnor U25789 (N_25789,N_23933,N_21338);
nand U25790 (N_25790,N_23276,N_21220);
or U25791 (N_25791,N_23094,N_23601);
nand U25792 (N_25792,N_22831,N_21336);
nand U25793 (N_25793,N_22184,N_23610);
nor U25794 (N_25794,N_23511,N_22211);
xnor U25795 (N_25795,N_21312,N_21380);
or U25796 (N_25796,N_22163,N_23177);
and U25797 (N_25797,N_21129,N_21809);
nor U25798 (N_25798,N_23303,N_23600);
nor U25799 (N_25799,N_22028,N_21116);
nor U25800 (N_25800,N_21847,N_23215);
and U25801 (N_25801,N_22887,N_21869);
and U25802 (N_25802,N_22085,N_22420);
xnor U25803 (N_25803,N_22106,N_21970);
nor U25804 (N_25804,N_22299,N_22559);
nor U25805 (N_25805,N_22567,N_21957);
xnor U25806 (N_25806,N_21909,N_22635);
and U25807 (N_25807,N_21087,N_23637);
nor U25808 (N_25808,N_23928,N_22484);
and U25809 (N_25809,N_22768,N_22651);
nand U25810 (N_25810,N_22662,N_21460);
nand U25811 (N_25811,N_22664,N_22957);
or U25812 (N_25812,N_21749,N_21211);
or U25813 (N_25813,N_21888,N_22137);
or U25814 (N_25814,N_22061,N_22999);
nand U25815 (N_25815,N_22636,N_21381);
nor U25816 (N_25816,N_23984,N_23630);
or U25817 (N_25817,N_21366,N_22637);
nor U25818 (N_25818,N_22726,N_22930);
nand U25819 (N_25819,N_23078,N_22152);
and U25820 (N_25820,N_22744,N_22559);
or U25821 (N_25821,N_22546,N_22572);
nand U25822 (N_25822,N_22403,N_22985);
nand U25823 (N_25823,N_23659,N_22143);
xor U25824 (N_25824,N_22977,N_21471);
nand U25825 (N_25825,N_23502,N_22510);
nor U25826 (N_25826,N_21905,N_21060);
nand U25827 (N_25827,N_21262,N_23170);
and U25828 (N_25828,N_22980,N_23498);
nand U25829 (N_25829,N_22989,N_22209);
nor U25830 (N_25830,N_21812,N_23648);
nor U25831 (N_25831,N_22863,N_22209);
or U25832 (N_25832,N_22836,N_21725);
nand U25833 (N_25833,N_21583,N_22377);
or U25834 (N_25834,N_23510,N_22397);
nor U25835 (N_25835,N_23535,N_23200);
and U25836 (N_25836,N_22096,N_22142);
and U25837 (N_25837,N_23884,N_21049);
or U25838 (N_25838,N_22955,N_21537);
or U25839 (N_25839,N_22474,N_23746);
and U25840 (N_25840,N_21794,N_21313);
xor U25841 (N_25841,N_23884,N_22987);
or U25842 (N_25842,N_22878,N_23982);
nor U25843 (N_25843,N_21497,N_23091);
nor U25844 (N_25844,N_22755,N_21509);
nor U25845 (N_25845,N_22233,N_22161);
nor U25846 (N_25846,N_22592,N_23545);
nand U25847 (N_25847,N_21403,N_22569);
nand U25848 (N_25848,N_21240,N_22360);
xnor U25849 (N_25849,N_23031,N_22188);
nor U25850 (N_25850,N_21853,N_23339);
xnor U25851 (N_25851,N_22924,N_22108);
nor U25852 (N_25852,N_23109,N_23685);
xor U25853 (N_25853,N_21752,N_21258);
nor U25854 (N_25854,N_21730,N_23952);
nand U25855 (N_25855,N_21785,N_22602);
nor U25856 (N_25856,N_23221,N_22682);
and U25857 (N_25857,N_21284,N_21307);
nand U25858 (N_25858,N_22028,N_21523);
xor U25859 (N_25859,N_21075,N_21543);
nand U25860 (N_25860,N_23717,N_22025);
nor U25861 (N_25861,N_21885,N_23217);
or U25862 (N_25862,N_22837,N_22750);
nor U25863 (N_25863,N_21066,N_23367);
xnor U25864 (N_25864,N_22462,N_22686);
and U25865 (N_25865,N_23070,N_22417);
xnor U25866 (N_25866,N_21603,N_21308);
and U25867 (N_25867,N_22024,N_21494);
xnor U25868 (N_25868,N_23004,N_23884);
nor U25869 (N_25869,N_21090,N_23999);
xor U25870 (N_25870,N_23545,N_22591);
nor U25871 (N_25871,N_23314,N_21690);
and U25872 (N_25872,N_23336,N_23895);
or U25873 (N_25873,N_23568,N_23621);
nand U25874 (N_25874,N_21180,N_22428);
or U25875 (N_25875,N_21153,N_21857);
or U25876 (N_25876,N_23212,N_22933);
nor U25877 (N_25877,N_21192,N_22610);
xor U25878 (N_25878,N_21869,N_22740);
nand U25879 (N_25879,N_23964,N_21524);
nand U25880 (N_25880,N_23589,N_22601);
xor U25881 (N_25881,N_22064,N_23309);
nor U25882 (N_25882,N_22170,N_22184);
and U25883 (N_25883,N_21908,N_22625);
xor U25884 (N_25884,N_22718,N_21507);
nand U25885 (N_25885,N_23883,N_21846);
nand U25886 (N_25886,N_21141,N_22029);
and U25887 (N_25887,N_22696,N_22953);
nand U25888 (N_25888,N_21920,N_21147);
nand U25889 (N_25889,N_21666,N_22498);
or U25890 (N_25890,N_23815,N_23187);
or U25891 (N_25891,N_23242,N_23659);
and U25892 (N_25892,N_21764,N_23304);
nor U25893 (N_25893,N_21195,N_21043);
nand U25894 (N_25894,N_22040,N_21267);
and U25895 (N_25895,N_22658,N_23958);
xnor U25896 (N_25896,N_21778,N_23007);
xnor U25897 (N_25897,N_23081,N_23709);
nor U25898 (N_25898,N_22501,N_21615);
nor U25899 (N_25899,N_23647,N_21634);
and U25900 (N_25900,N_21045,N_21543);
nand U25901 (N_25901,N_21188,N_22728);
nand U25902 (N_25902,N_23074,N_22969);
or U25903 (N_25903,N_21027,N_23281);
nor U25904 (N_25904,N_21757,N_22482);
nand U25905 (N_25905,N_21468,N_21136);
or U25906 (N_25906,N_21011,N_22952);
and U25907 (N_25907,N_22529,N_22176);
or U25908 (N_25908,N_23122,N_21205);
and U25909 (N_25909,N_22091,N_23301);
and U25910 (N_25910,N_23805,N_22255);
xor U25911 (N_25911,N_23841,N_22947);
or U25912 (N_25912,N_22743,N_21419);
nand U25913 (N_25913,N_23286,N_23358);
and U25914 (N_25914,N_21791,N_22462);
and U25915 (N_25915,N_22998,N_22264);
xnor U25916 (N_25916,N_22778,N_23132);
and U25917 (N_25917,N_22097,N_23899);
and U25918 (N_25918,N_23392,N_23878);
xnor U25919 (N_25919,N_23622,N_22164);
xnor U25920 (N_25920,N_23015,N_21879);
nor U25921 (N_25921,N_21186,N_23956);
xnor U25922 (N_25922,N_21776,N_22951);
xor U25923 (N_25923,N_23590,N_21350);
nand U25924 (N_25924,N_22311,N_23667);
nor U25925 (N_25925,N_21268,N_22688);
or U25926 (N_25926,N_23878,N_21848);
or U25927 (N_25927,N_23979,N_22175);
nor U25928 (N_25928,N_22961,N_21444);
nand U25929 (N_25929,N_22938,N_23264);
and U25930 (N_25930,N_23638,N_22290);
nand U25931 (N_25931,N_21100,N_22209);
xnor U25932 (N_25932,N_21942,N_21998);
or U25933 (N_25933,N_23800,N_21773);
and U25934 (N_25934,N_21755,N_21022);
nand U25935 (N_25935,N_22570,N_22440);
or U25936 (N_25936,N_21171,N_23668);
nand U25937 (N_25937,N_21058,N_23791);
xnor U25938 (N_25938,N_23575,N_21784);
xnor U25939 (N_25939,N_22880,N_21187);
nand U25940 (N_25940,N_21878,N_23829);
xnor U25941 (N_25941,N_22440,N_21404);
nor U25942 (N_25942,N_21577,N_21874);
and U25943 (N_25943,N_23908,N_21650);
or U25944 (N_25944,N_23349,N_22126);
or U25945 (N_25945,N_23105,N_21539);
nand U25946 (N_25946,N_22954,N_21275);
and U25947 (N_25947,N_22032,N_21932);
nor U25948 (N_25948,N_21468,N_22896);
and U25949 (N_25949,N_22466,N_22702);
or U25950 (N_25950,N_23562,N_21973);
xnor U25951 (N_25951,N_21932,N_23916);
or U25952 (N_25952,N_23067,N_23381);
nor U25953 (N_25953,N_22483,N_22487);
nor U25954 (N_25954,N_21112,N_23000);
nand U25955 (N_25955,N_22438,N_21254);
nor U25956 (N_25956,N_21028,N_23695);
and U25957 (N_25957,N_21926,N_22778);
xnor U25958 (N_25958,N_21609,N_23850);
nand U25959 (N_25959,N_23440,N_23059);
nor U25960 (N_25960,N_21452,N_21533);
or U25961 (N_25961,N_23012,N_21502);
and U25962 (N_25962,N_23559,N_23299);
nand U25963 (N_25963,N_21723,N_21211);
xor U25964 (N_25964,N_21192,N_23117);
xor U25965 (N_25965,N_22526,N_22467);
nand U25966 (N_25966,N_23798,N_23377);
nor U25967 (N_25967,N_21577,N_21836);
nand U25968 (N_25968,N_22514,N_21845);
or U25969 (N_25969,N_22466,N_21835);
or U25970 (N_25970,N_22969,N_22279);
nand U25971 (N_25971,N_23892,N_23484);
and U25972 (N_25972,N_23071,N_22344);
nor U25973 (N_25973,N_21949,N_21193);
and U25974 (N_25974,N_22135,N_22693);
xor U25975 (N_25975,N_21200,N_22853);
nor U25976 (N_25976,N_23088,N_22070);
xnor U25977 (N_25977,N_23394,N_21823);
or U25978 (N_25978,N_21715,N_21066);
nand U25979 (N_25979,N_23571,N_22386);
nor U25980 (N_25980,N_23121,N_22497);
or U25981 (N_25981,N_22288,N_21504);
nand U25982 (N_25982,N_22440,N_23324);
or U25983 (N_25983,N_23908,N_23608);
nor U25984 (N_25984,N_21772,N_21763);
nor U25985 (N_25985,N_21794,N_21215);
nand U25986 (N_25986,N_22480,N_22871);
nand U25987 (N_25987,N_23386,N_22841);
nor U25988 (N_25988,N_22835,N_22683);
nand U25989 (N_25989,N_21276,N_22030);
and U25990 (N_25990,N_23445,N_22313);
xnor U25991 (N_25991,N_21209,N_23384);
and U25992 (N_25992,N_23194,N_21965);
or U25993 (N_25993,N_21649,N_21940);
or U25994 (N_25994,N_22369,N_23332);
and U25995 (N_25995,N_22838,N_22335);
nand U25996 (N_25996,N_23908,N_23323);
nand U25997 (N_25997,N_21559,N_23343);
xnor U25998 (N_25998,N_23248,N_23169);
or U25999 (N_25999,N_21012,N_22816);
xnor U26000 (N_26000,N_23158,N_21432);
nand U26001 (N_26001,N_23389,N_23959);
or U26002 (N_26002,N_23781,N_21675);
nand U26003 (N_26003,N_21538,N_22028);
xnor U26004 (N_26004,N_21895,N_21783);
or U26005 (N_26005,N_23831,N_21126);
nand U26006 (N_26006,N_22554,N_22796);
and U26007 (N_26007,N_22075,N_22431);
and U26008 (N_26008,N_21495,N_22284);
nor U26009 (N_26009,N_22198,N_21291);
nor U26010 (N_26010,N_23268,N_23734);
or U26011 (N_26011,N_23948,N_23428);
nand U26012 (N_26012,N_23961,N_23116);
xnor U26013 (N_26013,N_23022,N_21355);
and U26014 (N_26014,N_22685,N_23815);
nand U26015 (N_26015,N_21708,N_21555);
nor U26016 (N_26016,N_22268,N_21930);
nand U26017 (N_26017,N_23482,N_23876);
nand U26018 (N_26018,N_21103,N_22100);
nand U26019 (N_26019,N_22307,N_22578);
nor U26020 (N_26020,N_23297,N_23944);
nor U26021 (N_26021,N_21087,N_22117);
nor U26022 (N_26022,N_23021,N_22109);
or U26023 (N_26023,N_21063,N_23005);
xnor U26024 (N_26024,N_22721,N_23262);
or U26025 (N_26025,N_22982,N_21422);
and U26026 (N_26026,N_22849,N_22341);
nor U26027 (N_26027,N_23484,N_21224);
or U26028 (N_26028,N_23558,N_23721);
and U26029 (N_26029,N_21840,N_21729);
or U26030 (N_26030,N_23033,N_21726);
nand U26031 (N_26031,N_21453,N_22653);
or U26032 (N_26032,N_23227,N_23490);
nor U26033 (N_26033,N_21868,N_21565);
nor U26034 (N_26034,N_21425,N_21299);
nand U26035 (N_26035,N_22729,N_21859);
nor U26036 (N_26036,N_21951,N_23388);
xnor U26037 (N_26037,N_21124,N_21201);
or U26038 (N_26038,N_21587,N_21723);
nand U26039 (N_26039,N_22656,N_21753);
or U26040 (N_26040,N_23251,N_22147);
xnor U26041 (N_26041,N_21538,N_21156);
and U26042 (N_26042,N_23684,N_22877);
or U26043 (N_26043,N_22852,N_23842);
xnor U26044 (N_26044,N_23906,N_23150);
and U26045 (N_26045,N_21611,N_21103);
nand U26046 (N_26046,N_22280,N_22498);
and U26047 (N_26047,N_22103,N_22201);
or U26048 (N_26048,N_21451,N_22369);
nor U26049 (N_26049,N_22846,N_23791);
and U26050 (N_26050,N_23208,N_22894);
nand U26051 (N_26051,N_22378,N_22333);
nor U26052 (N_26052,N_21403,N_21226);
nor U26053 (N_26053,N_23722,N_22760);
nor U26054 (N_26054,N_22924,N_23730);
and U26055 (N_26055,N_22405,N_22376);
nor U26056 (N_26056,N_21909,N_22425);
and U26057 (N_26057,N_22806,N_23740);
nand U26058 (N_26058,N_22484,N_23305);
nor U26059 (N_26059,N_23071,N_21594);
or U26060 (N_26060,N_21563,N_23467);
nand U26061 (N_26061,N_23254,N_22579);
xnor U26062 (N_26062,N_21142,N_23829);
or U26063 (N_26063,N_23383,N_21270);
nor U26064 (N_26064,N_22962,N_22048);
xnor U26065 (N_26065,N_21462,N_23165);
and U26066 (N_26066,N_23566,N_22395);
nor U26067 (N_26067,N_22168,N_23818);
xor U26068 (N_26068,N_22450,N_21215);
or U26069 (N_26069,N_23738,N_21341);
or U26070 (N_26070,N_21936,N_23232);
xor U26071 (N_26071,N_23282,N_21795);
nand U26072 (N_26072,N_22723,N_23215);
and U26073 (N_26073,N_23740,N_21285);
nand U26074 (N_26074,N_22489,N_22318);
or U26075 (N_26075,N_23864,N_23248);
nor U26076 (N_26076,N_22760,N_21088);
xnor U26077 (N_26077,N_23543,N_22044);
xnor U26078 (N_26078,N_23214,N_22594);
nand U26079 (N_26079,N_21544,N_22931);
nor U26080 (N_26080,N_21017,N_22055);
nand U26081 (N_26081,N_23675,N_23511);
nand U26082 (N_26082,N_22779,N_23985);
nor U26083 (N_26083,N_22914,N_22745);
nor U26084 (N_26084,N_21743,N_23388);
or U26085 (N_26085,N_23777,N_23831);
nor U26086 (N_26086,N_22542,N_21664);
and U26087 (N_26087,N_23415,N_21750);
and U26088 (N_26088,N_21479,N_22252);
nand U26089 (N_26089,N_22212,N_21074);
nor U26090 (N_26090,N_23649,N_23265);
nand U26091 (N_26091,N_22744,N_23721);
and U26092 (N_26092,N_23547,N_22883);
nand U26093 (N_26093,N_23584,N_21787);
xor U26094 (N_26094,N_22398,N_22620);
nor U26095 (N_26095,N_21993,N_23845);
nor U26096 (N_26096,N_23948,N_22085);
nand U26097 (N_26097,N_21349,N_22224);
nor U26098 (N_26098,N_22933,N_23039);
and U26099 (N_26099,N_22003,N_21070);
nor U26100 (N_26100,N_21127,N_22524);
and U26101 (N_26101,N_23234,N_22957);
or U26102 (N_26102,N_23976,N_22319);
nor U26103 (N_26103,N_23992,N_22915);
and U26104 (N_26104,N_21002,N_23369);
nor U26105 (N_26105,N_22133,N_21830);
xor U26106 (N_26106,N_21989,N_23024);
or U26107 (N_26107,N_23278,N_21502);
xnor U26108 (N_26108,N_21480,N_23189);
nor U26109 (N_26109,N_23667,N_23595);
or U26110 (N_26110,N_21531,N_22924);
nand U26111 (N_26111,N_22624,N_22563);
nand U26112 (N_26112,N_22709,N_22680);
or U26113 (N_26113,N_21510,N_23470);
or U26114 (N_26114,N_23037,N_23584);
or U26115 (N_26115,N_23488,N_21514);
nor U26116 (N_26116,N_21186,N_23353);
or U26117 (N_26117,N_21332,N_23302);
xnor U26118 (N_26118,N_23494,N_21061);
xor U26119 (N_26119,N_22147,N_23274);
nand U26120 (N_26120,N_23001,N_22900);
xnor U26121 (N_26121,N_22380,N_22338);
or U26122 (N_26122,N_23620,N_23003);
xnor U26123 (N_26123,N_22840,N_21834);
xor U26124 (N_26124,N_22219,N_21116);
and U26125 (N_26125,N_22256,N_22210);
nor U26126 (N_26126,N_23230,N_21258);
nor U26127 (N_26127,N_22726,N_21551);
and U26128 (N_26128,N_21560,N_22665);
and U26129 (N_26129,N_21717,N_23615);
and U26130 (N_26130,N_23409,N_21645);
nand U26131 (N_26131,N_22493,N_22246);
or U26132 (N_26132,N_22616,N_23323);
nor U26133 (N_26133,N_21676,N_21242);
and U26134 (N_26134,N_21304,N_21397);
nand U26135 (N_26135,N_21211,N_23589);
or U26136 (N_26136,N_23631,N_23849);
nand U26137 (N_26137,N_23965,N_22374);
nor U26138 (N_26138,N_22074,N_22073);
nor U26139 (N_26139,N_23464,N_23442);
nand U26140 (N_26140,N_21295,N_23968);
xnor U26141 (N_26141,N_21042,N_22173);
nand U26142 (N_26142,N_21281,N_22613);
nand U26143 (N_26143,N_21479,N_22800);
or U26144 (N_26144,N_22467,N_22260);
xnor U26145 (N_26145,N_22331,N_22178);
or U26146 (N_26146,N_21444,N_23166);
or U26147 (N_26147,N_22204,N_21357);
and U26148 (N_26148,N_21234,N_23996);
and U26149 (N_26149,N_22661,N_22046);
and U26150 (N_26150,N_22604,N_21495);
or U26151 (N_26151,N_23573,N_22809);
xor U26152 (N_26152,N_22823,N_21443);
nor U26153 (N_26153,N_22823,N_21681);
or U26154 (N_26154,N_22147,N_22220);
nand U26155 (N_26155,N_22986,N_23704);
or U26156 (N_26156,N_21583,N_22155);
and U26157 (N_26157,N_21960,N_23356);
and U26158 (N_26158,N_22474,N_21872);
nor U26159 (N_26159,N_21571,N_23002);
nand U26160 (N_26160,N_21778,N_23364);
xnor U26161 (N_26161,N_21325,N_23465);
or U26162 (N_26162,N_21680,N_22387);
or U26163 (N_26163,N_22463,N_22974);
xor U26164 (N_26164,N_22998,N_23699);
nand U26165 (N_26165,N_23972,N_23488);
nand U26166 (N_26166,N_23582,N_21968);
xor U26167 (N_26167,N_23512,N_21707);
nand U26168 (N_26168,N_21908,N_22870);
xor U26169 (N_26169,N_23332,N_21646);
and U26170 (N_26170,N_21020,N_23828);
or U26171 (N_26171,N_23814,N_22949);
or U26172 (N_26172,N_23792,N_21753);
nand U26173 (N_26173,N_21217,N_23808);
and U26174 (N_26174,N_23629,N_22435);
or U26175 (N_26175,N_22775,N_22470);
nand U26176 (N_26176,N_21620,N_21723);
or U26177 (N_26177,N_22191,N_21036);
nor U26178 (N_26178,N_23198,N_21077);
nor U26179 (N_26179,N_22768,N_21719);
nand U26180 (N_26180,N_22092,N_23101);
xnor U26181 (N_26181,N_21932,N_22611);
nor U26182 (N_26182,N_22272,N_22360);
nand U26183 (N_26183,N_21665,N_22695);
xor U26184 (N_26184,N_21968,N_22052);
nor U26185 (N_26185,N_21225,N_21719);
nand U26186 (N_26186,N_22789,N_21787);
and U26187 (N_26187,N_22017,N_22670);
and U26188 (N_26188,N_22925,N_21417);
xnor U26189 (N_26189,N_22363,N_23172);
or U26190 (N_26190,N_23387,N_22786);
or U26191 (N_26191,N_22040,N_22016);
and U26192 (N_26192,N_21666,N_22084);
or U26193 (N_26193,N_21448,N_22231);
or U26194 (N_26194,N_21540,N_21886);
and U26195 (N_26195,N_22741,N_23240);
and U26196 (N_26196,N_23156,N_21132);
nand U26197 (N_26197,N_22711,N_22846);
nand U26198 (N_26198,N_23007,N_22339);
and U26199 (N_26199,N_22810,N_23408);
or U26200 (N_26200,N_21496,N_22987);
and U26201 (N_26201,N_23376,N_21169);
and U26202 (N_26202,N_21695,N_21120);
and U26203 (N_26203,N_21519,N_22982);
nor U26204 (N_26204,N_21054,N_21860);
xor U26205 (N_26205,N_22277,N_23008);
or U26206 (N_26206,N_23358,N_22685);
xor U26207 (N_26207,N_23820,N_22352);
nor U26208 (N_26208,N_21292,N_22637);
xnor U26209 (N_26209,N_22074,N_23263);
xor U26210 (N_26210,N_22809,N_23759);
and U26211 (N_26211,N_21797,N_21856);
or U26212 (N_26212,N_21798,N_21038);
or U26213 (N_26213,N_22437,N_22546);
or U26214 (N_26214,N_21234,N_23987);
or U26215 (N_26215,N_23639,N_23046);
or U26216 (N_26216,N_22523,N_21847);
and U26217 (N_26217,N_22764,N_21713);
nand U26218 (N_26218,N_22362,N_22070);
xnor U26219 (N_26219,N_22911,N_21092);
and U26220 (N_26220,N_23517,N_22294);
nand U26221 (N_26221,N_21045,N_23150);
nand U26222 (N_26222,N_22112,N_22021);
or U26223 (N_26223,N_21139,N_23570);
nand U26224 (N_26224,N_23917,N_22735);
nor U26225 (N_26225,N_21414,N_22732);
nand U26226 (N_26226,N_21755,N_22959);
nor U26227 (N_26227,N_23103,N_23572);
nor U26228 (N_26228,N_23670,N_23229);
xor U26229 (N_26229,N_21748,N_23919);
xor U26230 (N_26230,N_23434,N_23465);
or U26231 (N_26231,N_23577,N_22332);
and U26232 (N_26232,N_21537,N_23155);
or U26233 (N_26233,N_21478,N_22734);
xor U26234 (N_26234,N_21002,N_21436);
nand U26235 (N_26235,N_21439,N_21483);
nor U26236 (N_26236,N_23928,N_23674);
xor U26237 (N_26237,N_22472,N_23679);
xnor U26238 (N_26238,N_22990,N_23515);
and U26239 (N_26239,N_22519,N_23599);
nor U26240 (N_26240,N_21358,N_23998);
nand U26241 (N_26241,N_23832,N_21991);
and U26242 (N_26242,N_22947,N_23328);
and U26243 (N_26243,N_23204,N_21254);
nor U26244 (N_26244,N_23502,N_23083);
nor U26245 (N_26245,N_21541,N_22880);
nor U26246 (N_26246,N_21798,N_22548);
nand U26247 (N_26247,N_22062,N_21654);
xnor U26248 (N_26248,N_22367,N_23925);
nor U26249 (N_26249,N_23363,N_23648);
and U26250 (N_26250,N_23310,N_21326);
xor U26251 (N_26251,N_22701,N_22139);
or U26252 (N_26252,N_21180,N_21095);
and U26253 (N_26253,N_21235,N_22392);
or U26254 (N_26254,N_23646,N_21438);
and U26255 (N_26255,N_23153,N_22392);
xor U26256 (N_26256,N_21562,N_22777);
nor U26257 (N_26257,N_21429,N_23743);
xor U26258 (N_26258,N_22571,N_21906);
and U26259 (N_26259,N_23952,N_21796);
nand U26260 (N_26260,N_23796,N_21739);
xor U26261 (N_26261,N_21913,N_23318);
nand U26262 (N_26262,N_21088,N_21987);
nor U26263 (N_26263,N_22154,N_21708);
and U26264 (N_26264,N_21372,N_23124);
xnor U26265 (N_26265,N_23033,N_22583);
xor U26266 (N_26266,N_22984,N_23501);
nor U26267 (N_26267,N_23485,N_21661);
or U26268 (N_26268,N_22556,N_23412);
xnor U26269 (N_26269,N_21223,N_23467);
xor U26270 (N_26270,N_23627,N_23540);
nand U26271 (N_26271,N_23679,N_22844);
or U26272 (N_26272,N_21184,N_23551);
nor U26273 (N_26273,N_21613,N_23746);
and U26274 (N_26274,N_22757,N_21719);
and U26275 (N_26275,N_21153,N_23698);
xnor U26276 (N_26276,N_21468,N_21037);
and U26277 (N_26277,N_23492,N_23082);
or U26278 (N_26278,N_23550,N_21110);
nand U26279 (N_26279,N_22890,N_23964);
or U26280 (N_26280,N_22785,N_23670);
nor U26281 (N_26281,N_23635,N_23209);
xor U26282 (N_26282,N_23948,N_22468);
nor U26283 (N_26283,N_22898,N_23228);
nor U26284 (N_26284,N_22084,N_22189);
or U26285 (N_26285,N_21521,N_21256);
and U26286 (N_26286,N_21562,N_22066);
xor U26287 (N_26287,N_22491,N_21120);
nand U26288 (N_26288,N_21790,N_21972);
nand U26289 (N_26289,N_23457,N_21068);
nand U26290 (N_26290,N_22502,N_21936);
nand U26291 (N_26291,N_21724,N_22296);
nor U26292 (N_26292,N_23809,N_21050);
nor U26293 (N_26293,N_23624,N_23795);
nor U26294 (N_26294,N_23553,N_22539);
nor U26295 (N_26295,N_23404,N_23130);
nor U26296 (N_26296,N_21903,N_21932);
nand U26297 (N_26297,N_22822,N_22082);
and U26298 (N_26298,N_22894,N_21316);
nand U26299 (N_26299,N_22588,N_23689);
and U26300 (N_26300,N_21657,N_23112);
xnor U26301 (N_26301,N_22008,N_21297);
xor U26302 (N_26302,N_21144,N_22841);
xor U26303 (N_26303,N_22675,N_21134);
xnor U26304 (N_26304,N_23817,N_22445);
nand U26305 (N_26305,N_22804,N_23830);
xnor U26306 (N_26306,N_22779,N_21200);
nand U26307 (N_26307,N_23426,N_23358);
or U26308 (N_26308,N_21005,N_22278);
nor U26309 (N_26309,N_23103,N_22618);
nor U26310 (N_26310,N_22771,N_22874);
nand U26311 (N_26311,N_22091,N_22102);
or U26312 (N_26312,N_23209,N_23824);
nand U26313 (N_26313,N_23083,N_21783);
nor U26314 (N_26314,N_23024,N_22610);
and U26315 (N_26315,N_22470,N_22993);
and U26316 (N_26316,N_21820,N_23065);
nand U26317 (N_26317,N_21540,N_23911);
or U26318 (N_26318,N_23299,N_23186);
nor U26319 (N_26319,N_21568,N_21922);
or U26320 (N_26320,N_23673,N_21383);
xnor U26321 (N_26321,N_23689,N_22231);
nand U26322 (N_26322,N_23279,N_21539);
nand U26323 (N_26323,N_21672,N_23578);
nand U26324 (N_26324,N_21316,N_23908);
nor U26325 (N_26325,N_21573,N_21478);
xor U26326 (N_26326,N_22205,N_21180);
nand U26327 (N_26327,N_21977,N_23490);
xor U26328 (N_26328,N_23445,N_22513);
or U26329 (N_26329,N_23276,N_21156);
or U26330 (N_26330,N_21522,N_21162);
nor U26331 (N_26331,N_22819,N_23069);
and U26332 (N_26332,N_21687,N_23880);
or U26333 (N_26333,N_22181,N_22329);
xor U26334 (N_26334,N_23774,N_22382);
and U26335 (N_26335,N_22064,N_23803);
xnor U26336 (N_26336,N_22963,N_22893);
and U26337 (N_26337,N_23182,N_22486);
nor U26338 (N_26338,N_23400,N_23633);
xor U26339 (N_26339,N_22645,N_21146);
nand U26340 (N_26340,N_22645,N_21228);
xor U26341 (N_26341,N_21567,N_21155);
nand U26342 (N_26342,N_21125,N_23961);
or U26343 (N_26343,N_23695,N_23864);
and U26344 (N_26344,N_21730,N_22624);
xnor U26345 (N_26345,N_22936,N_22706);
and U26346 (N_26346,N_23250,N_23712);
xor U26347 (N_26347,N_21587,N_22471);
xor U26348 (N_26348,N_21090,N_23402);
or U26349 (N_26349,N_23355,N_21401);
nor U26350 (N_26350,N_22028,N_23693);
xor U26351 (N_26351,N_21750,N_21454);
or U26352 (N_26352,N_22237,N_23461);
or U26353 (N_26353,N_22166,N_22704);
and U26354 (N_26354,N_21203,N_23104);
nand U26355 (N_26355,N_23605,N_21539);
nor U26356 (N_26356,N_22072,N_21156);
and U26357 (N_26357,N_21796,N_22800);
or U26358 (N_26358,N_21151,N_23134);
or U26359 (N_26359,N_22972,N_21153);
nand U26360 (N_26360,N_21260,N_22445);
and U26361 (N_26361,N_22794,N_22996);
and U26362 (N_26362,N_22400,N_23257);
or U26363 (N_26363,N_22761,N_22805);
and U26364 (N_26364,N_23128,N_23127);
nor U26365 (N_26365,N_23999,N_21591);
nand U26366 (N_26366,N_23002,N_21573);
xnor U26367 (N_26367,N_21572,N_22317);
xnor U26368 (N_26368,N_23209,N_23758);
or U26369 (N_26369,N_22420,N_21956);
or U26370 (N_26370,N_21801,N_23344);
xor U26371 (N_26371,N_23121,N_21350);
xnor U26372 (N_26372,N_23306,N_22641);
nor U26373 (N_26373,N_22713,N_23922);
and U26374 (N_26374,N_21064,N_23255);
nand U26375 (N_26375,N_21959,N_22688);
or U26376 (N_26376,N_22160,N_23145);
nor U26377 (N_26377,N_23641,N_23900);
nor U26378 (N_26378,N_21748,N_21518);
or U26379 (N_26379,N_22223,N_23416);
xor U26380 (N_26380,N_21082,N_23857);
xor U26381 (N_26381,N_21582,N_23590);
xor U26382 (N_26382,N_21979,N_21017);
and U26383 (N_26383,N_21099,N_22961);
nand U26384 (N_26384,N_22018,N_22887);
xor U26385 (N_26385,N_23471,N_23342);
or U26386 (N_26386,N_22687,N_23116);
nor U26387 (N_26387,N_23997,N_22748);
nand U26388 (N_26388,N_21720,N_23496);
xnor U26389 (N_26389,N_23921,N_21051);
and U26390 (N_26390,N_22193,N_21228);
xnor U26391 (N_26391,N_21281,N_22846);
nand U26392 (N_26392,N_23876,N_22986);
or U26393 (N_26393,N_23772,N_23497);
nand U26394 (N_26394,N_23712,N_21120);
nand U26395 (N_26395,N_22475,N_22582);
and U26396 (N_26396,N_21594,N_23843);
and U26397 (N_26397,N_22697,N_21331);
nand U26398 (N_26398,N_22194,N_21180);
nor U26399 (N_26399,N_23441,N_22419);
xnor U26400 (N_26400,N_22394,N_23632);
nor U26401 (N_26401,N_21270,N_21086);
nand U26402 (N_26402,N_21816,N_22806);
nor U26403 (N_26403,N_23276,N_23872);
nor U26404 (N_26404,N_21711,N_21373);
and U26405 (N_26405,N_21279,N_22681);
xnor U26406 (N_26406,N_22543,N_22343);
and U26407 (N_26407,N_22506,N_23787);
or U26408 (N_26408,N_22520,N_21479);
nor U26409 (N_26409,N_23290,N_22221);
or U26410 (N_26410,N_22303,N_21908);
or U26411 (N_26411,N_21580,N_21407);
nand U26412 (N_26412,N_22448,N_21904);
xnor U26413 (N_26413,N_21087,N_21455);
or U26414 (N_26414,N_22218,N_23743);
nand U26415 (N_26415,N_23039,N_21961);
and U26416 (N_26416,N_22153,N_22456);
nor U26417 (N_26417,N_21320,N_21033);
nor U26418 (N_26418,N_23822,N_23201);
nor U26419 (N_26419,N_22506,N_23688);
xnor U26420 (N_26420,N_23803,N_21718);
nand U26421 (N_26421,N_21943,N_22372);
or U26422 (N_26422,N_21327,N_21318);
nand U26423 (N_26423,N_22617,N_23730);
nor U26424 (N_26424,N_21023,N_22587);
or U26425 (N_26425,N_22551,N_22183);
nand U26426 (N_26426,N_22915,N_21001);
nand U26427 (N_26427,N_23397,N_21482);
and U26428 (N_26428,N_21025,N_22572);
nand U26429 (N_26429,N_22651,N_21501);
nor U26430 (N_26430,N_21298,N_21637);
xor U26431 (N_26431,N_21939,N_23818);
nand U26432 (N_26432,N_23794,N_21901);
nand U26433 (N_26433,N_22196,N_22763);
or U26434 (N_26434,N_21457,N_23623);
and U26435 (N_26435,N_23258,N_22347);
and U26436 (N_26436,N_21210,N_23756);
and U26437 (N_26437,N_23598,N_22393);
nand U26438 (N_26438,N_21175,N_22919);
xnor U26439 (N_26439,N_22139,N_22440);
xnor U26440 (N_26440,N_23487,N_23225);
nand U26441 (N_26441,N_22069,N_21510);
nand U26442 (N_26442,N_22277,N_21318);
nor U26443 (N_26443,N_21211,N_22445);
xor U26444 (N_26444,N_23810,N_23059);
and U26445 (N_26445,N_22233,N_22121);
nand U26446 (N_26446,N_22186,N_21849);
or U26447 (N_26447,N_23194,N_23476);
xor U26448 (N_26448,N_22013,N_23421);
or U26449 (N_26449,N_22019,N_22221);
xnor U26450 (N_26450,N_21541,N_21547);
xnor U26451 (N_26451,N_22592,N_22597);
and U26452 (N_26452,N_21238,N_21836);
nor U26453 (N_26453,N_23555,N_23694);
nand U26454 (N_26454,N_23306,N_21565);
and U26455 (N_26455,N_22362,N_23947);
nor U26456 (N_26456,N_22084,N_22553);
nor U26457 (N_26457,N_21004,N_23726);
or U26458 (N_26458,N_21287,N_22970);
or U26459 (N_26459,N_21979,N_22036);
or U26460 (N_26460,N_21984,N_21484);
xor U26461 (N_26461,N_22845,N_22194);
xor U26462 (N_26462,N_21053,N_22211);
nand U26463 (N_26463,N_21031,N_21599);
or U26464 (N_26464,N_21511,N_21205);
and U26465 (N_26465,N_23842,N_21310);
nor U26466 (N_26466,N_21994,N_21466);
and U26467 (N_26467,N_22673,N_21638);
nand U26468 (N_26468,N_21422,N_23135);
and U26469 (N_26469,N_23657,N_22512);
nand U26470 (N_26470,N_22468,N_23124);
or U26471 (N_26471,N_22440,N_22967);
xnor U26472 (N_26472,N_21379,N_21022);
and U26473 (N_26473,N_22553,N_22383);
or U26474 (N_26474,N_21404,N_23909);
xor U26475 (N_26475,N_21721,N_21648);
nor U26476 (N_26476,N_23049,N_22397);
and U26477 (N_26477,N_21944,N_23819);
and U26478 (N_26478,N_22903,N_23055);
or U26479 (N_26479,N_22336,N_23887);
nor U26480 (N_26480,N_23986,N_23016);
or U26481 (N_26481,N_23933,N_21982);
or U26482 (N_26482,N_22914,N_23213);
nand U26483 (N_26483,N_22464,N_22325);
nand U26484 (N_26484,N_22908,N_22630);
xor U26485 (N_26485,N_22168,N_21467);
nand U26486 (N_26486,N_22306,N_23241);
and U26487 (N_26487,N_21449,N_23952);
nor U26488 (N_26488,N_23096,N_22842);
and U26489 (N_26489,N_21153,N_23946);
and U26490 (N_26490,N_21707,N_21074);
xor U26491 (N_26491,N_21475,N_21232);
or U26492 (N_26492,N_22843,N_23845);
or U26493 (N_26493,N_22675,N_22035);
nor U26494 (N_26494,N_23358,N_21631);
nor U26495 (N_26495,N_21082,N_23358);
nor U26496 (N_26496,N_21187,N_22149);
nand U26497 (N_26497,N_22674,N_23833);
and U26498 (N_26498,N_21346,N_21101);
or U26499 (N_26499,N_21227,N_23111);
or U26500 (N_26500,N_23348,N_22507);
and U26501 (N_26501,N_22009,N_23535);
or U26502 (N_26502,N_21934,N_22944);
and U26503 (N_26503,N_22243,N_21702);
nand U26504 (N_26504,N_21930,N_21332);
nor U26505 (N_26505,N_21134,N_23082);
or U26506 (N_26506,N_22650,N_21559);
nand U26507 (N_26507,N_21427,N_21829);
nand U26508 (N_26508,N_22303,N_21183);
nand U26509 (N_26509,N_21394,N_23654);
nor U26510 (N_26510,N_22752,N_21081);
and U26511 (N_26511,N_22934,N_22463);
and U26512 (N_26512,N_22730,N_21304);
xnor U26513 (N_26513,N_23030,N_23804);
xnor U26514 (N_26514,N_23650,N_22588);
nor U26515 (N_26515,N_21807,N_23496);
and U26516 (N_26516,N_22571,N_23098);
nor U26517 (N_26517,N_21722,N_21699);
xor U26518 (N_26518,N_21723,N_23549);
or U26519 (N_26519,N_23427,N_23292);
or U26520 (N_26520,N_21894,N_21706);
xnor U26521 (N_26521,N_23365,N_23149);
or U26522 (N_26522,N_21410,N_21481);
nand U26523 (N_26523,N_23576,N_23454);
nor U26524 (N_26524,N_21504,N_22094);
nand U26525 (N_26525,N_23392,N_23500);
nor U26526 (N_26526,N_23739,N_22774);
and U26527 (N_26527,N_22994,N_21133);
nand U26528 (N_26528,N_23435,N_21444);
and U26529 (N_26529,N_23092,N_23855);
xnor U26530 (N_26530,N_23784,N_21095);
xor U26531 (N_26531,N_22019,N_23134);
nand U26532 (N_26532,N_21843,N_21269);
and U26533 (N_26533,N_23469,N_21411);
and U26534 (N_26534,N_22433,N_21925);
nor U26535 (N_26535,N_22467,N_21957);
xor U26536 (N_26536,N_22886,N_22811);
or U26537 (N_26537,N_22636,N_21400);
xnor U26538 (N_26538,N_23663,N_23729);
xor U26539 (N_26539,N_21404,N_21860);
and U26540 (N_26540,N_23559,N_21071);
nor U26541 (N_26541,N_21257,N_22099);
nor U26542 (N_26542,N_22807,N_23964);
and U26543 (N_26543,N_23156,N_23111);
or U26544 (N_26544,N_22148,N_23729);
nor U26545 (N_26545,N_21056,N_23527);
and U26546 (N_26546,N_23596,N_22586);
and U26547 (N_26547,N_22345,N_23223);
and U26548 (N_26548,N_22518,N_21586);
nor U26549 (N_26549,N_23171,N_23840);
and U26550 (N_26550,N_23598,N_21267);
and U26551 (N_26551,N_21726,N_21542);
nor U26552 (N_26552,N_23454,N_22336);
nand U26553 (N_26553,N_23618,N_21852);
xnor U26554 (N_26554,N_22315,N_21059);
and U26555 (N_26555,N_23577,N_23540);
or U26556 (N_26556,N_21444,N_21218);
or U26557 (N_26557,N_22062,N_22514);
or U26558 (N_26558,N_22922,N_23966);
or U26559 (N_26559,N_22419,N_22464);
and U26560 (N_26560,N_21206,N_23755);
or U26561 (N_26561,N_23062,N_22394);
or U26562 (N_26562,N_21592,N_21080);
nor U26563 (N_26563,N_23646,N_21629);
nand U26564 (N_26564,N_21553,N_23534);
nand U26565 (N_26565,N_22984,N_22966);
nand U26566 (N_26566,N_22048,N_21574);
nor U26567 (N_26567,N_21629,N_21052);
xnor U26568 (N_26568,N_21666,N_21339);
nand U26569 (N_26569,N_23373,N_23020);
nand U26570 (N_26570,N_22659,N_21412);
or U26571 (N_26571,N_22034,N_21072);
xor U26572 (N_26572,N_21470,N_22418);
xor U26573 (N_26573,N_23929,N_22648);
nand U26574 (N_26574,N_23920,N_23401);
and U26575 (N_26575,N_22236,N_23935);
nor U26576 (N_26576,N_22151,N_23308);
and U26577 (N_26577,N_22393,N_22635);
nor U26578 (N_26578,N_23073,N_22871);
nor U26579 (N_26579,N_23445,N_23388);
and U26580 (N_26580,N_21450,N_23945);
nor U26581 (N_26581,N_23477,N_21405);
xor U26582 (N_26582,N_22646,N_22308);
nand U26583 (N_26583,N_21512,N_23746);
nor U26584 (N_26584,N_23513,N_23125);
or U26585 (N_26585,N_21306,N_22073);
or U26586 (N_26586,N_21779,N_21682);
and U26587 (N_26587,N_21101,N_22220);
nand U26588 (N_26588,N_23636,N_21360);
and U26589 (N_26589,N_22307,N_22946);
and U26590 (N_26590,N_23941,N_22618);
or U26591 (N_26591,N_21392,N_22754);
and U26592 (N_26592,N_22375,N_21166);
xor U26593 (N_26593,N_21159,N_23935);
nor U26594 (N_26594,N_21515,N_21178);
nor U26595 (N_26595,N_23644,N_21581);
nand U26596 (N_26596,N_22385,N_21961);
and U26597 (N_26597,N_21686,N_21280);
xor U26598 (N_26598,N_22299,N_23846);
xor U26599 (N_26599,N_21126,N_23133);
xnor U26600 (N_26600,N_21152,N_22352);
nor U26601 (N_26601,N_23920,N_23313);
xor U26602 (N_26602,N_22608,N_21232);
and U26603 (N_26603,N_21460,N_21230);
nor U26604 (N_26604,N_22331,N_23929);
or U26605 (N_26605,N_22625,N_22655);
nor U26606 (N_26606,N_21683,N_21268);
and U26607 (N_26607,N_21399,N_23050);
nand U26608 (N_26608,N_22051,N_21532);
nor U26609 (N_26609,N_22630,N_21748);
nor U26610 (N_26610,N_22900,N_23716);
and U26611 (N_26611,N_22561,N_22596);
nand U26612 (N_26612,N_22002,N_22396);
xnor U26613 (N_26613,N_21065,N_22801);
xnor U26614 (N_26614,N_22370,N_23596);
nand U26615 (N_26615,N_21986,N_21533);
or U26616 (N_26616,N_22080,N_21603);
nand U26617 (N_26617,N_23589,N_21650);
or U26618 (N_26618,N_22599,N_21918);
xor U26619 (N_26619,N_22035,N_23673);
and U26620 (N_26620,N_21441,N_23124);
nand U26621 (N_26621,N_23524,N_21151);
nand U26622 (N_26622,N_21185,N_22221);
xor U26623 (N_26623,N_21929,N_21384);
xnor U26624 (N_26624,N_22284,N_23808);
or U26625 (N_26625,N_22283,N_22915);
nand U26626 (N_26626,N_22688,N_22390);
nand U26627 (N_26627,N_22447,N_21394);
xnor U26628 (N_26628,N_21142,N_21881);
xor U26629 (N_26629,N_22344,N_21249);
and U26630 (N_26630,N_23285,N_21174);
nor U26631 (N_26631,N_23463,N_23178);
and U26632 (N_26632,N_23373,N_21129);
and U26633 (N_26633,N_21922,N_21650);
xor U26634 (N_26634,N_23701,N_23355);
or U26635 (N_26635,N_22104,N_21372);
nand U26636 (N_26636,N_23402,N_21648);
nand U26637 (N_26637,N_22096,N_23628);
xnor U26638 (N_26638,N_23723,N_22994);
xor U26639 (N_26639,N_21282,N_23610);
and U26640 (N_26640,N_22080,N_23971);
nor U26641 (N_26641,N_23094,N_22434);
or U26642 (N_26642,N_22631,N_23950);
and U26643 (N_26643,N_22190,N_23855);
nor U26644 (N_26644,N_22601,N_22605);
or U26645 (N_26645,N_22815,N_22692);
or U26646 (N_26646,N_22036,N_22896);
xor U26647 (N_26647,N_23070,N_21793);
nor U26648 (N_26648,N_21136,N_22163);
nand U26649 (N_26649,N_22731,N_22780);
nand U26650 (N_26650,N_23176,N_22332);
nand U26651 (N_26651,N_22827,N_22338);
or U26652 (N_26652,N_23098,N_23458);
nand U26653 (N_26653,N_22965,N_21625);
or U26654 (N_26654,N_22154,N_23225);
or U26655 (N_26655,N_22111,N_23299);
xnor U26656 (N_26656,N_23650,N_22148);
nor U26657 (N_26657,N_22162,N_23877);
xor U26658 (N_26658,N_22957,N_22436);
xnor U26659 (N_26659,N_21775,N_23100);
nand U26660 (N_26660,N_21340,N_22835);
xor U26661 (N_26661,N_22435,N_22584);
nand U26662 (N_26662,N_22714,N_23617);
or U26663 (N_26663,N_23598,N_21575);
xnor U26664 (N_26664,N_23922,N_23197);
xor U26665 (N_26665,N_21083,N_21764);
or U26666 (N_26666,N_21619,N_23202);
or U26667 (N_26667,N_22500,N_23530);
or U26668 (N_26668,N_23160,N_22828);
nand U26669 (N_26669,N_21347,N_21278);
or U26670 (N_26670,N_22781,N_21961);
or U26671 (N_26671,N_21426,N_22911);
nand U26672 (N_26672,N_22139,N_21294);
nor U26673 (N_26673,N_21604,N_22484);
nand U26674 (N_26674,N_22461,N_23074);
nor U26675 (N_26675,N_21069,N_23471);
and U26676 (N_26676,N_23747,N_22470);
or U26677 (N_26677,N_21683,N_23052);
nand U26678 (N_26678,N_22587,N_21034);
and U26679 (N_26679,N_22911,N_22591);
nand U26680 (N_26680,N_22503,N_21385);
and U26681 (N_26681,N_23275,N_22966);
or U26682 (N_26682,N_22667,N_23781);
nand U26683 (N_26683,N_22311,N_22481);
nor U26684 (N_26684,N_23485,N_23505);
nor U26685 (N_26685,N_22620,N_23277);
xor U26686 (N_26686,N_22075,N_22743);
and U26687 (N_26687,N_21912,N_23240);
nor U26688 (N_26688,N_21610,N_22347);
and U26689 (N_26689,N_22130,N_22891);
or U26690 (N_26690,N_23742,N_21446);
or U26691 (N_26691,N_22471,N_22588);
or U26692 (N_26692,N_22130,N_23684);
or U26693 (N_26693,N_22337,N_21496);
xnor U26694 (N_26694,N_22352,N_23096);
nand U26695 (N_26695,N_22295,N_22091);
nor U26696 (N_26696,N_23599,N_22615);
nor U26697 (N_26697,N_23769,N_23894);
and U26698 (N_26698,N_22660,N_21799);
nand U26699 (N_26699,N_23700,N_23558);
or U26700 (N_26700,N_22697,N_22225);
nand U26701 (N_26701,N_23214,N_21991);
nand U26702 (N_26702,N_22830,N_22871);
or U26703 (N_26703,N_21241,N_23896);
or U26704 (N_26704,N_21876,N_23636);
nand U26705 (N_26705,N_21102,N_23053);
and U26706 (N_26706,N_21003,N_22802);
and U26707 (N_26707,N_22165,N_23269);
xor U26708 (N_26708,N_23875,N_21627);
nor U26709 (N_26709,N_21990,N_21886);
nand U26710 (N_26710,N_23712,N_22507);
nand U26711 (N_26711,N_22759,N_23227);
xor U26712 (N_26712,N_23233,N_22396);
or U26713 (N_26713,N_21982,N_23723);
and U26714 (N_26714,N_22185,N_21896);
xor U26715 (N_26715,N_23379,N_23030);
nor U26716 (N_26716,N_21962,N_21089);
nand U26717 (N_26717,N_22110,N_22460);
nor U26718 (N_26718,N_22062,N_22231);
xor U26719 (N_26719,N_21471,N_23767);
and U26720 (N_26720,N_21713,N_23016);
xor U26721 (N_26721,N_23552,N_23026);
nand U26722 (N_26722,N_23506,N_22196);
nand U26723 (N_26723,N_23248,N_21150);
nor U26724 (N_26724,N_22161,N_23671);
or U26725 (N_26725,N_21473,N_23175);
nand U26726 (N_26726,N_21457,N_21169);
xnor U26727 (N_26727,N_23601,N_21479);
xor U26728 (N_26728,N_22415,N_21426);
or U26729 (N_26729,N_22590,N_22090);
xor U26730 (N_26730,N_21956,N_23933);
or U26731 (N_26731,N_23647,N_22797);
xor U26732 (N_26732,N_23754,N_22450);
and U26733 (N_26733,N_21041,N_21896);
xnor U26734 (N_26734,N_23855,N_22666);
and U26735 (N_26735,N_21610,N_22565);
and U26736 (N_26736,N_21990,N_22988);
nor U26737 (N_26737,N_22974,N_22856);
and U26738 (N_26738,N_22381,N_23385);
xor U26739 (N_26739,N_23545,N_23113);
and U26740 (N_26740,N_22347,N_22642);
and U26741 (N_26741,N_23010,N_21074);
or U26742 (N_26742,N_23707,N_21578);
and U26743 (N_26743,N_21737,N_21989);
or U26744 (N_26744,N_23532,N_23033);
nand U26745 (N_26745,N_22546,N_21519);
xnor U26746 (N_26746,N_22360,N_23480);
nor U26747 (N_26747,N_23543,N_21348);
nor U26748 (N_26748,N_23638,N_22159);
nor U26749 (N_26749,N_21177,N_21643);
nor U26750 (N_26750,N_21494,N_23495);
nand U26751 (N_26751,N_23933,N_21325);
nor U26752 (N_26752,N_23559,N_21023);
or U26753 (N_26753,N_21511,N_22707);
xnor U26754 (N_26754,N_22852,N_21207);
nand U26755 (N_26755,N_21856,N_21379);
or U26756 (N_26756,N_22120,N_22679);
and U26757 (N_26757,N_21945,N_22872);
nand U26758 (N_26758,N_21145,N_23765);
xnor U26759 (N_26759,N_21482,N_23692);
xnor U26760 (N_26760,N_22752,N_21577);
or U26761 (N_26761,N_23783,N_22542);
xnor U26762 (N_26762,N_22614,N_22026);
and U26763 (N_26763,N_21470,N_21712);
and U26764 (N_26764,N_21855,N_21425);
nand U26765 (N_26765,N_21618,N_22953);
nand U26766 (N_26766,N_22485,N_23934);
nor U26767 (N_26767,N_23075,N_22451);
and U26768 (N_26768,N_23092,N_22001);
and U26769 (N_26769,N_21447,N_21327);
and U26770 (N_26770,N_21008,N_22217);
xor U26771 (N_26771,N_21027,N_21902);
or U26772 (N_26772,N_22104,N_21172);
xor U26773 (N_26773,N_23020,N_22467);
or U26774 (N_26774,N_22526,N_22432);
xor U26775 (N_26775,N_23573,N_23024);
or U26776 (N_26776,N_22836,N_22797);
nand U26777 (N_26777,N_21300,N_21010);
nor U26778 (N_26778,N_23989,N_23344);
and U26779 (N_26779,N_23626,N_23821);
or U26780 (N_26780,N_22667,N_22644);
nand U26781 (N_26781,N_21988,N_22618);
or U26782 (N_26782,N_23840,N_22740);
and U26783 (N_26783,N_22894,N_22310);
xnor U26784 (N_26784,N_22891,N_22408);
nor U26785 (N_26785,N_23974,N_21692);
or U26786 (N_26786,N_22127,N_23221);
xnor U26787 (N_26787,N_23081,N_21077);
xnor U26788 (N_26788,N_23055,N_23342);
or U26789 (N_26789,N_23048,N_22690);
nor U26790 (N_26790,N_22721,N_23666);
or U26791 (N_26791,N_22002,N_22615);
nor U26792 (N_26792,N_21010,N_23695);
or U26793 (N_26793,N_22148,N_23018);
xor U26794 (N_26794,N_22222,N_21768);
nand U26795 (N_26795,N_22099,N_23144);
xor U26796 (N_26796,N_21018,N_21701);
nand U26797 (N_26797,N_22404,N_22157);
xor U26798 (N_26798,N_21762,N_23657);
xor U26799 (N_26799,N_23305,N_23081);
xnor U26800 (N_26800,N_23422,N_21254);
xor U26801 (N_26801,N_21489,N_23311);
or U26802 (N_26802,N_23289,N_22579);
nand U26803 (N_26803,N_23400,N_21264);
nor U26804 (N_26804,N_22656,N_23278);
xnor U26805 (N_26805,N_23675,N_22332);
or U26806 (N_26806,N_22259,N_21246);
nand U26807 (N_26807,N_23659,N_22913);
xnor U26808 (N_26808,N_21885,N_22096);
nand U26809 (N_26809,N_22815,N_21299);
xnor U26810 (N_26810,N_21521,N_21970);
and U26811 (N_26811,N_23525,N_21936);
nand U26812 (N_26812,N_23727,N_21300);
xnor U26813 (N_26813,N_21877,N_23336);
nand U26814 (N_26814,N_22712,N_21249);
or U26815 (N_26815,N_23916,N_22285);
nand U26816 (N_26816,N_23949,N_21838);
nand U26817 (N_26817,N_22415,N_23584);
nand U26818 (N_26818,N_23055,N_21351);
nor U26819 (N_26819,N_21061,N_22942);
xor U26820 (N_26820,N_21004,N_22422);
xor U26821 (N_26821,N_22292,N_22999);
and U26822 (N_26822,N_23955,N_22174);
nand U26823 (N_26823,N_21310,N_22220);
nor U26824 (N_26824,N_23113,N_23490);
nand U26825 (N_26825,N_23475,N_21482);
or U26826 (N_26826,N_23326,N_21422);
nand U26827 (N_26827,N_22729,N_22378);
nor U26828 (N_26828,N_21843,N_23303);
or U26829 (N_26829,N_23068,N_21888);
nor U26830 (N_26830,N_22703,N_21537);
or U26831 (N_26831,N_21749,N_21691);
and U26832 (N_26832,N_22484,N_23064);
xor U26833 (N_26833,N_22253,N_22712);
nor U26834 (N_26834,N_21084,N_23364);
nand U26835 (N_26835,N_21629,N_21102);
nor U26836 (N_26836,N_21468,N_23645);
nor U26837 (N_26837,N_22947,N_23737);
nor U26838 (N_26838,N_21292,N_21684);
xnor U26839 (N_26839,N_23865,N_22086);
nand U26840 (N_26840,N_23216,N_23448);
nand U26841 (N_26841,N_22738,N_21577);
xnor U26842 (N_26842,N_23955,N_23912);
and U26843 (N_26843,N_23589,N_21594);
or U26844 (N_26844,N_21464,N_23688);
or U26845 (N_26845,N_23529,N_22948);
nand U26846 (N_26846,N_21996,N_23594);
nor U26847 (N_26847,N_22798,N_23169);
or U26848 (N_26848,N_23814,N_22649);
nor U26849 (N_26849,N_23609,N_21967);
nor U26850 (N_26850,N_22762,N_21919);
nand U26851 (N_26851,N_23114,N_23845);
nor U26852 (N_26852,N_21744,N_22029);
xnor U26853 (N_26853,N_22963,N_22525);
xnor U26854 (N_26854,N_22424,N_21650);
or U26855 (N_26855,N_22771,N_21940);
nand U26856 (N_26856,N_21849,N_23628);
nand U26857 (N_26857,N_21493,N_22785);
and U26858 (N_26858,N_22764,N_23976);
nand U26859 (N_26859,N_22806,N_23247);
nand U26860 (N_26860,N_21501,N_22345);
nor U26861 (N_26861,N_21835,N_21066);
nand U26862 (N_26862,N_22541,N_23445);
and U26863 (N_26863,N_22568,N_22659);
or U26864 (N_26864,N_23456,N_23742);
or U26865 (N_26865,N_23530,N_23967);
or U26866 (N_26866,N_21894,N_21361);
xnor U26867 (N_26867,N_23816,N_23326);
and U26868 (N_26868,N_21997,N_21488);
xnor U26869 (N_26869,N_22543,N_23069);
nand U26870 (N_26870,N_23552,N_22508);
or U26871 (N_26871,N_22189,N_23316);
or U26872 (N_26872,N_23996,N_21658);
nor U26873 (N_26873,N_23828,N_23803);
xnor U26874 (N_26874,N_21846,N_22696);
nand U26875 (N_26875,N_22772,N_22728);
and U26876 (N_26876,N_21873,N_22840);
xor U26877 (N_26877,N_22780,N_22939);
nand U26878 (N_26878,N_21984,N_21233);
nor U26879 (N_26879,N_22555,N_21356);
nand U26880 (N_26880,N_21809,N_21198);
or U26881 (N_26881,N_21334,N_22293);
xor U26882 (N_26882,N_21033,N_22684);
and U26883 (N_26883,N_21292,N_23446);
or U26884 (N_26884,N_21701,N_23264);
nand U26885 (N_26885,N_23133,N_21802);
or U26886 (N_26886,N_22660,N_21279);
nand U26887 (N_26887,N_23992,N_22130);
nor U26888 (N_26888,N_21752,N_21111);
or U26889 (N_26889,N_21845,N_22575);
nor U26890 (N_26890,N_23166,N_21349);
and U26891 (N_26891,N_22046,N_23337);
xor U26892 (N_26892,N_21840,N_23856);
xnor U26893 (N_26893,N_22613,N_23705);
nor U26894 (N_26894,N_21346,N_23047);
or U26895 (N_26895,N_22978,N_22422);
xnor U26896 (N_26896,N_21357,N_23579);
nor U26897 (N_26897,N_23848,N_21577);
or U26898 (N_26898,N_22739,N_22638);
nand U26899 (N_26899,N_23900,N_21433);
and U26900 (N_26900,N_21341,N_21243);
nand U26901 (N_26901,N_22491,N_21642);
nor U26902 (N_26902,N_23352,N_22585);
or U26903 (N_26903,N_22803,N_23960);
and U26904 (N_26904,N_23192,N_23327);
nand U26905 (N_26905,N_22950,N_23820);
and U26906 (N_26906,N_22361,N_22558);
nand U26907 (N_26907,N_22608,N_23257);
nand U26908 (N_26908,N_21642,N_23979);
nand U26909 (N_26909,N_21489,N_23256);
and U26910 (N_26910,N_21005,N_22841);
nor U26911 (N_26911,N_21188,N_21467);
nor U26912 (N_26912,N_23641,N_21817);
or U26913 (N_26913,N_21119,N_21252);
nor U26914 (N_26914,N_21618,N_23902);
and U26915 (N_26915,N_21555,N_22379);
or U26916 (N_26916,N_23377,N_22849);
nand U26917 (N_26917,N_21957,N_22366);
xor U26918 (N_26918,N_22978,N_23870);
xnor U26919 (N_26919,N_22611,N_21704);
and U26920 (N_26920,N_22918,N_21051);
nand U26921 (N_26921,N_23426,N_21417);
or U26922 (N_26922,N_21845,N_22680);
and U26923 (N_26923,N_21134,N_23958);
nand U26924 (N_26924,N_22097,N_21566);
nor U26925 (N_26925,N_23144,N_23518);
and U26926 (N_26926,N_23149,N_21734);
nand U26927 (N_26927,N_23107,N_22800);
nor U26928 (N_26928,N_22419,N_21323);
and U26929 (N_26929,N_22323,N_22173);
and U26930 (N_26930,N_23705,N_23906);
nand U26931 (N_26931,N_21140,N_22544);
and U26932 (N_26932,N_21147,N_21324);
xnor U26933 (N_26933,N_21475,N_22630);
nand U26934 (N_26934,N_23658,N_23944);
xnor U26935 (N_26935,N_22985,N_22913);
nand U26936 (N_26936,N_21144,N_23031);
nor U26937 (N_26937,N_23060,N_21690);
xor U26938 (N_26938,N_22130,N_22685);
or U26939 (N_26939,N_22452,N_23306);
nand U26940 (N_26940,N_22227,N_21981);
nand U26941 (N_26941,N_23516,N_21021);
and U26942 (N_26942,N_23636,N_23891);
or U26943 (N_26943,N_22540,N_22097);
nor U26944 (N_26944,N_23478,N_21602);
nand U26945 (N_26945,N_22501,N_21894);
nand U26946 (N_26946,N_21035,N_22627);
nor U26947 (N_26947,N_23297,N_21935);
xnor U26948 (N_26948,N_22368,N_21240);
nor U26949 (N_26949,N_22829,N_22509);
nor U26950 (N_26950,N_22164,N_22091);
or U26951 (N_26951,N_21555,N_22863);
nand U26952 (N_26952,N_22037,N_22418);
xor U26953 (N_26953,N_21758,N_21018);
and U26954 (N_26954,N_23135,N_23530);
and U26955 (N_26955,N_23694,N_23707);
nand U26956 (N_26956,N_23309,N_22579);
and U26957 (N_26957,N_23748,N_22481);
xnor U26958 (N_26958,N_22314,N_22382);
or U26959 (N_26959,N_23968,N_22818);
nand U26960 (N_26960,N_22562,N_22541);
or U26961 (N_26961,N_22305,N_21783);
xnor U26962 (N_26962,N_21340,N_23670);
and U26963 (N_26963,N_23242,N_23731);
and U26964 (N_26964,N_21900,N_21046);
and U26965 (N_26965,N_23930,N_22206);
and U26966 (N_26966,N_22906,N_23402);
xnor U26967 (N_26967,N_23714,N_22583);
nand U26968 (N_26968,N_23221,N_23392);
or U26969 (N_26969,N_22490,N_22081);
nor U26970 (N_26970,N_21930,N_22377);
nand U26971 (N_26971,N_22192,N_22846);
nor U26972 (N_26972,N_22899,N_21656);
nand U26973 (N_26973,N_21554,N_22304);
and U26974 (N_26974,N_23802,N_22285);
or U26975 (N_26975,N_22537,N_21552);
nor U26976 (N_26976,N_23110,N_22915);
nor U26977 (N_26977,N_21580,N_23008);
or U26978 (N_26978,N_23891,N_22082);
nand U26979 (N_26979,N_22212,N_22462);
nor U26980 (N_26980,N_22550,N_23699);
and U26981 (N_26981,N_22456,N_23515);
and U26982 (N_26982,N_22467,N_23134);
or U26983 (N_26983,N_23027,N_23228);
xnor U26984 (N_26984,N_21166,N_22170);
nand U26985 (N_26985,N_21316,N_21613);
xor U26986 (N_26986,N_21808,N_22031);
nand U26987 (N_26987,N_21975,N_22753);
nor U26988 (N_26988,N_23647,N_21793);
xor U26989 (N_26989,N_22589,N_22514);
xnor U26990 (N_26990,N_21456,N_23333);
and U26991 (N_26991,N_23056,N_22184);
or U26992 (N_26992,N_22294,N_22241);
xnor U26993 (N_26993,N_23990,N_21423);
xnor U26994 (N_26994,N_21975,N_21546);
or U26995 (N_26995,N_23335,N_21583);
xor U26996 (N_26996,N_22315,N_23223);
or U26997 (N_26997,N_21916,N_22777);
or U26998 (N_26998,N_23465,N_22323);
nor U26999 (N_26999,N_23244,N_21963);
nor U27000 (N_27000,N_25684,N_26606);
or U27001 (N_27001,N_24214,N_24242);
or U27002 (N_27002,N_25677,N_24460);
xnor U27003 (N_27003,N_25175,N_25533);
nand U27004 (N_27004,N_26694,N_26894);
or U27005 (N_27005,N_26443,N_25129);
nor U27006 (N_27006,N_24355,N_25247);
nor U27007 (N_27007,N_25358,N_25315);
xor U27008 (N_27008,N_24522,N_25950);
or U27009 (N_27009,N_24891,N_24649);
and U27010 (N_27010,N_26773,N_25923);
or U27011 (N_27011,N_26793,N_26088);
nor U27012 (N_27012,N_25423,N_25110);
xnor U27013 (N_27013,N_25203,N_24695);
nor U27014 (N_27014,N_24055,N_24640);
nor U27015 (N_27015,N_24863,N_24995);
nand U27016 (N_27016,N_24105,N_26833);
nand U27017 (N_27017,N_24315,N_25820);
and U27018 (N_27018,N_25137,N_26180);
or U27019 (N_27019,N_26242,N_26387);
or U27020 (N_27020,N_26811,N_25683);
nand U27021 (N_27021,N_26484,N_26726);
or U27022 (N_27022,N_26255,N_25335);
xor U27023 (N_27023,N_26620,N_26917);
nand U27024 (N_27024,N_26536,N_26083);
nor U27025 (N_27025,N_25093,N_25316);
or U27026 (N_27026,N_24630,N_25706);
or U27027 (N_27027,N_24339,N_26452);
or U27028 (N_27028,N_24674,N_24685);
or U27029 (N_27029,N_24171,N_26377);
or U27030 (N_27030,N_25492,N_25141);
or U27031 (N_27031,N_26134,N_25027);
nor U27032 (N_27032,N_25859,N_26265);
xnor U27033 (N_27033,N_24837,N_25135);
nand U27034 (N_27034,N_25075,N_24806);
and U27035 (N_27035,N_25696,N_25451);
nor U27036 (N_27036,N_24835,N_26270);
xnor U27037 (N_27037,N_25576,N_25650);
nor U27038 (N_27038,N_26640,N_25794);
nor U27039 (N_27039,N_26900,N_26130);
nor U27040 (N_27040,N_26167,N_26149);
and U27041 (N_27041,N_25305,N_26815);
nand U27042 (N_27042,N_26925,N_24956);
xor U27043 (N_27043,N_26355,N_26003);
nor U27044 (N_27044,N_25026,N_25810);
and U27045 (N_27045,N_24512,N_25345);
nand U27046 (N_27046,N_26450,N_24049);
or U27047 (N_27047,N_24363,N_26277);
nor U27048 (N_27048,N_25762,N_25140);
and U27049 (N_27049,N_26874,N_26405);
xor U27050 (N_27050,N_25513,N_25227);
or U27051 (N_27051,N_24789,N_24286);
nor U27052 (N_27052,N_25441,N_26161);
nand U27053 (N_27053,N_24553,N_26986);
or U27054 (N_27054,N_25694,N_26120);
and U27055 (N_27055,N_26549,N_25914);
nand U27056 (N_27056,N_25021,N_25465);
nor U27057 (N_27057,N_24318,N_25056);
or U27058 (N_27058,N_24575,N_26220);
nand U27059 (N_27059,N_24807,N_26350);
and U27060 (N_27060,N_24222,N_24074);
and U27061 (N_27061,N_25809,N_26827);
nor U27062 (N_27062,N_26859,N_26704);
or U27063 (N_27063,N_24111,N_25937);
nand U27064 (N_27064,N_26197,N_24491);
nor U27065 (N_27065,N_24713,N_26399);
or U27066 (N_27066,N_24381,N_24569);
xnor U27067 (N_27067,N_24767,N_24482);
xor U27068 (N_27068,N_24913,N_24675);
nor U27069 (N_27069,N_24751,N_24324);
nor U27070 (N_27070,N_24211,N_25414);
nor U27071 (N_27071,N_26800,N_26666);
or U27072 (N_27072,N_25210,N_24106);
nand U27073 (N_27073,N_25898,N_25867);
or U27074 (N_27074,N_25198,N_24504);
nand U27075 (N_27075,N_24215,N_25631);
and U27076 (N_27076,N_24953,N_26433);
or U27077 (N_27077,N_26706,N_24694);
or U27078 (N_27078,N_25364,N_26464);
nand U27079 (N_27079,N_26119,N_24579);
and U27080 (N_27080,N_25878,N_24130);
or U27081 (N_27081,N_26692,N_24975);
or U27082 (N_27082,N_26232,N_24673);
nand U27083 (N_27083,N_26324,N_26626);
nor U27084 (N_27084,N_26345,N_25385);
xor U27085 (N_27085,N_24808,N_24972);
and U27086 (N_27086,N_24800,N_26979);
xor U27087 (N_27087,N_25469,N_26117);
nand U27088 (N_27088,N_24245,N_26871);
or U27089 (N_27089,N_25061,N_26691);
or U27090 (N_27090,N_24422,N_26305);
nor U27091 (N_27091,N_25107,N_25427);
or U27092 (N_27092,N_26516,N_24534);
and U27093 (N_27093,N_26506,N_26982);
and U27094 (N_27094,N_24583,N_26720);
and U27095 (N_27095,N_26375,N_24322);
or U27096 (N_27096,N_25037,N_25174);
and U27097 (N_27097,N_26022,N_26998);
xnor U27098 (N_27098,N_24388,N_24719);
or U27099 (N_27099,N_26632,N_24533);
xor U27100 (N_27100,N_25556,N_25235);
and U27101 (N_27101,N_25970,N_24804);
xor U27102 (N_27102,N_25119,N_25813);
or U27103 (N_27103,N_26140,N_25639);
and U27104 (N_27104,N_24763,N_26674);
and U27105 (N_27105,N_25742,N_24276);
or U27106 (N_27106,N_24416,N_26832);
nand U27107 (N_27107,N_26478,N_25952);
xor U27108 (N_27108,N_25184,N_24759);
or U27109 (N_27109,N_25442,N_25875);
xnor U27110 (N_27110,N_26207,N_24476);
nor U27111 (N_27111,N_25515,N_25429);
xor U27112 (N_27112,N_26202,N_24177);
or U27113 (N_27113,N_24964,N_24717);
nor U27114 (N_27114,N_26658,N_26384);
or U27115 (N_27115,N_24186,N_25504);
and U27116 (N_27116,N_24449,N_25409);
and U27117 (N_27117,N_25740,N_26089);
and U27118 (N_27118,N_24791,N_25873);
nor U27119 (N_27119,N_24384,N_24969);
and U27120 (N_27120,N_26802,N_24907);
xnor U27121 (N_27121,N_24587,N_26957);
nand U27122 (N_27122,N_25499,N_26079);
nand U27123 (N_27123,N_24656,N_24357);
and U27124 (N_27124,N_24951,N_26586);
or U27125 (N_27125,N_24586,N_24684);
nand U27126 (N_27126,N_24300,N_26583);
xor U27127 (N_27127,N_26990,N_24524);
and U27128 (N_27128,N_24678,N_24742);
or U27129 (N_27129,N_25579,N_24838);
nand U27130 (N_27130,N_25930,N_26053);
and U27131 (N_27131,N_26701,N_25488);
or U27132 (N_27132,N_25042,N_26145);
nor U27133 (N_27133,N_24520,N_24884);
nor U27134 (N_27134,N_24262,N_24366);
nor U27135 (N_27135,N_26535,N_25539);
or U27136 (N_27136,N_25361,N_24367);
and U27137 (N_27137,N_25017,N_24990);
or U27138 (N_27138,N_24264,N_24474);
xor U27139 (N_27139,N_25909,N_24383);
nand U27140 (N_27140,N_25980,N_24195);
nand U27141 (N_27141,N_24902,N_24644);
and U27142 (N_27142,N_25298,N_26058);
nand U27143 (N_27143,N_26109,N_26192);
and U27144 (N_27144,N_24825,N_26373);
or U27145 (N_27145,N_25926,N_25092);
xor U27146 (N_27146,N_24768,N_25991);
nor U27147 (N_27147,N_24549,N_24481);
xnor U27148 (N_27148,N_24319,N_24773);
or U27149 (N_27149,N_25992,N_26633);
nand U27150 (N_27150,N_25167,N_24034);
nand U27151 (N_27151,N_24395,N_24918);
and U27152 (N_27152,N_24680,N_26427);
nor U27153 (N_27153,N_25691,N_24589);
xor U27154 (N_27154,N_24976,N_26534);
and U27155 (N_27155,N_24858,N_25645);
or U27156 (N_27156,N_25240,N_25490);
nor U27157 (N_27157,N_24620,N_25132);
or U27158 (N_27158,N_24280,N_24496);
and U27159 (N_27159,N_24090,N_25053);
nand U27160 (N_27160,N_24303,N_26042);
xnor U27161 (N_27161,N_25517,N_24354);
nand U27162 (N_27162,N_26245,N_26411);
xor U27163 (N_27163,N_24250,N_25965);
nand U27164 (N_27164,N_26863,N_26764);
nor U27165 (N_27165,N_25201,N_26592);
nand U27166 (N_27166,N_25857,N_26974);
or U27167 (N_27167,N_24957,N_24545);
nor U27168 (N_27168,N_25014,N_25864);
xor U27169 (N_27169,N_25125,N_26178);
xor U27170 (N_27170,N_26498,N_25601);
or U27171 (N_27171,N_25322,N_25729);
xnor U27172 (N_27172,N_25756,N_25597);
nor U27173 (N_27173,N_25976,N_24997);
or U27174 (N_27174,N_25714,N_25336);
xor U27175 (N_27175,N_24919,N_24169);
nand U27176 (N_27176,N_24839,N_26223);
xor U27177 (N_27177,N_25447,N_26014);
and U27178 (N_27178,N_25654,N_24076);
and U27179 (N_27179,N_26654,N_25372);
nand U27180 (N_27180,N_26047,N_26241);
and U27181 (N_27181,N_25790,N_24755);
and U27182 (N_27182,N_25332,N_24636);
nor U27183 (N_27183,N_24993,N_25877);
nor U27184 (N_27184,N_25757,N_24448);
xnor U27185 (N_27185,N_25557,N_24100);
xnor U27186 (N_27186,N_25282,N_25846);
or U27187 (N_27187,N_26881,N_26699);
nor U27188 (N_27188,N_26960,N_24567);
nor U27189 (N_27189,N_25252,N_25560);
or U27190 (N_27190,N_26458,N_25010);
xor U27191 (N_27191,N_26422,N_24885);
and U27192 (N_27192,N_26712,N_26789);
xnor U27193 (N_27193,N_25885,N_24928);
nor U27194 (N_27194,N_26337,N_26934);
and U27195 (N_27195,N_25470,N_24723);
nand U27196 (N_27196,N_25329,N_26989);
and U27197 (N_27197,N_26273,N_25530);
or U27198 (N_27198,N_25972,N_24610);
nand U27199 (N_27199,N_25866,N_25544);
xnor U27200 (N_27200,N_25593,N_26737);
or U27201 (N_27201,N_24651,N_26573);
nand U27202 (N_27202,N_24653,N_25013);
or U27203 (N_27203,N_26641,N_24781);
nand U27204 (N_27204,N_25884,N_26814);
nor U27205 (N_27205,N_25031,N_25931);
nor U27206 (N_27206,N_25398,N_26939);
or U27207 (N_27207,N_25102,N_24469);
nor U27208 (N_27208,N_24382,N_26812);
nand U27209 (N_27209,N_24871,N_26486);
nand U27210 (N_27210,N_25718,N_24041);
nand U27211 (N_27211,N_26985,N_26770);
nand U27212 (N_27212,N_25253,N_25025);
nor U27213 (N_27213,N_25467,N_25719);
xor U27214 (N_27214,N_24862,N_24220);
and U27215 (N_27215,N_25892,N_25432);
and U27216 (N_27216,N_24240,N_24943);
or U27217 (N_27217,N_26447,N_24281);
xnor U27218 (N_27218,N_24502,N_24187);
nor U27219 (N_27219,N_24356,N_24135);
xor U27220 (N_27220,N_25443,N_26781);
nand U27221 (N_27221,N_25891,N_26166);
or U27222 (N_27222,N_24253,N_25495);
nand U27223 (N_27223,N_24278,N_25351);
nand U27224 (N_27224,N_26496,N_26276);
xor U27225 (N_27225,N_24470,N_25917);
and U27226 (N_27226,N_26956,N_26791);
nor U27227 (N_27227,N_26217,N_25573);
xnor U27228 (N_27228,N_26578,N_26211);
nor U27229 (N_27229,N_24981,N_24013);
nor U27230 (N_27230,N_24398,N_24299);
nand U27231 (N_27231,N_25549,N_26988);
or U27232 (N_27232,N_26279,N_26016);
xnor U27233 (N_27233,N_25977,N_25774);
nand U27234 (N_27234,N_24103,N_25642);
nor U27235 (N_27235,N_25095,N_25637);
or U27236 (N_27236,N_25510,N_25344);
and U27237 (N_27237,N_26258,N_25254);
and U27238 (N_27238,N_25094,N_24988);
and U27239 (N_27239,N_25060,N_24657);
or U27240 (N_27240,N_25307,N_24937);
and U27241 (N_27241,N_24691,N_26214);
or U27242 (N_27242,N_25151,N_26772);
and U27243 (N_27243,N_24766,N_26926);
or U27244 (N_27244,N_24002,N_26903);
and U27245 (N_27245,N_26436,N_24731);
xor U27246 (N_27246,N_25904,N_26456);
or U27247 (N_27247,N_26133,N_26707);
nor U27248 (N_27248,N_26541,N_24181);
and U27249 (N_27249,N_26967,N_25120);
or U27250 (N_27250,N_24308,N_26479);
nand U27251 (N_27251,N_24447,N_25889);
and U27252 (N_27252,N_26191,N_24554);
nor U27253 (N_27253,N_26181,N_26336);
and U27254 (N_27254,N_26520,N_26840);
and U27255 (N_27255,N_24389,N_24904);
or U27256 (N_27256,N_24999,N_24899);
or U27257 (N_27257,N_25540,N_25265);
xnor U27258 (N_27258,N_24908,N_25730);
and U27259 (N_27259,N_26308,N_26844);
xor U27260 (N_27260,N_24805,N_26895);
and U27261 (N_27261,N_26096,N_24754);
xor U27262 (N_27262,N_26210,N_24246);
nand U27263 (N_27263,N_24815,N_25039);
nor U27264 (N_27264,N_25697,N_25801);
xor U27265 (N_27265,N_24927,N_26554);
or U27266 (N_27266,N_24374,N_25956);
xnor U27267 (N_27267,N_26280,N_25401);
nor U27268 (N_27268,N_24349,N_24683);
nor U27269 (N_27269,N_25695,N_25478);
or U27270 (N_27270,N_26582,N_26567);
nor U27271 (N_27271,N_24306,N_26911);
or U27272 (N_27272,N_26103,N_25353);
xor U27273 (N_27273,N_26027,N_25365);
and U27274 (N_27274,N_25479,N_24600);
xnor U27275 (N_27275,N_25395,N_26804);
nor U27276 (N_27276,N_24778,N_24711);
xnor U27277 (N_27277,N_26910,N_25708);
and U27278 (N_27278,N_25362,N_25237);
xnor U27279 (N_27279,N_25958,N_25481);
nor U27280 (N_27280,N_26118,N_26327);
nor U27281 (N_27281,N_24637,N_25787);
or U27282 (N_27282,N_26050,N_24393);
nor U27283 (N_27283,N_26501,N_25966);
and U27284 (N_27284,N_26170,N_24727);
or U27285 (N_27285,N_26169,N_24216);
nor U27286 (N_27286,N_26719,N_24741);
nand U27287 (N_27287,N_25837,N_26543);
or U27288 (N_27288,N_24598,N_25131);
or U27289 (N_27289,N_25897,N_26460);
nand U27290 (N_27290,N_24340,N_25245);
nor U27291 (N_27291,N_26751,N_25734);
xor U27292 (N_27292,N_24551,N_25461);
or U27293 (N_27293,N_25653,N_25630);
and U27294 (N_27294,N_24980,N_24793);
nor U27295 (N_27295,N_25701,N_26524);
xor U27296 (N_27296,N_24328,N_26184);
or U27297 (N_27297,N_25200,N_25272);
or U27298 (N_27298,N_24992,N_25249);
xor U27299 (N_27299,N_25916,N_25072);
xnor U27300 (N_27300,N_24629,N_25584);
and U27301 (N_27301,N_25769,N_25887);
or U27302 (N_27302,N_24477,N_24313);
nor U27303 (N_27303,N_26285,N_24570);
nand U27304 (N_27304,N_26463,N_26841);
or U27305 (N_27305,N_24700,N_25699);
nor U27306 (N_27306,N_24233,N_25802);
nand U27307 (N_27307,N_24542,N_26610);
xnor U27308 (N_27308,N_24056,N_25005);
or U27309 (N_27309,N_25062,N_25389);
nand U27310 (N_27310,N_24952,N_24025);
nor U27311 (N_27311,N_24503,N_26205);
or U27312 (N_27312,N_26189,N_26051);
nand U27313 (N_27313,N_25647,N_26935);
xor U27314 (N_27314,N_25503,N_26835);
and U27315 (N_27315,N_26830,N_25070);
or U27316 (N_27316,N_24312,N_25301);
nor U27317 (N_27317,N_25686,N_26745);
nor U27318 (N_27318,N_24059,N_24495);
nand U27319 (N_27319,N_26519,N_26522);
or U27320 (N_27320,N_25759,N_24922);
or U27321 (N_27321,N_24267,N_24406);
or U27322 (N_27322,N_26010,N_25177);
and U27323 (N_27323,N_25360,N_24429);
xnor U27324 (N_27324,N_25143,N_25920);
nor U27325 (N_27325,N_24046,N_25948);
and U27326 (N_27326,N_24027,N_24175);
nor U27327 (N_27327,N_26465,N_26670);
and U27328 (N_27328,N_26158,N_24962);
and U27329 (N_27329,N_26787,N_25894);
nor U27330 (N_27330,N_24627,N_26099);
nor U27331 (N_27331,N_25633,N_24439);
and U27332 (N_27332,N_24794,N_25933);
xor U27333 (N_27333,N_25999,N_24369);
nor U27334 (N_27334,N_26195,N_24911);
nand U27335 (N_27335,N_25388,N_25725);
nand U27336 (N_27336,N_24184,N_24061);
xnor U27337 (N_27337,N_25773,N_25420);
xor U27338 (N_27338,N_26819,N_24564);
nor U27339 (N_27339,N_24402,N_26796);
and U27340 (N_27340,N_25314,N_24084);
and U27341 (N_27341,N_25196,N_24213);
and U27342 (N_27342,N_25793,N_25747);
and U27343 (N_27343,N_24415,N_26663);
nor U27344 (N_27344,N_25994,N_25772);
nand U27345 (N_27345,N_24836,N_24133);
and U27346 (N_27346,N_24334,N_24841);
nor U27347 (N_27347,N_24715,N_25962);
nand U27348 (N_27348,N_24436,N_24378);
and U27349 (N_27349,N_26453,N_26061);
and U27350 (N_27350,N_24803,N_25460);
nand U27351 (N_27351,N_26514,N_26239);
nand U27352 (N_27352,N_25007,N_24151);
xor U27353 (N_27353,N_25571,N_25840);
nand U27354 (N_27354,N_26817,N_25792);
nand U27355 (N_27355,N_25274,N_26024);
xnor U27356 (N_27356,N_24613,N_25279);
or U27357 (N_27357,N_25852,N_24621);
nor U27358 (N_27358,N_24706,N_24182);
xor U27359 (N_27359,N_25752,N_25375);
and U27360 (N_27360,N_25074,N_26993);
and U27361 (N_27361,N_26927,N_25055);
nor U27362 (N_27362,N_24769,N_24050);
nand U27363 (N_27363,N_24287,N_24652);
and U27364 (N_27364,N_24882,N_24265);
nand U27365 (N_27365,N_25160,N_26698);
or U27366 (N_27366,N_25812,N_24110);
xor U27367 (N_27367,N_24386,N_26898);
xnor U27368 (N_27368,N_26365,N_25331);
nor U27369 (N_27369,N_24592,N_25625);
and U27370 (N_27370,N_24757,N_25346);
or U27371 (N_27371,N_25811,N_26397);
and U27372 (N_27372,N_25303,N_25258);
nand U27373 (N_27373,N_24903,N_26293);
nand U27374 (N_27374,N_25324,N_24289);
xnor U27375 (N_27375,N_26015,N_25266);
xnor U27376 (N_27376,N_26380,N_24284);
nand U27377 (N_27377,N_25671,N_25121);
or U27378 (N_27378,N_26052,N_24126);
or U27379 (N_27379,N_24905,N_26937);
nand U27380 (N_27380,N_24607,N_25673);
or U27381 (N_27381,N_25596,N_25393);
or U27382 (N_27382,N_25555,N_26401);
nor U27383 (N_27383,N_26304,N_25417);
and U27384 (N_27384,N_26563,N_25700);
xnor U27385 (N_27385,N_24792,N_24261);
or U27386 (N_27386,N_25180,N_24647);
nor U27387 (N_27387,N_24221,N_24880);
or U27388 (N_27388,N_26556,N_25286);
nand U27389 (N_27389,N_26338,N_24007);
or U27390 (N_27390,N_25624,N_26424);
and U27391 (N_27391,N_26750,N_26282);
and U27392 (N_27392,N_26150,N_26389);
and U27393 (N_27393,N_24405,N_24115);
nand U27394 (N_27394,N_24774,N_26660);
xnor U27395 (N_27395,N_25538,N_24206);
nor U27396 (N_27396,N_25040,N_24896);
or U27397 (N_27397,N_24643,N_25384);
and U27398 (N_27398,N_26264,N_26063);
xnor U27399 (N_27399,N_26421,N_26951);
xnor U27400 (N_27400,N_26742,N_24628);
or U27401 (N_27401,N_26477,N_26652);
xnor U27402 (N_27402,N_24557,N_26066);
nand U27403 (N_27403,N_24698,N_25494);
nand U27404 (N_27404,N_25776,N_24174);
and U27405 (N_27405,N_24305,N_24568);
nor U27406 (N_27406,N_24832,N_26488);
and U27407 (N_27407,N_25739,N_24822);
xor U27408 (N_27408,N_25862,N_25320);
or U27409 (N_27409,N_25951,N_26919);
xor U27410 (N_27410,N_26417,N_25064);
xnor U27411 (N_27411,N_26574,N_24736);
nor U27412 (N_27412,N_24492,N_26952);
nor U27413 (N_27413,N_24664,N_24204);
nor U27414 (N_27414,N_25750,N_24234);
xor U27415 (N_27415,N_25230,N_26286);
nand U27416 (N_27416,N_26560,N_24812);
xor U27417 (N_27417,N_24301,N_26624);
nand U27418 (N_27418,N_25374,N_25041);
or U27419 (N_27419,N_26728,N_25907);
nor U27420 (N_27420,N_24501,N_24087);
and U27421 (N_27421,N_26295,N_24671);
nand U27422 (N_27422,N_25083,N_26748);
and U27423 (N_27423,N_26598,N_26201);
or U27424 (N_27424,N_24722,N_25103);
nand U27425 (N_27425,N_25439,N_26693);
xor U27426 (N_27426,N_25118,N_26267);
nor U27427 (N_27427,N_25693,N_25921);
xor U27428 (N_27428,N_26568,N_25246);
or U27429 (N_27429,N_26126,N_24965);
xor U27430 (N_27430,N_25682,N_24817);
nand U27431 (N_27431,N_24977,N_25339);
and U27432 (N_27432,N_24856,N_24833);
and U27433 (N_27433,N_25674,N_24726);
nand U27434 (N_27434,N_25832,N_25638);
and U27435 (N_27435,N_25391,N_26713);
nor U27436 (N_27436,N_24693,N_24931);
or U27437 (N_27437,N_24982,N_25194);
nand U27438 (N_27438,N_24071,N_26495);
or U27439 (N_27439,N_26576,N_24940);
xnor U27440 (N_27440,N_24200,N_24085);
or U27441 (N_27441,N_24323,N_26087);
nand U27442 (N_27442,N_26984,N_26138);
xor U27443 (N_27443,N_25532,N_25438);
nor U27444 (N_27444,N_26879,N_24619);
and U27445 (N_27445,N_26437,N_24310);
xnor U27446 (N_27446,N_26132,N_26648);
nor U27447 (N_27447,N_25436,N_25715);
nor U27448 (N_27448,N_24971,N_26946);
xnor U27449 (N_27449,N_25173,N_24454);
nor U27450 (N_27450,N_26733,N_25164);
or U27451 (N_27451,N_24617,N_26932);
nand U27452 (N_27452,N_24597,N_25081);
and U27453 (N_27453,N_25090,N_24738);
or U27454 (N_27454,N_24946,N_25520);
nor U27455 (N_27455,N_26376,N_24249);
xnor U27456 (N_27456,N_25968,N_24037);
nor U27457 (N_27457,N_25248,N_26129);
nor U27458 (N_27458,N_24942,N_25291);
xor U27459 (N_27459,N_25692,N_26596);
xor U27460 (N_27460,N_25942,N_25285);
xor U27461 (N_27461,N_25574,N_26512);
nand U27462 (N_27462,N_25868,N_26313);
and U27463 (N_27463,N_25241,N_26729);
nand U27464 (N_27464,N_24075,N_26559);
xnor U27465 (N_27465,N_24418,N_25676);
and U27466 (N_27466,N_24121,N_25034);
nor U27467 (N_27467,N_25284,N_26155);
nand U27468 (N_27468,N_25707,N_26601);
nand U27469 (N_27469,N_24933,N_24983);
and U27470 (N_27470,N_24162,N_24089);
or U27471 (N_27471,N_25987,N_25830);
xnor U27472 (N_27472,N_26271,N_24232);
xor U27473 (N_27473,N_24869,N_26775);
and U27474 (N_27474,N_24332,N_26395);
nor U27475 (N_27475,N_24536,N_24887);
or U27476 (N_27476,N_25611,N_26144);
and U27477 (N_27477,N_25943,N_26480);
nand U27478 (N_27478,N_24463,N_26839);
nor U27479 (N_27479,N_24662,N_24252);
nor U27480 (N_27480,N_26386,N_25233);
or U27481 (N_27481,N_26758,N_25150);
and U27482 (N_27482,N_26941,N_26351);
nand U27483 (N_27483,N_25704,N_25100);
nor U27484 (N_27484,N_24909,N_24102);
nor U27485 (N_27485,N_25957,N_25588);
and U27486 (N_27486,N_25870,N_25507);
or U27487 (N_27487,N_24954,N_26084);
and U27488 (N_27488,N_25226,N_26690);
nor U27489 (N_27489,N_24779,N_25455);
nor U27490 (N_27490,N_25640,N_24578);
xnor U27491 (N_27491,N_26403,N_25908);
and U27492 (N_27492,N_26906,N_24203);
and U27493 (N_27493,N_24523,N_26617);
nor U27494 (N_27494,N_24006,N_26646);
or U27495 (N_27495,N_25257,N_24104);
nand U27496 (N_27496,N_26807,N_24042);
nand U27497 (N_27497,N_26888,N_26423);
and U27498 (N_27498,N_24527,N_26216);
nand U27499 (N_27499,N_24556,N_25424);
nor U27500 (N_27500,N_24588,N_24134);
nor U27501 (N_27501,N_24263,N_25903);
and U27502 (N_27502,N_25146,N_24202);
or U27503 (N_27503,N_25101,N_25768);
and U27504 (N_27504,N_25416,N_25359);
or U27505 (N_27505,N_25403,N_24044);
xnor U27506 (N_27506,N_25263,N_26928);
and U27507 (N_27507,N_26182,N_24867);
nand U27508 (N_27508,N_26838,N_26208);
or U27509 (N_27509,N_26920,N_25978);
and U27510 (N_27510,N_24420,N_24165);
or U27511 (N_27511,N_24770,N_24337);
nor U27512 (N_27512,N_26428,N_24031);
xnor U27513 (N_27513,N_26072,N_25981);
and U27514 (N_27514,N_26174,N_26025);
nor U27515 (N_27515,N_25002,N_25913);
nor U27516 (N_27516,N_25526,N_24499);
nand U27517 (N_27517,N_26860,N_25924);
nand U27518 (N_27518,N_26709,N_26101);
and U27519 (N_27519,N_24820,N_24963);
nor U27520 (N_27520,N_26569,N_26873);
nand U27521 (N_27521,N_25860,N_25592);
xor U27522 (N_27522,N_25755,N_25437);
and U27523 (N_27523,N_24543,N_24047);
xnor U27524 (N_27524,N_24236,N_25749);
or U27525 (N_27525,N_26756,N_25669);
nand U27526 (N_27526,N_26526,N_25415);
nand U27527 (N_27527,N_24599,N_25554);
or U27528 (N_27528,N_26971,N_26857);
nor U27529 (N_27529,N_26315,N_26968);
or U27530 (N_27530,N_26850,N_24168);
and U27531 (N_27531,N_24444,N_26039);
nand U27532 (N_27532,N_24430,N_26121);
nor U27533 (N_27533,N_25032,N_26600);
and U27534 (N_27534,N_24414,N_24178);
xor U27535 (N_27535,N_26431,N_25829);
nor U27536 (N_27536,N_24924,N_26222);
and U27537 (N_27537,N_26322,N_24417);
nand U27538 (N_27538,N_25463,N_26981);
xnor U27539 (N_27539,N_24073,N_26425);
and U27540 (N_27540,N_25606,N_26092);
nor U27541 (N_27541,N_24648,N_24734);
and U27542 (N_27542,N_26100,N_25019);
or U27543 (N_27543,N_24272,N_26969);
nand U27544 (N_27544,N_26317,N_26959);
or U27545 (N_27545,N_24452,N_25452);
nand U27546 (N_27546,N_25142,N_24573);
and U27547 (N_27547,N_25216,N_25281);
xnor U27548 (N_27548,N_26198,N_24266);
xnor U27549 (N_27549,N_26876,N_25097);
and U27550 (N_27550,N_26366,N_24285);
xnor U27551 (N_27551,N_25197,N_26912);
and U27552 (N_27552,N_25628,N_24091);
or U27553 (N_27553,N_26485,N_24164);
nand U27554 (N_27554,N_26246,N_26330);
xor U27555 (N_27555,N_25543,N_25670);
and U27556 (N_27556,N_24844,N_25577);
nor U27557 (N_27557,N_26771,N_25569);
xnor U27558 (N_27558,N_24784,N_24748);
xor U27559 (N_27559,N_26203,N_24852);
nor U27560 (N_27560,N_26782,N_26339);
nand U27561 (N_27561,N_25893,N_24538);
nor U27562 (N_27562,N_25352,N_26344);
nand U27563 (N_27563,N_24786,N_26153);
nor U27564 (N_27564,N_25564,N_26383);
nor U27565 (N_27565,N_24403,N_24912);
nor U27566 (N_27566,N_24860,N_25199);
nor U27567 (N_27567,N_25761,N_24521);
and U27568 (N_27568,N_26272,N_26943);
or U27569 (N_27569,N_25890,N_25827);
nand U27570 (N_27570,N_26602,N_25482);
xnor U27571 (N_27571,N_25220,N_25928);
nand U27572 (N_27572,N_25484,N_24331);
and U27573 (N_27573,N_26635,N_24478);
nand U27574 (N_27574,N_24193,N_26502);
or U27575 (N_27575,N_24910,N_26562);
and U27576 (N_27576,N_26075,N_25551);
xor U27577 (N_27577,N_25480,N_26749);
or U27578 (N_27578,N_25168,N_26595);
nand U27579 (N_27579,N_26009,N_26049);
and U27580 (N_27580,N_26725,N_25089);
or U27581 (N_27581,N_26518,N_26627);
nor U27582 (N_27582,N_26767,N_25008);
and U27583 (N_27583,N_26128,N_25833);
or U27584 (N_27584,N_26080,N_24535);
nor U27585 (N_27585,N_25516,N_24144);
xnor U27586 (N_27586,N_25067,N_25371);
or U27587 (N_27587,N_24487,N_24433);
xor U27588 (N_27588,N_26259,N_24304);
or U27589 (N_27589,N_25161,N_24605);
or U27590 (N_27590,N_24847,N_26176);
nand U27591 (N_27591,N_25675,N_24294);
and U27592 (N_27592,N_25000,N_25251);
xnor U27593 (N_27593,N_24532,N_24681);
nand U27594 (N_27594,N_24205,N_24488);
or U27595 (N_27595,N_26157,N_26675);
xor U27596 (N_27596,N_24935,N_25155);
xor U27597 (N_27597,N_25182,N_26580);
xnor U27598 (N_27598,N_26552,N_26151);
xor U27599 (N_27599,N_26257,N_26146);
or U27600 (N_27600,N_26848,N_24373);
nor U27601 (N_27601,N_24517,N_25572);
xnor U27602 (N_27602,N_26513,N_24048);
nand U27603 (N_27603,N_25679,N_24650);
nor U27604 (N_27604,N_26855,N_26160);
nand U27605 (N_27605,N_25458,N_25152);
nand U27606 (N_27606,N_25086,N_24485);
nand U27607 (N_27607,N_24525,N_24137);
or U27608 (N_27608,N_24079,N_26135);
and U27609 (N_27609,N_25954,N_25687);
xor U27610 (N_27610,N_25413,N_26352);
nand U27611 (N_27611,N_24270,N_26183);
nand U27612 (N_27612,N_24777,N_24358);
and U27613 (N_27613,N_25133,N_24875);
nand U27614 (N_27614,N_26179,N_24054);
or U27615 (N_27615,N_24167,N_26228);
nor U27616 (N_27616,N_24923,N_26064);
nor U27617 (N_27617,N_26468,N_25190);
nand U27618 (N_27618,N_24413,N_24020);
and U27619 (N_27619,N_24690,N_26829);
nand U27620 (N_27620,N_26736,N_24003);
xnor U27621 (N_27621,N_26115,N_25844);
nand U27622 (N_27622,N_26538,N_26593);
nand U27623 (N_27623,N_26816,N_24631);
nand U27624 (N_27624,N_26372,N_25825);
or U27625 (N_27625,N_24017,N_25287);
nor U27626 (N_27626,N_24368,N_25386);
nor U27627 (N_27627,N_26613,N_25971);
nand U27628 (N_27628,N_25052,N_25188);
and U27629 (N_27629,N_26091,N_25404);
nand U27630 (N_27630,N_25607,N_26426);
xor U27631 (N_27631,N_24709,N_26639);
and U27632 (N_27632,N_25434,N_24064);
xor U27633 (N_27633,N_26950,N_24850);
and U27634 (N_27634,N_24026,N_26212);
and U27635 (N_27635,N_26676,N_24890);
or U27636 (N_27636,N_24594,N_25453);
nor U27637 (N_27637,N_24258,N_24341);
xnor U27638 (N_27638,N_26976,N_24223);
xor U27639 (N_27639,N_26114,N_25528);
nor U27640 (N_27640,N_24883,N_24776);
xnor U27641 (N_27641,N_26904,N_24859);
nand U27642 (N_27642,N_25422,N_25029);
nor U27643 (N_27643,N_24707,N_24494);
nor U27644 (N_27644,N_24926,N_25221);
nor U27645 (N_27645,N_24625,N_26021);
and U27646 (N_27646,N_26219,N_26321);
or U27647 (N_27647,N_24490,N_26415);
nor U27648 (N_27648,N_26493,N_24771);
nand U27649 (N_27649,N_24895,N_26788);
and U27650 (N_27650,N_24347,N_24959);
and U27651 (N_27651,N_25678,N_26685);
and U27652 (N_27652,N_25491,N_26869);
xnor U27653 (N_27653,N_26306,N_24172);
or U27654 (N_27654,N_24515,N_24889);
nor U27655 (N_27655,N_25475,N_24455);
or U27656 (N_27656,N_26899,N_25057);
nor U27657 (N_27657,N_26999,N_24375);
nand U27658 (N_27658,N_24518,N_26766);
nor U27659 (N_27659,N_25936,N_24798);
nor U27660 (N_27660,N_26056,N_25319);
xor U27661 (N_27661,N_24122,N_24898);
nor U27662 (N_27662,N_25895,N_25855);
or U27663 (N_27663,N_24288,N_25511);
nor U27664 (N_27664,N_25514,N_24623);
nand U27665 (N_27665,N_24427,N_26227);
nor U27666 (N_27666,N_24855,N_24466);
or U27667 (N_27667,N_25944,N_25583);
nand U27668 (N_27668,N_25836,N_26283);
nor U27669 (N_27669,N_26284,N_25421);
or U27670 (N_27670,N_24611,N_24635);
or U27671 (N_27671,N_25466,N_26067);
nor U27672 (N_27672,N_24699,N_26269);
and U27673 (N_27673,N_25407,N_24780);
xnor U27674 (N_27674,N_25798,N_24752);
or U27675 (N_27675,N_25938,N_24155);
nor U27676 (N_27676,N_26379,N_25586);
xor U27677 (N_27677,N_25553,N_25341);
nand U27678 (N_27678,N_26448,N_24066);
or U27679 (N_27679,N_26082,N_26604);
and U27680 (N_27680,N_26499,N_24446);
xnor U27681 (N_27681,N_25289,N_26889);
or U27682 (N_27682,N_25799,N_25073);
or U27683 (N_27683,N_26172,N_24376);
nor U27684 (N_27684,N_26851,N_24029);
and U27685 (N_27685,N_26882,N_24733);
and U27686 (N_27686,N_25390,N_26555);
or U27687 (N_27687,N_24001,N_24936);
and U27688 (N_27688,N_25874,N_24385);
or U27689 (N_27689,N_25911,N_24109);
and U27690 (N_27690,N_24019,N_24326);
xnor U27691 (N_27691,N_24978,N_24051);
xnor U27692 (N_27692,N_26497,N_24677);
nor U27693 (N_27693,N_25213,N_26996);
and U27694 (N_27694,N_26312,N_25474);
nand U27695 (N_27695,N_24058,N_24785);
nor U27696 (N_27696,N_24513,N_26972);
nand U27697 (N_27697,N_25815,N_25736);
xnor U27698 (N_27698,N_25807,N_25295);
xor U27699 (N_27699,N_24330,N_25049);
nor U27700 (N_27700,N_24821,N_25030);
and U27701 (N_27701,N_24566,N_25912);
nor U27702 (N_27702,N_24493,N_25419);
xnor U27703 (N_27703,N_26193,N_24148);
nor U27704 (N_27704,N_24425,N_26980);
or U27705 (N_27705,N_24131,N_24641);
or U27706 (N_27706,N_25412,N_26244);
or U27707 (N_27707,N_24317,N_26102);
nor U27708 (N_27708,N_25983,N_25854);
nand U27709 (N_27709,N_24189,N_24140);
and U27710 (N_27710,N_25751,N_25099);
xnor U27711 (N_27711,N_26341,N_26856);
xnor U27712 (N_27712,N_25082,N_25264);
xnor U27713 (N_27713,N_26462,N_25006);
and U27714 (N_27714,N_25716,N_26074);
nand U27715 (N_27715,N_26571,N_26681);
or U27716 (N_27716,N_24765,N_24740);
nand U27717 (N_27717,N_24560,N_26011);
nand U27718 (N_27718,N_26715,N_26921);
and U27719 (N_27719,N_26962,N_24509);
and U27720 (N_27720,N_25603,N_26786);
xor U27721 (N_27721,N_24892,N_26162);
nand U27722 (N_27722,N_26892,N_26215);
xor U27723 (N_27723,N_26509,N_26615);
or U27724 (N_27724,N_24387,N_25268);
or U27725 (N_27725,N_24445,N_26474);
and U27726 (N_27726,N_24606,N_26607);
xnor U27727 (N_27727,N_26071,N_26300);
nand U27728 (N_27728,N_25111,N_25366);
or U27729 (N_27729,N_25218,N_26533);
and U27730 (N_27730,N_26185,N_25805);
and U27731 (N_27731,N_25986,N_24925);
or U27732 (N_27732,N_24424,N_24540);
and U27733 (N_27733,N_25448,N_25781);
or U27734 (N_27734,N_26008,N_25929);
nand U27735 (N_27735,N_24702,N_24823);
or U27736 (N_27736,N_24435,N_24298);
nand U27737 (N_27737,N_24149,N_24329);
and U27738 (N_27738,N_26249,N_24949);
nor U27739 (N_27739,N_24008,N_24170);
and U27740 (N_27740,N_26234,N_24516);
nor U27741 (N_27741,N_26095,N_26643);
xnor U27742 (N_27742,N_26340,N_26581);
and U27743 (N_27743,N_24746,N_25963);
and U27744 (N_27744,N_25778,N_26525);
nand U27745 (N_27745,N_26890,N_26429);
xnor U27746 (N_27746,N_25735,N_24921);
and U27747 (N_27747,N_26187,N_25489);
and U27748 (N_27748,N_26537,N_24271);
and U27749 (N_27749,N_24840,N_24714);
xor U27750 (N_27750,N_24199,N_25559);
and U27751 (N_27751,N_26634,N_26550);
or U27752 (N_27752,N_26472,N_24945);
or U27753 (N_27753,N_24582,N_26507);
nor U27754 (N_27754,N_24580,N_24099);
or U27755 (N_27755,N_25524,N_26877);
or U27756 (N_27756,N_26168,N_26741);
xor U27757 (N_27757,N_26356,N_24442);
nand U27758 (N_27758,N_24257,N_24687);
and U27759 (N_27759,N_25789,N_26029);
nand U27760 (N_27760,N_26069,N_25737);
nand U27761 (N_27761,N_25047,N_24361);
nand U27762 (N_27762,N_24309,N_24450);
and U27763 (N_27763,N_24014,N_26759);
and U27764 (N_27764,N_24639,N_26290);
xnor U27765 (N_27765,N_24666,N_24114);
nor U27766 (N_27766,N_26018,N_26746);
nand U27767 (N_27767,N_26662,N_25162);
and U27768 (N_27768,N_24201,N_26371);
and U27769 (N_27769,N_26252,N_25299);
nand U27770 (N_27770,N_24724,N_25519);
or U27771 (N_27771,N_26459,N_25428);
nor U27772 (N_27772,N_26449,N_26298);
or U27773 (N_27773,N_25387,N_25657);
and U27774 (N_27774,N_24826,N_25178);
xnor U27775 (N_27775,N_24467,N_25450);
nand U27776 (N_27776,N_24660,N_26037);
and U27777 (N_27777,N_24244,N_26301);
nand U27778 (N_27778,N_26716,N_25501);
nand U27779 (N_27779,N_24998,N_26686);
nor U27780 (N_27780,N_25804,N_25535);
or U27781 (N_27781,N_26046,N_24546);
and U27782 (N_27782,N_26026,N_24679);
xor U27783 (N_27783,N_25300,N_26137);
nor U27784 (N_27784,N_25626,N_24194);
and U27785 (N_27785,N_25293,N_24739);
xnor U27786 (N_27786,N_26467,N_24283);
nor U27787 (N_27787,N_24505,N_24604);
and U27788 (N_27788,N_25896,N_25702);
and U27789 (N_27789,N_25242,N_24343);
or U27790 (N_27790,N_24400,N_26661);
or U27791 (N_27791,N_25821,N_26164);
nor U27792 (N_27792,N_25974,N_24077);
xor U27793 (N_27793,N_24072,N_24802);
xor U27794 (N_27794,N_26924,N_25239);
nand U27795 (N_27795,N_26329,N_25782);
nor U27796 (N_27796,N_25456,N_24248);
or U27797 (N_27797,N_26445,N_26826);
nand U27798 (N_27798,N_24851,N_25045);
nor U27799 (N_27799,N_24128,N_26695);
nor U27800 (N_27800,N_25468,N_26945);
nor U27801 (N_27801,N_26093,N_26997);
nor U27802 (N_27802,N_24161,N_25995);
nand U27803 (N_27803,N_26868,N_25785);
nand U27804 (N_27804,N_25157,N_26905);
or U27805 (N_27805,N_25613,N_24480);
nand U27806 (N_27806,N_25932,N_24934);
nand U27807 (N_27807,N_24735,N_24831);
nand U27808 (N_27808,N_24848,N_25236);
and U27809 (N_27809,N_24878,N_26689);
nand U27810 (N_27810,N_26846,N_26152);
nand U27811 (N_27811,N_24682,N_24316);
nor U27812 (N_27812,N_26795,N_25947);
nand U27813 (N_27813,N_24854,N_26048);
nor U27814 (N_27814,N_24721,N_25509);
or U27815 (N_27815,N_25496,N_24642);
or U27816 (N_27816,N_26907,N_26457);
xor U27817 (N_27817,N_26887,N_26253);
and U27818 (N_27818,N_24255,N_24514);
nor U27819 (N_27819,N_24247,N_24379);
nand U27820 (N_27820,N_26041,N_26803);
and U27821 (N_27821,N_26319,N_26708);
xor U27822 (N_27822,N_24086,N_24336);
xor U27823 (N_27823,N_25990,N_25536);
nand U27824 (N_27824,N_26579,N_26206);
nor U27825 (N_27825,N_24431,N_26975);
xor U27826 (N_27826,N_25123,N_26531);
and U27827 (N_27827,N_26836,N_24229);
and U27828 (N_27828,N_26209,N_26310);
nor U27829 (N_27829,N_26113,N_25663);
xnor U27830 (N_27830,N_24783,N_26494);
and U27831 (N_27831,N_24461,N_25270);
nor U27832 (N_27832,N_25834,N_25065);
or U27833 (N_27833,N_26978,N_26631);
and U27834 (N_27834,N_25605,N_25280);
nor U27835 (N_27835,N_25195,N_26853);
nand U27836 (N_27836,N_25668,N_26994);
or U27837 (N_27837,N_25338,N_26461);
and U27838 (N_27838,N_25753,N_25582);
nor U27839 (N_27839,N_24083,N_26302);
xor U27840 (N_27840,N_24471,N_24670);
and U27841 (N_27841,N_24725,N_24302);
xor U27842 (N_27842,N_25084,N_24320);
and U27843 (N_27843,N_26045,N_26299);
nand U27844 (N_27844,N_26682,N_24401);
nand U27845 (N_27845,N_26572,N_25138);
or U27846 (N_27846,N_25208,N_26636);
and U27847 (N_27847,N_26618,N_26558);
nor U27848 (N_27848,N_24069,N_26398);
and U27849 (N_27849,N_26085,N_25408);
or U27850 (N_27850,N_24608,N_24750);
and U27851 (N_27851,N_26915,N_26947);
or U27852 (N_27852,N_24021,N_25011);
or U27853 (N_27853,N_25325,N_24489);
xnor U27854 (N_27854,N_25015,N_25440);
xor U27855 (N_27855,N_24274,N_25229);
nor U27856 (N_27856,N_25996,N_25728);
xor U27857 (N_27857,N_25269,N_26703);
or U27858 (N_27858,N_25435,N_26619);
nor U27859 (N_27859,N_25215,N_26492);
xnor U27860 (N_27860,N_26668,N_25158);
nand U27861 (N_27861,N_25283,N_26801);
or U27862 (N_27862,N_24873,N_24160);
xor U27863 (N_27863,N_25059,N_26291);
nand U27864 (N_27864,N_24879,N_26400);
nand U27865 (N_27865,N_24018,N_24390);
nand U27866 (N_27866,N_26238,N_25845);
xor U27867 (N_27867,N_26747,N_25627);
nand U27868 (N_27868,N_24009,N_24897);
nand U27869 (N_27869,N_24365,N_26256);
nor U27870 (N_27870,N_26861,N_24372);
and U27871 (N_27871,N_26303,N_24849);
nand U27872 (N_27872,N_26842,N_25882);
nor U27873 (N_27873,N_25363,N_25116);
nand U27874 (N_27874,N_25426,N_24602);
xnor U27875 (N_27875,N_26837,N_24166);
nor U27876 (N_27876,N_26778,N_25652);
xor U27877 (N_27877,N_24377,N_25078);
nor U27878 (N_27878,N_25122,N_25445);
and U27879 (N_27879,N_26028,N_24015);
and U27880 (N_27880,N_25717,N_25054);
xor U27881 (N_27881,N_26139,N_26240);
or U27882 (N_27882,N_24230,N_26722);
nor U27883 (N_27883,N_24295,N_25327);
or U27884 (N_27884,N_26281,N_25959);
xor U27885 (N_27885,N_24624,N_25425);
and U27886 (N_27886,N_25343,N_24985);
nand U27887 (N_27887,N_24947,N_26862);
xor U27888 (N_27888,N_24581,N_26287);
and U27889 (N_27889,N_24915,N_26954);
nand U27890 (N_27890,N_26588,N_26515);
nor U27891 (N_27891,N_25727,N_25087);
xor U27892 (N_27892,N_25849,N_26551);
or U27893 (N_27893,N_24237,N_25795);
xor U27894 (N_27894,N_24828,N_25508);
xor U27895 (N_27895,N_24024,N_24097);
and U27896 (N_27896,N_26831,N_25879);
nand U27897 (N_27897,N_25368,N_26944);
nand U27898 (N_27898,N_26235,N_26843);
or U27899 (N_27899,N_25910,N_25159);
nand U27900 (N_27900,N_25317,N_24325);
nand U27901 (N_27901,N_26584,N_25126);
xnor U27902 (N_27902,N_26723,N_25193);
nand U27903 (N_27903,N_24584,N_24227);
or U27904 (N_27904,N_25212,N_25109);
xnor U27905 (N_27905,N_26823,N_26653);
nor U27906 (N_27906,N_24095,N_25886);
xnor U27907 (N_27907,N_25711,N_26369);
or U27908 (N_27908,N_26597,N_24809);
and U27909 (N_27909,N_26872,N_24101);
nor U27910 (N_27910,N_26570,N_26032);
nand U27911 (N_27911,N_26326,N_26940);
nand U27912 (N_27912,N_25745,N_24327);
and U27913 (N_27913,N_25457,N_26896);
nand U27914 (N_27914,N_26734,N_24371);
xor U27915 (N_27915,N_26483,N_24364);
and U27916 (N_27916,N_24930,N_26385);
xnor U27917 (N_27917,N_25713,N_25915);
nand U27918 (N_27918,N_25367,N_25326);
and U27919 (N_27919,N_24440,N_25527);
or U27920 (N_27920,N_25863,N_25839);
nor U27921 (N_27921,N_24728,N_24254);
and U27922 (N_27922,N_24173,N_24348);
xnor U27923 (N_27923,N_26517,N_26625);
nand U27924 (N_27924,N_26236,N_26738);
xnor U27925 (N_27925,N_25400,N_25681);
nor U27926 (N_27926,N_25883,N_26504);
xor U27927 (N_27927,N_25587,N_24117);
nor U27928 (N_27928,N_24342,N_24035);
and U27929 (N_27929,N_24321,N_26665);
or U27930 (N_27930,N_26642,N_26473);
or U27931 (N_27931,N_25826,N_24269);
nor U27932 (N_27932,N_25348,N_26866);
xor U27933 (N_27933,N_26481,N_24955);
or U27934 (N_27934,N_26755,N_25192);
nand U27935 (N_27935,N_25934,N_25741);
xor U27936 (N_27936,N_24139,N_26394);
or U27937 (N_27937,N_25552,N_26491);
xnor U27938 (N_27938,N_25373,N_24562);
nand U27939 (N_27939,N_26822,N_25558);
xnor U27940 (N_27940,N_26001,N_24591);
and U27941 (N_27941,N_25204,N_24796);
nand U27942 (N_27942,N_24544,N_25232);
xnor U27943 (N_27943,N_26732,N_26740);
xor U27944 (N_27944,N_26225,N_24659);
nand U27945 (N_27945,N_26254,N_25383);
and U27946 (N_27946,N_26333,N_26098);
and U27947 (N_27947,N_26702,N_26724);
nor U27948 (N_27948,N_26163,N_25777);
or U27949 (N_27949,N_25817,N_25823);
nor U27950 (N_27950,N_24437,N_26154);
xor U27951 (N_27951,N_26768,N_26797);
nor U27952 (N_27952,N_24893,N_26466);
xnor U27953 (N_27953,N_26331,N_25405);
and U27954 (N_27954,N_24472,N_24338);
nand U27955 (N_27955,N_26004,N_25337);
nand U27956 (N_27956,N_25271,N_26930);
and U27957 (N_27957,N_26171,N_24335);
xnor U27958 (N_27958,N_24843,N_25397);
or U27959 (N_27959,N_25620,N_25720);
nor U27960 (N_27960,N_26034,N_26783);
and U27961 (N_27961,N_26849,N_26487);
and U27962 (N_27962,N_24209,N_26353);
xnor U27963 (N_27963,N_25418,N_24756);
or U27964 (N_27964,N_24190,N_24507);
xor U27965 (N_27965,N_26361,N_26710);
nor U27966 (N_27966,N_25080,N_25113);
nor U27967 (N_27967,N_25069,N_25537);
nor U27968 (N_27968,N_26110,N_24154);
and U27969 (N_27969,N_26381,N_25698);
and U27970 (N_27970,N_26913,N_26510);
and U27971 (N_27971,N_25127,N_25634);
xor U27972 (N_27972,N_25796,N_26575);
nand U27973 (N_27973,N_26226,N_25748);
nor U27974 (N_27974,N_25148,N_26288);
xor U27975 (N_27975,N_25098,N_25872);
nor U27976 (N_27976,N_26360,N_25672);
xor U27977 (N_27977,N_24158,N_26432);
nand U27978 (N_27978,N_26673,N_25770);
nand U27979 (N_27979,N_24428,N_26412);
nand U27980 (N_27980,N_24626,N_26539);
nor U27981 (N_27981,N_26864,N_26500);
nor U27982 (N_27982,N_25848,N_26669);
nor U27983 (N_27983,N_25732,N_26414);
and U27984 (N_27984,N_24138,N_24458);
nor U27985 (N_27985,N_26818,N_24256);
or U27986 (N_27986,N_24273,N_26186);
xnor U27987 (N_27987,N_24464,N_25918);
nor U27988 (N_27988,N_24196,N_24638);
nor U27989 (N_27989,N_24136,N_26809);
nor U27990 (N_27990,N_26033,N_24483);
xor U27991 (N_27991,N_24729,N_25615);
xor U27992 (N_27992,N_25304,N_26992);
nor U27993 (N_27993,N_24665,N_24689);
and U27994 (N_27994,N_24479,N_25170);
nand U27995 (N_27995,N_26435,N_26243);
nor U27996 (N_27996,N_25788,N_26323);
xor U27997 (N_27997,N_25806,N_24225);
nand U27998 (N_27998,N_25881,N_25472);
xnor U27999 (N_27999,N_26810,N_26970);
or U28000 (N_28000,N_24022,N_26388);
or U28001 (N_28001,N_25310,N_26328);
nand U28002 (N_28002,N_24459,N_26054);
nand U28003 (N_28003,N_25187,N_25901);
and U28004 (N_28004,N_24498,N_25294);
xor U28005 (N_28005,N_25459,N_26175);
or U28006 (N_28006,N_25144,N_25071);
nor U28007 (N_28007,N_24618,N_24410);
nor U28008 (N_28008,N_25171,N_26752);
and U28009 (N_28009,N_24646,N_24814);
nand U28010 (N_28010,N_25722,N_25822);
xor U28011 (N_28011,N_26204,N_24241);
and U28012 (N_28012,N_25771,N_24124);
nor U28013 (N_28013,N_26532,N_25841);
and U28014 (N_28014,N_24350,N_25710);
and U28015 (N_28015,N_24259,N_24816);
and U28016 (N_28016,N_26349,N_26434);
nor U28017 (N_28017,N_24645,N_26370);
xnor U28018 (N_28018,N_26880,N_24529);
xor U28019 (N_28019,N_26374,N_24708);
and U28020 (N_28020,N_25985,N_24108);
xnor U28021 (N_28021,N_26438,N_24984);
and U28022 (N_28022,N_26948,N_25018);
nand U28023 (N_28023,N_25505,N_24795);
nand U28024 (N_28024,N_25354,N_26585);
and U28025 (N_28025,N_26060,N_26929);
nor U28026 (N_28026,N_26318,N_26505);
and U28027 (N_28027,N_24712,N_26718);
nor U28028 (N_28028,N_24043,N_25128);
nor U28029 (N_28029,N_24519,N_25328);
nand U28030 (N_28030,N_25900,N_24634);
xor U28031 (N_28031,N_25369,N_25800);
and U28032 (N_28032,N_25608,N_25803);
nor U28033 (N_28033,N_25705,N_24268);
and U28034 (N_28034,N_24547,N_26805);
or U28035 (N_28035,N_25665,N_26780);
and U28036 (N_28036,N_25043,N_24829);
nor U28037 (N_28037,N_25267,N_26188);
xnor U28038 (N_28038,N_26106,N_24362);
nor U28039 (N_28039,N_26440,N_25105);
nor U28040 (N_28040,N_26623,N_26553);
xnor U28041 (N_28041,N_24548,N_26420);
and U28042 (N_28042,N_25635,N_24654);
or U28043 (N_28043,N_26936,N_26609);
xnor U28044 (N_28044,N_25523,N_25085);
or U28045 (N_28045,N_25975,N_25446);
nor U28046 (N_28046,N_25114,N_25149);
nand U28047 (N_28047,N_24143,N_24810);
and U28048 (N_28048,N_25048,N_26131);
or U28049 (N_28049,N_26070,N_24192);
xnor U28050 (N_28050,N_25202,N_24967);
or U28051 (N_28051,N_25243,N_24703);
and U28052 (N_28052,N_25166,N_24764);
and U28053 (N_28053,N_26757,N_26278);
or U28054 (N_28054,N_26094,N_26250);
xor U28055 (N_28055,N_26599,N_26224);
or U28056 (N_28056,N_26870,N_25244);
or U28057 (N_28057,N_25473,N_26777);
and U28058 (N_28058,N_25112,N_26199);
xor U28059 (N_28059,N_25808,N_25260);
xor U28060 (N_28060,N_24958,N_24028);
or U28061 (N_28061,N_24861,N_24053);
and U28062 (N_28062,N_26030,N_25602);
nand U28063 (N_28063,N_26390,N_25641);
nand U28064 (N_28064,N_26367,N_25356);
nand U28065 (N_28065,N_26847,N_24572);
and U28066 (N_28066,N_26002,N_24096);
nand U28067 (N_28067,N_24082,N_24830);
nand U28068 (N_28068,N_26404,N_25997);
xnor U28069 (N_28069,N_24775,N_26754);
nand U28070 (N_28070,N_24563,N_24874);
nand U28071 (N_28071,N_26688,N_24088);
nand U28072 (N_28072,N_26953,N_26565);
xor U28073 (N_28073,N_26875,N_24411);
nand U28074 (N_28074,N_26608,N_26961);
nand U28075 (N_28075,N_25108,N_26825);
nand U28076 (N_28076,N_26076,N_25656);
or U28077 (N_28077,N_26813,N_26116);
and U28078 (N_28078,N_26785,N_25927);
nor U28079 (N_28079,N_24391,N_26678);
and U28080 (N_28080,N_26419,N_26523);
nor U28081 (N_28081,N_24465,N_26908);
and U28082 (N_28082,N_24419,N_26262);
xor U28083 (N_28083,N_24333,N_25275);
nand U28084 (N_28084,N_26123,N_26314);
and U28085 (N_28085,N_26901,N_26878);
xor U28086 (N_28086,N_25667,N_24392);
and U28087 (N_28087,N_26590,N_24152);
nand U28088 (N_28088,N_24868,N_25256);
and U28089 (N_28089,N_25165,N_24842);
xor U28090 (N_28090,N_24595,N_24970);
or U28091 (N_28091,N_24758,N_25483);
and U28092 (N_28092,N_26808,N_24127);
nand U28093 (N_28093,N_24291,N_25685);
and U28094 (N_28094,N_24157,N_24528);
or U28095 (N_28095,N_24811,N_25738);
and U28096 (N_28096,N_25518,N_24062);
xor U28097 (N_28097,N_26612,N_24986);
or U28098 (N_28098,N_25766,N_25462);
nor U28099 (N_28099,N_25023,N_26995);
nand U28100 (N_28100,N_24745,N_26638);
nor U28101 (N_28101,N_26922,N_25433);
and U28102 (N_28102,N_24040,N_24212);
and U28103 (N_28103,N_26774,N_25853);
or U28104 (N_28104,N_25619,N_25758);
xnor U28105 (N_28105,N_24667,N_25381);
nand U28106 (N_28106,N_25658,N_24818);
nor U28107 (N_28107,N_25945,N_25312);
or U28108 (N_28108,N_24068,N_26540);
nor U28109 (N_28109,N_25621,N_26897);
nand U28110 (N_28110,N_24948,N_25321);
nand U28111 (N_28111,N_26730,N_25004);
xnor U28112 (N_28112,N_25406,N_24210);
nor U28113 (N_28113,N_26820,N_24092);
xnor U28114 (N_28114,N_26006,N_24622);
xnor U28115 (N_28115,N_25297,N_26977);
nor U28116 (N_28116,N_25534,N_25207);
or U28117 (N_28117,N_24078,N_24744);
or U28118 (N_28118,N_25760,N_26883);
nor U28119 (N_28119,N_26261,N_24118);
or U28120 (N_28120,N_24872,N_25106);
and U28121 (N_28121,N_24888,N_24453);
and U28122 (N_28122,N_24394,N_24813);
xor U28123 (N_28123,N_24881,N_26090);
nor U28124 (N_28124,N_24297,N_24782);
xor U28125 (N_28125,N_26700,N_26891);
nor U28126 (N_28126,N_24692,N_24486);
nand U28127 (N_28127,N_24511,N_25568);
nand U28128 (N_28128,N_24010,N_24142);
nand U28129 (N_28129,N_25124,N_25580);
nor U28130 (N_28130,N_24508,N_24565);
nor U28131 (N_28131,N_25529,N_24761);
nor U28132 (N_28132,N_25431,N_26332);
xor U28133 (N_28133,N_25578,N_25953);
and U28134 (N_28134,N_25205,N_25278);
xnor U28135 (N_28135,N_25764,N_24183);
and U28136 (N_28136,N_25396,N_25561);
xor U28137 (N_28137,N_25003,N_26040);
nand U28138 (N_28138,N_25906,N_24036);
xnor U28139 (N_28139,N_25506,N_26790);
xor U28140 (N_28140,N_26806,N_25225);
nor U28141 (N_28141,N_25313,N_24426);
and U28142 (N_28142,N_26611,N_25522);
nand U28143 (N_28143,N_26446,N_24672);
nand U28144 (N_28144,N_25333,N_24603);
nor U28145 (N_28145,N_25276,N_26248);
or U28146 (N_28146,N_25843,N_24526);
and U28147 (N_28147,N_25973,N_25323);
nand U28148 (N_28148,N_24762,N_25392);
nor U28149 (N_28149,N_26711,N_25617);
xor U28150 (N_28150,N_24938,N_26916);
nor U28151 (N_28151,N_26294,N_24797);
and U28152 (N_28152,N_25096,N_26697);
nand U28153 (N_28153,N_26107,N_25399);
nand U28154 (N_28154,N_24906,N_24070);
xnor U28155 (N_28155,N_24468,N_25838);
and U28156 (N_28156,N_25744,N_25185);
and U28157 (N_28157,N_24000,N_26268);
nor U28158 (N_28158,N_25575,N_24432);
and U28159 (N_28159,N_25816,N_26148);
and U28160 (N_28160,N_26865,N_25306);
or U28161 (N_28161,N_24558,N_25655);
nand U28162 (N_28162,N_24290,N_25567);
or U28163 (N_28163,N_26143,N_25318);
xnor U28164 (N_28164,N_25444,N_26012);
or U28165 (N_28165,N_25648,N_25865);
or U28166 (N_28166,N_25850,N_26031);
nor U28167 (N_28167,N_26055,N_25688);
nor U28168 (N_28168,N_26407,N_24197);
nand U28169 (N_28169,N_25842,N_24585);
or U28170 (N_28170,N_25618,N_24696);
nand U28171 (N_28171,N_26591,N_25217);
and U28172 (N_28172,N_25598,N_25330);
nand U28173 (N_28173,N_26111,N_25661);
xnor U28174 (N_28174,N_24163,N_26649);
nor U28175 (N_28175,N_24787,N_24052);
xnor U28176 (N_28176,N_26651,N_25786);
xnor U28177 (N_28177,N_24067,N_25824);
xor U28178 (N_28178,N_25179,N_26221);
and U28179 (N_28179,N_25993,N_26963);
nand U28180 (N_28180,N_26357,N_25347);
and U28181 (N_28181,N_25690,N_25454);
and U28182 (N_28182,N_24156,N_26413);
nand U28183 (N_28183,N_25035,N_24686);
and U28184 (N_28184,N_26508,N_24251);
and U28185 (N_28185,N_26213,N_24760);
and U28186 (N_28186,N_25357,N_25172);
nand U28187 (N_28187,N_25181,N_26965);
and U28188 (N_28188,N_25022,N_25077);
and U28189 (N_28189,N_26991,N_25721);
xor U28190 (N_28190,N_24016,N_25545);
or U28191 (N_28191,N_26442,N_26078);
nand U28192 (N_28192,N_26470,N_24661);
and U28193 (N_28193,N_26798,N_25531);
and U28194 (N_28194,N_26547,N_24423);
xor U28195 (N_28195,N_26065,N_24057);
nor U28196 (N_28196,N_26057,N_26105);
nand U28197 (N_28197,N_24987,N_26307);
nor U28198 (N_28198,N_24260,N_24409);
and U28199 (N_28199,N_26343,N_26173);
xnor U28200 (N_28200,N_25566,N_25498);
xor U28201 (N_28201,N_24045,N_26973);
and U28202 (N_28202,N_25871,N_25009);
nand U28203 (N_28203,N_26762,N_26233);
nor U28204 (N_28204,N_26363,N_26721);
or U28205 (N_28205,N_24633,N_24023);
xor U28206 (N_28206,N_26490,N_25028);
xor U28207 (N_28207,N_24176,N_26902);
and U28208 (N_28208,N_25493,N_25659);
xor U28209 (N_28209,N_25308,N_24179);
xor U28210 (N_28210,N_25117,N_25189);
xor U28211 (N_28211,N_24716,N_25861);
nand U28212 (N_28212,N_26614,N_26637);
and U28213 (N_28213,N_26359,N_24033);
nand U28214 (N_28214,N_24060,N_24559);
nor U28215 (N_28215,N_26561,N_24443);
and U28216 (N_28216,N_24457,N_25998);
xnor U28217 (N_28217,N_25068,N_25612);
nand U28218 (N_28218,N_26735,N_26124);
and U28219 (N_28219,N_26645,N_26263);
and U28220 (N_28220,N_26696,N_24710);
nand U28221 (N_28221,N_26511,N_24701);
and U28222 (N_28222,N_24704,N_24396);
xnor U28223 (N_28223,N_26471,N_26629);
and U28224 (N_28224,N_25378,N_25223);
and U28225 (N_28225,N_25476,N_26035);
nand U28226 (N_28226,N_26023,N_25214);
xnor U28227 (N_28227,N_25651,N_24593);
xnor U28228 (N_28228,N_26622,N_24845);
or U28229 (N_28229,N_26949,N_25585);
xnor U28230 (N_28230,N_26983,N_24119);
nor U28231 (N_28231,N_25273,N_26159);
and U28232 (N_28232,N_25600,N_25046);
or U28233 (N_28233,N_26616,N_26503);
or U28234 (N_28234,N_24226,N_26824);
and U28235 (N_28235,N_24360,N_25471);
xor U28236 (N_28236,N_24730,N_26335);
or U28237 (N_28237,N_25919,N_26454);
and U28238 (N_28238,N_25562,N_26763);
xor U28239 (N_28239,N_24120,N_26469);
and U28240 (N_28240,N_25869,N_25044);
and U28241 (N_28241,N_24344,N_26292);
nand U28242 (N_28242,N_24484,N_25036);
nor U28243 (N_28243,N_25828,N_26297);
xnor U28244 (N_28244,N_25502,N_25292);
nand U28245 (N_28245,N_26714,N_25899);
and U28246 (N_28246,N_25541,N_24979);
nor U28247 (N_28247,N_25380,N_26274);
and U28248 (N_28248,N_25309,N_24944);
nand U28249 (N_28249,N_24866,N_25033);
nor U28250 (N_28250,N_24632,N_24113);
nand U28251 (N_28251,N_26296,N_25224);
or U28252 (N_28252,N_26603,N_25410);
xnor U28253 (N_28253,N_25349,N_25464);
nor U28254 (N_28254,N_24038,N_24864);
and U28255 (N_28255,N_25250,N_24577);
nand U28256 (N_28256,N_25430,N_24663);
nand U28257 (N_28257,N_26346,N_24345);
nor U28258 (N_28258,N_25984,N_25547);
nand U28259 (N_28259,N_26013,N_24749);
and U28260 (N_28260,N_26218,N_26086);
nor U28261 (N_28261,N_26753,N_25228);
and U28262 (N_28262,N_24601,N_26717);
xor U28263 (N_28263,N_26854,N_26739);
or U28264 (N_28264,N_25960,N_26020);
and U28265 (N_28265,N_26289,N_26439);
xor U28266 (N_28266,N_25206,N_25858);
nand U28267 (N_28267,N_24932,N_24039);
nand U28268 (N_28268,N_26451,N_24968);
nor U28269 (N_28269,N_25765,N_26557);
nor U28270 (N_28270,N_25288,N_26194);
xnor U28271 (N_28271,N_24989,N_24996);
xor U28272 (N_28272,N_24125,N_24870);
nand U28273 (N_28273,N_24462,N_24668);
nand U28274 (N_28274,N_25767,N_25163);
and U28275 (N_28275,N_25880,N_26104);
xor U28276 (N_28276,N_26529,N_25370);
or U28277 (N_28277,N_26577,N_26647);
nor U28278 (N_28278,N_26112,N_25831);
or U28279 (N_28279,N_24277,N_25001);
nor U28280 (N_28280,N_26347,N_24307);
xor U28281 (N_28281,N_24939,N_25402);
nand U28282 (N_28282,N_25818,N_26655);
nand U28283 (N_28283,N_26779,N_24960);
nor U28284 (N_28284,N_25754,N_26545);
xnor U28285 (N_28285,N_25209,N_26190);
or U28286 (N_28286,N_24185,N_24346);
nand U28287 (N_28287,N_24380,N_24153);
or U28288 (N_28288,N_26667,N_26542);
xor U28289 (N_28289,N_25334,N_24901);
nor U28290 (N_28290,N_25302,N_25486);
nor U28291 (N_28291,N_24705,N_24614);
xnor U28292 (N_28292,N_26316,N_26731);
or U28293 (N_28293,N_24655,N_26348);
or U28294 (N_28294,N_24612,N_24857);
xnor U28295 (N_28295,N_25680,N_26368);
xnor U28296 (N_28296,N_26141,N_24834);
xnor U28297 (N_28297,N_24063,N_26628);
nor U28298 (N_28298,N_26845,N_25565);
nand U28299 (N_28299,N_25296,N_25636);
or U28300 (N_28300,N_25940,N_24359);
nand U28301 (N_28301,N_25340,N_25497);
xor U28302 (N_28302,N_26406,N_26409);
or U28303 (N_28303,N_24218,N_24574);
nor U28304 (N_28304,N_24293,N_24550);
xnor U28305 (N_28305,N_25169,N_26884);
xnor U28306 (N_28306,N_24147,N_24180);
nand U28307 (N_28307,N_24920,N_24961);
xor U28308 (N_28308,N_26964,N_26320);
nor U28309 (N_28309,N_26792,N_25876);
or U28310 (N_28310,N_25487,N_24966);
xnor U28311 (N_28311,N_26077,N_24441);
nor U28312 (N_28312,N_25485,N_24616);
and U28313 (N_28313,N_25780,N_26885);
xor U28314 (N_28314,N_26677,N_26528);
nand U28315 (N_28315,N_25079,N_24351);
xor U28316 (N_28316,N_25644,N_26391);
or U28317 (N_28317,N_25156,N_25989);
or U28318 (N_28318,N_24112,N_26656);
and U28319 (N_28319,N_25091,N_24720);
nand U28320 (N_28320,N_26036,N_26476);
nand U28321 (N_28321,N_25377,N_24191);
or U28322 (N_28322,N_25610,N_24080);
or U28323 (N_28323,N_26564,N_24132);
and U28324 (N_28324,N_26923,N_26938);
nor U28325 (N_28325,N_26430,N_25058);
nor U28326 (N_28326,N_26589,N_26017);
or U28327 (N_28327,N_25623,N_24198);
and U28328 (N_28328,N_25733,N_25139);
nor U28329 (N_28329,N_24282,N_24093);
xor U28330 (N_28330,N_24788,N_24571);
xnor U28331 (N_28331,N_25594,N_24531);
and U28332 (N_28332,N_26043,N_25609);
or U28333 (N_28333,N_26097,N_25342);
nor U28334 (N_28334,N_26229,N_25038);
or U28335 (N_28335,N_26799,N_24950);
and U28336 (N_28336,N_24658,N_26566);
nor U28337 (N_28337,N_24407,N_24421);
or U28338 (N_28338,N_24188,N_24239);
xor U28339 (N_28339,N_26671,N_25783);
and U28340 (N_28340,N_26893,N_24541);
xor U28341 (N_28341,N_26230,N_25563);
and U28342 (N_28342,N_25222,N_26482);
nor U28343 (N_28343,N_25521,N_26073);
or U28344 (N_28344,N_26605,N_26237);
nor U28345 (N_28345,N_24718,N_25967);
and U28346 (N_28346,N_25922,N_24404);
xor U28347 (N_28347,N_24150,N_25726);
and U28348 (N_28348,N_25104,N_24530);
nor U28349 (N_28349,N_26000,N_25941);
nor U28350 (N_28350,N_25662,N_26062);
nor U28351 (N_28351,N_24753,N_25191);
or U28352 (N_28352,N_25955,N_24914);
nor U28353 (N_28353,N_24732,N_25176);
and U28354 (N_28354,N_26680,N_24098);
or U28355 (N_28355,N_25525,N_25905);
and U28356 (N_28356,N_24790,N_26621);
or U28357 (N_28357,N_25550,N_26769);
nor U28358 (N_28358,N_26630,N_25723);
xor U28359 (N_28359,N_25394,N_25542);
and U28360 (N_28360,N_26672,N_26416);
xor U28361 (N_28361,N_25988,N_25255);
xor U28362 (N_28362,N_26664,N_24473);
xor U28363 (N_28363,N_24146,N_25136);
or U28364 (N_28364,N_24004,N_24123);
nor U28365 (N_28365,N_25632,N_26914);
xor U28366 (N_28366,N_26530,N_25066);
nor U28367 (N_28367,N_25604,N_25614);
or U28368 (N_28368,N_24094,N_25946);
or U28369 (N_28369,N_26382,N_26687);
or U28370 (N_28370,N_26684,N_25234);
and U28371 (N_28371,N_25259,N_26594);
nor U28372 (N_28372,N_25643,N_25888);
xor U28373 (N_28373,N_26933,N_24352);
xnor U28374 (N_28374,N_25819,N_25703);
or U28375 (N_28375,N_25261,N_24370);
nor U28376 (N_28376,N_24116,N_26418);
or U28377 (N_28377,N_26266,N_24129);
nand U28378 (N_28378,N_25595,N_26828);
and U28379 (N_28379,N_25063,N_25145);
or U28380 (N_28380,N_24353,N_24397);
xnor U28381 (N_28381,N_26136,N_26396);
nand U28382 (N_28382,N_24224,N_26165);
xnor U28383 (N_28383,N_24011,N_26834);
and U28384 (N_28384,N_26038,N_25411);
xnor U28385 (N_28385,N_24408,N_24853);
nand U28386 (N_28386,N_26546,N_26408);
nor U28387 (N_28387,N_24399,N_25622);
or U28388 (N_28388,N_24561,N_25211);
xnor U28389 (N_28389,N_26765,N_25961);
nand U28390 (N_28390,N_25979,N_26958);
or U28391 (N_28391,N_24412,N_26125);
or U28392 (N_28392,N_25024,N_26260);
xnor U28393 (N_28393,N_26007,N_26544);
and U28394 (N_28394,N_25311,N_26364);
and U28395 (N_28395,N_25512,N_24676);
nor U28396 (N_28396,N_25379,N_25712);
nor U28397 (N_28397,N_24827,N_25775);
nor U28398 (N_28398,N_26019,N_26587);
and U28399 (N_28399,N_26309,N_25982);
and U28400 (N_28400,N_25016,N_24235);
nand U28401 (N_28401,N_25902,N_25548);
nand U28402 (N_28402,N_24275,N_26955);
nand U28403 (N_28403,N_26127,N_24590);
and U28404 (N_28404,N_26727,N_26987);
or U28405 (N_28405,N_25949,N_25709);
nand U28406 (N_28406,N_24609,N_24929);
nand U28407 (N_28407,N_24737,N_24451);
xor U28408 (N_28408,N_25939,N_26683);
xnor U28409 (N_28409,N_25779,N_25355);
nor U28410 (N_28410,N_24081,N_25847);
or U28411 (N_28411,N_25376,N_25589);
and U28412 (N_28412,N_24243,N_25797);
and U28413 (N_28413,N_26852,N_24846);
nand U28414 (N_28414,N_26393,N_24941);
and U28415 (N_28415,N_24994,N_26918);
nand U28416 (N_28416,N_26931,N_24107);
nor U28417 (N_28417,N_24555,N_24217);
or U28418 (N_28418,N_24537,N_24900);
and U28419 (N_28419,N_26059,N_24917);
xor U28420 (N_28420,N_25731,N_24065);
nor U28421 (N_28421,N_26744,N_25616);
and U28422 (N_28422,N_24669,N_26362);
nand U28423 (N_28423,N_26521,N_25130);
xnor U28424 (N_28424,N_25835,N_26402);
xor U28425 (N_28425,N_26068,N_25012);
or U28426 (N_28426,N_25115,N_25629);
or U28427 (N_28427,N_24894,N_26444);
or U28428 (N_28428,N_24219,N_25814);
nor U28429 (N_28429,N_24799,N_24500);
xnor U28430 (N_28430,N_24005,N_24886);
and U28431 (N_28431,N_25599,N_25660);
nand U28432 (N_28432,N_24030,N_26142);
nor U28433 (N_28433,N_26794,N_25925);
and U28434 (N_28434,N_25591,N_25134);
xnor U28435 (N_28435,N_25238,N_26548);
or U28436 (N_28436,N_24552,N_24697);
nand U28437 (N_28437,N_24141,N_25590);
or U28438 (N_28438,N_25277,N_24596);
nor U28439 (N_28439,N_24576,N_25743);
nor U28440 (N_28440,N_26942,N_24032);
nand U28441 (N_28441,N_24314,N_25382);
nand U28442 (N_28442,N_25153,N_25666);
nor U28443 (N_28443,N_25851,N_24292);
or U28444 (N_28444,N_25646,N_26679);
or U28445 (N_28445,N_24973,N_24877);
nand U28446 (N_28446,N_24688,N_24510);
nand U28447 (N_28447,N_26392,N_26659);
and U28448 (N_28448,N_24747,N_25649);
and U28449 (N_28449,N_26644,N_25500);
xor U28450 (N_28450,N_24865,N_26275);
and U28451 (N_28451,N_26784,N_26200);
nor U28452 (N_28452,N_26743,N_25581);
nor U28453 (N_28453,N_26177,N_24506);
nor U28454 (N_28454,N_25546,N_26441);
and U28455 (N_28455,N_24238,N_24615);
and U28456 (N_28456,N_26650,N_25477);
nor U28457 (N_28457,N_26867,N_26108);
nor U28458 (N_28458,N_26325,N_24208);
nand U28459 (N_28459,N_26334,N_25088);
xnor U28460 (N_28460,N_24801,N_26044);
nor U28461 (N_28461,N_24296,N_26005);
or U28462 (N_28462,N_25746,N_24819);
nand U28463 (N_28463,N_25051,N_26761);
nor U28464 (N_28464,N_25154,N_24876);
and U28465 (N_28465,N_24539,N_26378);
or U28466 (N_28466,N_25076,N_25350);
nor U28467 (N_28467,N_24456,N_25186);
or U28468 (N_28468,N_26147,N_26342);
or U28469 (N_28469,N_24145,N_24279);
or U28470 (N_28470,N_26909,N_26231);
nand U28471 (N_28471,N_25763,N_26821);
nor U28472 (N_28472,N_26776,N_26251);
xor U28473 (N_28473,N_25020,N_25724);
xnor U28474 (N_28474,N_26311,N_25664);
xor U28475 (N_28475,N_26858,N_26705);
and U28476 (N_28476,N_25969,N_24772);
and U28477 (N_28477,N_25689,N_24311);
or U28478 (N_28478,N_24916,N_25183);
nand U28479 (N_28479,N_24438,N_25231);
nor U28480 (N_28480,N_26247,N_25449);
or U28481 (N_28481,N_26966,N_24012);
nor U28482 (N_28482,N_26358,N_25935);
nand U28483 (N_28483,N_24991,N_26657);
nor U28484 (N_28484,N_24475,N_26455);
nand U28485 (N_28485,N_25147,N_25856);
xor U28486 (N_28486,N_25964,N_24497);
nor U28487 (N_28487,N_25570,N_25262);
and U28488 (N_28488,N_26354,N_24231);
and U28489 (N_28489,N_24824,N_26475);
xor U28490 (N_28490,N_26122,N_25290);
or U28491 (N_28491,N_26156,N_25791);
nand U28492 (N_28492,N_24743,N_25050);
nand U28493 (N_28493,N_26196,N_24434);
or U28494 (N_28494,N_26527,N_24207);
or U28495 (N_28495,N_26886,N_26489);
and U28496 (N_28496,N_26760,N_26410);
and U28497 (N_28497,N_24159,N_24228);
and U28498 (N_28498,N_25784,N_26081);
xor U28499 (N_28499,N_24974,N_25219);
and U28500 (N_28500,N_24676,N_25217);
and U28501 (N_28501,N_25758,N_24699);
nand U28502 (N_28502,N_26847,N_24245);
nand U28503 (N_28503,N_25265,N_25620);
xnor U28504 (N_28504,N_25692,N_26441);
or U28505 (N_28505,N_26221,N_24704);
or U28506 (N_28506,N_24279,N_24692);
or U28507 (N_28507,N_24456,N_24824);
or U28508 (N_28508,N_26072,N_26323);
and U28509 (N_28509,N_25511,N_25930);
nand U28510 (N_28510,N_26383,N_26647);
xor U28511 (N_28511,N_24243,N_26417);
nor U28512 (N_28512,N_24988,N_25293);
nand U28513 (N_28513,N_26910,N_26424);
and U28514 (N_28514,N_24440,N_25629);
nand U28515 (N_28515,N_25044,N_26748);
xnor U28516 (N_28516,N_25228,N_25129);
xor U28517 (N_28517,N_26421,N_24884);
xnor U28518 (N_28518,N_25941,N_25896);
and U28519 (N_28519,N_26316,N_25798);
nand U28520 (N_28520,N_25851,N_26269);
nand U28521 (N_28521,N_26413,N_26236);
and U28522 (N_28522,N_25123,N_24911);
nand U28523 (N_28523,N_24558,N_26994);
xnor U28524 (N_28524,N_24244,N_24605);
nand U28525 (N_28525,N_25450,N_24816);
xnor U28526 (N_28526,N_24850,N_26880);
nand U28527 (N_28527,N_24481,N_24259);
nand U28528 (N_28528,N_26466,N_26705);
or U28529 (N_28529,N_25670,N_25036);
and U28530 (N_28530,N_24853,N_26457);
xnor U28531 (N_28531,N_24994,N_26658);
nand U28532 (N_28532,N_26717,N_26322);
nand U28533 (N_28533,N_25924,N_26614);
or U28534 (N_28534,N_26215,N_24070);
nand U28535 (N_28535,N_25434,N_25979);
nor U28536 (N_28536,N_25414,N_24429);
and U28537 (N_28537,N_24866,N_26402);
xor U28538 (N_28538,N_24422,N_24694);
xor U28539 (N_28539,N_25027,N_26716);
or U28540 (N_28540,N_24469,N_26807);
nor U28541 (N_28541,N_26674,N_24101);
and U28542 (N_28542,N_24115,N_24947);
nor U28543 (N_28543,N_26488,N_26596);
and U28544 (N_28544,N_26030,N_26263);
xnor U28545 (N_28545,N_24589,N_25197);
and U28546 (N_28546,N_26886,N_24924);
nand U28547 (N_28547,N_25332,N_26968);
nand U28548 (N_28548,N_25433,N_25326);
and U28549 (N_28549,N_26247,N_25415);
nor U28550 (N_28550,N_26774,N_25288);
and U28551 (N_28551,N_25587,N_25916);
nor U28552 (N_28552,N_25033,N_24455);
or U28553 (N_28553,N_24374,N_26612);
xnor U28554 (N_28554,N_26473,N_25435);
xnor U28555 (N_28555,N_25322,N_24595);
nor U28556 (N_28556,N_24583,N_26224);
and U28557 (N_28557,N_25160,N_26970);
xor U28558 (N_28558,N_24201,N_26401);
or U28559 (N_28559,N_25745,N_26610);
nand U28560 (N_28560,N_24427,N_25374);
xor U28561 (N_28561,N_24974,N_25730);
nor U28562 (N_28562,N_25679,N_24026);
or U28563 (N_28563,N_25572,N_24886);
and U28564 (N_28564,N_25362,N_24992);
xor U28565 (N_28565,N_25971,N_25241);
nor U28566 (N_28566,N_26152,N_24630);
or U28567 (N_28567,N_25601,N_26263);
nor U28568 (N_28568,N_25266,N_25713);
or U28569 (N_28569,N_25599,N_26146);
and U28570 (N_28570,N_25488,N_25386);
and U28571 (N_28571,N_25893,N_24661);
or U28572 (N_28572,N_25773,N_26499);
nand U28573 (N_28573,N_26621,N_25729);
and U28574 (N_28574,N_24048,N_26573);
xnor U28575 (N_28575,N_25859,N_24010);
or U28576 (N_28576,N_25781,N_26498);
nand U28577 (N_28577,N_26757,N_24771);
nor U28578 (N_28578,N_26146,N_24780);
xnor U28579 (N_28579,N_25492,N_26130);
xor U28580 (N_28580,N_26269,N_26489);
and U28581 (N_28581,N_26794,N_24469);
nand U28582 (N_28582,N_24067,N_24459);
and U28583 (N_28583,N_26656,N_26047);
nand U28584 (N_28584,N_24480,N_26764);
nor U28585 (N_28585,N_24333,N_24348);
nand U28586 (N_28586,N_26517,N_25545);
nor U28587 (N_28587,N_25034,N_25330);
nor U28588 (N_28588,N_24782,N_26855);
nand U28589 (N_28589,N_26690,N_25071);
and U28590 (N_28590,N_25978,N_26774);
xor U28591 (N_28591,N_25283,N_24293);
xor U28592 (N_28592,N_26655,N_26339);
or U28593 (N_28593,N_25599,N_26598);
or U28594 (N_28594,N_26194,N_25905);
or U28595 (N_28595,N_24871,N_26334);
nor U28596 (N_28596,N_24124,N_26236);
nand U28597 (N_28597,N_26964,N_26924);
and U28598 (N_28598,N_26076,N_26773);
xor U28599 (N_28599,N_24223,N_24944);
or U28600 (N_28600,N_24203,N_25485);
and U28601 (N_28601,N_25277,N_24726);
and U28602 (N_28602,N_25330,N_25015);
and U28603 (N_28603,N_26040,N_24057);
and U28604 (N_28604,N_24929,N_25453);
nor U28605 (N_28605,N_25355,N_26253);
nand U28606 (N_28606,N_25614,N_26345);
or U28607 (N_28607,N_25464,N_25223);
nand U28608 (N_28608,N_26949,N_26749);
nand U28609 (N_28609,N_26379,N_25702);
nor U28610 (N_28610,N_25340,N_24985);
nor U28611 (N_28611,N_26193,N_24542);
nor U28612 (N_28612,N_24420,N_24657);
nand U28613 (N_28613,N_26370,N_24276);
or U28614 (N_28614,N_25719,N_24702);
and U28615 (N_28615,N_25651,N_25469);
nor U28616 (N_28616,N_25881,N_24181);
xor U28617 (N_28617,N_24001,N_26788);
nand U28618 (N_28618,N_25672,N_26362);
nand U28619 (N_28619,N_26387,N_26420);
nor U28620 (N_28620,N_26173,N_25211);
xnor U28621 (N_28621,N_26682,N_26310);
and U28622 (N_28622,N_25800,N_25774);
nor U28623 (N_28623,N_26418,N_25265);
or U28624 (N_28624,N_26937,N_24580);
nor U28625 (N_28625,N_25971,N_25023);
nand U28626 (N_28626,N_26145,N_24675);
or U28627 (N_28627,N_26125,N_24377);
xnor U28628 (N_28628,N_26505,N_24689);
or U28629 (N_28629,N_24415,N_26656);
nand U28630 (N_28630,N_25406,N_26251);
and U28631 (N_28631,N_26147,N_26188);
nor U28632 (N_28632,N_26599,N_25996);
nor U28633 (N_28633,N_24858,N_26407);
or U28634 (N_28634,N_25417,N_26305);
xnor U28635 (N_28635,N_26232,N_25695);
nand U28636 (N_28636,N_26992,N_24823);
nand U28637 (N_28637,N_24413,N_24870);
nor U28638 (N_28638,N_24988,N_25252);
and U28639 (N_28639,N_24832,N_26659);
xnor U28640 (N_28640,N_25686,N_26765);
or U28641 (N_28641,N_25424,N_24162);
xor U28642 (N_28642,N_25464,N_24651);
nor U28643 (N_28643,N_26138,N_24851);
or U28644 (N_28644,N_24224,N_26426);
nor U28645 (N_28645,N_25191,N_25876);
nand U28646 (N_28646,N_26559,N_26742);
nand U28647 (N_28647,N_25757,N_25362);
or U28648 (N_28648,N_25201,N_24047);
or U28649 (N_28649,N_25450,N_24929);
nor U28650 (N_28650,N_26362,N_26864);
or U28651 (N_28651,N_26893,N_26854);
and U28652 (N_28652,N_24381,N_26928);
and U28653 (N_28653,N_25624,N_25692);
nand U28654 (N_28654,N_26187,N_24440);
or U28655 (N_28655,N_26092,N_25398);
xor U28656 (N_28656,N_26735,N_26367);
xnor U28657 (N_28657,N_24957,N_25292);
nor U28658 (N_28658,N_24211,N_24218);
xor U28659 (N_28659,N_25483,N_26052);
or U28660 (N_28660,N_24652,N_26479);
xor U28661 (N_28661,N_26791,N_26224);
nand U28662 (N_28662,N_25326,N_26562);
xnor U28663 (N_28663,N_24698,N_24075);
or U28664 (N_28664,N_24692,N_26533);
nor U28665 (N_28665,N_24404,N_24275);
xor U28666 (N_28666,N_25422,N_24426);
xnor U28667 (N_28667,N_25976,N_25164);
nor U28668 (N_28668,N_26998,N_24329);
xor U28669 (N_28669,N_26095,N_24233);
or U28670 (N_28670,N_25139,N_25058);
nand U28671 (N_28671,N_25220,N_26598);
and U28672 (N_28672,N_25830,N_25483);
nor U28673 (N_28673,N_24697,N_26194);
or U28674 (N_28674,N_25917,N_25359);
nor U28675 (N_28675,N_25702,N_24159);
xnor U28676 (N_28676,N_24488,N_26883);
nor U28677 (N_28677,N_26716,N_26134);
nor U28678 (N_28678,N_24105,N_25749);
nand U28679 (N_28679,N_26199,N_25361);
nor U28680 (N_28680,N_25568,N_24741);
nor U28681 (N_28681,N_26253,N_25964);
nor U28682 (N_28682,N_25980,N_24438);
or U28683 (N_28683,N_24665,N_26760);
nand U28684 (N_28684,N_26439,N_24573);
nand U28685 (N_28685,N_26746,N_26201);
and U28686 (N_28686,N_24844,N_24426);
nand U28687 (N_28687,N_25210,N_26944);
or U28688 (N_28688,N_24691,N_25077);
and U28689 (N_28689,N_26847,N_24521);
and U28690 (N_28690,N_25169,N_25421);
xor U28691 (N_28691,N_24074,N_25988);
or U28692 (N_28692,N_24364,N_24762);
and U28693 (N_28693,N_24861,N_26986);
or U28694 (N_28694,N_24767,N_26271);
nand U28695 (N_28695,N_25771,N_25527);
or U28696 (N_28696,N_26223,N_26544);
nor U28697 (N_28697,N_25768,N_24751);
or U28698 (N_28698,N_25322,N_24581);
or U28699 (N_28699,N_26439,N_25610);
nor U28700 (N_28700,N_24158,N_25984);
nand U28701 (N_28701,N_26943,N_24005);
or U28702 (N_28702,N_25315,N_26939);
or U28703 (N_28703,N_25224,N_24787);
xnor U28704 (N_28704,N_26489,N_25949);
or U28705 (N_28705,N_26110,N_25507);
nand U28706 (N_28706,N_24489,N_25574);
and U28707 (N_28707,N_26090,N_25798);
and U28708 (N_28708,N_24787,N_26067);
nand U28709 (N_28709,N_25557,N_25810);
xnor U28710 (N_28710,N_26164,N_24207);
xnor U28711 (N_28711,N_25095,N_25834);
or U28712 (N_28712,N_24948,N_26489);
xnor U28713 (N_28713,N_24712,N_25864);
nor U28714 (N_28714,N_24548,N_26675);
and U28715 (N_28715,N_25737,N_25889);
nand U28716 (N_28716,N_25784,N_24708);
or U28717 (N_28717,N_25299,N_24152);
or U28718 (N_28718,N_25080,N_26597);
nand U28719 (N_28719,N_26006,N_26746);
nand U28720 (N_28720,N_26915,N_26842);
nor U28721 (N_28721,N_24043,N_26907);
nand U28722 (N_28722,N_24624,N_24476);
xnor U28723 (N_28723,N_24671,N_24255);
or U28724 (N_28724,N_26169,N_24040);
and U28725 (N_28725,N_26463,N_25310);
xnor U28726 (N_28726,N_25767,N_26195);
nand U28727 (N_28727,N_24177,N_25260);
nor U28728 (N_28728,N_24612,N_24927);
nand U28729 (N_28729,N_24019,N_25225);
or U28730 (N_28730,N_25391,N_26908);
nand U28731 (N_28731,N_25898,N_25048);
xor U28732 (N_28732,N_24699,N_24870);
and U28733 (N_28733,N_24252,N_25863);
and U28734 (N_28734,N_26762,N_26185);
nor U28735 (N_28735,N_25645,N_25315);
or U28736 (N_28736,N_25285,N_26279);
or U28737 (N_28737,N_24126,N_26073);
and U28738 (N_28738,N_26731,N_24534);
nand U28739 (N_28739,N_24070,N_25736);
nor U28740 (N_28740,N_25519,N_26121);
and U28741 (N_28741,N_24097,N_26943);
and U28742 (N_28742,N_24377,N_25757);
nand U28743 (N_28743,N_25681,N_26874);
nand U28744 (N_28744,N_24116,N_26939);
xor U28745 (N_28745,N_26209,N_24791);
or U28746 (N_28746,N_24377,N_25696);
nand U28747 (N_28747,N_24059,N_25876);
and U28748 (N_28748,N_24533,N_25070);
nand U28749 (N_28749,N_25656,N_24151);
and U28750 (N_28750,N_25136,N_26382);
nor U28751 (N_28751,N_24837,N_25170);
nand U28752 (N_28752,N_25575,N_26256);
nor U28753 (N_28753,N_26405,N_26720);
nor U28754 (N_28754,N_24515,N_24465);
and U28755 (N_28755,N_26034,N_25954);
or U28756 (N_28756,N_26620,N_25757);
and U28757 (N_28757,N_24126,N_25341);
or U28758 (N_28758,N_26479,N_25450);
xnor U28759 (N_28759,N_26801,N_24918);
nand U28760 (N_28760,N_24853,N_25577);
nand U28761 (N_28761,N_24632,N_26456);
or U28762 (N_28762,N_26049,N_25191);
nand U28763 (N_28763,N_26748,N_25293);
or U28764 (N_28764,N_26363,N_26755);
xnor U28765 (N_28765,N_24907,N_25236);
nand U28766 (N_28766,N_25218,N_24131);
nand U28767 (N_28767,N_24304,N_24830);
or U28768 (N_28768,N_24221,N_25042);
and U28769 (N_28769,N_26387,N_25320);
nor U28770 (N_28770,N_25748,N_24070);
or U28771 (N_28771,N_25691,N_24604);
and U28772 (N_28772,N_24283,N_24543);
nand U28773 (N_28773,N_26147,N_26274);
and U28774 (N_28774,N_25058,N_26625);
nor U28775 (N_28775,N_26180,N_25046);
xor U28776 (N_28776,N_24908,N_24916);
and U28777 (N_28777,N_26417,N_25515);
nand U28778 (N_28778,N_25589,N_26788);
xnor U28779 (N_28779,N_24791,N_24331);
xor U28780 (N_28780,N_26669,N_26824);
xnor U28781 (N_28781,N_24157,N_26167);
and U28782 (N_28782,N_26542,N_24758);
and U28783 (N_28783,N_26703,N_26441);
or U28784 (N_28784,N_25841,N_26627);
or U28785 (N_28785,N_24028,N_25042);
nand U28786 (N_28786,N_25503,N_24044);
and U28787 (N_28787,N_25194,N_25792);
nand U28788 (N_28788,N_24314,N_25014);
nor U28789 (N_28789,N_26646,N_24896);
and U28790 (N_28790,N_26413,N_26448);
or U28791 (N_28791,N_26820,N_25759);
or U28792 (N_28792,N_25210,N_24716);
nor U28793 (N_28793,N_24238,N_25049);
and U28794 (N_28794,N_24567,N_24225);
and U28795 (N_28795,N_26238,N_26386);
xnor U28796 (N_28796,N_25055,N_25693);
nand U28797 (N_28797,N_24982,N_24425);
and U28798 (N_28798,N_25984,N_25045);
xor U28799 (N_28799,N_25349,N_26956);
or U28800 (N_28800,N_25157,N_24855);
xnor U28801 (N_28801,N_25266,N_25002);
or U28802 (N_28802,N_24114,N_24251);
xor U28803 (N_28803,N_25506,N_25613);
or U28804 (N_28804,N_24860,N_26775);
or U28805 (N_28805,N_24752,N_26591);
xor U28806 (N_28806,N_24227,N_25438);
xor U28807 (N_28807,N_24779,N_26167);
or U28808 (N_28808,N_26808,N_25206);
nand U28809 (N_28809,N_26892,N_26711);
nand U28810 (N_28810,N_25820,N_24317);
nand U28811 (N_28811,N_25031,N_24934);
and U28812 (N_28812,N_25262,N_24282);
xnor U28813 (N_28813,N_25489,N_26881);
nor U28814 (N_28814,N_24922,N_24712);
xnor U28815 (N_28815,N_24625,N_24752);
xnor U28816 (N_28816,N_24875,N_26861);
nor U28817 (N_28817,N_24084,N_24274);
or U28818 (N_28818,N_24470,N_26166);
xnor U28819 (N_28819,N_26866,N_26702);
nand U28820 (N_28820,N_25112,N_24186);
xnor U28821 (N_28821,N_25070,N_24947);
xnor U28822 (N_28822,N_25965,N_24621);
and U28823 (N_28823,N_26439,N_25002);
or U28824 (N_28824,N_24040,N_25309);
nand U28825 (N_28825,N_25268,N_25662);
nand U28826 (N_28826,N_26210,N_25159);
or U28827 (N_28827,N_25763,N_26994);
xnor U28828 (N_28828,N_26306,N_25047);
nor U28829 (N_28829,N_26474,N_25656);
nand U28830 (N_28830,N_26066,N_25827);
and U28831 (N_28831,N_26943,N_26781);
and U28832 (N_28832,N_24372,N_25937);
and U28833 (N_28833,N_26829,N_24105);
nand U28834 (N_28834,N_25546,N_24789);
or U28835 (N_28835,N_25189,N_25087);
nand U28836 (N_28836,N_26141,N_24156);
nor U28837 (N_28837,N_26770,N_24603);
nand U28838 (N_28838,N_25528,N_24000);
and U28839 (N_28839,N_25102,N_26163);
xor U28840 (N_28840,N_26463,N_24071);
and U28841 (N_28841,N_25100,N_26724);
xor U28842 (N_28842,N_25592,N_26862);
xnor U28843 (N_28843,N_24887,N_25173);
nand U28844 (N_28844,N_26004,N_25008);
nor U28845 (N_28845,N_25114,N_25513);
or U28846 (N_28846,N_26672,N_25225);
nand U28847 (N_28847,N_26762,N_25529);
xnor U28848 (N_28848,N_24491,N_25903);
or U28849 (N_28849,N_25643,N_25352);
xor U28850 (N_28850,N_24833,N_24422);
xnor U28851 (N_28851,N_24706,N_25338);
and U28852 (N_28852,N_24832,N_26166);
nor U28853 (N_28853,N_25153,N_24879);
xor U28854 (N_28854,N_26182,N_24689);
and U28855 (N_28855,N_26025,N_26077);
or U28856 (N_28856,N_25096,N_25537);
and U28857 (N_28857,N_25436,N_25358);
and U28858 (N_28858,N_26039,N_25167);
nand U28859 (N_28859,N_26584,N_26218);
or U28860 (N_28860,N_24937,N_24031);
nor U28861 (N_28861,N_26301,N_25576);
nand U28862 (N_28862,N_26089,N_25147);
nand U28863 (N_28863,N_25492,N_24136);
and U28864 (N_28864,N_24110,N_25636);
nand U28865 (N_28865,N_24266,N_25618);
nand U28866 (N_28866,N_26291,N_24487);
and U28867 (N_28867,N_25300,N_24737);
xor U28868 (N_28868,N_24438,N_26458);
nor U28869 (N_28869,N_25444,N_26970);
xor U28870 (N_28870,N_25932,N_25848);
nand U28871 (N_28871,N_25387,N_25896);
xor U28872 (N_28872,N_24863,N_26907);
xor U28873 (N_28873,N_24937,N_26465);
nor U28874 (N_28874,N_25301,N_24611);
xnor U28875 (N_28875,N_25334,N_26309);
nor U28876 (N_28876,N_26806,N_25791);
nor U28877 (N_28877,N_26902,N_24310);
or U28878 (N_28878,N_24130,N_24384);
nor U28879 (N_28879,N_26127,N_25150);
xnor U28880 (N_28880,N_24965,N_26036);
and U28881 (N_28881,N_24922,N_26339);
or U28882 (N_28882,N_25459,N_24463);
xnor U28883 (N_28883,N_25727,N_26358);
xnor U28884 (N_28884,N_25775,N_24020);
xor U28885 (N_28885,N_24219,N_25747);
nand U28886 (N_28886,N_25999,N_25290);
xnor U28887 (N_28887,N_24274,N_24863);
or U28888 (N_28888,N_26396,N_24080);
nor U28889 (N_28889,N_24978,N_26719);
xnor U28890 (N_28890,N_25000,N_24574);
xor U28891 (N_28891,N_26554,N_25310);
or U28892 (N_28892,N_24893,N_26785);
nor U28893 (N_28893,N_26419,N_26936);
xor U28894 (N_28894,N_25974,N_24682);
xor U28895 (N_28895,N_26619,N_24967);
and U28896 (N_28896,N_26508,N_24313);
nand U28897 (N_28897,N_26508,N_26018);
nor U28898 (N_28898,N_25607,N_25538);
or U28899 (N_28899,N_24751,N_25766);
and U28900 (N_28900,N_26269,N_26712);
nand U28901 (N_28901,N_24067,N_25795);
xnor U28902 (N_28902,N_25417,N_24876);
xor U28903 (N_28903,N_24468,N_26454);
nand U28904 (N_28904,N_25394,N_24817);
xnor U28905 (N_28905,N_24282,N_25696);
or U28906 (N_28906,N_24496,N_25421);
or U28907 (N_28907,N_24441,N_25845);
or U28908 (N_28908,N_25723,N_25500);
xnor U28909 (N_28909,N_26245,N_26747);
nor U28910 (N_28910,N_26853,N_26844);
xnor U28911 (N_28911,N_24461,N_24550);
xnor U28912 (N_28912,N_24590,N_26698);
nor U28913 (N_28913,N_25009,N_26432);
nor U28914 (N_28914,N_24118,N_26538);
nor U28915 (N_28915,N_25203,N_26271);
nand U28916 (N_28916,N_26323,N_25666);
nand U28917 (N_28917,N_24795,N_24024);
nor U28918 (N_28918,N_24690,N_24240);
and U28919 (N_28919,N_24764,N_25645);
or U28920 (N_28920,N_25552,N_24551);
nand U28921 (N_28921,N_25040,N_25195);
xnor U28922 (N_28922,N_24153,N_26107);
nand U28923 (N_28923,N_25273,N_26901);
and U28924 (N_28924,N_26428,N_26317);
nand U28925 (N_28925,N_25649,N_24020);
or U28926 (N_28926,N_25877,N_26151);
nand U28927 (N_28927,N_26219,N_26510);
or U28928 (N_28928,N_25986,N_25969);
nor U28929 (N_28929,N_26305,N_26151);
or U28930 (N_28930,N_26427,N_25718);
and U28931 (N_28931,N_26462,N_25148);
and U28932 (N_28932,N_26940,N_26955);
and U28933 (N_28933,N_24089,N_25767);
nand U28934 (N_28934,N_25078,N_25443);
and U28935 (N_28935,N_25217,N_25010);
nand U28936 (N_28936,N_25526,N_24518);
nand U28937 (N_28937,N_25108,N_24069);
or U28938 (N_28938,N_24437,N_26448);
xnor U28939 (N_28939,N_25549,N_25518);
nor U28940 (N_28940,N_26183,N_25804);
xor U28941 (N_28941,N_25944,N_26548);
nor U28942 (N_28942,N_24858,N_24062);
xor U28943 (N_28943,N_26082,N_25174);
or U28944 (N_28944,N_26601,N_24847);
xor U28945 (N_28945,N_25933,N_25414);
and U28946 (N_28946,N_26999,N_26926);
xor U28947 (N_28947,N_26336,N_25244);
nor U28948 (N_28948,N_25849,N_25187);
nor U28949 (N_28949,N_25723,N_25372);
nand U28950 (N_28950,N_25424,N_24400);
or U28951 (N_28951,N_24097,N_26621);
xnor U28952 (N_28952,N_26144,N_25984);
nor U28953 (N_28953,N_26718,N_25672);
and U28954 (N_28954,N_25362,N_24896);
nor U28955 (N_28955,N_26272,N_26596);
nand U28956 (N_28956,N_25191,N_24414);
or U28957 (N_28957,N_25424,N_24695);
nand U28958 (N_28958,N_24432,N_26184);
or U28959 (N_28959,N_26271,N_26651);
xnor U28960 (N_28960,N_26555,N_25231);
xnor U28961 (N_28961,N_26037,N_25125);
xor U28962 (N_28962,N_26597,N_24636);
nand U28963 (N_28963,N_26769,N_24100);
and U28964 (N_28964,N_24150,N_26837);
nor U28965 (N_28965,N_24844,N_24090);
nor U28966 (N_28966,N_25903,N_24151);
nand U28967 (N_28967,N_24607,N_25449);
or U28968 (N_28968,N_24971,N_25244);
nand U28969 (N_28969,N_26844,N_26843);
or U28970 (N_28970,N_25729,N_25253);
nor U28971 (N_28971,N_25415,N_25964);
nand U28972 (N_28972,N_25137,N_24696);
xor U28973 (N_28973,N_25765,N_24615);
nand U28974 (N_28974,N_25761,N_26221);
nor U28975 (N_28975,N_25788,N_24375);
xnor U28976 (N_28976,N_26532,N_26885);
nor U28977 (N_28977,N_24882,N_26540);
and U28978 (N_28978,N_26620,N_24645);
and U28979 (N_28979,N_25916,N_26350);
nor U28980 (N_28980,N_26480,N_25279);
and U28981 (N_28981,N_25630,N_26978);
and U28982 (N_28982,N_24644,N_25969);
nor U28983 (N_28983,N_25006,N_25657);
nor U28984 (N_28984,N_26276,N_26294);
nor U28985 (N_28985,N_25714,N_26170);
and U28986 (N_28986,N_26636,N_24036);
or U28987 (N_28987,N_25736,N_25302);
and U28988 (N_28988,N_25220,N_24103);
or U28989 (N_28989,N_25485,N_26053);
nand U28990 (N_28990,N_26578,N_24901);
or U28991 (N_28991,N_24928,N_26331);
xor U28992 (N_28992,N_26149,N_26687);
and U28993 (N_28993,N_24319,N_26277);
or U28994 (N_28994,N_26243,N_26293);
nand U28995 (N_28995,N_24575,N_26391);
or U28996 (N_28996,N_25224,N_26049);
nand U28997 (N_28997,N_24864,N_25062);
nor U28998 (N_28998,N_26988,N_25354);
or U28999 (N_28999,N_25062,N_25697);
or U29000 (N_29000,N_24009,N_25426);
nor U29001 (N_29001,N_26643,N_24321);
nor U29002 (N_29002,N_26579,N_24794);
nor U29003 (N_29003,N_26504,N_25290);
nor U29004 (N_29004,N_24102,N_24806);
nand U29005 (N_29005,N_24018,N_25941);
xnor U29006 (N_29006,N_26819,N_24279);
nor U29007 (N_29007,N_24407,N_24949);
xor U29008 (N_29008,N_26849,N_25613);
and U29009 (N_29009,N_25684,N_25798);
and U29010 (N_29010,N_26430,N_24802);
nand U29011 (N_29011,N_25842,N_26380);
xor U29012 (N_29012,N_26285,N_25230);
xor U29013 (N_29013,N_25641,N_24638);
nor U29014 (N_29014,N_24145,N_24404);
and U29015 (N_29015,N_26931,N_26331);
and U29016 (N_29016,N_26526,N_25661);
or U29017 (N_29017,N_26950,N_26813);
or U29018 (N_29018,N_24961,N_26467);
and U29019 (N_29019,N_25204,N_24977);
and U29020 (N_29020,N_25729,N_25215);
nand U29021 (N_29021,N_24122,N_24585);
xnor U29022 (N_29022,N_25071,N_25278);
and U29023 (N_29023,N_24398,N_24919);
and U29024 (N_29024,N_26481,N_26364);
or U29025 (N_29025,N_24839,N_25750);
nand U29026 (N_29026,N_24060,N_24781);
xor U29027 (N_29027,N_24001,N_25343);
xnor U29028 (N_29028,N_26844,N_26407);
and U29029 (N_29029,N_25680,N_24691);
and U29030 (N_29030,N_26403,N_26688);
nor U29031 (N_29031,N_24800,N_26591);
xor U29032 (N_29032,N_24171,N_25125);
xor U29033 (N_29033,N_24430,N_26168);
nand U29034 (N_29034,N_25474,N_24807);
xnor U29035 (N_29035,N_24085,N_26295);
xor U29036 (N_29036,N_25434,N_25507);
xnor U29037 (N_29037,N_26964,N_26230);
and U29038 (N_29038,N_25608,N_26609);
or U29039 (N_29039,N_25286,N_25791);
and U29040 (N_29040,N_26944,N_26254);
or U29041 (N_29041,N_24340,N_26018);
nand U29042 (N_29042,N_25956,N_24624);
or U29043 (N_29043,N_24920,N_26740);
or U29044 (N_29044,N_26281,N_24029);
nor U29045 (N_29045,N_25410,N_25715);
and U29046 (N_29046,N_26075,N_26486);
nand U29047 (N_29047,N_25874,N_25071);
nand U29048 (N_29048,N_26548,N_25509);
or U29049 (N_29049,N_26024,N_25951);
xnor U29050 (N_29050,N_26968,N_24649);
and U29051 (N_29051,N_25490,N_25541);
or U29052 (N_29052,N_24205,N_26794);
nand U29053 (N_29053,N_25277,N_26045);
or U29054 (N_29054,N_26996,N_25089);
nor U29055 (N_29055,N_24259,N_24508);
nor U29056 (N_29056,N_26901,N_24437);
xnor U29057 (N_29057,N_25836,N_26235);
xnor U29058 (N_29058,N_25904,N_24367);
xnor U29059 (N_29059,N_25411,N_25437);
xor U29060 (N_29060,N_25782,N_25766);
nand U29061 (N_29061,N_26923,N_25031);
xnor U29062 (N_29062,N_26902,N_26618);
and U29063 (N_29063,N_24155,N_24325);
nand U29064 (N_29064,N_24476,N_26890);
xor U29065 (N_29065,N_25000,N_26271);
nor U29066 (N_29066,N_25122,N_25625);
nor U29067 (N_29067,N_24241,N_26484);
and U29068 (N_29068,N_24960,N_24244);
or U29069 (N_29069,N_24071,N_24946);
and U29070 (N_29070,N_26799,N_26118);
or U29071 (N_29071,N_25700,N_26101);
nand U29072 (N_29072,N_25746,N_25071);
nor U29073 (N_29073,N_24769,N_26265);
nor U29074 (N_29074,N_24726,N_26917);
or U29075 (N_29075,N_26491,N_24394);
and U29076 (N_29076,N_26480,N_26066);
nand U29077 (N_29077,N_25341,N_24880);
nand U29078 (N_29078,N_26652,N_24307);
xor U29079 (N_29079,N_24091,N_25495);
or U29080 (N_29080,N_24411,N_25796);
nor U29081 (N_29081,N_25567,N_24279);
nor U29082 (N_29082,N_26483,N_26307);
nand U29083 (N_29083,N_26488,N_24109);
and U29084 (N_29084,N_24628,N_25458);
or U29085 (N_29085,N_24842,N_25702);
nand U29086 (N_29086,N_24567,N_24538);
nor U29087 (N_29087,N_24940,N_26806);
and U29088 (N_29088,N_25914,N_24407);
xnor U29089 (N_29089,N_25775,N_26232);
and U29090 (N_29090,N_25106,N_26010);
or U29091 (N_29091,N_24328,N_26453);
nand U29092 (N_29092,N_25230,N_26739);
nor U29093 (N_29093,N_24146,N_24176);
or U29094 (N_29094,N_25519,N_26005);
nand U29095 (N_29095,N_25069,N_24256);
nor U29096 (N_29096,N_24796,N_25410);
or U29097 (N_29097,N_26468,N_24427);
nor U29098 (N_29098,N_24007,N_26981);
xnor U29099 (N_29099,N_25597,N_24946);
or U29100 (N_29100,N_26592,N_24583);
xnor U29101 (N_29101,N_26436,N_24333);
and U29102 (N_29102,N_24350,N_26977);
xor U29103 (N_29103,N_24275,N_26134);
nor U29104 (N_29104,N_24784,N_25307);
xnor U29105 (N_29105,N_26794,N_25960);
and U29106 (N_29106,N_24025,N_26449);
nand U29107 (N_29107,N_26857,N_25415);
nor U29108 (N_29108,N_26573,N_26184);
or U29109 (N_29109,N_24197,N_24539);
nor U29110 (N_29110,N_25158,N_25431);
nor U29111 (N_29111,N_25588,N_26440);
xor U29112 (N_29112,N_26049,N_26825);
and U29113 (N_29113,N_24126,N_25393);
xnor U29114 (N_29114,N_24153,N_25947);
and U29115 (N_29115,N_25623,N_24301);
or U29116 (N_29116,N_26900,N_25177);
nand U29117 (N_29117,N_25981,N_25841);
xnor U29118 (N_29118,N_26764,N_24850);
or U29119 (N_29119,N_26598,N_24369);
nand U29120 (N_29120,N_26108,N_25591);
xor U29121 (N_29121,N_26391,N_26123);
and U29122 (N_29122,N_25980,N_25775);
or U29123 (N_29123,N_24864,N_26809);
nand U29124 (N_29124,N_24438,N_26623);
or U29125 (N_29125,N_25306,N_26105);
nor U29126 (N_29126,N_24817,N_26530);
or U29127 (N_29127,N_26680,N_25202);
or U29128 (N_29128,N_26743,N_26850);
or U29129 (N_29129,N_24016,N_24742);
nand U29130 (N_29130,N_26825,N_24066);
or U29131 (N_29131,N_25539,N_25205);
and U29132 (N_29132,N_25853,N_24060);
nor U29133 (N_29133,N_26217,N_25454);
and U29134 (N_29134,N_26848,N_24788);
or U29135 (N_29135,N_26066,N_25537);
xnor U29136 (N_29136,N_24620,N_25456);
nor U29137 (N_29137,N_25779,N_24705);
xnor U29138 (N_29138,N_25886,N_25855);
or U29139 (N_29139,N_26159,N_24449);
or U29140 (N_29140,N_25711,N_25125);
nor U29141 (N_29141,N_26375,N_25358);
or U29142 (N_29142,N_26862,N_26447);
nor U29143 (N_29143,N_25388,N_26538);
xnor U29144 (N_29144,N_25492,N_26248);
nand U29145 (N_29145,N_25290,N_26392);
and U29146 (N_29146,N_24537,N_25435);
or U29147 (N_29147,N_24331,N_24245);
or U29148 (N_29148,N_24421,N_25123);
or U29149 (N_29149,N_26039,N_25776);
and U29150 (N_29150,N_25198,N_26380);
nor U29151 (N_29151,N_25807,N_25291);
nand U29152 (N_29152,N_25502,N_26112);
nand U29153 (N_29153,N_25681,N_26433);
xnor U29154 (N_29154,N_25764,N_26222);
and U29155 (N_29155,N_25316,N_26434);
and U29156 (N_29156,N_25446,N_26883);
or U29157 (N_29157,N_25972,N_25511);
nand U29158 (N_29158,N_24280,N_24274);
or U29159 (N_29159,N_26911,N_26711);
nor U29160 (N_29160,N_25313,N_24606);
nor U29161 (N_29161,N_24234,N_24411);
nor U29162 (N_29162,N_25323,N_24289);
nand U29163 (N_29163,N_24905,N_26101);
nor U29164 (N_29164,N_24848,N_26377);
nand U29165 (N_29165,N_24289,N_25865);
or U29166 (N_29166,N_25789,N_24321);
nand U29167 (N_29167,N_25075,N_25589);
nor U29168 (N_29168,N_26428,N_26514);
xor U29169 (N_29169,N_26974,N_26908);
nor U29170 (N_29170,N_26236,N_25623);
and U29171 (N_29171,N_25850,N_26739);
xnor U29172 (N_29172,N_24436,N_26525);
and U29173 (N_29173,N_24532,N_24342);
nand U29174 (N_29174,N_24028,N_26233);
and U29175 (N_29175,N_25806,N_24408);
nand U29176 (N_29176,N_26173,N_24834);
nand U29177 (N_29177,N_26443,N_25914);
xor U29178 (N_29178,N_25379,N_24364);
and U29179 (N_29179,N_25683,N_24759);
or U29180 (N_29180,N_25739,N_26007);
xor U29181 (N_29181,N_24777,N_25182);
nor U29182 (N_29182,N_25483,N_26259);
nor U29183 (N_29183,N_25937,N_26400);
xor U29184 (N_29184,N_24740,N_24480);
nand U29185 (N_29185,N_26086,N_26142);
nand U29186 (N_29186,N_24523,N_24392);
xor U29187 (N_29187,N_25711,N_25485);
nor U29188 (N_29188,N_24060,N_24589);
or U29189 (N_29189,N_25064,N_24051);
nand U29190 (N_29190,N_24921,N_26388);
nor U29191 (N_29191,N_25464,N_26560);
and U29192 (N_29192,N_24751,N_24168);
nand U29193 (N_29193,N_25874,N_25309);
xor U29194 (N_29194,N_25516,N_26761);
xnor U29195 (N_29195,N_25493,N_24952);
nor U29196 (N_29196,N_25969,N_25196);
nand U29197 (N_29197,N_25915,N_26800);
nor U29198 (N_29198,N_24828,N_26269);
and U29199 (N_29199,N_24493,N_25537);
nand U29200 (N_29200,N_24258,N_26283);
nand U29201 (N_29201,N_24758,N_24324);
or U29202 (N_29202,N_26882,N_25935);
xnor U29203 (N_29203,N_26073,N_26680);
nor U29204 (N_29204,N_26564,N_25608);
nand U29205 (N_29205,N_25080,N_25548);
or U29206 (N_29206,N_24809,N_24954);
nor U29207 (N_29207,N_25974,N_24921);
nand U29208 (N_29208,N_24430,N_26245);
or U29209 (N_29209,N_24955,N_24551);
nor U29210 (N_29210,N_25957,N_26831);
nand U29211 (N_29211,N_25095,N_26604);
xor U29212 (N_29212,N_25827,N_26236);
or U29213 (N_29213,N_25405,N_25776);
nand U29214 (N_29214,N_24319,N_26211);
nor U29215 (N_29215,N_25591,N_26127);
nand U29216 (N_29216,N_26398,N_26765);
nand U29217 (N_29217,N_26302,N_25835);
nand U29218 (N_29218,N_26872,N_26855);
nor U29219 (N_29219,N_26473,N_25116);
nand U29220 (N_29220,N_25783,N_26635);
and U29221 (N_29221,N_26369,N_25598);
or U29222 (N_29222,N_24894,N_25385);
xor U29223 (N_29223,N_24940,N_24939);
nand U29224 (N_29224,N_24955,N_24712);
and U29225 (N_29225,N_25780,N_26368);
or U29226 (N_29226,N_24096,N_25507);
and U29227 (N_29227,N_24625,N_25055);
xor U29228 (N_29228,N_24047,N_25964);
xor U29229 (N_29229,N_24146,N_24005);
and U29230 (N_29230,N_24087,N_24022);
nor U29231 (N_29231,N_25034,N_25835);
and U29232 (N_29232,N_26782,N_24161);
nand U29233 (N_29233,N_24275,N_26522);
nand U29234 (N_29234,N_26607,N_25461);
nand U29235 (N_29235,N_26927,N_24854);
and U29236 (N_29236,N_24057,N_25704);
and U29237 (N_29237,N_24150,N_26736);
xor U29238 (N_29238,N_26027,N_24203);
nor U29239 (N_29239,N_26969,N_24687);
and U29240 (N_29240,N_26073,N_25596);
nor U29241 (N_29241,N_25860,N_26308);
nor U29242 (N_29242,N_25286,N_26691);
nor U29243 (N_29243,N_24636,N_24746);
and U29244 (N_29244,N_24446,N_26874);
and U29245 (N_29245,N_26125,N_24319);
xnor U29246 (N_29246,N_24296,N_26029);
nor U29247 (N_29247,N_26809,N_26581);
nand U29248 (N_29248,N_26095,N_26550);
xnor U29249 (N_29249,N_24553,N_24349);
or U29250 (N_29250,N_24693,N_25291);
nor U29251 (N_29251,N_25563,N_26770);
xor U29252 (N_29252,N_26009,N_24532);
or U29253 (N_29253,N_25919,N_24596);
and U29254 (N_29254,N_24524,N_25016);
and U29255 (N_29255,N_24914,N_24550);
xnor U29256 (N_29256,N_24000,N_26685);
or U29257 (N_29257,N_25389,N_25186);
nor U29258 (N_29258,N_25320,N_24124);
and U29259 (N_29259,N_25320,N_25030);
xor U29260 (N_29260,N_26219,N_26601);
nor U29261 (N_29261,N_24992,N_26580);
xor U29262 (N_29262,N_25387,N_24526);
nor U29263 (N_29263,N_25981,N_26205);
xor U29264 (N_29264,N_24973,N_26833);
nand U29265 (N_29265,N_25944,N_24245);
nand U29266 (N_29266,N_24961,N_24229);
or U29267 (N_29267,N_24902,N_26446);
xor U29268 (N_29268,N_26780,N_26810);
nor U29269 (N_29269,N_25509,N_25598);
xor U29270 (N_29270,N_24941,N_26332);
or U29271 (N_29271,N_25992,N_24086);
xnor U29272 (N_29272,N_24402,N_25267);
or U29273 (N_29273,N_26743,N_25692);
nor U29274 (N_29274,N_25367,N_26591);
or U29275 (N_29275,N_26008,N_24174);
xor U29276 (N_29276,N_25663,N_25524);
nor U29277 (N_29277,N_24176,N_24288);
nand U29278 (N_29278,N_25164,N_25769);
nand U29279 (N_29279,N_24880,N_25734);
or U29280 (N_29280,N_25489,N_26906);
nor U29281 (N_29281,N_24553,N_25294);
and U29282 (N_29282,N_26195,N_26286);
xnor U29283 (N_29283,N_26941,N_25897);
and U29284 (N_29284,N_24240,N_24812);
or U29285 (N_29285,N_26253,N_26622);
nand U29286 (N_29286,N_24086,N_24803);
xnor U29287 (N_29287,N_25337,N_24175);
and U29288 (N_29288,N_25137,N_24486);
and U29289 (N_29289,N_25185,N_24388);
xnor U29290 (N_29290,N_26202,N_26062);
or U29291 (N_29291,N_24957,N_25504);
xor U29292 (N_29292,N_25280,N_26906);
or U29293 (N_29293,N_24975,N_26043);
nor U29294 (N_29294,N_24891,N_26187);
or U29295 (N_29295,N_25752,N_26970);
or U29296 (N_29296,N_25415,N_26664);
or U29297 (N_29297,N_25246,N_25149);
nor U29298 (N_29298,N_26200,N_25521);
nand U29299 (N_29299,N_24478,N_26816);
xnor U29300 (N_29300,N_25738,N_25345);
or U29301 (N_29301,N_26918,N_25127);
nand U29302 (N_29302,N_26680,N_24385);
or U29303 (N_29303,N_26765,N_26108);
xor U29304 (N_29304,N_25141,N_25530);
or U29305 (N_29305,N_26797,N_26155);
nor U29306 (N_29306,N_26559,N_26274);
nand U29307 (N_29307,N_25649,N_24561);
xnor U29308 (N_29308,N_24797,N_26102);
nand U29309 (N_29309,N_26146,N_25576);
and U29310 (N_29310,N_25721,N_24735);
or U29311 (N_29311,N_26710,N_26768);
nand U29312 (N_29312,N_26715,N_26838);
nor U29313 (N_29313,N_25623,N_26256);
or U29314 (N_29314,N_26373,N_26043);
or U29315 (N_29315,N_26948,N_26060);
or U29316 (N_29316,N_25657,N_26876);
nor U29317 (N_29317,N_26763,N_24120);
or U29318 (N_29318,N_24343,N_24728);
nand U29319 (N_29319,N_26833,N_26541);
and U29320 (N_29320,N_26355,N_24959);
nand U29321 (N_29321,N_26026,N_26908);
nand U29322 (N_29322,N_24962,N_26376);
and U29323 (N_29323,N_26978,N_25640);
and U29324 (N_29324,N_26359,N_25930);
and U29325 (N_29325,N_25022,N_25727);
nor U29326 (N_29326,N_24622,N_26644);
xor U29327 (N_29327,N_24027,N_26507);
or U29328 (N_29328,N_24349,N_25293);
and U29329 (N_29329,N_26736,N_26745);
nor U29330 (N_29330,N_24304,N_25908);
or U29331 (N_29331,N_24280,N_24101);
and U29332 (N_29332,N_26509,N_26164);
or U29333 (N_29333,N_25712,N_25101);
or U29334 (N_29334,N_26408,N_24265);
nand U29335 (N_29335,N_26031,N_26960);
nor U29336 (N_29336,N_26316,N_24712);
nor U29337 (N_29337,N_26558,N_26513);
or U29338 (N_29338,N_24315,N_24312);
nand U29339 (N_29339,N_24921,N_25007);
and U29340 (N_29340,N_26731,N_25816);
nor U29341 (N_29341,N_26244,N_24577);
and U29342 (N_29342,N_25441,N_26157);
or U29343 (N_29343,N_26755,N_25495);
xnor U29344 (N_29344,N_25814,N_24297);
nor U29345 (N_29345,N_24058,N_26665);
nand U29346 (N_29346,N_25040,N_25266);
or U29347 (N_29347,N_25830,N_26338);
xor U29348 (N_29348,N_25795,N_25365);
or U29349 (N_29349,N_25206,N_26717);
xnor U29350 (N_29350,N_25545,N_25578);
xor U29351 (N_29351,N_24673,N_24940);
and U29352 (N_29352,N_26054,N_26255);
nand U29353 (N_29353,N_24682,N_24267);
and U29354 (N_29354,N_24182,N_26007);
or U29355 (N_29355,N_26873,N_24037);
nor U29356 (N_29356,N_24497,N_24893);
and U29357 (N_29357,N_26977,N_26669);
and U29358 (N_29358,N_26404,N_24682);
nand U29359 (N_29359,N_26317,N_26089);
and U29360 (N_29360,N_25530,N_25119);
nor U29361 (N_29361,N_26282,N_24862);
nor U29362 (N_29362,N_26294,N_24017);
nor U29363 (N_29363,N_24192,N_26975);
and U29364 (N_29364,N_26375,N_24729);
xor U29365 (N_29365,N_24648,N_26668);
nand U29366 (N_29366,N_24294,N_25852);
xnor U29367 (N_29367,N_25866,N_24156);
and U29368 (N_29368,N_24356,N_25110);
nor U29369 (N_29369,N_26966,N_26082);
nor U29370 (N_29370,N_26567,N_24285);
nand U29371 (N_29371,N_25470,N_24532);
nand U29372 (N_29372,N_26698,N_26888);
nor U29373 (N_29373,N_24887,N_25550);
xor U29374 (N_29374,N_25520,N_24086);
and U29375 (N_29375,N_24642,N_25056);
or U29376 (N_29376,N_25457,N_26771);
nand U29377 (N_29377,N_26724,N_24226);
nand U29378 (N_29378,N_25747,N_26896);
nand U29379 (N_29379,N_24211,N_25902);
nand U29380 (N_29380,N_25332,N_24471);
nor U29381 (N_29381,N_25023,N_26726);
nor U29382 (N_29382,N_24334,N_25650);
or U29383 (N_29383,N_25152,N_26392);
and U29384 (N_29384,N_25770,N_24060);
nand U29385 (N_29385,N_26523,N_25595);
nand U29386 (N_29386,N_25300,N_25067);
nand U29387 (N_29387,N_25262,N_26290);
nand U29388 (N_29388,N_26637,N_26131);
nor U29389 (N_29389,N_26098,N_25329);
nand U29390 (N_29390,N_25832,N_26760);
nor U29391 (N_29391,N_25661,N_25907);
or U29392 (N_29392,N_26691,N_25606);
nand U29393 (N_29393,N_24064,N_26722);
or U29394 (N_29394,N_25693,N_26110);
xor U29395 (N_29395,N_25247,N_25729);
or U29396 (N_29396,N_24170,N_25087);
xor U29397 (N_29397,N_24447,N_26380);
nand U29398 (N_29398,N_25278,N_25324);
or U29399 (N_29399,N_24716,N_25317);
or U29400 (N_29400,N_24362,N_26666);
nand U29401 (N_29401,N_24894,N_24946);
nor U29402 (N_29402,N_26656,N_26705);
nand U29403 (N_29403,N_26479,N_24515);
nor U29404 (N_29404,N_26687,N_25985);
nand U29405 (N_29405,N_25857,N_25442);
and U29406 (N_29406,N_25795,N_24017);
or U29407 (N_29407,N_26810,N_25896);
and U29408 (N_29408,N_25520,N_24658);
and U29409 (N_29409,N_25803,N_26843);
nor U29410 (N_29410,N_26285,N_26388);
and U29411 (N_29411,N_24629,N_24673);
xor U29412 (N_29412,N_26576,N_26757);
nand U29413 (N_29413,N_24467,N_25608);
nor U29414 (N_29414,N_24726,N_26328);
or U29415 (N_29415,N_24468,N_26696);
nor U29416 (N_29416,N_25553,N_26518);
or U29417 (N_29417,N_25352,N_26329);
nand U29418 (N_29418,N_26551,N_26879);
or U29419 (N_29419,N_24963,N_24663);
nand U29420 (N_29420,N_24655,N_24183);
nor U29421 (N_29421,N_26243,N_25229);
and U29422 (N_29422,N_25202,N_25749);
and U29423 (N_29423,N_25934,N_24507);
xnor U29424 (N_29424,N_24628,N_25632);
nand U29425 (N_29425,N_25623,N_25486);
xnor U29426 (N_29426,N_25686,N_26696);
nor U29427 (N_29427,N_25059,N_25624);
and U29428 (N_29428,N_25045,N_24313);
nand U29429 (N_29429,N_25868,N_26482);
or U29430 (N_29430,N_25413,N_26721);
nand U29431 (N_29431,N_26363,N_24842);
and U29432 (N_29432,N_24522,N_24594);
and U29433 (N_29433,N_25878,N_24749);
or U29434 (N_29434,N_25544,N_26926);
or U29435 (N_29435,N_24380,N_26188);
nor U29436 (N_29436,N_25948,N_24832);
or U29437 (N_29437,N_26704,N_24718);
nand U29438 (N_29438,N_24479,N_25744);
and U29439 (N_29439,N_25950,N_24516);
nand U29440 (N_29440,N_25018,N_24157);
or U29441 (N_29441,N_25019,N_25281);
or U29442 (N_29442,N_24932,N_24791);
and U29443 (N_29443,N_24472,N_26179);
nor U29444 (N_29444,N_25662,N_26748);
nor U29445 (N_29445,N_24258,N_25504);
or U29446 (N_29446,N_24209,N_25104);
and U29447 (N_29447,N_25775,N_24907);
nor U29448 (N_29448,N_25134,N_25951);
xnor U29449 (N_29449,N_25777,N_26468);
or U29450 (N_29450,N_24432,N_24318);
nor U29451 (N_29451,N_25199,N_25937);
or U29452 (N_29452,N_24916,N_25013);
or U29453 (N_29453,N_24479,N_26636);
xor U29454 (N_29454,N_24245,N_24237);
nor U29455 (N_29455,N_24639,N_24866);
nand U29456 (N_29456,N_25989,N_25149);
xor U29457 (N_29457,N_26613,N_26413);
nor U29458 (N_29458,N_24447,N_25788);
and U29459 (N_29459,N_24201,N_25532);
or U29460 (N_29460,N_24437,N_24323);
nor U29461 (N_29461,N_25655,N_25020);
and U29462 (N_29462,N_25847,N_26366);
nor U29463 (N_29463,N_26709,N_26165);
nor U29464 (N_29464,N_25941,N_26110);
nand U29465 (N_29465,N_24535,N_26089);
nor U29466 (N_29466,N_24580,N_26802);
xor U29467 (N_29467,N_24607,N_26125);
or U29468 (N_29468,N_26265,N_26160);
and U29469 (N_29469,N_25212,N_25842);
xor U29470 (N_29470,N_24894,N_26152);
xor U29471 (N_29471,N_26649,N_25421);
or U29472 (N_29472,N_25682,N_26822);
nand U29473 (N_29473,N_25502,N_25368);
and U29474 (N_29474,N_24980,N_26075);
and U29475 (N_29475,N_26336,N_24915);
nand U29476 (N_29476,N_26912,N_26106);
xnor U29477 (N_29477,N_26287,N_26097);
and U29478 (N_29478,N_26684,N_24376);
nor U29479 (N_29479,N_25283,N_24807);
or U29480 (N_29480,N_24977,N_24142);
nor U29481 (N_29481,N_24634,N_24010);
or U29482 (N_29482,N_25850,N_24740);
xor U29483 (N_29483,N_26344,N_26112);
and U29484 (N_29484,N_26758,N_25411);
or U29485 (N_29485,N_26220,N_24981);
and U29486 (N_29486,N_25288,N_26413);
nor U29487 (N_29487,N_24154,N_25034);
and U29488 (N_29488,N_24891,N_25215);
nand U29489 (N_29489,N_26448,N_26514);
nand U29490 (N_29490,N_24963,N_25645);
or U29491 (N_29491,N_24729,N_25857);
nand U29492 (N_29492,N_25192,N_24727);
or U29493 (N_29493,N_26758,N_24951);
xor U29494 (N_29494,N_24018,N_24578);
xor U29495 (N_29495,N_25592,N_24791);
and U29496 (N_29496,N_24091,N_24921);
nand U29497 (N_29497,N_25638,N_26605);
nor U29498 (N_29498,N_25991,N_26366);
and U29499 (N_29499,N_24295,N_26038);
nor U29500 (N_29500,N_24380,N_26207);
or U29501 (N_29501,N_26024,N_25368);
or U29502 (N_29502,N_25955,N_24875);
or U29503 (N_29503,N_25402,N_25908);
and U29504 (N_29504,N_26092,N_26196);
xor U29505 (N_29505,N_26477,N_25060);
nand U29506 (N_29506,N_25371,N_26599);
xor U29507 (N_29507,N_26009,N_24233);
and U29508 (N_29508,N_25213,N_26987);
or U29509 (N_29509,N_26215,N_26592);
xor U29510 (N_29510,N_24659,N_26516);
nor U29511 (N_29511,N_25725,N_26421);
and U29512 (N_29512,N_25023,N_24069);
and U29513 (N_29513,N_25264,N_25343);
and U29514 (N_29514,N_26538,N_26934);
xor U29515 (N_29515,N_26589,N_25263);
xnor U29516 (N_29516,N_25127,N_26028);
xor U29517 (N_29517,N_25594,N_25325);
xor U29518 (N_29518,N_24049,N_26884);
xor U29519 (N_29519,N_26776,N_25847);
or U29520 (N_29520,N_26013,N_25344);
xor U29521 (N_29521,N_24955,N_24097);
xnor U29522 (N_29522,N_26786,N_25886);
xnor U29523 (N_29523,N_25145,N_26583);
and U29524 (N_29524,N_26192,N_24862);
and U29525 (N_29525,N_24024,N_24398);
or U29526 (N_29526,N_24703,N_24255);
and U29527 (N_29527,N_24723,N_26977);
or U29528 (N_29528,N_24023,N_24876);
nor U29529 (N_29529,N_26861,N_25138);
nor U29530 (N_29530,N_26133,N_26773);
nor U29531 (N_29531,N_26687,N_24840);
nand U29532 (N_29532,N_26134,N_26929);
xnor U29533 (N_29533,N_24366,N_26044);
xor U29534 (N_29534,N_24619,N_24166);
xnor U29535 (N_29535,N_25292,N_26013);
and U29536 (N_29536,N_24036,N_25399);
or U29537 (N_29537,N_24857,N_24373);
xor U29538 (N_29538,N_26263,N_24029);
and U29539 (N_29539,N_24193,N_26313);
nor U29540 (N_29540,N_25358,N_26202);
and U29541 (N_29541,N_25975,N_26030);
nor U29542 (N_29542,N_26350,N_25709);
xnor U29543 (N_29543,N_24395,N_26105);
xor U29544 (N_29544,N_25446,N_25995);
nor U29545 (N_29545,N_24836,N_24569);
xor U29546 (N_29546,N_24520,N_25080);
xnor U29547 (N_29547,N_25282,N_24814);
nand U29548 (N_29548,N_26129,N_25689);
and U29549 (N_29549,N_26840,N_24752);
xor U29550 (N_29550,N_26019,N_24839);
nor U29551 (N_29551,N_25310,N_25765);
xor U29552 (N_29552,N_26544,N_25406);
or U29553 (N_29553,N_24466,N_26827);
and U29554 (N_29554,N_25160,N_25199);
xor U29555 (N_29555,N_26064,N_25964);
and U29556 (N_29556,N_25259,N_24538);
nor U29557 (N_29557,N_26817,N_25551);
and U29558 (N_29558,N_26781,N_25893);
nor U29559 (N_29559,N_25558,N_24474);
and U29560 (N_29560,N_26593,N_24255);
xnor U29561 (N_29561,N_26757,N_26333);
nand U29562 (N_29562,N_25322,N_24145);
or U29563 (N_29563,N_24821,N_24750);
or U29564 (N_29564,N_25182,N_24017);
or U29565 (N_29565,N_26803,N_26624);
xor U29566 (N_29566,N_26105,N_24038);
and U29567 (N_29567,N_26450,N_26385);
or U29568 (N_29568,N_26597,N_25260);
nand U29569 (N_29569,N_25508,N_24521);
or U29570 (N_29570,N_24312,N_26891);
and U29571 (N_29571,N_26486,N_26888);
or U29572 (N_29572,N_25329,N_24629);
and U29573 (N_29573,N_26148,N_24797);
and U29574 (N_29574,N_26094,N_26862);
xor U29575 (N_29575,N_26629,N_26080);
xor U29576 (N_29576,N_25449,N_24010);
xnor U29577 (N_29577,N_26052,N_25021);
or U29578 (N_29578,N_24760,N_25128);
nor U29579 (N_29579,N_26892,N_24572);
nand U29580 (N_29580,N_26186,N_24443);
xnor U29581 (N_29581,N_25211,N_25624);
xnor U29582 (N_29582,N_25587,N_25646);
nand U29583 (N_29583,N_24634,N_25438);
xnor U29584 (N_29584,N_25285,N_26372);
and U29585 (N_29585,N_26000,N_25388);
or U29586 (N_29586,N_26036,N_25730);
nor U29587 (N_29587,N_25885,N_26733);
xor U29588 (N_29588,N_25775,N_25168);
nand U29589 (N_29589,N_25582,N_25656);
nand U29590 (N_29590,N_24352,N_26209);
nor U29591 (N_29591,N_26456,N_25124);
nor U29592 (N_29592,N_24409,N_24992);
nor U29593 (N_29593,N_24461,N_25027);
or U29594 (N_29594,N_26082,N_25767);
and U29595 (N_29595,N_24291,N_24557);
or U29596 (N_29596,N_25691,N_26067);
xor U29597 (N_29597,N_24210,N_24321);
and U29598 (N_29598,N_26646,N_25458);
or U29599 (N_29599,N_26124,N_26697);
and U29600 (N_29600,N_26882,N_24001);
or U29601 (N_29601,N_26680,N_26190);
nand U29602 (N_29602,N_25561,N_26437);
nand U29603 (N_29603,N_25921,N_25312);
nor U29604 (N_29604,N_25482,N_24810);
or U29605 (N_29605,N_24356,N_26714);
and U29606 (N_29606,N_26212,N_26708);
and U29607 (N_29607,N_24485,N_25352);
and U29608 (N_29608,N_24038,N_25311);
xnor U29609 (N_29609,N_26619,N_26666);
nor U29610 (N_29610,N_25205,N_26269);
xnor U29611 (N_29611,N_24147,N_24626);
xor U29612 (N_29612,N_24057,N_24436);
xnor U29613 (N_29613,N_24437,N_24460);
and U29614 (N_29614,N_25362,N_26975);
nand U29615 (N_29615,N_26508,N_26635);
nor U29616 (N_29616,N_24544,N_24582);
nor U29617 (N_29617,N_25329,N_26149);
nor U29618 (N_29618,N_26830,N_25555);
nor U29619 (N_29619,N_24092,N_24368);
nand U29620 (N_29620,N_24813,N_24571);
or U29621 (N_29621,N_24300,N_26196);
nor U29622 (N_29622,N_24353,N_25435);
nor U29623 (N_29623,N_25054,N_25208);
nor U29624 (N_29624,N_24875,N_26344);
nand U29625 (N_29625,N_24384,N_25334);
or U29626 (N_29626,N_26807,N_26238);
nand U29627 (N_29627,N_24057,N_24765);
nor U29628 (N_29628,N_26815,N_24767);
nand U29629 (N_29629,N_26523,N_26345);
nor U29630 (N_29630,N_26180,N_26274);
xor U29631 (N_29631,N_25035,N_25087);
or U29632 (N_29632,N_25200,N_24388);
nand U29633 (N_29633,N_26345,N_24982);
nand U29634 (N_29634,N_26442,N_26993);
xnor U29635 (N_29635,N_25549,N_24046);
nor U29636 (N_29636,N_24555,N_26408);
nand U29637 (N_29637,N_24726,N_25346);
or U29638 (N_29638,N_24816,N_25038);
or U29639 (N_29639,N_26761,N_25617);
and U29640 (N_29640,N_24564,N_24626);
and U29641 (N_29641,N_24076,N_25630);
and U29642 (N_29642,N_26695,N_26530);
or U29643 (N_29643,N_26960,N_25583);
and U29644 (N_29644,N_24345,N_24982);
and U29645 (N_29645,N_24946,N_26122);
nand U29646 (N_29646,N_25016,N_26481);
nor U29647 (N_29647,N_25003,N_26631);
nand U29648 (N_29648,N_25521,N_25831);
xor U29649 (N_29649,N_25279,N_26384);
and U29650 (N_29650,N_24199,N_25848);
nand U29651 (N_29651,N_24143,N_25294);
nand U29652 (N_29652,N_24204,N_24636);
and U29653 (N_29653,N_25068,N_25143);
or U29654 (N_29654,N_25537,N_25563);
and U29655 (N_29655,N_25484,N_26142);
or U29656 (N_29656,N_25471,N_26245);
nor U29657 (N_29657,N_24043,N_24346);
xnor U29658 (N_29658,N_24201,N_25328);
and U29659 (N_29659,N_24280,N_25382);
nand U29660 (N_29660,N_26234,N_24529);
xor U29661 (N_29661,N_26235,N_25123);
nor U29662 (N_29662,N_24026,N_25232);
and U29663 (N_29663,N_25197,N_26631);
nor U29664 (N_29664,N_25320,N_24378);
and U29665 (N_29665,N_25336,N_25619);
nor U29666 (N_29666,N_26750,N_26984);
nand U29667 (N_29667,N_26180,N_26967);
xor U29668 (N_29668,N_25982,N_26442);
or U29669 (N_29669,N_26950,N_25714);
nand U29670 (N_29670,N_25970,N_24724);
xnor U29671 (N_29671,N_26137,N_26015);
nor U29672 (N_29672,N_26446,N_25966);
nand U29673 (N_29673,N_25229,N_24749);
nand U29674 (N_29674,N_26507,N_26036);
nor U29675 (N_29675,N_26706,N_26052);
nand U29676 (N_29676,N_24303,N_26022);
nand U29677 (N_29677,N_25719,N_24436);
nand U29678 (N_29678,N_24623,N_26993);
or U29679 (N_29679,N_26378,N_24921);
xor U29680 (N_29680,N_25305,N_26299);
or U29681 (N_29681,N_24993,N_26271);
nor U29682 (N_29682,N_24259,N_25681);
and U29683 (N_29683,N_25330,N_24620);
xor U29684 (N_29684,N_25063,N_26560);
nor U29685 (N_29685,N_25223,N_26023);
nor U29686 (N_29686,N_25774,N_24412);
nor U29687 (N_29687,N_26420,N_26970);
xnor U29688 (N_29688,N_25617,N_24692);
nor U29689 (N_29689,N_25218,N_26266);
nand U29690 (N_29690,N_25318,N_25050);
xor U29691 (N_29691,N_25280,N_25363);
nand U29692 (N_29692,N_25052,N_26635);
nor U29693 (N_29693,N_24789,N_25249);
nand U29694 (N_29694,N_26882,N_26175);
and U29695 (N_29695,N_25490,N_26873);
nor U29696 (N_29696,N_24315,N_24139);
and U29697 (N_29697,N_24576,N_24022);
nand U29698 (N_29698,N_25645,N_25711);
or U29699 (N_29699,N_25126,N_26668);
nor U29700 (N_29700,N_25610,N_25799);
nor U29701 (N_29701,N_24889,N_24958);
and U29702 (N_29702,N_25933,N_25671);
xnor U29703 (N_29703,N_26512,N_26062);
nor U29704 (N_29704,N_25849,N_24462);
xor U29705 (N_29705,N_24080,N_26846);
xnor U29706 (N_29706,N_26333,N_26004);
or U29707 (N_29707,N_24617,N_25421);
nand U29708 (N_29708,N_26116,N_24666);
and U29709 (N_29709,N_26981,N_24882);
and U29710 (N_29710,N_25902,N_26526);
or U29711 (N_29711,N_26665,N_24349);
or U29712 (N_29712,N_26000,N_26996);
nor U29713 (N_29713,N_25678,N_26555);
nand U29714 (N_29714,N_25737,N_25735);
and U29715 (N_29715,N_24902,N_26442);
xor U29716 (N_29716,N_25039,N_26461);
and U29717 (N_29717,N_26348,N_26009);
and U29718 (N_29718,N_24602,N_26982);
xor U29719 (N_29719,N_26467,N_24577);
and U29720 (N_29720,N_26478,N_26886);
and U29721 (N_29721,N_25209,N_25363);
xor U29722 (N_29722,N_24267,N_24439);
and U29723 (N_29723,N_25594,N_26426);
nand U29724 (N_29724,N_24123,N_24684);
and U29725 (N_29725,N_24332,N_25001);
nor U29726 (N_29726,N_25675,N_26662);
nand U29727 (N_29727,N_24849,N_24393);
nor U29728 (N_29728,N_24028,N_26149);
nor U29729 (N_29729,N_24690,N_25484);
xor U29730 (N_29730,N_25684,N_24111);
and U29731 (N_29731,N_24609,N_24288);
and U29732 (N_29732,N_25587,N_25619);
or U29733 (N_29733,N_24068,N_24305);
and U29734 (N_29734,N_26483,N_24106);
and U29735 (N_29735,N_26797,N_24597);
nor U29736 (N_29736,N_24167,N_26093);
or U29737 (N_29737,N_25039,N_26046);
nand U29738 (N_29738,N_24664,N_26604);
nor U29739 (N_29739,N_26590,N_24974);
nor U29740 (N_29740,N_24970,N_24556);
nand U29741 (N_29741,N_25982,N_26410);
nor U29742 (N_29742,N_26495,N_26129);
or U29743 (N_29743,N_24450,N_24673);
nand U29744 (N_29744,N_24644,N_24352);
and U29745 (N_29745,N_25385,N_26580);
or U29746 (N_29746,N_25865,N_24681);
xnor U29747 (N_29747,N_25480,N_26842);
nor U29748 (N_29748,N_25410,N_26119);
and U29749 (N_29749,N_25875,N_26685);
or U29750 (N_29750,N_25272,N_24108);
nor U29751 (N_29751,N_26210,N_24926);
xnor U29752 (N_29752,N_26291,N_26672);
or U29753 (N_29753,N_24813,N_24759);
nand U29754 (N_29754,N_26763,N_25168);
xor U29755 (N_29755,N_26070,N_24482);
xnor U29756 (N_29756,N_25391,N_25251);
nor U29757 (N_29757,N_24370,N_26007);
nor U29758 (N_29758,N_24423,N_26073);
xor U29759 (N_29759,N_26981,N_26791);
nor U29760 (N_29760,N_26972,N_24456);
and U29761 (N_29761,N_24103,N_25560);
nor U29762 (N_29762,N_26181,N_25246);
nand U29763 (N_29763,N_26721,N_26286);
or U29764 (N_29764,N_25566,N_26611);
or U29765 (N_29765,N_24272,N_26799);
nand U29766 (N_29766,N_26596,N_26747);
or U29767 (N_29767,N_25948,N_25334);
or U29768 (N_29768,N_26553,N_25270);
and U29769 (N_29769,N_24629,N_24815);
nor U29770 (N_29770,N_24030,N_25837);
xnor U29771 (N_29771,N_26397,N_26148);
xor U29772 (N_29772,N_26481,N_24460);
and U29773 (N_29773,N_26983,N_24994);
or U29774 (N_29774,N_25709,N_26272);
nor U29775 (N_29775,N_24435,N_25847);
or U29776 (N_29776,N_25390,N_24001);
xor U29777 (N_29777,N_26188,N_26289);
or U29778 (N_29778,N_26997,N_25756);
xnor U29779 (N_29779,N_26432,N_25240);
and U29780 (N_29780,N_24970,N_24329);
xor U29781 (N_29781,N_25561,N_26263);
or U29782 (N_29782,N_25698,N_24536);
and U29783 (N_29783,N_25123,N_24880);
or U29784 (N_29784,N_26329,N_25896);
nand U29785 (N_29785,N_24340,N_25421);
and U29786 (N_29786,N_26601,N_26446);
nand U29787 (N_29787,N_25013,N_24388);
or U29788 (N_29788,N_24692,N_24757);
or U29789 (N_29789,N_24625,N_26194);
nand U29790 (N_29790,N_26988,N_26851);
or U29791 (N_29791,N_25069,N_25771);
or U29792 (N_29792,N_24877,N_24739);
or U29793 (N_29793,N_25861,N_24074);
nor U29794 (N_29794,N_26096,N_25848);
nand U29795 (N_29795,N_24985,N_24286);
and U29796 (N_29796,N_25101,N_24723);
nand U29797 (N_29797,N_26215,N_26907);
and U29798 (N_29798,N_25077,N_24826);
and U29799 (N_29799,N_25186,N_24954);
and U29800 (N_29800,N_25984,N_26474);
and U29801 (N_29801,N_26729,N_25080);
nand U29802 (N_29802,N_24917,N_26176);
xor U29803 (N_29803,N_26222,N_24925);
and U29804 (N_29804,N_25013,N_26767);
nand U29805 (N_29805,N_24313,N_26048);
nor U29806 (N_29806,N_24029,N_25563);
xnor U29807 (N_29807,N_26749,N_24744);
xnor U29808 (N_29808,N_24663,N_25403);
and U29809 (N_29809,N_25311,N_26581);
nor U29810 (N_29810,N_26388,N_26275);
xnor U29811 (N_29811,N_25856,N_24399);
nor U29812 (N_29812,N_26565,N_24689);
or U29813 (N_29813,N_25163,N_26519);
or U29814 (N_29814,N_24992,N_24087);
xnor U29815 (N_29815,N_25241,N_26893);
xnor U29816 (N_29816,N_26732,N_25102);
or U29817 (N_29817,N_26841,N_26160);
xnor U29818 (N_29818,N_26316,N_24230);
nor U29819 (N_29819,N_24789,N_25833);
nand U29820 (N_29820,N_24765,N_26335);
and U29821 (N_29821,N_25469,N_25611);
nand U29822 (N_29822,N_26818,N_24797);
nand U29823 (N_29823,N_25691,N_26092);
or U29824 (N_29824,N_25517,N_26841);
or U29825 (N_29825,N_24424,N_26521);
nand U29826 (N_29826,N_26683,N_24492);
and U29827 (N_29827,N_25969,N_24477);
xnor U29828 (N_29828,N_26696,N_25837);
and U29829 (N_29829,N_26509,N_26992);
and U29830 (N_29830,N_24610,N_25432);
or U29831 (N_29831,N_26344,N_25955);
nand U29832 (N_29832,N_25250,N_24122);
or U29833 (N_29833,N_26357,N_24989);
nor U29834 (N_29834,N_25041,N_24240);
nor U29835 (N_29835,N_26378,N_25209);
xnor U29836 (N_29836,N_24498,N_25447);
nor U29837 (N_29837,N_25608,N_24942);
or U29838 (N_29838,N_26737,N_26185);
and U29839 (N_29839,N_26546,N_25180);
xnor U29840 (N_29840,N_25342,N_26219);
nand U29841 (N_29841,N_24808,N_26651);
nand U29842 (N_29842,N_26971,N_26340);
or U29843 (N_29843,N_26002,N_26172);
or U29844 (N_29844,N_24681,N_25052);
xor U29845 (N_29845,N_25244,N_24428);
and U29846 (N_29846,N_26670,N_26520);
nand U29847 (N_29847,N_24714,N_24604);
nor U29848 (N_29848,N_25251,N_25696);
xnor U29849 (N_29849,N_26001,N_25359);
and U29850 (N_29850,N_24951,N_25143);
nand U29851 (N_29851,N_24685,N_26292);
nor U29852 (N_29852,N_24017,N_26249);
nor U29853 (N_29853,N_24010,N_26592);
or U29854 (N_29854,N_24341,N_26224);
or U29855 (N_29855,N_26513,N_24626);
or U29856 (N_29856,N_26315,N_24990);
and U29857 (N_29857,N_24608,N_25162);
xor U29858 (N_29858,N_25652,N_26512);
nand U29859 (N_29859,N_24621,N_25895);
or U29860 (N_29860,N_24031,N_24132);
nor U29861 (N_29861,N_26563,N_25881);
and U29862 (N_29862,N_24978,N_26165);
nor U29863 (N_29863,N_25853,N_26637);
and U29864 (N_29864,N_25177,N_24341);
and U29865 (N_29865,N_25191,N_24948);
nand U29866 (N_29866,N_25043,N_24289);
nor U29867 (N_29867,N_25498,N_25394);
xor U29868 (N_29868,N_26898,N_24013);
nand U29869 (N_29869,N_26285,N_25060);
or U29870 (N_29870,N_25077,N_24979);
or U29871 (N_29871,N_26471,N_26594);
nor U29872 (N_29872,N_26609,N_24675);
and U29873 (N_29873,N_24239,N_25295);
nor U29874 (N_29874,N_26986,N_25309);
and U29875 (N_29875,N_24942,N_24110);
and U29876 (N_29876,N_26775,N_25933);
xor U29877 (N_29877,N_25152,N_26887);
xnor U29878 (N_29878,N_26823,N_24779);
nor U29879 (N_29879,N_26268,N_26940);
or U29880 (N_29880,N_24511,N_24143);
nand U29881 (N_29881,N_26941,N_26374);
nand U29882 (N_29882,N_24884,N_25926);
xor U29883 (N_29883,N_25740,N_26087);
and U29884 (N_29884,N_26265,N_26872);
nor U29885 (N_29885,N_25052,N_26211);
xor U29886 (N_29886,N_24693,N_26693);
or U29887 (N_29887,N_26078,N_26069);
nand U29888 (N_29888,N_25807,N_24672);
nand U29889 (N_29889,N_25129,N_24804);
nand U29890 (N_29890,N_25157,N_24178);
nand U29891 (N_29891,N_24768,N_26899);
xnor U29892 (N_29892,N_26515,N_26109);
xor U29893 (N_29893,N_25972,N_25914);
and U29894 (N_29894,N_25333,N_25113);
or U29895 (N_29895,N_26041,N_24738);
nand U29896 (N_29896,N_24341,N_24655);
and U29897 (N_29897,N_26116,N_25538);
and U29898 (N_29898,N_25836,N_25351);
nand U29899 (N_29899,N_25215,N_24346);
xor U29900 (N_29900,N_26493,N_24309);
nor U29901 (N_29901,N_25735,N_25961);
nor U29902 (N_29902,N_25341,N_26633);
xor U29903 (N_29903,N_24475,N_24296);
xor U29904 (N_29904,N_25124,N_24075);
nand U29905 (N_29905,N_24912,N_25632);
xor U29906 (N_29906,N_25798,N_26195);
nor U29907 (N_29907,N_25042,N_25015);
nor U29908 (N_29908,N_24652,N_24759);
or U29909 (N_29909,N_24294,N_24421);
nor U29910 (N_29910,N_25252,N_26931);
nor U29911 (N_29911,N_26350,N_24432);
and U29912 (N_29912,N_24223,N_24842);
and U29913 (N_29913,N_24079,N_26693);
or U29914 (N_29914,N_24702,N_25999);
or U29915 (N_29915,N_25711,N_26133);
nor U29916 (N_29916,N_25952,N_25042);
nor U29917 (N_29917,N_26696,N_25340);
nand U29918 (N_29918,N_24116,N_25490);
nor U29919 (N_29919,N_24926,N_24966);
nor U29920 (N_29920,N_25607,N_25319);
and U29921 (N_29921,N_24074,N_26412);
nand U29922 (N_29922,N_26336,N_25650);
or U29923 (N_29923,N_24516,N_26446);
xnor U29924 (N_29924,N_26484,N_24141);
and U29925 (N_29925,N_25457,N_24592);
nor U29926 (N_29926,N_25264,N_24515);
nand U29927 (N_29927,N_25324,N_25954);
or U29928 (N_29928,N_26845,N_26990);
nor U29929 (N_29929,N_24536,N_24379);
nand U29930 (N_29930,N_26443,N_26852);
or U29931 (N_29931,N_26870,N_26089);
xnor U29932 (N_29932,N_25920,N_26385);
nand U29933 (N_29933,N_26912,N_26983);
and U29934 (N_29934,N_25773,N_26841);
nor U29935 (N_29935,N_24721,N_25210);
xor U29936 (N_29936,N_26482,N_24592);
xnor U29937 (N_29937,N_26568,N_25262);
or U29938 (N_29938,N_26227,N_24347);
and U29939 (N_29939,N_25962,N_24686);
or U29940 (N_29940,N_24434,N_25003);
nor U29941 (N_29941,N_25532,N_25933);
nor U29942 (N_29942,N_24233,N_25394);
xnor U29943 (N_29943,N_25351,N_25891);
xnor U29944 (N_29944,N_24796,N_26602);
nor U29945 (N_29945,N_24351,N_24074);
xnor U29946 (N_29946,N_26426,N_24500);
nor U29947 (N_29947,N_24272,N_25922);
xor U29948 (N_29948,N_24503,N_25517);
or U29949 (N_29949,N_25653,N_24882);
nand U29950 (N_29950,N_25179,N_24868);
nand U29951 (N_29951,N_25205,N_24029);
and U29952 (N_29952,N_26344,N_25573);
nor U29953 (N_29953,N_26247,N_26262);
xor U29954 (N_29954,N_26110,N_24433);
and U29955 (N_29955,N_25699,N_24724);
nor U29956 (N_29956,N_26399,N_26281);
nor U29957 (N_29957,N_25468,N_25177);
xnor U29958 (N_29958,N_26236,N_25840);
xnor U29959 (N_29959,N_26435,N_25143);
nor U29960 (N_29960,N_25844,N_24375);
and U29961 (N_29961,N_26345,N_26267);
xor U29962 (N_29962,N_24910,N_25438);
nor U29963 (N_29963,N_24240,N_25876);
and U29964 (N_29964,N_24839,N_25058);
or U29965 (N_29965,N_25615,N_24981);
or U29966 (N_29966,N_25929,N_24627);
and U29967 (N_29967,N_25017,N_25637);
nor U29968 (N_29968,N_26644,N_26197);
nor U29969 (N_29969,N_26071,N_25708);
xor U29970 (N_29970,N_24999,N_24663);
nand U29971 (N_29971,N_24206,N_24116);
nand U29972 (N_29972,N_25626,N_26394);
or U29973 (N_29973,N_25963,N_25076);
nand U29974 (N_29974,N_26786,N_25211);
nor U29975 (N_29975,N_26191,N_26584);
nor U29976 (N_29976,N_24484,N_25622);
nor U29977 (N_29977,N_24722,N_25971);
nor U29978 (N_29978,N_24656,N_25299);
nor U29979 (N_29979,N_24484,N_24703);
nand U29980 (N_29980,N_24195,N_24462);
or U29981 (N_29981,N_25690,N_24716);
or U29982 (N_29982,N_26201,N_26714);
and U29983 (N_29983,N_25229,N_26642);
and U29984 (N_29984,N_26359,N_24542);
xor U29985 (N_29985,N_25519,N_24379);
nor U29986 (N_29986,N_24469,N_26949);
xnor U29987 (N_29987,N_25227,N_25095);
nor U29988 (N_29988,N_26972,N_25126);
xor U29989 (N_29989,N_26970,N_25512);
or U29990 (N_29990,N_24795,N_24802);
xnor U29991 (N_29991,N_25631,N_24177);
or U29992 (N_29992,N_26731,N_26877);
nor U29993 (N_29993,N_26371,N_24081);
nand U29994 (N_29994,N_25347,N_24334);
or U29995 (N_29995,N_24388,N_24120);
xnor U29996 (N_29996,N_25547,N_24479);
or U29997 (N_29997,N_25658,N_25145);
and U29998 (N_29998,N_24597,N_24515);
nand U29999 (N_29999,N_24239,N_26147);
and UO_0 (O_0,N_27510,N_28039);
or UO_1 (O_1,N_29021,N_28523);
xor UO_2 (O_2,N_29009,N_28483);
or UO_3 (O_3,N_28732,N_29340);
or UO_4 (O_4,N_29850,N_27972);
xor UO_5 (O_5,N_29064,N_28647);
or UO_6 (O_6,N_28591,N_28715);
and UO_7 (O_7,N_29041,N_29610);
nor UO_8 (O_8,N_29981,N_29651);
and UO_9 (O_9,N_28883,N_27818);
nor UO_10 (O_10,N_27762,N_29298);
and UO_11 (O_11,N_28313,N_28756);
xor UO_12 (O_12,N_29055,N_28652);
nand UO_13 (O_13,N_28747,N_29915);
xnor UO_14 (O_14,N_29505,N_27354);
xor UO_15 (O_15,N_29276,N_29986);
and UO_16 (O_16,N_29988,N_27504);
and UO_17 (O_17,N_27142,N_27618);
and UO_18 (O_18,N_29196,N_28571);
and UO_19 (O_19,N_29702,N_27473);
xor UO_20 (O_20,N_28551,N_27283);
xor UO_21 (O_21,N_27434,N_28418);
xnor UO_22 (O_22,N_27946,N_27969);
nor UO_23 (O_23,N_28734,N_29176);
nor UO_24 (O_24,N_29096,N_28504);
and UO_25 (O_25,N_29539,N_29907);
or UO_26 (O_26,N_27833,N_28339);
and UO_27 (O_27,N_27140,N_27882);
or UO_28 (O_28,N_29343,N_27416);
and UO_29 (O_29,N_29679,N_29958);
xor UO_30 (O_30,N_28770,N_29730);
or UO_31 (O_31,N_29297,N_28806);
and UO_32 (O_32,N_27633,N_27942);
nand UO_33 (O_33,N_29594,N_29857);
xor UO_34 (O_34,N_29847,N_29131);
nor UO_35 (O_35,N_29127,N_29576);
xnor UO_36 (O_36,N_27229,N_28998);
xor UO_37 (O_37,N_27502,N_27739);
nand UO_38 (O_38,N_27317,N_29320);
or UO_39 (O_39,N_28866,N_29919);
nand UO_40 (O_40,N_27609,N_29295);
xnor UO_41 (O_41,N_29444,N_29689);
and UO_42 (O_42,N_27951,N_29338);
xnor UO_43 (O_43,N_29564,N_28073);
nand UO_44 (O_44,N_28091,N_28423);
or UO_45 (O_45,N_27993,N_27826);
and UO_46 (O_46,N_27567,N_27742);
xor UO_47 (O_47,N_27613,N_27412);
nor UO_48 (O_48,N_27827,N_28597);
or UO_49 (O_49,N_29242,N_28171);
xnor UO_50 (O_50,N_27121,N_29043);
xor UO_51 (O_51,N_29912,N_28297);
nor UO_52 (O_52,N_28559,N_29114);
nor UO_53 (O_53,N_28102,N_27281);
xnor UO_54 (O_54,N_28582,N_27374);
nand UO_55 (O_55,N_29223,N_27278);
and UO_56 (O_56,N_27484,N_27053);
nor UO_57 (O_57,N_29992,N_27854);
or UO_58 (O_58,N_28285,N_28244);
xor UO_59 (O_59,N_29602,N_29659);
xor UO_60 (O_60,N_29721,N_28872);
and UO_61 (O_61,N_28728,N_29120);
xnor UO_62 (O_62,N_28749,N_27287);
and UO_63 (O_63,N_29948,N_29140);
or UO_64 (O_64,N_27883,N_27390);
xor UO_65 (O_65,N_27286,N_28602);
and UO_66 (O_66,N_28304,N_29648);
nor UO_67 (O_67,N_28019,N_27380);
xnor UO_68 (O_68,N_29169,N_28381);
nand UO_69 (O_69,N_27839,N_29201);
and UO_70 (O_70,N_28624,N_29759);
and UO_71 (O_71,N_27204,N_27789);
and UO_72 (O_72,N_27713,N_27772);
or UO_73 (O_73,N_28942,N_29813);
or UO_74 (O_74,N_27940,N_27754);
xor UO_75 (O_75,N_27632,N_28158);
nor UO_76 (O_76,N_27903,N_27989);
xnor UO_77 (O_77,N_28511,N_28917);
and UO_78 (O_78,N_27312,N_29612);
and UO_79 (O_79,N_27191,N_27125);
and UO_80 (O_80,N_29931,N_29153);
and UO_81 (O_81,N_28393,N_27824);
or UO_82 (O_82,N_28710,N_29553);
nand UO_83 (O_83,N_27999,N_28856);
xnor UO_84 (O_84,N_28242,N_28277);
and UO_85 (O_85,N_27406,N_28167);
xnor UO_86 (O_86,N_29381,N_28996);
xnor UO_87 (O_87,N_28676,N_27072);
nand UO_88 (O_88,N_28343,N_29882);
nor UO_89 (O_89,N_29229,N_29782);
and UO_90 (O_90,N_27738,N_28447);
nor UO_91 (O_91,N_28601,N_27345);
nor UO_92 (O_92,N_29846,N_28028);
and UO_93 (O_93,N_28805,N_29536);
nor UO_94 (O_94,N_27667,N_29371);
nor UO_95 (O_95,N_27049,N_27555);
nand UO_96 (O_96,N_28508,N_28605);
nor UO_97 (O_97,N_29160,N_29796);
nor UO_98 (O_98,N_28411,N_28791);
nor UO_99 (O_99,N_29439,N_29415);
or UO_100 (O_100,N_27933,N_27367);
or UO_101 (O_101,N_29109,N_28684);
nor UO_102 (O_102,N_27780,N_27112);
xnor UO_103 (O_103,N_29188,N_28045);
nor UO_104 (O_104,N_29815,N_29657);
or UO_105 (O_105,N_29995,N_29750);
nor UO_106 (O_106,N_28301,N_27706);
xnor UO_107 (O_107,N_28214,N_28786);
xor UO_108 (O_108,N_29472,N_29511);
and UO_109 (O_109,N_29218,N_28930);
xor UO_110 (O_110,N_28207,N_27359);
nand UO_111 (O_111,N_28925,N_28215);
nor UO_112 (O_112,N_29943,N_27261);
or UO_113 (O_113,N_27990,N_29577);
nor UO_114 (O_114,N_29865,N_27619);
or UO_115 (O_115,N_29829,N_27331);
nand UO_116 (O_116,N_28595,N_29888);
xor UO_117 (O_117,N_27055,N_29823);
and UO_118 (O_118,N_27977,N_29929);
nor UO_119 (O_119,N_29962,N_27936);
and UO_120 (O_120,N_29524,N_27321);
or UO_121 (O_121,N_29037,N_29321);
nand UO_122 (O_122,N_29604,N_28357);
or UO_123 (O_123,N_27277,N_27436);
nor UO_124 (O_124,N_28132,N_27100);
and UO_125 (O_125,N_27135,N_28789);
and UO_126 (O_126,N_29640,N_27469);
and UO_127 (O_127,N_28702,N_27293);
xnor UO_128 (O_128,N_27298,N_27852);
and UO_129 (O_129,N_27651,N_27997);
xor UO_130 (O_130,N_29296,N_27604);
nor UO_131 (O_131,N_29938,N_28193);
nand UO_132 (O_132,N_29325,N_27703);
and UO_133 (O_133,N_27655,N_27902);
nor UO_134 (O_134,N_27475,N_28034);
or UO_135 (O_135,N_29151,N_28318);
xor UO_136 (O_136,N_29706,N_29362);
or UO_137 (O_137,N_29384,N_29336);
nand UO_138 (O_138,N_27147,N_28468);
and UO_139 (O_139,N_28562,N_28858);
xnor UO_140 (O_140,N_28644,N_28363);
and UO_141 (O_141,N_28754,N_27245);
nor UO_142 (O_142,N_29906,N_27673);
and UO_143 (O_143,N_27167,N_29061);
or UO_144 (O_144,N_27478,N_29805);
xnor UO_145 (O_145,N_28076,N_27560);
or UO_146 (O_146,N_29816,N_29356);
xnor UO_147 (O_147,N_27953,N_27527);
nand UO_148 (O_148,N_29693,N_29313);
nand UO_149 (O_149,N_28181,N_29082);
nand UO_150 (O_150,N_27741,N_29486);
nand UO_151 (O_151,N_28894,N_28051);
or UO_152 (O_152,N_29467,N_29567);
nand UO_153 (O_153,N_27526,N_28315);
nand UO_154 (O_154,N_27222,N_28914);
nor UO_155 (O_155,N_27230,N_27982);
nor UO_156 (O_156,N_28573,N_27077);
and UO_157 (O_157,N_28809,N_29044);
or UO_158 (O_158,N_27348,N_28302);
or UO_159 (O_159,N_27492,N_28299);
and UO_160 (O_160,N_27728,N_29790);
xor UO_161 (O_161,N_29345,N_28906);
xor UO_162 (O_162,N_27155,N_27482);
or UO_163 (O_163,N_27404,N_29433);
nor UO_164 (O_164,N_27507,N_27929);
xnor UO_165 (O_165,N_28609,N_27564);
nor UO_166 (O_166,N_29435,N_27980);
nand UO_167 (O_167,N_28712,N_29093);
and UO_168 (O_168,N_27524,N_29214);
nand UO_169 (O_169,N_27102,N_27097);
and UO_170 (O_170,N_29589,N_28837);
xor UO_171 (O_171,N_28953,N_27377);
nand UO_172 (O_172,N_28482,N_29423);
nand UO_173 (O_173,N_28638,N_27050);
or UO_174 (O_174,N_29330,N_28096);
nand UO_175 (O_175,N_27038,N_29068);
xor UO_176 (O_176,N_28216,N_29828);
and UO_177 (O_177,N_27921,N_28918);
xor UO_178 (O_178,N_28373,N_27584);
nor UO_179 (O_179,N_27640,N_27376);
xnor UO_180 (O_180,N_28556,N_27546);
and UO_181 (O_181,N_28135,N_27722);
nand UO_182 (O_182,N_27361,N_29278);
and UO_183 (O_183,N_27771,N_29143);
nor UO_184 (O_184,N_29848,N_29440);
nor UO_185 (O_185,N_29746,N_28099);
and UO_186 (O_186,N_28531,N_28070);
nor UO_187 (O_187,N_27319,N_29102);
nand UO_188 (O_188,N_27547,N_28913);
nand UO_189 (O_189,N_27196,N_29489);
nand UO_190 (O_190,N_29797,N_28166);
or UO_191 (O_191,N_29798,N_27681);
or UO_192 (O_192,N_28966,N_27817);
and UO_193 (O_193,N_29243,N_27645);
or UO_194 (O_194,N_29711,N_27508);
nor UO_195 (O_195,N_29953,N_29185);
or UO_196 (O_196,N_28127,N_28397);
nand UO_197 (O_197,N_28820,N_29993);
and UO_198 (O_198,N_28265,N_27694);
and UO_199 (O_199,N_28170,N_27787);
nor UO_200 (O_200,N_28103,N_28148);
xor UO_201 (O_201,N_28328,N_29255);
xor UO_202 (O_202,N_28500,N_27840);
nor UO_203 (O_203,N_28368,N_28125);
nand UO_204 (O_204,N_28143,N_28367);
and UO_205 (O_205,N_27616,N_27923);
nor UO_206 (O_206,N_27012,N_27160);
xor UO_207 (O_207,N_29890,N_28063);
or UO_208 (O_208,N_27201,N_29292);
nor UO_209 (O_209,N_29033,N_28420);
xnor UO_210 (O_210,N_28570,N_29507);
nand UO_211 (O_211,N_27540,N_28832);
or UO_212 (O_212,N_29838,N_29914);
and UO_213 (O_213,N_28341,N_28566);
nor UO_214 (O_214,N_29720,N_27601);
xnor UO_215 (O_215,N_28290,N_27005);
nor UO_216 (O_216,N_28174,N_28100);
nor UO_217 (O_217,N_29527,N_28704);
xnor UO_218 (O_218,N_27864,N_27543);
or UO_219 (O_219,N_28067,N_28741);
xnor UO_220 (O_220,N_29603,N_27476);
nor UO_221 (O_221,N_29053,N_29944);
or UO_222 (O_222,N_29119,N_29479);
and UO_223 (O_223,N_28776,N_27426);
or UO_224 (O_224,N_27028,N_28812);
and UO_225 (O_225,N_29641,N_28399);
xnor UO_226 (O_226,N_29462,N_28678);
and UO_227 (O_227,N_28928,N_27205);
and UO_228 (O_228,N_28187,N_28830);
and UO_229 (O_229,N_27731,N_29876);
and UO_230 (O_230,N_29608,N_29949);
or UO_231 (O_231,N_29743,N_29245);
xor UO_232 (O_232,N_27967,N_28921);
nor UO_233 (O_233,N_27985,N_27075);
nand UO_234 (O_234,N_28853,N_29581);
nand UO_235 (O_235,N_28105,N_27806);
nand UO_236 (O_236,N_28435,N_27291);
nor UO_237 (O_237,N_27627,N_28616);
xnor UO_238 (O_238,N_29360,N_27580);
or UO_239 (O_239,N_29474,N_28464);
nand UO_240 (O_240,N_29509,N_28873);
nand UO_241 (O_241,N_28669,N_29510);
xor UO_242 (O_242,N_28311,N_29309);
or UO_243 (O_243,N_28247,N_29911);
xnor UO_244 (O_244,N_28842,N_29873);
xnor UO_245 (O_245,N_27491,N_27411);
xor UO_246 (O_246,N_29476,N_27232);
nor UO_247 (O_247,N_29725,N_28692);
or UO_248 (O_248,N_28623,N_29565);
xor UO_249 (O_249,N_28541,N_29046);
nor UO_250 (O_250,N_27581,N_28845);
nor UO_251 (O_251,N_28092,N_28807);
nor UO_252 (O_252,N_27332,N_28200);
or UO_253 (O_253,N_27170,N_28991);
or UO_254 (O_254,N_28753,N_28862);
xor UO_255 (O_255,N_27586,N_27877);
nand UO_256 (O_256,N_27193,N_29773);
nand UO_257 (O_257,N_28267,N_28436);
or UO_258 (O_258,N_27221,N_29606);
or UO_259 (O_259,N_27151,N_27895);
or UO_260 (O_260,N_28658,N_27335);
nand UO_261 (O_261,N_28748,N_28186);
xnor UO_262 (O_262,N_28033,N_27407);
xor UO_263 (O_263,N_29686,N_28321);
nor UO_264 (O_264,N_29187,N_28960);
nor UO_265 (O_265,N_27711,N_27156);
nand UO_266 (O_266,N_29585,N_27884);
xor UO_267 (O_267,N_29056,N_29443);
nor UO_268 (O_268,N_27626,N_27941);
nand UO_269 (O_269,N_29729,N_29060);
xor UO_270 (O_270,N_29379,N_28564);
nand UO_271 (O_271,N_28988,N_27369);
or UO_272 (O_272,N_27860,N_29395);
nand UO_273 (O_273,N_28861,N_28160);
nor UO_274 (O_274,N_27401,N_29791);
nor UO_275 (O_275,N_29801,N_28516);
nand UO_276 (O_276,N_28956,N_29566);
xor UO_277 (O_277,N_29783,N_27347);
and UO_278 (O_278,N_28633,N_29735);
nor UO_279 (O_279,N_29979,N_29206);
xor UO_280 (O_280,N_28413,N_28173);
and UO_281 (O_281,N_28314,N_27386);
and UO_282 (O_282,N_28698,N_27919);
and UO_283 (O_283,N_29233,N_28263);
or UO_284 (O_284,N_28926,N_27957);
and UO_285 (O_285,N_28934,N_29437);
nand UO_286 (O_286,N_29353,N_27018);
nor UO_287 (O_287,N_28162,N_28876);
or UO_288 (O_288,N_27509,N_28241);
or UO_289 (O_289,N_27814,N_29818);
or UO_290 (O_290,N_27594,N_27538);
xor UO_291 (O_291,N_27449,N_28625);
and UO_292 (O_292,N_27966,N_29372);
nor UO_293 (O_293,N_28911,N_28117);
or UO_294 (O_294,N_28046,N_27668);
xor UO_295 (O_295,N_27719,N_28032);
nor UO_296 (O_296,N_28249,N_29552);
nor UO_297 (O_297,N_29727,N_27863);
xnor UO_298 (O_298,N_29035,N_28533);
nor UO_299 (O_299,N_28642,N_29207);
nor UO_300 (O_300,N_29701,N_27529);
and UO_301 (O_301,N_27216,N_29349);
or UO_302 (O_302,N_29067,N_29925);
nor UO_303 (O_303,N_28498,N_27745);
nor UO_304 (O_304,N_29312,N_29972);
and UO_305 (O_305,N_28177,N_28686);
nand UO_306 (O_306,N_27709,N_28355);
nor UO_307 (O_307,N_29316,N_28048);
and UO_308 (O_308,N_28963,N_27682);
or UO_309 (O_309,N_27753,N_27887);
nor UO_310 (O_310,N_29685,N_29090);
or UO_311 (O_311,N_28058,N_29454);
nor UO_312 (O_312,N_28864,N_29652);
xnor UO_313 (O_313,N_29083,N_28746);
and UO_314 (O_314,N_27777,N_27625);
nor UO_315 (O_315,N_27382,N_28385);
or UO_316 (O_316,N_28643,N_29677);
or UO_317 (O_317,N_29387,N_27458);
xor UO_318 (O_318,N_29731,N_27384);
or UO_319 (O_319,N_28990,N_28544);
or UO_320 (O_320,N_28600,N_29238);
nor UO_321 (O_321,N_27774,N_29352);
nor UO_322 (O_322,N_28524,N_29665);
and UO_323 (O_323,N_27341,N_28026);
and UO_324 (O_324,N_28316,N_27794);
and UO_325 (O_325,N_28675,N_28717);
xor UO_326 (O_326,N_28414,N_28374);
nor UO_327 (O_327,N_29253,N_28222);
and UO_328 (O_328,N_28952,N_27130);
and UO_329 (O_329,N_29990,N_27062);
nand UO_330 (O_330,N_28361,N_27336);
xnor UO_331 (O_331,N_27083,N_27006);
and UO_332 (O_332,N_29582,N_29583);
or UO_333 (O_333,N_28164,N_27074);
and UO_334 (O_334,N_27260,N_27172);
and UO_335 (O_335,N_29817,N_28887);
xor UO_336 (O_336,N_29942,N_27263);
and UO_337 (O_337,N_28064,N_29249);
nand UO_338 (O_338,N_28388,N_29441);
or UO_339 (O_339,N_29103,N_28350);
and UO_340 (O_340,N_28788,N_29259);
nand UO_341 (O_341,N_28172,N_28787);
nand UO_342 (O_342,N_29742,N_29241);
xnor UO_343 (O_343,N_27450,N_27605);
nand UO_344 (O_344,N_28632,N_29767);
and UO_345 (O_345,N_27497,N_28804);
nand UO_346 (O_346,N_27391,N_27836);
xnor UO_347 (O_347,N_27733,N_27813);
xnor UO_348 (O_348,N_29300,N_28446);
or UO_349 (O_349,N_29057,N_29733);
or UO_350 (O_350,N_27243,N_28936);
nand UO_351 (O_351,N_29363,N_27356);
nand UO_352 (O_352,N_29804,N_29947);
and UO_353 (O_353,N_29048,N_29521);
or UO_354 (O_354,N_27025,N_27849);
or UO_355 (O_355,N_28855,N_28257);
nor UO_356 (O_356,N_27421,N_29718);
nor UO_357 (O_357,N_29770,N_29787);
nor UO_358 (O_358,N_27660,N_28922);
or UO_359 (O_359,N_29551,N_29460);
nand UO_360 (O_360,N_29264,N_29409);
and UO_361 (O_361,N_27435,N_27402);
or UO_362 (O_362,N_29753,N_28395);
xor UO_363 (O_363,N_28425,N_27965);
nand UO_364 (O_364,N_28613,N_27051);
nor UO_365 (O_365,N_28370,N_27577);
nand UO_366 (O_366,N_27646,N_28098);
and UO_367 (O_367,N_28543,N_28795);
and UO_368 (O_368,N_29323,N_29200);
nor UO_369 (O_369,N_27381,N_29869);
or UO_370 (O_370,N_29755,N_28443);
and UO_371 (O_371,N_27372,N_28226);
nor UO_372 (O_372,N_28722,N_27512);
and UO_373 (O_373,N_27858,N_27859);
xor UO_374 (O_374,N_28324,N_27415);
and UO_375 (O_375,N_29715,N_28975);
nor UO_376 (O_376,N_28358,N_28416);
or UO_377 (O_377,N_29210,N_29646);
nand UO_378 (O_378,N_27506,N_29649);
or UO_379 (O_379,N_28954,N_28586);
xnor UO_380 (O_380,N_27375,N_28774);
nor UO_381 (O_381,N_29724,N_28920);
nor UO_382 (O_382,N_28977,N_27750);
or UO_383 (O_383,N_27596,N_29311);
nor UO_384 (O_384,N_28518,N_27477);
xnor UO_385 (O_385,N_28775,N_27187);
nor UO_386 (O_386,N_28352,N_27650);
nor UO_387 (O_387,N_27893,N_29969);
nand UO_388 (O_388,N_29453,N_27108);
xnor UO_389 (O_389,N_29705,N_28945);
nor UO_390 (O_390,N_28283,N_28421);
xnor UO_391 (O_391,N_29645,N_28036);
or UO_392 (O_392,N_27471,N_29698);
or UO_393 (O_393,N_28535,N_28122);
xor UO_394 (O_394,N_29156,N_27315);
xor UO_395 (O_395,N_29588,N_28107);
nand UO_396 (O_396,N_29690,N_29910);
nor UO_397 (O_397,N_29483,N_28427);
nand UO_398 (O_398,N_28915,N_29824);
and UO_399 (O_399,N_27498,N_28965);
nand UO_400 (O_400,N_27240,N_29076);
nor UO_401 (O_401,N_27909,N_29244);
nand UO_402 (O_402,N_27644,N_27761);
or UO_403 (O_403,N_29547,N_28950);
nor UO_404 (O_404,N_28927,N_27290);
nor UO_405 (O_405,N_29182,N_27368);
and UO_406 (O_406,N_29936,N_27330);
xor UO_407 (O_407,N_27662,N_28197);
or UO_408 (O_408,N_28041,N_27505);
and UO_409 (O_409,N_29215,N_27178);
nand UO_410 (O_410,N_27314,N_27521);
nor UO_411 (O_411,N_29870,N_28345);
xnor UO_412 (O_412,N_27885,N_29028);
nand UO_413 (O_413,N_29470,N_27614);
xnor UO_414 (O_414,N_27360,N_28583);
xor UO_415 (O_415,N_29175,N_29161);
nand UO_416 (O_416,N_27173,N_28163);
or UO_417 (O_417,N_29157,N_28506);
nand UO_418 (O_418,N_29933,N_29403);
or UO_419 (O_419,N_29261,N_27743);
nand UO_420 (O_420,N_28889,N_28069);
nor UO_421 (O_421,N_28394,N_28923);
xnor UO_422 (O_422,N_29416,N_29534);
and UO_423 (O_423,N_27755,N_29851);
and UO_424 (O_424,N_29811,N_28386);
and UO_425 (O_425,N_29456,N_27163);
or UO_426 (O_426,N_28580,N_29913);
and UO_427 (O_427,N_27866,N_28094);
nor UO_428 (O_428,N_29568,N_28621);
or UO_429 (O_429,N_27091,N_28007);
nor UO_430 (O_430,N_28310,N_27448);
nand UO_431 (O_431,N_27064,N_27530);
nor UO_432 (O_432,N_27392,N_29898);
nand UO_433 (O_433,N_29579,N_28588);
or UO_434 (O_434,N_27621,N_27769);
nand UO_435 (O_435,N_29973,N_28880);
nor UO_436 (O_436,N_27158,N_29736);
and UO_437 (O_437,N_29726,N_29704);
and UO_438 (O_438,N_29573,N_28834);
or UO_439 (O_439,N_27904,N_29142);
or UO_440 (O_440,N_28690,N_28472);
nor UO_441 (O_441,N_28138,N_27566);
nand UO_442 (O_442,N_27723,N_27259);
xor UO_443 (O_443,N_27549,N_27623);
nor UO_444 (O_444,N_29110,N_28821);
and UO_445 (O_445,N_29054,N_29283);
nor UO_446 (O_446,N_29199,N_29655);
nor UO_447 (O_447,N_27144,N_28037);
nor UO_448 (O_448,N_29130,N_28453);
xor UO_449 (O_449,N_29100,N_27974);
nand UO_450 (O_450,N_27831,N_28088);
nand UO_451 (O_451,N_29637,N_29830);
or UO_452 (O_452,N_28294,N_28874);
and UO_453 (O_453,N_28617,N_27154);
and UO_454 (O_454,N_29978,N_29291);
nand UO_455 (O_455,N_27052,N_29985);
and UO_456 (O_456,N_29596,N_28881);
xor UO_457 (O_457,N_28799,N_27848);
nand UO_458 (O_458,N_29508,N_27013);
or UO_459 (O_459,N_28090,N_28626);
nor UO_460 (O_460,N_27307,N_28841);
nor UO_461 (O_461,N_29181,N_27945);
nand UO_462 (O_462,N_28256,N_29485);
or UO_463 (O_463,N_29920,N_29469);
nor UO_464 (O_464,N_29112,N_28455);
nand UO_465 (O_465,N_27656,N_27034);
nor UO_466 (O_466,N_27759,N_29827);
nand UO_467 (O_467,N_28180,N_29417);
and UO_468 (O_468,N_28179,N_27019);
nand UO_469 (O_469,N_29688,N_28797);
nor UO_470 (O_470,N_29557,N_29744);
or UO_471 (O_471,N_27846,N_27862);
nor UO_472 (O_472,N_28085,N_29964);
or UO_473 (O_473,N_27608,N_28015);
and UO_474 (O_474,N_29436,N_29662);
or UO_475 (O_475,N_29516,N_28228);
nand UO_476 (O_476,N_28232,N_27054);
xnor UO_477 (O_477,N_27791,N_27732);
nand UO_478 (O_478,N_29871,N_29051);
xor UO_479 (O_479,N_28452,N_27907);
nand UO_480 (O_480,N_27023,N_29197);
nor UO_481 (O_481,N_28970,N_29438);
nand UO_482 (O_482,N_28599,N_29808);
nor UO_483 (O_483,N_27462,N_27429);
xor UO_484 (O_484,N_29361,N_29088);
nand UO_485 (O_485,N_29248,N_27423);
and UO_486 (O_486,N_27855,N_28496);
xnor UO_487 (O_487,N_27394,N_28477);
or UO_488 (O_488,N_28489,N_29760);
nand UO_489 (O_489,N_27906,N_29834);
nand UO_490 (O_490,N_28630,N_28705);
nand UO_491 (O_491,N_29713,N_29193);
nor UO_492 (O_492,N_28415,N_27269);
xor UO_493 (O_493,N_29289,N_28332);
and UO_494 (O_494,N_27692,N_27169);
or UO_495 (O_495,N_29987,N_29708);
nand UO_496 (O_496,N_28817,N_27103);
xor UO_497 (O_497,N_29094,N_27044);
and UO_498 (O_498,N_28196,N_27607);
and UO_499 (O_499,N_27007,N_28641);
and UO_500 (O_500,N_27063,N_28844);
and UO_501 (O_501,N_29231,N_28542);
nand UO_502 (O_502,N_27760,N_27697);
and UO_503 (O_503,N_27934,N_29393);
xnor UO_504 (O_504,N_27796,N_27778);
or UO_505 (O_505,N_27254,N_28818);
xor UO_506 (O_506,N_28391,N_28681);
nor UO_507 (O_507,N_29217,N_27873);
and UO_508 (O_508,N_29219,N_28825);
and UO_509 (O_509,N_29137,N_27136);
nor UO_510 (O_510,N_27273,N_27552);
or UO_511 (O_511,N_28546,N_27689);
or UO_512 (O_512,N_27400,N_27788);
or UO_513 (O_513,N_29115,N_27120);
and UO_514 (O_514,N_27268,N_29333);
xor UO_515 (O_515,N_28879,N_29785);
nand UO_516 (O_516,N_27838,N_27930);
nand UO_517 (O_517,N_28929,N_29877);
or UO_518 (O_518,N_27237,N_27122);
xnor UO_519 (O_519,N_28731,N_27410);
xnor UO_520 (O_520,N_27996,N_27365);
nor UO_521 (O_521,N_29779,N_27445);
xnor UO_522 (O_522,N_28027,N_28860);
nand UO_523 (O_523,N_29937,N_27490);
nand UO_524 (O_524,N_29202,N_28843);
xnor UO_525 (O_525,N_28522,N_29183);
or UO_526 (O_526,N_28065,N_29146);
nand UO_527 (O_527,N_28900,N_27088);
nand UO_528 (O_528,N_28501,N_27020);
and UO_529 (O_529,N_28461,N_28114);
nand UO_530 (O_530,N_28985,N_28334);
nand UO_531 (O_531,N_27968,N_28329);
or UO_532 (O_532,N_27118,N_29676);
nand UO_533 (O_533,N_28376,N_27603);
nor UO_534 (O_534,N_29996,N_27617);
or UO_535 (O_535,N_27915,N_28142);
and UO_536 (O_536,N_29232,N_28145);
nand UO_537 (O_537,N_29040,N_27556);
nor UO_538 (O_538,N_27595,N_29968);
or UO_539 (O_539,N_27296,N_28480);
xnor UO_540 (O_540,N_27010,N_28018);
and UO_541 (O_541,N_29466,N_28157);
nand UO_542 (O_542,N_28178,N_28398);
nand UO_543 (O_543,N_27797,N_27825);
nor UO_544 (O_544,N_29895,N_28706);
nand UO_545 (O_545,N_28944,N_27004);
nor UO_546 (O_546,N_29419,N_27440);
xor UO_547 (O_547,N_27652,N_29792);
or UO_548 (O_548,N_28109,N_27393);
or UO_549 (O_549,N_28406,N_27249);
nor UO_550 (O_550,N_28782,N_29319);
and UO_551 (O_551,N_29464,N_28777);
nor UO_552 (O_552,N_27961,N_28495);
nand UO_553 (O_553,N_29134,N_28155);
or UO_554 (O_554,N_27081,N_28882);
xor UO_555 (O_555,N_27984,N_28487);
and UO_556 (O_556,N_29475,N_27835);
and UO_557 (O_557,N_27422,N_29903);
or UO_558 (O_558,N_29224,N_28387);
nand UO_559 (O_559,N_28380,N_29840);
or UO_560 (O_560,N_27775,N_29418);
xor UO_561 (O_561,N_28878,N_28919);
nand UO_562 (O_562,N_28475,N_28454);
or UO_563 (O_563,N_28869,N_27579);
or UO_564 (O_564,N_27337,N_27363);
or UO_565 (O_565,N_27080,N_27258);
nand UO_566 (O_566,N_29752,N_27878);
xor UO_567 (O_567,N_27533,N_27133);
and UO_568 (O_568,N_28939,N_27869);
xor UO_569 (O_569,N_29329,N_29273);
nor UO_570 (O_570,N_29620,N_29468);
xnor UO_571 (O_571,N_27801,N_29406);
nand UO_572 (O_572,N_27472,N_28209);
nand UO_573 (O_573,N_28300,N_29473);
or UO_574 (O_574,N_29642,N_28176);
nor UO_575 (O_575,N_28723,N_28794);
nand UO_576 (O_576,N_28892,N_28188);
or UO_577 (O_577,N_29050,N_28439);
or UO_578 (O_578,N_29085,N_29010);
xnor UO_579 (O_579,N_29806,N_29591);
nand UO_580 (O_580,N_28640,N_28971);
or UO_581 (O_581,N_27721,N_28890);
xnor UO_582 (O_582,N_27535,N_29692);
and UO_583 (O_583,N_29322,N_28751);
nand UO_584 (O_584,N_28700,N_28204);
nand UO_585 (O_585,N_27113,N_27073);
or UO_586 (O_586,N_27834,N_28412);
nor UO_587 (O_587,N_27520,N_29212);
nor UO_588 (O_588,N_27956,N_29570);
xor UO_589 (O_589,N_29487,N_29814);
nor UO_590 (O_590,N_29571,N_29290);
and UO_591 (O_591,N_29147,N_29880);
or UO_592 (O_592,N_28441,N_29004);
and UO_593 (O_593,N_28606,N_29983);
nand UO_594 (O_594,N_29909,N_28667);
xnor UO_595 (O_595,N_28592,N_27804);
nor UO_596 (O_596,N_28935,N_29145);
or UO_597 (O_597,N_27532,N_29864);
nor UO_598 (O_598,N_27767,N_29886);
and UO_599 (O_599,N_29793,N_29997);
or UO_600 (O_600,N_29459,N_28560);
nor UO_601 (O_601,N_28254,N_29221);
nor UO_602 (O_602,N_29697,N_28671);
nand UO_603 (O_603,N_27418,N_28307);
or UO_604 (O_604,N_28319,N_28270);
nand UO_605 (O_605,N_29449,N_29271);
or UO_606 (O_606,N_28000,N_27599);
nand UO_607 (O_607,N_29584,N_28729);
nand UO_608 (O_608,N_29956,N_29019);
and UO_609 (O_609,N_28479,N_27043);
and UO_610 (O_610,N_27973,N_28949);
nor UO_611 (O_611,N_28614,N_29399);
and UO_612 (O_612,N_29989,N_29537);
nand UO_613 (O_613,N_27868,N_27199);
xor UO_614 (O_614,N_29855,N_27438);
nand UO_615 (O_615,N_27795,N_29687);
nand UO_616 (O_616,N_27557,N_27385);
or UO_617 (O_617,N_27021,N_29775);
and UO_618 (O_618,N_28868,N_27294);
xor UO_619 (O_619,N_27582,N_29905);
and UO_620 (O_620,N_28095,N_28909);
and UO_621 (O_621,N_29493,N_29656);
and UO_622 (O_622,N_29307,N_28432);
xor UO_623 (O_623,N_27563,N_27894);
nor UO_624 (O_624,N_27197,N_28716);
nor UO_625 (O_625,N_27698,N_29719);
and UO_626 (O_626,N_29737,N_29982);
nor UO_627 (O_627,N_28780,N_29892);
xnor UO_628 (O_628,N_27408,N_28382);
and UO_629 (O_629,N_29980,N_29150);
nand UO_630 (O_630,N_29263,N_29703);
or UO_631 (O_631,N_27031,N_27499);
xor UO_632 (O_632,N_29446,N_28903);
nor UO_633 (O_633,N_29005,N_29764);
and UO_634 (O_634,N_27297,N_28211);
or UO_635 (O_635,N_28833,N_28810);
or UO_636 (O_636,N_29402,N_29001);
nor UO_637 (O_637,N_29481,N_28126);
or UO_638 (O_638,N_29228,N_27235);
nand UO_639 (O_639,N_28964,N_28767);
and UO_640 (O_640,N_29364,N_29900);
and UO_641 (O_641,N_28718,N_27405);
and UO_642 (O_642,N_27724,N_29434);
nand UO_643 (O_643,N_27174,N_28445);
or UO_644 (O_644,N_27664,N_28072);
nor UO_645 (O_645,N_29385,N_27606);
xor UO_646 (O_646,N_27017,N_27643);
nand UO_647 (O_647,N_29500,N_27124);
or UO_648 (O_648,N_29543,N_28612);
nor UO_649 (O_649,N_28282,N_28940);
nor UO_650 (O_650,N_28665,N_29673);
xor UO_651 (O_651,N_29382,N_27215);
xnor UO_652 (O_652,N_28210,N_29772);
or UO_653 (O_653,N_27735,N_28907);
or UO_654 (O_654,N_28460,N_28693);
nor UO_655 (O_655,N_27045,N_28779);
or UO_656 (O_656,N_29634,N_28896);
and UO_657 (O_657,N_27798,N_28003);
xor UO_658 (O_658,N_29887,N_28875);
or UO_659 (O_659,N_27234,N_28973);
xor UO_660 (O_660,N_29695,N_29699);
and UO_661 (O_661,N_27675,N_28673);
or UO_662 (O_662,N_28151,N_27218);
nor UO_663 (O_663,N_28049,N_27161);
and UO_664 (O_664,N_28989,N_28618);
nor UO_665 (O_665,N_29063,N_27489);
nor UO_666 (O_666,N_27592,N_29749);
and UO_667 (O_667,N_28116,N_27181);
and UO_668 (O_668,N_27035,N_27569);
nand UO_669 (O_669,N_29532,N_27955);
or UO_670 (O_670,N_28469,N_29494);
xnor UO_671 (O_671,N_27781,N_28349);
or UO_672 (O_672,N_28735,N_27048);
and UO_673 (O_673,N_28499,N_29032);
nor UO_674 (O_674,N_27587,N_29800);
nand UO_675 (O_675,N_29429,N_29674);
xor UO_676 (O_676,N_28937,N_27099);
xnor UO_677 (O_677,N_29407,N_28778);
nand UO_678 (O_678,N_27981,N_28938);
and UO_679 (O_679,N_29519,N_29334);
xnor UO_680 (O_680,N_29951,N_28983);
and UO_681 (O_681,N_27496,N_28947);
or UO_682 (O_682,N_28273,N_27111);
nand UO_683 (O_683,N_28545,N_28271);
nand UO_684 (O_684,N_29148,N_27288);
xor UO_685 (O_685,N_28742,N_28353);
xnor UO_686 (O_686,N_27131,N_29267);
nand UO_687 (O_687,N_27480,N_29367);
and UO_688 (O_688,N_28908,N_29039);
nor UO_689 (O_689,N_28781,N_29863);
xnor UO_690 (O_690,N_29672,N_28916);
xor UO_691 (O_691,N_27880,N_28250);
and UO_692 (O_692,N_29784,N_27545);
nand UO_693 (O_693,N_27239,N_28462);
xnor UO_694 (O_694,N_27452,N_27439);
nand UO_695 (O_695,N_28272,N_29526);
and UO_696 (O_696,N_29448,N_28195);
nor UO_697 (O_697,N_28994,N_28035);
and UO_698 (O_698,N_29810,N_29716);
nand UO_699 (O_699,N_28456,N_27208);
and UO_700 (O_700,N_28243,N_27139);
nand UO_701 (O_701,N_29562,N_29087);
nand UO_702 (O_702,N_27403,N_28389);
nand UO_703 (O_703,N_28932,N_28682);
nor UO_704 (O_704,N_29952,N_28849);
or UO_705 (O_705,N_29831,N_27227);
and UO_706 (O_706,N_27430,N_27171);
nand UO_707 (O_707,N_29748,N_29763);
and UO_708 (O_708,N_27890,N_28013);
xnor UO_709 (O_709,N_29946,N_29502);
and UO_710 (O_710,N_28968,N_28974);
or UO_711 (O_711,N_28354,N_27548);
nand UO_712 (O_712,N_28851,N_29546);
or UO_713 (O_713,N_29369,N_28593);
xnor UO_714 (O_714,N_28054,N_28514);
xor UO_715 (O_715,N_27225,N_29265);
nand UO_716 (O_716,N_28814,N_29839);
nor UO_717 (O_717,N_29023,N_27432);
nor UO_718 (O_718,N_27334,N_27802);
nand UO_719 (O_719,N_28333,N_27865);
xnor UO_720 (O_720,N_29129,N_28958);
and UO_721 (O_721,N_29081,N_27327);
or UO_722 (O_722,N_28689,N_27657);
and UO_723 (O_723,N_28899,N_28549);
nand UO_724 (O_724,N_29111,N_27622);
xor UO_725 (O_725,N_28409,N_28342);
or UO_726 (O_726,N_28106,N_28002);
and UO_727 (O_727,N_29136,N_27714);
or UO_728 (O_728,N_29609,N_28169);
nand UO_729 (O_729,N_29999,N_27282);
or UO_730 (O_730,N_27576,N_29165);
nor UO_731 (O_731,N_28182,N_28645);
and UO_732 (O_732,N_29404,N_28258);
nor UO_733 (O_733,N_27800,N_28631);
xor UO_734 (O_734,N_27518,N_29540);
nand UO_735 (O_735,N_27395,N_27264);
or UO_736 (O_736,N_27937,N_28870);
or UO_737 (O_737,N_29178,N_27553);
and UO_738 (O_738,N_29632,N_28685);
or UO_739 (O_739,N_28604,N_27085);
nand UO_740 (O_740,N_28683,N_29514);
nor UO_741 (O_741,N_27255,N_28962);
nand UO_742 (O_742,N_28802,N_29326);
nor UO_743 (O_743,N_29897,N_27931);
nand UO_744 (O_744,N_29495,N_29751);
and UO_745 (O_745,N_29966,N_29504);
or UO_746 (O_746,N_28699,N_28590);
nor UO_747 (O_747,N_29710,N_27220);
nand UO_748 (O_748,N_28112,N_27203);
nand UO_749 (O_749,N_29162,N_27701);
nand UO_750 (O_750,N_29563,N_29965);
and UO_751 (O_751,N_29559,N_29501);
nor UO_752 (O_752,N_28865,N_28951);
or UO_753 (O_753,N_29556,N_27925);
xnor UO_754 (O_754,N_28709,N_29961);
or UO_755 (O_755,N_27364,N_27792);
or UO_756 (O_756,N_29149,N_29015);
and UO_757 (O_757,N_29927,N_27217);
or UO_758 (O_758,N_28371,N_29896);
xor UO_759 (O_759,N_27285,N_28895);
and UO_760 (O_760,N_29774,N_29213);
nor UO_761 (O_761,N_28596,N_28955);
or UO_762 (O_762,N_27634,N_27685);
xor UO_763 (O_763,N_27329,N_29133);
and UO_764 (O_764,N_27150,N_27528);
and UO_765 (O_765,N_27069,N_29314);
nand UO_766 (O_766,N_27342,N_27026);
and UO_767 (O_767,N_28351,N_27078);
or UO_768 (O_768,N_28639,N_28071);
xor UO_769 (O_769,N_28083,N_29139);
nor UO_770 (O_770,N_28736,N_27068);
nand UO_771 (O_771,N_27128,N_28637);
nand UO_772 (O_772,N_28218,N_28724);
or UO_773 (O_773,N_29458,N_29550);
xor UO_774 (O_774,N_29128,N_28442);
nand UO_775 (O_775,N_29593,N_27861);
and UO_776 (O_776,N_27808,N_28847);
and UO_777 (O_777,N_29928,N_28291);
xnor UO_778 (O_778,N_29059,N_28528);
or UO_779 (O_779,N_29881,N_29154);
nor UO_780 (O_780,N_28459,N_29661);
nand UO_781 (O_781,N_28292,N_28403);
and UO_782 (O_782,N_27690,N_27736);
nand UO_783 (O_783,N_27419,N_27016);
and UO_784 (O_784,N_28838,N_28568);
xnor UO_785 (O_785,N_28061,N_29205);
xor UO_786 (O_786,N_27897,N_28082);
or UO_787 (O_787,N_29615,N_29302);
and UO_788 (O_788,N_28796,N_28230);
xor UO_789 (O_789,N_29889,N_27250);
nand UO_790 (O_790,N_29078,N_27207);
and UO_791 (O_791,N_27832,N_29239);
nor UO_792 (O_792,N_27971,N_27857);
xor UO_793 (O_793,N_29006,N_29621);
xnor UO_794 (O_794,N_28997,N_27976);
xor UO_795 (O_795,N_29158,N_27001);
nand UO_796 (O_796,N_27695,N_29587);
nand UO_797 (O_797,N_28219,N_28505);
nand UO_798 (O_798,N_28030,N_29541);
nor UO_799 (O_799,N_27598,N_28274);
xnor UO_800 (O_800,N_29732,N_29155);
and UO_801 (O_801,N_28987,N_29611);
nor UO_802 (O_802,N_29179,N_28565);
nand UO_803 (O_803,N_29344,N_28813);
or UO_804 (O_804,N_27636,N_27461);
xnor UO_805 (O_805,N_28055,N_27093);
nor UO_806 (O_806,N_27149,N_27176);
and UO_807 (O_807,N_27558,N_29924);
nand UO_808 (O_808,N_28650,N_27958);
nand UO_809 (O_809,N_29020,N_28133);
and UO_810 (O_810,N_27109,N_29280);
nor UO_811 (O_811,N_28149,N_27446);
xor UO_812 (O_812,N_27899,N_29086);
nor UO_813 (O_813,N_28336,N_28755);
or UO_814 (O_814,N_28521,N_27988);
xnor UO_815 (O_815,N_28168,N_28784);
nor UO_816 (O_816,N_29625,N_29833);
nor UO_817 (O_817,N_28150,N_27565);
and UO_818 (O_818,N_29230,N_28808);
or UO_819 (O_819,N_27485,N_27561);
or UO_820 (O_820,N_28721,N_29601);
and UO_821 (O_821,N_27612,N_27837);
and UO_822 (O_822,N_29293,N_27588);
or UO_823 (O_823,N_29845,N_29497);
nand UO_824 (O_824,N_29251,N_28372);
or UO_825 (O_825,N_27090,N_28800);
nor UO_826 (O_826,N_27823,N_28999);
or UO_827 (O_827,N_29227,N_29899);
nor UO_828 (O_828,N_27790,N_29837);
nor UO_829 (O_829,N_28719,N_27233);
nand UO_830 (O_830,N_28976,N_27040);
nand UO_831 (O_831,N_27289,N_27488);
or UO_832 (O_832,N_28961,N_28369);
nand UO_833 (O_833,N_28713,N_29916);
nor UO_834 (O_834,N_27455,N_27117);
xor UO_835 (O_835,N_29802,N_29535);
nand UO_836 (O_836,N_27641,N_27746);
or UO_837 (O_837,N_28785,N_29350);
or UO_838 (O_838,N_29065,N_29670);
xnor UO_839 (O_839,N_27370,N_29954);
xnor UO_840 (O_840,N_28129,N_27842);
nand UO_841 (O_841,N_27666,N_28765);
nor UO_842 (O_842,N_28430,N_29018);
xor UO_843 (O_843,N_29026,N_29971);
or UO_844 (O_844,N_27302,N_27413);
or UO_845 (O_845,N_27299,N_27030);
xnor UO_846 (O_846,N_29821,N_27932);
nor UO_847 (O_847,N_28009,N_27649);
or UO_848 (O_848,N_27098,N_28128);
nand UO_849 (O_849,N_29104,N_28897);
and UO_850 (O_850,N_27479,N_29034);
nand UO_851 (O_851,N_29681,N_27070);
xor UO_852 (O_852,N_27542,N_27912);
xor UO_853 (O_853,N_29520,N_29803);
and UO_854 (O_854,N_28437,N_28248);
and UO_855 (O_855,N_28124,N_29079);
nor UO_856 (O_856,N_28526,N_27554);
and UO_857 (O_857,N_29893,N_28733);
and UO_858 (O_858,N_28594,N_29884);
xor UO_859 (O_859,N_27986,N_27357);
or UO_860 (O_860,N_29401,N_29849);
nand UO_861 (O_861,N_29123,N_27782);
or UO_862 (O_862,N_27162,N_29776);
and UO_863 (O_863,N_28006,N_27346);
nand UO_864 (O_864,N_28298,N_29627);
and UO_865 (O_865,N_29561,N_27212);
nor UO_866 (O_866,N_29922,N_28296);
and UO_867 (O_867,N_29465,N_29598);
xor UO_868 (O_868,N_27570,N_28714);
nand UO_869 (O_869,N_28694,N_27635);
or UO_870 (O_870,N_29545,N_28761);
nor UO_871 (O_871,N_27252,N_28245);
and UO_872 (O_872,N_28760,N_29107);
or UO_873 (O_873,N_27853,N_28745);
nand UO_874 (O_874,N_28010,N_28338);
nand UO_875 (O_875,N_28080,N_28619);
or UO_876 (O_876,N_27057,N_29091);
and UO_877 (O_877,N_29597,N_29712);
xnor UO_878 (O_878,N_27242,N_29762);
or UO_879 (O_879,N_27067,N_29375);
nor UO_880 (O_880,N_28816,N_28240);
and UO_881 (O_881,N_27637,N_28419);
nand UO_882 (O_882,N_28017,N_27366);
xor UO_883 (O_883,N_29318,N_27079);
and UO_884 (O_884,N_27511,N_29062);
xor UO_885 (O_885,N_28097,N_27793);
nand UO_886 (O_886,N_27141,N_29769);
xor UO_887 (O_887,N_28772,N_27847);
or UO_888 (O_888,N_29159,N_27568);
or UO_889 (O_889,N_27486,N_29410);
xor UO_890 (O_890,N_29549,N_28227);
nor UO_891 (O_891,N_28485,N_28536);
nand UO_892 (O_892,N_27305,N_27015);
nand UO_893 (O_893,N_29663,N_29780);
and UO_894 (O_894,N_27039,N_27148);
xnor UO_895 (O_895,N_27841,N_29272);
or UO_896 (O_896,N_27935,N_29294);
nand UO_897 (O_897,N_27047,N_28891);
nor UO_898 (O_898,N_27467,N_29778);
nand UO_899 (O_899,N_29923,N_29807);
and UO_900 (O_900,N_29812,N_28803);
and UO_901 (O_901,N_28674,N_27822);
xor UO_902 (O_902,N_29492,N_28050);
or UO_903 (O_903,N_29168,N_28677);
xnor UO_904 (O_904,N_28986,N_28636);
nor UO_905 (O_905,N_29258,N_27247);
nor UO_906 (O_906,N_27152,N_27744);
and UO_907 (O_907,N_27962,N_27631);
nand UO_908 (O_908,N_28831,N_27730);
nor UO_909 (O_909,N_28444,N_27351);
nand UO_910 (O_910,N_28040,N_28023);
or UO_911 (O_911,N_27638,N_29635);
nand UO_912 (O_912,N_27226,N_29745);
nor UO_913 (O_913,N_27195,N_29254);
or UO_914 (O_914,N_27892,N_29117);
and UO_915 (O_915,N_27378,N_29339);
xnor UO_916 (O_916,N_28969,N_28287);
and UO_917 (O_917,N_29586,N_27153);
and UO_918 (O_918,N_27628,N_28750);
and UO_919 (O_919,N_28466,N_29683);
or UO_920 (O_920,N_29957,N_28852);
nor UO_921 (O_921,N_29377,N_27326);
and UO_922 (O_922,N_28159,N_28893);
nand UO_923 (O_923,N_29069,N_28203);
xnor UO_924 (O_924,N_29452,N_27198);
or UO_925 (O_925,N_29503,N_27373);
nor UO_926 (O_926,N_29412,N_27495);
nand UO_927 (O_927,N_27428,N_28762);
nand UO_928 (O_928,N_29513,N_27014);
nand UO_929 (O_929,N_28234,N_27427);
and UO_930 (O_930,N_28199,N_28662);
nor UO_931 (O_931,N_28212,N_29171);
or UO_932 (O_932,N_27454,N_28659);
nand UO_933 (O_933,N_28408,N_29191);
nor UO_934 (O_934,N_28165,N_27094);
nand UO_935 (O_935,N_27830,N_28783);
nor UO_936 (O_936,N_28004,N_29631);
nand UO_937 (O_937,N_28192,N_29723);
xor UO_938 (O_938,N_27747,N_28768);
nand UO_939 (O_939,N_28379,N_27874);
or UO_940 (O_940,N_28433,N_29861);
or UO_941 (O_941,N_27944,N_28737);
nand UO_942 (O_942,N_28364,N_27654);
xnor UO_943 (O_943,N_28440,N_27716);
or UO_944 (O_944,N_29327,N_27350);
and UO_945 (O_945,N_29647,N_29757);
xnor UO_946 (O_946,N_27318,N_29560);
and UO_947 (O_947,N_29707,N_27749);
nand UO_948 (O_948,N_28553,N_28236);
nor UO_949 (O_949,N_29786,N_29341);
and UO_950 (O_950,N_27304,N_29991);
nand UO_951 (O_951,N_28980,N_28902);
nand UO_952 (O_952,N_28235,N_28068);
nor UO_953 (O_953,N_27963,N_28221);
nand UO_954 (O_954,N_28491,N_27311);
and UO_955 (O_955,N_27441,N_27251);
xor UO_956 (O_956,N_27500,N_28488);
nor UO_957 (O_957,N_29843,N_28801);
or UO_958 (O_958,N_29098,N_28362);
nand UO_959 (O_959,N_27076,N_27879);
or UO_960 (O_960,N_29216,N_28154);
or UO_961 (O_961,N_27523,N_27889);
or UO_962 (O_962,N_29390,N_28840);
nand UO_963 (O_963,N_29852,N_27995);
nand UO_964 (O_964,N_29106,N_27024);
and UO_965 (O_965,N_27926,N_29386);
and UO_966 (O_966,N_29926,N_27089);
and UO_967 (O_967,N_28752,N_28467);
nand UO_968 (O_968,N_28815,N_28486);
xor UO_969 (O_969,N_28322,N_29097);
nand UO_970 (O_970,N_29172,N_29700);
or UO_971 (O_971,N_29883,N_28829);
or UO_972 (O_972,N_29491,N_29976);
nor UO_973 (O_973,N_29220,N_29653);
xnor UO_974 (O_974,N_29346,N_28077);
or UO_975 (O_975,N_29768,N_28043);
nor UO_976 (O_976,N_27189,N_29262);
or UO_977 (O_977,N_27310,N_29058);
nand UO_978 (O_978,N_29844,N_29684);
nor UO_979 (O_979,N_27922,N_29126);
or UO_980 (O_980,N_27115,N_27236);
and UO_981 (O_981,N_29694,N_29427);
and UO_982 (O_982,N_28134,N_28264);
or UO_983 (O_983,N_27474,N_29630);
nand UO_984 (O_984,N_29138,N_28021);
nand UO_985 (O_985,N_29173,N_29008);
or UO_986 (O_986,N_28303,N_27042);
xnor UO_987 (O_987,N_29722,N_27444);
or UO_988 (O_988,N_29378,N_27306);
xor UO_989 (O_989,N_28509,N_27202);
and UO_990 (O_990,N_29252,N_29348);
nor UO_991 (O_991,N_29682,N_27924);
nor UO_992 (O_992,N_27200,N_29045);
xnor UO_993 (O_993,N_27503,N_29451);
or UO_994 (O_994,N_27465,N_29337);
or UO_995 (O_995,N_29623,N_27443);
and UO_996 (O_996,N_29368,N_28557);
xnor UO_997 (O_997,N_27810,N_27257);
or UO_998 (O_998,N_29841,N_29317);
and UO_999 (O_999,N_28769,N_29135);
xor UO_1000 (O_1000,N_27262,N_28111);
xor UO_1001 (O_1001,N_28056,N_28390);
nor UO_1002 (O_1002,N_29618,N_29959);
or UO_1003 (O_1003,N_29638,N_29960);
nor UO_1004 (O_1004,N_29190,N_27630);
nand UO_1005 (O_1005,N_27525,N_29799);
xor UO_1006 (O_1006,N_29605,N_27686);
xnor UO_1007 (O_1007,N_27522,N_27950);
and UO_1008 (O_1008,N_28572,N_27593);
nor UO_1009 (O_1009,N_29538,N_28957);
or UO_1010 (O_1010,N_28401,N_28136);
nor UO_1011 (O_1011,N_28146,N_28744);
nor UO_1012 (O_1012,N_29669,N_29257);
nor UO_1013 (O_1013,N_27309,N_27143);
nand UO_1014 (O_1014,N_28312,N_28610);
nand UO_1015 (O_1015,N_29858,N_27539);
nor UO_1016 (O_1016,N_27320,N_27301);
nor UO_1017 (O_1017,N_27424,N_27513);
xnor UO_1018 (O_1018,N_29932,N_27620);
nand UO_1019 (O_1019,N_27705,N_27629);
nand UO_1020 (O_1020,N_29939,N_28086);
xnor UO_1021 (O_1021,N_27066,N_29374);
or UO_1022 (O_1022,N_28670,N_28147);
xor UO_1023 (O_1023,N_29771,N_29945);
nor UO_1024 (O_1024,N_28758,N_29141);
or UO_1025 (O_1025,N_29644,N_28220);
or UO_1026 (O_1026,N_28484,N_27086);
nor UO_1027 (O_1027,N_29287,N_28532);
nand UO_1028 (O_1028,N_29184,N_27101);
nor UO_1029 (O_1029,N_28253,N_27891);
or UO_1030 (O_1030,N_27881,N_29380);
nand UO_1031 (O_1031,N_28317,N_27362);
xor UO_1032 (O_1032,N_28239,N_29414);
nor UO_1033 (O_1033,N_27704,N_27253);
xor UO_1034 (O_1034,N_29600,N_29554);
nor UO_1035 (O_1035,N_28793,N_29222);
nor UO_1036 (O_1036,N_29118,N_29599);
nor UO_1037 (O_1037,N_28141,N_28340);
or UO_1038 (O_1038,N_29301,N_28478);
and UO_1039 (O_1039,N_29075,N_27514);
or UO_1040 (O_1040,N_29522,N_27585);
or UO_1041 (O_1041,N_28335,N_29709);
or UO_1042 (O_1042,N_28703,N_28276);
xor UO_1043 (O_1043,N_27693,N_28827);
nor UO_1044 (O_1044,N_27699,N_28757);
or UO_1045 (O_1045,N_27751,N_28404);
and UO_1046 (O_1046,N_29955,N_28967);
nand UO_1047 (O_1047,N_27770,N_28493);
or UO_1048 (O_1048,N_29741,N_28577);
or UO_1049 (O_1049,N_28463,N_29675);
and UO_1050 (O_1050,N_29528,N_27138);
nor UO_1051 (O_1051,N_27765,N_27717);
xor UO_1052 (O_1052,N_29575,N_27388);
nand UO_1053 (O_1053,N_28697,N_29761);
or UO_1054 (O_1054,N_27805,N_27280);
xnor UO_1055 (O_1055,N_28087,N_27888);
xor UO_1056 (O_1056,N_28739,N_28857);
and UO_1057 (O_1057,N_29868,N_27752);
or UO_1058 (O_1058,N_29950,N_29204);
xor UO_1059 (O_1059,N_28707,N_29167);
xor UO_1060 (O_1060,N_28848,N_27084);
or UO_1061 (O_1061,N_28279,N_27313);
xor UO_1062 (O_1062,N_27970,N_27756);
and UO_1063 (O_1063,N_29795,N_29121);
or UO_1064 (O_1064,N_28548,N_27417);
and UO_1065 (O_1065,N_27126,N_28269);
xnor UO_1066 (O_1066,N_27870,N_28024);
nand UO_1067 (O_1067,N_29299,N_27328);
and UO_1068 (O_1068,N_29011,N_27493);
and UO_1069 (O_1069,N_27457,N_29891);
or UO_1070 (O_1070,N_28031,N_27185);
nor UO_1071 (O_1071,N_29809,N_27551);
nor UO_1072 (O_1072,N_29246,N_28608);
xnor UO_1073 (O_1073,N_28537,N_28293);
nor UO_1074 (O_1074,N_27727,N_27184);
and UO_1075 (O_1075,N_29490,N_28375);
nor UO_1076 (O_1076,N_27483,N_28101);
nor UO_1077 (O_1077,N_28044,N_28503);
nand UO_1078 (O_1078,N_29030,N_27720);
and UO_1079 (O_1079,N_27850,N_27896);
or UO_1080 (O_1080,N_28672,N_28554);
and UO_1081 (O_1081,N_27979,N_27611);
nor UO_1082 (O_1082,N_28198,N_27908);
nor UO_1083 (O_1083,N_28585,N_29714);
and UO_1084 (O_1084,N_29397,N_28053);
nor UO_1085 (O_1085,N_27927,N_29036);
xnor UO_1086 (O_1086,N_29766,N_27964);
xnor UO_1087 (O_1087,N_29268,N_28981);
and UO_1088 (O_1088,N_27300,N_28470);
and UO_1089 (O_1089,N_29874,N_27011);
nand UO_1090 (O_1090,N_27843,N_28666);
nor UO_1091 (O_1091,N_28598,N_29144);
xor UO_1092 (O_1092,N_28202,N_29691);
nand UO_1093 (O_1093,N_28451,N_28428);
or UO_1094 (O_1094,N_29921,N_28190);
xnor UO_1095 (O_1095,N_27768,N_27918);
nor UO_1096 (O_1096,N_28011,N_29304);
xor UO_1097 (O_1097,N_28798,N_28587);
nand UO_1098 (O_1098,N_27398,N_28025);
nor UO_1099 (O_1099,N_27132,N_27146);
or UO_1100 (O_1100,N_27876,N_29678);
nand UO_1101 (O_1101,N_27464,N_29424);
nand UO_1102 (O_1102,N_29084,N_28708);
nor UO_1103 (O_1103,N_27270,N_28189);
or UO_1104 (O_1104,N_27192,N_29967);
or UO_1105 (O_1105,N_28653,N_27758);
xnor UO_1106 (O_1106,N_27648,N_29580);
xnor UO_1107 (O_1107,N_29286,N_28213);
nor UO_1108 (O_1108,N_28725,N_29237);
nor UO_1109 (O_1109,N_27578,N_29310);
or UO_1110 (O_1110,N_28575,N_29071);
or UO_1111 (O_1111,N_27256,N_27002);
or UO_1112 (O_1112,N_27572,N_29506);
and UO_1113 (O_1113,N_28850,N_29014);
nor UO_1114 (O_1114,N_27168,N_29862);
or UO_1115 (O_1115,N_28979,N_28835);
or UO_1116 (O_1116,N_29878,N_28120);
or UO_1117 (O_1117,N_28552,N_27816);
or UO_1118 (O_1118,N_29366,N_28656);
and UO_1119 (O_1119,N_27036,N_27214);
and UO_1120 (O_1120,N_29496,N_27095);
xor UO_1121 (O_1121,N_28550,N_27710);
nor UO_1122 (O_1122,N_29354,N_29024);
nor UO_1123 (O_1123,N_29902,N_29122);
and UO_1124 (O_1124,N_27032,N_29643);
nand UO_1125 (O_1125,N_27776,N_29578);
and UO_1126 (O_1126,N_29042,N_28288);
xor UO_1127 (O_1127,N_27665,N_28246);
nand UO_1128 (O_1128,N_29853,N_29331);
nand UO_1129 (O_1129,N_29324,N_27271);
or UO_1130 (O_1130,N_29860,N_27105);
or UO_1131 (O_1131,N_28262,N_29025);
or UO_1132 (O_1132,N_28284,N_29820);
nor UO_1133 (O_1133,N_27574,N_27702);
or UO_1134 (O_1134,N_29066,N_28383);
nor UO_1135 (O_1135,N_28062,N_28431);
or UO_1136 (O_1136,N_27071,N_28450);
nand UO_1137 (O_1137,N_27316,N_27029);
xnor UO_1138 (O_1138,N_28137,N_28438);
nand UO_1139 (O_1139,N_29872,N_29288);
nand UO_1140 (O_1140,N_29335,N_28519);
and UO_1141 (O_1141,N_27550,N_28005);
xnor UO_1142 (O_1142,N_29370,N_28020);
or UO_1143 (O_1143,N_27779,N_29544);
nand UO_1144 (O_1144,N_27992,N_27583);
and UO_1145 (O_1145,N_29639,N_29355);
or UO_1146 (O_1146,N_27983,N_29866);
xor UO_1147 (O_1147,N_28492,N_28309);
or UO_1148 (O_1148,N_27349,N_29984);
and UO_1149 (O_1149,N_28898,N_27687);
nor UO_1150 (O_1150,N_28701,N_28251);
or UO_1151 (O_1151,N_28603,N_29080);
nor UO_1152 (O_1152,N_28323,N_29208);
nand UO_1153 (O_1153,N_27324,N_27534);
and UO_1154 (O_1154,N_28885,N_28854);
nand UO_1155 (O_1155,N_27209,N_29525);
and UO_1156 (O_1156,N_29789,N_28663);
xnor UO_1157 (O_1157,N_28396,N_28664);
or UO_1158 (O_1158,N_27116,N_28563);
xnor UO_1159 (O_1159,N_28407,N_29092);
xor UO_1160 (O_1160,N_29822,N_27938);
nor UO_1161 (O_1161,N_29408,N_28634);
nand UO_1162 (O_1162,N_28943,N_27387);
xnor UO_1163 (O_1163,N_29717,N_27905);
nor UO_1164 (O_1164,N_29908,N_28130);
and UO_1165 (O_1165,N_27210,N_28790);
and UO_1166 (O_1166,N_27470,N_29854);
xnor UO_1167 (O_1167,N_27292,N_28558);
xnor UO_1168 (O_1168,N_28607,N_29116);
xor UO_1169 (O_1169,N_29445,N_28515);
nand UO_1170 (O_1170,N_27338,N_28655);
xnor UO_1171 (O_1171,N_29405,N_29269);
xnor UO_1172 (O_1172,N_28581,N_27447);
or UO_1173 (O_1173,N_27683,N_29373);
xor UO_1174 (O_1174,N_27763,N_28510);
and UO_1175 (O_1175,N_27379,N_27468);
nor UO_1176 (O_1176,N_29003,N_29398);
and UO_1177 (O_1177,N_27684,N_27145);
nor UO_1178 (O_1178,N_27845,N_29740);
or UO_1179 (O_1179,N_28366,N_29867);
xnor UO_1180 (O_1180,N_28278,N_29624);
and UO_1181 (O_1181,N_29070,N_29636);
nand UO_1182 (O_1182,N_27943,N_29617);
nor UO_1183 (O_1183,N_27059,N_27913);
nand UO_1184 (O_1184,N_29234,N_29590);
xnor UO_1185 (O_1185,N_27159,N_27647);
xnor UO_1186 (O_1186,N_29918,N_29622);
nand UO_1187 (O_1187,N_27190,N_29747);
xnor UO_1188 (O_1188,N_28252,N_29457);
xor UO_1189 (O_1189,N_28654,N_29499);
nand UO_1190 (O_1190,N_29530,N_28651);
and UO_1191 (O_1191,N_27784,N_28578);
nand UO_1192 (O_1192,N_28206,N_29282);
nor UO_1193 (O_1193,N_27670,N_29431);
nor UO_1194 (O_1194,N_29211,N_27180);
or UO_1195 (O_1195,N_27246,N_28904);
and UO_1196 (O_1196,N_27248,N_28152);
and UO_1197 (O_1197,N_29478,N_28308);
nand UO_1198 (O_1198,N_27420,N_27994);
and UO_1199 (O_1199,N_27939,N_27399);
nor UO_1200 (O_1200,N_29765,N_27186);
nand UO_1201 (O_1201,N_27773,N_29012);
and UO_1202 (O_1202,N_28763,N_29095);
and UO_1203 (O_1203,N_29728,N_28720);
and UO_1204 (O_1204,N_28059,N_27463);
nor UO_1205 (O_1205,N_27228,N_28635);
xor UO_1206 (O_1206,N_28348,N_29396);
and UO_1207 (O_1207,N_28567,N_28223);
or UO_1208 (O_1208,N_28140,N_27134);
and UO_1209 (O_1209,N_27672,N_27658);
nor UO_1210 (O_1210,N_29975,N_29671);
nor UO_1211 (O_1211,N_29328,N_28052);
nor UO_1212 (O_1212,N_28118,N_29616);
nor UO_1213 (O_1213,N_27851,N_28584);
nor UO_1214 (O_1214,N_29007,N_29788);
and UO_1215 (O_1215,N_28764,N_28320);
nand UO_1216 (O_1216,N_29523,N_27541);
and UO_1217 (O_1217,N_28628,N_28711);
nor UO_1218 (O_1218,N_29592,N_28205);
or UO_1219 (O_1219,N_27562,N_29970);
or UO_1220 (O_1220,N_29626,N_27948);
nor UO_1221 (O_1221,N_28066,N_27515);
nand UO_1222 (O_1222,N_28194,N_27536);
and UO_1223 (O_1223,N_29225,N_28208);
or UO_1224 (O_1224,N_29934,N_29518);
nand UO_1225 (O_1225,N_28078,N_28238);
and UO_1226 (O_1226,N_27600,N_28305);
nor UO_1227 (O_1227,N_29574,N_27487);
xnor UO_1228 (O_1228,N_29274,N_28434);
xor UO_1229 (O_1229,N_28365,N_29013);
nor UO_1230 (O_1230,N_29977,N_28360);
and UO_1231 (O_1231,N_27886,N_29754);
nand UO_1232 (O_1232,N_29781,N_29512);
xnor UO_1233 (O_1233,N_27409,N_28286);
and UO_1234 (O_1234,N_27807,N_28224);
xor UO_1235 (O_1235,N_27033,N_28766);
nand UO_1236 (O_1236,N_29247,N_29315);
or UO_1237 (O_1237,N_27466,N_29660);
and UO_1238 (O_1238,N_29101,N_29073);
nand UO_1239 (O_1239,N_28661,N_27041);
or UO_1240 (O_1240,N_28859,N_29447);
xnor UO_1241 (O_1241,N_27707,N_28471);
or UO_1242 (O_1242,N_27265,N_29284);
nand UO_1243 (O_1243,N_28392,N_28084);
and UO_1244 (O_1244,N_28948,N_29266);
and UO_1245 (O_1245,N_28123,N_28839);
nor UO_1246 (O_1246,N_27114,N_27819);
and UO_1247 (O_1247,N_28984,N_28405);
and UO_1248 (O_1248,N_29016,N_28422);
nor UO_1249 (O_1249,N_28759,N_29195);
and UO_1250 (O_1250,N_28527,N_27353);
nor UO_1251 (O_1251,N_29358,N_28281);
nand UO_1252 (O_1252,N_29017,N_29613);
or UO_1253 (O_1253,N_28726,N_29038);
and UO_1254 (O_1254,N_28513,N_27481);
nand UO_1255 (O_1255,N_29383,N_28057);
nor UO_1256 (O_1256,N_27333,N_27531);
nand UO_1257 (O_1257,N_29825,N_27809);
nand UO_1258 (O_1258,N_27129,N_27177);
or UO_1259 (O_1259,N_29480,N_29027);
and UO_1260 (O_1260,N_27663,N_27284);
nand UO_1261 (O_1261,N_27056,N_27729);
or UO_1262 (O_1262,N_29277,N_29667);
and UO_1263 (O_1263,N_29072,N_28089);
xnor UO_1264 (O_1264,N_27046,N_28611);
and UO_1265 (O_1265,N_28931,N_27872);
nand UO_1266 (O_1266,N_27610,N_27718);
or UO_1267 (O_1267,N_28022,N_28229);
nand UO_1268 (O_1268,N_28792,N_27679);
or UO_1269 (O_1269,N_27954,N_27414);
nor UO_1270 (O_1270,N_27537,N_29000);
and UO_1271 (O_1271,N_29306,N_28629);
xor UO_1272 (O_1272,N_27911,N_27166);
nor UO_1273 (O_1273,N_27820,N_28555);
nor UO_1274 (O_1274,N_27815,N_27659);
xnor UO_1275 (O_1275,N_29450,N_29186);
xor UO_1276 (O_1276,N_28108,N_28377);
nor UO_1277 (O_1277,N_29305,N_27947);
nand UO_1278 (O_1278,N_29859,N_27003);
or UO_1279 (O_1279,N_29113,N_27712);
nor UO_1280 (O_1280,N_27708,N_28113);
or UO_1281 (O_1281,N_28836,N_27575);
nand UO_1282 (O_1282,N_27516,N_27437);
nor UO_1283 (O_1283,N_27696,N_27589);
xor UO_1284 (O_1284,N_27799,N_29430);
xor UO_1285 (O_1285,N_27978,N_27355);
xnor UO_1286 (O_1286,N_28561,N_29391);
or UO_1287 (O_1287,N_29531,N_29572);
nand UO_1288 (O_1288,N_27900,N_27653);
nand UO_1289 (O_1289,N_27431,N_29332);
nor UO_1290 (O_1290,N_28497,N_29389);
nor UO_1291 (O_1291,N_27104,N_28280);
nand UO_1292 (O_1292,N_29963,N_27451);
nand UO_1293 (O_1293,N_27241,N_27786);
or UO_1294 (O_1294,N_28476,N_29917);
and UO_1295 (O_1295,N_28846,N_29484);
or UO_1296 (O_1296,N_28465,N_28344);
nand UO_1297 (O_1297,N_28912,N_28331);
and UO_1298 (O_1298,N_27725,N_29180);
xor UO_1299 (O_1299,N_29124,N_27358);
nor UO_1300 (O_1300,N_29654,N_28081);
and UO_1301 (O_1301,N_29935,N_27060);
and UO_1302 (O_1302,N_29904,N_28104);
nor UO_1303 (O_1303,N_28867,N_29029);
and UO_1304 (O_1304,N_28161,N_28184);
and UO_1305 (O_1305,N_27590,N_27272);
and UO_1306 (O_1306,N_28131,N_28481);
and UO_1307 (O_1307,N_27179,N_27022);
and UO_1308 (O_1308,N_27266,N_29628);
or UO_1309 (O_1309,N_28525,N_28529);
or UO_1310 (O_1310,N_27910,N_28047);
and UO_1311 (O_1311,N_27092,N_27517);
or UO_1312 (O_1312,N_27182,N_28627);
nand UO_1313 (O_1313,N_29836,N_27206);
and UO_1314 (O_1314,N_27987,N_29108);
and UO_1315 (O_1315,N_28275,N_27680);
or UO_1316 (O_1316,N_27602,N_29517);
or UO_1317 (O_1317,N_29515,N_29696);
nand UO_1318 (O_1318,N_28268,N_28346);
xor UO_1319 (O_1319,N_27661,N_28993);
xnor UO_1320 (O_1320,N_28038,N_29351);
or UO_1321 (O_1321,N_28959,N_27519);
xor UO_1322 (O_1322,N_27211,N_29189);
and UO_1323 (O_1323,N_29256,N_29052);
nand UO_1324 (O_1324,N_29974,N_27061);
nor UO_1325 (O_1325,N_29629,N_27087);
nand UO_1326 (O_1326,N_27785,N_28201);
or UO_1327 (O_1327,N_28183,N_29856);
and UO_1328 (O_1328,N_27501,N_27783);
and UO_1329 (O_1329,N_29392,N_28473);
nand UO_1330 (O_1330,N_27811,N_29125);
and UO_1331 (O_1331,N_29164,N_28540);
nor UO_1332 (O_1332,N_28457,N_29471);
xor UO_1333 (O_1333,N_28225,N_27639);
nor UO_1334 (O_1334,N_28410,N_28325);
xnor UO_1335 (O_1335,N_28905,N_27340);
nor UO_1336 (O_1336,N_28426,N_28771);
nor UO_1337 (O_1337,N_27119,N_28888);
nand UO_1338 (O_1338,N_28576,N_27856);
nand UO_1339 (O_1339,N_29432,N_28356);
and UO_1340 (O_1340,N_29666,N_27096);
nand UO_1341 (O_1341,N_28886,N_29758);
or UO_1342 (O_1342,N_29413,N_28730);
xor UO_1343 (O_1343,N_29940,N_29777);
and UO_1344 (O_1344,N_29177,N_27157);
and UO_1345 (O_1345,N_28429,N_28185);
nand UO_1346 (O_1346,N_28512,N_28093);
xnor UO_1347 (O_1347,N_28494,N_29308);
nor UO_1348 (O_1348,N_29285,N_29426);
xor UO_1349 (O_1349,N_27188,N_27875);
or UO_1350 (O_1350,N_28901,N_27339);
or UO_1351 (O_1351,N_29461,N_28502);
xnor UO_1352 (O_1352,N_27276,N_28121);
nor UO_1353 (O_1353,N_28384,N_27383);
xor UO_1354 (O_1354,N_28153,N_29394);
nor UO_1355 (O_1355,N_28657,N_28359);
or UO_1356 (O_1356,N_29347,N_28982);
or UO_1357 (O_1357,N_28144,N_27224);
or UO_1358 (O_1358,N_27867,N_27916);
nand UO_1359 (O_1359,N_29022,N_27352);
nand UO_1360 (O_1360,N_27688,N_28679);
or UO_1361 (O_1361,N_28191,N_27219);
nor UO_1362 (O_1362,N_29203,N_29002);
nor UO_1363 (O_1363,N_27274,N_29650);
xnor UO_1364 (O_1364,N_28042,N_29236);
nand UO_1365 (O_1365,N_27615,N_29047);
and UO_1366 (O_1366,N_29425,N_28819);
or UO_1367 (O_1367,N_27425,N_28649);
or UO_1368 (O_1368,N_28871,N_28327);
nand UO_1369 (O_1369,N_28569,N_28828);
nor UO_1370 (O_1370,N_27674,N_27920);
or UO_1371 (O_1371,N_28695,N_29174);
or UO_1372 (O_1372,N_27275,N_28579);
and UO_1373 (O_1373,N_28458,N_28547);
and UO_1374 (O_1374,N_29376,N_27183);
nand UO_1375 (O_1375,N_27748,N_27460);
and UO_1376 (O_1376,N_28260,N_29832);
nand UO_1377 (O_1377,N_27571,N_29569);
xnor UO_1378 (O_1378,N_29901,N_29198);
and UO_1379 (O_1379,N_29529,N_27898);
nor UO_1380 (O_1380,N_28016,N_27677);
nand UO_1381 (O_1381,N_29359,N_28995);
or UO_1382 (O_1382,N_29463,N_27065);
and UO_1383 (O_1383,N_27642,N_27110);
nand UO_1384 (O_1384,N_29658,N_29279);
and UO_1385 (O_1385,N_28727,N_27917);
xor UO_1386 (O_1386,N_29099,N_28534);
or UO_1387 (O_1387,N_29595,N_28306);
and UO_1388 (O_1388,N_28424,N_28691);
and UO_1389 (O_1389,N_28217,N_28615);
nor UO_1390 (O_1390,N_29170,N_27691);
xor UO_1391 (O_1391,N_28012,N_27597);
or UO_1392 (O_1392,N_28326,N_27700);
nor UO_1393 (O_1393,N_28330,N_29074);
nand UO_1394 (O_1394,N_27175,N_27975);
and UO_1395 (O_1395,N_29819,N_29619);
xor UO_1396 (O_1396,N_28490,N_28233);
nand UO_1397 (O_1397,N_28079,N_28811);
nor UO_1398 (O_1398,N_28992,N_28075);
nor UO_1399 (O_1399,N_28449,N_28574);
xnor UO_1400 (O_1400,N_27295,N_27991);
nor UO_1401 (O_1401,N_29400,N_27678);
xnor UO_1402 (O_1402,N_27952,N_28520);
xor UO_1403 (O_1403,N_28530,N_27082);
nand UO_1404 (O_1404,N_27676,N_28255);
xor UO_1405 (O_1405,N_27123,N_29885);
and UO_1406 (O_1406,N_29226,N_29555);
nor UO_1407 (O_1407,N_28978,N_29739);
and UO_1408 (O_1408,N_27343,N_27127);
nor UO_1409 (O_1409,N_29163,N_28448);
or UO_1410 (O_1410,N_29668,N_27928);
xnor UO_1411 (O_1411,N_29275,N_29105);
nand UO_1412 (O_1412,N_27901,N_29482);
nor UO_1413 (O_1413,N_28680,N_28622);
and UO_1414 (O_1414,N_28175,N_27325);
nand UO_1415 (O_1415,N_28822,N_27494);
or UO_1416 (O_1416,N_27389,N_27821);
or UO_1417 (O_1417,N_27106,N_28295);
xor UO_1418 (O_1418,N_28266,N_29421);
nand UO_1419 (O_1419,N_28910,N_29941);
and UO_1420 (O_1420,N_29879,N_27267);
xnor UO_1421 (O_1421,N_28688,N_29734);
xnor UO_1422 (O_1422,N_28029,N_28402);
nor UO_1423 (O_1423,N_29756,N_28924);
xnor UO_1424 (O_1424,N_27456,N_28646);
and UO_1425 (O_1425,N_27397,N_27914);
nand UO_1426 (O_1426,N_28946,N_28941);
or UO_1427 (O_1427,N_27344,N_28110);
and UO_1428 (O_1428,N_28060,N_27544);
and UO_1429 (O_1429,N_27459,N_29250);
or UO_1430 (O_1430,N_29240,N_29388);
or UO_1431 (O_1431,N_27308,N_28877);
and UO_1432 (O_1432,N_29894,N_29077);
nand UO_1433 (O_1433,N_29303,N_27137);
nor UO_1434 (O_1434,N_27433,N_29270);
xnor UO_1435 (O_1435,N_27037,N_29488);
or UO_1436 (O_1436,N_27764,N_29031);
nor UO_1437 (O_1437,N_27194,N_29192);
or UO_1438 (O_1438,N_28589,N_27959);
and UO_1439 (O_1439,N_27165,N_28474);
or UO_1440 (O_1440,N_27009,N_27000);
and UO_1441 (O_1441,N_27726,N_29260);
xor UO_1442 (O_1442,N_28826,N_27871);
nand UO_1443 (O_1443,N_27371,N_27453);
nor UO_1444 (O_1444,N_27396,N_29875);
or UO_1445 (O_1445,N_29794,N_27303);
nand UO_1446 (O_1446,N_27008,N_29281);
or UO_1447 (O_1447,N_29365,N_29498);
or UO_1448 (O_1448,N_27829,N_28231);
or UO_1449 (O_1449,N_27238,N_28139);
nand UO_1450 (O_1450,N_27734,N_28824);
nor UO_1451 (O_1451,N_27671,N_28972);
xnor UO_1452 (O_1452,N_27960,N_29664);
nor UO_1453 (O_1453,N_27164,N_27107);
or UO_1454 (O_1454,N_28823,N_28738);
or UO_1455 (O_1455,N_27766,N_29533);
and UO_1456 (O_1456,N_28259,N_29826);
nor UO_1457 (O_1457,N_29738,N_28620);
nor UO_1458 (O_1458,N_29477,N_28933);
xor UO_1459 (O_1459,N_27213,N_28740);
or UO_1460 (O_1460,N_29357,N_29132);
and UO_1461 (O_1461,N_29633,N_27715);
nor UO_1462 (O_1462,N_27803,N_29614);
xnor UO_1463 (O_1463,N_29420,N_29235);
nand UO_1464 (O_1464,N_29422,N_28743);
xnor UO_1465 (O_1465,N_27322,N_28237);
nor UO_1466 (O_1466,N_28115,N_29548);
and UO_1467 (O_1467,N_28517,N_27624);
nand UO_1468 (O_1468,N_27323,N_29411);
nand UO_1469 (O_1469,N_29558,N_28687);
or UO_1470 (O_1470,N_28156,N_27442);
and UO_1471 (O_1471,N_28668,N_29998);
or UO_1472 (O_1472,N_27998,N_27828);
or UO_1473 (O_1473,N_29089,N_28378);
nand UO_1474 (O_1474,N_27757,N_29835);
nand UO_1475 (O_1475,N_27591,N_29680);
nor UO_1476 (O_1476,N_27223,N_27669);
xnor UO_1477 (O_1477,N_27244,N_28014);
or UO_1478 (O_1478,N_28884,N_29994);
xor UO_1479 (O_1479,N_29455,N_28660);
xor UO_1480 (O_1480,N_28400,N_28337);
xnor UO_1481 (O_1481,N_28538,N_27740);
nor UO_1482 (O_1482,N_27058,N_28119);
or UO_1483 (O_1483,N_28773,N_29930);
nor UO_1484 (O_1484,N_27279,N_27844);
nand UO_1485 (O_1485,N_29049,N_27812);
nand UO_1486 (O_1486,N_28074,N_27573);
and UO_1487 (O_1487,N_27231,N_28261);
xor UO_1488 (O_1488,N_28417,N_29428);
xor UO_1489 (O_1489,N_28001,N_29152);
xnor UO_1490 (O_1490,N_28289,N_28648);
or UO_1491 (O_1491,N_29842,N_28507);
and UO_1492 (O_1492,N_28008,N_28347);
xor UO_1493 (O_1493,N_29442,N_28863);
nor UO_1494 (O_1494,N_27737,N_29194);
nor UO_1495 (O_1495,N_27559,N_29342);
or UO_1496 (O_1496,N_29209,N_27949);
or UO_1497 (O_1497,N_27027,N_28696);
nor UO_1498 (O_1498,N_29542,N_29166);
and UO_1499 (O_1499,N_28539,N_29607);
and UO_1500 (O_1500,N_27057,N_29747);
nand UO_1501 (O_1501,N_27587,N_28583);
or UO_1502 (O_1502,N_27373,N_28007);
xor UO_1503 (O_1503,N_27848,N_28875);
or UO_1504 (O_1504,N_27372,N_27486);
nor UO_1505 (O_1505,N_28437,N_29179);
and UO_1506 (O_1506,N_29941,N_29279);
and UO_1507 (O_1507,N_27116,N_27067);
xnor UO_1508 (O_1508,N_28843,N_28402);
or UO_1509 (O_1509,N_28738,N_29826);
nor UO_1510 (O_1510,N_27616,N_29053);
or UO_1511 (O_1511,N_29455,N_28117);
nor UO_1512 (O_1512,N_27759,N_29093);
or UO_1513 (O_1513,N_28072,N_29438);
and UO_1514 (O_1514,N_29790,N_28507);
nor UO_1515 (O_1515,N_29689,N_29695);
and UO_1516 (O_1516,N_29332,N_28371);
or UO_1517 (O_1517,N_27375,N_27563);
nand UO_1518 (O_1518,N_27388,N_28124);
xor UO_1519 (O_1519,N_29787,N_28045);
xnor UO_1520 (O_1520,N_29409,N_28429);
nand UO_1521 (O_1521,N_28483,N_29189);
or UO_1522 (O_1522,N_27391,N_28457);
nor UO_1523 (O_1523,N_27991,N_29660);
xnor UO_1524 (O_1524,N_27643,N_28923);
xor UO_1525 (O_1525,N_29981,N_29801);
or UO_1526 (O_1526,N_27135,N_29810);
nor UO_1527 (O_1527,N_29889,N_27537);
nand UO_1528 (O_1528,N_27961,N_28594);
or UO_1529 (O_1529,N_29500,N_27319);
or UO_1530 (O_1530,N_29646,N_29999);
and UO_1531 (O_1531,N_29831,N_29638);
xnor UO_1532 (O_1532,N_28799,N_28387);
nor UO_1533 (O_1533,N_29700,N_28413);
nor UO_1534 (O_1534,N_28117,N_28551);
and UO_1535 (O_1535,N_27106,N_27922);
xor UO_1536 (O_1536,N_28973,N_29711);
or UO_1537 (O_1537,N_28807,N_28933);
or UO_1538 (O_1538,N_29975,N_28066);
nor UO_1539 (O_1539,N_28142,N_27255);
nor UO_1540 (O_1540,N_27710,N_27168);
or UO_1541 (O_1541,N_29835,N_28487);
and UO_1542 (O_1542,N_28475,N_28917);
or UO_1543 (O_1543,N_27967,N_29943);
nand UO_1544 (O_1544,N_27581,N_28416);
nand UO_1545 (O_1545,N_28169,N_27557);
nor UO_1546 (O_1546,N_29011,N_28558);
nand UO_1547 (O_1547,N_27382,N_27656);
xnor UO_1548 (O_1548,N_28552,N_27821);
nand UO_1549 (O_1549,N_28713,N_27076);
nand UO_1550 (O_1550,N_28207,N_28254);
nor UO_1551 (O_1551,N_29491,N_28740);
nand UO_1552 (O_1552,N_29651,N_28664);
and UO_1553 (O_1553,N_29485,N_27141);
nor UO_1554 (O_1554,N_28589,N_29880);
and UO_1555 (O_1555,N_27072,N_28237);
and UO_1556 (O_1556,N_29303,N_28698);
nand UO_1557 (O_1557,N_27698,N_29076);
nor UO_1558 (O_1558,N_28424,N_29467);
and UO_1559 (O_1559,N_27189,N_28373);
xnor UO_1560 (O_1560,N_28780,N_27477);
nor UO_1561 (O_1561,N_28102,N_27726);
and UO_1562 (O_1562,N_27946,N_27289);
xnor UO_1563 (O_1563,N_29347,N_27478);
xnor UO_1564 (O_1564,N_27386,N_28823);
xnor UO_1565 (O_1565,N_28117,N_28056);
xnor UO_1566 (O_1566,N_27123,N_28825);
xnor UO_1567 (O_1567,N_28554,N_28182);
nand UO_1568 (O_1568,N_28879,N_27971);
nand UO_1569 (O_1569,N_27360,N_27275);
nor UO_1570 (O_1570,N_27503,N_27555);
or UO_1571 (O_1571,N_29882,N_28572);
nand UO_1572 (O_1572,N_28036,N_28422);
or UO_1573 (O_1573,N_28379,N_29809);
and UO_1574 (O_1574,N_29250,N_29607);
nor UO_1575 (O_1575,N_28720,N_27882);
or UO_1576 (O_1576,N_29209,N_29373);
xor UO_1577 (O_1577,N_29428,N_27177);
or UO_1578 (O_1578,N_28350,N_28272);
or UO_1579 (O_1579,N_27143,N_29903);
or UO_1580 (O_1580,N_27031,N_27358);
or UO_1581 (O_1581,N_28785,N_28721);
nand UO_1582 (O_1582,N_27739,N_29672);
nor UO_1583 (O_1583,N_29837,N_29042);
and UO_1584 (O_1584,N_27054,N_28704);
and UO_1585 (O_1585,N_28787,N_29243);
and UO_1586 (O_1586,N_27459,N_28345);
xor UO_1587 (O_1587,N_29836,N_27449);
nand UO_1588 (O_1588,N_29431,N_27495);
xor UO_1589 (O_1589,N_28741,N_28085);
or UO_1590 (O_1590,N_28343,N_27662);
nand UO_1591 (O_1591,N_27459,N_27747);
or UO_1592 (O_1592,N_28015,N_29151);
or UO_1593 (O_1593,N_27583,N_28812);
or UO_1594 (O_1594,N_27257,N_28506);
nor UO_1595 (O_1595,N_27292,N_29983);
nor UO_1596 (O_1596,N_28135,N_29177);
nor UO_1597 (O_1597,N_29710,N_27323);
or UO_1598 (O_1598,N_29598,N_28438);
nand UO_1599 (O_1599,N_27899,N_27133);
nand UO_1600 (O_1600,N_28844,N_28565);
nand UO_1601 (O_1601,N_29806,N_28407);
and UO_1602 (O_1602,N_28617,N_27588);
and UO_1603 (O_1603,N_28832,N_29921);
and UO_1604 (O_1604,N_27461,N_29696);
or UO_1605 (O_1605,N_27438,N_27667);
nor UO_1606 (O_1606,N_27671,N_28453);
nor UO_1607 (O_1607,N_29804,N_28278);
and UO_1608 (O_1608,N_28418,N_29918);
nand UO_1609 (O_1609,N_27792,N_27935);
nor UO_1610 (O_1610,N_28475,N_28048);
nand UO_1611 (O_1611,N_27769,N_28867);
or UO_1612 (O_1612,N_29360,N_27841);
xor UO_1613 (O_1613,N_28471,N_27430);
nor UO_1614 (O_1614,N_29446,N_27733);
and UO_1615 (O_1615,N_29449,N_27266);
xnor UO_1616 (O_1616,N_29026,N_27530);
xnor UO_1617 (O_1617,N_28893,N_28892);
nor UO_1618 (O_1618,N_28392,N_29636);
and UO_1619 (O_1619,N_28114,N_27024);
xnor UO_1620 (O_1620,N_29118,N_27811);
nor UO_1621 (O_1621,N_29485,N_28813);
or UO_1622 (O_1622,N_27487,N_28960);
xor UO_1623 (O_1623,N_27439,N_29577);
or UO_1624 (O_1624,N_28498,N_29382);
xnor UO_1625 (O_1625,N_27243,N_29992);
xor UO_1626 (O_1626,N_27788,N_29655);
nor UO_1627 (O_1627,N_28049,N_29653);
nor UO_1628 (O_1628,N_28532,N_29769);
nand UO_1629 (O_1629,N_29916,N_29839);
xor UO_1630 (O_1630,N_27679,N_28513);
or UO_1631 (O_1631,N_28010,N_29216);
nor UO_1632 (O_1632,N_27234,N_29338);
nand UO_1633 (O_1633,N_28096,N_29459);
nor UO_1634 (O_1634,N_27106,N_28715);
or UO_1635 (O_1635,N_28549,N_27923);
xnor UO_1636 (O_1636,N_27465,N_27428);
or UO_1637 (O_1637,N_27390,N_28869);
xor UO_1638 (O_1638,N_29134,N_27754);
and UO_1639 (O_1639,N_28444,N_28125);
nor UO_1640 (O_1640,N_29268,N_28537);
and UO_1641 (O_1641,N_29472,N_28292);
and UO_1642 (O_1642,N_28979,N_28887);
nor UO_1643 (O_1643,N_27978,N_28105);
xnor UO_1644 (O_1644,N_28416,N_28907);
and UO_1645 (O_1645,N_27692,N_28661);
xor UO_1646 (O_1646,N_29096,N_28796);
nor UO_1647 (O_1647,N_28681,N_27642);
nand UO_1648 (O_1648,N_28100,N_28830);
xnor UO_1649 (O_1649,N_27946,N_28329);
nand UO_1650 (O_1650,N_29215,N_28961);
and UO_1651 (O_1651,N_27766,N_28505);
xnor UO_1652 (O_1652,N_29711,N_27449);
xor UO_1653 (O_1653,N_29645,N_27295);
or UO_1654 (O_1654,N_29958,N_29998);
nand UO_1655 (O_1655,N_29718,N_28248);
xor UO_1656 (O_1656,N_29763,N_27370);
nor UO_1657 (O_1657,N_29554,N_27792);
and UO_1658 (O_1658,N_27597,N_28825);
or UO_1659 (O_1659,N_29069,N_29142);
and UO_1660 (O_1660,N_29670,N_27059);
xnor UO_1661 (O_1661,N_29243,N_28669);
and UO_1662 (O_1662,N_28476,N_27881);
and UO_1663 (O_1663,N_29578,N_27625);
or UO_1664 (O_1664,N_28873,N_27344);
nor UO_1665 (O_1665,N_27933,N_28201);
nand UO_1666 (O_1666,N_27811,N_29822);
nand UO_1667 (O_1667,N_27144,N_28323);
xor UO_1668 (O_1668,N_28120,N_27029);
nor UO_1669 (O_1669,N_27721,N_29657);
xnor UO_1670 (O_1670,N_29828,N_28258);
xnor UO_1671 (O_1671,N_27404,N_28335);
xor UO_1672 (O_1672,N_29206,N_28037);
nand UO_1673 (O_1673,N_29401,N_28482);
xnor UO_1674 (O_1674,N_29723,N_27794);
xnor UO_1675 (O_1675,N_28275,N_29545);
nand UO_1676 (O_1676,N_27745,N_28526);
or UO_1677 (O_1677,N_29120,N_28806);
nor UO_1678 (O_1678,N_27967,N_29455);
or UO_1679 (O_1679,N_29473,N_27736);
or UO_1680 (O_1680,N_27348,N_28714);
xnor UO_1681 (O_1681,N_29256,N_29197);
and UO_1682 (O_1682,N_27589,N_29728);
and UO_1683 (O_1683,N_27113,N_28062);
nor UO_1684 (O_1684,N_29890,N_29102);
and UO_1685 (O_1685,N_29933,N_29114);
nor UO_1686 (O_1686,N_27793,N_27835);
or UO_1687 (O_1687,N_29041,N_28706);
xnor UO_1688 (O_1688,N_27055,N_27070);
and UO_1689 (O_1689,N_27158,N_28563);
and UO_1690 (O_1690,N_27549,N_29880);
nand UO_1691 (O_1691,N_28175,N_29179);
nand UO_1692 (O_1692,N_27660,N_28641);
and UO_1693 (O_1693,N_29198,N_29409);
xnor UO_1694 (O_1694,N_28645,N_27940);
nand UO_1695 (O_1695,N_28716,N_29688);
nor UO_1696 (O_1696,N_29905,N_28478);
and UO_1697 (O_1697,N_28484,N_29011);
xnor UO_1698 (O_1698,N_27440,N_28363);
and UO_1699 (O_1699,N_29120,N_28219);
or UO_1700 (O_1700,N_29069,N_27800);
nand UO_1701 (O_1701,N_28130,N_28280);
nand UO_1702 (O_1702,N_27700,N_27111);
and UO_1703 (O_1703,N_27620,N_29244);
xnor UO_1704 (O_1704,N_29111,N_28877);
nor UO_1705 (O_1705,N_29738,N_27537);
nor UO_1706 (O_1706,N_28065,N_29973);
nor UO_1707 (O_1707,N_27983,N_28787);
xnor UO_1708 (O_1708,N_29947,N_28816);
and UO_1709 (O_1709,N_29225,N_27020);
and UO_1710 (O_1710,N_28419,N_28305);
and UO_1711 (O_1711,N_29391,N_27830);
nor UO_1712 (O_1712,N_29331,N_27240);
nor UO_1713 (O_1713,N_27313,N_29746);
nand UO_1714 (O_1714,N_27677,N_28615);
or UO_1715 (O_1715,N_27944,N_29618);
nor UO_1716 (O_1716,N_28578,N_28892);
nor UO_1717 (O_1717,N_27036,N_29486);
or UO_1718 (O_1718,N_28161,N_29567);
and UO_1719 (O_1719,N_28959,N_28169);
nor UO_1720 (O_1720,N_29486,N_27490);
or UO_1721 (O_1721,N_29677,N_29675);
nand UO_1722 (O_1722,N_28197,N_27724);
and UO_1723 (O_1723,N_28256,N_27017);
and UO_1724 (O_1724,N_28842,N_27203);
and UO_1725 (O_1725,N_27012,N_29135);
and UO_1726 (O_1726,N_29128,N_28032);
nand UO_1727 (O_1727,N_27464,N_29947);
nor UO_1728 (O_1728,N_28688,N_28372);
nand UO_1729 (O_1729,N_29803,N_27386);
nand UO_1730 (O_1730,N_28417,N_29951);
xnor UO_1731 (O_1731,N_27278,N_27848);
nor UO_1732 (O_1732,N_27253,N_27196);
nand UO_1733 (O_1733,N_29838,N_29054);
nor UO_1734 (O_1734,N_29971,N_28958);
xor UO_1735 (O_1735,N_28115,N_27559);
or UO_1736 (O_1736,N_29456,N_27715);
nor UO_1737 (O_1737,N_29899,N_28247);
nor UO_1738 (O_1738,N_27803,N_28627);
and UO_1739 (O_1739,N_28729,N_29904);
xnor UO_1740 (O_1740,N_27105,N_27345);
or UO_1741 (O_1741,N_28446,N_27753);
nand UO_1742 (O_1742,N_29359,N_29912);
and UO_1743 (O_1743,N_27592,N_27851);
and UO_1744 (O_1744,N_28023,N_27792);
xnor UO_1745 (O_1745,N_27219,N_28222);
and UO_1746 (O_1746,N_27796,N_28760);
and UO_1747 (O_1747,N_29628,N_28791);
and UO_1748 (O_1748,N_28137,N_29287);
nand UO_1749 (O_1749,N_28435,N_28644);
nor UO_1750 (O_1750,N_29900,N_29390);
and UO_1751 (O_1751,N_29084,N_29199);
and UO_1752 (O_1752,N_27495,N_29646);
and UO_1753 (O_1753,N_29832,N_28670);
nand UO_1754 (O_1754,N_28698,N_29057);
nor UO_1755 (O_1755,N_29140,N_28947);
nor UO_1756 (O_1756,N_27547,N_29936);
nand UO_1757 (O_1757,N_27595,N_29857);
and UO_1758 (O_1758,N_27810,N_29096);
and UO_1759 (O_1759,N_29140,N_29688);
and UO_1760 (O_1760,N_29682,N_27954);
nor UO_1761 (O_1761,N_29766,N_29153);
xor UO_1762 (O_1762,N_28646,N_27639);
nor UO_1763 (O_1763,N_28899,N_29402);
nand UO_1764 (O_1764,N_29339,N_27372);
or UO_1765 (O_1765,N_29258,N_28082);
xor UO_1766 (O_1766,N_27034,N_28955);
or UO_1767 (O_1767,N_27352,N_29897);
nor UO_1768 (O_1768,N_28653,N_27310);
or UO_1769 (O_1769,N_28250,N_29959);
and UO_1770 (O_1770,N_28174,N_28796);
nor UO_1771 (O_1771,N_28714,N_29563);
nor UO_1772 (O_1772,N_29868,N_27019);
nor UO_1773 (O_1773,N_28878,N_27007);
xnor UO_1774 (O_1774,N_29886,N_29035);
xnor UO_1775 (O_1775,N_27213,N_27146);
and UO_1776 (O_1776,N_27483,N_28499);
or UO_1777 (O_1777,N_27244,N_28515);
nand UO_1778 (O_1778,N_27922,N_28531);
nand UO_1779 (O_1779,N_28666,N_27990);
xor UO_1780 (O_1780,N_27841,N_29584);
or UO_1781 (O_1781,N_28044,N_28188);
xor UO_1782 (O_1782,N_29134,N_29006);
xnor UO_1783 (O_1783,N_27937,N_28791);
nand UO_1784 (O_1784,N_29643,N_29273);
or UO_1785 (O_1785,N_27406,N_28127);
nor UO_1786 (O_1786,N_29956,N_28871);
and UO_1787 (O_1787,N_29353,N_28407);
xnor UO_1788 (O_1788,N_29583,N_27683);
nor UO_1789 (O_1789,N_27136,N_27084);
xor UO_1790 (O_1790,N_28819,N_27259);
xnor UO_1791 (O_1791,N_28553,N_28722);
xor UO_1792 (O_1792,N_28166,N_28293);
or UO_1793 (O_1793,N_27692,N_28428);
nand UO_1794 (O_1794,N_29009,N_27729);
nand UO_1795 (O_1795,N_28134,N_27372);
xor UO_1796 (O_1796,N_28879,N_28392);
and UO_1797 (O_1797,N_28876,N_28060);
nand UO_1798 (O_1798,N_28143,N_28134);
nor UO_1799 (O_1799,N_27842,N_28931);
nand UO_1800 (O_1800,N_28899,N_29522);
nand UO_1801 (O_1801,N_28462,N_27622);
or UO_1802 (O_1802,N_27569,N_29629);
nand UO_1803 (O_1803,N_28595,N_27977);
nand UO_1804 (O_1804,N_27386,N_27228);
or UO_1805 (O_1805,N_27658,N_28495);
or UO_1806 (O_1806,N_27411,N_28633);
and UO_1807 (O_1807,N_27907,N_27136);
nand UO_1808 (O_1808,N_28909,N_27101);
and UO_1809 (O_1809,N_28211,N_27786);
and UO_1810 (O_1810,N_29707,N_27092);
nand UO_1811 (O_1811,N_28450,N_29667);
nand UO_1812 (O_1812,N_28708,N_27019);
xnor UO_1813 (O_1813,N_27111,N_28988);
nand UO_1814 (O_1814,N_29050,N_29433);
nand UO_1815 (O_1815,N_29155,N_28341);
and UO_1816 (O_1816,N_27131,N_29818);
nand UO_1817 (O_1817,N_27692,N_29068);
or UO_1818 (O_1818,N_28080,N_29856);
and UO_1819 (O_1819,N_28426,N_29332);
and UO_1820 (O_1820,N_27566,N_27198);
and UO_1821 (O_1821,N_28106,N_28563);
nand UO_1822 (O_1822,N_29369,N_27641);
and UO_1823 (O_1823,N_29378,N_28607);
or UO_1824 (O_1824,N_28297,N_29512);
nand UO_1825 (O_1825,N_28377,N_29966);
and UO_1826 (O_1826,N_27577,N_29187);
or UO_1827 (O_1827,N_27536,N_27740);
nor UO_1828 (O_1828,N_28247,N_27653);
nand UO_1829 (O_1829,N_29655,N_28082);
nor UO_1830 (O_1830,N_29402,N_29031);
or UO_1831 (O_1831,N_27440,N_28001);
nand UO_1832 (O_1832,N_27917,N_29607);
xor UO_1833 (O_1833,N_28143,N_28205);
nor UO_1834 (O_1834,N_27112,N_29386);
xnor UO_1835 (O_1835,N_29125,N_27691);
and UO_1836 (O_1836,N_27244,N_29315);
and UO_1837 (O_1837,N_29983,N_27384);
xor UO_1838 (O_1838,N_28613,N_27034);
xor UO_1839 (O_1839,N_28200,N_27271);
and UO_1840 (O_1840,N_28800,N_27233);
or UO_1841 (O_1841,N_28633,N_28725);
xnor UO_1842 (O_1842,N_27208,N_28913);
and UO_1843 (O_1843,N_27430,N_28035);
nor UO_1844 (O_1844,N_28391,N_29561);
xnor UO_1845 (O_1845,N_29749,N_28716);
xor UO_1846 (O_1846,N_27087,N_28754);
and UO_1847 (O_1847,N_27793,N_29726);
nor UO_1848 (O_1848,N_27964,N_28002);
or UO_1849 (O_1849,N_28699,N_28625);
or UO_1850 (O_1850,N_28483,N_27688);
and UO_1851 (O_1851,N_27677,N_27714);
and UO_1852 (O_1852,N_28760,N_28720);
or UO_1853 (O_1853,N_29598,N_28843);
or UO_1854 (O_1854,N_27163,N_27222);
nor UO_1855 (O_1855,N_27995,N_27926);
or UO_1856 (O_1856,N_29465,N_28447);
and UO_1857 (O_1857,N_29847,N_29035);
or UO_1858 (O_1858,N_28754,N_28266);
nor UO_1859 (O_1859,N_29012,N_28452);
or UO_1860 (O_1860,N_28425,N_28118);
and UO_1861 (O_1861,N_29718,N_29912);
and UO_1862 (O_1862,N_27645,N_29668);
nand UO_1863 (O_1863,N_27917,N_29471);
nor UO_1864 (O_1864,N_28031,N_29217);
xnor UO_1865 (O_1865,N_27119,N_29072);
and UO_1866 (O_1866,N_28769,N_27355);
or UO_1867 (O_1867,N_27495,N_27569);
or UO_1868 (O_1868,N_27350,N_27524);
nor UO_1869 (O_1869,N_27755,N_27216);
or UO_1870 (O_1870,N_28594,N_28898);
nand UO_1871 (O_1871,N_29085,N_28753);
nand UO_1872 (O_1872,N_27183,N_27789);
and UO_1873 (O_1873,N_27787,N_28381);
xnor UO_1874 (O_1874,N_27139,N_28536);
nand UO_1875 (O_1875,N_29888,N_29996);
nand UO_1876 (O_1876,N_28085,N_28608);
nand UO_1877 (O_1877,N_28745,N_29995);
nand UO_1878 (O_1878,N_28696,N_27959);
nand UO_1879 (O_1879,N_27129,N_28436);
xor UO_1880 (O_1880,N_29040,N_28163);
nand UO_1881 (O_1881,N_29165,N_29393);
nor UO_1882 (O_1882,N_29041,N_29592);
nor UO_1883 (O_1883,N_28703,N_28734);
or UO_1884 (O_1884,N_27232,N_27002);
nor UO_1885 (O_1885,N_27801,N_27419);
or UO_1886 (O_1886,N_29457,N_27721);
or UO_1887 (O_1887,N_29896,N_29269);
nor UO_1888 (O_1888,N_27748,N_29016);
and UO_1889 (O_1889,N_29104,N_29342);
xor UO_1890 (O_1890,N_29536,N_29232);
or UO_1891 (O_1891,N_28820,N_29293);
and UO_1892 (O_1892,N_29822,N_28375);
or UO_1893 (O_1893,N_28845,N_29576);
and UO_1894 (O_1894,N_27147,N_28401);
xnor UO_1895 (O_1895,N_29253,N_27660);
xnor UO_1896 (O_1896,N_29913,N_29153);
or UO_1897 (O_1897,N_27150,N_29328);
or UO_1898 (O_1898,N_29023,N_27909);
nand UO_1899 (O_1899,N_29550,N_29170);
nor UO_1900 (O_1900,N_27127,N_28416);
nand UO_1901 (O_1901,N_27696,N_27950);
nand UO_1902 (O_1902,N_27304,N_29020);
nand UO_1903 (O_1903,N_27190,N_29881);
nor UO_1904 (O_1904,N_29445,N_27754);
and UO_1905 (O_1905,N_27662,N_29662);
or UO_1906 (O_1906,N_27028,N_27364);
and UO_1907 (O_1907,N_29585,N_28394);
nor UO_1908 (O_1908,N_29267,N_28269);
nor UO_1909 (O_1909,N_29331,N_29437);
xnor UO_1910 (O_1910,N_29243,N_29811);
and UO_1911 (O_1911,N_29762,N_27859);
nand UO_1912 (O_1912,N_28877,N_29888);
and UO_1913 (O_1913,N_27615,N_29489);
xnor UO_1914 (O_1914,N_29205,N_29031);
nand UO_1915 (O_1915,N_27162,N_29439);
or UO_1916 (O_1916,N_29876,N_28389);
xnor UO_1917 (O_1917,N_27452,N_29491);
xnor UO_1918 (O_1918,N_28592,N_29766);
xnor UO_1919 (O_1919,N_28871,N_28320);
or UO_1920 (O_1920,N_29360,N_29909);
and UO_1921 (O_1921,N_27917,N_27222);
xor UO_1922 (O_1922,N_28668,N_28291);
or UO_1923 (O_1923,N_28126,N_27953);
and UO_1924 (O_1924,N_28832,N_27096);
nand UO_1925 (O_1925,N_29753,N_27850);
xor UO_1926 (O_1926,N_29475,N_29098);
nand UO_1927 (O_1927,N_27879,N_29918);
and UO_1928 (O_1928,N_28614,N_28394);
and UO_1929 (O_1929,N_27293,N_27659);
xnor UO_1930 (O_1930,N_29632,N_29362);
nand UO_1931 (O_1931,N_29819,N_29773);
and UO_1932 (O_1932,N_27925,N_29050);
xnor UO_1933 (O_1933,N_27990,N_28253);
or UO_1934 (O_1934,N_29770,N_29293);
nand UO_1935 (O_1935,N_27279,N_27044);
nor UO_1936 (O_1936,N_29205,N_28171);
nor UO_1937 (O_1937,N_29487,N_28327);
or UO_1938 (O_1938,N_28858,N_27424);
and UO_1939 (O_1939,N_29757,N_28021);
nand UO_1940 (O_1940,N_28874,N_29947);
or UO_1941 (O_1941,N_27965,N_28653);
or UO_1942 (O_1942,N_29833,N_28555);
nand UO_1943 (O_1943,N_28954,N_28244);
and UO_1944 (O_1944,N_28816,N_29706);
or UO_1945 (O_1945,N_28914,N_29856);
nor UO_1946 (O_1946,N_27675,N_28998);
and UO_1947 (O_1947,N_28267,N_29451);
nand UO_1948 (O_1948,N_27015,N_28260);
nand UO_1949 (O_1949,N_28147,N_27955);
nor UO_1950 (O_1950,N_29077,N_27850);
xnor UO_1951 (O_1951,N_28922,N_28543);
xor UO_1952 (O_1952,N_28038,N_29718);
xnor UO_1953 (O_1953,N_29573,N_28047);
xor UO_1954 (O_1954,N_29111,N_28217);
or UO_1955 (O_1955,N_27071,N_28115);
nand UO_1956 (O_1956,N_27999,N_28035);
or UO_1957 (O_1957,N_28499,N_27194);
and UO_1958 (O_1958,N_28573,N_28096);
nor UO_1959 (O_1959,N_28895,N_28942);
nor UO_1960 (O_1960,N_28734,N_28382);
or UO_1961 (O_1961,N_27535,N_29635);
or UO_1962 (O_1962,N_29417,N_27731);
and UO_1963 (O_1963,N_27573,N_29193);
nor UO_1964 (O_1964,N_28907,N_28501);
and UO_1965 (O_1965,N_28453,N_29839);
xor UO_1966 (O_1966,N_28964,N_27161);
nand UO_1967 (O_1967,N_28313,N_27824);
and UO_1968 (O_1968,N_27090,N_29956);
or UO_1969 (O_1969,N_28721,N_27226);
or UO_1970 (O_1970,N_29697,N_28907);
xnor UO_1971 (O_1971,N_27604,N_28483);
or UO_1972 (O_1972,N_27205,N_29750);
or UO_1973 (O_1973,N_28468,N_29237);
xnor UO_1974 (O_1974,N_27042,N_27209);
and UO_1975 (O_1975,N_29806,N_28662);
or UO_1976 (O_1976,N_28172,N_27649);
nand UO_1977 (O_1977,N_27515,N_28385);
nor UO_1978 (O_1978,N_29919,N_29732);
xnor UO_1979 (O_1979,N_27415,N_28389);
nand UO_1980 (O_1980,N_29172,N_29187);
or UO_1981 (O_1981,N_29680,N_28484);
xnor UO_1982 (O_1982,N_29475,N_27793);
nand UO_1983 (O_1983,N_27023,N_28607);
xnor UO_1984 (O_1984,N_29533,N_29911);
nor UO_1985 (O_1985,N_27353,N_27166);
nand UO_1986 (O_1986,N_28371,N_27449);
and UO_1987 (O_1987,N_27874,N_29064);
nand UO_1988 (O_1988,N_27230,N_28594);
xor UO_1989 (O_1989,N_28179,N_27237);
xnor UO_1990 (O_1990,N_28828,N_29802);
and UO_1991 (O_1991,N_27504,N_29330);
nand UO_1992 (O_1992,N_28607,N_28200);
nand UO_1993 (O_1993,N_28392,N_27925);
nor UO_1994 (O_1994,N_27433,N_28592);
and UO_1995 (O_1995,N_28437,N_28979);
and UO_1996 (O_1996,N_28167,N_27562);
xnor UO_1997 (O_1997,N_27148,N_27095);
or UO_1998 (O_1998,N_28167,N_28627);
nor UO_1999 (O_1999,N_27455,N_27033);
xor UO_2000 (O_2000,N_27913,N_27163);
nor UO_2001 (O_2001,N_28026,N_29797);
xor UO_2002 (O_2002,N_27770,N_29973);
xnor UO_2003 (O_2003,N_28618,N_29457);
and UO_2004 (O_2004,N_27917,N_29606);
and UO_2005 (O_2005,N_28779,N_27532);
and UO_2006 (O_2006,N_27101,N_28659);
nor UO_2007 (O_2007,N_29408,N_29753);
nand UO_2008 (O_2008,N_27487,N_28989);
and UO_2009 (O_2009,N_28392,N_29346);
and UO_2010 (O_2010,N_27956,N_27551);
nand UO_2011 (O_2011,N_28079,N_28785);
nand UO_2012 (O_2012,N_27061,N_29635);
nor UO_2013 (O_2013,N_29820,N_29287);
nand UO_2014 (O_2014,N_28913,N_27832);
xnor UO_2015 (O_2015,N_29324,N_29232);
nor UO_2016 (O_2016,N_29214,N_29017);
nand UO_2017 (O_2017,N_27466,N_27793);
nor UO_2018 (O_2018,N_29488,N_28322);
and UO_2019 (O_2019,N_28221,N_27968);
or UO_2020 (O_2020,N_29297,N_28412);
or UO_2021 (O_2021,N_28364,N_28761);
xnor UO_2022 (O_2022,N_28313,N_27888);
nor UO_2023 (O_2023,N_28237,N_27145);
xnor UO_2024 (O_2024,N_28806,N_29019);
nor UO_2025 (O_2025,N_29169,N_28639);
nor UO_2026 (O_2026,N_27250,N_28980);
and UO_2027 (O_2027,N_29909,N_27654);
and UO_2028 (O_2028,N_29181,N_29644);
xor UO_2029 (O_2029,N_29379,N_29989);
or UO_2030 (O_2030,N_27249,N_28043);
nand UO_2031 (O_2031,N_27736,N_29685);
nor UO_2032 (O_2032,N_29939,N_29508);
nand UO_2033 (O_2033,N_29541,N_27233);
nand UO_2034 (O_2034,N_27799,N_29814);
nor UO_2035 (O_2035,N_27135,N_28145);
xnor UO_2036 (O_2036,N_29316,N_28036);
and UO_2037 (O_2037,N_29906,N_27897);
nand UO_2038 (O_2038,N_29338,N_27327);
xnor UO_2039 (O_2039,N_29055,N_28985);
or UO_2040 (O_2040,N_28037,N_27217);
nor UO_2041 (O_2041,N_28390,N_27836);
xor UO_2042 (O_2042,N_28042,N_27288);
and UO_2043 (O_2043,N_27982,N_28362);
nand UO_2044 (O_2044,N_27846,N_27525);
nand UO_2045 (O_2045,N_27267,N_28081);
and UO_2046 (O_2046,N_28693,N_27189);
or UO_2047 (O_2047,N_28218,N_29565);
nand UO_2048 (O_2048,N_29632,N_27830);
or UO_2049 (O_2049,N_27777,N_28290);
and UO_2050 (O_2050,N_27438,N_28124);
or UO_2051 (O_2051,N_27706,N_29810);
nand UO_2052 (O_2052,N_28788,N_28852);
or UO_2053 (O_2053,N_27951,N_27016);
xnor UO_2054 (O_2054,N_28328,N_29257);
nor UO_2055 (O_2055,N_29811,N_28923);
xnor UO_2056 (O_2056,N_28751,N_28780);
nor UO_2057 (O_2057,N_28883,N_28955);
or UO_2058 (O_2058,N_28647,N_28567);
nand UO_2059 (O_2059,N_27016,N_29607);
xor UO_2060 (O_2060,N_27131,N_27161);
nor UO_2061 (O_2061,N_29977,N_29193);
nor UO_2062 (O_2062,N_28600,N_27463);
and UO_2063 (O_2063,N_27171,N_27753);
and UO_2064 (O_2064,N_29870,N_29194);
and UO_2065 (O_2065,N_27462,N_29390);
xor UO_2066 (O_2066,N_29213,N_27311);
xnor UO_2067 (O_2067,N_28529,N_27020);
and UO_2068 (O_2068,N_29477,N_29372);
nor UO_2069 (O_2069,N_27375,N_27525);
nand UO_2070 (O_2070,N_29563,N_27354);
and UO_2071 (O_2071,N_29264,N_28203);
or UO_2072 (O_2072,N_27278,N_28541);
and UO_2073 (O_2073,N_28606,N_29018);
xnor UO_2074 (O_2074,N_27495,N_28224);
nand UO_2075 (O_2075,N_29861,N_29981);
nand UO_2076 (O_2076,N_28181,N_28589);
and UO_2077 (O_2077,N_28429,N_28621);
xor UO_2078 (O_2078,N_27784,N_28208);
and UO_2079 (O_2079,N_29435,N_29688);
and UO_2080 (O_2080,N_27243,N_29053);
and UO_2081 (O_2081,N_27689,N_27432);
nor UO_2082 (O_2082,N_28378,N_29162);
nand UO_2083 (O_2083,N_27782,N_28681);
nand UO_2084 (O_2084,N_28674,N_27811);
nand UO_2085 (O_2085,N_27296,N_29056);
nand UO_2086 (O_2086,N_29529,N_29675);
nand UO_2087 (O_2087,N_27462,N_28128);
and UO_2088 (O_2088,N_27063,N_27876);
nor UO_2089 (O_2089,N_29444,N_28523);
xnor UO_2090 (O_2090,N_27405,N_28367);
and UO_2091 (O_2091,N_28357,N_29204);
nand UO_2092 (O_2092,N_27241,N_28811);
nand UO_2093 (O_2093,N_28646,N_28088);
or UO_2094 (O_2094,N_28086,N_27408);
nand UO_2095 (O_2095,N_29327,N_29350);
nor UO_2096 (O_2096,N_28287,N_27692);
xor UO_2097 (O_2097,N_29062,N_28852);
xor UO_2098 (O_2098,N_29275,N_27146);
or UO_2099 (O_2099,N_29925,N_28503);
xor UO_2100 (O_2100,N_27370,N_28494);
nand UO_2101 (O_2101,N_29628,N_28304);
nand UO_2102 (O_2102,N_28126,N_28621);
or UO_2103 (O_2103,N_27255,N_28508);
nand UO_2104 (O_2104,N_28947,N_27086);
nand UO_2105 (O_2105,N_27881,N_29034);
or UO_2106 (O_2106,N_27820,N_27202);
nand UO_2107 (O_2107,N_27348,N_28595);
nor UO_2108 (O_2108,N_27019,N_29141);
nand UO_2109 (O_2109,N_28131,N_28911);
and UO_2110 (O_2110,N_29866,N_27575);
nor UO_2111 (O_2111,N_29894,N_29954);
nand UO_2112 (O_2112,N_27383,N_29505);
xnor UO_2113 (O_2113,N_29248,N_28535);
and UO_2114 (O_2114,N_28602,N_29888);
xnor UO_2115 (O_2115,N_29034,N_27996);
nor UO_2116 (O_2116,N_29422,N_29583);
and UO_2117 (O_2117,N_28353,N_27010);
nor UO_2118 (O_2118,N_28916,N_29675);
nand UO_2119 (O_2119,N_27120,N_28682);
or UO_2120 (O_2120,N_27641,N_27864);
and UO_2121 (O_2121,N_29156,N_29556);
nand UO_2122 (O_2122,N_28830,N_27280);
nor UO_2123 (O_2123,N_29329,N_29901);
nor UO_2124 (O_2124,N_29028,N_29288);
or UO_2125 (O_2125,N_28247,N_29759);
xnor UO_2126 (O_2126,N_28393,N_29023);
nand UO_2127 (O_2127,N_28426,N_28455);
nand UO_2128 (O_2128,N_27692,N_28994);
or UO_2129 (O_2129,N_27625,N_27072);
nor UO_2130 (O_2130,N_27547,N_28096);
nor UO_2131 (O_2131,N_28431,N_29579);
xor UO_2132 (O_2132,N_27204,N_27373);
or UO_2133 (O_2133,N_29606,N_28483);
nand UO_2134 (O_2134,N_27417,N_28970);
or UO_2135 (O_2135,N_28743,N_29063);
nand UO_2136 (O_2136,N_29445,N_28511);
or UO_2137 (O_2137,N_28538,N_27547);
or UO_2138 (O_2138,N_28646,N_28650);
nand UO_2139 (O_2139,N_27932,N_29578);
nor UO_2140 (O_2140,N_28587,N_28342);
or UO_2141 (O_2141,N_27274,N_29266);
and UO_2142 (O_2142,N_27483,N_27671);
nor UO_2143 (O_2143,N_27447,N_29412);
and UO_2144 (O_2144,N_27788,N_28948);
nand UO_2145 (O_2145,N_27554,N_28618);
xnor UO_2146 (O_2146,N_27820,N_27519);
and UO_2147 (O_2147,N_28773,N_28631);
xor UO_2148 (O_2148,N_27150,N_27208);
and UO_2149 (O_2149,N_28729,N_28467);
nor UO_2150 (O_2150,N_29111,N_27791);
nor UO_2151 (O_2151,N_28500,N_29056);
and UO_2152 (O_2152,N_29417,N_28536);
nor UO_2153 (O_2153,N_28778,N_27517);
xor UO_2154 (O_2154,N_28257,N_27975);
or UO_2155 (O_2155,N_29039,N_27627);
nand UO_2156 (O_2156,N_28045,N_27858);
nor UO_2157 (O_2157,N_28454,N_29174);
and UO_2158 (O_2158,N_29205,N_29712);
nand UO_2159 (O_2159,N_27042,N_29161);
and UO_2160 (O_2160,N_29598,N_27665);
xor UO_2161 (O_2161,N_28994,N_29117);
nand UO_2162 (O_2162,N_29839,N_29941);
xor UO_2163 (O_2163,N_29509,N_29036);
or UO_2164 (O_2164,N_27686,N_27079);
nor UO_2165 (O_2165,N_28006,N_27434);
nor UO_2166 (O_2166,N_27030,N_27726);
and UO_2167 (O_2167,N_29275,N_29313);
nor UO_2168 (O_2168,N_29057,N_29475);
xnor UO_2169 (O_2169,N_29691,N_28671);
or UO_2170 (O_2170,N_27603,N_28765);
xnor UO_2171 (O_2171,N_29801,N_27976);
xor UO_2172 (O_2172,N_28038,N_27914);
nand UO_2173 (O_2173,N_27316,N_28777);
nor UO_2174 (O_2174,N_28241,N_29905);
nand UO_2175 (O_2175,N_27033,N_27026);
nand UO_2176 (O_2176,N_27719,N_29165);
or UO_2177 (O_2177,N_27838,N_28392);
or UO_2178 (O_2178,N_27429,N_29378);
nand UO_2179 (O_2179,N_29957,N_27038);
xor UO_2180 (O_2180,N_29921,N_28233);
xnor UO_2181 (O_2181,N_29068,N_28259);
nand UO_2182 (O_2182,N_29667,N_27463);
nand UO_2183 (O_2183,N_27547,N_29971);
or UO_2184 (O_2184,N_28461,N_29958);
and UO_2185 (O_2185,N_27191,N_27613);
or UO_2186 (O_2186,N_28690,N_29508);
nor UO_2187 (O_2187,N_28029,N_27947);
and UO_2188 (O_2188,N_28285,N_27919);
nand UO_2189 (O_2189,N_29529,N_27380);
nor UO_2190 (O_2190,N_29844,N_28939);
nor UO_2191 (O_2191,N_27021,N_28347);
or UO_2192 (O_2192,N_29713,N_28602);
nor UO_2193 (O_2193,N_29877,N_29663);
xnor UO_2194 (O_2194,N_29486,N_27541);
or UO_2195 (O_2195,N_27934,N_29477);
nor UO_2196 (O_2196,N_28409,N_28567);
nor UO_2197 (O_2197,N_29648,N_29129);
nand UO_2198 (O_2198,N_27622,N_28963);
xor UO_2199 (O_2199,N_27322,N_27890);
nand UO_2200 (O_2200,N_29900,N_29893);
xor UO_2201 (O_2201,N_27725,N_29353);
nand UO_2202 (O_2202,N_29957,N_29337);
and UO_2203 (O_2203,N_27378,N_27832);
nor UO_2204 (O_2204,N_27400,N_28140);
xnor UO_2205 (O_2205,N_29188,N_29130);
nor UO_2206 (O_2206,N_28199,N_27970);
nor UO_2207 (O_2207,N_29529,N_27312);
xor UO_2208 (O_2208,N_28945,N_29924);
xnor UO_2209 (O_2209,N_28600,N_28312);
nand UO_2210 (O_2210,N_29693,N_28389);
nor UO_2211 (O_2211,N_29808,N_27667);
and UO_2212 (O_2212,N_27504,N_28592);
xor UO_2213 (O_2213,N_28351,N_28857);
xnor UO_2214 (O_2214,N_27938,N_28922);
nor UO_2215 (O_2215,N_28469,N_27582);
and UO_2216 (O_2216,N_27136,N_27262);
and UO_2217 (O_2217,N_27473,N_29428);
nand UO_2218 (O_2218,N_28786,N_29561);
or UO_2219 (O_2219,N_29770,N_27646);
nand UO_2220 (O_2220,N_29517,N_27286);
and UO_2221 (O_2221,N_29909,N_28905);
or UO_2222 (O_2222,N_27314,N_28443);
or UO_2223 (O_2223,N_29420,N_28669);
xnor UO_2224 (O_2224,N_27501,N_28192);
and UO_2225 (O_2225,N_29751,N_27343);
or UO_2226 (O_2226,N_27023,N_27051);
and UO_2227 (O_2227,N_27173,N_27721);
and UO_2228 (O_2228,N_28662,N_29992);
xor UO_2229 (O_2229,N_27444,N_27107);
xnor UO_2230 (O_2230,N_27529,N_27151);
nand UO_2231 (O_2231,N_28574,N_29765);
and UO_2232 (O_2232,N_27371,N_27689);
nand UO_2233 (O_2233,N_27860,N_29549);
xnor UO_2234 (O_2234,N_29832,N_28125);
nand UO_2235 (O_2235,N_27792,N_27776);
nand UO_2236 (O_2236,N_28167,N_27899);
xor UO_2237 (O_2237,N_27623,N_28700);
xnor UO_2238 (O_2238,N_29805,N_28740);
nor UO_2239 (O_2239,N_28707,N_28353);
or UO_2240 (O_2240,N_27240,N_29175);
xnor UO_2241 (O_2241,N_27943,N_28425);
xnor UO_2242 (O_2242,N_29929,N_29164);
nand UO_2243 (O_2243,N_28880,N_29783);
or UO_2244 (O_2244,N_27401,N_28913);
xor UO_2245 (O_2245,N_27893,N_27318);
or UO_2246 (O_2246,N_29741,N_27395);
nand UO_2247 (O_2247,N_27117,N_27254);
or UO_2248 (O_2248,N_29043,N_29209);
nor UO_2249 (O_2249,N_27684,N_28380);
nor UO_2250 (O_2250,N_27391,N_27866);
nand UO_2251 (O_2251,N_27366,N_28788);
xor UO_2252 (O_2252,N_28550,N_28015);
nand UO_2253 (O_2253,N_29880,N_27356);
or UO_2254 (O_2254,N_28257,N_28976);
xor UO_2255 (O_2255,N_27054,N_28729);
and UO_2256 (O_2256,N_27004,N_29263);
xnor UO_2257 (O_2257,N_27076,N_28327);
nand UO_2258 (O_2258,N_28098,N_27078);
nor UO_2259 (O_2259,N_29247,N_29096);
and UO_2260 (O_2260,N_29946,N_28106);
and UO_2261 (O_2261,N_28602,N_27162);
or UO_2262 (O_2262,N_29212,N_28997);
nor UO_2263 (O_2263,N_29228,N_27778);
nor UO_2264 (O_2264,N_29760,N_28495);
nor UO_2265 (O_2265,N_28411,N_28819);
or UO_2266 (O_2266,N_28015,N_27961);
nor UO_2267 (O_2267,N_29928,N_28456);
or UO_2268 (O_2268,N_29649,N_27403);
xnor UO_2269 (O_2269,N_28491,N_28401);
nor UO_2270 (O_2270,N_28660,N_28720);
xnor UO_2271 (O_2271,N_27420,N_28064);
nor UO_2272 (O_2272,N_28971,N_28906);
nor UO_2273 (O_2273,N_29273,N_29602);
nor UO_2274 (O_2274,N_27782,N_27406);
nand UO_2275 (O_2275,N_27249,N_28569);
xnor UO_2276 (O_2276,N_28055,N_29065);
and UO_2277 (O_2277,N_27103,N_29202);
nor UO_2278 (O_2278,N_27230,N_28501);
and UO_2279 (O_2279,N_27532,N_29201);
or UO_2280 (O_2280,N_28376,N_27873);
xnor UO_2281 (O_2281,N_27038,N_27008);
and UO_2282 (O_2282,N_28201,N_29069);
and UO_2283 (O_2283,N_29562,N_27716);
nor UO_2284 (O_2284,N_27656,N_29331);
xnor UO_2285 (O_2285,N_27017,N_27834);
and UO_2286 (O_2286,N_28711,N_28102);
nand UO_2287 (O_2287,N_29008,N_27119);
or UO_2288 (O_2288,N_27061,N_27646);
nor UO_2289 (O_2289,N_27519,N_27270);
xor UO_2290 (O_2290,N_27997,N_28902);
and UO_2291 (O_2291,N_29834,N_28883);
xor UO_2292 (O_2292,N_28543,N_27895);
or UO_2293 (O_2293,N_28447,N_28580);
nor UO_2294 (O_2294,N_29243,N_28677);
nor UO_2295 (O_2295,N_29230,N_27111);
or UO_2296 (O_2296,N_28718,N_27627);
nor UO_2297 (O_2297,N_27732,N_29302);
xnor UO_2298 (O_2298,N_28818,N_28156);
nor UO_2299 (O_2299,N_28362,N_28013);
xnor UO_2300 (O_2300,N_29877,N_28435);
nor UO_2301 (O_2301,N_27621,N_29554);
nor UO_2302 (O_2302,N_27045,N_28156);
xnor UO_2303 (O_2303,N_29641,N_29103);
nand UO_2304 (O_2304,N_29152,N_27339);
or UO_2305 (O_2305,N_27731,N_28494);
or UO_2306 (O_2306,N_27159,N_28626);
and UO_2307 (O_2307,N_27244,N_29973);
xor UO_2308 (O_2308,N_27721,N_27003);
nor UO_2309 (O_2309,N_27464,N_27486);
or UO_2310 (O_2310,N_28813,N_29438);
nand UO_2311 (O_2311,N_28935,N_29819);
or UO_2312 (O_2312,N_27642,N_28476);
nor UO_2313 (O_2313,N_28792,N_27673);
nor UO_2314 (O_2314,N_28271,N_28503);
xor UO_2315 (O_2315,N_29666,N_27642);
and UO_2316 (O_2316,N_27691,N_29081);
nor UO_2317 (O_2317,N_27229,N_29872);
nand UO_2318 (O_2318,N_28619,N_27891);
or UO_2319 (O_2319,N_29854,N_29011);
xor UO_2320 (O_2320,N_27730,N_29829);
and UO_2321 (O_2321,N_29480,N_28456);
or UO_2322 (O_2322,N_29953,N_27245);
and UO_2323 (O_2323,N_29388,N_29582);
xnor UO_2324 (O_2324,N_28572,N_28490);
xnor UO_2325 (O_2325,N_28534,N_29698);
xor UO_2326 (O_2326,N_28698,N_27296);
nor UO_2327 (O_2327,N_27554,N_29445);
xnor UO_2328 (O_2328,N_29019,N_28291);
nand UO_2329 (O_2329,N_29874,N_27939);
or UO_2330 (O_2330,N_27698,N_27897);
nand UO_2331 (O_2331,N_28939,N_28698);
and UO_2332 (O_2332,N_28178,N_28064);
xor UO_2333 (O_2333,N_29155,N_29339);
nor UO_2334 (O_2334,N_29805,N_29228);
nand UO_2335 (O_2335,N_28194,N_27037);
or UO_2336 (O_2336,N_29440,N_28881);
and UO_2337 (O_2337,N_28612,N_28573);
xnor UO_2338 (O_2338,N_28921,N_29956);
xor UO_2339 (O_2339,N_28249,N_29976);
xor UO_2340 (O_2340,N_29287,N_27250);
or UO_2341 (O_2341,N_29009,N_29311);
or UO_2342 (O_2342,N_28385,N_27937);
and UO_2343 (O_2343,N_28932,N_27842);
nand UO_2344 (O_2344,N_29754,N_27524);
nor UO_2345 (O_2345,N_29624,N_29723);
nand UO_2346 (O_2346,N_27916,N_27074);
nand UO_2347 (O_2347,N_27082,N_27872);
and UO_2348 (O_2348,N_29456,N_27316);
or UO_2349 (O_2349,N_29684,N_29517);
and UO_2350 (O_2350,N_28529,N_27297);
xor UO_2351 (O_2351,N_28278,N_29936);
or UO_2352 (O_2352,N_29544,N_29322);
or UO_2353 (O_2353,N_29105,N_29129);
nand UO_2354 (O_2354,N_27023,N_28632);
nand UO_2355 (O_2355,N_28208,N_27320);
and UO_2356 (O_2356,N_28345,N_29022);
xnor UO_2357 (O_2357,N_27902,N_28801);
xnor UO_2358 (O_2358,N_28699,N_29181);
and UO_2359 (O_2359,N_29701,N_28819);
nand UO_2360 (O_2360,N_28377,N_28884);
or UO_2361 (O_2361,N_27721,N_28067);
xnor UO_2362 (O_2362,N_28007,N_29120);
or UO_2363 (O_2363,N_29930,N_27621);
and UO_2364 (O_2364,N_29168,N_29181);
xnor UO_2365 (O_2365,N_28402,N_27739);
or UO_2366 (O_2366,N_28160,N_29412);
xor UO_2367 (O_2367,N_28820,N_27560);
xnor UO_2368 (O_2368,N_27513,N_29368);
and UO_2369 (O_2369,N_28429,N_28840);
xnor UO_2370 (O_2370,N_29992,N_29845);
nor UO_2371 (O_2371,N_27038,N_28350);
and UO_2372 (O_2372,N_27784,N_27463);
nand UO_2373 (O_2373,N_29904,N_28660);
and UO_2374 (O_2374,N_28562,N_29787);
and UO_2375 (O_2375,N_28961,N_27589);
nor UO_2376 (O_2376,N_27360,N_28368);
and UO_2377 (O_2377,N_28210,N_27220);
nor UO_2378 (O_2378,N_28544,N_28315);
or UO_2379 (O_2379,N_29493,N_29481);
and UO_2380 (O_2380,N_29173,N_28152);
nor UO_2381 (O_2381,N_28197,N_27293);
or UO_2382 (O_2382,N_28248,N_28427);
nand UO_2383 (O_2383,N_29965,N_28719);
nand UO_2384 (O_2384,N_28543,N_29812);
nand UO_2385 (O_2385,N_27231,N_27867);
nor UO_2386 (O_2386,N_28292,N_29209);
nor UO_2387 (O_2387,N_27808,N_27629);
nor UO_2388 (O_2388,N_27248,N_29939);
and UO_2389 (O_2389,N_29203,N_27409);
nand UO_2390 (O_2390,N_28512,N_29979);
and UO_2391 (O_2391,N_28508,N_28573);
or UO_2392 (O_2392,N_27045,N_29296);
nand UO_2393 (O_2393,N_27736,N_29846);
nor UO_2394 (O_2394,N_28829,N_27193);
and UO_2395 (O_2395,N_29639,N_28268);
xnor UO_2396 (O_2396,N_28932,N_29205);
nand UO_2397 (O_2397,N_29531,N_28131);
and UO_2398 (O_2398,N_28104,N_28990);
xnor UO_2399 (O_2399,N_29073,N_29233);
xor UO_2400 (O_2400,N_27082,N_27115);
nor UO_2401 (O_2401,N_27110,N_28105);
nand UO_2402 (O_2402,N_27059,N_27609);
or UO_2403 (O_2403,N_28781,N_27646);
or UO_2404 (O_2404,N_28309,N_28152);
and UO_2405 (O_2405,N_28837,N_27440);
nor UO_2406 (O_2406,N_27735,N_29650);
and UO_2407 (O_2407,N_28032,N_29410);
nor UO_2408 (O_2408,N_29177,N_29616);
and UO_2409 (O_2409,N_27634,N_27077);
or UO_2410 (O_2410,N_29347,N_28503);
nand UO_2411 (O_2411,N_27578,N_28696);
and UO_2412 (O_2412,N_28443,N_27775);
xor UO_2413 (O_2413,N_27198,N_27088);
nor UO_2414 (O_2414,N_27081,N_27281);
or UO_2415 (O_2415,N_27227,N_27498);
nor UO_2416 (O_2416,N_28662,N_28687);
xnor UO_2417 (O_2417,N_28655,N_27192);
nand UO_2418 (O_2418,N_29618,N_28163);
nor UO_2419 (O_2419,N_27085,N_28848);
or UO_2420 (O_2420,N_27028,N_28626);
and UO_2421 (O_2421,N_28342,N_28785);
nand UO_2422 (O_2422,N_27148,N_29358);
and UO_2423 (O_2423,N_27897,N_27247);
or UO_2424 (O_2424,N_27624,N_28501);
nand UO_2425 (O_2425,N_29806,N_29390);
xnor UO_2426 (O_2426,N_27401,N_27594);
nand UO_2427 (O_2427,N_29324,N_27214);
nand UO_2428 (O_2428,N_27251,N_29563);
or UO_2429 (O_2429,N_29420,N_28960);
xor UO_2430 (O_2430,N_29854,N_27611);
nand UO_2431 (O_2431,N_29394,N_28544);
or UO_2432 (O_2432,N_29106,N_29578);
and UO_2433 (O_2433,N_29796,N_28773);
nor UO_2434 (O_2434,N_28588,N_29148);
xnor UO_2435 (O_2435,N_29418,N_27765);
or UO_2436 (O_2436,N_29108,N_27902);
xor UO_2437 (O_2437,N_28596,N_29630);
and UO_2438 (O_2438,N_28702,N_27045);
nor UO_2439 (O_2439,N_28019,N_28327);
nor UO_2440 (O_2440,N_29065,N_27125);
or UO_2441 (O_2441,N_27760,N_28939);
or UO_2442 (O_2442,N_28249,N_29432);
xnor UO_2443 (O_2443,N_28538,N_29750);
or UO_2444 (O_2444,N_28422,N_27997);
or UO_2445 (O_2445,N_28158,N_28071);
or UO_2446 (O_2446,N_29448,N_27041);
or UO_2447 (O_2447,N_28920,N_27895);
nand UO_2448 (O_2448,N_28138,N_29575);
or UO_2449 (O_2449,N_29905,N_28055);
and UO_2450 (O_2450,N_27061,N_27925);
xor UO_2451 (O_2451,N_28277,N_29431);
nor UO_2452 (O_2452,N_28239,N_28990);
nor UO_2453 (O_2453,N_27253,N_27463);
and UO_2454 (O_2454,N_27285,N_29178);
or UO_2455 (O_2455,N_27153,N_27680);
nand UO_2456 (O_2456,N_27059,N_27417);
xor UO_2457 (O_2457,N_27590,N_28398);
xnor UO_2458 (O_2458,N_27076,N_29605);
and UO_2459 (O_2459,N_29094,N_28816);
and UO_2460 (O_2460,N_29755,N_28180);
or UO_2461 (O_2461,N_29064,N_27991);
or UO_2462 (O_2462,N_28365,N_27572);
and UO_2463 (O_2463,N_29385,N_28119);
and UO_2464 (O_2464,N_28207,N_27491);
xor UO_2465 (O_2465,N_27857,N_27267);
nor UO_2466 (O_2466,N_29683,N_29716);
nor UO_2467 (O_2467,N_29766,N_27809);
xnor UO_2468 (O_2468,N_28785,N_29200);
or UO_2469 (O_2469,N_27169,N_28324);
nand UO_2470 (O_2470,N_28657,N_27090);
and UO_2471 (O_2471,N_28409,N_29367);
and UO_2472 (O_2472,N_29445,N_28901);
and UO_2473 (O_2473,N_29764,N_27423);
nor UO_2474 (O_2474,N_29179,N_28389);
nand UO_2475 (O_2475,N_27401,N_29146);
and UO_2476 (O_2476,N_29860,N_28880);
xnor UO_2477 (O_2477,N_27535,N_27772);
xnor UO_2478 (O_2478,N_29224,N_29287);
or UO_2479 (O_2479,N_28344,N_28449);
nor UO_2480 (O_2480,N_27701,N_28703);
and UO_2481 (O_2481,N_27488,N_28924);
or UO_2482 (O_2482,N_28995,N_27298);
xor UO_2483 (O_2483,N_28384,N_27552);
or UO_2484 (O_2484,N_29966,N_27683);
or UO_2485 (O_2485,N_27067,N_29285);
or UO_2486 (O_2486,N_28790,N_27571);
nor UO_2487 (O_2487,N_29080,N_28983);
or UO_2488 (O_2488,N_29131,N_29489);
and UO_2489 (O_2489,N_27485,N_29315);
xor UO_2490 (O_2490,N_29035,N_28811);
nand UO_2491 (O_2491,N_28282,N_29017);
nand UO_2492 (O_2492,N_28075,N_27239);
xor UO_2493 (O_2493,N_27057,N_28202);
nand UO_2494 (O_2494,N_29913,N_28519);
or UO_2495 (O_2495,N_28132,N_29062);
and UO_2496 (O_2496,N_28675,N_29315);
nor UO_2497 (O_2497,N_28548,N_28242);
nand UO_2498 (O_2498,N_27525,N_27677);
nor UO_2499 (O_2499,N_27260,N_28007);
and UO_2500 (O_2500,N_27250,N_29477);
or UO_2501 (O_2501,N_27481,N_28615);
nand UO_2502 (O_2502,N_28203,N_28188);
or UO_2503 (O_2503,N_29360,N_28809);
or UO_2504 (O_2504,N_29826,N_27058);
or UO_2505 (O_2505,N_28355,N_29417);
or UO_2506 (O_2506,N_28874,N_28278);
and UO_2507 (O_2507,N_29941,N_27972);
nor UO_2508 (O_2508,N_29566,N_29379);
nand UO_2509 (O_2509,N_28921,N_29303);
xnor UO_2510 (O_2510,N_29445,N_27059);
or UO_2511 (O_2511,N_29041,N_27225);
nand UO_2512 (O_2512,N_27705,N_27797);
nand UO_2513 (O_2513,N_29265,N_28926);
or UO_2514 (O_2514,N_28179,N_27809);
and UO_2515 (O_2515,N_28308,N_28047);
nand UO_2516 (O_2516,N_29998,N_29155);
nand UO_2517 (O_2517,N_29939,N_27132);
nor UO_2518 (O_2518,N_29811,N_28293);
xor UO_2519 (O_2519,N_27219,N_29084);
nand UO_2520 (O_2520,N_28225,N_27510);
and UO_2521 (O_2521,N_29608,N_29000);
or UO_2522 (O_2522,N_28996,N_29765);
xor UO_2523 (O_2523,N_27952,N_28066);
and UO_2524 (O_2524,N_27976,N_27387);
or UO_2525 (O_2525,N_29634,N_27013);
or UO_2526 (O_2526,N_27281,N_27993);
xor UO_2527 (O_2527,N_27546,N_27504);
nor UO_2528 (O_2528,N_29745,N_29187);
nor UO_2529 (O_2529,N_29693,N_28379);
or UO_2530 (O_2530,N_29644,N_27123);
and UO_2531 (O_2531,N_27747,N_28324);
xnor UO_2532 (O_2532,N_28696,N_29055);
and UO_2533 (O_2533,N_29543,N_27865);
and UO_2534 (O_2534,N_28187,N_27977);
xnor UO_2535 (O_2535,N_27075,N_27225);
nand UO_2536 (O_2536,N_28082,N_27999);
or UO_2537 (O_2537,N_29919,N_29971);
nand UO_2538 (O_2538,N_27586,N_28405);
and UO_2539 (O_2539,N_27251,N_28881);
xor UO_2540 (O_2540,N_27774,N_29229);
nand UO_2541 (O_2541,N_27319,N_29256);
or UO_2542 (O_2542,N_29268,N_27808);
and UO_2543 (O_2543,N_27320,N_28437);
or UO_2544 (O_2544,N_29187,N_29039);
or UO_2545 (O_2545,N_28178,N_27763);
nand UO_2546 (O_2546,N_28988,N_29073);
nor UO_2547 (O_2547,N_27794,N_29985);
nor UO_2548 (O_2548,N_27480,N_27196);
and UO_2549 (O_2549,N_27042,N_28117);
nor UO_2550 (O_2550,N_29165,N_27431);
xor UO_2551 (O_2551,N_28741,N_28059);
nor UO_2552 (O_2552,N_27670,N_28072);
nand UO_2553 (O_2553,N_27886,N_27566);
nand UO_2554 (O_2554,N_27652,N_28223);
and UO_2555 (O_2555,N_28174,N_27803);
nand UO_2556 (O_2556,N_28362,N_27817);
xnor UO_2557 (O_2557,N_27296,N_27983);
xnor UO_2558 (O_2558,N_29082,N_29488);
nand UO_2559 (O_2559,N_29189,N_29222);
xnor UO_2560 (O_2560,N_28841,N_29141);
xnor UO_2561 (O_2561,N_28448,N_28088);
nor UO_2562 (O_2562,N_28934,N_27273);
or UO_2563 (O_2563,N_29208,N_27046);
and UO_2564 (O_2564,N_29176,N_28849);
or UO_2565 (O_2565,N_29117,N_27797);
nor UO_2566 (O_2566,N_27350,N_29539);
nor UO_2567 (O_2567,N_27826,N_28393);
xor UO_2568 (O_2568,N_28462,N_28563);
nand UO_2569 (O_2569,N_28005,N_29824);
xor UO_2570 (O_2570,N_27904,N_27502);
xor UO_2571 (O_2571,N_28393,N_29803);
xor UO_2572 (O_2572,N_28609,N_29043);
nand UO_2573 (O_2573,N_29500,N_27449);
nand UO_2574 (O_2574,N_27985,N_28571);
or UO_2575 (O_2575,N_27851,N_27729);
xnor UO_2576 (O_2576,N_28923,N_27467);
and UO_2577 (O_2577,N_29847,N_29049);
nand UO_2578 (O_2578,N_28665,N_28621);
or UO_2579 (O_2579,N_27677,N_29105);
and UO_2580 (O_2580,N_27348,N_28863);
xor UO_2581 (O_2581,N_27385,N_27775);
nor UO_2582 (O_2582,N_29544,N_29942);
or UO_2583 (O_2583,N_28131,N_29739);
xor UO_2584 (O_2584,N_28287,N_27349);
nor UO_2585 (O_2585,N_27153,N_29819);
nor UO_2586 (O_2586,N_29616,N_27514);
xnor UO_2587 (O_2587,N_28600,N_29876);
and UO_2588 (O_2588,N_28239,N_28485);
nand UO_2589 (O_2589,N_29381,N_28665);
nand UO_2590 (O_2590,N_29562,N_27552);
or UO_2591 (O_2591,N_27071,N_28754);
nor UO_2592 (O_2592,N_27107,N_27841);
xnor UO_2593 (O_2593,N_29822,N_29334);
nand UO_2594 (O_2594,N_28225,N_29565);
and UO_2595 (O_2595,N_28659,N_27899);
and UO_2596 (O_2596,N_27712,N_28863);
and UO_2597 (O_2597,N_28554,N_28383);
nor UO_2598 (O_2598,N_28736,N_27417);
or UO_2599 (O_2599,N_28236,N_27149);
nor UO_2600 (O_2600,N_29262,N_27587);
xnor UO_2601 (O_2601,N_27976,N_29809);
or UO_2602 (O_2602,N_27984,N_29750);
nor UO_2603 (O_2603,N_29824,N_29108);
xor UO_2604 (O_2604,N_29038,N_27593);
xnor UO_2605 (O_2605,N_28905,N_28363);
nor UO_2606 (O_2606,N_28695,N_27721);
xnor UO_2607 (O_2607,N_28531,N_28877);
nor UO_2608 (O_2608,N_28418,N_29421);
and UO_2609 (O_2609,N_27913,N_28289);
nor UO_2610 (O_2610,N_29201,N_29216);
or UO_2611 (O_2611,N_27966,N_28497);
or UO_2612 (O_2612,N_27895,N_27562);
nor UO_2613 (O_2613,N_29203,N_27238);
or UO_2614 (O_2614,N_29125,N_28561);
nand UO_2615 (O_2615,N_29786,N_29077);
nand UO_2616 (O_2616,N_29219,N_29227);
nor UO_2617 (O_2617,N_27050,N_28534);
and UO_2618 (O_2618,N_28361,N_27098);
xnor UO_2619 (O_2619,N_27780,N_28941);
xor UO_2620 (O_2620,N_28960,N_29821);
nor UO_2621 (O_2621,N_28366,N_29105);
xnor UO_2622 (O_2622,N_28323,N_29277);
or UO_2623 (O_2623,N_27422,N_27832);
xor UO_2624 (O_2624,N_28758,N_27169);
nor UO_2625 (O_2625,N_27434,N_27010);
nor UO_2626 (O_2626,N_28862,N_29664);
or UO_2627 (O_2627,N_27473,N_28454);
nand UO_2628 (O_2628,N_27806,N_29395);
nor UO_2629 (O_2629,N_27269,N_27717);
or UO_2630 (O_2630,N_28517,N_29389);
xor UO_2631 (O_2631,N_27451,N_29797);
nand UO_2632 (O_2632,N_27509,N_28366);
or UO_2633 (O_2633,N_29549,N_28138);
xnor UO_2634 (O_2634,N_29167,N_28108);
xnor UO_2635 (O_2635,N_29713,N_27582);
nor UO_2636 (O_2636,N_27178,N_29990);
or UO_2637 (O_2637,N_27150,N_29198);
nand UO_2638 (O_2638,N_29369,N_29348);
or UO_2639 (O_2639,N_29466,N_27907);
and UO_2640 (O_2640,N_29198,N_27383);
nor UO_2641 (O_2641,N_28816,N_27816);
or UO_2642 (O_2642,N_27994,N_29188);
and UO_2643 (O_2643,N_29705,N_28879);
nor UO_2644 (O_2644,N_28375,N_29466);
xnor UO_2645 (O_2645,N_27865,N_29245);
nand UO_2646 (O_2646,N_29618,N_29516);
xnor UO_2647 (O_2647,N_29725,N_28648);
nor UO_2648 (O_2648,N_28007,N_29108);
nand UO_2649 (O_2649,N_29581,N_28092);
and UO_2650 (O_2650,N_28547,N_29932);
xnor UO_2651 (O_2651,N_29444,N_27638);
nand UO_2652 (O_2652,N_27844,N_29177);
or UO_2653 (O_2653,N_27355,N_28528);
nand UO_2654 (O_2654,N_28300,N_28291);
and UO_2655 (O_2655,N_28032,N_27615);
and UO_2656 (O_2656,N_29491,N_28715);
or UO_2657 (O_2657,N_27171,N_27258);
xnor UO_2658 (O_2658,N_29147,N_28267);
xnor UO_2659 (O_2659,N_29219,N_29453);
nor UO_2660 (O_2660,N_27978,N_28501);
and UO_2661 (O_2661,N_27092,N_29614);
nand UO_2662 (O_2662,N_28737,N_27612);
nor UO_2663 (O_2663,N_27888,N_27666);
nor UO_2664 (O_2664,N_28134,N_27410);
or UO_2665 (O_2665,N_29347,N_27993);
and UO_2666 (O_2666,N_28504,N_27418);
or UO_2667 (O_2667,N_27047,N_27642);
nor UO_2668 (O_2668,N_27772,N_28699);
and UO_2669 (O_2669,N_29545,N_28581);
xnor UO_2670 (O_2670,N_27621,N_29552);
or UO_2671 (O_2671,N_29647,N_29402);
and UO_2672 (O_2672,N_28598,N_27433);
nand UO_2673 (O_2673,N_27562,N_29978);
or UO_2674 (O_2674,N_28865,N_27840);
nand UO_2675 (O_2675,N_29815,N_27626);
xnor UO_2676 (O_2676,N_28169,N_29076);
nand UO_2677 (O_2677,N_28216,N_27478);
and UO_2678 (O_2678,N_27733,N_29256);
xor UO_2679 (O_2679,N_27228,N_29857);
and UO_2680 (O_2680,N_29245,N_29003);
nand UO_2681 (O_2681,N_29496,N_29881);
and UO_2682 (O_2682,N_28889,N_29492);
nor UO_2683 (O_2683,N_29012,N_29948);
and UO_2684 (O_2684,N_28170,N_27002);
nor UO_2685 (O_2685,N_27456,N_28226);
xnor UO_2686 (O_2686,N_28577,N_27675);
nand UO_2687 (O_2687,N_29458,N_29907);
xor UO_2688 (O_2688,N_27689,N_28303);
nor UO_2689 (O_2689,N_27694,N_27454);
or UO_2690 (O_2690,N_29526,N_29327);
or UO_2691 (O_2691,N_29529,N_28989);
nand UO_2692 (O_2692,N_29479,N_27229);
nor UO_2693 (O_2693,N_29610,N_29031);
nand UO_2694 (O_2694,N_27964,N_27338);
or UO_2695 (O_2695,N_27835,N_28109);
xor UO_2696 (O_2696,N_28621,N_29629);
nor UO_2697 (O_2697,N_29511,N_29302);
xnor UO_2698 (O_2698,N_28370,N_27383);
or UO_2699 (O_2699,N_29380,N_29905);
nand UO_2700 (O_2700,N_28751,N_28102);
or UO_2701 (O_2701,N_28368,N_28245);
xnor UO_2702 (O_2702,N_28659,N_29053);
or UO_2703 (O_2703,N_28117,N_28887);
nand UO_2704 (O_2704,N_27931,N_29782);
xnor UO_2705 (O_2705,N_27923,N_28949);
xor UO_2706 (O_2706,N_29732,N_27523);
and UO_2707 (O_2707,N_29293,N_28247);
xor UO_2708 (O_2708,N_28945,N_28222);
and UO_2709 (O_2709,N_29794,N_27805);
xnor UO_2710 (O_2710,N_27135,N_29059);
xor UO_2711 (O_2711,N_29183,N_28998);
or UO_2712 (O_2712,N_29492,N_29259);
nand UO_2713 (O_2713,N_29801,N_28284);
nand UO_2714 (O_2714,N_28261,N_28085);
xnor UO_2715 (O_2715,N_29047,N_27783);
and UO_2716 (O_2716,N_29600,N_27995);
or UO_2717 (O_2717,N_28865,N_27152);
xor UO_2718 (O_2718,N_29510,N_27490);
xnor UO_2719 (O_2719,N_28741,N_27624);
and UO_2720 (O_2720,N_27349,N_27981);
nand UO_2721 (O_2721,N_28158,N_29485);
nand UO_2722 (O_2722,N_28119,N_28962);
nand UO_2723 (O_2723,N_28722,N_27058);
and UO_2724 (O_2724,N_29374,N_29132);
or UO_2725 (O_2725,N_28428,N_29767);
xnor UO_2726 (O_2726,N_28601,N_29947);
nand UO_2727 (O_2727,N_28037,N_28857);
and UO_2728 (O_2728,N_29561,N_27141);
nand UO_2729 (O_2729,N_27613,N_28599);
and UO_2730 (O_2730,N_27390,N_28493);
xor UO_2731 (O_2731,N_27133,N_28195);
and UO_2732 (O_2732,N_28849,N_28710);
or UO_2733 (O_2733,N_28371,N_29109);
or UO_2734 (O_2734,N_28029,N_28870);
or UO_2735 (O_2735,N_29246,N_27697);
xor UO_2736 (O_2736,N_27547,N_29454);
and UO_2737 (O_2737,N_27575,N_27728);
or UO_2738 (O_2738,N_28885,N_27663);
and UO_2739 (O_2739,N_29481,N_28560);
and UO_2740 (O_2740,N_28247,N_28244);
nand UO_2741 (O_2741,N_27203,N_28080);
xor UO_2742 (O_2742,N_28255,N_28485);
nand UO_2743 (O_2743,N_27874,N_27244);
and UO_2744 (O_2744,N_28287,N_29716);
xnor UO_2745 (O_2745,N_27664,N_29246);
and UO_2746 (O_2746,N_29262,N_28718);
and UO_2747 (O_2747,N_28849,N_28414);
xnor UO_2748 (O_2748,N_28926,N_28585);
and UO_2749 (O_2749,N_28019,N_28939);
and UO_2750 (O_2750,N_27895,N_29429);
xnor UO_2751 (O_2751,N_28956,N_29518);
and UO_2752 (O_2752,N_27183,N_28350);
xnor UO_2753 (O_2753,N_27364,N_28203);
xnor UO_2754 (O_2754,N_27067,N_28479);
or UO_2755 (O_2755,N_29200,N_29848);
nand UO_2756 (O_2756,N_28368,N_28803);
and UO_2757 (O_2757,N_27096,N_27005);
nor UO_2758 (O_2758,N_28243,N_27902);
or UO_2759 (O_2759,N_28681,N_29261);
nor UO_2760 (O_2760,N_29370,N_29273);
nor UO_2761 (O_2761,N_28321,N_29178);
or UO_2762 (O_2762,N_28572,N_28194);
nor UO_2763 (O_2763,N_29646,N_27948);
nand UO_2764 (O_2764,N_27389,N_28089);
nand UO_2765 (O_2765,N_29999,N_28844);
and UO_2766 (O_2766,N_27150,N_27655);
nor UO_2767 (O_2767,N_29098,N_29904);
nand UO_2768 (O_2768,N_27795,N_27218);
xor UO_2769 (O_2769,N_28813,N_29386);
xor UO_2770 (O_2770,N_27427,N_28464);
or UO_2771 (O_2771,N_27375,N_29480);
nor UO_2772 (O_2772,N_28738,N_29503);
nor UO_2773 (O_2773,N_28361,N_29860);
or UO_2774 (O_2774,N_27306,N_27694);
or UO_2775 (O_2775,N_27008,N_27373);
or UO_2776 (O_2776,N_29929,N_28486);
and UO_2777 (O_2777,N_27190,N_29367);
nor UO_2778 (O_2778,N_27330,N_27629);
nor UO_2779 (O_2779,N_29429,N_28019);
nand UO_2780 (O_2780,N_29008,N_28771);
nor UO_2781 (O_2781,N_28867,N_27881);
xnor UO_2782 (O_2782,N_29571,N_28716);
nor UO_2783 (O_2783,N_27529,N_29597);
nand UO_2784 (O_2784,N_28593,N_29462);
and UO_2785 (O_2785,N_27461,N_28338);
or UO_2786 (O_2786,N_28693,N_29891);
xor UO_2787 (O_2787,N_27474,N_29565);
xnor UO_2788 (O_2788,N_27320,N_29337);
nand UO_2789 (O_2789,N_27725,N_28075);
or UO_2790 (O_2790,N_28439,N_28309);
xnor UO_2791 (O_2791,N_28770,N_27929);
xnor UO_2792 (O_2792,N_27581,N_28559);
and UO_2793 (O_2793,N_27861,N_29039);
or UO_2794 (O_2794,N_29749,N_27442);
xor UO_2795 (O_2795,N_29949,N_28434);
or UO_2796 (O_2796,N_27750,N_27196);
nand UO_2797 (O_2797,N_27490,N_29242);
xor UO_2798 (O_2798,N_29043,N_28846);
nor UO_2799 (O_2799,N_28561,N_29749);
xnor UO_2800 (O_2800,N_28056,N_28968);
nor UO_2801 (O_2801,N_29260,N_29841);
nor UO_2802 (O_2802,N_29290,N_29503);
nor UO_2803 (O_2803,N_27960,N_27122);
or UO_2804 (O_2804,N_29431,N_29089);
and UO_2805 (O_2805,N_27841,N_27766);
or UO_2806 (O_2806,N_28091,N_28167);
and UO_2807 (O_2807,N_27917,N_29629);
and UO_2808 (O_2808,N_28054,N_28366);
and UO_2809 (O_2809,N_29006,N_29454);
xnor UO_2810 (O_2810,N_28308,N_27640);
nand UO_2811 (O_2811,N_29231,N_28596);
or UO_2812 (O_2812,N_28790,N_28223);
nand UO_2813 (O_2813,N_29864,N_29793);
nand UO_2814 (O_2814,N_29201,N_29657);
and UO_2815 (O_2815,N_28171,N_29105);
nand UO_2816 (O_2816,N_27226,N_27644);
nor UO_2817 (O_2817,N_29280,N_29523);
and UO_2818 (O_2818,N_28450,N_28691);
or UO_2819 (O_2819,N_29852,N_29619);
or UO_2820 (O_2820,N_28207,N_27189);
nor UO_2821 (O_2821,N_29951,N_28826);
nor UO_2822 (O_2822,N_28846,N_28309);
and UO_2823 (O_2823,N_29506,N_27336);
nor UO_2824 (O_2824,N_27382,N_27029);
xnor UO_2825 (O_2825,N_29563,N_29717);
xnor UO_2826 (O_2826,N_29885,N_28892);
or UO_2827 (O_2827,N_29131,N_28809);
and UO_2828 (O_2828,N_29342,N_28917);
or UO_2829 (O_2829,N_29923,N_27042);
and UO_2830 (O_2830,N_28499,N_27902);
nor UO_2831 (O_2831,N_29771,N_28798);
or UO_2832 (O_2832,N_27753,N_29132);
nor UO_2833 (O_2833,N_29849,N_28531);
nor UO_2834 (O_2834,N_27719,N_28196);
or UO_2835 (O_2835,N_27932,N_29303);
and UO_2836 (O_2836,N_28985,N_28652);
nand UO_2837 (O_2837,N_27811,N_27753);
nor UO_2838 (O_2838,N_28213,N_29283);
xor UO_2839 (O_2839,N_27115,N_27092);
and UO_2840 (O_2840,N_28374,N_28589);
and UO_2841 (O_2841,N_29190,N_29579);
and UO_2842 (O_2842,N_27847,N_29619);
or UO_2843 (O_2843,N_28395,N_28225);
xnor UO_2844 (O_2844,N_27839,N_28651);
xor UO_2845 (O_2845,N_27934,N_29579);
nor UO_2846 (O_2846,N_28289,N_28535);
and UO_2847 (O_2847,N_28321,N_27360);
nand UO_2848 (O_2848,N_27334,N_29327);
or UO_2849 (O_2849,N_27355,N_27379);
or UO_2850 (O_2850,N_28234,N_27014);
or UO_2851 (O_2851,N_29727,N_28445);
nand UO_2852 (O_2852,N_28093,N_28856);
nand UO_2853 (O_2853,N_28805,N_28005);
or UO_2854 (O_2854,N_28731,N_29288);
and UO_2855 (O_2855,N_29017,N_28184);
xor UO_2856 (O_2856,N_28975,N_28289);
or UO_2857 (O_2857,N_28395,N_28137);
nor UO_2858 (O_2858,N_28976,N_29797);
xnor UO_2859 (O_2859,N_27140,N_29692);
nor UO_2860 (O_2860,N_28476,N_29252);
xnor UO_2861 (O_2861,N_29768,N_28574);
xnor UO_2862 (O_2862,N_28810,N_28237);
nor UO_2863 (O_2863,N_28030,N_27818);
nor UO_2864 (O_2864,N_28395,N_28975);
or UO_2865 (O_2865,N_28660,N_29621);
or UO_2866 (O_2866,N_27720,N_29804);
nand UO_2867 (O_2867,N_27505,N_29906);
nor UO_2868 (O_2868,N_27394,N_27719);
nor UO_2869 (O_2869,N_27360,N_29332);
or UO_2870 (O_2870,N_28969,N_28457);
nand UO_2871 (O_2871,N_27604,N_29341);
nor UO_2872 (O_2872,N_28773,N_29530);
nand UO_2873 (O_2873,N_29503,N_27770);
nor UO_2874 (O_2874,N_27849,N_28649);
or UO_2875 (O_2875,N_27687,N_29944);
nor UO_2876 (O_2876,N_28783,N_28493);
and UO_2877 (O_2877,N_29474,N_29277);
or UO_2878 (O_2878,N_29685,N_28154);
nor UO_2879 (O_2879,N_28786,N_28696);
and UO_2880 (O_2880,N_27084,N_29537);
or UO_2881 (O_2881,N_27253,N_28717);
or UO_2882 (O_2882,N_28934,N_27758);
or UO_2883 (O_2883,N_27899,N_29371);
or UO_2884 (O_2884,N_28204,N_29220);
nand UO_2885 (O_2885,N_28500,N_28178);
or UO_2886 (O_2886,N_28319,N_27246);
xnor UO_2887 (O_2887,N_29697,N_28210);
and UO_2888 (O_2888,N_27390,N_28633);
xnor UO_2889 (O_2889,N_29067,N_28610);
xnor UO_2890 (O_2890,N_29284,N_29907);
xor UO_2891 (O_2891,N_29929,N_28831);
and UO_2892 (O_2892,N_29065,N_27447);
and UO_2893 (O_2893,N_27875,N_27906);
nor UO_2894 (O_2894,N_27797,N_28100);
or UO_2895 (O_2895,N_29705,N_27601);
or UO_2896 (O_2896,N_27865,N_29418);
nand UO_2897 (O_2897,N_29454,N_27822);
and UO_2898 (O_2898,N_27928,N_29528);
nor UO_2899 (O_2899,N_29859,N_28907);
or UO_2900 (O_2900,N_29050,N_28449);
or UO_2901 (O_2901,N_29263,N_28195);
nand UO_2902 (O_2902,N_28115,N_27799);
xnor UO_2903 (O_2903,N_29179,N_29150);
and UO_2904 (O_2904,N_27864,N_29062);
nand UO_2905 (O_2905,N_27954,N_29720);
nor UO_2906 (O_2906,N_28534,N_27325);
xnor UO_2907 (O_2907,N_28354,N_29792);
and UO_2908 (O_2908,N_27715,N_28284);
xnor UO_2909 (O_2909,N_28964,N_28642);
nor UO_2910 (O_2910,N_28135,N_28476);
nand UO_2911 (O_2911,N_28333,N_29929);
nand UO_2912 (O_2912,N_29932,N_28077);
nand UO_2913 (O_2913,N_29951,N_27662);
or UO_2914 (O_2914,N_28355,N_29662);
nand UO_2915 (O_2915,N_29281,N_29182);
and UO_2916 (O_2916,N_28147,N_28497);
nor UO_2917 (O_2917,N_28432,N_27741);
nand UO_2918 (O_2918,N_29283,N_29758);
xnor UO_2919 (O_2919,N_29694,N_27446);
nor UO_2920 (O_2920,N_28494,N_28830);
nor UO_2921 (O_2921,N_27157,N_29452);
nand UO_2922 (O_2922,N_29591,N_29709);
or UO_2923 (O_2923,N_28470,N_28519);
nand UO_2924 (O_2924,N_27715,N_29057);
and UO_2925 (O_2925,N_28580,N_27115);
or UO_2926 (O_2926,N_29842,N_27240);
nor UO_2927 (O_2927,N_29207,N_27422);
nand UO_2928 (O_2928,N_28432,N_28472);
nor UO_2929 (O_2929,N_29308,N_29591);
xor UO_2930 (O_2930,N_29387,N_27360);
or UO_2931 (O_2931,N_28923,N_27992);
or UO_2932 (O_2932,N_29092,N_27769);
nor UO_2933 (O_2933,N_29258,N_27780);
or UO_2934 (O_2934,N_29006,N_27364);
and UO_2935 (O_2935,N_29209,N_29121);
or UO_2936 (O_2936,N_28616,N_27270);
xor UO_2937 (O_2937,N_28698,N_27499);
nand UO_2938 (O_2938,N_28673,N_29606);
xnor UO_2939 (O_2939,N_28702,N_28651);
and UO_2940 (O_2940,N_28649,N_28377);
and UO_2941 (O_2941,N_28977,N_29453);
xor UO_2942 (O_2942,N_29643,N_28867);
xor UO_2943 (O_2943,N_27196,N_29268);
nor UO_2944 (O_2944,N_29192,N_29261);
or UO_2945 (O_2945,N_29907,N_28159);
xnor UO_2946 (O_2946,N_27579,N_28958);
nor UO_2947 (O_2947,N_29343,N_29302);
nand UO_2948 (O_2948,N_29938,N_28398);
or UO_2949 (O_2949,N_27970,N_27328);
xnor UO_2950 (O_2950,N_27328,N_29577);
nor UO_2951 (O_2951,N_27309,N_29112);
or UO_2952 (O_2952,N_27300,N_28384);
xor UO_2953 (O_2953,N_29153,N_28200);
xor UO_2954 (O_2954,N_29767,N_28873);
nor UO_2955 (O_2955,N_28583,N_28142);
xnor UO_2956 (O_2956,N_28630,N_29203);
or UO_2957 (O_2957,N_27177,N_28042);
or UO_2958 (O_2958,N_28096,N_29445);
nand UO_2959 (O_2959,N_27852,N_29109);
nand UO_2960 (O_2960,N_28073,N_27076);
nand UO_2961 (O_2961,N_29313,N_28800);
nand UO_2962 (O_2962,N_27689,N_27686);
xor UO_2963 (O_2963,N_27174,N_28493);
or UO_2964 (O_2964,N_29531,N_28769);
and UO_2965 (O_2965,N_27462,N_28583);
nand UO_2966 (O_2966,N_28278,N_28758);
xnor UO_2967 (O_2967,N_29363,N_28901);
nand UO_2968 (O_2968,N_28973,N_29699);
nand UO_2969 (O_2969,N_28549,N_29373);
nor UO_2970 (O_2970,N_28602,N_28251);
and UO_2971 (O_2971,N_28588,N_28652);
nor UO_2972 (O_2972,N_27326,N_28710);
and UO_2973 (O_2973,N_27824,N_28650);
or UO_2974 (O_2974,N_27664,N_28853);
xnor UO_2975 (O_2975,N_29405,N_28462);
nor UO_2976 (O_2976,N_29376,N_29176);
nor UO_2977 (O_2977,N_28382,N_27470);
or UO_2978 (O_2978,N_27908,N_28151);
nor UO_2979 (O_2979,N_27878,N_27318);
nor UO_2980 (O_2980,N_28901,N_27746);
nand UO_2981 (O_2981,N_27852,N_29200);
xnor UO_2982 (O_2982,N_27114,N_29368);
or UO_2983 (O_2983,N_27415,N_29186);
nand UO_2984 (O_2984,N_29565,N_29578);
xor UO_2985 (O_2985,N_28475,N_29369);
nor UO_2986 (O_2986,N_28247,N_27072);
nor UO_2987 (O_2987,N_29222,N_28691);
or UO_2988 (O_2988,N_29180,N_27156);
or UO_2989 (O_2989,N_28965,N_29244);
xor UO_2990 (O_2990,N_28914,N_29807);
nand UO_2991 (O_2991,N_28550,N_29703);
nor UO_2992 (O_2992,N_27450,N_29340);
or UO_2993 (O_2993,N_28713,N_29949);
nand UO_2994 (O_2994,N_29907,N_28697);
nand UO_2995 (O_2995,N_29459,N_28695);
nor UO_2996 (O_2996,N_27303,N_27711);
nand UO_2997 (O_2997,N_29986,N_27064);
nor UO_2998 (O_2998,N_27732,N_28406);
or UO_2999 (O_2999,N_27468,N_27828);
nand UO_3000 (O_3000,N_28459,N_28209);
and UO_3001 (O_3001,N_27040,N_29717);
and UO_3002 (O_3002,N_29335,N_27166);
xor UO_3003 (O_3003,N_29680,N_29974);
and UO_3004 (O_3004,N_29431,N_28394);
and UO_3005 (O_3005,N_27952,N_28673);
or UO_3006 (O_3006,N_28482,N_27621);
xnor UO_3007 (O_3007,N_27782,N_29008);
xnor UO_3008 (O_3008,N_27720,N_29831);
nor UO_3009 (O_3009,N_27989,N_29747);
nor UO_3010 (O_3010,N_28205,N_29716);
nor UO_3011 (O_3011,N_29031,N_29660);
and UO_3012 (O_3012,N_28839,N_27731);
nand UO_3013 (O_3013,N_27994,N_29735);
xor UO_3014 (O_3014,N_28175,N_27092);
and UO_3015 (O_3015,N_29950,N_28835);
nor UO_3016 (O_3016,N_28424,N_27825);
nand UO_3017 (O_3017,N_27856,N_27158);
nor UO_3018 (O_3018,N_27818,N_28685);
nor UO_3019 (O_3019,N_29571,N_29994);
xnor UO_3020 (O_3020,N_27050,N_27757);
nor UO_3021 (O_3021,N_29620,N_27992);
nor UO_3022 (O_3022,N_27911,N_29346);
xor UO_3023 (O_3023,N_27609,N_28652);
and UO_3024 (O_3024,N_28715,N_27812);
nand UO_3025 (O_3025,N_29696,N_28100);
and UO_3026 (O_3026,N_28996,N_27912);
and UO_3027 (O_3027,N_29193,N_29810);
xnor UO_3028 (O_3028,N_28455,N_27169);
or UO_3029 (O_3029,N_29589,N_28621);
nand UO_3030 (O_3030,N_28123,N_29057);
xnor UO_3031 (O_3031,N_27104,N_29159);
nor UO_3032 (O_3032,N_29964,N_28214);
or UO_3033 (O_3033,N_28633,N_27656);
xor UO_3034 (O_3034,N_28210,N_27458);
xor UO_3035 (O_3035,N_28941,N_27142);
or UO_3036 (O_3036,N_27926,N_27611);
and UO_3037 (O_3037,N_28406,N_28814);
nand UO_3038 (O_3038,N_27933,N_29225);
nor UO_3039 (O_3039,N_27479,N_27159);
xnor UO_3040 (O_3040,N_29603,N_29451);
nand UO_3041 (O_3041,N_29259,N_27509);
or UO_3042 (O_3042,N_29782,N_28003);
nor UO_3043 (O_3043,N_29481,N_27401);
nor UO_3044 (O_3044,N_29496,N_29395);
and UO_3045 (O_3045,N_28407,N_28447);
nand UO_3046 (O_3046,N_29182,N_29981);
nor UO_3047 (O_3047,N_29620,N_28785);
nand UO_3048 (O_3048,N_28652,N_28439);
nand UO_3049 (O_3049,N_29443,N_27073);
and UO_3050 (O_3050,N_28353,N_29898);
and UO_3051 (O_3051,N_28684,N_27100);
and UO_3052 (O_3052,N_29413,N_28339);
or UO_3053 (O_3053,N_28902,N_29068);
xnor UO_3054 (O_3054,N_29635,N_29590);
nand UO_3055 (O_3055,N_28096,N_27493);
nand UO_3056 (O_3056,N_27572,N_28937);
nor UO_3057 (O_3057,N_28863,N_29148);
nor UO_3058 (O_3058,N_27709,N_27617);
xor UO_3059 (O_3059,N_28878,N_29147);
xor UO_3060 (O_3060,N_28415,N_29299);
or UO_3061 (O_3061,N_28478,N_29575);
xnor UO_3062 (O_3062,N_27827,N_27473);
and UO_3063 (O_3063,N_28301,N_27114);
nand UO_3064 (O_3064,N_27508,N_27002);
xor UO_3065 (O_3065,N_29060,N_28421);
xor UO_3066 (O_3066,N_27163,N_27981);
or UO_3067 (O_3067,N_28693,N_29417);
and UO_3068 (O_3068,N_27900,N_27339);
nor UO_3069 (O_3069,N_28821,N_29919);
nor UO_3070 (O_3070,N_28896,N_28363);
or UO_3071 (O_3071,N_29506,N_28180);
nor UO_3072 (O_3072,N_28946,N_28319);
and UO_3073 (O_3073,N_29025,N_27224);
and UO_3074 (O_3074,N_29957,N_29489);
or UO_3075 (O_3075,N_29526,N_27093);
nand UO_3076 (O_3076,N_28954,N_29658);
or UO_3077 (O_3077,N_29198,N_28232);
nor UO_3078 (O_3078,N_29291,N_29013);
or UO_3079 (O_3079,N_27699,N_27280);
nand UO_3080 (O_3080,N_29618,N_28677);
nand UO_3081 (O_3081,N_29872,N_29130);
or UO_3082 (O_3082,N_28414,N_27072);
and UO_3083 (O_3083,N_27890,N_28589);
or UO_3084 (O_3084,N_28065,N_27408);
nor UO_3085 (O_3085,N_27935,N_27886);
or UO_3086 (O_3086,N_27094,N_29096);
and UO_3087 (O_3087,N_28999,N_28748);
or UO_3088 (O_3088,N_29370,N_28897);
and UO_3089 (O_3089,N_27826,N_27969);
nand UO_3090 (O_3090,N_27729,N_28733);
and UO_3091 (O_3091,N_28779,N_29019);
xnor UO_3092 (O_3092,N_28797,N_29231);
nor UO_3093 (O_3093,N_28227,N_28509);
nand UO_3094 (O_3094,N_29726,N_29998);
or UO_3095 (O_3095,N_29382,N_28770);
or UO_3096 (O_3096,N_28577,N_27227);
nor UO_3097 (O_3097,N_29170,N_27464);
xnor UO_3098 (O_3098,N_27581,N_29130);
nor UO_3099 (O_3099,N_29378,N_27596);
nand UO_3100 (O_3100,N_28888,N_29118);
and UO_3101 (O_3101,N_29397,N_29070);
nor UO_3102 (O_3102,N_29895,N_29376);
and UO_3103 (O_3103,N_28451,N_29596);
nor UO_3104 (O_3104,N_29407,N_28809);
xnor UO_3105 (O_3105,N_28598,N_28976);
and UO_3106 (O_3106,N_28461,N_29083);
nand UO_3107 (O_3107,N_27587,N_27311);
or UO_3108 (O_3108,N_29533,N_29393);
xnor UO_3109 (O_3109,N_28370,N_27367);
and UO_3110 (O_3110,N_27348,N_29195);
nand UO_3111 (O_3111,N_29657,N_27541);
nor UO_3112 (O_3112,N_29132,N_27957);
nand UO_3113 (O_3113,N_27498,N_29064);
or UO_3114 (O_3114,N_27302,N_29253);
and UO_3115 (O_3115,N_28167,N_27704);
or UO_3116 (O_3116,N_27427,N_28342);
or UO_3117 (O_3117,N_27541,N_28649);
xor UO_3118 (O_3118,N_27434,N_27528);
nand UO_3119 (O_3119,N_29862,N_29812);
nor UO_3120 (O_3120,N_28991,N_27824);
and UO_3121 (O_3121,N_27797,N_28010);
or UO_3122 (O_3122,N_27593,N_27633);
nor UO_3123 (O_3123,N_29656,N_29960);
nand UO_3124 (O_3124,N_27469,N_29833);
nor UO_3125 (O_3125,N_28560,N_28729);
or UO_3126 (O_3126,N_29686,N_29534);
and UO_3127 (O_3127,N_29731,N_27062);
nand UO_3128 (O_3128,N_27886,N_28633);
or UO_3129 (O_3129,N_28863,N_29445);
or UO_3130 (O_3130,N_29060,N_27809);
nor UO_3131 (O_3131,N_29616,N_29834);
nand UO_3132 (O_3132,N_29796,N_28100);
and UO_3133 (O_3133,N_27692,N_29459);
xor UO_3134 (O_3134,N_29906,N_28802);
nand UO_3135 (O_3135,N_27329,N_28814);
nand UO_3136 (O_3136,N_29802,N_29798);
and UO_3137 (O_3137,N_29811,N_28188);
nand UO_3138 (O_3138,N_27348,N_28889);
or UO_3139 (O_3139,N_29085,N_27705);
xnor UO_3140 (O_3140,N_27670,N_28640);
nor UO_3141 (O_3141,N_28538,N_29357);
nand UO_3142 (O_3142,N_28052,N_27835);
nand UO_3143 (O_3143,N_29962,N_29662);
and UO_3144 (O_3144,N_28061,N_28072);
and UO_3145 (O_3145,N_29540,N_29545);
or UO_3146 (O_3146,N_27229,N_29444);
nor UO_3147 (O_3147,N_27950,N_29690);
nor UO_3148 (O_3148,N_29662,N_29037);
nand UO_3149 (O_3149,N_27776,N_28735);
and UO_3150 (O_3150,N_27683,N_29520);
nand UO_3151 (O_3151,N_27185,N_29619);
nor UO_3152 (O_3152,N_27244,N_29282);
or UO_3153 (O_3153,N_28727,N_29004);
and UO_3154 (O_3154,N_28686,N_28414);
or UO_3155 (O_3155,N_29090,N_27323);
or UO_3156 (O_3156,N_29672,N_29970);
nand UO_3157 (O_3157,N_29007,N_29000);
nand UO_3158 (O_3158,N_28029,N_29193);
nand UO_3159 (O_3159,N_28551,N_28108);
xor UO_3160 (O_3160,N_29769,N_27311);
and UO_3161 (O_3161,N_27252,N_27796);
nor UO_3162 (O_3162,N_27247,N_28579);
xnor UO_3163 (O_3163,N_28382,N_29406);
or UO_3164 (O_3164,N_29583,N_27992);
xnor UO_3165 (O_3165,N_29967,N_29795);
nor UO_3166 (O_3166,N_27605,N_28624);
nand UO_3167 (O_3167,N_27265,N_27490);
nor UO_3168 (O_3168,N_29126,N_28931);
and UO_3169 (O_3169,N_27824,N_27313);
and UO_3170 (O_3170,N_28619,N_27129);
nand UO_3171 (O_3171,N_28833,N_27997);
and UO_3172 (O_3172,N_27872,N_27221);
xor UO_3173 (O_3173,N_29857,N_28106);
or UO_3174 (O_3174,N_29033,N_29362);
and UO_3175 (O_3175,N_27998,N_29773);
nand UO_3176 (O_3176,N_28957,N_28784);
and UO_3177 (O_3177,N_29136,N_29782);
xor UO_3178 (O_3178,N_28169,N_27576);
and UO_3179 (O_3179,N_28817,N_29128);
nand UO_3180 (O_3180,N_28070,N_28118);
xnor UO_3181 (O_3181,N_27841,N_29817);
xor UO_3182 (O_3182,N_28132,N_29138);
xnor UO_3183 (O_3183,N_28729,N_28526);
nand UO_3184 (O_3184,N_29287,N_27252);
nor UO_3185 (O_3185,N_29620,N_27553);
xor UO_3186 (O_3186,N_27945,N_27044);
or UO_3187 (O_3187,N_29017,N_29633);
xor UO_3188 (O_3188,N_29314,N_27219);
nor UO_3189 (O_3189,N_27249,N_27453);
or UO_3190 (O_3190,N_27355,N_28377);
and UO_3191 (O_3191,N_27891,N_29298);
nor UO_3192 (O_3192,N_29512,N_28819);
nand UO_3193 (O_3193,N_29541,N_28602);
or UO_3194 (O_3194,N_28981,N_29956);
and UO_3195 (O_3195,N_28196,N_29697);
or UO_3196 (O_3196,N_27872,N_27875);
xor UO_3197 (O_3197,N_27974,N_29528);
nor UO_3198 (O_3198,N_29811,N_29156);
nand UO_3199 (O_3199,N_28194,N_28677);
xnor UO_3200 (O_3200,N_29347,N_28642);
and UO_3201 (O_3201,N_29467,N_29962);
nor UO_3202 (O_3202,N_28852,N_28668);
and UO_3203 (O_3203,N_28138,N_27243);
xor UO_3204 (O_3204,N_27945,N_28920);
and UO_3205 (O_3205,N_29494,N_28636);
nand UO_3206 (O_3206,N_29544,N_27527);
nor UO_3207 (O_3207,N_27122,N_28717);
nor UO_3208 (O_3208,N_29424,N_27918);
and UO_3209 (O_3209,N_28283,N_28008);
and UO_3210 (O_3210,N_29185,N_27014);
or UO_3211 (O_3211,N_28759,N_29118);
nor UO_3212 (O_3212,N_27020,N_28435);
or UO_3213 (O_3213,N_27899,N_27931);
nand UO_3214 (O_3214,N_27117,N_29995);
nand UO_3215 (O_3215,N_27765,N_28627);
and UO_3216 (O_3216,N_28152,N_27065);
or UO_3217 (O_3217,N_29439,N_29243);
nor UO_3218 (O_3218,N_28914,N_27943);
or UO_3219 (O_3219,N_28537,N_29821);
nand UO_3220 (O_3220,N_29049,N_29989);
and UO_3221 (O_3221,N_27011,N_27429);
nor UO_3222 (O_3222,N_29667,N_29899);
nand UO_3223 (O_3223,N_27345,N_29609);
or UO_3224 (O_3224,N_27448,N_29978);
nand UO_3225 (O_3225,N_27730,N_27368);
and UO_3226 (O_3226,N_28273,N_29543);
nand UO_3227 (O_3227,N_27121,N_29576);
xor UO_3228 (O_3228,N_27607,N_29101);
and UO_3229 (O_3229,N_27989,N_29578);
nand UO_3230 (O_3230,N_27891,N_28442);
or UO_3231 (O_3231,N_29233,N_28240);
nand UO_3232 (O_3232,N_27557,N_28631);
and UO_3233 (O_3233,N_28461,N_29067);
nand UO_3234 (O_3234,N_27152,N_29596);
nor UO_3235 (O_3235,N_28346,N_29203);
nand UO_3236 (O_3236,N_28520,N_27182);
or UO_3237 (O_3237,N_27293,N_28038);
nand UO_3238 (O_3238,N_29432,N_27377);
xor UO_3239 (O_3239,N_27852,N_29446);
nor UO_3240 (O_3240,N_28721,N_29249);
or UO_3241 (O_3241,N_29292,N_27805);
xnor UO_3242 (O_3242,N_29537,N_27218);
xor UO_3243 (O_3243,N_29309,N_29468);
nor UO_3244 (O_3244,N_27671,N_29814);
or UO_3245 (O_3245,N_27450,N_27076);
nand UO_3246 (O_3246,N_29809,N_28166);
nor UO_3247 (O_3247,N_27565,N_27684);
or UO_3248 (O_3248,N_28670,N_28022);
nor UO_3249 (O_3249,N_29202,N_28020);
nand UO_3250 (O_3250,N_28740,N_28842);
nand UO_3251 (O_3251,N_28478,N_28280);
or UO_3252 (O_3252,N_27051,N_29827);
or UO_3253 (O_3253,N_27377,N_27417);
xor UO_3254 (O_3254,N_27888,N_28278);
xnor UO_3255 (O_3255,N_28253,N_29405);
nor UO_3256 (O_3256,N_27455,N_28015);
and UO_3257 (O_3257,N_28059,N_27707);
nand UO_3258 (O_3258,N_29833,N_29473);
nor UO_3259 (O_3259,N_29398,N_29474);
or UO_3260 (O_3260,N_29646,N_27630);
nand UO_3261 (O_3261,N_28116,N_29622);
xnor UO_3262 (O_3262,N_29336,N_27198);
and UO_3263 (O_3263,N_28079,N_28532);
nor UO_3264 (O_3264,N_27175,N_27318);
and UO_3265 (O_3265,N_27790,N_27106);
nand UO_3266 (O_3266,N_27892,N_27038);
or UO_3267 (O_3267,N_28691,N_28096);
nor UO_3268 (O_3268,N_28472,N_27343);
or UO_3269 (O_3269,N_27819,N_27075);
nand UO_3270 (O_3270,N_27330,N_28427);
and UO_3271 (O_3271,N_27506,N_29155);
nand UO_3272 (O_3272,N_27550,N_27948);
nand UO_3273 (O_3273,N_28739,N_28790);
and UO_3274 (O_3274,N_29499,N_27167);
nand UO_3275 (O_3275,N_28598,N_29169);
xor UO_3276 (O_3276,N_27587,N_28942);
nor UO_3277 (O_3277,N_27836,N_27036);
xor UO_3278 (O_3278,N_27062,N_28030);
nor UO_3279 (O_3279,N_29252,N_28063);
xor UO_3280 (O_3280,N_28189,N_27801);
xnor UO_3281 (O_3281,N_29007,N_27461);
nor UO_3282 (O_3282,N_27344,N_28130);
xnor UO_3283 (O_3283,N_27849,N_27861);
nor UO_3284 (O_3284,N_27331,N_27544);
and UO_3285 (O_3285,N_29009,N_28629);
xor UO_3286 (O_3286,N_27761,N_28743);
nand UO_3287 (O_3287,N_29409,N_29646);
nand UO_3288 (O_3288,N_28683,N_27467);
nor UO_3289 (O_3289,N_29861,N_27909);
nand UO_3290 (O_3290,N_29807,N_29088);
or UO_3291 (O_3291,N_27419,N_29659);
nor UO_3292 (O_3292,N_28060,N_29477);
or UO_3293 (O_3293,N_29696,N_27086);
xnor UO_3294 (O_3294,N_27193,N_27550);
nor UO_3295 (O_3295,N_27385,N_28910);
nor UO_3296 (O_3296,N_29829,N_29784);
xnor UO_3297 (O_3297,N_29648,N_29542);
nand UO_3298 (O_3298,N_27467,N_27154);
nor UO_3299 (O_3299,N_27909,N_27604);
nand UO_3300 (O_3300,N_27411,N_29047);
nor UO_3301 (O_3301,N_27903,N_28744);
nor UO_3302 (O_3302,N_28332,N_29880);
or UO_3303 (O_3303,N_27581,N_29825);
nand UO_3304 (O_3304,N_29047,N_28908);
or UO_3305 (O_3305,N_28726,N_27104);
or UO_3306 (O_3306,N_28736,N_28051);
or UO_3307 (O_3307,N_27961,N_29075);
and UO_3308 (O_3308,N_29050,N_29733);
or UO_3309 (O_3309,N_29155,N_27383);
nor UO_3310 (O_3310,N_28358,N_28215);
nor UO_3311 (O_3311,N_29128,N_29464);
nand UO_3312 (O_3312,N_29375,N_29522);
and UO_3313 (O_3313,N_27178,N_29963);
xor UO_3314 (O_3314,N_28545,N_27243);
or UO_3315 (O_3315,N_27076,N_28851);
and UO_3316 (O_3316,N_27952,N_28029);
nand UO_3317 (O_3317,N_29679,N_29362);
nand UO_3318 (O_3318,N_29975,N_29377);
nor UO_3319 (O_3319,N_29880,N_27820);
or UO_3320 (O_3320,N_29558,N_28301);
or UO_3321 (O_3321,N_29164,N_29357);
nand UO_3322 (O_3322,N_28718,N_28281);
nand UO_3323 (O_3323,N_28608,N_28941);
xor UO_3324 (O_3324,N_29807,N_27968);
nor UO_3325 (O_3325,N_27114,N_28210);
and UO_3326 (O_3326,N_29917,N_28878);
nand UO_3327 (O_3327,N_29694,N_27961);
or UO_3328 (O_3328,N_28570,N_29977);
or UO_3329 (O_3329,N_27161,N_28360);
xor UO_3330 (O_3330,N_29854,N_28011);
nand UO_3331 (O_3331,N_29614,N_29867);
nand UO_3332 (O_3332,N_27447,N_28007);
or UO_3333 (O_3333,N_28354,N_27213);
or UO_3334 (O_3334,N_29012,N_28139);
nand UO_3335 (O_3335,N_28461,N_27103);
xnor UO_3336 (O_3336,N_27541,N_29272);
or UO_3337 (O_3337,N_28303,N_28675);
or UO_3338 (O_3338,N_27343,N_28323);
and UO_3339 (O_3339,N_29958,N_27918);
nand UO_3340 (O_3340,N_28751,N_29246);
nand UO_3341 (O_3341,N_29534,N_27879);
or UO_3342 (O_3342,N_28684,N_28789);
xor UO_3343 (O_3343,N_29555,N_28530);
and UO_3344 (O_3344,N_27542,N_27744);
and UO_3345 (O_3345,N_27109,N_29307);
and UO_3346 (O_3346,N_29498,N_29139);
xnor UO_3347 (O_3347,N_27805,N_27927);
nand UO_3348 (O_3348,N_29261,N_29668);
or UO_3349 (O_3349,N_27450,N_29111);
xor UO_3350 (O_3350,N_29105,N_28858);
and UO_3351 (O_3351,N_27567,N_27766);
xnor UO_3352 (O_3352,N_27353,N_27630);
nor UO_3353 (O_3353,N_29228,N_27883);
nor UO_3354 (O_3354,N_27692,N_29012);
nand UO_3355 (O_3355,N_27007,N_28645);
or UO_3356 (O_3356,N_29967,N_29379);
and UO_3357 (O_3357,N_27656,N_27621);
or UO_3358 (O_3358,N_28948,N_28451);
or UO_3359 (O_3359,N_28489,N_29899);
xnor UO_3360 (O_3360,N_29535,N_28670);
nor UO_3361 (O_3361,N_28760,N_28602);
nor UO_3362 (O_3362,N_28961,N_29179);
or UO_3363 (O_3363,N_27914,N_29957);
nand UO_3364 (O_3364,N_29467,N_29087);
or UO_3365 (O_3365,N_27636,N_28800);
or UO_3366 (O_3366,N_27857,N_29208);
nor UO_3367 (O_3367,N_28724,N_28635);
and UO_3368 (O_3368,N_27052,N_28995);
nor UO_3369 (O_3369,N_29518,N_29929);
nand UO_3370 (O_3370,N_27572,N_29093);
and UO_3371 (O_3371,N_28382,N_29919);
nor UO_3372 (O_3372,N_29771,N_29830);
or UO_3373 (O_3373,N_29274,N_29099);
or UO_3374 (O_3374,N_27997,N_28658);
or UO_3375 (O_3375,N_29293,N_28921);
nor UO_3376 (O_3376,N_27171,N_28014);
xnor UO_3377 (O_3377,N_28013,N_29798);
nor UO_3378 (O_3378,N_28404,N_28744);
xnor UO_3379 (O_3379,N_27947,N_27892);
and UO_3380 (O_3380,N_29183,N_28767);
and UO_3381 (O_3381,N_29659,N_29962);
nand UO_3382 (O_3382,N_28712,N_27002);
and UO_3383 (O_3383,N_27492,N_29389);
nand UO_3384 (O_3384,N_27426,N_29037);
xnor UO_3385 (O_3385,N_27043,N_28836);
and UO_3386 (O_3386,N_29604,N_29880);
nand UO_3387 (O_3387,N_27039,N_27032);
nor UO_3388 (O_3388,N_27446,N_28700);
and UO_3389 (O_3389,N_29647,N_27311);
nand UO_3390 (O_3390,N_27653,N_29117);
xnor UO_3391 (O_3391,N_29825,N_27459);
xor UO_3392 (O_3392,N_28739,N_28997);
and UO_3393 (O_3393,N_28095,N_29921);
and UO_3394 (O_3394,N_27474,N_29611);
and UO_3395 (O_3395,N_28369,N_27288);
xor UO_3396 (O_3396,N_28945,N_29792);
nor UO_3397 (O_3397,N_28143,N_27495);
xor UO_3398 (O_3398,N_27579,N_27426);
nor UO_3399 (O_3399,N_29459,N_29571);
nand UO_3400 (O_3400,N_29582,N_29628);
or UO_3401 (O_3401,N_29095,N_27442);
and UO_3402 (O_3402,N_28818,N_28986);
or UO_3403 (O_3403,N_29367,N_28355);
or UO_3404 (O_3404,N_29114,N_27122);
and UO_3405 (O_3405,N_29915,N_27271);
and UO_3406 (O_3406,N_27506,N_29392);
nor UO_3407 (O_3407,N_29465,N_28154);
nand UO_3408 (O_3408,N_27353,N_27254);
or UO_3409 (O_3409,N_28972,N_27969);
xnor UO_3410 (O_3410,N_29291,N_29817);
nand UO_3411 (O_3411,N_27090,N_27748);
and UO_3412 (O_3412,N_27678,N_28596);
and UO_3413 (O_3413,N_29375,N_27712);
nor UO_3414 (O_3414,N_28253,N_27378);
xnor UO_3415 (O_3415,N_29789,N_27923);
or UO_3416 (O_3416,N_28928,N_28441);
and UO_3417 (O_3417,N_27383,N_27403);
xnor UO_3418 (O_3418,N_27787,N_27943);
and UO_3419 (O_3419,N_27556,N_27040);
nand UO_3420 (O_3420,N_27577,N_27968);
and UO_3421 (O_3421,N_29239,N_29719);
nor UO_3422 (O_3422,N_29890,N_27645);
xor UO_3423 (O_3423,N_28133,N_29186);
and UO_3424 (O_3424,N_27752,N_29211);
or UO_3425 (O_3425,N_29206,N_29704);
nor UO_3426 (O_3426,N_28788,N_28228);
and UO_3427 (O_3427,N_29752,N_29086);
and UO_3428 (O_3428,N_29327,N_27328);
nand UO_3429 (O_3429,N_27319,N_29764);
xor UO_3430 (O_3430,N_27462,N_28056);
xor UO_3431 (O_3431,N_29730,N_28703);
and UO_3432 (O_3432,N_29940,N_29254);
nor UO_3433 (O_3433,N_28924,N_27739);
or UO_3434 (O_3434,N_29619,N_29198);
or UO_3435 (O_3435,N_28581,N_29795);
nor UO_3436 (O_3436,N_28963,N_29418);
and UO_3437 (O_3437,N_28955,N_27877);
and UO_3438 (O_3438,N_28972,N_27164);
or UO_3439 (O_3439,N_28880,N_28498);
xor UO_3440 (O_3440,N_29409,N_28995);
nor UO_3441 (O_3441,N_27836,N_28736);
or UO_3442 (O_3442,N_27937,N_29854);
and UO_3443 (O_3443,N_28914,N_28435);
nand UO_3444 (O_3444,N_27116,N_29795);
and UO_3445 (O_3445,N_27031,N_29651);
nor UO_3446 (O_3446,N_27332,N_27815);
and UO_3447 (O_3447,N_27963,N_29726);
nor UO_3448 (O_3448,N_28220,N_28479);
and UO_3449 (O_3449,N_27048,N_29002);
xor UO_3450 (O_3450,N_27942,N_29301);
nor UO_3451 (O_3451,N_27976,N_28303);
nand UO_3452 (O_3452,N_28219,N_29874);
nor UO_3453 (O_3453,N_29303,N_27036);
and UO_3454 (O_3454,N_29009,N_29426);
nand UO_3455 (O_3455,N_28043,N_28771);
nand UO_3456 (O_3456,N_28554,N_28666);
nor UO_3457 (O_3457,N_27860,N_28066);
or UO_3458 (O_3458,N_27155,N_29677);
or UO_3459 (O_3459,N_27328,N_27252);
xnor UO_3460 (O_3460,N_28575,N_29986);
nor UO_3461 (O_3461,N_27959,N_28752);
or UO_3462 (O_3462,N_28840,N_28451);
and UO_3463 (O_3463,N_29839,N_27053);
nand UO_3464 (O_3464,N_27921,N_29571);
and UO_3465 (O_3465,N_27587,N_27843);
and UO_3466 (O_3466,N_28267,N_29432);
nand UO_3467 (O_3467,N_27634,N_29736);
and UO_3468 (O_3468,N_28575,N_27543);
and UO_3469 (O_3469,N_28705,N_29252);
or UO_3470 (O_3470,N_29063,N_28713);
nor UO_3471 (O_3471,N_29551,N_27980);
nand UO_3472 (O_3472,N_27235,N_28172);
and UO_3473 (O_3473,N_27434,N_27102);
nand UO_3474 (O_3474,N_28962,N_29381);
or UO_3475 (O_3475,N_28594,N_28743);
nand UO_3476 (O_3476,N_27009,N_27569);
or UO_3477 (O_3477,N_29687,N_27644);
or UO_3478 (O_3478,N_27454,N_29130);
and UO_3479 (O_3479,N_29348,N_28760);
and UO_3480 (O_3480,N_27227,N_28998);
and UO_3481 (O_3481,N_29247,N_28911);
and UO_3482 (O_3482,N_27879,N_29983);
xor UO_3483 (O_3483,N_29593,N_28751);
nand UO_3484 (O_3484,N_27598,N_27968);
nand UO_3485 (O_3485,N_29261,N_27544);
xnor UO_3486 (O_3486,N_27414,N_29259);
xor UO_3487 (O_3487,N_29914,N_29643);
xor UO_3488 (O_3488,N_28180,N_29385);
nand UO_3489 (O_3489,N_27248,N_29134);
nand UO_3490 (O_3490,N_28293,N_27603);
and UO_3491 (O_3491,N_29891,N_29736);
xor UO_3492 (O_3492,N_28495,N_27292);
xnor UO_3493 (O_3493,N_29809,N_28177);
nand UO_3494 (O_3494,N_27461,N_27806);
xnor UO_3495 (O_3495,N_29502,N_29600);
xor UO_3496 (O_3496,N_29292,N_27066);
xor UO_3497 (O_3497,N_27958,N_27474);
nor UO_3498 (O_3498,N_29659,N_29573);
nand UO_3499 (O_3499,N_28314,N_27688);
endmodule