module basic_1500_15000_2000_5_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1028,In_146);
or U1 (N_1,In_1246,In_910);
nand U2 (N_2,In_788,In_992);
or U3 (N_3,In_50,In_1442);
nor U4 (N_4,In_1334,In_204);
nand U5 (N_5,In_22,In_16);
nor U6 (N_6,In_449,In_1040);
and U7 (N_7,In_969,In_809);
nor U8 (N_8,In_859,In_678);
nor U9 (N_9,In_1431,In_1187);
nand U10 (N_10,In_822,In_1109);
and U11 (N_11,In_1020,In_1);
and U12 (N_12,In_128,In_780);
and U13 (N_13,In_573,In_1116);
nand U14 (N_14,In_4,In_464);
nor U15 (N_15,In_173,In_530);
or U16 (N_16,In_946,In_862);
nand U17 (N_17,In_1151,In_781);
nor U18 (N_18,In_91,In_219);
nand U19 (N_19,In_268,In_262);
or U20 (N_20,In_792,In_1421);
and U21 (N_21,In_585,In_1093);
nor U22 (N_22,In_479,In_510);
or U23 (N_23,In_1495,In_309);
and U24 (N_24,In_1244,In_160);
and U25 (N_25,In_166,In_796);
and U26 (N_26,In_737,In_676);
nand U27 (N_27,In_328,In_88);
nor U28 (N_28,In_360,In_306);
or U29 (N_29,In_847,In_416);
or U30 (N_30,In_887,In_1272);
or U31 (N_31,In_1285,In_916);
and U32 (N_32,In_1132,In_839);
nor U33 (N_33,In_1158,In_388);
or U34 (N_34,In_1145,In_816);
nor U35 (N_35,In_455,In_611);
or U36 (N_36,In_801,In_852);
nand U37 (N_37,In_1265,In_866);
or U38 (N_38,In_55,In_448);
or U39 (N_39,In_123,In_130);
and U40 (N_40,In_831,In_138);
nand U41 (N_41,In_52,In_948);
nor U42 (N_42,In_263,In_951);
nand U43 (N_43,In_548,In_1408);
and U44 (N_44,In_1192,In_1140);
and U45 (N_45,In_243,In_1300);
or U46 (N_46,In_925,In_1181);
and U47 (N_47,In_715,In_1363);
nor U48 (N_48,In_979,In_838);
nand U49 (N_49,In_1423,In_987);
and U50 (N_50,In_407,In_963);
or U51 (N_51,In_217,In_1100);
and U52 (N_52,In_1207,In_352);
nand U53 (N_53,In_1266,In_1152);
nand U54 (N_54,In_1235,In_332);
nor U55 (N_55,In_149,In_1030);
nand U56 (N_56,In_1455,In_1149);
and U57 (N_57,In_708,In_711);
nor U58 (N_58,In_865,In_1464);
nor U59 (N_59,In_1419,In_1232);
nor U60 (N_60,In_895,In_919);
or U61 (N_61,In_1446,In_1163);
nand U62 (N_62,In_73,In_197);
and U63 (N_63,In_494,In_1198);
nor U64 (N_64,In_528,In_795);
nor U65 (N_65,In_356,In_329);
or U66 (N_66,In_325,In_456);
nor U67 (N_67,In_616,In_646);
nor U68 (N_68,In_1254,In_114);
and U69 (N_69,In_1486,In_286);
or U70 (N_70,In_1379,In_1171);
and U71 (N_71,In_391,In_512);
or U72 (N_72,In_480,In_421);
and U73 (N_73,In_302,In_563);
nand U74 (N_74,In_897,In_984);
or U75 (N_75,In_482,In_1064);
nand U76 (N_76,In_1258,In_470);
nor U77 (N_77,In_782,In_1425);
or U78 (N_78,In_1104,In_505);
and U79 (N_79,In_1186,In_888);
or U80 (N_80,In_769,In_1305);
nand U81 (N_81,In_1147,In_837);
or U82 (N_82,In_434,In_675);
nor U83 (N_83,In_1141,In_843);
nor U84 (N_84,In_600,In_1036);
nor U85 (N_85,In_1302,In_808);
and U86 (N_86,In_833,In_350);
nor U87 (N_87,In_1216,In_314);
nand U88 (N_88,In_1352,In_459);
and U89 (N_89,In_593,In_1470);
nand U90 (N_90,In_1007,In_376);
nor U91 (N_91,In_1489,In_1197);
nor U92 (N_92,In_107,In_1436);
and U93 (N_93,In_661,In_1347);
and U94 (N_94,In_962,In_763);
nor U95 (N_95,In_1478,In_1017);
nand U96 (N_96,In_518,In_985);
and U97 (N_97,In_829,In_1349);
nor U98 (N_98,In_275,In_519);
or U99 (N_99,In_187,In_1061);
nand U100 (N_100,In_484,In_1124);
or U101 (N_101,In_909,In_719);
or U102 (N_102,In_1125,In_259);
and U103 (N_103,In_31,In_136);
nor U104 (N_104,In_681,In_750);
or U105 (N_105,In_111,In_1103);
and U106 (N_106,In_1319,In_1062);
and U107 (N_107,In_604,In_72);
and U108 (N_108,In_1076,In_647);
nor U109 (N_109,In_30,In_165);
and U110 (N_110,In_569,In_1405);
and U111 (N_111,In_1383,In_522);
nand U112 (N_112,In_958,In_695);
or U113 (N_113,In_728,In_1251);
or U114 (N_114,In_23,In_297);
nand U115 (N_115,In_1194,In_1069);
nand U116 (N_116,In_981,In_747);
or U117 (N_117,In_516,In_1358);
or U118 (N_118,In_825,In_1080);
nor U119 (N_119,In_1282,In_742);
and U120 (N_120,In_806,In_924);
nand U121 (N_121,In_377,In_1038);
or U122 (N_122,In_1448,In_730);
nor U123 (N_123,In_1267,In_1435);
nand U124 (N_124,In_269,In_33);
or U125 (N_125,In_1023,In_367);
and U126 (N_126,In_1083,In_819);
and U127 (N_127,In_180,In_227);
or U128 (N_128,In_267,In_403);
nand U129 (N_129,In_353,In_755);
nor U130 (N_130,In_790,In_1430);
nand U131 (N_131,In_1463,In_1049);
nor U132 (N_132,In_1052,In_1137);
nand U133 (N_133,In_12,In_1233);
nor U134 (N_134,In_62,In_186);
or U135 (N_135,In_135,In_1362);
or U136 (N_136,In_282,In_236);
or U137 (N_137,In_95,In_599);
and U138 (N_138,In_1477,In_629);
nand U139 (N_139,In_734,In_64);
or U140 (N_140,In_882,In_840);
nand U141 (N_141,In_883,In_894);
and U142 (N_142,In_1184,In_460);
nor U143 (N_143,In_1086,In_504);
nand U144 (N_144,In_875,In_1209);
or U145 (N_145,In_454,In_818);
nor U146 (N_146,In_3,In_435);
nor U147 (N_147,In_1324,In_784);
nor U148 (N_148,In_145,In_982);
and U149 (N_149,In_553,In_1382);
and U150 (N_150,In_0,In_1058);
nand U151 (N_151,In_513,In_858);
nor U152 (N_152,In_190,In_581);
nor U153 (N_153,In_439,In_625);
or U154 (N_154,In_326,In_1240);
and U155 (N_155,In_1466,In_1013);
and U156 (N_156,In_1303,In_736);
and U157 (N_157,In_1097,In_85);
or U158 (N_158,In_1113,In_817);
or U159 (N_159,In_230,In_463);
and U160 (N_160,In_975,In_968);
or U161 (N_161,In_457,In_1139);
nor U162 (N_162,In_805,In_368);
or U163 (N_163,In_1433,In_578);
nor U164 (N_164,In_127,In_944);
nand U165 (N_165,In_891,In_1434);
nor U166 (N_166,In_498,In_1268);
nand U167 (N_167,In_500,In_557);
nand U168 (N_168,In_497,In_26);
nor U169 (N_169,In_802,In_659);
nor U170 (N_170,In_1066,In_966);
nand U171 (N_171,In_1160,In_890);
nor U172 (N_172,In_1351,In_879);
nand U173 (N_173,In_1111,In_66);
nand U174 (N_174,In_1309,In_154);
nand U175 (N_175,In_807,In_1173);
or U176 (N_176,In_233,In_687);
or U177 (N_177,In_184,In_405);
or U178 (N_178,In_697,In_287);
nand U179 (N_179,In_1467,In_1196);
or U180 (N_180,In_1420,In_797);
or U181 (N_181,In_168,In_1261);
and U182 (N_182,In_841,In_382);
nand U183 (N_183,In_637,In_252);
nand U184 (N_184,In_641,In_1317);
and U185 (N_185,In_560,In_598);
nand U186 (N_186,In_928,In_876);
and U187 (N_187,In_735,In_1475);
or U188 (N_188,In_359,In_621);
and U189 (N_189,In_874,In_814);
and U190 (N_190,In_1494,In_372);
nand U191 (N_191,In_904,In_108);
or U192 (N_192,In_1422,In_1117);
nor U193 (N_193,In_1273,In_583);
nor U194 (N_194,In_872,In_1380);
nor U195 (N_195,In_999,In_491);
nand U196 (N_196,In_1226,In_499);
or U197 (N_197,In_371,In_603);
nand U198 (N_198,In_1390,In_112);
nor U199 (N_199,In_358,In_1188);
nor U200 (N_200,In_644,In_988);
and U201 (N_201,In_972,In_273);
or U202 (N_202,In_922,In_673);
nand U203 (N_203,In_424,In_1174);
and U204 (N_204,In_1452,In_1316);
or U205 (N_205,In_82,In_486);
and U206 (N_206,In_1177,In_413);
nand U207 (N_207,In_532,In_59);
nor U208 (N_208,In_1329,In_726);
nand U209 (N_209,In_1264,In_634);
nand U210 (N_210,In_1243,In_283);
nand U211 (N_211,In_558,In_472);
nor U212 (N_212,In_467,In_250);
or U213 (N_213,In_447,In_947);
nor U214 (N_214,In_159,In_1195);
and U215 (N_215,In_871,In_1156);
or U216 (N_216,In_1108,In_1374);
nor U217 (N_217,In_257,In_907);
or U218 (N_218,In_1248,In_823);
nor U219 (N_219,In_1077,In_986);
nor U220 (N_220,In_789,In_773);
and U221 (N_221,In_702,In_465);
and U222 (N_222,In_760,In_1215);
or U223 (N_223,In_1284,In_76);
and U224 (N_224,In_244,In_713);
or U225 (N_225,In_543,In_152);
or U226 (N_226,In_1112,In_1450);
and U227 (N_227,In_1499,In_775);
and U228 (N_228,In_856,In_1353);
nand U229 (N_229,In_889,In_541);
or U230 (N_230,In_1418,In_520);
and U231 (N_231,In_638,In_1409);
and U232 (N_232,In_1260,In_693);
and U233 (N_233,In_620,In_1364);
and U234 (N_234,In_125,In_939);
nand U235 (N_235,In_1301,In_777);
nand U236 (N_236,In_949,In_361);
or U237 (N_237,In_1392,In_746);
or U238 (N_238,In_650,In_1288);
and U239 (N_239,In_234,In_635);
nor U240 (N_240,In_670,In_1332);
nor U241 (N_241,In_756,In_1231);
or U242 (N_242,In_835,In_1496);
or U243 (N_243,In_980,In_1126);
nor U244 (N_244,In_1131,In_1047);
and U245 (N_245,In_893,In_1255);
and U246 (N_246,In_140,In_663);
and U247 (N_247,In_177,In_60);
nor U248 (N_248,In_1032,In_1339);
nand U249 (N_249,In_442,In_1024);
nor U250 (N_250,In_685,In_926);
and U251 (N_251,In_509,In_526);
nand U252 (N_252,In_401,In_727);
and U253 (N_253,In_1458,In_546);
nor U254 (N_254,In_487,In_432);
or U255 (N_255,In_1414,In_853);
nand U256 (N_256,In_978,In_241);
and U257 (N_257,In_1019,In_343);
nor U258 (N_258,In_607,In_815);
nand U259 (N_259,In_716,In_1236);
nor U260 (N_260,In_478,In_799);
nor U261 (N_261,In_1468,In_1445);
or U262 (N_262,In_418,In_587);
nand U263 (N_263,In_993,In_100);
and U264 (N_264,In_1333,In_1043);
or U265 (N_265,In_1003,In_1089);
or U266 (N_266,In_458,In_193);
and U267 (N_267,In_515,In_1493);
nor U268 (N_268,In_466,In_864);
nor U269 (N_269,In_517,In_1189);
nand U270 (N_270,In_934,In_229);
and U271 (N_271,In_183,In_918);
nand U272 (N_272,In_813,In_395);
and U273 (N_273,In_28,In_9);
or U274 (N_274,In_115,In_1009);
nor U275 (N_275,In_609,In_586);
nor U276 (N_276,In_34,In_1081);
nor U277 (N_277,In_535,In_626);
and U278 (N_278,In_983,In_303);
nand U279 (N_279,In_249,In_613);
and U280 (N_280,In_1136,In_1110);
and U281 (N_281,In_161,In_1432);
and U282 (N_282,In_684,In_757);
nand U283 (N_283,In_57,In_741);
nor U284 (N_284,In_1277,In_355);
nand U285 (N_285,In_223,In_433);
nand U286 (N_286,In_696,In_568);
nand U287 (N_287,In_899,In_1296);
and U288 (N_288,In_246,In_631);
and U289 (N_289,In_1252,In_740);
and U290 (N_290,In_301,In_139);
or U291 (N_291,In_1087,In_554);
or U292 (N_292,In_25,In_1298);
or U293 (N_293,In_794,In_956);
nor U294 (N_294,In_492,In_102);
nor U295 (N_295,In_1299,In_271);
nor U296 (N_296,In_580,In_902);
and U297 (N_297,In_428,In_1487);
nor U298 (N_298,In_1008,In_1340);
or U299 (N_299,In_1403,In_1343);
or U300 (N_300,In_385,In_1262);
or U301 (N_301,In_1229,In_1391);
nor U302 (N_302,In_485,In_121);
nand U303 (N_303,In_1336,In_1142);
and U304 (N_304,In_258,In_1085);
and U305 (N_305,In_1063,In_61);
or U306 (N_306,In_1146,In_1004);
nand U307 (N_307,In_1135,In_288);
and U308 (N_308,In_1022,In_225);
or U309 (N_309,In_294,In_1201);
or U310 (N_310,In_253,In_1133);
nand U311 (N_311,In_1441,In_452);
and U312 (N_312,In_534,In_1401);
or U313 (N_313,In_821,In_63);
nand U314 (N_314,In_1016,In_1461);
and U315 (N_315,In_1230,In_590);
and U316 (N_316,In_200,In_1095);
or U317 (N_317,In_1031,In_148);
nor U318 (N_318,In_545,In_917);
and U319 (N_319,In_1393,In_251);
or U320 (N_320,In_991,In_705);
nor U321 (N_321,In_1271,In_654);
nor U322 (N_322,In_1479,In_1001);
and U323 (N_323,In_502,In_1480);
or U324 (N_324,In_709,In_1057);
and U325 (N_325,In_295,In_284);
nor U326 (N_326,In_83,In_364);
nand U327 (N_327,In_357,In_679);
or U328 (N_328,In_1078,In_1002);
nand U329 (N_329,In_1315,In_885);
nand U330 (N_330,In_1213,In_231);
nor U331 (N_331,In_1387,In_1015);
and U332 (N_332,In_778,In_164);
or U333 (N_333,In_1321,In_937);
or U334 (N_334,In_1042,In_701);
and U335 (N_335,In_1328,In_1119);
nand U336 (N_336,In_155,In_550);
nor U337 (N_337,In_195,In_722);
nor U338 (N_338,In_1044,In_1338);
nand U339 (N_339,In_768,In_717);
and U340 (N_340,In_221,In_908);
nand U341 (N_341,In_1386,In_44);
and U342 (N_342,In_666,In_913);
and U343 (N_343,In_338,In_1247);
and U344 (N_344,In_1313,In_1278);
and U345 (N_345,In_199,In_514);
or U346 (N_346,In_35,In_105);
nor U347 (N_347,In_1027,In_1400);
nor U348 (N_348,In_591,In_566);
or U349 (N_349,In_74,In_863);
nand U350 (N_350,In_191,In_1099);
and U351 (N_351,In_1384,In_386);
nor U352 (N_352,In_860,In_1484);
nand U353 (N_353,In_324,In_929);
or U354 (N_354,In_109,In_878);
or U355 (N_355,In_394,In_800);
xor U356 (N_356,In_451,In_436);
or U357 (N_357,In_540,In_1257);
nor U358 (N_358,In_213,In_1396);
and U359 (N_359,In_98,In_1227);
nand U360 (N_360,In_976,In_767);
nand U361 (N_361,In_335,In_559);
nor U362 (N_362,In_417,In_1105);
and U363 (N_363,In_627,In_153);
nand U364 (N_364,In_461,In_1449);
nor U365 (N_365,In_144,In_1394);
nand U366 (N_366,In_1465,In_349);
or U367 (N_367,In_1413,In_1385);
or U368 (N_368,In_653,In_363);
nor U369 (N_369,In_298,In_99);
or U370 (N_370,In_477,In_274);
and U371 (N_371,In_618,In_390);
and U372 (N_372,In_920,In_1367);
nor U373 (N_373,In_163,In_997);
nand U374 (N_374,In_1378,In_592);
nand U375 (N_375,In_1491,In_1217);
and U376 (N_376,In_345,In_1169);
and U377 (N_377,In_1033,In_998);
or U378 (N_378,In_495,In_201);
nand U379 (N_379,In_1327,In_48);
nor U380 (N_380,In_1427,In_446);
and U381 (N_381,In_1070,In_245);
nor U382 (N_382,In_1350,In_425);
nor U383 (N_383,In_232,In_277);
and U384 (N_384,In_1025,In_1286);
nor U385 (N_385,In_772,In_380);
and U386 (N_386,In_718,In_488);
or U387 (N_387,In_348,In_218);
and U388 (N_388,In_104,In_765);
nand U389 (N_389,In_450,In_84);
nor U390 (N_390,In_1256,In_178);
or U391 (N_391,In_1490,In_224);
xnor U392 (N_392,In_660,In_409);
or U393 (N_393,In_786,In_651);
nand U394 (N_394,In_1294,In_331);
nand U395 (N_395,In_158,In_1287);
or U396 (N_396,In_255,In_601);
nor U397 (N_397,In_266,In_444);
nor U398 (N_398,In_272,In_279);
or U399 (N_399,In_397,In_577);
and U400 (N_400,In_1498,In_851);
and U401 (N_401,In_720,In_933);
nand U402 (N_402,In_322,In_415);
nor U403 (N_403,In_898,In_336);
nor U404 (N_404,In_915,In_1344);
xnor U405 (N_405,In_539,In_285);
and U406 (N_406,In_13,In_776);
nand U407 (N_407,In_536,In_1457);
nand U408 (N_408,In_691,In_914);
and U409 (N_409,In_850,In_935);
or U410 (N_410,In_995,In_1325);
nand U411 (N_411,In_1067,In_1179);
nand U412 (N_412,In_698,In_1159);
nor U413 (N_413,In_174,In_855);
or U414 (N_414,In_1245,In_70);
and U415 (N_415,In_11,In_490);
nand U416 (N_416,In_1094,In_901);
nand U417 (N_417,In_443,In_1293);
or U418 (N_418,In_873,In_575);
and U419 (N_419,In_1492,In_1218);
or U420 (N_420,In_384,In_665);
nor U421 (N_421,In_402,In_633);
nor U422 (N_422,In_208,In_215);
nor U423 (N_423,In_207,In_688);
or U424 (N_424,In_316,In_533);
nor U425 (N_425,In_475,In_476);
or U426 (N_426,In_440,In_1454);
and U427 (N_427,In_45,In_1357);
or U428 (N_428,In_1118,In_759);
nor U429 (N_429,In_237,In_738);
nor U430 (N_430,In_1091,In_923);
or U431 (N_431,In_340,In_38);
nand U432 (N_432,In_1371,In_32);
and U433 (N_433,In_1395,In_18);
or U434 (N_434,In_1259,In_351);
nand U435 (N_435,In_643,In_552);
and U436 (N_436,In_751,In_724);
and U437 (N_437,In_496,In_1444);
nor U438 (N_438,In_1205,In_289);
or U439 (N_439,In_1176,In_181);
and U440 (N_440,In_753,In_315);
nand U441 (N_441,In_27,In_419);
nand U442 (N_442,In_1106,In_117);
xnor U443 (N_443,In_212,In_1279);
nor U444 (N_444,In_1138,In_20);
nand U445 (N_445,In_1134,In_828);
nor U446 (N_446,In_942,In_147);
or U447 (N_447,In_431,In_43);
nor U448 (N_448,In_206,In_375);
and U449 (N_449,In_39,In_820);
nor U450 (N_450,In_732,In_1453);
or U451 (N_451,In_1473,In_381);
nand U452 (N_452,In_1006,In_680);
or U453 (N_453,In_1308,In_1199);
or U454 (N_454,In_1055,In_523);
xor U455 (N_455,In_574,In_1084);
and U456 (N_456,In_589,In_369);
nand U457 (N_457,In_683,In_198);
nor U458 (N_458,In_967,In_378);
nor U459 (N_459,In_1148,In_555);
nand U460 (N_460,In_1348,In_1443);
nor U461 (N_461,In_1429,In_134);
nand U462 (N_462,In_414,In_1221);
nor U463 (N_463,In_1381,In_1045);
or U464 (N_464,In_320,In_542);
nor U465 (N_465,In_832,In_595);
nor U466 (N_466,In_1389,In_1053);
nor U467 (N_467,In_1424,In_362);
and U468 (N_468,In_672,In_1211);
nand U469 (N_469,In_1098,In_572);
and U470 (N_470,In_1361,In_779);
nor U471 (N_471,In_75,In_1191);
nand U472 (N_472,In_1280,In_119);
or U473 (N_473,In_1250,In_179);
nand U474 (N_474,In_132,In_994);
nand U475 (N_475,In_1356,In_1092);
and U476 (N_476,In_748,In_260);
nand U477 (N_477,In_1185,In_671);
nand U478 (N_478,In_1481,In_649);
nor U479 (N_479,In_81,In_142);
nand U480 (N_480,In_170,In_754);
nor U481 (N_481,In_1460,In_1346);
or U482 (N_482,In_202,In_655);
nand U483 (N_483,In_1406,In_1474);
nand U484 (N_484,In_1178,In_989);
nand U485 (N_485,In_196,In_133);
nand U486 (N_486,In_869,In_692);
nand U487 (N_487,In_971,In_339);
and U488 (N_488,In_667,In_596);
or U489 (N_489,In_1082,In_842);
and U490 (N_490,In_1456,In_86);
nand U491 (N_491,In_93,In_87);
nand U492 (N_492,In_602,In_1407);
nor U493 (N_493,In_588,In_80);
nand U494 (N_494,In_608,In_471);
and U495 (N_495,In_766,In_422);
nor U496 (N_496,In_892,In_867);
or U497 (N_497,In_468,In_1410);
nand U498 (N_498,In_830,In_1114);
xor U499 (N_499,In_764,In_712);
or U500 (N_500,In_549,In_96);
xor U501 (N_501,In_1129,In_5);
or U502 (N_502,In_323,In_1161);
and U503 (N_503,In_521,In_441);
nor U504 (N_504,In_725,In_406);
nor U505 (N_505,In_49,In_785);
or U506 (N_506,In_40,In_977);
or U507 (N_507,In_699,In_694);
and U508 (N_508,In_189,In_996);
nand U509 (N_509,In_974,In_636);
and U510 (N_510,In_1203,In_8);
and U511 (N_511,In_1154,In_1018);
nor U512 (N_512,In_551,In_1375);
or U513 (N_513,In_674,In_544);
or U514 (N_514,In_561,In_957);
nor U515 (N_515,In_1182,In_836);
nand U516 (N_516,In_228,In_392);
nand U517 (N_517,In_1297,In_354);
nand U518 (N_518,In_118,In_1295);
and U519 (N_519,In_365,In_1121);
nor U520 (N_520,In_167,In_143);
and U521 (N_521,In_1402,In_1289);
or U522 (N_522,In_597,In_664);
or U523 (N_523,In_46,In_296);
and U524 (N_524,In_749,In_743);
nand U525 (N_525,In_582,In_194);
or U526 (N_526,In_810,In_1497);
nor U527 (N_527,In_721,In_226);
or U528 (N_528,In_1071,In_529);
nor U529 (N_529,In_886,In_940);
or U530 (N_530,In_1214,In_71);
nand U531 (N_531,In_317,In_305);
and U532 (N_532,In_379,In_906);
nand U533 (N_533,In_10,In_411);
or U534 (N_534,In_19,In_176);
and U535 (N_535,In_1220,In_141);
nor U536 (N_536,In_739,In_921);
nand U537 (N_537,In_576,In_280);
nor U538 (N_538,In_952,In_579);
nand U539 (N_539,In_240,In_1360);
nor U540 (N_540,In_427,In_290);
nor U541 (N_541,In_68,In_1005);
nand U542 (N_542,In_622,In_483);
nor U543 (N_543,In_1276,In_333);
nor U544 (N_544,In_1482,In_826);
and U545 (N_545,In_489,In_56);
or U546 (N_546,In_430,In_344);
nor U547 (N_547,In_1090,In_1241);
nor U548 (N_548,In_399,In_1228);
or U549 (N_549,In_834,In_525);
nand U550 (N_550,In_758,In_624);
nand U551 (N_551,In_248,In_677);
and U552 (N_552,In_547,In_162);
or U553 (N_553,In_29,In_404);
nor U554 (N_554,In_564,In_945);
nor U555 (N_555,In_936,In_700);
and U556 (N_556,In_1167,In_17);
nor U557 (N_557,In_185,In_1370);
nor U558 (N_558,In_857,In_1404);
or U559 (N_559,In_222,In_106);
nand U560 (N_560,In_1292,In_1162);
or U561 (N_561,In_1000,In_1059);
nand U562 (N_562,In_53,In_733);
and U563 (N_563,In_209,In_1041);
nor U564 (N_564,In_1366,In_771);
nor U565 (N_565,In_1060,In_1183);
xnor U566 (N_566,In_342,In_689);
nor U567 (N_567,In_1314,In_192);
and U568 (N_568,In_1210,In_300);
and U569 (N_569,In_965,In_1311);
nor U570 (N_570,In_1029,In_437);
nor U571 (N_571,In_824,In_462);
nand U572 (N_572,In_304,In_723);
and U573 (N_573,In_1234,In_783);
and U574 (N_574,In_1107,In_126);
nor U575 (N_575,In_1281,In_1168);
and U576 (N_576,In_570,In_538);
nor U577 (N_577,In_710,In_1200);
or U578 (N_578,In_950,In_383);
or U579 (N_579,In_877,In_1075);
or U580 (N_580,In_931,In_341);
nand U581 (N_581,In_310,In_1068);
nor U582 (N_582,In_1373,In_150);
nor U583 (N_583,In_429,In_524);
or U584 (N_584,In_744,In_151);
or U585 (N_585,In_1144,In_51);
nor U586 (N_586,In_1337,In_1253);
and U587 (N_587,In_930,In_1291);
nand U588 (N_588,In_265,In_1331);
nor U589 (N_589,In_205,In_630);
nand U590 (N_590,In_619,In_506);
nor U591 (N_591,In_1415,In_129);
and U592 (N_592,In_1322,In_973);
xor U593 (N_593,In_400,In_270);
nand U594 (N_594,In_1115,In_1355);
nor U595 (N_595,In_188,In_242);
or U596 (N_596,In_256,In_426);
and U597 (N_597,In_1354,In_169);
nor U598 (N_598,In_849,In_1225);
nor U599 (N_599,In_1050,In_327);
nand U600 (N_600,In_238,In_182);
nand U601 (N_601,In_493,In_1485);
and U602 (N_602,In_903,In_157);
and U603 (N_603,In_374,In_373);
nand U604 (N_604,In_1438,In_1072);
nor U605 (N_605,In_1368,In_276);
nor U606 (N_606,In_941,In_1310);
nand U607 (N_607,In_884,In_1440);
or U608 (N_608,In_501,In_642);
nand U609 (N_609,In_77,In_1014);
nand U610 (N_610,In_905,In_704);
nor U611 (N_611,In_1306,In_1073);
nor U612 (N_612,In_299,In_1372);
nor U613 (N_613,In_214,In_1054);
or U614 (N_614,In_706,In_210);
and U615 (N_615,In_658,In_292);
or U616 (N_616,In_628,In_1170);
nor U617 (N_617,In_669,In_1462);
or U618 (N_618,In_1439,In_247);
nor U619 (N_619,In_1102,In_278);
or U620 (N_620,In_211,In_932);
nor U621 (N_621,In_110,In_752);
and U622 (N_622,In_1039,In_1483);
nand U623 (N_623,In_330,In_36);
nor U624 (N_624,In_1012,In_714);
and U625 (N_625,In_1312,In_1369);
and U626 (N_626,In_798,In_175);
nand U627 (N_627,In_645,In_1065);
or U628 (N_628,In_6,In_1239);
and U629 (N_629,In_1208,In_707);
nand U630 (N_630,In_396,In_1304);
nor U631 (N_631,In_648,In_97);
nand U632 (N_632,In_24,In_313);
or U633 (N_633,In_662,In_762);
xor U634 (N_634,In_1101,In_1175);
nor U635 (N_635,In_481,In_1342);
or U636 (N_636,In_1153,In_1204);
nand U637 (N_637,In_1290,In_565);
xnor U638 (N_638,In_293,In_1283);
nor U639 (N_639,In_900,In_1172);
and U640 (N_640,In_1451,In_594);
or U641 (N_641,In_235,In_1488);
nor U642 (N_642,In_1193,In_868);
or U643 (N_643,In_511,In_1237);
and U644 (N_644,In_1224,In_632);
and U645 (N_645,In_116,In_1021);
or U646 (N_646,In_961,In_1471);
and U647 (N_647,In_562,In_531);
and U648 (N_648,In_47,In_21);
and U649 (N_649,In_571,In_408);
nand U650 (N_650,In_387,In_473);
or U651 (N_651,In_346,In_870);
or U652 (N_652,In_1164,In_682);
and U653 (N_653,In_281,In_970);
nor U654 (N_654,In_1096,In_438);
nand U655 (N_655,In_845,In_1426);
and U656 (N_656,In_1128,In_1143);
nand U657 (N_657,In_612,In_1472);
nand U658 (N_658,In_1051,In_291);
nor U659 (N_659,In_774,In_453);
and U660 (N_660,In_1377,In_803);
nand U661 (N_661,In_261,In_124);
or U662 (N_662,In_7,In_912);
nor U663 (N_663,In_171,In_527);
or U664 (N_664,In_1155,In_469);
and U665 (N_665,In_605,In_2);
nand U666 (N_666,In_854,In_94);
nor U667 (N_667,In_122,In_445);
nor U668 (N_668,In_321,In_1242);
or U669 (N_669,In_761,In_37);
and U670 (N_670,In_308,In_1165);
or U671 (N_671,In_953,In_990);
or U672 (N_672,In_41,In_54);
or U673 (N_673,In_1341,In_312);
nand U674 (N_674,In_1323,In_65);
or U675 (N_675,In_264,In_927);
or U676 (N_676,In_216,In_307);
and U677 (N_677,In_1202,In_423);
nand U678 (N_678,In_793,In_337);
or U679 (N_679,In_861,In_652);
xor U680 (N_680,In_896,In_334);
or U681 (N_681,In_311,In_1222);
and U682 (N_682,In_614,In_955);
nor U683 (N_683,In_319,In_1330);
nor U684 (N_684,In_1447,In_1411);
nand U685 (N_685,In_318,In_610);
nand U686 (N_686,In_69,In_880);
and U687 (N_687,In_1011,In_556);
and U688 (N_688,In_156,In_812);
or U689 (N_689,In_1270,In_1223);
nor U690 (N_690,In_1326,In_881);
or U691 (N_691,In_960,In_729);
nor U692 (N_692,In_615,In_811);
nand U693 (N_693,In_1249,In_656);
and U694 (N_694,In_393,In_1010);
or U695 (N_695,In_1398,In_92);
nand U696 (N_696,In_254,In_58);
nor U697 (N_697,In_567,In_389);
nor U698 (N_698,In_639,In_1088);
and U699 (N_699,In_137,In_791);
and U700 (N_700,In_1476,In_15);
or U701 (N_701,In_938,In_1034);
and U702 (N_702,In_943,In_67);
nor U703 (N_703,In_347,In_1238);
or U704 (N_704,In_103,In_1219);
nor U705 (N_705,In_1275,In_1026);
nand U706 (N_706,In_846,In_420);
nor U707 (N_707,In_844,In_1274);
and U708 (N_708,In_78,In_1166);
or U709 (N_709,In_101,In_537);
and U710 (N_710,In_370,In_113);
or U711 (N_711,In_640,In_1376);
nor U712 (N_712,In_1157,In_398);
nor U713 (N_713,In_686,In_1035);
nand U714 (N_714,In_827,In_954);
and U715 (N_715,In_1190,In_1345);
nand U716 (N_716,In_203,In_42);
nor U717 (N_717,In_1318,In_657);
or U718 (N_718,In_1417,In_90);
or U719 (N_719,In_1048,In_1335);
and U720 (N_720,In_120,In_1359);
or U721 (N_721,In_131,In_220);
nor U722 (N_722,In_1469,In_239);
or U723 (N_723,In_1037,In_1046);
or U724 (N_724,In_1123,In_508);
nor U725 (N_725,In_14,In_1130);
or U726 (N_726,In_412,In_503);
nand U727 (N_727,In_911,In_1120);
and U728 (N_728,In_1180,In_1399);
or U729 (N_729,In_507,In_1365);
nor U730 (N_730,In_1269,In_668);
nand U731 (N_731,In_606,In_731);
or U732 (N_732,In_79,In_1459);
and U733 (N_733,In_1212,In_964);
or U734 (N_734,In_617,In_172);
or U735 (N_735,In_1079,In_623);
or U736 (N_736,In_1206,In_690);
and U737 (N_737,In_1307,In_1074);
and U738 (N_738,In_366,In_770);
nand U739 (N_739,In_1388,In_959);
nand U740 (N_740,In_584,In_1428);
nand U741 (N_741,In_1397,In_804);
and U742 (N_742,In_787,In_1412);
nand U743 (N_743,In_1127,In_1437);
nand U744 (N_744,In_1150,In_848);
and U745 (N_745,In_410,In_1416);
or U746 (N_746,In_89,In_474);
and U747 (N_747,In_1320,In_703);
or U748 (N_748,In_745,In_1056);
nand U749 (N_749,In_1122,In_1263);
or U750 (N_750,In_86,In_322);
or U751 (N_751,In_1321,In_877);
nand U752 (N_752,In_328,In_789);
nor U753 (N_753,In_671,In_1148);
and U754 (N_754,In_1045,In_896);
nor U755 (N_755,In_51,In_819);
nor U756 (N_756,In_690,In_551);
nand U757 (N_757,In_534,In_214);
or U758 (N_758,In_982,In_109);
nor U759 (N_759,In_485,In_994);
nand U760 (N_760,In_130,In_254);
nor U761 (N_761,In_583,In_506);
or U762 (N_762,In_1311,In_984);
and U763 (N_763,In_1041,In_248);
nand U764 (N_764,In_709,In_779);
nor U765 (N_765,In_1002,In_1339);
or U766 (N_766,In_1366,In_1130);
nand U767 (N_767,In_1319,In_479);
nor U768 (N_768,In_42,In_179);
and U769 (N_769,In_794,In_363);
or U770 (N_770,In_1399,In_385);
nand U771 (N_771,In_255,In_684);
and U772 (N_772,In_583,In_965);
nor U773 (N_773,In_980,In_622);
nor U774 (N_774,In_1012,In_1317);
or U775 (N_775,In_840,In_26);
nor U776 (N_776,In_57,In_1074);
and U777 (N_777,In_635,In_1472);
nor U778 (N_778,In_1303,In_1467);
or U779 (N_779,In_234,In_947);
xor U780 (N_780,In_1162,In_917);
or U781 (N_781,In_653,In_218);
or U782 (N_782,In_1082,In_86);
or U783 (N_783,In_1192,In_618);
nor U784 (N_784,In_919,In_552);
and U785 (N_785,In_422,In_92);
and U786 (N_786,In_1372,In_1035);
and U787 (N_787,In_363,In_465);
nor U788 (N_788,In_184,In_1193);
and U789 (N_789,In_943,In_1467);
nand U790 (N_790,In_984,In_538);
nand U791 (N_791,In_517,In_1260);
and U792 (N_792,In_1371,In_1122);
xnor U793 (N_793,In_885,In_1426);
nor U794 (N_794,In_1365,In_477);
and U795 (N_795,In_589,In_961);
nor U796 (N_796,In_425,In_26);
or U797 (N_797,In_1424,In_1073);
nor U798 (N_798,In_215,In_1017);
nand U799 (N_799,In_881,In_504);
nor U800 (N_800,In_1228,In_696);
and U801 (N_801,In_1443,In_638);
nor U802 (N_802,In_386,In_979);
or U803 (N_803,In_814,In_676);
or U804 (N_804,In_121,In_709);
or U805 (N_805,In_46,In_723);
nor U806 (N_806,In_752,In_305);
nand U807 (N_807,In_256,In_1421);
and U808 (N_808,In_1456,In_1331);
nor U809 (N_809,In_712,In_6);
or U810 (N_810,In_1343,In_504);
nand U811 (N_811,In_1152,In_360);
and U812 (N_812,In_395,In_748);
nor U813 (N_813,In_663,In_1391);
nor U814 (N_814,In_438,In_83);
or U815 (N_815,In_497,In_1144);
nor U816 (N_816,In_781,In_898);
and U817 (N_817,In_948,In_1209);
nand U818 (N_818,In_545,In_838);
nor U819 (N_819,In_540,In_1361);
or U820 (N_820,In_871,In_1146);
and U821 (N_821,In_1173,In_1169);
or U822 (N_822,In_815,In_759);
nand U823 (N_823,In_235,In_1147);
and U824 (N_824,In_365,In_1304);
nand U825 (N_825,In_1306,In_372);
nand U826 (N_826,In_45,In_1235);
xnor U827 (N_827,In_789,In_1105);
nand U828 (N_828,In_1384,In_1377);
nor U829 (N_829,In_1094,In_1233);
nor U830 (N_830,In_464,In_90);
xnor U831 (N_831,In_371,In_597);
and U832 (N_832,In_640,In_420);
nor U833 (N_833,In_1294,In_718);
nand U834 (N_834,In_211,In_642);
and U835 (N_835,In_531,In_701);
and U836 (N_836,In_1305,In_1417);
nor U837 (N_837,In_687,In_244);
and U838 (N_838,In_707,In_514);
or U839 (N_839,In_585,In_569);
or U840 (N_840,In_850,In_1018);
or U841 (N_841,In_303,In_564);
nand U842 (N_842,In_282,In_391);
nand U843 (N_843,In_33,In_603);
or U844 (N_844,In_131,In_1056);
and U845 (N_845,In_712,In_770);
and U846 (N_846,In_516,In_66);
nand U847 (N_847,In_688,In_405);
nor U848 (N_848,In_970,In_393);
nor U849 (N_849,In_572,In_701);
or U850 (N_850,In_56,In_962);
and U851 (N_851,In_1009,In_151);
or U852 (N_852,In_431,In_0);
nand U853 (N_853,In_274,In_543);
or U854 (N_854,In_697,In_1044);
nand U855 (N_855,In_1150,In_873);
or U856 (N_856,In_358,In_309);
nand U857 (N_857,In_1110,In_426);
or U858 (N_858,In_1394,In_476);
nand U859 (N_859,In_883,In_1474);
nand U860 (N_860,In_1013,In_731);
and U861 (N_861,In_441,In_722);
or U862 (N_862,In_1401,In_1245);
nor U863 (N_863,In_1077,In_537);
and U864 (N_864,In_759,In_1478);
or U865 (N_865,In_1347,In_0);
nand U866 (N_866,In_665,In_460);
and U867 (N_867,In_611,In_476);
nand U868 (N_868,In_356,In_1431);
and U869 (N_869,In_886,In_1018);
nand U870 (N_870,In_790,In_1451);
or U871 (N_871,In_1385,In_1005);
or U872 (N_872,In_383,In_1281);
or U873 (N_873,In_445,In_1007);
nand U874 (N_874,In_1333,In_1265);
nor U875 (N_875,In_1400,In_685);
or U876 (N_876,In_717,In_313);
or U877 (N_877,In_1278,In_507);
nor U878 (N_878,In_1030,In_410);
or U879 (N_879,In_998,In_174);
nand U880 (N_880,In_254,In_136);
and U881 (N_881,In_5,In_756);
nand U882 (N_882,In_615,In_358);
and U883 (N_883,In_1065,In_1150);
nor U884 (N_884,In_644,In_304);
nand U885 (N_885,In_525,In_93);
or U886 (N_886,In_1000,In_117);
and U887 (N_887,In_424,In_1164);
nand U888 (N_888,In_729,In_696);
nand U889 (N_889,In_362,In_1328);
nand U890 (N_890,In_1045,In_1480);
or U891 (N_891,In_20,In_789);
or U892 (N_892,In_1091,In_811);
nand U893 (N_893,In_563,In_739);
and U894 (N_894,In_498,In_1055);
and U895 (N_895,In_446,In_126);
nor U896 (N_896,In_985,In_945);
nand U897 (N_897,In_248,In_280);
nor U898 (N_898,In_463,In_1338);
nand U899 (N_899,In_1305,In_491);
and U900 (N_900,In_1353,In_21);
and U901 (N_901,In_869,In_861);
or U902 (N_902,In_750,In_1239);
nand U903 (N_903,In_939,In_754);
or U904 (N_904,In_281,In_788);
or U905 (N_905,In_8,In_1253);
nand U906 (N_906,In_160,In_866);
and U907 (N_907,In_771,In_844);
nand U908 (N_908,In_341,In_1397);
and U909 (N_909,In_1393,In_1001);
or U910 (N_910,In_1497,In_229);
nor U911 (N_911,In_315,In_1496);
or U912 (N_912,In_3,In_389);
nand U913 (N_913,In_15,In_1357);
or U914 (N_914,In_557,In_534);
nor U915 (N_915,In_507,In_460);
nor U916 (N_916,In_1408,In_1464);
nor U917 (N_917,In_810,In_598);
nand U918 (N_918,In_1361,In_1009);
nand U919 (N_919,In_549,In_1317);
nand U920 (N_920,In_60,In_229);
or U921 (N_921,In_764,In_706);
nand U922 (N_922,In_200,In_34);
nor U923 (N_923,In_164,In_496);
nand U924 (N_924,In_1490,In_745);
or U925 (N_925,In_1132,In_307);
or U926 (N_926,In_1067,In_955);
and U927 (N_927,In_1253,In_676);
nand U928 (N_928,In_1090,In_593);
or U929 (N_929,In_580,In_949);
nand U930 (N_930,In_368,In_950);
and U931 (N_931,In_89,In_958);
nor U932 (N_932,In_1233,In_1303);
or U933 (N_933,In_117,In_795);
and U934 (N_934,In_115,In_470);
nor U935 (N_935,In_358,In_465);
nor U936 (N_936,In_924,In_49);
or U937 (N_937,In_1265,In_779);
nand U938 (N_938,In_366,In_1144);
nor U939 (N_939,In_383,In_262);
nor U940 (N_940,In_824,In_217);
or U941 (N_941,In_393,In_1316);
or U942 (N_942,In_1415,In_220);
nor U943 (N_943,In_75,In_2);
or U944 (N_944,In_970,In_969);
or U945 (N_945,In_166,In_379);
nand U946 (N_946,In_924,In_423);
xor U947 (N_947,In_1228,In_1372);
nor U948 (N_948,In_288,In_812);
and U949 (N_949,In_324,In_155);
and U950 (N_950,In_108,In_1020);
or U951 (N_951,In_156,In_118);
nor U952 (N_952,In_983,In_1483);
or U953 (N_953,In_1371,In_649);
or U954 (N_954,In_855,In_319);
and U955 (N_955,In_1309,In_733);
and U956 (N_956,In_51,In_1463);
nor U957 (N_957,In_601,In_436);
nor U958 (N_958,In_529,In_45);
and U959 (N_959,In_496,In_197);
or U960 (N_960,In_476,In_698);
and U961 (N_961,In_1017,In_591);
nand U962 (N_962,In_1137,In_26);
nor U963 (N_963,In_574,In_1491);
nor U964 (N_964,In_1098,In_1115);
and U965 (N_965,In_1223,In_935);
or U966 (N_966,In_992,In_1245);
nor U967 (N_967,In_1269,In_808);
nor U968 (N_968,In_108,In_1044);
or U969 (N_969,In_625,In_1314);
nand U970 (N_970,In_340,In_353);
or U971 (N_971,In_832,In_472);
or U972 (N_972,In_588,In_199);
nor U973 (N_973,In_999,In_424);
nor U974 (N_974,In_1294,In_179);
nand U975 (N_975,In_260,In_77);
and U976 (N_976,In_1026,In_1283);
nand U977 (N_977,In_381,In_977);
and U978 (N_978,In_657,In_388);
and U979 (N_979,In_54,In_1153);
or U980 (N_980,In_199,In_179);
nand U981 (N_981,In_661,In_615);
and U982 (N_982,In_1086,In_939);
nand U983 (N_983,In_1486,In_546);
and U984 (N_984,In_805,In_678);
nor U985 (N_985,In_92,In_335);
and U986 (N_986,In_655,In_1243);
nor U987 (N_987,In_76,In_666);
or U988 (N_988,In_1233,In_819);
or U989 (N_989,In_373,In_1149);
xor U990 (N_990,In_342,In_642);
and U991 (N_991,In_231,In_973);
or U992 (N_992,In_328,In_574);
or U993 (N_993,In_21,In_1322);
nor U994 (N_994,In_178,In_607);
and U995 (N_995,In_1468,In_49);
and U996 (N_996,In_1470,In_861);
nor U997 (N_997,In_271,In_485);
or U998 (N_998,In_849,In_939);
nand U999 (N_999,In_318,In_591);
nor U1000 (N_1000,In_617,In_682);
nand U1001 (N_1001,In_761,In_50);
and U1002 (N_1002,In_313,In_790);
or U1003 (N_1003,In_999,In_1198);
or U1004 (N_1004,In_973,In_1051);
or U1005 (N_1005,In_1010,In_1028);
or U1006 (N_1006,In_971,In_682);
and U1007 (N_1007,In_548,In_728);
nand U1008 (N_1008,In_421,In_89);
nand U1009 (N_1009,In_1193,In_710);
nand U1010 (N_1010,In_400,In_135);
nand U1011 (N_1011,In_869,In_263);
nand U1012 (N_1012,In_802,In_1457);
and U1013 (N_1013,In_427,In_330);
and U1014 (N_1014,In_946,In_58);
or U1015 (N_1015,In_269,In_912);
nor U1016 (N_1016,In_215,In_464);
or U1017 (N_1017,In_673,In_785);
and U1018 (N_1018,In_1053,In_324);
and U1019 (N_1019,In_913,In_1193);
nor U1020 (N_1020,In_370,In_1025);
nand U1021 (N_1021,In_373,In_1256);
and U1022 (N_1022,In_631,In_479);
or U1023 (N_1023,In_39,In_552);
nand U1024 (N_1024,In_962,In_447);
or U1025 (N_1025,In_458,In_785);
nor U1026 (N_1026,In_549,In_1262);
nor U1027 (N_1027,In_902,In_1260);
and U1028 (N_1028,In_1426,In_403);
and U1029 (N_1029,In_1114,In_1451);
or U1030 (N_1030,In_280,In_921);
or U1031 (N_1031,In_1294,In_691);
nor U1032 (N_1032,In_1315,In_40);
and U1033 (N_1033,In_481,In_1409);
and U1034 (N_1034,In_13,In_1151);
nor U1035 (N_1035,In_888,In_582);
nand U1036 (N_1036,In_628,In_211);
nand U1037 (N_1037,In_1493,In_822);
nor U1038 (N_1038,In_753,In_490);
and U1039 (N_1039,In_915,In_380);
and U1040 (N_1040,In_187,In_1426);
and U1041 (N_1041,In_327,In_656);
nand U1042 (N_1042,In_97,In_1155);
nor U1043 (N_1043,In_456,In_622);
nand U1044 (N_1044,In_1133,In_701);
or U1045 (N_1045,In_625,In_63);
nand U1046 (N_1046,In_492,In_521);
and U1047 (N_1047,In_572,In_371);
nor U1048 (N_1048,In_1055,In_843);
nor U1049 (N_1049,In_1287,In_349);
and U1050 (N_1050,In_99,In_933);
nand U1051 (N_1051,In_210,In_75);
or U1052 (N_1052,In_1037,In_483);
nor U1053 (N_1053,In_985,In_1096);
and U1054 (N_1054,In_397,In_607);
nand U1055 (N_1055,In_280,In_886);
xor U1056 (N_1056,In_1068,In_1471);
and U1057 (N_1057,In_458,In_1364);
nor U1058 (N_1058,In_520,In_939);
or U1059 (N_1059,In_348,In_709);
and U1060 (N_1060,In_264,In_225);
nor U1061 (N_1061,In_1038,In_27);
nand U1062 (N_1062,In_411,In_4);
nor U1063 (N_1063,In_455,In_1330);
or U1064 (N_1064,In_1259,In_1019);
and U1065 (N_1065,In_822,In_1080);
nand U1066 (N_1066,In_711,In_571);
or U1067 (N_1067,In_1070,In_326);
or U1068 (N_1068,In_279,In_1103);
nand U1069 (N_1069,In_333,In_965);
and U1070 (N_1070,In_746,In_666);
nor U1071 (N_1071,In_845,In_1211);
and U1072 (N_1072,In_457,In_507);
or U1073 (N_1073,In_908,In_983);
nand U1074 (N_1074,In_763,In_200);
nor U1075 (N_1075,In_1370,In_158);
nand U1076 (N_1076,In_1449,In_1038);
and U1077 (N_1077,In_1213,In_835);
nor U1078 (N_1078,In_1472,In_517);
nand U1079 (N_1079,In_850,In_1036);
nor U1080 (N_1080,In_494,In_1448);
or U1081 (N_1081,In_310,In_697);
and U1082 (N_1082,In_184,In_108);
nor U1083 (N_1083,In_876,In_552);
and U1084 (N_1084,In_1464,In_445);
or U1085 (N_1085,In_413,In_1130);
or U1086 (N_1086,In_671,In_1259);
nor U1087 (N_1087,In_371,In_1379);
nor U1088 (N_1088,In_314,In_1328);
nand U1089 (N_1089,In_1337,In_1071);
or U1090 (N_1090,In_1257,In_823);
or U1091 (N_1091,In_1201,In_552);
nor U1092 (N_1092,In_779,In_914);
and U1093 (N_1093,In_1337,In_1447);
and U1094 (N_1094,In_546,In_438);
or U1095 (N_1095,In_352,In_1142);
or U1096 (N_1096,In_365,In_306);
and U1097 (N_1097,In_336,In_225);
nor U1098 (N_1098,In_903,In_944);
and U1099 (N_1099,In_233,In_103);
nor U1100 (N_1100,In_790,In_235);
nand U1101 (N_1101,In_807,In_200);
or U1102 (N_1102,In_182,In_1080);
nor U1103 (N_1103,In_371,In_386);
nor U1104 (N_1104,In_1495,In_1042);
or U1105 (N_1105,In_484,In_1260);
nor U1106 (N_1106,In_1193,In_888);
or U1107 (N_1107,In_1442,In_269);
nor U1108 (N_1108,In_1287,In_1009);
or U1109 (N_1109,In_661,In_117);
and U1110 (N_1110,In_932,In_1210);
and U1111 (N_1111,In_246,In_706);
or U1112 (N_1112,In_722,In_342);
or U1113 (N_1113,In_1040,In_53);
or U1114 (N_1114,In_405,In_243);
and U1115 (N_1115,In_451,In_990);
nand U1116 (N_1116,In_33,In_260);
xor U1117 (N_1117,In_514,In_1444);
nor U1118 (N_1118,In_87,In_802);
nor U1119 (N_1119,In_745,In_1475);
and U1120 (N_1120,In_1341,In_274);
nand U1121 (N_1121,In_133,In_1073);
and U1122 (N_1122,In_881,In_1443);
or U1123 (N_1123,In_1366,In_662);
xnor U1124 (N_1124,In_1087,In_385);
nor U1125 (N_1125,In_1249,In_724);
nand U1126 (N_1126,In_258,In_376);
nand U1127 (N_1127,In_1261,In_1440);
nor U1128 (N_1128,In_1484,In_786);
and U1129 (N_1129,In_186,In_183);
nand U1130 (N_1130,In_693,In_1444);
nand U1131 (N_1131,In_828,In_1312);
nor U1132 (N_1132,In_132,In_873);
and U1133 (N_1133,In_717,In_1011);
and U1134 (N_1134,In_530,In_571);
and U1135 (N_1135,In_802,In_1329);
nor U1136 (N_1136,In_422,In_511);
and U1137 (N_1137,In_1410,In_1154);
nand U1138 (N_1138,In_1277,In_1484);
or U1139 (N_1139,In_1357,In_1390);
or U1140 (N_1140,In_1023,In_965);
or U1141 (N_1141,In_1417,In_1166);
nand U1142 (N_1142,In_1296,In_608);
nor U1143 (N_1143,In_220,In_638);
or U1144 (N_1144,In_616,In_676);
nor U1145 (N_1145,In_1303,In_560);
or U1146 (N_1146,In_621,In_1213);
nor U1147 (N_1147,In_391,In_313);
or U1148 (N_1148,In_1435,In_462);
or U1149 (N_1149,In_333,In_398);
and U1150 (N_1150,In_752,In_1005);
nand U1151 (N_1151,In_421,In_558);
nand U1152 (N_1152,In_1318,In_310);
and U1153 (N_1153,In_683,In_150);
nand U1154 (N_1154,In_444,In_467);
nand U1155 (N_1155,In_341,In_1327);
and U1156 (N_1156,In_980,In_991);
nand U1157 (N_1157,In_317,In_901);
nor U1158 (N_1158,In_1396,In_1144);
nor U1159 (N_1159,In_1281,In_977);
nor U1160 (N_1160,In_559,In_903);
and U1161 (N_1161,In_57,In_262);
or U1162 (N_1162,In_1189,In_578);
or U1163 (N_1163,In_403,In_1274);
nand U1164 (N_1164,In_1412,In_1308);
nand U1165 (N_1165,In_119,In_365);
and U1166 (N_1166,In_1252,In_709);
and U1167 (N_1167,In_265,In_271);
nand U1168 (N_1168,In_575,In_530);
and U1169 (N_1169,In_1249,In_1008);
and U1170 (N_1170,In_629,In_1284);
or U1171 (N_1171,In_986,In_1038);
nor U1172 (N_1172,In_82,In_786);
and U1173 (N_1173,In_293,In_1382);
and U1174 (N_1174,In_1340,In_975);
nor U1175 (N_1175,In_79,In_66);
and U1176 (N_1176,In_906,In_861);
or U1177 (N_1177,In_534,In_899);
and U1178 (N_1178,In_1052,In_977);
nand U1179 (N_1179,In_918,In_1295);
and U1180 (N_1180,In_12,In_787);
nand U1181 (N_1181,In_1028,In_765);
and U1182 (N_1182,In_926,In_615);
nand U1183 (N_1183,In_1339,In_593);
nand U1184 (N_1184,In_553,In_382);
nand U1185 (N_1185,In_335,In_1264);
nand U1186 (N_1186,In_1268,In_591);
nor U1187 (N_1187,In_1134,In_1262);
nand U1188 (N_1188,In_1267,In_115);
nor U1189 (N_1189,In_44,In_152);
or U1190 (N_1190,In_1213,In_657);
nand U1191 (N_1191,In_820,In_874);
nand U1192 (N_1192,In_1443,In_582);
nor U1193 (N_1193,In_1361,In_1407);
nand U1194 (N_1194,In_511,In_507);
or U1195 (N_1195,In_832,In_429);
nor U1196 (N_1196,In_862,In_527);
nand U1197 (N_1197,In_408,In_1460);
or U1198 (N_1198,In_522,In_488);
or U1199 (N_1199,In_1402,In_943);
nor U1200 (N_1200,In_758,In_383);
nand U1201 (N_1201,In_1218,In_259);
or U1202 (N_1202,In_71,In_1005);
or U1203 (N_1203,In_1195,In_956);
or U1204 (N_1204,In_984,In_736);
nand U1205 (N_1205,In_635,In_1143);
nand U1206 (N_1206,In_703,In_791);
or U1207 (N_1207,In_1300,In_1088);
nand U1208 (N_1208,In_157,In_1430);
nor U1209 (N_1209,In_617,In_598);
nand U1210 (N_1210,In_116,In_17);
and U1211 (N_1211,In_1189,In_468);
nand U1212 (N_1212,In_899,In_318);
or U1213 (N_1213,In_1081,In_744);
nand U1214 (N_1214,In_114,In_1170);
nor U1215 (N_1215,In_1397,In_1340);
or U1216 (N_1216,In_100,In_104);
or U1217 (N_1217,In_809,In_748);
or U1218 (N_1218,In_518,In_7);
nand U1219 (N_1219,In_397,In_399);
nor U1220 (N_1220,In_150,In_947);
nand U1221 (N_1221,In_402,In_1368);
nand U1222 (N_1222,In_1377,In_104);
and U1223 (N_1223,In_621,In_655);
or U1224 (N_1224,In_294,In_1295);
or U1225 (N_1225,In_145,In_731);
and U1226 (N_1226,In_112,In_455);
or U1227 (N_1227,In_1477,In_79);
or U1228 (N_1228,In_1338,In_330);
nor U1229 (N_1229,In_787,In_604);
or U1230 (N_1230,In_784,In_1013);
or U1231 (N_1231,In_117,In_88);
nor U1232 (N_1232,In_346,In_999);
and U1233 (N_1233,In_42,In_181);
nand U1234 (N_1234,In_917,In_852);
or U1235 (N_1235,In_524,In_1211);
or U1236 (N_1236,In_365,In_678);
nor U1237 (N_1237,In_428,In_319);
nand U1238 (N_1238,In_528,In_1004);
and U1239 (N_1239,In_670,In_190);
nor U1240 (N_1240,In_172,In_1239);
nor U1241 (N_1241,In_904,In_57);
nor U1242 (N_1242,In_819,In_336);
nor U1243 (N_1243,In_466,In_400);
and U1244 (N_1244,In_413,In_997);
nand U1245 (N_1245,In_1159,In_1483);
nor U1246 (N_1246,In_1378,In_636);
nor U1247 (N_1247,In_876,In_428);
or U1248 (N_1248,In_1366,In_234);
nor U1249 (N_1249,In_682,In_440);
or U1250 (N_1250,In_496,In_564);
or U1251 (N_1251,In_904,In_1434);
or U1252 (N_1252,In_37,In_38);
or U1253 (N_1253,In_181,In_484);
nand U1254 (N_1254,In_114,In_854);
nand U1255 (N_1255,In_728,In_692);
nor U1256 (N_1256,In_261,In_620);
nor U1257 (N_1257,In_1479,In_430);
nand U1258 (N_1258,In_1434,In_1336);
nor U1259 (N_1259,In_1087,In_661);
or U1260 (N_1260,In_1450,In_1198);
and U1261 (N_1261,In_575,In_395);
or U1262 (N_1262,In_606,In_1360);
xor U1263 (N_1263,In_361,In_49);
nand U1264 (N_1264,In_211,In_1069);
nor U1265 (N_1265,In_879,In_812);
nor U1266 (N_1266,In_1005,In_1207);
nand U1267 (N_1267,In_26,In_181);
or U1268 (N_1268,In_8,In_186);
nand U1269 (N_1269,In_987,In_387);
nand U1270 (N_1270,In_887,In_238);
nand U1271 (N_1271,In_1148,In_1064);
or U1272 (N_1272,In_996,In_1270);
or U1273 (N_1273,In_23,In_1178);
or U1274 (N_1274,In_1049,In_1210);
nand U1275 (N_1275,In_705,In_942);
nor U1276 (N_1276,In_1270,In_1146);
and U1277 (N_1277,In_59,In_698);
and U1278 (N_1278,In_1137,In_254);
and U1279 (N_1279,In_46,In_279);
and U1280 (N_1280,In_529,In_519);
or U1281 (N_1281,In_1230,In_179);
and U1282 (N_1282,In_239,In_1390);
or U1283 (N_1283,In_61,In_429);
and U1284 (N_1284,In_1008,In_1369);
nand U1285 (N_1285,In_92,In_1108);
nor U1286 (N_1286,In_16,In_675);
nand U1287 (N_1287,In_1370,In_904);
nor U1288 (N_1288,In_802,In_974);
or U1289 (N_1289,In_435,In_310);
nor U1290 (N_1290,In_555,In_1269);
nand U1291 (N_1291,In_627,In_2);
and U1292 (N_1292,In_1078,In_255);
and U1293 (N_1293,In_109,In_679);
or U1294 (N_1294,In_1301,In_1432);
nand U1295 (N_1295,In_190,In_233);
and U1296 (N_1296,In_1133,In_920);
or U1297 (N_1297,In_575,In_89);
or U1298 (N_1298,In_547,In_8);
nor U1299 (N_1299,In_189,In_896);
nor U1300 (N_1300,In_1315,In_901);
and U1301 (N_1301,In_1116,In_184);
or U1302 (N_1302,In_1337,In_123);
or U1303 (N_1303,In_397,In_1032);
nand U1304 (N_1304,In_1,In_938);
nand U1305 (N_1305,In_499,In_1068);
and U1306 (N_1306,In_290,In_219);
and U1307 (N_1307,In_1186,In_920);
nor U1308 (N_1308,In_161,In_1026);
nor U1309 (N_1309,In_1305,In_322);
nor U1310 (N_1310,In_819,In_203);
or U1311 (N_1311,In_1433,In_1442);
nand U1312 (N_1312,In_330,In_883);
nor U1313 (N_1313,In_1120,In_1286);
nand U1314 (N_1314,In_745,In_1198);
or U1315 (N_1315,In_98,In_65);
or U1316 (N_1316,In_311,In_126);
or U1317 (N_1317,In_310,In_829);
nor U1318 (N_1318,In_385,In_1164);
nor U1319 (N_1319,In_752,In_288);
nor U1320 (N_1320,In_285,In_1298);
nor U1321 (N_1321,In_1400,In_1028);
nand U1322 (N_1322,In_61,In_17);
or U1323 (N_1323,In_902,In_937);
nand U1324 (N_1324,In_1003,In_140);
nor U1325 (N_1325,In_525,In_944);
xor U1326 (N_1326,In_472,In_1229);
nor U1327 (N_1327,In_600,In_1268);
nor U1328 (N_1328,In_361,In_716);
nor U1329 (N_1329,In_1120,In_367);
or U1330 (N_1330,In_37,In_693);
xnor U1331 (N_1331,In_951,In_954);
and U1332 (N_1332,In_997,In_890);
nor U1333 (N_1333,In_844,In_215);
or U1334 (N_1334,In_194,In_1328);
or U1335 (N_1335,In_568,In_76);
or U1336 (N_1336,In_839,In_788);
nand U1337 (N_1337,In_752,In_320);
nand U1338 (N_1338,In_1213,In_1136);
and U1339 (N_1339,In_1336,In_1246);
nor U1340 (N_1340,In_439,In_84);
and U1341 (N_1341,In_562,In_175);
and U1342 (N_1342,In_193,In_550);
nor U1343 (N_1343,In_1108,In_1263);
xnor U1344 (N_1344,In_882,In_1485);
nor U1345 (N_1345,In_1179,In_1203);
nand U1346 (N_1346,In_215,In_1477);
nand U1347 (N_1347,In_139,In_75);
and U1348 (N_1348,In_140,In_989);
nand U1349 (N_1349,In_761,In_128);
nor U1350 (N_1350,In_249,In_1141);
and U1351 (N_1351,In_323,In_772);
nor U1352 (N_1352,In_1340,In_1401);
nor U1353 (N_1353,In_470,In_1345);
nor U1354 (N_1354,In_1223,In_1063);
and U1355 (N_1355,In_1397,In_963);
or U1356 (N_1356,In_250,In_118);
nor U1357 (N_1357,In_779,In_304);
nand U1358 (N_1358,In_1423,In_7);
or U1359 (N_1359,In_878,In_1203);
nor U1360 (N_1360,In_137,In_1440);
and U1361 (N_1361,In_777,In_409);
nor U1362 (N_1362,In_258,In_9);
or U1363 (N_1363,In_859,In_699);
or U1364 (N_1364,In_465,In_838);
or U1365 (N_1365,In_1498,In_227);
xnor U1366 (N_1366,In_553,In_1298);
or U1367 (N_1367,In_1285,In_1092);
nor U1368 (N_1368,In_808,In_1266);
nand U1369 (N_1369,In_425,In_1385);
nor U1370 (N_1370,In_875,In_1398);
nand U1371 (N_1371,In_395,In_297);
and U1372 (N_1372,In_323,In_1237);
nand U1373 (N_1373,In_444,In_181);
and U1374 (N_1374,In_1430,In_1170);
or U1375 (N_1375,In_1390,In_1275);
nand U1376 (N_1376,In_894,In_1322);
nor U1377 (N_1377,In_1000,In_1131);
or U1378 (N_1378,In_1422,In_851);
nand U1379 (N_1379,In_318,In_675);
nand U1380 (N_1380,In_34,In_622);
or U1381 (N_1381,In_1359,In_383);
and U1382 (N_1382,In_470,In_937);
or U1383 (N_1383,In_795,In_842);
nand U1384 (N_1384,In_111,In_1077);
nor U1385 (N_1385,In_782,In_38);
nor U1386 (N_1386,In_1298,In_1172);
nand U1387 (N_1387,In_707,In_541);
nor U1388 (N_1388,In_1348,In_313);
or U1389 (N_1389,In_231,In_194);
nand U1390 (N_1390,In_798,In_832);
or U1391 (N_1391,In_996,In_1150);
nand U1392 (N_1392,In_1363,In_155);
nand U1393 (N_1393,In_587,In_572);
nand U1394 (N_1394,In_1054,In_68);
and U1395 (N_1395,In_752,In_347);
and U1396 (N_1396,In_1209,In_1124);
nand U1397 (N_1397,In_462,In_197);
and U1398 (N_1398,In_329,In_948);
nor U1399 (N_1399,In_1320,In_411);
and U1400 (N_1400,In_961,In_787);
nand U1401 (N_1401,In_741,In_399);
nand U1402 (N_1402,In_435,In_538);
nor U1403 (N_1403,In_243,In_339);
nand U1404 (N_1404,In_962,In_847);
xor U1405 (N_1405,In_184,In_570);
and U1406 (N_1406,In_1033,In_918);
nor U1407 (N_1407,In_1356,In_280);
nor U1408 (N_1408,In_49,In_1270);
nand U1409 (N_1409,In_1395,In_1323);
nand U1410 (N_1410,In_202,In_567);
and U1411 (N_1411,In_210,In_1119);
or U1412 (N_1412,In_1312,In_534);
xor U1413 (N_1413,In_94,In_1097);
or U1414 (N_1414,In_68,In_1350);
or U1415 (N_1415,In_30,In_553);
nand U1416 (N_1416,In_486,In_1091);
nand U1417 (N_1417,In_55,In_1139);
and U1418 (N_1418,In_276,In_777);
nand U1419 (N_1419,In_613,In_131);
nand U1420 (N_1420,In_247,In_1209);
nor U1421 (N_1421,In_507,In_1043);
nand U1422 (N_1422,In_972,In_1438);
nand U1423 (N_1423,In_53,In_1239);
nand U1424 (N_1424,In_1095,In_1435);
or U1425 (N_1425,In_1438,In_1082);
and U1426 (N_1426,In_944,In_27);
and U1427 (N_1427,In_520,In_1103);
nand U1428 (N_1428,In_1414,In_230);
and U1429 (N_1429,In_769,In_411);
nor U1430 (N_1430,In_1196,In_1027);
nand U1431 (N_1431,In_1062,In_775);
and U1432 (N_1432,In_272,In_715);
nor U1433 (N_1433,In_1233,In_1122);
or U1434 (N_1434,In_993,In_547);
nor U1435 (N_1435,In_885,In_227);
or U1436 (N_1436,In_231,In_352);
nand U1437 (N_1437,In_1237,In_720);
or U1438 (N_1438,In_662,In_851);
nor U1439 (N_1439,In_148,In_669);
or U1440 (N_1440,In_1427,In_1133);
and U1441 (N_1441,In_1076,In_175);
nand U1442 (N_1442,In_1116,In_657);
or U1443 (N_1443,In_604,In_929);
and U1444 (N_1444,In_861,In_1120);
and U1445 (N_1445,In_558,In_770);
or U1446 (N_1446,In_835,In_1302);
nand U1447 (N_1447,In_70,In_246);
or U1448 (N_1448,In_828,In_1104);
or U1449 (N_1449,In_1272,In_672);
or U1450 (N_1450,In_1450,In_797);
nand U1451 (N_1451,In_596,In_1467);
nor U1452 (N_1452,In_1006,In_132);
and U1453 (N_1453,In_992,In_1481);
and U1454 (N_1454,In_830,In_123);
and U1455 (N_1455,In_1100,In_826);
nor U1456 (N_1456,In_14,In_107);
nor U1457 (N_1457,In_392,In_514);
and U1458 (N_1458,In_255,In_494);
nand U1459 (N_1459,In_394,In_1390);
or U1460 (N_1460,In_60,In_681);
and U1461 (N_1461,In_860,In_496);
and U1462 (N_1462,In_1342,In_849);
nor U1463 (N_1463,In_615,In_676);
or U1464 (N_1464,In_288,In_607);
nor U1465 (N_1465,In_1395,In_194);
nor U1466 (N_1466,In_826,In_799);
nor U1467 (N_1467,In_1362,In_508);
nand U1468 (N_1468,In_1173,In_224);
xnor U1469 (N_1469,In_827,In_341);
or U1470 (N_1470,In_311,In_50);
or U1471 (N_1471,In_385,In_1001);
and U1472 (N_1472,In_746,In_199);
and U1473 (N_1473,In_707,In_376);
or U1474 (N_1474,In_1031,In_117);
or U1475 (N_1475,In_1181,In_646);
nor U1476 (N_1476,In_276,In_1325);
nor U1477 (N_1477,In_1085,In_323);
nor U1478 (N_1478,In_836,In_820);
or U1479 (N_1479,In_107,In_226);
nand U1480 (N_1480,In_774,In_548);
nor U1481 (N_1481,In_783,In_177);
nand U1482 (N_1482,In_1209,In_69);
or U1483 (N_1483,In_252,In_819);
nor U1484 (N_1484,In_402,In_354);
nand U1485 (N_1485,In_1254,In_192);
and U1486 (N_1486,In_620,In_548);
or U1487 (N_1487,In_52,In_946);
and U1488 (N_1488,In_920,In_984);
nor U1489 (N_1489,In_5,In_99);
nor U1490 (N_1490,In_1364,In_14);
nand U1491 (N_1491,In_497,In_390);
nand U1492 (N_1492,In_876,In_1029);
nor U1493 (N_1493,In_768,In_1248);
nor U1494 (N_1494,In_34,In_1460);
and U1495 (N_1495,In_495,In_1126);
nor U1496 (N_1496,In_1163,In_48);
and U1497 (N_1497,In_274,In_986);
and U1498 (N_1498,In_1116,In_1333);
and U1499 (N_1499,In_747,In_387);
nor U1500 (N_1500,In_927,In_247);
nor U1501 (N_1501,In_1028,In_1072);
nand U1502 (N_1502,In_293,In_125);
and U1503 (N_1503,In_406,In_604);
nor U1504 (N_1504,In_969,In_1342);
nand U1505 (N_1505,In_44,In_790);
nand U1506 (N_1506,In_780,In_288);
nor U1507 (N_1507,In_689,In_484);
nor U1508 (N_1508,In_1197,In_309);
or U1509 (N_1509,In_1160,In_1218);
nand U1510 (N_1510,In_1425,In_379);
or U1511 (N_1511,In_1110,In_391);
and U1512 (N_1512,In_362,In_561);
or U1513 (N_1513,In_856,In_427);
nor U1514 (N_1514,In_581,In_4);
and U1515 (N_1515,In_1376,In_986);
nor U1516 (N_1516,In_973,In_1279);
nor U1517 (N_1517,In_29,In_1275);
or U1518 (N_1518,In_762,In_80);
nor U1519 (N_1519,In_1027,In_981);
and U1520 (N_1520,In_358,In_39);
nor U1521 (N_1521,In_1206,In_906);
and U1522 (N_1522,In_361,In_1108);
nor U1523 (N_1523,In_955,In_180);
or U1524 (N_1524,In_1351,In_190);
nand U1525 (N_1525,In_1056,In_409);
and U1526 (N_1526,In_332,In_573);
nand U1527 (N_1527,In_469,In_500);
and U1528 (N_1528,In_1289,In_1141);
nor U1529 (N_1529,In_41,In_1268);
or U1530 (N_1530,In_149,In_284);
and U1531 (N_1531,In_697,In_1205);
nor U1532 (N_1532,In_1334,In_565);
or U1533 (N_1533,In_1440,In_863);
and U1534 (N_1534,In_847,In_209);
nand U1535 (N_1535,In_724,In_1301);
nor U1536 (N_1536,In_1438,In_366);
or U1537 (N_1537,In_844,In_579);
and U1538 (N_1538,In_714,In_914);
nand U1539 (N_1539,In_992,In_4);
nand U1540 (N_1540,In_1190,In_180);
nand U1541 (N_1541,In_599,In_199);
nor U1542 (N_1542,In_1273,In_1018);
nand U1543 (N_1543,In_376,In_683);
or U1544 (N_1544,In_788,In_1416);
nand U1545 (N_1545,In_1343,In_762);
nand U1546 (N_1546,In_772,In_568);
nor U1547 (N_1547,In_549,In_57);
nand U1548 (N_1548,In_568,In_331);
xnor U1549 (N_1549,In_992,In_93);
or U1550 (N_1550,In_441,In_134);
and U1551 (N_1551,In_608,In_152);
nor U1552 (N_1552,In_767,In_511);
nand U1553 (N_1553,In_765,In_733);
nand U1554 (N_1554,In_519,In_564);
or U1555 (N_1555,In_818,In_1443);
nor U1556 (N_1556,In_446,In_287);
and U1557 (N_1557,In_865,In_41);
nand U1558 (N_1558,In_724,In_226);
and U1559 (N_1559,In_249,In_878);
nor U1560 (N_1560,In_1153,In_986);
nor U1561 (N_1561,In_657,In_1148);
xnor U1562 (N_1562,In_1245,In_115);
or U1563 (N_1563,In_288,In_1219);
nand U1564 (N_1564,In_195,In_1253);
or U1565 (N_1565,In_1195,In_1293);
and U1566 (N_1566,In_601,In_1139);
nor U1567 (N_1567,In_449,In_377);
nor U1568 (N_1568,In_597,In_48);
and U1569 (N_1569,In_838,In_609);
nand U1570 (N_1570,In_1144,In_1352);
nor U1571 (N_1571,In_153,In_1415);
nor U1572 (N_1572,In_363,In_1321);
and U1573 (N_1573,In_852,In_686);
or U1574 (N_1574,In_290,In_639);
and U1575 (N_1575,In_1282,In_338);
nor U1576 (N_1576,In_308,In_426);
or U1577 (N_1577,In_1272,In_1216);
and U1578 (N_1578,In_1269,In_1455);
and U1579 (N_1579,In_815,In_1276);
nor U1580 (N_1580,In_1109,In_1439);
or U1581 (N_1581,In_1366,In_811);
and U1582 (N_1582,In_86,In_1378);
or U1583 (N_1583,In_1247,In_22);
or U1584 (N_1584,In_404,In_974);
or U1585 (N_1585,In_550,In_1487);
nor U1586 (N_1586,In_335,In_330);
nand U1587 (N_1587,In_669,In_589);
nand U1588 (N_1588,In_587,In_334);
nand U1589 (N_1589,In_374,In_645);
xor U1590 (N_1590,In_186,In_1039);
nor U1591 (N_1591,In_636,In_583);
or U1592 (N_1592,In_1373,In_439);
or U1593 (N_1593,In_110,In_753);
or U1594 (N_1594,In_497,In_356);
nor U1595 (N_1595,In_1180,In_208);
nor U1596 (N_1596,In_1141,In_128);
nor U1597 (N_1597,In_357,In_569);
or U1598 (N_1598,In_559,In_53);
or U1599 (N_1599,In_298,In_486);
nor U1600 (N_1600,In_148,In_189);
or U1601 (N_1601,In_461,In_760);
nand U1602 (N_1602,In_1077,In_116);
xor U1603 (N_1603,In_78,In_1339);
and U1604 (N_1604,In_218,In_822);
nand U1605 (N_1605,In_366,In_279);
or U1606 (N_1606,In_1010,In_1447);
and U1607 (N_1607,In_949,In_740);
nor U1608 (N_1608,In_1366,In_1024);
nor U1609 (N_1609,In_412,In_281);
or U1610 (N_1610,In_66,In_1020);
nand U1611 (N_1611,In_821,In_52);
or U1612 (N_1612,In_723,In_627);
nor U1613 (N_1613,In_512,In_1150);
or U1614 (N_1614,In_1074,In_313);
nand U1615 (N_1615,In_1428,In_712);
nor U1616 (N_1616,In_1093,In_1142);
nand U1617 (N_1617,In_541,In_1444);
nand U1618 (N_1618,In_1062,In_764);
and U1619 (N_1619,In_119,In_379);
or U1620 (N_1620,In_1327,In_1260);
nand U1621 (N_1621,In_571,In_462);
nand U1622 (N_1622,In_1499,In_200);
nand U1623 (N_1623,In_605,In_239);
nand U1624 (N_1624,In_261,In_1072);
and U1625 (N_1625,In_786,In_231);
or U1626 (N_1626,In_1160,In_13);
nand U1627 (N_1627,In_934,In_1125);
nand U1628 (N_1628,In_971,In_137);
nor U1629 (N_1629,In_954,In_538);
or U1630 (N_1630,In_272,In_692);
nor U1631 (N_1631,In_1036,In_572);
nor U1632 (N_1632,In_457,In_56);
nor U1633 (N_1633,In_1240,In_11);
or U1634 (N_1634,In_102,In_995);
nor U1635 (N_1635,In_1279,In_63);
and U1636 (N_1636,In_1252,In_783);
nor U1637 (N_1637,In_534,In_1053);
xnor U1638 (N_1638,In_1175,In_1381);
or U1639 (N_1639,In_177,In_1358);
nand U1640 (N_1640,In_568,In_1256);
or U1641 (N_1641,In_993,In_448);
nor U1642 (N_1642,In_1139,In_1172);
and U1643 (N_1643,In_1342,In_981);
and U1644 (N_1644,In_843,In_260);
nor U1645 (N_1645,In_1201,In_894);
and U1646 (N_1646,In_587,In_371);
and U1647 (N_1647,In_250,In_988);
nor U1648 (N_1648,In_1053,In_147);
and U1649 (N_1649,In_475,In_1336);
nor U1650 (N_1650,In_657,In_273);
nor U1651 (N_1651,In_1075,In_1393);
or U1652 (N_1652,In_485,In_15);
or U1653 (N_1653,In_1306,In_361);
nand U1654 (N_1654,In_967,In_563);
nand U1655 (N_1655,In_1199,In_1478);
or U1656 (N_1656,In_1499,In_668);
or U1657 (N_1657,In_554,In_513);
and U1658 (N_1658,In_416,In_584);
nand U1659 (N_1659,In_958,In_857);
and U1660 (N_1660,In_738,In_881);
and U1661 (N_1661,In_1486,In_383);
nor U1662 (N_1662,In_1267,In_438);
nand U1663 (N_1663,In_1157,In_367);
or U1664 (N_1664,In_968,In_1283);
nand U1665 (N_1665,In_1096,In_946);
and U1666 (N_1666,In_1038,In_689);
nand U1667 (N_1667,In_809,In_771);
nor U1668 (N_1668,In_161,In_403);
or U1669 (N_1669,In_332,In_988);
nor U1670 (N_1670,In_396,In_1443);
or U1671 (N_1671,In_933,In_16);
nor U1672 (N_1672,In_791,In_948);
and U1673 (N_1673,In_239,In_1492);
and U1674 (N_1674,In_911,In_1201);
and U1675 (N_1675,In_135,In_8);
and U1676 (N_1676,In_484,In_864);
or U1677 (N_1677,In_899,In_1118);
nand U1678 (N_1678,In_605,In_1343);
nand U1679 (N_1679,In_1066,In_73);
nand U1680 (N_1680,In_1181,In_1013);
xor U1681 (N_1681,In_404,In_1134);
or U1682 (N_1682,In_881,In_779);
nor U1683 (N_1683,In_716,In_175);
nand U1684 (N_1684,In_50,In_493);
and U1685 (N_1685,In_80,In_957);
and U1686 (N_1686,In_1095,In_651);
or U1687 (N_1687,In_326,In_622);
nand U1688 (N_1688,In_1331,In_18);
or U1689 (N_1689,In_38,In_1428);
nand U1690 (N_1690,In_914,In_1469);
and U1691 (N_1691,In_585,In_625);
nand U1692 (N_1692,In_501,In_282);
nor U1693 (N_1693,In_325,In_198);
and U1694 (N_1694,In_1429,In_1453);
and U1695 (N_1695,In_517,In_2);
nor U1696 (N_1696,In_340,In_107);
or U1697 (N_1697,In_103,In_949);
and U1698 (N_1698,In_387,In_110);
nor U1699 (N_1699,In_1247,In_221);
and U1700 (N_1700,In_214,In_693);
and U1701 (N_1701,In_1255,In_1273);
or U1702 (N_1702,In_777,In_1247);
nor U1703 (N_1703,In_414,In_484);
or U1704 (N_1704,In_881,In_839);
nor U1705 (N_1705,In_1489,In_1483);
or U1706 (N_1706,In_877,In_545);
xor U1707 (N_1707,In_851,In_13);
and U1708 (N_1708,In_557,In_63);
nand U1709 (N_1709,In_603,In_778);
and U1710 (N_1710,In_1283,In_482);
nand U1711 (N_1711,In_120,In_335);
and U1712 (N_1712,In_512,In_362);
and U1713 (N_1713,In_1319,In_25);
and U1714 (N_1714,In_1070,In_996);
nor U1715 (N_1715,In_713,In_223);
or U1716 (N_1716,In_1173,In_709);
xnor U1717 (N_1717,In_1346,In_4);
nand U1718 (N_1718,In_711,In_1272);
and U1719 (N_1719,In_936,In_1416);
nor U1720 (N_1720,In_131,In_698);
nor U1721 (N_1721,In_744,In_322);
and U1722 (N_1722,In_673,In_1164);
nor U1723 (N_1723,In_446,In_284);
and U1724 (N_1724,In_75,In_86);
nor U1725 (N_1725,In_995,In_317);
or U1726 (N_1726,In_321,In_408);
and U1727 (N_1727,In_399,In_502);
nor U1728 (N_1728,In_857,In_1186);
or U1729 (N_1729,In_1218,In_868);
nor U1730 (N_1730,In_1345,In_308);
nor U1731 (N_1731,In_1484,In_1428);
and U1732 (N_1732,In_943,In_729);
nor U1733 (N_1733,In_700,In_1396);
or U1734 (N_1734,In_599,In_1087);
nor U1735 (N_1735,In_1023,In_1259);
nor U1736 (N_1736,In_1428,In_1110);
or U1737 (N_1737,In_730,In_976);
and U1738 (N_1738,In_553,In_235);
xnor U1739 (N_1739,In_114,In_726);
or U1740 (N_1740,In_1296,In_168);
or U1741 (N_1741,In_875,In_1337);
and U1742 (N_1742,In_212,In_388);
and U1743 (N_1743,In_209,In_46);
nor U1744 (N_1744,In_1166,In_695);
nor U1745 (N_1745,In_1178,In_482);
nand U1746 (N_1746,In_261,In_1052);
or U1747 (N_1747,In_42,In_271);
nand U1748 (N_1748,In_900,In_424);
nor U1749 (N_1749,In_144,In_376);
and U1750 (N_1750,In_1335,In_382);
or U1751 (N_1751,In_884,In_1411);
and U1752 (N_1752,In_849,In_2);
nor U1753 (N_1753,In_623,In_1340);
or U1754 (N_1754,In_275,In_1277);
or U1755 (N_1755,In_1431,In_767);
or U1756 (N_1756,In_1226,In_357);
or U1757 (N_1757,In_543,In_994);
or U1758 (N_1758,In_1292,In_1080);
or U1759 (N_1759,In_1008,In_1187);
nand U1760 (N_1760,In_397,In_1363);
nor U1761 (N_1761,In_196,In_1324);
and U1762 (N_1762,In_30,In_1039);
or U1763 (N_1763,In_734,In_1402);
nand U1764 (N_1764,In_482,In_1189);
nor U1765 (N_1765,In_582,In_1410);
nand U1766 (N_1766,In_222,In_81);
or U1767 (N_1767,In_77,In_93);
or U1768 (N_1768,In_1482,In_670);
or U1769 (N_1769,In_187,In_67);
and U1770 (N_1770,In_1404,In_437);
nand U1771 (N_1771,In_727,In_1006);
nor U1772 (N_1772,In_399,In_1065);
nor U1773 (N_1773,In_492,In_1364);
xnor U1774 (N_1774,In_661,In_645);
and U1775 (N_1775,In_812,In_484);
xnor U1776 (N_1776,In_762,In_792);
nor U1777 (N_1777,In_1393,In_456);
or U1778 (N_1778,In_1042,In_237);
or U1779 (N_1779,In_77,In_568);
xnor U1780 (N_1780,In_1004,In_1315);
and U1781 (N_1781,In_1420,In_1098);
and U1782 (N_1782,In_149,In_361);
nand U1783 (N_1783,In_138,In_1426);
or U1784 (N_1784,In_147,In_770);
and U1785 (N_1785,In_1103,In_1131);
nand U1786 (N_1786,In_1352,In_1179);
nand U1787 (N_1787,In_1173,In_1317);
nand U1788 (N_1788,In_1101,In_1275);
or U1789 (N_1789,In_996,In_1400);
and U1790 (N_1790,In_475,In_757);
and U1791 (N_1791,In_396,In_39);
and U1792 (N_1792,In_1036,In_78);
or U1793 (N_1793,In_1012,In_755);
and U1794 (N_1794,In_211,In_361);
or U1795 (N_1795,In_651,In_1176);
or U1796 (N_1796,In_979,In_247);
nor U1797 (N_1797,In_553,In_1105);
or U1798 (N_1798,In_677,In_1350);
nand U1799 (N_1799,In_479,In_686);
and U1800 (N_1800,In_409,In_354);
nand U1801 (N_1801,In_959,In_1160);
and U1802 (N_1802,In_671,In_584);
nor U1803 (N_1803,In_408,In_825);
nand U1804 (N_1804,In_915,In_744);
nor U1805 (N_1805,In_1305,In_924);
nor U1806 (N_1806,In_1384,In_1380);
nor U1807 (N_1807,In_598,In_125);
and U1808 (N_1808,In_902,In_342);
or U1809 (N_1809,In_1253,In_1310);
or U1810 (N_1810,In_1182,In_266);
and U1811 (N_1811,In_723,In_911);
nand U1812 (N_1812,In_1491,In_870);
nand U1813 (N_1813,In_181,In_48);
nand U1814 (N_1814,In_96,In_1447);
nand U1815 (N_1815,In_1182,In_734);
nor U1816 (N_1816,In_437,In_230);
or U1817 (N_1817,In_197,In_132);
and U1818 (N_1818,In_86,In_406);
or U1819 (N_1819,In_517,In_1349);
nand U1820 (N_1820,In_166,In_157);
or U1821 (N_1821,In_647,In_669);
nor U1822 (N_1822,In_431,In_115);
or U1823 (N_1823,In_1223,In_524);
nor U1824 (N_1824,In_1087,In_344);
nand U1825 (N_1825,In_906,In_192);
or U1826 (N_1826,In_499,In_138);
nor U1827 (N_1827,In_409,In_1152);
or U1828 (N_1828,In_1384,In_1028);
and U1829 (N_1829,In_1249,In_436);
and U1830 (N_1830,In_811,In_788);
or U1831 (N_1831,In_1212,In_995);
and U1832 (N_1832,In_471,In_1193);
nand U1833 (N_1833,In_824,In_887);
and U1834 (N_1834,In_761,In_424);
nor U1835 (N_1835,In_264,In_412);
or U1836 (N_1836,In_252,In_919);
and U1837 (N_1837,In_1344,In_568);
or U1838 (N_1838,In_390,In_1073);
nor U1839 (N_1839,In_1062,In_291);
or U1840 (N_1840,In_358,In_1255);
nor U1841 (N_1841,In_1317,In_1402);
nor U1842 (N_1842,In_458,In_333);
and U1843 (N_1843,In_677,In_172);
and U1844 (N_1844,In_1270,In_1302);
nor U1845 (N_1845,In_800,In_1360);
and U1846 (N_1846,In_714,In_796);
nor U1847 (N_1847,In_1104,In_1037);
nand U1848 (N_1848,In_725,In_1337);
nand U1849 (N_1849,In_291,In_121);
nand U1850 (N_1850,In_1471,In_1046);
and U1851 (N_1851,In_1133,In_835);
or U1852 (N_1852,In_1328,In_312);
or U1853 (N_1853,In_775,In_1044);
nor U1854 (N_1854,In_1462,In_1006);
nand U1855 (N_1855,In_441,In_308);
nand U1856 (N_1856,In_1336,In_1059);
nor U1857 (N_1857,In_1096,In_1380);
and U1858 (N_1858,In_41,In_738);
and U1859 (N_1859,In_591,In_428);
and U1860 (N_1860,In_1069,In_559);
nand U1861 (N_1861,In_941,In_1454);
nand U1862 (N_1862,In_863,In_1330);
nand U1863 (N_1863,In_793,In_194);
and U1864 (N_1864,In_1376,In_516);
nand U1865 (N_1865,In_1143,In_54);
or U1866 (N_1866,In_153,In_1445);
nand U1867 (N_1867,In_802,In_559);
nand U1868 (N_1868,In_936,In_897);
and U1869 (N_1869,In_711,In_820);
nor U1870 (N_1870,In_21,In_873);
nor U1871 (N_1871,In_1096,In_959);
and U1872 (N_1872,In_1043,In_1367);
and U1873 (N_1873,In_127,In_1055);
nor U1874 (N_1874,In_251,In_137);
nor U1875 (N_1875,In_222,In_1437);
nand U1876 (N_1876,In_783,In_432);
or U1877 (N_1877,In_490,In_1185);
nor U1878 (N_1878,In_1360,In_1123);
nor U1879 (N_1879,In_904,In_128);
nor U1880 (N_1880,In_1491,In_623);
or U1881 (N_1881,In_282,In_99);
nand U1882 (N_1882,In_840,In_833);
and U1883 (N_1883,In_110,In_89);
nor U1884 (N_1884,In_1089,In_790);
nand U1885 (N_1885,In_244,In_178);
and U1886 (N_1886,In_1381,In_1161);
nand U1887 (N_1887,In_220,In_269);
or U1888 (N_1888,In_524,In_1154);
nand U1889 (N_1889,In_944,In_1426);
and U1890 (N_1890,In_357,In_1494);
nor U1891 (N_1891,In_1428,In_891);
and U1892 (N_1892,In_966,In_1087);
nor U1893 (N_1893,In_802,In_1090);
nor U1894 (N_1894,In_620,In_679);
nand U1895 (N_1895,In_790,In_585);
nand U1896 (N_1896,In_1412,In_1032);
and U1897 (N_1897,In_1395,In_1438);
or U1898 (N_1898,In_1255,In_646);
and U1899 (N_1899,In_1230,In_351);
nor U1900 (N_1900,In_1351,In_1181);
or U1901 (N_1901,In_171,In_60);
or U1902 (N_1902,In_474,In_1202);
nor U1903 (N_1903,In_1048,In_1201);
or U1904 (N_1904,In_1320,In_32);
nand U1905 (N_1905,In_579,In_123);
and U1906 (N_1906,In_849,In_927);
nor U1907 (N_1907,In_759,In_737);
nor U1908 (N_1908,In_121,In_655);
nand U1909 (N_1909,In_601,In_1464);
and U1910 (N_1910,In_331,In_89);
nand U1911 (N_1911,In_888,In_127);
or U1912 (N_1912,In_1356,In_136);
or U1913 (N_1913,In_57,In_1387);
and U1914 (N_1914,In_812,In_1112);
nand U1915 (N_1915,In_963,In_616);
and U1916 (N_1916,In_21,In_620);
nand U1917 (N_1917,In_1287,In_742);
or U1918 (N_1918,In_830,In_1323);
nand U1919 (N_1919,In_1234,In_1452);
xnor U1920 (N_1920,In_723,In_491);
or U1921 (N_1921,In_781,In_1446);
nor U1922 (N_1922,In_66,In_882);
and U1923 (N_1923,In_531,In_1219);
nor U1924 (N_1924,In_20,In_121);
and U1925 (N_1925,In_510,In_972);
and U1926 (N_1926,In_1133,In_166);
nor U1927 (N_1927,In_530,In_1038);
nor U1928 (N_1928,In_632,In_601);
and U1929 (N_1929,In_1269,In_23);
nand U1930 (N_1930,In_1300,In_510);
nor U1931 (N_1931,In_1105,In_1302);
and U1932 (N_1932,In_339,In_867);
or U1933 (N_1933,In_1215,In_389);
nor U1934 (N_1934,In_1488,In_409);
nor U1935 (N_1935,In_1272,In_479);
nor U1936 (N_1936,In_103,In_1248);
and U1937 (N_1937,In_583,In_1036);
nand U1938 (N_1938,In_920,In_1292);
or U1939 (N_1939,In_953,In_44);
and U1940 (N_1940,In_1460,In_287);
and U1941 (N_1941,In_49,In_230);
xnor U1942 (N_1942,In_50,In_222);
nand U1943 (N_1943,In_995,In_1041);
nor U1944 (N_1944,In_1123,In_850);
nor U1945 (N_1945,In_1477,In_995);
or U1946 (N_1946,In_1034,In_1332);
nand U1947 (N_1947,In_1170,In_1267);
or U1948 (N_1948,In_114,In_196);
nor U1949 (N_1949,In_492,In_1176);
and U1950 (N_1950,In_1008,In_417);
xnor U1951 (N_1951,In_445,In_605);
nor U1952 (N_1952,In_1251,In_93);
nand U1953 (N_1953,In_277,In_1192);
nor U1954 (N_1954,In_740,In_702);
nor U1955 (N_1955,In_146,In_568);
or U1956 (N_1956,In_604,In_359);
nor U1957 (N_1957,In_946,In_470);
nand U1958 (N_1958,In_638,In_1415);
nor U1959 (N_1959,In_535,In_793);
or U1960 (N_1960,In_370,In_766);
and U1961 (N_1961,In_736,In_1055);
nor U1962 (N_1962,In_954,In_372);
or U1963 (N_1963,In_1458,In_531);
and U1964 (N_1964,In_1355,In_1149);
and U1965 (N_1965,In_396,In_516);
nand U1966 (N_1966,In_1163,In_1283);
or U1967 (N_1967,In_953,In_357);
or U1968 (N_1968,In_442,In_250);
and U1969 (N_1969,In_608,In_1290);
nor U1970 (N_1970,In_136,In_40);
nor U1971 (N_1971,In_111,In_1150);
nor U1972 (N_1972,In_621,In_428);
or U1973 (N_1973,In_1095,In_846);
and U1974 (N_1974,In_1172,In_1286);
or U1975 (N_1975,In_133,In_1254);
nor U1976 (N_1976,In_193,In_685);
nor U1977 (N_1977,In_358,In_735);
and U1978 (N_1978,In_262,In_304);
nand U1979 (N_1979,In_813,In_1065);
nand U1980 (N_1980,In_835,In_650);
and U1981 (N_1981,In_590,In_1081);
and U1982 (N_1982,In_1474,In_756);
nor U1983 (N_1983,In_760,In_1223);
nor U1984 (N_1984,In_716,In_221);
nor U1985 (N_1985,In_352,In_906);
nor U1986 (N_1986,In_294,In_1271);
nor U1987 (N_1987,In_958,In_1145);
or U1988 (N_1988,In_946,In_831);
nor U1989 (N_1989,In_85,In_947);
nor U1990 (N_1990,In_1234,In_667);
and U1991 (N_1991,In_339,In_1421);
nor U1992 (N_1992,In_340,In_915);
or U1993 (N_1993,In_127,In_117);
and U1994 (N_1994,In_601,In_1185);
nor U1995 (N_1995,In_1100,In_632);
nand U1996 (N_1996,In_1078,In_1497);
and U1997 (N_1997,In_688,In_194);
and U1998 (N_1998,In_259,In_261);
and U1999 (N_1999,In_440,In_1134);
nand U2000 (N_2000,In_1183,In_774);
nor U2001 (N_2001,In_1465,In_1245);
or U2002 (N_2002,In_717,In_574);
nor U2003 (N_2003,In_86,In_769);
or U2004 (N_2004,In_1086,In_627);
or U2005 (N_2005,In_1123,In_753);
nor U2006 (N_2006,In_1277,In_967);
nand U2007 (N_2007,In_752,In_1086);
nand U2008 (N_2008,In_457,In_597);
xor U2009 (N_2009,In_1100,In_7);
and U2010 (N_2010,In_400,In_157);
or U2011 (N_2011,In_1203,In_58);
and U2012 (N_2012,In_928,In_429);
nand U2013 (N_2013,In_1297,In_437);
or U2014 (N_2014,In_484,In_172);
and U2015 (N_2015,In_747,In_1497);
nand U2016 (N_2016,In_351,In_1375);
and U2017 (N_2017,In_1249,In_101);
or U2018 (N_2018,In_964,In_1080);
nor U2019 (N_2019,In_150,In_1232);
nand U2020 (N_2020,In_1357,In_473);
and U2021 (N_2021,In_617,In_1046);
nand U2022 (N_2022,In_1396,In_59);
nand U2023 (N_2023,In_19,In_594);
or U2024 (N_2024,In_1395,In_35);
and U2025 (N_2025,In_1161,In_704);
nand U2026 (N_2026,In_535,In_818);
nand U2027 (N_2027,In_556,In_199);
nor U2028 (N_2028,In_1123,In_188);
nor U2029 (N_2029,In_801,In_541);
nor U2030 (N_2030,In_1209,In_1425);
and U2031 (N_2031,In_766,In_652);
and U2032 (N_2032,In_47,In_1305);
or U2033 (N_2033,In_983,In_1138);
nor U2034 (N_2034,In_984,In_698);
nor U2035 (N_2035,In_343,In_16);
and U2036 (N_2036,In_500,In_1114);
nand U2037 (N_2037,In_1438,In_1379);
or U2038 (N_2038,In_198,In_938);
nand U2039 (N_2039,In_1033,In_759);
nand U2040 (N_2040,In_1141,In_15);
or U2041 (N_2041,In_1316,In_1429);
and U2042 (N_2042,In_1432,In_1445);
nor U2043 (N_2043,In_791,In_1055);
and U2044 (N_2044,In_448,In_587);
nand U2045 (N_2045,In_1036,In_327);
and U2046 (N_2046,In_213,In_101);
nand U2047 (N_2047,In_81,In_1156);
nand U2048 (N_2048,In_1057,In_415);
nor U2049 (N_2049,In_709,In_1216);
and U2050 (N_2050,In_518,In_787);
and U2051 (N_2051,In_1017,In_1294);
or U2052 (N_2052,In_876,In_572);
nor U2053 (N_2053,In_899,In_1145);
nor U2054 (N_2054,In_747,In_695);
and U2055 (N_2055,In_803,In_189);
and U2056 (N_2056,In_1195,In_1097);
or U2057 (N_2057,In_907,In_1046);
or U2058 (N_2058,In_1234,In_298);
and U2059 (N_2059,In_910,In_231);
or U2060 (N_2060,In_1042,In_1033);
and U2061 (N_2061,In_555,In_458);
or U2062 (N_2062,In_909,In_727);
nand U2063 (N_2063,In_1167,In_176);
or U2064 (N_2064,In_918,In_1451);
nor U2065 (N_2065,In_738,In_586);
and U2066 (N_2066,In_1227,In_819);
or U2067 (N_2067,In_1375,In_1172);
or U2068 (N_2068,In_990,In_1229);
or U2069 (N_2069,In_222,In_1235);
nor U2070 (N_2070,In_1465,In_1234);
nand U2071 (N_2071,In_1190,In_1356);
or U2072 (N_2072,In_575,In_1063);
and U2073 (N_2073,In_357,In_456);
nor U2074 (N_2074,In_1000,In_1176);
or U2075 (N_2075,In_847,In_443);
or U2076 (N_2076,In_1226,In_412);
and U2077 (N_2077,In_584,In_949);
nand U2078 (N_2078,In_201,In_168);
and U2079 (N_2079,In_768,In_688);
or U2080 (N_2080,In_206,In_120);
nor U2081 (N_2081,In_84,In_97);
or U2082 (N_2082,In_792,In_689);
nand U2083 (N_2083,In_891,In_508);
and U2084 (N_2084,In_1465,In_591);
xnor U2085 (N_2085,In_249,In_969);
and U2086 (N_2086,In_343,In_1017);
and U2087 (N_2087,In_1259,In_976);
nor U2088 (N_2088,In_132,In_1339);
or U2089 (N_2089,In_1116,In_1170);
and U2090 (N_2090,In_575,In_848);
and U2091 (N_2091,In_642,In_1224);
or U2092 (N_2092,In_512,In_1486);
and U2093 (N_2093,In_829,In_170);
and U2094 (N_2094,In_726,In_381);
nand U2095 (N_2095,In_676,In_451);
or U2096 (N_2096,In_298,In_625);
and U2097 (N_2097,In_1246,In_1186);
or U2098 (N_2098,In_1070,In_28);
nand U2099 (N_2099,In_596,In_419);
or U2100 (N_2100,In_270,In_87);
or U2101 (N_2101,In_44,In_458);
and U2102 (N_2102,In_1401,In_1223);
and U2103 (N_2103,In_1233,In_1442);
nand U2104 (N_2104,In_829,In_399);
or U2105 (N_2105,In_34,In_1364);
or U2106 (N_2106,In_989,In_711);
xnor U2107 (N_2107,In_71,In_795);
nand U2108 (N_2108,In_1004,In_591);
or U2109 (N_2109,In_1152,In_871);
and U2110 (N_2110,In_1449,In_736);
nor U2111 (N_2111,In_1495,In_7);
nor U2112 (N_2112,In_1158,In_1175);
or U2113 (N_2113,In_1392,In_761);
nor U2114 (N_2114,In_93,In_851);
nor U2115 (N_2115,In_639,In_1358);
nor U2116 (N_2116,In_1408,In_951);
or U2117 (N_2117,In_774,In_1338);
nand U2118 (N_2118,In_1413,In_700);
nor U2119 (N_2119,In_244,In_364);
nor U2120 (N_2120,In_1114,In_986);
and U2121 (N_2121,In_1332,In_268);
and U2122 (N_2122,In_1409,In_82);
and U2123 (N_2123,In_36,In_561);
nor U2124 (N_2124,In_848,In_790);
or U2125 (N_2125,In_795,In_1092);
nor U2126 (N_2126,In_10,In_1105);
nand U2127 (N_2127,In_1023,In_385);
nor U2128 (N_2128,In_186,In_152);
and U2129 (N_2129,In_321,In_8);
and U2130 (N_2130,In_392,In_652);
nor U2131 (N_2131,In_116,In_863);
and U2132 (N_2132,In_586,In_1391);
nand U2133 (N_2133,In_170,In_490);
or U2134 (N_2134,In_913,In_724);
and U2135 (N_2135,In_1075,In_1262);
and U2136 (N_2136,In_1342,In_884);
and U2137 (N_2137,In_415,In_1150);
and U2138 (N_2138,In_688,In_469);
nand U2139 (N_2139,In_1428,In_1104);
nor U2140 (N_2140,In_957,In_822);
nand U2141 (N_2141,In_1043,In_811);
and U2142 (N_2142,In_805,In_390);
or U2143 (N_2143,In_721,In_1131);
or U2144 (N_2144,In_430,In_1419);
nand U2145 (N_2145,In_926,In_632);
or U2146 (N_2146,In_1139,In_468);
nand U2147 (N_2147,In_71,In_957);
or U2148 (N_2148,In_947,In_22);
and U2149 (N_2149,In_1036,In_612);
nor U2150 (N_2150,In_569,In_696);
or U2151 (N_2151,In_122,In_444);
and U2152 (N_2152,In_568,In_1394);
nor U2153 (N_2153,In_1399,In_645);
and U2154 (N_2154,In_834,In_632);
and U2155 (N_2155,In_1320,In_902);
nor U2156 (N_2156,In_1104,In_745);
or U2157 (N_2157,In_1204,In_121);
nor U2158 (N_2158,In_1399,In_987);
nand U2159 (N_2159,In_744,In_945);
nor U2160 (N_2160,In_1466,In_1030);
nor U2161 (N_2161,In_855,In_956);
nand U2162 (N_2162,In_1423,In_1497);
nor U2163 (N_2163,In_1241,In_1073);
and U2164 (N_2164,In_378,In_1175);
or U2165 (N_2165,In_729,In_822);
nor U2166 (N_2166,In_803,In_1338);
nand U2167 (N_2167,In_447,In_682);
nand U2168 (N_2168,In_769,In_627);
and U2169 (N_2169,In_748,In_688);
nor U2170 (N_2170,In_444,In_1093);
and U2171 (N_2171,In_1120,In_848);
nor U2172 (N_2172,In_862,In_860);
nor U2173 (N_2173,In_699,In_1129);
or U2174 (N_2174,In_664,In_485);
nand U2175 (N_2175,In_987,In_278);
or U2176 (N_2176,In_1130,In_127);
and U2177 (N_2177,In_1148,In_1206);
or U2178 (N_2178,In_1325,In_29);
and U2179 (N_2179,In_22,In_313);
nor U2180 (N_2180,In_156,In_1417);
nor U2181 (N_2181,In_112,In_771);
or U2182 (N_2182,In_1364,In_638);
or U2183 (N_2183,In_1100,In_402);
or U2184 (N_2184,In_1144,In_140);
nand U2185 (N_2185,In_862,In_1114);
nor U2186 (N_2186,In_353,In_78);
and U2187 (N_2187,In_984,In_918);
xor U2188 (N_2188,In_1048,In_646);
or U2189 (N_2189,In_1086,In_1351);
nor U2190 (N_2190,In_698,In_1333);
or U2191 (N_2191,In_499,In_647);
nand U2192 (N_2192,In_953,In_367);
nor U2193 (N_2193,In_220,In_1027);
nor U2194 (N_2194,In_1362,In_299);
and U2195 (N_2195,In_1218,In_1234);
and U2196 (N_2196,In_517,In_1415);
nand U2197 (N_2197,In_972,In_339);
and U2198 (N_2198,In_848,In_556);
nand U2199 (N_2199,In_834,In_615);
nor U2200 (N_2200,In_1094,In_566);
or U2201 (N_2201,In_432,In_26);
nor U2202 (N_2202,In_1440,In_1012);
and U2203 (N_2203,In_1120,In_637);
or U2204 (N_2204,In_49,In_683);
and U2205 (N_2205,In_270,In_472);
or U2206 (N_2206,In_123,In_181);
nand U2207 (N_2207,In_514,In_1087);
or U2208 (N_2208,In_1344,In_815);
and U2209 (N_2209,In_509,In_365);
and U2210 (N_2210,In_89,In_1454);
and U2211 (N_2211,In_231,In_473);
or U2212 (N_2212,In_1086,In_553);
or U2213 (N_2213,In_507,In_989);
and U2214 (N_2214,In_327,In_745);
nand U2215 (N_2215,In_83,In_403);
and U2216 (N_2216,In_1098,In_1391);
and U2217 (N_2217,In_1257,In_1170);
nor U2218 (N_2218,In_431,In_492);
nand U2219 (N_2219,In_1436,In_113);
or U2220 (N_2220,In_41,In_1213);
nor U2221 (N_2221,In_696,In_970);
and U2222 (N_2222,In_826,In_481);
nand U2223 (N_2223,In_864,In_216);
nor U2224 (N_2224,In_313,In_13);
nor U2225 (N_2225,In_537,In_1054);
or U2226 (N_2226,In_1197,In_818);
nor U2227 (N_2227,In_236,In_1270);
nand U2228 (N_2228,In_1396,In_770);
nor U2229 (N_2229,In_778,In_1303);
nor U2230 (N_2230,In_972,In_52);
nor U2231 (N_2231,In_1063,In_112);
xnor U2232 (N_2232,In_1476,In_1331);
or U2233 (N_2233,In_1235,In_517);
and U2234 (N_2234,In_962,In_898);
and U2235 (N_2235,In_1022,In_351);
nor U2236 (N_2236,In_443,In_921);
nand U2237 (N_2237,In_705,In_313);
nor U2238 (N_2238,In_893,In_1043);
or U2239 (N_2239,In_1327,In_91);
nand U2240 (N_2240,In_874,In_749);
nand U2241 (N_2241,In_1048,In_256);
or U2242 (N_2242,In_1181,In_932);
or U2243 (N_2243,In_72,In_1392);
or U2244 (N_2244,In_381,In_243);
and U2245 (N_2245,In_671,In_1036);
nand U2246 (N_2246,In_597,In_1089);
and U2247 (N_2247,In_515,In_1035);
nor U2248 (N_2248,In_7,In_1195);
nor U2249 (N_2249,In_923,In_1310);
nor U2250 (N_2250,In_402,In_801);
and U2251 (N_2251,In_537,In_432);
nor U2252 (N_2252,In_1390,In_535);
or U2253 (N_2253,In_1204,In_665);
and U2254 (N_2254,In_460,In_986);
or U2255 (N_2255,In_1249,In_471);
and U2256 (N_2256,In_921,In_413);
or U2257 (N_2257,In_1447,In_107);
or U2258 (N_2258,In_1446,In_1179);
nand U2259 (N_2259,In_1402,In_255);
and U2260 (N_2260,In_251,In_365);
and U2261 (N_2261,In_711,In_1398);
nor U2262 (N_2262,In_592,In_721);
and U2263 (N_2263,In_721,In_1228);
nand U2264 (N_2264,In_860,In_886);
nor U2265 (N_2265,In_406,In_1384);
nand U2266 (N_2266,In_830,In_664);
or U2267 (N_2267,In_853,In_989);
nand U2268 (N_2268,In_328,In_278);
and U2269 (N_2269,In_1050,In_570);
nor U2270 (N_2270,In_1222,In_977);
nand U2271 (N_2271,In_689,In_1335);
and U2272 (N_2272,In_175,In_936);
or U2273 (N_2273,In_548,In_45);
and U2274 (N_2274,In_752,In_524);
or U2275 (N_2275,In_1285,In_971);
and U2276 (N_2276,In_267,In_772);
and U2277 (N_2277,In_1378,In_581);
nand U2278 (N_2278,In_1499,In_734);
nor U2279 (N_2279,In_504,In_675);
or U2280 (N_2280,In_863,In_934);
nand U2281 (N_2281,In_1450,In_630);
xor U2282 (N_2282,In_1262,In_745);
and U2283 (N_2283,In_455,In_513);
nor U2284 (N_2284,In_959,In_305);
nor U2285 (N_2285,In_1154,In_422);
and U2286 (N_2286,In_123,In_1115);
and U2287 (N_2287,In_757,In_664);
or U2288 (N_2288,In_458,In_394);
or U2289 (N_2289,In_586,In_868);
nand U2290 (N_2290,In_1030,In_1209);
or U2291 (N_2291,In_873,In_1416);
nand U2292 (N_2292,In_36,In_729);
nor U2293 (N_2293,In_74,In_1360);
or U2294 (N_2294,In_112,In_1097);
nand U2295 (N_2295,In_1452,In_260);
or U2296 (N_2296,In_1050,In_726);
nor U2297 (N_2297,In_1407,In_1281);
nand U2298 (N_2298,In_691,In_91);
nor U2299 (N_2299,In_656,In_1394);
or U2300 (N_2300,In_743,In_919);
and U2301 (N_2301,In_611,In_1490);
nor U2302 (N_2302,In_1390,In_658);
or U2303 (N_2303,In_1247,In_1005);
nor U2304 (N_2304,In_924,In_1113);
and U2305 (N_2305,In_1426,In_1031);
nor U2306 (N_2306,In_1480,In_520);
nor U2307 (N_2307,In_1072,In_190);
nor U2308 (N_2308,In_939,In_311);
and U2309 (N_2309,In_1485,In_1173);
and U2310 (N_2310,In_629,In_639);
nor U2311 (N_2311,In_1173,In_1034);
nand U2312 (N_2312,In_1449,In_1046);
nand U2313 (N_2313,In_502,In_674);
nor U2314 (N_2314,In_899,In_967);
xnor U2315 (N_2315,In_347,In_1167);
nand U2316 (N_2316,In_50,In_534);
nand U2317 (N_2317,In_1339,In_0);
nor U2318 (N_2318,In_444,In_1367);
or U2319 (N_2319,In_309,In_15);
nor U2320 (N_2320,In_1304,In_1232);
nor U2321 (N_2321,In_78,In_1009);
and U2322 (N_2322,In_234,In_1410);
and U2323 (N_2323,In_734,In_288);
nor U2324 (N_2324,In_92,In_1357);
nand U2325 (N_2325,In_823,In_936);
or U2326 (N_2326,In_645,In_186);
and U2327 (N_2327,In_702,In_522);
nor U2328 (N_2328,In_5,In_479);
nand U2329 (N_2329,In_1400,In_261);
nor U2330 (N_2330,In_901,In_516);
or U2331 (N_2331,In_1397,In_656);
or U2332 (N_2332,In_521,In_1040);
or U2333 (N_2333,In_130,In_584);
xnor U2334 (N_2334,In_1360,In_919);
nand U2335 (N_2335,In_47,In_888);
or U2336 (N_2336,In_525,In_9);
or U2337 (N_2337,In_338,In_1142);
or U2338 (N_2338,In_580,In_441);
or U2339 (N_2339,In_535,In_69);
nor U2340 (N_2340,In_434,In_703);
nand U2341 (N_2341,In_1391,In_1420);
or U2342 (N_2342,In_217,In_1010);
or U2343 (N_2343,In_132,In_719);
or U2344 (N_2344,In_1142,In_349);
nor U2345 (N_2345,In_1173,In_1175);
or U2346 (N_2346,In_1274,In_709);
and U2347 (N_2347,In_964,In_1273);
and U2348 (N_2348,In_838,In_853);
nor U2349 (N_2349,In_293,In_1172);
nor U2350 (N_2350,In_1270,In_986);
nand U2351 (N_2351,In_845,In_264);
nor U2352 (N_2352,In_585,In_57);
and U2353 (N_2353,In_1446,In_626);
and U2354 (N_2354,In_1101,In_967);
nor U2355 (N_2355,In_1496,In_1444);
or U2356 (N_2356,In_244,In_1323);
nor U2357 (N_2357,In_864,In_1385);
nor U2358 (N_2358,In_1444,In_477);
or U2359 (N_2359,In_345,In_1378);
xor U2360 (N_2360,In_980,In_1130);
nor U2361 (N_2361,In_534,In_44);
and U2362 (N_2362,In_618,In_1209);
nand U2363 (N_2363,In_815,In_272);
nor U2364 (N_2364,In_799,In_750);
or U2365 (N_2365,In_689,In_833);
nand U2366 (N_2366,In_1018,In_788);
and U2367 (N_2367,In_1496,In_336);
or U2368 (N_2368,In_291,In_838);
or U2369 (N_2369,In_1083,In_1406);
and U2370 (N_2370,In_872,In_93);
nand U2371 (N_2371,In_514,In_110);
or U2372 (N_2372,In_1313,In_332);
nor U2373 (N_2373,In_767,In_980);
or U2374 (N_2374,In_318,In_242);
and U2375 (N_2375,In_1308,In_1216);
or U2376 (N_2376,In_168,In_268);
nor U2377 (N_2377,In_1098,In_342);
or U2378 (N_2378,In_980,In_499);
nor U2379 (N_2379,In_134,In_959);
nor U2380 (N_2380,In_425,In_102);
and U2381 (N_2381,In_150,In_161);
xnor U2382 (N_2382,In_1236,In_1449);
nor U2383 (N_2383,In_291,In_7);
nor U2384 (N_2384,In_179,In_1144);
and U2385 (N_2385,In_99,In_646);
or U2386 (N_2386,In_1163,In_643);
or U2387 (N_2387,In_1231,In_1253);
nor U2388 (N_2388,In_1011,In_670);
nor U2389 (N_2389,In_362,In_1211);
nor U2390 (N_2390,In_641,In_1295);
or U2391 (N_2391,In_1022,In_974);
and U2392 (N_2392,In_8,In_1103);
and U2393 (N_2393,In_1280,In_201);
or U2394 (N_2394,In_426,In_552);
and U2395 (N_2395,In_580,In_996);
nand U2396 (N_2396,In_627,In_1263);
nand U2397 (N_2397,In_735,In_814);
nand U2398 (N_2398,In_1206,In_438);
nor U2399 (N_2399,In_158,In_1145);
nor U2400 (N_2400,In_609,In_667);
nand U2401 (N_2401,In_104,In_1212);
nand U2402 (N_2402,In_886,In_236);
or U2403 (N_2403,In_628,In_560);
or U2404 (N_2404,In_536,In_1194);
nor U2405 (N_2405,In_1404,In_1138);
nor U2406 (N_2406,In_646,In_304);
and U2407 (N_2407,In_1361,In_662);
nor U2408 (N_2408,In_528,In_849);
nand U2409 (N_2409,In_1256,In_288);
nand U2410 (N_2410,In_1065,In_165);
nor U2411 (N_2411,In_877,In_895);
and U2412 (N_2412,In_153,In_954);
nor U2413 (N_2413,In_1236,In_546);
or U2414 (N_2414,In_487,In_406);
nor U2415 (N_2415,In_225,In_1048);
nor U2416 (N_2416,In_62,In_567);
nand U2417 (N_2417,In_60,In_975);
and U2418 (N_2418,In_88,In_615);
nor U2419 (N_2419,In_1311,In_1192);
and U2420 (N_2420,In_159,In_472);
nor U2421 (N_2421,In_639,In_213);
nor U2422 (N_2422,In_700,In_910);
nor U2423 (N_2423,In_1041,In_526);
nand U2424 (N_2424,In_935,In_644);
nand U2425 (N_2425,In_848,In_264);
nor U2426 (N_2426,In_1488,In_690);
nand U2427 (N_2427,In_868,In_838);
and U2428 (N_2428,In_66,In_256);
nor U2429 (N_2429,In_298,In_1010);
and U2430 (N_2430,In_1108,In_114);
nor U2431 (N_2431,In_815,In_330);
nand U2432 (N_2432,In_396,In_562);
nor U2433 (N_2433,In_978,In_608);
or U2434 (N_2434,In_6,In_236);
nor U2435 (N_2435,In_1139,In_748);
and U2436 (N_2436,In_719,In_1020);
or U2437 (N_2437,In_134,In_1358);
nand U2438 (N_2438,In_680,In_98);
nand U2439 (N_2439,In_1095,In_997);
nor U2440 (N_2440,In_1346,In_995);
or U2441 (N_2441,In_63,In_1448);
and U2442 (N_2442,In_1090,In_759);
nor U2443 (N_2443,In_1103,In_1445);
nor U2444 (N_2444,In_874,In_492);
nor U2445 (N_2445,In_302,In_1227);
nor U2446 (N_2446,In_904,In_120);
and U2447 (N_2447,In_488,In_956);
nand U2448 (N_2448,In_482,In_1244);
and U2449 (N_2449,In_562,In_1221);
and U2450 (N_2450,In_15,In_1423);
and U2451 (N_2451,In_155,In_841);
nand U2452 (N_2452,In_688,In_1201);
and U2453 (N_2453,In_1252,In_854);
nand U2454 (N_2454,In_365,In_689);
nor U2455 (N_2455,In_278,In_1062);
nand U2456 (N_2456,In_1458,In_379);
xnor U2457 (N_2457,In_1389,In_992);
and U2458 (N_2458,In_946,In_354);
or U2459 (N_2459,In_865,In_1296);
nor U2460 (N_2460,In_64,In_950);
nand U2461 (N_2461,In_164,In_1160);
nor U2462 (N_2462,In_1168,In_943);
and U2463 (N_2463,In_147,In_869);
or U2464 (N_2464,In_469,In_1275);
or U2465 (N_2465,In_65,In_985);
nor U2466 (N_2466,In_1178,In_1257);
or U2467 (N_2467,In_871,In_327);
nor U2468 (N_2468,In_295,In_719);
nor U2469 (N_2469,In_588,In_1049);
nor U2470 (N_2470,In_536,In_1099);
nor U2471 (N_2471,In_1414,In_512);
or U2472 (N_2472,In_777,In_900);
nand U2473 (N_2473,In_878,In_331);
or U2474 (N_2474,In_221,In_260);
nor U2475 (N_2475,In_1345,In_802);
nand U2476 (N_2476,In_860,In_507);
nand U2477 (N_2477,In_1138,In_535);
or U2478 (N_2478,In_316,In_697);
nand U2479 (N_2479,In_922,In_1444);
nand U2480 (N_2480,In_462,In_551);
nand U2481 (N_2481,In_787,In_914);
nor U2482 (N_2482,In_670,In_106);
and U2483 (N_2483,In_766,In_125);
nor U2484 (N_2484,In_1366,In_869);
or U2485 (N_2485,In_154,In_692);
or U2486 (N_2486,In_1039,In_1212);
and U2487 (N_2487,In_1180,In_1261);
nor U2488 (N_2488,In_1384,In_170);
nor U2489 (N_2489,In_682,In_912);
and U2490 (N_2490,In_1037,In_185);
and U2491 (N_2491,In_783,In_1125);
and U2492 (N_2492,In_348,In_533);
nor U2493 (N_2493,In_801,In_649);
and U2494 (N_2494,In_1355,In_1323);
nand U2495 (N_2495,In_752,In_1489);
or U2496 (N_2496,In_1163,In_1038);
and U2497 (N_2497,In_745,In_440);
nor U2498 (N_2498,In_504,In_1312);
and U2499 (N_2499,In_566,In_98);
or U2500 (N_2500,In_538,In_1175);
nand U2501 (N_2501,In_901,In_372);
or U2502 (N_2502,In_782,In_255);
or U2503 (N_2503,In_441,In_626);
nor U2504 (N_2504,In_719,In_1313);
or U2505 (N_2505,In_1450,In_1319);
and U2506 (N_2506,In_756,In_897);
nor U2507 (N_2507,In_346,In_1258);
and U2508 (N_2508,In_1348,In_1078);
nor U2509 (N_2509,In_1034,In_1202);
and U2510 (N_2510,In_210,In_389);
nand U2511 (N_2511,In_1231,In_1084);
or U2512 (N_2512,In_1348,In_1417);
or U2513 (N_2513,In_432,In_1096);
nand U2514 (N_2514,In_295,In_440);
nand U2515 (N_2515,In_229,In_726);
nor U2516 (N_2516,In_999,In_598);
or U2517 (N_2517,In_1177,In_765);
nor U2518 (N_2518,In_1216,In_642);
nor U2519 (N_2519,In_1422,In_229);
or U2520 (N_2520,In_507,In_985);
or U2521 (N_2521,In_1327,In_863);
and U2522 (N_2522,In_690,In_90);
or U2523 (N_2523,In_830,In_811);
and U2524 (N_2524,In_475,In_602);
and U2525 (N_2525,In_417,In_57);
and U2526 (N_2526,In_1317,In_1076);
nor U2527 (N_2527,In_988,In_1429);
nand U2528 (N_2528,In_898,In_600);
nor U2529 (N_2529,In_931,In_949);
nand U2530 (N_2530,In_1412,In_437);
nand U2531 (N_2531,In_1493,In_566);
nand U2532 (N_2532,In_678,In_380);
or U2533 (N_2533,In_354,In_73);
nor U2534 (N_2534,In_33,In_191);
nand U2535 (N_2535,In_444,In_527);
and U2536 (N_2536,In_673,In_744);
and U2537 (N_2537,In_935,In_905);
nor U2538 (N_2538,In_749,In_1286);
and U2539 (N_2539,In_247,In_81);
or U2540 (N_2540,In_1231,In_788);
nor U2541 (N_2541,In_229,In_46);
or U2542 (N_2542,In_404,In_1480);
nor U2543 (N_2543,In_517,In_324);
xnor U2544 (N_2544,In_1451,In_789);
nand U2545 (N_2545,In_560,In_289);
nor U2546 (N_2546,In_1230,In_1318);
and U2547 (N_2547,In_157,In_530);
nand U2548 (N_2548,In_159,In_156);
and U2549 (N_2549,In_1351,In_1037);
nor U2550 (N_2550,In_91,In_269);
nand U2551 (N_2551,In_726,In_1123);
nor U2552 (N_2552,In_539,In_1441);
nor U2553 (N_2553,In_263,In_1270);
nor U2554 (N_2554,In_823,In_669);
and U2555 (N_2555,In_28,In_1433);
or U2556 (N_2556,In_1379,In_985);
and U2557 (N_2557,In_1188,In_567);
and U2558 (N_2558,In_513,In_1456);
nand U2559 (N_2559,In_167,In_252);
nand U2560 (N_2560,In_739,In_1324);
nor U2561 (N_2561,In_113,In_1238);
and U2562 (N_2562,In_1480,In_1194);
or U2563 (N_2563,In_340,In_1461);
nand U2564 (N_2564,In_214,In_434);
nand U2565 (N_2565,In_242,In_897);
nor U2566 (N_2566,In_285,In_1052);
or U2567 (N_2567,In_75,In_603);
nand U2568 (N_2568,In_489,In_1016);
or U2569 (N_2569,In_1119,In_354);
nor U2570 (N_2570,In_385,In_399);
nor U2571 (N_2571,In_133,In_1433);
or U2572 (N_2572,In_406,In_1269);
nor U2573 (N_2573,In_1001,In_1079);
or U2574 (N_2574,In_377,In_1386);
or U2575 (N_2575,In_1082,In_1147);
or U2576 (N_2576,In_359,In_759);
nor U2577 (N_2577,In_546,In_980);
and U2578 (N_2578,In_1360,In_899);
and U2579 (N_2579,In_497,In_852);
or U2580 (N_2580,In_88,In_324);
nor U2581 (N_2581,In_684,In_1232);
or U2582 (N_2582,In_625,In_977);
nor U2583 (N_2583,In_60,In_516);
and U2584 (N_2584,In_1115,In_1247);
or U2585 (N_2585,In_788,In_608);
or U2586 (N_2586,In_495,In_922);
nor U2587 (N_2587,In_483,In_513);
or U2588 (N_2588,In_849,In_1061);
nand U2589 (N_2589,In_174,In_984);
and U2590 (N_2590,In_1084,In_1129);
and U2591 (N_2591,In_231,In_1471);
and U2592 (N_2592,In_525,In_1231);
or U2593 (N_2593,In_723,In_168);
and U2594 (N_2594,In_216,In_575);
and U2595 (N_2595,In_794,In_732);
nor U2596 (N_2596,In_1074,In_445);
or U2597 (N_2597,In_1036,In_943);
and U2598 (N_2598,In_1160,In_289);
nand U2599 (N_2599,In_427,In_259);
or U2600 (N_2600,In_132,In_726);
or U2601 (N_2601,In_1337,In_562);
and U2602 (N_2602,In_489,In_808);
and U2603 (N_2603,In_43,In_255);
and U2604 (N_2604,In_224,In_1014);
nand U2605 (N_2605,In_1077,In_282);
or U2606 (N_2606,In_1158,In_1193);
nor U2607 (N_2607,In_217,In_792);
and U2608 (N_2608,In_1084,In_1203);
and U2609 (N_2609,In_126,In_1079);
nand U2610 (N_2610,In_1173,In_234);
and U2611 (N_2611,In_687,In_926);
or U2612 (N_2612,In_544,In_181);
or U2613 (N_2613,In_313,In_249);
nand U2614 (N_2614,In_763,In_372);
nor U2615 (N_2615,In_124,In_63);
nand U2616 (N_2616,In_524,In_1179);
nor U2617 (N_2617,In_952,In_216);
nor U2618 (N_2618,In_964,In_517);
nand U2619 (N_2619,In_135,In_94);
nor U2620 (N_2620,In_1100,In_1156);
nand U2621 (N_2621,In_833,In_1312);
or U2622 (N_2622,In_1183,In_174);
and U2623 (N_2623,In_183,In_1071);
nand U2624 (N_2624,In_708,In_1466);
or U2625 (N_2625,In_776,In_570);
and U2626 (N_2626,In_1082,In_787);
and U2627 (N_2627,In_1228,In_520);
nand U2628 (N_2628,In_85,In_1474);
nor U2629 (N_2629,In_1193,In_384);
and U2630 (N_2630,In_1346,In_346);
nand U2631 (N_2631,In_18,In_1381);
and U2632 (N_2632,In_287,In_1357);
or U2633 (N_2633,In_232,In_1349);
nor U2634 (N_2634,In_908,In_827);
nand U2635 (N_2635,In_1089,In_1432);
nor U2636 (N_2636,In_1408,In_271);
and U2637 (N_2637,In_152,In_501);
or U2638 (N_2638,In_844,In_654);
or U2639 (N_2639,In_1212,In_290);
nand U2640 (N_2640,In_145,In_904);
or U2641 (N_2641,In_1373,In_131);
nand U2642 (N_2642,In_735,In_964);
and U2643 (N_2643,In_839,In_954);
nand U2644 (N_2644,In_686,In_970);
nor U2645 (N_2645,In_713,In_37);
and U2646 (N_2646,In_813,In_529);
nor U2647 (N_2647,In_1484,In_336);
and U2648 (N_2648,In_1462,In_427);
nor U2649 (N_2649,In_874,In_178);
nand U2650 (N_2650,In_1160,In_1167);
nor U2651 (N_2651,In_907,In_402);
and U2652 (N_2652,In_636,In_305);
nand U2653 (N_2653,In_12,In_1211);
xnor U2654 (N_2654,In_1398,In_639);
nor U2655 (N_2655,In_177,In_676);
or U2656 (N_2656,In_1101,In_1465);
nor U2657 (N_2657,In_806,In_527);
nor U2658 (N_2658,In_661,In_981);
nand U2659 (N_2659,In_208,In_333);
xnor U2660 (N_2660,In_1380,In_640);
and U2661 (N_2661,In_1322,In_410);
and U2662 (N_2662,In_1255,In_1317);
nand U2663 (N_2663,In_307,In_439);
nand U2664 (N_2664,In_351,In_575);
nand U2665 (N_2665,In_1287,In_402);
nand U2666 (N_2666,In_332,In_562);
nand U2667 (N_2667,In_1010,In_812);
nor U2668 (N_2668,In_1063,In_1065);
nand U2669 (N_2669,In_136,In_714);
and U2670 (N_2670,In_1024,In_890);
nor U2671 (N_2671,In_1196,In_420);
nand U2672 (N_2672,In_179,In_697);
or U2673 (N_2673,In_323,In_701);
and U2674 (N_2674,In_1331,In_769);
and U2675 (N_2675,In_873,In_420);
nand U2676 (N_2676,In_694,In_129);
nand U2677 (N_2677,In_1048,In_1197);
nand U2678 (N_2678,In_1370,In_22);
and U2679 (N_2679,In_532,In_931);
or U2680 (N_2680,In_112,In_529);
and U2681 (N_2681,In_490,In_430);
and U2682 (N_2682,In_730,In_750);
nor U2683 (N_2683,In_426,In_1482);
and U2684 (N_2684,In_937,In_1432);
or U2685 (N_2685,In_1089,In_168);
and U2686 (N_2686,In_1230,In_146);
or U2687 (N_2687,In_280,In_1156);
nor U2688 (N_2688,In_1045,In_546);
nor U2689 (N_2689,In_438,In_1424);
nor U2690 (N_2690,In_1264,In_1358);
or U2691 (N_2691,In_95,In_323);
and U2692 (N_2692,In_37,In_1484);
or U2693 (N_2693,In_1046,In_701);
and U2694 (N_2694,In_16,In_540);
nand U2695 (N_2695,In_215,In_1373);
nor U2696 (N_2696,In_686,In_727);
nand U2697 (N_2697,In_1203,In_65);
nand U2698 (N_2698,In_1065,In_1208);
and U2699 (N_2699,In_874,In_773);
nor U2700 (N_2700,In_59,In_38);
nand U2701 (N_2701,In_444,In_1495);
xor U2702 (N_2702,In_107,In_378);
and U2703 (N_2703,In_1076,In_88);
or U2704 (N_2704,In_373,In_121);
and U2705 (N_2705,In_1057,In_734);
or U2706 (N_2706,In_813,In_116);
or U2707 (N_2707,In_17,In_591);
nand U2708 (N_2708,In_898,In_50);
nor U2709 (N_2709,In_1222,In_181);
and U2710 (N_2710,In_772,In_102);
nand U2711 (N_2711,In_1437,In_1274);
and U2712 (N_2712,In_805,In_815);
and U2713 (N_2713,In_1425,In_778);
nor U2714 (N_2714,In_1008,In_579);
nor U2715 (N_2715,In_532,In_1247);
or U2716 (N_2716,In_1254,In_371);
and U2717 (N_2717,In_835,In_934);
or U2718 (N_2718,In_1407,In_1030);
and U2719 (N_2719,In_1,In_509);
nor U2720 (N_2720,In_1481,In_1326);
and U2721 (N_2721,In_31,In_3);
and U2722 (N_2722,In_527,In_1043);
or U2723 (N_2723,In_190,In_407);
nor U2724 (N_2724,In_100,In_72);
xor U2725 (N_2725,In_631,In_1007);
and U2726 (N_2726,In_452,In_412);
nand U2727 (N_2727,In_1107,In_183);
or U2728 (N_2728,In_314,In_1353);
nor U2729 (N_2729,In_685,In_213);
nor U2730 (N_2730,In_919,In_23);
or U2731 (N_2731,In_1142,In_1106);
and U2732 (N_2732,In_1464,In_983);
nand U2733 (N_2733,In_689,In_848);
nor U2734 (N_2734,In_214,In_96);
or U2735 (N_2735,In_1192,In_38);
and U2736 (N_2736,In_628,In_652);
nand U2737 (N_2737,In_731,In_922);
nor U2738 (N_2738,In_292,In_642);
and U2739 (N_2739,In_1497,In_1294);
or U2740 (N_2740,In_709,In_205);
or U2741 (N_2741,In_193,In_689);
nand U2742 (N_2742,In_1157,In_1231);
nand U2743 (N_2743,In_446,In_77);
nor U2744 (N_2744,In_153,In_1359);
and U2745 (N_2745,In_1047,In_4);
and U2746 (N_2746,In_192,In_111);
and U2747 (N_2747,In_743,In_124);
nor U2748 (N_2748,In_593,In_119);
nor U2749 (N_2749,In_10,In_1351);
nor U2750 (N_2750,In_375,In_1289);
nand U2751 (N_2751,In_545,In_391);
and U2752 (N_2752,In_1407,In_1451);
or U2753 (N_2753,In_670,In_831);
and U2754 (N_2754,In_390,In_367);
or U2755 (N_2755,In_939,In_1124);
and U2756 (N_2756,In_599,In_737);
or U2757 (N_2757,In_574,In_666);
nand U2758 (N_2758,In_1349,In_767);
nor U2759 (N_2759,In_952,In_242);
or U2760 (N_2760,In_663,In_780);
nand U2761 (N_2761,In_1482,In_1191);
and U2762 (N_2762,In_942,In_90);
nor U2763 (N_2763,In_1405,In_432);
and U2764 (N_2764,In_1473,In_1424);
or U2765 (N_2765,In_735,In_372);
or U2766 (N_2766,In_734,In_530);
or U2767 (N_2767,In_301,In_128);
and U2768 (N_2768,In_686,In_879);
nor U2769 (N_2769,In_339,In_398);
nand U2770 (N_2770,In_829,In_500);
nor U2771 (N_2771,In_1395,In_1266);
or U2772 (N_2772,In_83,In_513);
or U2773 (N_2773,In_1336,In_1074);
or U2774 (N_2774,In_617,In_1062);
and U2775 (N_2775,In_894,In_638);
nor U2776 (N_2776,In_523,In_260);
or U2777 (N_2777,In_729,In_23);
and U2778 (N_2778,In_575,In_1140);
or U2779 (N_2779,In_765,In_55);
nand U2780 (N_2780,In_462,In_28);
nand U2781 (N_2781,In_290,In_622);
or U2782 (N_2782,In_703,In_1452);
nand U2783 (N_2783,In_1171,In_582);
nor U2784 (N_2784,In_1398,In_292);
nand U2785 (N_2785,In_1411,In_1460);
nand U2786 (N_2786,In_929,In_1250);
nor U2787 (N_2787,In_1127,In_1244);
nand U2788 (N_2788,In_656,In_1270);
nand U2789 (N_2789,In_1260,In_1389);
nand U2790 (N_2790,In_875,In_391);
xnor U2791 (N_2791,In_58,In_351);
nor U2792 (N_2792,In_1294,In_873);
nand U2793 (N_2793,In_433,In_762);
or U2794 (N_2794,In_808,In_705);
and U2795 (N_2795,In_757,In_764);
or U2796 (N_2796,In_96,In_1040);
and U2797 (N_2797,In_1416,In_1066);
or U2798 (N_2798,In_900,In_756);
nor U2799 (N_2799,In_116,In_896);
nor U2800 (N_2800,In_432,In_1161);
or U2801 (N_2801,In_863,In_509);
and U2802 (N_2802,In_974,In_297);
nor U2803 (N_2803,In_1382,In_359);
nand U2804 (N_2804,In_578,In_334);
or U2805 (N_2805,In_684,In_1314);
nand U2806 (N_2806,In_754,In_17);
nor U2807 (N_2807,In_1003,In_54);
and U2808 (N_2808,In_659,In_900);
or U2809 (N_2809,In_530,In_1421);
xnor U2810 (N_2810,In_930,In_678);
nor U2811 (N_2811,In_1319,In_594);
and U2812 (N_2812,In_1143,In_505);
and U2813 (N_2813,In_960,In_1498);
and U2814 (N_2814,In_871,In_979);
or U2815 (N_2815,In_1364,In_163);
nor U2816 (N_2816,In_210,In_130);
nand U2817 (N_2817,In_583,In_883);
and U2818 (N_2818,In_213,In_671);
and U2819 (N_2819,In_607,In_104);
or U2820 (N_2820,In_996,In_213);
or U2821 (N_2821,In_505,In_818);
nand U2822 (N_2822,In_62,In_1257);
nand U2823 (N_2823,In_971,In_369);
and U2824 (N_2824,In_1108,In_10);
and U2825 (N_2825,In_940,In_107);
and U2826 (N_2826,In_251,In_1376);
and U2827 (N_2827,In_1,In_1201);
and U2828 (N_2828,In_1357,In_102);
nor U2829 (N_2829,In_797,In_531);
nand U2830 (N_2830,In_427,In_653);
nor U2831 (N_2831,In_1325,In_1081);
nor U2832 (N_2832,In_452,In_1348);
nor U2833 (N_2833,In_260,In_431);
and U2834 (N_2834,In_1288,In_585);
and U2835 (N_2835,In_155,In_1488);
xor U2836 (N_2836,In_1395,In_305);
or U2837 (N_2837,In_329,In_1488);
nand U2838 (N_2838,In_553,In_689);
and U2839 (N_2839,In_1420,In_317);
and U2840 (N_2840,In_1420,In_93);
and U2841 (N_2841,In_234,In_475);
or U2842 (N_2842,In_555,In_217);
nand U2843 (N_2843,In_868,In_106);
xor U2844 (N_2844,In_686,In_71);
nand U2845 (N_2845,In_281,In_521);
and U2846 (N_2846,In_699,In_1391);
and U2847 (N_2847,In_1367,In_1285);
or U2848 (N_2848,In_1126,In_168);
and U2849 (N_2849,In_26,In_1420);
nor U2850 (N_2850,In_1000,In_959);
nand U2851 (N_2851,In_561,In_45);
nor U2852 (N_2852,In_699,In_1068);
nand U2853 (N_2853,In_1020,In_206);
nor U2854 (N_2854,In_596,In_194);
or U2855 (N_2855,In_1028,In_229);
and U2856 (N_2856,In_1279,In_49);
nor U2857 (N_2857,In_516,In_1433);
nor U2858 (N_2858,In_515,In_915);
and U2859 (N_2859,In_1414,In_301);
or U2860 (N_2860,In_188,In_922);
or U2861 (N_2861,In_1290,In_1422);
and U2862 (N_2862,In_606,In_459);
and U2863 (N_2863,In_1425,In_146);
and U2864 (N_2864,In_1037,In_247);
nand U2865 (N_2865,In_210,In_563);
nand U2866 (N_2866,In_372,In_607);
nand U2867 (N_2867,In_587,In_1025);
and U2868 (N_2868,In_221,In_152);
nor U2869 (N_2869,In_1455,In_1481);
and U2870 (N_2870,In_1052,In_108);
nor U2871 (N_2871,In_1267,In_199);
xnor U2872 (N_2872,In_1145,In_694);
or U2873 (N_2873,In_711,In_384);
nor U2874 (N_2874,In_311,In_154);
nor U2875 (N_2875,In_1051,In_812);
nand U2876 (N_2876,In_632,In_1478);
or U2877 (N_2877,In_738,In_1212);
nand U2878 (N_2878,In_877,In_1070);
nor U2879 (N_2879,In_801,In_1468);
nand U2880 (N_2880,In_274,In_346);
and U2881 (N_2881,In_1,In_474);
and U2882 (N_2882,In_419,In_454);
nor U2883 (N_2883,In_460,In_1051);
and U2884 (N_2884,In_878,In_791);
nor U2885 (N_2885,In_845,In_1092);
and U2886 (N_2886,In_477,In_141);
and U2887 (N_2887,In_832,In_346);
and U2888 (N_2888,In_307,In_186);
and U2889 (N_2889,In_286,In_568);
nor U2890 (N_2890,In_600,In_525);
or U2891 (N_2891,In_250,In_119);
nand U2892 (N_2892,In_1499,In_70);
nand U2893 (N_2893,In_1148,In_196);
nand U2894 (N_2894,In_163,In_1057);
or U2895 (N_2895,In_991,In_977);
nor U2896 (N_2896,In_100,In_18);
nand U2897 (N_2897,In_1409,In_767);
and U2898 (N_2898,In_610,In_389);
nand U2899 (N_2899,In_1360,In_136);
or U2900 (N_2900,In_1228,In_973);
and U2901 (N_2901,In_482,In_804);
and U2902 (N_2902,In_59,In_1387);
nand U2903 (N_2903,In_433,In_1148);
nand U2904 (N_2904,In_1362,In_1101);
nand U2905 (N_2905,In_1310,In_386);
and U2906 (N_2906,In_16,In_718);
and U2907 (N_2907,In_92,In_756);
nor U2908 (N_2908,In_601,In_28);
or U2909 (N_2909,In_1204,In_729);
nand U2910 (N_2910,In_561,In_818);
nand U2911 (N_2911,In_218,In_331);
nand U2912 (N_2912,In_181,In_464);
nand U2913 (N_2913,In_824,In_1461);
or U2914 (N_2914,In_721,In_895);
or U2915 (N_2915,In_666,In_343);
nand U2916 (N_2916,In_987,In_110);
nand U2917 (N_2917,In_1488,In_719);
and U2918 (N_2918,In_827,In_1146);
or U2919 (N_2919,In_550,In_444);
and U2920 (N_2920,In_924,In_1378);
or U2921 (N_2921,In_25,In_374);
nor U2922 (N_2922,In_1234,In_799);
or U2923 (N_2923,In_73,In_881);
nor U2924 (N_2924,In_1288,In_790);
nor U2925 (N_2925,In_796,In_867);
nand U2926 (N_2926,In_1008,In_922);
nor U2927 (N_2927,In_1436,In_1396);
nor U2928 (N_2928,In_273,In_1262);
or U2929 (N_2929,In_1152,In_844);
and U2930 (N_2930,In_478,In_362);
or U2931 (N_2931,In_796,In_822);
and U2932 (N_2932,In_1163,In_410);
nor U2933 (N_2933,In_314,In_220);
and U2934 (N_2934,In_1123,In_349);
nor U2935 (N_2935,In_883,In_1142);
and U2936 (N_2936,In_788,In_1093);
and U2937 (N_2937,In_812,In_1465);
and U2938 (N_2938,In_585,In_462);
nor U2939 (N_2939,In_1001,In_345);
and U2940 (N_2940,In_335,In_1131);
nand U2941 (N_2941,In_1409,In_1402);
nor U2942 (N_2942,In_981,In_934);
nand U2943 (N_2943,In_887,In_806);
nor U2944 (N_2944,In_1014,In_267);
nor U2945 (N_2945,In_817,In_726);
or U2946 (N_2946,In_1133,In_742);
nor U2947 (N_2947,In_1236,In_324);
nand U2948 (N_2948,In_1175,In_25);
nor U2949 (N_2949,In_409,In_1409);
nor U2950 (N_2950,In_1199,In_1079);
and U2951 (N_2951,In_470,In_1308);
nor U2952 (N_2952,In_1190,In_36);
nor U2953 (N_2953,In_1431,In_316);
or U2954 (N_2954,In_32,In_301);
and U2955 (N_2955,In_512,In_1476);
nand U2956 (N_2956,In_271,In_980);
nand U2957 (N_2957,In_901,In_124);
or U2958 (N_2958,In_185,In_1276);
nand U2959 (N_2959,In_1102,In_878);
or U2960 (N_2960,In_1059,In_49);
and U2961 (N_2961,In_655,In_1250);
nor U2962 (N_2962,In_909,In_448);
and U2963 (N_2963,In_268,In_152);
or U2964 (N_2964,In_490,In_716);
and U2965 (N_2965,In_284,In_389);
nor U2966 (N_2966,In_108,In_414);
nand U2967 (N_2967,In_23,In_1229);
and U2968 (N_2968,In_225,In_893);
nand U2969 (N_2969,In_1292,In_1442);
nand U2970 (N_2970,In_1173,In_1392);
nor U2971 (N_2971,In_741,In_145);
nand U2972 (N_2972,In_603,In_803);
and U2973 (N_2973,In_369,In_308);
nand U2974 (N_2974,In_221,In_599);
nand U2975 (N_2975,In_597,In_337);
and U2976 (N_2976,In_998,In_601);
and U2977 (N_2977,In_616,In_615);
nor U2978 (N_2978,In_758,In_1467);
nor U2979 (N_2979,In_1033,In_753);
or U2980 (N_2980,In_126,In_1164);
nand U2981 (N_2981,In_901,In_1488);
or U2982 (N_2982,In_415,In_1048);
and U2983 (N_2983,In_1182,In_596);
and U2984 (N_2984,In_45,In_771);
nor U2985 (N_2985,In_936,In_560);
and U2986 (N_2986,In_239,In_1447);
and U2987 (N_2987,In_728,In_695);
and U2988 (N_2988,In_422,In_1128);
nor U2989 (N_2989,In_500,In_142);
or U2990 (N_2990,In_386,In_12);
nor U2991 (N_2991,In_528,In_437);
nor U2992 (N_2992,In_940,In_1177);
nand U2993 (N_2993,In_507,In_1301);
nor U2994 (N_2994,In_58,In_1321);
or U2995 (N_2995,In_898,In_67);
nor U2996 (N_2996,In_568,In_386);
nand U2997 (N_2997,In_1364,In_265);
nor U2998 (N_2998,In_211,In_1296);
and U2999 (N_2999,In_240,In_174);
nor U3000 (N_3000,N_505,N_1417);
nor U3001 (N_3001,N_1840,N_482);
nor U3002 (N_3002,N_916,N_2269);
and U3003 (N_3003,N_1055,N_2775);
or U3004 (N_3004,N_926,N_530);
nand U3005 (N_3005,N_577,N_2914);
nor U3006 (N_3006,N_2151,N_984);
nand U3007 (N_3007,N_2366,N_1328);
nor U3008 (N_3008,N_150,N_2224);
nand U3009 (N_3009,N_1160,N_526);
and U3010 (N_3010,N_822,N_1660);
nor U3011 (N_3011,N_2799,N_1941);
nor U3012 (N_3012,N_1420,N_2465);
nor U3013 (N_3013,N_2476,N_120);
and U3014 (N_3014,N_764,N_1281);
nor U3015 (N_3015,N_2433,N_2412);
nor U3016 (N_3016,N_207,N_2895);
and U3017 (N_3017,N_581,N_614);
nand U3018 (N_3018,N_1183,N_1344);
xor U3019 (N_3019,N_1916,N_2184);
nand U3020 (N_3020,N_672,N_2674);
or U3021 (N_3021,N_1887,N_1307);
or U3022 (N_3022,N_2445,N_1630);
or U3023 (N_3023,N_771,N_2611);
and U3024 (N_3024,N_204,N_2940);
or U3025 (N_3025,N_912,N_1925);
nand U3026 (N_3026,N_1047,N_939);
nor U3027 (N_3027,N_1108,N_1746);
nor U3028 (N_3028,N_1681,N_411);
nor U3029 (N_3029,N_2804,N_814);
nand U3030 (N_3030,N_1111,N_2342);
or U3031 (N_3031,N_677,N_1121);
and U3032 (N_3032,N_1751,N_1566);
nor U3033 (N_3033,N_2540,N_2932);
or U3034 (N_3034,N_1377,N_1778);
and U3035 (N_3035,N_626,N_2163);
or U3036 (N_3036,N_2519,N_515);
and U3037 (N_3037,N_2573,N_1653);
or U3038 (N_3038,N_32,N_293);
and U3039 (N_3039,N_354,N_1277);
or U3040 (N_3040,N_1764,N_1644);
nor U3041 (N_3041,N_2138,N_365);
and U3042 (N_3042,N_195,N_2904);
or U3043 (N_3043,N_656,N_848);
and U3044 (N_3044,N_211,N_2650);
nand U3045 (N_3045,N_981,N_2442);
or U3046 (N_3046,N_798,N_527);
or U3047 (N_3047,N_1187,N_2222);
or U3048 (N_3048,N_683,N_2305);
nor U3049 (N_3049,N_2190,N_2318);
nor U3050 (N_3050,N_2927,N_2352);
nand U3051 (N_3051,N_2238,N_2763);
or U3052 (N_3052,N_2531,N_1898);
nand U3053 (N_3053,N_2434,N_478);
or U3054 (N_3054,N_2427,N_2438);
and U3055 (N_3055,N_1174,N_2529);
and U3056 (N_3056,N_1118,N_47);
or U3057 (N_3057,N_2871,N_933);
nor U3058 (N_3058,N_2546,N_215);
or U3059 (N_3059,N_2994,N_276);
nor U3060 (N_3060,N_2217,N_209);
nor U3061 (N_3061,N_1970,N_2992);
and U3062 (N_3062,N_1415,N_1383);
nand U3063 (N_3063,N_2309,N_746);
nand U3064 (N_3064,N_2512,N_2172);
nand U3065 (N_3065,N_494,N_2507);
nor U3066 (N_3066,N_1028,N_579);
and U3067 (N_3067,N_2637,N_2951);
nor U3068 (N_3068,N_2379,N_1019);
nor U3069 (N_3069,N_1608,N_2153);
and U3070 (N_3070,N_444,N_2171);
nand U3071 (N_3071,N_1255,N_1731);
or U3072 (N_3072,N_452,N_1928);
nor U3073 (N_3073,N_287,N_1797);
and U3074 (N_3074,N_689,N_2450);
nor U3075 (N_3075,N_1526,N_2387);
nor U3076 (N_3076,N_2235,N_2487);
and U3077 (N_3077,N_1318,N_1992);
nor U3078 (N_3078,N_2866,N_615);
or U3079 (N_3079,N_1037,N_156);
and U3080 (N_3080,N_2346,N_599);
and U3081 (N_3081,N_387,N_1379);
and U3082 (N_3082,N_2197,N_2758);
nand U3083 (N_3083,N_954,N_2586);
nor U3084 (N_3084,N_1408,N_1400);
and U3085 (N_3085,N_731,N_1575);
or U3086 (N_3086,N_2266,N_2214);
nand U3087 (N_3087,N_261,N_2762);
nor U3088 (N_3088,N_1842,N_2623);
nor U3089 (N_3089,N_1975,N_1150);
and U3090 (N_3090,N_2317,N_886);
or U3091 (N_3091,N_2769,N_236);
and U3092 (N_3092,N_659,N_1624);
nor U3093 (N_3093,N_1686,N_25);
nand U3094 (N_3094,N_2009,N_199);
nor U3095 (N_3095,N_2005,N_950);
or U3096 (N_3096,N_2626,N_2274);
or U3097 (N_3097,N_888,N_1169);
nor U3098 (N_3098,N_1509,N_1489);
or U3099 (N_3099,N_314,N_1772);
or U3100 (N_3100,N_319,N_2714);
nand U3101 (N_3101,N_1292,N_1996);
nor U3102 (N_3102,N_73,N_2661);
nor U3103 (N_3103,N_2015,N_2500);
and U3104 (N_3104,N_2035,N_832);
nor U3105 (N_3105,N_2863,N_2618);
or U3106 (N_3106,N_968,N_84);
nor U3107 (N_3107,N_1560,N_2948);
nand U3108 (N_3108,N_1597,N_1508);
or U3109 (N_3109,N_343,N_2440);
nand U3110 (N_3110,N_38,N_1079);
or U3111 (N_3111,N_1395,N_1024);
nand U3112 (N_3112,N_959,N_1533);
or U3113 (N_3113,N_2400,N_2303);
nand U3114 (N_3114,N_177,N_2826);
nor U3115 (N_3115,N_192,N_938);
and U3116 (N_3116,N_213,N_2415);
xnor U3117 (N_3117,N_1014,N_2162);
and U3118 (N_3118,N_961,N_486);
and U3119 (N_3119,N_1218,N_1359);
nand U3120 (N_3120,N_2959,N_1333);
nand U3121 (N_3121,N_2552,N_2955);
nand U3122 (N_3122,N_131,N_2845);
and U3123 (N_3123,N_812,N_106);
nor U3124 (N_3124,N_1213,N_2745);
and U3125 (N_3125,N_2501,N_2472);
nor U3126 (N_3126,N_2380,N_2348);
nand U3127 (N_3127,N_2407,N_949);
nand U3128 (N_3128,N_989,N_1286);
or U3129 (N_3129,N_250,N_540);
or U3130 (N_3130,N_1211,N_2215);
nand U3131 (N_3131,N_2046,N_1003);
nor U3132 (N_3132,N_1242,N_191);
and U3133 (N_3133,N_45,N_2810);
or U3134 (N_3134,N_266,N_2700);
and U3135 (N_3135,N_2879,N_562);
nor U3136 (N_3136,N_841,N_2524);
and U3137 (N_3137,N_90,N_2135);
nor U3138 (N_3138,N_2658,N_248);
or U3139 (N_3139,N_49,N_1651);
nor U3140 (N_3140,N_2202,N_1029);
nand U3141 (N_3141,N_1872,N_2926);
or U3142 (N_3142,N_2513,N_1205);
nor U3143 (N_3143,N_818,N_684);
nand U3144 (N_3144,N_1511,N_1816);
or U3145 (N_3145,N_2456,N_847);
nand U3146 (N_3146,N_2329,N_1084);
and U3147 (N_3147,N_2613,N_1865);
and U3148 (N_3148,N_870,N_2690);
nor U3149 (N_3149,N_1409,N_1969);
nand U3150 (N_3150,N_1188,N_747);
and U3151 (N_3151,N_617,N_291);
or U3152 (N_3152,N_1806,N_2699);
or U3153 (N_3153,N_2185,N_2575);
or U3154 (N_3154,N_176,N_2917);
or U3155 (N_3155,N_2077,N_558);
nor U3156 (N_3156,N_2654,N_2752);
and U3157 (N_3157,N_2390,N_2891);
nand U3158 (N_3158,N_2378,N_76);
and U3159 (N_3159,N_1684,N_2023);
nor U3160 (N_3160,N_2635,N_1190);
and U3161 (N_3161,N_2156,N_2727);
and U3162 (N_3162,N_16,N_113);
or U3163 (N_3163,N_1454,N_1294);
nor U3164 (N_3164,N_1912,N_260);
or U3165 (N_3165,N_749,N_1008);
and U3166 (N_3166,N_1657,N_2045);
and U3167 (N_3167,N_1885,N_2027);
nor U3168 (N_3168,N_1354,N_2330);
and U3169 (N_3169,N_1064,N_2053);
nor U3170 (N_3170,N_1607,N_1752);
nand U3171 (N_3171,N_2502,N_2285);
nand U3172 (N_3172,N_1500,N_552);
or U3173 (N_3173,N_1675,N_1894);
or U3174 (N_3174,N_2398,N_2681);
or U3175 (N_3175,N_869,N_362);
nor U3176 (N_3176,N_2278,N_1423);
or U3177 (N_3177,N_519,N_671);
nor U3178 (N_3178,N_2569,N_1131);
nor U3179 (N_3179,N_1601,N_448);
nand U3180 (N_3180,N_393,N_1663);
nor U3181 (N_3181,N_2292,N_0);
nor U3182 (N_3182,N_1957,N_1987);
nand U3183 (N_3183,N_418,N_190);
nand U3184 (N_3184,N_1800,N_1234);
or U3185 (N_3185,N_2017,N_842);
nand U3186 (N_3186,N_1151,N_2242);
or U3187 (N_3187,N_12,N_1319);
and U3188 (N_3188,N_2978,N_2470);
and U3189 (N_3189,N_1228,N_2832);
and U3190 (N_3190,N_2028,N_602);
and U3191 (N_3191,N_69,N_2272);
and U3192 (N_3192,N_435,N_43);
nand U3193 (N_3193,N_955,N_1133);
or U3194 (N_3194,N_2413,N_2559);
nor U3195 (N_3195,N_854,N_2038);
or U3196 (N_3196,N_681,N_1632);
and U3197 (N_3197,N_244,N_1273);
nand U3198 (N_3198,N_1459,N_2852);
nand U3199 (N_3199,N_2283,N_1949);
and U3200 (N_3200,N_1737,N_1378);
or U3201 (N_3201,N_2980,N_2902);
and U3202 (N_3202,N_1787,N_1367);
or U3203 (N_3203,N_117,N_1452);
nor U3204 (N_3204,N_2882,N_1026);
nor U3205 (N_3205,N_705,N_1506);
nor U3206 (N_3206,N_1515,N_1586);
and U3207 (N_3207,N_1253,N_1936);
nor U3208 (N_3208,N_2706,N_2818);
nand U3209 (N_3209,N_1443,N_2289);
and U3210 (N_3210,N_1411,N_502);
nand U3211 (N_3211,N_1860,N_1825);
nand U3212 (N_3212,N_2008,N_1775);
nor U3213 (N_3213,N_2414,N_2191);
nand U3214 (N_3214,N_161,N_256);
nand U3215 (N_3215,N_1375,N_2454);
and U3216 (N_3216,N_422,N_918);
nand U3217 (N_3217,N_971,N_1082);
xor U3218 (N_3218,N_594,N_2733);
or U3219 (N_3219,N_688,N_2155);
nand U3220 (N_3220,N_2543,N_722);
or U3221 (N_3221,N_605,N_126);
or U3222 (N_3222,N_2622,N_229);
nand U3223 (N_3223,N_2482,N_2725);
nand U3224 (N_3224,N_275,N_1274);
nor U3225 (N_3225,N_1126,N_2560);
nor U3226 (N_3226,N_1493,N_2312);
nor U3227 (N_3227,N_568,N_2234);
nand U3228 (N_3228,N_2843,N_1695);
nand U3229 (N_3229,N_2423,N_392);
xnor U3230 (N_3230,N_887,N_1611);
nand U3231 (N_3231,N_1226,N_995);
nor U3232 (N_3232,N_274,N_1603);
nor U3233 (N_3233,N_1818,N_980);
and U3234 (N_3234,N_2511,N_167);
nor U3235 (N_3235,N_1374,N_1680);
or U3236 (N_3236,N_144,N_2987);
nor U3237 (N_3237,N_1052,N_1606);
or U3238 (N_3238,N_1640,N_368);
nand U3239 (N_3239,N_1262,N_1462);
nand U3240 (N_3240,N_311,N_181);
and U3241 (N_3241,N_62,N_1753);
and U3242 (N_3242,N_1291,N_1537);
nor U3243 (N_3243,N_1312,N_2273);
or U3244 (N_3244,N_2416,N_2912);
and U3245 (N_3245,N_2182,N_1336);
or U3246 (N_3246,N_2319,N_1756);
nand U3247 (N_3247,N_456,N_2750);
nand U3248 (N_3248,N_442,N_833);
nand U3249 (N_3249,N_59,N_1155);
nor U3250 (N_3250,N_99,N_598);
nor U3251 (N_3251,N_129,N_1967);
nand U3252 (N_3252,N_2030,N_258);
nor U3253 (N_3253,N_1296,N_2647);
or U3254 (N_3254,N_2279,N_619);
and U3255 (N_3255,N_541,N_44);
nor U3256 (N_3256,N_2006,N_2213);
nand U3257 (N_3257,N_212,N_1505);
and U3258 (N_3258,N_2024,N_1889);
or U3259 (N_3259,N_2111,N_109);
nand U3260 (N_3260,N_1143,N_2694);
nand U3261 (N_3261,N_667,N_537);
or U3262 (N_3262,N_1195,N_1596);
nor U3263 (N_3263,N_42,N_1365);
and U3264 (N_3264,N_1757,N_1884);
and U3265 (N_3265,N_240,N_2859);
or U3266 (N_3266,N_769,N_1159);
and U3267 (N_3267,N_1634,N_1231);
nand U3268 (N_3268,N_139,N_481);
or U3269 (N_3269,N_2241,N_1387);
nand U3270 (N_3270,N_1943,N_533);
or U3271 (N_3271,N_100,N_158);
or U3272 (N_3272,N_1820,N_1981);
nand U3273 (N_3273,N_2148,N_1774);
nand U3274 (N_3274,N_1050,N_1869);
and U3275 (N_3275,N_2475,N_264);
nand U3276 (N_3276,N_2328,N_2106);
and U3277 (N_3277,N_2239,N_650);
nand U3278 (N_3278,N_2154,N_1385);
nor U3279 (N_3279,N_2965,N_2625);
nor U3280 (N_3280,N_1587,N_2287);
and U3281 (N_3281,N_1892,N_2291);
nand U3282 (N_3282,N_2459,N_378);
or U3283 (N_3283,N_1549,N_346);
nor U3284 (N_3284,N_2517,N_535);
nand U3285 (N_3285,N_2515,N_903);
or U3286 (N_3286,N_2789,N_2933);
nor U3287 (N_3287,N_1341,N_151);
nor U3288 (N_3288,N_1132,N_1594);
and U3289 (N_3289,N_1067,N_1538);
or U3290 (N_3290,N_2064,N_1573);
and U3291 (N_3291,N_2439,N_408);
or U3292 (N_3292,N_1267,N_432);
or U3293 (N_3293,N_1781,N_1283);
or U3294 (N_3294,N_600,N_409);
and U3295 (N_3295,N_678,N_445);
nand U3296 (N_3296,N_2572,N_509);
and U3297 (N_3297,N_2549,N_71);
and U3298 (N_3298,N_2334,N_18);
nor U3299 (N_3299,N_267,N_1995);
and U3300 (N_3300,N_107,N_2907);
or U3301 (N_3301,N_2911,N_1355);
and U3302 (N_3302,N_2816,N_1202);
nor U3303 (N_3303,N_786,N_1481);
or U3304 (N_3304,N_761,N_2688);
nand U3305 (N_3305,N_273,N_1112);
or U3306 (N_3306,N_2353,N_2276);
nor U3307 (N_3307,N_2254,N_1435);
and U3308 (N_3308,N_2748,N_2704);
nand U3309 (N_3309,N_676,N_1652);
and U3310 (N_3310,N_585,N_404);
and U3311 (N_3311,N_24,N_196);
and U3312 (N_3312,N_825,N_1373);
nor U3313 (N_3313,N_2297,N_936);
nor U3314 (N_3314,N_1043,N_8);
nand U3315 (N_3315,N_1641,N_410);
and U3316 (N_3316,N_200,N_88);
nand U3317 (N_3317,N_2211,N_1572);
or U3318 (N_3318,N_119,N_1440);
and U3319 (N_3319,N_1470,N_490);
nand U3320 (N_3320,N_2055,N_1280);
and U3321 (N_3321,N_1331,N_2447);
nor U3322 (N_3322,N_782,N_203);
or U3323 (N_3323,N_1361,N_155);
nand U3324 (N_3324,N_367,N_1215);
and U3325 (N_3325,N_2127,N_2856);
and U3326 (N_3326,N_1540,N_403);
nor U3327 (N_3327,N_114,N_2836);
or U3328 (N_3328,N_1703,N_2842);
nand U3329 (N_3329,N_172,N_1713);
and U3330 (N_3330,N_1144,N_564);
or U3331 (N_3331,N_852,N_2264);
nor U3332 (N_3332,N_1780,N_2033);
nor U3333 (N_3333,N_2644,N_1600);
nor U3334 (N_3334,N_2263,N_1918);
and U3335 (N_3335,N_92,N_1707);
and U3336 (N_3336,N_280,N_2553);
or U3337 (N_3337,N_2953,N_2288);
nor U3338 (N_3338,N_592,N_546);
or U3339 (N_3339,N_1221,N_2490);
and U3340 (N_3340,N_2558,N_773);
nand U3341 (N_3341,N_1716,N_2503);
nand U3342 (N_3342,N_1418,N_2275);
or U3343 (N_3343,N_2041,N_2599);
and U3344 (N_3344,N_2983,N_2831);
and U3345 (N_3345,N_727,N_840);
or U3346 (N_3346,N_1033,N_883);
xor U3347 (N_3347,N_1140,N_2117);
or U3348 (N_3348,N_2938,N_2884);
nor U3349 (N_3349,N_737,N_2099);
nor U3350 (N_3350,N_1313,N_2228);
nand U3351 (N_3351,N_1123,N_2510);
nand U3352 (N_3352,N_508,N_1117);
or U3353 (N_3353,N_1935,N_2491);
nor U3354 (N_3354,N_1798,N_1946);
nor U3355 (N_3355,N_2641,N_2528);
or U3356 (N_3356,N_548,N_1185);
or U3357 (N_3357,N_122,N_2666);
nand U3358 (N_3358,N_610,N_2136);
or U3359 (N_3359,N_1182,N_189);
nor U3360 (N_3360,N_2170,N_874);
nor U3361 (N_3361,N_1839,N_2537);
nor U3362 (N_3362,N_728,N_159);
nor U3363 (N_3363,N_2853,N_2662);
nand U3364 (N_3364,N_770,N_1930);
nor U3365 (N_3365,N_2794,N_1261);
nor U3366 (N_3366,N_538,N_1002);
nor U3367 (N_3367,N_231,N_1334);
nand U3368 (N_3368,N_2243,N_796);
and U3369 (N_3369,N_2449,N_2967);
or U3370 (N_3370,N_1929,N_2361);
nand U3371 (N_3371,N_1295,N_2555);
nand U3372 (N_3372,N_1623,N_2092);
or U3373 (N_3373,N_111,N_463);
nor U3374 (N_3374,N_2075,N_2091);
and U3375 (N_3375,N_911,N_487);
nor U3376 (N_3376,N_1525,N_462);
or U3377 (N_3377,N_1063,N_1069);
nor U3378 (N_3378,N_68,N_868);
nand U3379 (N_3379,N_2350,N_182);
nor U3380 (N_3380,N_1460,N_2749);
or U3381 (N_3381,N_1348,N_2939);
nor U3382 (N_3382,N_2682,N_294);
nand U3383 (N_3383,N_2963,N_66);
nor U3384 (N_3384,N_664,N_2742);
nand U3385 (N_3385,N_1167,N_1768);
and U3386 (N_3386,N_709,N_976);
nor U3387 (N_3387,N_1206,N_2869);
nor U3388 (N_3388,N_265,N_2444);
nor U3389 (N_3389,N_531,N_2129);
nor U3390 (N_3390,N_1832,N_867);
nand U3391 (N_3391,N_823,N_687);
or U3392 (N_3392,N_363,N_501);
or U3393 (N_3393,N_757,N_458);
or U3394 (N_3394,N_2498,N_1306);
nand U3395 (N_3395,N_2893,N_1471);
nor U3396 (N_3396,N_1396,N_986);
nor U3397 (N_3397,N_2889,N_2088);
nand U3398 (N_3398,N_1837,N_1672);
or U3399 (N_3399,N_464,N_1258);
and U3400 (N_3400,N_1044,N_72);
or U3401 (N_3401,N_227,N_732);
nor U3402 (N_3402,N_2801,N_93);
or U3403 (N_3403,N_2399,N_1626);
nor U3404 (N_3404,N_108,N_1848);
nor U3405 (N_3405,N_1032,N_712);
nor U3406 (N_3406,N_1197,N_1137);
or U3407 (N_3407,N_2245,N_64);
nand U3408 (N_3408,N_2771,N_551);
or U3409 (N_3409,N_1490,N_194);
nor U3410 (N_3410,N_2474,N_202);
and U3411 (N_3411,N_1475,N_1308);
or U3412 (N_3412,N_1220,N_919);
nand U3413 (N_3413,N_1807,N_5);
or U3414 (N_3414,N_510,N_729);
or U3415 (N_3415,N_2014,N_2726);
nand U3416 (N_3416,N_2640,N_948);
nand U3417 (N_3417,N_1156,N_1759);
xor U3418 (N_3418,N_2548,N_629);
nor U3419 (N_3419,N_1543,N_471);
and U3420 (N_3420,N_717,N_1507);
and U3421 (N_3421,N_1789,N_815);
nand U3422 (N_3422,N_2071,N_1429);
and U3423 (N_3423,N_2128,N_1605);
nor U3424 (N_3424,N_1804,N_1610);
or U3425 (N_3425,N_2057,N_216);
or U3426 (N_3426,N_2974,N_574);
nor U3427 (N_3427,N_2945,N_1698);
nand U3428 (N_3428,N_1254,N_1547);
and U3429 (N_3429,N_1722,N_2047);
nor U3430 (N_3430,N_193,N_1399);
and U3431 (N_3431,N_576,N_2885);
xnor U3432 (N_3432,N_760,N_801);
nand U3433 (N_3433,N_1243,N_2499);
nor U3434 (N_3434,N_357,N_921);
nand U3435 (N_3435,N_377,N_1908);
nor U3436 (N_3436,N_1322,N_891);
nand U3437 (N_3437,N_1670,N_2477);
nor U3438 (N_3438,N_2850,N_1776);
or U3439 (N_3439,N_1467,N_2374);
or U3440 (N_3440,N_2429,N_1593);
or U3441 (N_3441,N_1934,N_1521);
or U3442 (N_3442,N_2061,N_1915);
nor U3443 (N_3443,N_2918,N_1369);
nand U3444 (N_3444,N_1676,N_2478);
nand U3445 (N_3445,N_2149,N_1227);
nand U3446 (N_3446,N_457,N_2356);
nor U3447 (N_3447,N_30,N_178);
nor U3448 (N_3448,N_384,N_292);
nand U3449 (N_3449,N_329,N_97);
xor U3450 (N_3450,N_2073,N_1158);
nor U3451 (N_3451,N_1057,N_1141);
or U3452 (N_3452,N_517,N_696);
nor U3453 (N_3453,N_2814,N_1788);
nand U3454 (N_3454,N_305,N_221);
and U3455 (N_3455,N_2109,N_1583);
nand U3456 (N_3456,N_2695,N_1455);
and U3457 (N_3457,N_2645,N_1579);
or U3458 (N_3458,N_957,N_2591);
nor U3459 (N_3459,N_1413,N_612);
and U3460 (N_3460,N_2737,N_2257);
nand U3461 (N_3461,N_1422,N_1472);
nor U3462 (N_3462,N_1072,N_210);
and U3463 (N_3463,N_1961,N_246);
nand U3464 (N_3464,N_1629,N_1609);
and U3465 (N_3465,N_2739,N_2971);
and U3466 (N_3466,N_2324,N_2589);
and U3467 (N_3467,N_2382,N_1222);
nand U3468 (N_3468,N_616,N_2942);
or U3469 (N_3469,N_2880,N_2315);
and U3470 (N_3470,N_2797,N_2004);
and U3471 (N_3471,N_1666,N_2188);
xnor U3472 (N_3472,N_2335,N_2039);
and U3473 (N_3473,N_2410,N_865);
or U3474 (N_3474,N_2620,N_2115);
nor U3475 (N_3475,N_2158,N_2998);
nand U3476 (N_3476,N_2604,N_2805);
nand U3477 (N_3477,N_927,N_2541);
and U3478 (N_3478,N_2208,N_372);
nor U3479 (N_3479,N_2034,N_660);
nor U3480 (N_3480,N_861,N_1199);
nand U3481 (N_3481,N_1264,N_1794);
nand U3482 (N_3482,N_647,N_1351);
and U3483 (N_3483,N_1165,N_1633);
nor U3484 (N_3484,N_2143,N_2327);
nor U3485 (N_3485,N_914,N_78);
nor U3486 (N_3486,N_469,N_682);
and U3487 (N_3487,N_1450,N_904);
and U3488 (N_3488,N_1311,N_850);
or U3489 (N_3489,N_613,N_834);
and U3490 (N_3490,N_1053,N_2890);
or U3491 (N_3491,N_2878,N_1551);
nand U3492 (N_3492,N_1958,N_803);
nor U3493 (N_3493,N_2584,N_2874);
nand U3494 (N_3494,N_358,N_1042);
nand U3495 (N_3495,N_811,N_75);
nand U3496 (N_3496,N_966,N_2977);
and U3497 (N_3497,N_450,N_1092);
and U3498 (N_3498,N_1007,N_2731);
and U3499 (N_3499,N_2081,N_931);
nand U3500 (N_3500,N_2082,N_2743);
and U3501 (N_3501,N_2137,N_839);
and U3502 (N_3502,N_2146,N_2363);
nor U3503 (N_3503,N_2962,N_1643);
or U3504 (N_3504,N_36,N_1799);
nand U3505 (N_3505,N_2935,N_2673);
and U3506 (N_3506,N_2322,N_2621);
and U3507 (N_3507,N_2282,N_1457);
nand U3508 (N_3508,N_2209,N_1530);
and U3509 (N_3509,N_440,N_928);
or U3510 (N_3510,N_2226,N_2761);
nor U3511 (N_3511,N_649,N_1847);
and U3512 (N_3512,N_2493,N_6);
nand U3513 (N_3513,N_2397,N_166);
and U3514 (N_3514,N_956,N_1714);
and U3515 (N_3515,N_1923,N_744);
and U3516 (N_3516,N_2747,N_1699);
or U3517 (N_3517,N_313,N_1817);
nand U3518 (N_3518,N_1099,N_521);
or U3519 (N_3519,N_1927,N_2059);
nor U3520 (N_3520,N_2248,N_371);
and U3521 (N_3521,N_2565,N_853);
nor U3522 (N_3522,N_560,N_2516);
nand U3523 (N_3523,N_2594,N_1906);
or U3524 (N_3524,N_2424,N_1993);
or U3525 (N_3525,N_695,N_396);
or U3526 (N_3526,N_1136,N_2691);
or U3527 (N_3527,N_1284,N_1726);
nand U3528 (N_3528,N_37,N_673);
or U3529 (N_3529,N_2409,N_439);
nor U3530 (N_3530,N_2609,N_896);
nand U3531 (N_3531,N_1896,N_2360);
nand U3532 (N_3532,N_54,N_550);
nor U3533 (N_3533,N_174,N_2396);
nand U3534 (N_3534,N_1683,N_31);
xnor U3535 (N_3535,N_1074,N_2568);
or U3536 (N_3536,N_366,N_1562);
and U3537 (N_3537,N_2815,N_1671);
nor U3538 (N_3538,N_1661,N_2394);
and U3539 (N_3539,N_1461,N_230);
or U3540 (N_3540,N_297,N_2970);
nand U3541 (N_3541,N_56,N_972);
nor U3542 (N_3542,N_1882,N_1363);
or U3543 (N_3543,N_937,N_2132);
or U3544 (N_3544,N_2612,N_436);
and U3545 (N_3545,N_2007,N_2633);
or U3546 (N_3546,N_762,N_1687);
nand U3547 (N_3547,N_2139,N_413);
or U3548 (N_3548,N_2657,N_1679);
nor U3549 (N_3549,N_1001,N_2509);
nand U3550 (N_3550,N_1548,N_2002);
nor U3551 (N_3551,N_1658,N_698);
or U3552 (N_3552,N_2649,N_1576);
nand U3553 (N_3553,N_2876,N_2103);
nor U3554 (N_3554,N_2323,N_1040);
or U3555 (N_3555,N_2984,N_2125);
or U3556 (N_3556,N_2958,N_1942);
nor U3557 (N_3557,N_1948,N_2692);
nand U3558 (N_3558,N_829,N_943);
nor U3559 (N_3559,N_1479,N_2683);
nor U3560 (N_3560,N_958,N_699);
nor U3561 (N_3561,N_2430,N_431);
nor U3562 (N_3562,N_1071,N_742);
and U3563 (N_3563,N_1394,N_1636);
nor U3564 (N_3564,N_352,N_1054);
nand U3565 (N_3565,N_2908,N_645);
nor U3566 (N_3566,N_1316,N_589);
or U3567 (N_3567,N_1477,N_2240);
and U3568 (N_3568,N_2693,N_270);
and U3569 (N_3569,N_70,N_2147);
nand U3570 (N_3570,N_2044,N_233);
nand U3571 (N_3571,N_2,N_991);
or U3572 (N_3572,N_2710,N_2364);
nor U3573 (N_3573,N_944,N_2999);
and U3574 (N_3574,N_1592,N_720);
or U3575 (N_3575,N_845,N_1482);
nor U3576 (N_3576,N_1905,N_1762);
or U3577 (N_3577,N_2587,N_488);
and U3578 (N_3578,N_2299,N_1203);
and U3579 (N_3579,N_655,N_670);
or U3580 (N_3580,N_2066,N_2756);
nand U3581 (N_3581,N_2376,N_1810);
nand U3582 (N_3582,N_1401,N_1251);
nand U3583 (N_3583,N_434,N_1667);
nor U3584 (N_3584,N_666,N_1888);
nand U3585 (N_3585,N_1720,N_637);
and U3586 (N_3586,N_994,N_2165);
nand U3587 (N_3587,N_85,N_2422);
and U3588 (N_3588,N_1285,N_259);
nor U3589 (N_3589,N_1747,N_1956);
or U3590 (N_3590,N_2578,N_996);
and U3591 (N_3591,N_2957,N_2574);
and U3592 (N_3592,N_2892,N_1718);
nand U3593 (N_3593,N_2065,N_1602);
and U3594 (N_3594,N_1162,N_1559);
nor U3595 (N_3595,N_2603,N_1436);
and U3596 (N_3596,N_566,N_1648);
nor U3597 (N_3597,N_1910,N_2233);
or U3598 (N_3598,N_2684,N_1094);
nor U3599 (N_3599,N_2123,N_1012);
nor U3600 (N_3600,N_417,N_1104);
nor U3601 (N_3601,N_1402,N_859);
nand U3602 (N_3602,N_1058,N_1542);
nor U3603 (N_3603,N_809,N_1763);
nor U3604 (N_3604,N_1109,N_1971);
nand U3605 (N_3605,N_553,N_824);
nor U3606 (N_3606,N_1899,N_1940);
nor U3607 (N_3607,N_2913,N_2915);
nor U3608 (N_3608,N_2943,N_2544);
nand U3609 (N_3609,N_2773,N_2563);
nor U3610 (N_3610,N_2484,N_2670);
nor U3611 (N_3611,N_1580,N_1729);
or U3612 (N_3612,N_1755,N_391);
and U3613 (N_3613,N_2837,N_880);
and U3614 (N_3614,N_1968,N_2950);
or U3615 (N_3615,N_1909,N_118);
nor U3616 (N_3616,N_152,N_573);
nor U3617 (N_3617,N_480,N_2766);
nand U3618 (N_3618,N_1965,N_1004);
and U3619 (N_3619,N_2451,N_940);
nor U3620 (N_3620,N_703,N_1513);
or U3621 (N_3621,N_2417,N_1225);
nand U3622 (N_3622,N_1265,N_473);
and U3623 (N_3623,N_285,N_154);
and U3624 (N_3624,N_2483,N_1510);
or U3625 (N_3625,N_46,N_1237);
nand U3626 (N_3626,N_1767,N_1142);
or U3627 (N_3627,N_2952,N_340);
or U3628 (N_3628,N_1921,N_40);
or U3629 (N_3629,N_2802,N_288);
nor U3630 (N_3630,N_2403,N_1239);
nand U3631 (N_3631,N_2753,N_479);
and U3632 (N_3632,N_2672,N_843);
nor U3633 (N_3633,N_415,N_544);
and U3634 (N_3634,N_350,N_1438);
nor U3635 (N_3635,N_1372,N_751);
or U3636 (N_3636,N_449,N_2277);
and U3637 (N_3637,N_1276,N_2598);
or U3638 (N_3638,N_962,N_795);
or U3639 (N_3639,N_290,N_427);
or U3640 (N_3640,N_788,N_2697);
or U3641 (N_3641,N_1858,N_1193);
and U3642 (N_3642,N_2250,N_249);
or U3643 (N_3643,N_628,N_1326);
nor U3644 (N_3644,N_2218,N_772);
or U3645 (N_3645,N_1476,N_718);
nor U3646 (N_3646,N_2085,N_1782);
nor U3647 (N_3647,N_1442,N_2833);
nor U3648 (N_3648,N_945,N_1883);
nor U3649 (N_3649,N_2679,N_1432);
nor U3650 (N_3650,N_1080,N_1900);
and U3651 (N_3651,N_635,N_2189);
nand U3652 (N_3652,N_1289,N_1783);
or U3653 (N_3653,N_2705,N_2261);
nand U3654 (N_3654,N_2734,N_1880);
nand U3655 (N_3655,N_2441,N_1495);
nand U3656 (N_3656,N_1127,N_20);
nor U3657 (N_3657,N_1717,N_810);
nand U3658 (N_3658,N_1618,N_1520);
and U3659 (N_3659,N_2779,N_138);
nor U3660 (N_3660,N_1332,N_1320);
and U3661 (N_3661,N_730,N_702);
and U3662 (N_3662,N_125,N_778);
nor U3663 (N_3663,N_2131,N_1678);
and U3664 (N_3664,N_1911,N_1161);
nand U3665 (N_3665,N_2080,N_2855);
or U3666 (N_3666,N_1487,N_2112);
nor U3667 (N_3667,N_608,N_451);
nor U3668 (N_3668,N_121,N_2956);
or U3669 (N_3669,N_1544,N_302);
or U3670 (N_3670,N_1163,N_2486);
nor U3671 (N_3671,N_1639,N_2419);
and U3672 (N_3672,N_2341,N_2037);
nand U3673 (N_3673,N_2227,N_2386);
and U3674 (N_3674,N_334,N_498);
or U3675 (N_3675,N_15,N_1146);
and U3676 (N_3676,N_653,N_2471);
nor U3677 (N_3677,N_1769,N_2296);
or U3678 (N_3678,N_421,N_1179);
or U3679 (N_3679,N_1129,N_1330);
nand U3680 (N_3680,N_103,N_1913);
and U3681 (N_3681,N_2489,N_2058);
or U3682 (N_3682,N_2492,N_1447);
or U3683 (N_3683,N_1122,N_1512);
and U3684 (N_3684,N_2910,N_2995);
nand U3685 (N_3685,N_1113,N_269);
or U3686 (N_3686,N_1299,N_2851);
nand U3687 (N_3687,N_2997,N_2068);
nor U3688 (N_3688,N_461,N_819);
nand U3689 (N_3689,N_1492,N_247);
nor U3690 (N_3690,N_1335,N_733);
or U3691 (N_3691,N_2777,N_206);
nor U3692 (N_3692,N_1514,N_1719);
nand U3693 (N_3693,N_2659,N_1863);
nor U3694 (N_3694,N_680,N_1115);
nand U3695 (N_3695,N_443,N_2113);
nor U3696 (N_3696,N_1979,N_1293);
or U3697 (N_3697,N_224,N_2530);
nor U3698 (N_3698,N_2596,N_783);
nand U3699 (N_3699,N_9,N_1083);
nor U3700 (N_3700,N_2698,N_2122);
or U3701 (N_3701,N_2094,N_2839);
and U3702 (N_3702,N_754,N_489);
or U3703 (N_3703,N_2104,N_1469);
and U3704 (N_3704,N_1743,N_1250);
or U3705 (N_3705,N_793,N_557);
and U3706 (N_3706,N_1749,N_95);
or U3707 (N_3707,N_1392,N_1890);
nand U3708 (N_3708,N_807,N_2947);
and U3709 (N_3709,N_1194,N_2772);
or U3710 (N_3710,N_390,N_308);
nor U3711 (N_3711,N_1453,N_2174);
nand U3712 (N_3712,N_2899,N_663);
and U3713 (N_3713,N_1920,N_779);
nand U3714 (N_3714,N_2642,N_2554);
or U3715 (N_3715,N_1868,N_2086);
nor U3716 (N_3716,N_2982,N_1516);
and U3717 (N_3717,N_741,N_1616);
nor U3718 (N_3718,N_112,N_1473);
nor U3719 (N_3719,N_1070,N_2898);
and U3720 (N_3720,N_2067,N_2542);
nor U3721 (N_3721,N_2126,N_2368);
and U3722 (N_3722,N_765,N_2457);
nor U3723 (N_3723,N_547,N_1534);
and U3724 (N_3724,N_2321,N_534);
or U3725 (N_3725,N_993,N_171);
and U3726 (N_3726,N_715,N_484);
and U3727 (N_3727,N_1497,N_299);
nand U3728 (N_3728,N_838,N_2677);
xor U3729 (N_3729,N_1649,N_2383);
or U3730 (N_3730,N_388,N_644);
or U3731 (N_3731,N_1824,N_2668);
nor U3732 (N_3732,N_135,N_2032);
and U3733 (N_3733,N_2954,N_271);
nand U3734 (N_3734,N_2916,N_2258);
and U3735 (N_3735,N_905,N_2703);
nand U3736 (N_3736,N_1430,N_1902);
and U3737 (N_3737,N_982,N_679);
or U3738 (N_3738,N_1009,N_2337);
and U3739 (N_3739,N_2781,N_639);
and U3740 (N_3740,N_2225,N_127);
nor U3741 (N_3741,N_137,N_2116);
or U3742 (N_3742,N_2373,N_724);
and U3743 (N_3743,N_1451,N_1939);
or U3744 (N_3744,N_569,N_465);
nor U3745 (N_3745,N_2358,N_52);
nor U3746 (N_3746,N_1315,N_2968);
nand U3747 (N_3747,N_322,N_2887);
nor U3748 (N_3748,N_500,N_1668);
nand U3749 (N_3749,N_2629,N_1134);
nand U3750 (N_3750,N_1371,N_523);
nor U3751 (N_3751,N_992,N_1750);
nand U3752 (N_3752,N_797,N_1924);
or U3753 (N_3753,N_145,N_2481);
or U3754 (N_3754,N_225,N_740);
nand U3755 (N_3755,N_2678,N_1546);
nand U3756 (N_3756,N_1362,N_837);
nor U3757 (N_3757,N_910,N_979);
nand U3758 (N_3758,N_1006,N_2875);
nand U3759 (N_3759,N_101,N_2255);
and U3760 (N_3760,N_554,N_2768);
nor U3761 (N_3761,N_2359,N_785);
nor U3762 (N_3762,N_634,N_2944);
and U3763 (N_3763,N_512,N_1503);
or U3764 (N_3764,N_973,N_1771);
nor U3765 (N_3765,N_2790,N_960);
nand U3766 (N_3766,N_794,N_359);
and U3767 (N_3767,N_665,N_2873);
nand U3768 (N_3768,N_2848,N_438);
and U3769 (N_3769,N_1728,N_336);
or U3770 (N_3770,N_1098,N_726);
and U3771 (N_3771,N_2259,N_1851);
nand U3772 (N_3772,N_10,N_693);
and U3773 (N_3773,N_520,N_1244);
or U3774 (N_3774,N_1483,N_1011);
or U3775 (N_3775,N_375,N_2949);
and U3776 (N_3776,N_692,N_701);
or U3777 (N_3777,N_906,N_1272);
nand U3778 (N_3778,N_2302,N_1448);
nand U3779 (N_3779,N_397,N_1217);
or U3780 (N_3780,N_2124,N_1407);
and U3781 (N_3781,N_1157,N_475);
nor U3782 (N_3782,N_2347,N_1831);
xnor U3783 (N_3783,N_2607,N_1236);
or U3784 (N_3784,N_2793,N_1130);
nand U3785 (N_3785,N_631,N_162);
nand U3786 (N_3786,N_739,N_831);
or U3787 (N_3787,N_513,N_2159);
and U3788 (N_3788,N_1013,N_401);
and U3789 (N_3789,N_1010,N_1690);
nand U3790 (N_3790,N_2494,N_691);
nand U3791 (N_3791,N_232,N_601);
or U3792 (N_3792,N_640,N_2301);
nor U3793 (N_3793,N_96,N_2220);
nand U3794 (N_3794,N_2286,N_1897);
nand U3795 (N_3795,N_337,N_990);
or U3796 (N_3796,N_2660,N_1232);
and U3797 (N_3797,N_2362,N_2830);
nor U3798 (N_3798,N_603,N_583);
nor U3799 (N_3799,N_1087,N_835);
and U3800 (N_3800,N_755,N_975);
or U3801 (N_3801,N_799,N_2435);
or U3802 (N_3802,N_1715,N_1859);
and U3803 (N_3803,N_2820,N_1536);
nor U3804 (N_3804,N_767,N_17);
or U3805 (N_3805,N_1700,N_1711);
or U3806 (N_3806,N_2561,N_186);
nand U3807 (N_3807,N_1598,N_1517);
nand U3808 (N_3808,N_2157,N_414);
nor U3809 (N_3809,N_2936,N_321);
nor U3810 (N_3810,N_312,N_1154);
nand U3811 (N_3811,N_1705,N_2425);
nor U3812 (N_3812,N_1673,N_1691);
and U3813 (N_3813,N_518,N_149);
nor U3814 (N_3814,N_2715,N_1390);
nand U3815 (N_3815,N_1389,N_998);
nand U3816 (N_3816,N_2671,N_2877);
and U3817 (N_3817,N_2534,N_1021);
xor U3818 (N_3818,N_1175,N_2201);
and U3819 (N_3819,N_1721,N_1382);
and U3820 (N_3820,N_2786,N_1496);
nor U3821 (N_3821,N_349,N_516);
nand U3822 (N_3822,N_528,N_356);
or U3823 (N_3823,N_257,N_1740);
nor U3824 (N_3824,N_163,N_766);
nor U3825 (N_3825,N_2175,N_1219);
nor U3826 (N_3826,N_750,N_1529);
nand U3827 (N_3827,N_374,N_472);
nand U3828 (N_3828,N_2436,N_89);
nor U3829 (N_3829,N_1570,N_2426);
or U3830 (N_3830,N_2648,N_2713);
nor U3831 (N_3831,N_1739,N_2751);
or U3832 (N_3832,N_197,N_1654);
nand U3833 (N_3833,N_1871,N_2314);
nand U3834 (N_3834,N_2316,N_373);
nand U3835 (N_3835,N_86,N_1552);
or U3836 (N_3836,N_621,N_1531);
nor U3837 (N_3837,N_1114,N_476);
nand U3838 (N_3838,N_1209,N_338);
or U3839 (N_3839,N_556,N_303);
or U3840 (N_3840,N_268,N_882);
nor U3841 (N_3841,N_597,N_2187);
and U3842 (N_3842,N_19,N_978);
nor U3843 (N_3843,N_2160,N_985);
nand U3844 (N_3844,N_428,N_2181);
nor U3845 (N_3845,N_23,N_1841);
nor U3846 (N_3846,N_65,N_908);
and U3847 (N_3847,N_800,N_774);
or U3848 (N_3848,N_2886,N_2167);
or U3849 (N_3849,N_2003,N_2521);
and U3850 (N_3850,N_723,N_91);
nand U3851 (N_3851,N_1353,N_1642);
or U3852 (N_3852,N_2078,N_584);
or U3853 (N_3853,N_862,N_2420);
nand U3854 (N_3854,N_1612,N_283);
or U3855 (N_3855,N_947,N_892);
or U3856 (N_3856,N_295,N_987);
nor U3857 (N_3857,N_170,N_67);
nand U3858 (N_3858,N_1822,N_1269);
or U3859 (N_3859,N_1338,N_2372);
or U3860 (N_3860,N_2052,N_115);
or U3861 (N_3861,N_2576,N_1901);
or U3862 (N_3862,N_2216,N_2306);
nand U3863 (N_3863,N_239,N_226);
nand U3864 (N_3864,N_1177,N_2728);
nand U3865 (N_3865,N_1419,N_2437);
nand U3866 (N_3866,N_2290,N_881);
nand U3867 (N_3867,N_1445,N_333);
nor U3868 (N_3868,N_900,N_1659);
nor U3869 (N_3869,N_967,N_567);
or U3870 (N_3870,N_2212,N_661);
nand U3871 (N_3871,N_2566,N_1813);
or U3872 (N_3872,N_1833,N_909);
nor U3873 (N_3873,N_1761,N_817);
nor U3874 (N_3874,N_2150,N_1017);
or U3875 (N_3875,N_136,N_902);
or U3876 (N_3876,N_1091,N_437);
nor U3877 (N_3877,N_1766,N_632);
and U3878 (N_3878,N_1301,N_228);
or U3879 (N_3879,N_332,N_1270);
nand U3880 (N_3880,N_453,N_1305);
nand U3881 (N_3881,N_1826,N_2042);
nor U3882 (N_3882,N_2221,N_1770);
and U3883 (N_3883,N_342,N_2408);
nand U3884 (N_3884,N_2377,N_2536);
nor U3885 (N_3885,N_198,N_1323);
or U3886 (N_3886,N_2525,N_1303);
or U3887 (N_3887,N_2340,N_969);
or U3888 (N_3888,N_495,N_2229);
nand U3889 (N_3889,N_668,N_1801);
or U3890 (N_3890,N_1416,N_1288);
or U3891 (N_3891,N_425,N_2102);
nand U3892 (N_3892,N_1171,N_1410);
and U3893 (N_3893,N_1034,N_2819);
nor U3894 (N_3894,N_2247,N_2313);
and U3895 (N_3895,N_863,N_360);
and U3896 (N_3896,N_2702,N_2929);
or U3897 (N_3897,N_2446,N_580);
nand U3898 (N_3898,N_2628,N_157);
and U3899 (N_3899,N_300,N_2070);
nor U3900 (N_3900,N_2354,N_2195);
and U3901 (N_3901,N_344,N_657);
nor U3902 (N_3902,N_1595,N_493);
or U3903 (N_3903,N_901,N_2636);
nor U3904 (N_3904,N_2054,N_2371);
nand U3905 (N_3905,N_1357,N_1785);
or U3906 (N_3906,N_1674,N_1662);
or U3907 (N_3907,N_1524,N_1031);
and U3908 (N_3908,N_1214,N_316);
nand U3909 (N_3909,N_2631,N_2924);
or U3910 (N_3910,N_836,N_1795);
nor U3911 (N_3911,N_1186,N_1105);
and U3912 (N_3912,N_2193,N_2829);
or U3913 (N_3913,N_1238,N_325);
nor U3914 (N_3914,N_81,N_361);
nor U3915 (N_3915,N_1656,N_2097);
xnor U3916 (N_3916,N_1823,N_2395);
nor U3917 (N_3917,N_1938,N_2656);
nand U3918 (N_3918,N_1518,N_2114);
nand U3919 (N_3919,N_296,N_2767);
or U3920 (N_3920,N_1845,N_497);
nor U3921 (N_3921,N_2724,N_14);
and U3922 (N_3922,N_1499,N_1984);
or U3923 (N_3923,N_2355,N_2411);
nand U3924 (N_3924,N_2083,N_1081);
nor U3925 (N_3925,N_326,N_2246);
or U3926 (N_3926,N_674,N_29);
nor U3927 (N_3927,N_278,N_2326);
or U3928 (N_3928,N_1107,N_132);
nand U3929 (N_3929,N_2567,N_1433);
or U3930 (N_3930,N_2905,N_1844);
or U3931 (N_3931,N_2550,N_609);
nor U3932 (N_3932,N_2021,N_1953);
nand U3933 (N_3933,N_1404,N_2782);
and U3934 (N_3934,N_1954,N_382);
or U3935 (N_3935,N_2976,N_2236);
nand U3936 (N_3936,N_2320,N_1393);
nand U3937 (N_3937,N_1904,N_1545);
or U3938 (N_3938,N_2811,N_763);
nand U3939 (N_3939,N_347,N_894);
or U3940 (N_3940,N_2194,N_2051);
nor U3941 (N_3941,N_1501,N_1862);
and U3942 (N_3942,N_2667,N_1327);
or U3943 (N_3943,N_1738,N_743);
and U3944 (N_3944,N_2712,N_1298);
or U3945 (N_3945,N_1886,N_890);
or U3946 (N_3946,N_2740,N_2931);
or U3947 (N_3947,N_1317,N_1864);
xor U3948 (N_3948,N_185,N_1439);
or U3949 (N_3949,N_2011,N_389);
nand U3950 (N_3950,N_400,N_2089);
nor U3951 (N_3951,N_348,N_1444);
or U3952 (N_3952,N_1147,N_2675);
nor U3953 (N_3953,N_77,N_2909);
or U3954 (N_3954,N_2508,N_307);
and U3955 (N_3955,N_719,N_134);
or U3956 (N_3956,N_1758,N_1877);
nand U3957 (N_3957,N_2669,N_2770);
and U3958 (N_3958,N_1278,N_1577);
nand U3959 (N_3959,N_1078,N_2110);
and U3960 (N_3960,N_173,N_1030);
nand U3961 (N_3961,N_1207,N_369);
nor U3962 (N_3962,N_2570,N_930);
nor U3963 (N_3963,N_1431,N_1181);
nor U3964 (N_3964,N_565,N_142);
nand U3965 (N_3965,N_2784,N_620);
nand U3966 (N_3966,N_355,N_879);
or U3967 (N_3967,N_1805,N_2680);
or U3968 (N_3968,N_1685,N_1412);
nand U3969 (N_3969,N_1850,N_561);
nor U3970 (N_3970,N_459,N_430);
or U3971 (N_3971,N_1819,N_1170);
or U3972 (N_3972,N_2592,N_2651);
nor U3973 (N_3973,N_590,N_789);
and U3974 (N_3974,N_2144,N_11);
nor U3975 (N_3975,N_1791,N_2230);
and U3976 (N_3976,N_1964,N_1152);
nand U3977 (N_3977,N_2495,N_2785);
nor U3978 (N_3978,N_1985,N_2920);
nand U3979 (N_3979,N_235,N_492);
or U3980 (N_3980,N_1669,N_1733);
nand U3981 (N_3981,N_2343,N_2653);
and U3982 (N_3982,N_1200,N_237);
nor U3983 (N_3983,N_2870,N_2806);
and U3984 (N_3984,N_2973,N_934);
or U3985 (N_3985,N_2562,N_913);
and U3986 (N_3986,N_1574,N_1340);
nand U3987 (N_3987,N_1491,N_1068);
or U3988 (N_3988,N_1352,N_1201);
nand U3989 (N_3989,N_1838,N_1631);
or U3990 (N_3990,N_219,N_1625);
and U3991 (N_3991,N_1637,N_2580);
or U3992 (N_3992,N_1252,N_218);
nand U3993 (N_3993,N_147,N_895);
and U3994 (N_3994,N_1023,N_2012);
and U3995 (N_3995,N_1742,N_483);
and U3996 (N_3996,N_130,N_460);
nor U3997 (N_3997,N_143,N_2854);
or U3998 (N_3998,N_2979,N_587);
nand U3999 (N_3999,N_2333,N_685);
or U4000 (N_4000,N_1486,N_1849);
nand U4001 (N_4001,N_1732,N_2506);
nor U4002 (N_4002,N_2860,N_1589);
and U4003 (N_4003,N_1077,N_2934);
nor U4004 (N_4004,N_941,N_1802);
and U4005 (N_4005,N_1271,N_1650);
and U4006 (N_4006,N_1955,N_2825);
and U4007 (N_4007,N_1347,N_2432);
and U4008 (N_4008,N_1727,N_2252);
and U4009 (N_4009,N_596,N_2632);
and U4010 (N_4010,N_877,N_970);
or U4011 (N_4011,N_2237,N_545);
nor U4012 (N_4012,N_2686,N_339);
nand U4013 (N_4013,N_1263,N_2043);
nor U4014 (N_4014,N_1089,N_1246);
and U4015 (N_4015,N_2602,N_1998);
or U4016 (N_4016,N_1474,N_2293);
nor U4017 (N_4017,N_2862,N_2389);
nand U4018 (N_4018,N_2223,N_1689);
nor U4019 (N_4019,N_2590,N_2741);
nor U4020 (N_4020,N_2310,N_2019);
and U4021 (N_4021,N_2813,N_2022);
xor U4022 (N_4022,N_2461,N_2655);
nand U4023 (N_4023,N_2267,N_898);
nor U4024 (N_4024,N_2168,N_1230);
or U4025 (N_4025,N_2545,N_2581);
and U4026 (N_4026,N_2634,N_1466);
nand U4027 (N_4027,N_2888,N_858);
or U4028 (N_4028,N_141,N_1000);
or U4029 (N_4029,N_208,N_2867);
nand U4030 (N_4030,N_2972,N_1176);
nor U4031 (N_4031,N_1568,N_1614);
or U4032 (N_4032,N_2872,N_1697);
and U4033 (N_4033,N_2919,N_897);
nor U4034 (N_4034,N_570,N_2120);
or U4035 (N_4035,N_849,N_1919);
and U4036 (N_4036,N_2101,N_2864);
nand U4037 (N_4037,N_1464,N_1815);
nand U4038 (N_4038,N_2338,N_2760);
or U4039 (N_4039,N_735,N_2391);
nand U4040 (N_4040,N_1102,N_2961);
nand U4041 (N_4041,N_2401,N_2169);
or U4042 (N_4042,N_2251,N_1314);
and U4043 (N_4043,N_1426,N_2405);
or U4044 (N_4044,N_1463,N_1830);
nand U4045 (N_4045,N_2564,N_405);
nor U4046 (N_4046,N_324,N_776);
or U4047 (N_4047,N_255,N_2460);
nor U4048 (N_4048,N_1297,N_1712);
and U4049 (N_4049,N_2518,N_2930);
nand U4050 (N_4050,N_2200,N_1039);
nand U4051 (N_4051,N_1620,N_780);
and U4052 (N_4052,N_395,N_353);
or U4053 (N_4053,N_1049,N_380);
nor U4054 (N_4054,N_201,N_781);
nor U4055 (N_4055,N_2210,N_2488);
nand U4056 (N_4056,N_2735,N_1343);
xor U4057 (N_4057,N_2527,N_1535);
nor U4058 (N_4058,N_2206,N_98);
or U4059 (N_4059,N_320,N_1976);
and U4060 (N_4060,N_643,N_623);
nand U4061 (N_4061,N_2601,N_133);
nor U4062 (N_4062,N_543,N_499);
nand U4063 (N_4063,N_2993,N_1212);
or U4064 (N_4064,N_1829,N_385);
nand U4065 (N_4065,N_485,N_1977);
nand U4066 (N_4066,N_2803,N_2260);
and U4067 (N_4067,N_1245,N_816);
nand U4068 (N_4068,N_1424,N_1275);
or U4069 (N_4069,N_1843,N_2231);
nor U4070 (N_4070,N_752,N_1812);
and U4071 (N_4071,N_1397,N_1793);
and U4072 (N_4072,N_1061,N_1364);
nor U4073 (N_4073,N_1441,N_1688);
and U4074 (N_4074,N_447,N_104);
and U4075 (N_4075,N_1932,N_586);
nand U4076 (N_4076,N_2822,N_2090);
or U4077 (N_4077,N_997,N_2452);
nor U4078 (N_4078,N_2925,N_2270);
or U4079 (N_4079,N_1814,N_1982);
and U4080 (N_4080,N_802,N_1391);
or U4081 (N_4081,N_2685,N_188);
xor U4082 (N_4082,N_2462,N_1224);
and U4083 (N_4083,N_804,N_3);
nand U4084 (N_4084,N_1556,N_1456);
or U4085 (N_4085,N_2711,N_2093);
nand U4086 (N_4086,N_707,N_1119);
or U4087 (N_4087,N_2505,N_1765);
or U4088 (N_4088,N_857,N_2466);
nand U4089 (N_4089,N_21,N_128);
and U4090 (N_4090,N_1149,N_1638);
nand U4091 (N_4091,N_2664,N_2736);
or U4092 (N_4092,N_123,N_2774);
and U4093 (N_4093,N_1342,N_2025);
nor U4094 (N_4094,N_1635,N_223);
and U4095 (N_4095,N_2988,N_83);
nand U4096 (N_4096,N_1437,N_1584);
nand U4097 (N_4097,N_1519,N_253);
or U4098 (N_4098,N_641,N_2738);
and U4099 (N_4099,N_1627,N_2244);
nor U4100 (N_4100,N_690,N_522);
nand U4101 (N_4101,N_2646,N_662);
nand U4102 (N_4102,N_2588,N_2778);
xor U4103 (N_4103,N_242,N_1875);
nor U4104 (N_4104,N_51,N_1895);
nand U4105 (N_4105,N_263,N_2048);
and U4106 (N_4106,N_306,N_1016);
or U4107 (N_4107,N_923,N_2178);
or U4108 (N_4108,N_759,N_2838);
and U4109 (N_4109,N_604,N_2013);
nor U4110 (N_4110,N_57,N_2720);
nand U4111 (N_4111,N_1406,N_1085);
and U4112 (N_4112,N_826,N_2937);
nand U4113 (N_4113,N_424,N_1527);
or U4114 (N_4114,N_1405,N_2729);
nand U4115 (N_4115,N_58,N_7);
and U4116 (N_4116,N_1428,N_652);
and U4117 (N_4117,N_529,N_1878);
and U4118 (N_4118,N_1693,N_1062);
nor U4119 (N_4119,N_524,N_262);
nor U4120 (N_4120,N_116,N_175);
nor U4121 (N_4121,N_1060,N_2865);
or U4122 (N_4122,N_1696,N_827);
and U4123 (N_4123,N_2922,N_2351);
nand U4124 (N_4124,N_884,N_426);
nand U4125 (N_4125,N_642,N_2141);
and U4126 (N_4126,N_622,N_2331);
or U4127 (N_4127,N_2619,N_2198);
nand U4128 (N_4128,N_1056,N_284);
or U4129 (N_4129,N_1790,N_1893);
and U4130 (N_4130,N_1972,N_813);
nor U4131 (N_4131,N_309,N_2345);
or U4132 (N_4132,N_2381,N_2219);
nor U4133 (N_4133,N_146,N_1223);
and U4134 (N_4134,N_1088,N_1180);
nand U4135 (N_4135,N_183,N_988);
nor U4136 (N_4136,N_2701,N_2161);
nor U4137 (N_4137,N_1784,N_588);
nor U4138 (N_4138,N_2497,N_2268);
nor U4139 (N_4139,N_1022,N_2551);
and U4140 (N_4140,N_1249,N_1360);
or U4141 (N_4141,N_2857,N_899);
nand U4142 (N_4142,N_2232,N_1458);
nor U4143 (N_4143,N_1557,N_1235);
nor U4144 (N_4144,N_1282,N_2130);
nand U4145 (N_4145,N_1358,N_2370);
nand U4146 (N_4146,N_1796,N_2406);
nor U4147 (N_4147,N_866,N_2539);
nor U4148 (N_4148,N_2473,N_1926);
nor U4149 (N_4149,N_1027,N_301);
nand U4150 (N_4150,N_1846,N_1309);
or U4151 (N_4151,N_140,N_542);
and U4152 (N_4152,N_1139,N_1523);
and U4153 (N_4153,N_1106,N_1599);
nor U4154 (N_4154,N_925,N_1494);
or U4155 (N_4155,N_2365,N_1005);
nand U4156 (N_4156,N_1986,N_2585);
nand U4157 (N_4157,N_2787,N_180);
nand U4158 (N_4158,N_1613,N_1966);
and U4159 (N_4159,N_2896,N_184);
nor U4160 (N_4160,N_1198,N_2617);
nand U4161 (N_4161,N_1541,N_160);
nor U4162 (N_4162,N_2339,N_2177);
and U4163 (N_4163,N_1532,N_2791);
nor U4164 (N_4164,N_2624,N_2464);
and U4165 (N_4165,N_2060,N_80);
or U4166 (N_4166,N_407,N_713);
or U4167 (N_4167,N_2020,N_1555);
nor U4168 (N_4168,N_1240,N_446);
or U4169 (N_4169,N_1999,N_1891);
or U4170 (N_4170,N_1356,N_74);
and U4171 (N_4171,N_187,N_331);
nor U4172 (N_4172,N_2765,N_234);
and U4173 (N_4173,N_506,N_1528);
nor U4174 (N_4174,N_1370,N_1827);
nand U4175 (N_4175,N_1744,N_2759);
nand U4176 (N_4176,N_1702,N_398);
nor U4177 (N_4177,N_2375,N_791);
nand U4178 (N_4178,N_1321,N_406);
or U4179 (N_4179,N_1325,N_514);
xnor U4180 (N_4180,N_806,N_2795);
nand U4181 (N_4181,N_2180,N_277);
nand U4182 (N_4182,N_279,N_419);
nand U4183 (N_4183,N_153,N_1554);
or U4184 (N_4184,N_217,N_2717);
nand U4185 (N_4185,N_864,N_477);
or U4186 (N_4186,N_205,N_2523);
or U4187 (N_4187,N_2369,N_1561);
nor U4188 (N_4188,N_2844,N_2986);
and U4189 (N_4189,N_790,N_1991);
nand U4190 (N_4190,N_2196,N_1035);
and U4191 (N_4191,N_351,N_1741);
nand U4192 (N_4192,N_1368,N_1914);
and U4193 (N_4193,N_165,N_2969);
nor U4194 (N_4194,N_1421,N_572);
or U4195 (N_4195,N_1138,N_694);
and U4196 (N_4196,N_2026,N_1349);
nand U4197 (N_4197,N_1931,N_1398);
and U4198 (N_4198,N_907,N_1403);
nand U4199 (N_4199,N_1196,N_2164);
nand U4200 (N_4200,N_1952,N_1339);
and U4201 (N_4201,N_2861,N_808);
nand U4202 (N_4202,N_1345,N_536);
or U4203 (N_4203,N_399,N_328);
and U4204 (N_4204,N_304,N_2556);
or U4205 (N_4205,N_792,N_1978);
nand U4206 (N_4206,N_963,N_2514);
nand U4207 (N_4207,N_758,N_63);
nand U4208 (N_4208,N_41,N_1018);
and U4209 (N_4209,N_624,N_2532);
nor U4210 (N_4210,N_736,N_929);
or U4211 (N_4211,N_87,N_402);
and U4212 (N_4212,N_364,N_1803);
nor U4213 (N_4213,N_1384,N_474);
or U4214 (N_4214,N_341,N_539);
nand U4215 (N_4215,N_455,N_2265);
or U4216 (N_4216,N_756,N_317);
and U4217 (N_4217,N_1048,N_50);
and U4218 (N_4218,N_2485,N_315);
nor U4219 (N_4219,N_2776,N_999);
nand U4220 (N_4220,N_2207,N_2463);
or U4221 (N_4221,N_1853,N_1539);
and U4222 (N_4222,N_2600,N_697);
nand U4223 (N_4223,N_1997,N_2384);
nand U4224 (N_4224,N_559,N_525);
and U4225 (N_4225,N_2946,N_2828);
or U4226 (N_4226,N_310,N_2199);
or U4227 (N_4227,N_2788,N_1917);
nand U4228 (N_4228,N_2357,N_1100);
or U4229 (N_4229,N_1933,N_254);
or U4230 (N_4230,N_872,N_2687);
or U4231 (N_4231,N_2203,N_935);
nand U4232 (N_4232,N_953,N_1066);
nor U4233 (N_4233,N_1745,N_611);
or U4234 (N_4234,N_1937,N_2431);
or U4235 (N_4235,N_511,N_1621);
nand U4236 (N_4236,N_2121,N_1488);
or U4237 (N_4237,N_282,N_1870);
nand U4238 (N_4238,N_2096,N_917);
or U4239 (N_4239,N_2280,N_1480);
and U4240 (N_4240,N_1522,N_2906);
nand U4241 (N_4241,N_281,N_532);
nor U4242 (N_4242,N_1828,N_1792);
nor U4243 (N_4243,N_13,N_2652);
and U4244 (N_4244,N_2985,N_951);
and U4245 (N_4245,N_4,N_169);
nor U4246 (N_4246,N_238,N_429);
nand U4247 (N_4247,N_2074,N_2145);
nor U4248 (N_4248,N_1090,N_2792);
or U4249 (N_4249,N_2522,N_1645);
nand U4250 (N_4250,N_2467,N_2056);
or U4251 (N_4251,N_1329,N_1553);
and U4252 (N_4252,N_1854,N_582);
and U4253 (N_4253,N_1164,N_2284);
and U4254 (N_4254,N_2421,N_1038);
and U4255 (N_4255,N_1811,N_1874);
and U4256 (N_4256,N_555,N_784);
nand U4257 (N_4257,N_1730,N_625);
or U4258 (N_4258,N_686,N_1095);
nor U4259 (N_4259,N_1287,N_2084);
or U4260 (N_4260,N_2722,N_1376);
and U4261 (N_4261,N_2807,N_1708);
nand U4262 (N_4262,N_2571,N_2062);
nand U4263 (N_4263,N_571,N_1148);
nor U4264 (N_4264,N_2709,N_1073);
and U4265 (N_4265,N_2583,N_376);
nor U4266 (N_4266,N_1346,N_2307);
or U4267 (N_4267,N_2133,N_1563);
nand U4268 (N_4268,N_1617,N_1947);
nor U4269 (N_4269,N_658,N_245);
nor U4270 (N_4270,N_2665,N_648);
nand U4271 (N_4271,N_1302,N_2300);
nand U4272 (N_4272,N_289,N_2107);
or U4273 (N_4273,N_179,N_2744);
and U4274 (N_4274,N_2079,N_1268);
and U4275 (N_4275,N_2186,N_1619);
and U4276 (N_4276,N_2069,N_2095);
nand U4277 (N_4277,N_1036,N_507);
nor U4278 (N_4278,N_1582,N_2344);
and U4279 (N_4279,N_2087,N_856);
nand U4280 (N_4280,N_1096,N_2204);
nand U4281 (N_4281,N_1701,N_1434);
nor U4282 (N_4282,N_2253,N_1709);
nor U4283 (N_4283,N_1647,N_1425);
nand U4284 (N_4284,N_1665,N_1388);
and U4285 (N_4285,N_830,N_327);
and U4286 (N_4286,N_2577,N_578);
nand U4287 (N_4287,N_563,N_1852);
nor U4288 (N_4288,N_2001,N_2140);
or U4289 (N_4289,N_2840,N_2063);
nor U4290 (N_4290,N_423,N_606);
nor U4291 (N_4291,N_965,N_370);
and U4292 (N_4292,N_1723,N_2176);
nor U4293 (N_4293,N_441,N_433);
and U4294 (N_4294,N_28,N_1876);
nand U4295 (N_4295,N_454,N_466);
or U4296 (N_4296,N_1337,N_79);
xor U4297 (N_4297,N_102,N_286);
nor U4298 (N_4298,N_2881,N_298);
nor U4299 (N_4299,N_1881,N_2393);
nand U4300 (N_4300,N_1247,N_2547);
and U4301 (N_4301,N_394,N_330);
and U4302 (N_4302,N_654,N_675);
or U4303 (N_4303,N_1103,N_2746);
nor U4304 (N_4304,N_2455,N_2192);
nand U4305 (N_4305,N_1963,N_878);
or U4306 (N_4306,N_61,N_1725);
nand U4307 (N_4307,N_2639,N_549);
or U4308 (N_4308,N_2614,N_1706);
and U4309 (N_4309,N_2031,N_2385);
and U4310 (N_4310,N_1427,N_2597);
nand U4311 (N_4311,N_820,N_345);
nor U4312 (N_4312,N_871,N_2311);
or U4313 (N_4313,N_2271,N_1734);
nand U4314 (N_4314,N_2010,N_1414);
nor U4315 (N_4315,N_2721,N_323);
or U4316 (N_4316,N_222,N_1604);
nand U4317 (N_4317,N_1581,N_2205);
nand U4318 (N_4318,N_48,N_1836);
and U4319 (N_4319,N_1867,N_2249);
nand U4320 (N_4320,N_1622,N_591);
nand U4321 (N_4321,N_2755,N_2719);
nand U4322 (N_4322,N_2897,N_2989);
or U4323 (N_4323,N_1989,N_2723);
and U4324 (N_4324,N_1704,N_932);
nand U4325 (N_4325,N_753,N_2538);
nand U4326 (N_4326,N_1855,N_2029);
or U4327 (N_4327,N_1324,N_1550);
nand U4328 (N_4328,N_1101,N_2676);
and U4329 (N_4329,N_1233,N_922);
nor U4330 (N_4330,N_55,N_22);
nor U4331 (N_4331,N_1178,N_2050);
or U4332 (N_4332,N_383,N_1310);
and U4333 (N_4333,N_748,N_2118);
nand U4334 (N_4334,N_1983,N_734);
nor U4335 (N_4335,N_2256,N_2049);
xor U4336 (N_4336,N_1682,N_2823);
nand U4337 (N_4337,N_1694,N_1567);
or U4338 (N_4338,N_2780,N_1478);
nor U4339 (N_4339,N_1075,N_1779);
or U4340 (N_4340,N_2496,N_942);
nor U4341 (N_4341,N_1773,N_2615);
nand U4342 (N_4342,N_412,N_164);
xor U4343 (N_4343,N_2923,N_468);
or U4344 (N_4344,N_2308,N_873);
or U4345 (N_4345,N_381,N_920);
and U4346 (N_4346,N_2817,N_2894);
xnor U4347 (N_4347,N_2336,N_2730);
and U4348 (N_4348,N_470,N_1168);
nand U4349 (N_4349,N_1692,N_1980);
and U4350 (N_4350,N_2966,N_2643);
nor U4351 (N_4351,N_2964,N_889);
nand U4352 (N_4352,N_768,N_2800);
or U4353 (N_4353,N_2535,N_1777);
nor U4354 (N_4354,N_241,N_977);
and U4355 (N_4355,N_2448,N_1569);
or U4356 (N_4356,N_60,N_828);
and U4357 (N_4357,N_34,N_1907);
or U4358 (N_4358,N_1173,N_33);
and U4359 (N_4359,N_1257,N_2627);
and U4360 (N_4360,N_1959,N_1588);
nand U4361 (N_4361,N_1465,N_1059);
xor U4362 (N_4362,N_1809,N_669);
nand U4363 (N_4363,N_1834,N_1786);
and U4364 (N_4364,N_618,N_1748);
or U4365 (N_4365,N_1988,N_1191);
or U4366 (N_4366,N_2990,N_2018);
nand U4367 (N_4367,N_2173,N_1135);
and U4368 (N_4368,N_1153,N_1558);
or U4369 (N_4369,N_1994,N_651);
xnor U4370 (N_4370,N_251,N_964);
nand U4371 (N_4371,N_2821,N_2298);
nand U4372 (N_4372,N_1585,N_1866);
and U4373 (N_4373,N_1565,N_2960);
nand U4374 (N_4374,N_2036,N_1279);
and U4375 (N_4375,N_1973,N_595);
or U4376 (N_4376,N_851,N_725);
nor U4377 (N_4377,N_335,N_272);
nand U4378 (N_4378,N_2183,N_2841);
or U4379 (N_4379,N_2696,N_2098);
and U4380 (N_4380,N_1835,N_2294);
nand U4381 (N_4381,N_2689,N_124);
and U4382 (N_4382,N_646,N_2404);
nor U4383 (N_4383,N_2332,N_2707);
and U4384 (N_4384,N_2605,N_2798);
or U4385 (N_4385,N_1350,N_2595);
nor U4386 (N_4386,N_2903,N_2072);
nor U4387 (N_4387,N_716,N_2616);
nor U4388 (N_4388,N_983,N_1304);
and U4389 (N_4389,N_875,N_2504);
or U4390 (N_4390,N_2808,N_2152);
or U4391 (N_4391,N_2812,N_915);
or U4392 (N_4392,N_467,N_946);
nand U4393 (N_4393,N_2849,N_2119);
nand U4394 (N_4394,N_2834,N_1386);
nor U4395 (N_4395,N_1076,N_855);
nor U4396 (N_4396,N_2796,N_110);
nand U4397 (N_4397,N_2349,N_1300);
nor U4398 (N_4398,N_708,N_2040);
nor U4399 (N_4399,N_1724,N_2827);
or U4400 (N_4400,N_2325,N_2428);
nand U4401 (N_4401,N_2610,N_860);
or U4402 (N_4402,N_214,N_627);
nor U4403 (N_4403,N_1861,N_2847);
nand U4404 (N_4404,N_26,N_1591);
and U4405 (N_4405,N_2108,N_2757);
nor U4406 (N_4406,N_2304,N_2883);
nand U4407 (N_4407,N_2392,N_2835);
or U4408 (N_4408,N_974,N_1677);
or U4409 (N_4409,N_1046,N_924);
nand U4410 (N_4410,N_2557,N_2443);
nor U4411 (N_4411,N_2458,N_1086);
nand U4412 (N_4412,N_420,N_706);
and U4413 (N_4413,N_2809,N_1172);
nand U4414 (N_4414,N_2764,N_1446);
nor U4415 (N_4415,N_721,N_638);
or U4416 (N_4416,N_1128,N_952);
nor U4417 (N_4417,N_168,N_1944);
and U4418 (N_4418,N_2262,N_1);
or U4419 (N_4419,N_2754,N_714);
and U4420 (N_4420,N_1879,N_2418);
nor U4421 (N_4421,N_1110,N_1256);
or U4422 (N_4422,N_805,N_2076);
or U4423 (N_4423,N_496,N_35);
nor U4424 (N_4424,N_821,N_633);
nand U4425 (N_4425,N_1204,N_775);
nor U4426 (N_4426,N_1821,N_27);
nor U4427 (N_4427,N_1710,N_1504);
nand U4428 (N_4428,N_416,N_148);
and U4429 (N_4429,N_53,N_1903);
and U4430 (N_4430,N_2582,N_2732);
nor U4431 (N_4431,N_1166,N_2526);
and U4432 (N_4432,N_1449,N_2479);
or U4433 (N_4433,N_1564,N_252);
or U4434 (N_4434,N_2996,N_1945);
or U4435 (N_4435,N_1065,N_243);
nor U4436 (N_4436,N_1120,N_1216);
nor U4437 (N_4437,N_2179,N_1045);
nand U4438 (N_4438,N_1116,N_2016);
nand U4439 (N_4439,N_846,N_2166);
and U4440 (N_4440,N_1960,N_504);
or U4441 (N_4441,N_777,N_1192);
or U4442 (N_4442,N_1856,N_1259);
nor U4443 (N_4443,N_2708,N_607);
or U4444 (N_4444,N_1380,N_710);
nor U4445 (N_4445,N_2783,N_1628);
nand U4446 (N_4446,N_1290,N_2975);
and U4447 (N_4447,N_1922,N_1145);
nand U4448 (N_4448,N_39,N_503);
nor U4449 (N_4449,N_1990,N_1754);
and U4450 (N_4450,N_2981,N_1646);
nand U4451 (N_4451,N_876,N_1189);
and U4452 (N_4452,N_711,N_2900);
or U4453 (N_4453,N_1097,N_1020);
nor U4454 (N_4454,N_1498,N_1468);
nor U4455 (N_4455,N_1015,N_379);
nor U4456 (N_4456,N_1051,N_2868);
and U4457 (N_4457,N_2608,N_2858);
nand U4458 (N_4458,N_1590,N_2105);
nor U4459 (N_4459,N_1381,N_386);
nand U4460 (N_4460,N_2134,N_2367);
or U4461 (N_4461,N_2281,N_2000);
and U4462 (N_4462,N_2480,N_1241);
and U4463 (N_4463,N_1655,N_2991);
and U4464 (N_4464,N_2533,N_2593);
nor U4465 (N_4465,N_2941,N_1184);
nor U4466 (N_4466,N_2716,N_1484);
nor U4467 (N_4467,N_1248,N_1210);
or U4468 (N_4468,N_1760,N_2928);
nand U4469 (N_4469,N_1502,N_2295);
and U4470 (N_4470,N_1951,N_1025);
or U4471 (N_4471,N_1808,N_885);
nor U4472 (N_4472,N_787,N_893);
or U4473 (N_4473,N_220,N_2824);
nor U4474 (N_4474,N_318,N_844);
nand U4475 (N_4475,N_2638,N_636);
nand U4476 (N_4476,N_630,N_1873);
or U4477 (N_4477,N_2388,N_2453);
nor U4478 (N_4478,N_704,N_1664);
or U4479 (N_4479,N_745,N_1229);
nand U4480 (N_4480,N_2846,N_2630);
or U4481 (N_4481,N_593,N_2921);
and U4482 (N_4482,N_1124,N_1571);
nand U4483 (N_4483,N_1735,N_1962);
nor U4484 (N_4484,N_700,N_82);
nand U4485 (N_4485,N_1615,N_1041);
and U4486 (N_4486,N_1950,N_1125);
nor U4487 (N_4487,N_2579,N_1974);
nor U4488 (N_4488,N_2402,N_1208);
and U4489 (N_4489,N_1485,N_2663);
nand U4490 (N_4490,N_575,N_2718);
and U4491 (N_4491,N_2901,N_2100);
or U4492 (N_4492,N_2469,N_2520);
or U4493 (N_4493,N_1578,N_1366);
nand U4494 (N_4494,N_1857,N_1736);
nor U4495 (N_4495,N_738,N_1093);
or U4496 (N_4496,N_2606,N_1260);
and U4497 (N_4497,N_491,N_2142);
nand U4498 (N_4498,N_1266,N_105);
nor U4499 (N_4499,N_2468,N_94);
and U4500 (N_4500,N_355,N_1381);
nand U4501 (N_4501,N_670,N_185);
or U4502 (N_4502,N_2279,N_2550);
nand U4503 (N_4503,N_1562,N_2719);
nand U4504 (N_4504,N_2269,N_2835);
or U4505 (N_4505,N_2794,N_46);
nand U4506 (N_4506,N_2172,N_507);
nor U4507 (N_4507,N_1742,N_2567);
nor U4508 (N_4508,N_2274,N_315);
and U4509 (N_4509,N_1301,N_1002);
or U4510 (N_4510,N_601,N_150);
or U4511 (N_4511,N_2148,N_527);
nand U4512 (N_4512,N_1094,N_2518);
and U4513 (N_4513,N_347,N_2870);
or U4514 (N_4514,N_1386,N_166);
and U4515 (N_4515,N_371,N_220);
or U4516 (N_4516,N_2166,N_1195);
nand U4517 (N_4517,N_1478,N_933);
or U4518 (N_4518,N_2935,N_1055);
xnor U4519 (N_4519,N_2274,N_642);
or U4520 (N_4520,N_896,N_2377);
nor U4521 (N_4521,N_353,N_733);
nand U4522 (N_4522,N_1026,N_872);
nand U4523 (N_4523,N_1449,N_180);
and U4524 (N_4524,N_1168,N_490);
and U4525 (N_4525,N_160,N_1350);
or U4526 (N_4526,N_1264,N_25);
nand U4527 (N_4527,N_2831,N_2852);
and U4528 (N_4528,N_1496,N_1771);
nor U4529 (N_4529,N_690,N_2475);
or U4530 (N_4530,N_178,N_2543);
or U4531 (N_4531,N_2424,N_2460);
and U4532 (N_4532,N_1916,N_2903);
or U4533 (N_4533,N_1346,N_2013);
or U4534 (N_4534,N_1967,N_650);
nor U4535 (N_4535,N_1258,N_1829);
nor U4536 (N_4536,N_2316,N_132);
and U4537 (N_4537,N_987,N_1477);
nor U4538 (N_4538,N_1059,N_2303);
or U4539 (N_4539,N_367,N_2781);
or U4540 (N_4540,N_2234,N_157);
and U4541 (N_4541,N_1586,N_2594);
and U4542 (N_4542,N_1756,N_2600);
nand U4543 (N_4543,N_1344,N_1531);
and U4544 (N_4544,N_604,N_1449);
and U4545 (N_4545,N_1468,N_518);
and U4546 (N_4546,N_966,N_2610);
or U4547 (N_4547,N_671,N_1985);
nand U4548 (N_4548,N_2056,N_800);
nor U4549 (N_4549,N_614,N_836);
nand U4550 (N_4550,N_1589,N_2164);
and U4551 (N_4551,N_2501,N_524);
and U4552 (N_4552,N_1,N_2813);
or U4553 (N_4553,N_1260,N_2180);
nand U4554 (N_4554,N_1589,N_2825);
or U4555 (N_4555,N_1714,N_1051);
nand U4556 (N_4556,N_1356,N_449);
nand U4557 (N_4557,N_1093,N_902);
and U4558 (N_4558,N_2652,N_2066);
and U4559 (N_4559,N_1990,N_1901);
nand U4560 (N_4560,N_2304,N_2170);
or U4561 (N_4561,N_2140,N_1360);
or U4562 (N_4562,N_547,N_2822);
nand U4563 (N_4563,N_2588,N_801);
or U4564 (N_4564,N_252,N_207);
or U4565 (N_4565,N_1410,N_349);
or U4566 (N_4566,N_2515,N_1455);
nor U4567 (N_4567,N_2265,N_845);
nand U4568 (N_4568,N_905,N_1876);
nor U4569 (N_4569,N_45,N_81);
and U4570 (N_4570,N_1330,N_2699);
nor U4571 (N_4571,N_2770,N_2992);
nor U4572 (N_4572,N_362,N_439);
nand U4573 (N_4573,N_1910,N_2853);
and U4574 (N_4574,N_2552,N_716);
nand U4575 (N_4575,N_2002,N_1842);
nand U4576 (N_4576,N_962,N_2377);
and U4577 (N_4577,N_1417,N_2065);
and U4578 (N_4578,N_103,N_2758);
or U4579 (N_4579,N_771,N_1926);
and U4580 (N_4580,N_2582,N_616);
xor U4581 (N_4581,N_1442,N_323);
nand U4582 (N_4582,N_824,N_621);
and U4583 (N_4583,N_2102,N_832);
nor U4584 (N_4584,N_2171,N_2049);
nand U4585 (N_4585,N_1693,N_254);
nand U4586 (N_4586,N_2631,N_51);
or U4587 (N_4587,N_2002,N_1110);
nor U4588 (N_4588,N_1425,N_2359);
nand U4589 (N_4589,N_2836,N_872);
nor U4590 (N_4590,N_2028,N_519);
and U4591 (N_4591,N_648,N_2516);
and U4592 (N_4592,N_960,N_281);
nor U4593 (N_4593,N_2785,N_2888);
nor U4594 (N_4594,N_2189,N_161);
nand U4595 (N_4595,N_1204,N_1532);
and U4596 (N_4596,N_72,N_972);
nand U4597 (N_4597,N_2282,N_288);
nor U4598 (N_4598,N_1219,N_1804);
nor U4599 (N_4599,N_2214,N_555);
or U4600 (N_4600,N_2291,N_1916);
nand U4601 (N_4601,N_1884,N_1053);
nor U4602 (N_4602,N_2359,N_1107);
and U4603 (N_4603,N_1310,N_2948);
nand U4604 (N_4604,N_410,N_1535);
or U4605 (N_4605,N_930,N_598);
and U4606 (N_4606,N_1031,N_1654);
nand U4607 (N_4607,N_300,N_1685);
nor U4608 (N_4608,N_203,N_2241);
nand U4609 (N_4609,N_1446,N_2083);
and U4610 (N_4610,N_911,N_1804);
nand U4611 (N_4611,N_445,N_1064);
nor U4612 (N_4612,N_2255,N_1500);
and U4613 (N_4613,N_2628,N_171);
nand U4614 (N_4614,N_1920,N_46);
nand U4615 (N_4615,N_691,N_1560);
and U4616 (N_4616,N_1217,N_1849);
nand U4617 (N_4617,N_1074,N_701);
and U4618 (N_4618,N_327,N_2054);
nand U4619 (N_4619,N_1163,N_1847);
nor U4620 (N_4620,N_15,N_1621);
nor U4621 (N_4621,N_2713,N_848);
or U4622 (N_4622,N_528,N_1436);
or U4623 (N_4623,N_2276,N_2458);
nor U4624 (N_4624,N_1603,N_2775);
nand U4625 (N_4625,N_1477,N_2940);
or U4626 (N_4626,N_761,N_241);
and U4627 (N_4627,N_2352,N_2331);
and U4628 (N_4628,N_1765,N_834);
nor U4629 (N_4629,N_926,N_2948);
nand U4630 (N_4630,N_2002,N_2958);
nor U4631 (N_4631,N_2560,N_1548);
nor U4632 (N_4632,N_563,N_1361);
nor U4633 (N_4633,N_2438,N_1364);
or U4634 (N_4634,N_1615,N_1255);
nor U4635 (N_4635,N_2662,N_379);
or U4636 (N_4636,N_2712,N_2849);
xor U4637 (N_4637,N_902,N_2292);
nor U4638 (N_4638,N_1236,N_1906);
and U4639 (N_4639,N_1056,N_2265);
and U4640 (N_4640,N_2911,N_88);
or U4641 (N_4641,N_551,N_188);
nor U4642 (N_4642,N_1712,N_2929);
or U4643 (N_4643,N_2252,N_2895);
nor U4644 (N_4644,N_292,N_2549);
and U4645 (N_4645,N_2022,N_1148);
nor U4646 (N_4646,N_2173,N_1705);
nor U4647 (N_4647,N_2372,N_2351);
and U4648 (N_4648,N_457,N_2874);
or U4649 (N_4649,N_2730,N_1836);
and U4650 (N_4650,N_1090,N_2073);
nand U4651 (N_4651,N_2076,N_2514);
nand U4652 (N_4652,N_29,N_2529);
or U4653 (N_4653,N_1022,N_2195);
and U4654 (N_4654,N_2254,N_1493);
xor U4655 (N_4655,N_1067,N_9);
nor U4656 (N_4656,N_919,N_2147);
nand U4657 (N_4657,N_2797,N_2670);
nor U4658 (N_4658,N_486,N_660);
and U4659 (N_4659,N_594,N_1222);
or U4660 (N_4660,N_434,N_2582);
or U4661 (N_4661,N_2515,N_701);
nand U4662 (N_4662,N_1322,N_1797);
or U4663 (N_4663,N_1387,N_2974);
and U4664 (N_4664,N_2597,N_1698);
nor U4665 (N_4665,N_2967,N_1989);
nor U4666 (N_4666,N_1479,N_478);
or U4667 (N_4667,N_1899,N_1438);
and U4668 (N_4668,N_1785,N_2747);
or U4669 (N_4669,N_1248,N_316);
or U4670 (N_4670,N_2516,N_799);
or U4671 (N_4671,N_2158,N_1715);
or U4672 (N_4672,N_2173,N_2392);
nand U4673 (N_4673,N_435,N_319);
nor U4674 (N_4674,N_79,N_1618);
or U4675 (N_4675,N_1718,N_1545);
or U4676 (N_4676,N_2848,N_2133);
or U4677 (N_4677,N_1532,N_1694);
nand U4678 (N_4678,N_1762,N_1600);
nor U4679 (N_4679,N_784,N_2410);
nor U4680 (N_4680,N_1093,N_1125);
nor U4681 (N_4681,N_318,N_1609);
or U4682 (N_4682,N_1294,N_1980);
nand U4683 (N_4683,N_1257,N_1643);
or U4684 (N_4684,N_2874,N_2430);
nand U4685 (N_4685,N_1410,N_2428);
or U4686 (N_4686,N_2998,N_245);
nand U4687 (N_4687,N_1770,N_338);
nor U4688 (N_4688,N_436,N_1557);
nand U4689 (N_4689,N_509,N_712);
xor U4690 (N_4690,N_2681,N_2878);
or U4691 (N_4691,N_1293,N_1699);
nand U4692 (N_4692,N_1874,N_607);
nand U4693 (N_4693,N_1678,N_1289);
and U4694 (N_4694,N_762,N_2550);
and U4695 (N_4695,N_993,N_2861);
or U4696 (N_4696,N_1594,N_2574);
nor U4697 (N_4697,N_844,N_2824);
nand U4698 (N_4698,N_1883,N_2601);
nand U4699 (N_4699,N_1869,N_2615);
nand U4700 (N_4700,N_1651,N_2665);
and U4701 (N_4701,N_1654,N_1090);
or U4702 (N_4702,N_1006,N_2665);
or U4703 (N_4703,N_2006,N_278);
and U4704 (N_4704,N_2294,N_211);
nand U4705 (N_4705,N_379,N_2542);
and U4706 (N_4706,N_1818,N_534);
nor U4707 (N_4707,N_2395,N_1718);
nand U4708 (N_4708,N_2443,N_1926);
nor U4709 (N_4709,N_572,N_473);
nor U4710 (N_4710,N_184,N_2784);
and U4711 (N_4711,N_1319,N_1559);
nand U4712 (N_4712,N_278,N_2429);
and U4713 (N_4713,N_476,N_1875);
and U4714 (N_4714,N_257,N_2518);
nand U4715 (N_4715,N_2549,N_2311);
and U4716 (N_4716,N_225,N_2756);
nor U4717 (N_4717,N_477,N_577);
or U4718 (N_4718,N_874,N_1342);
nand U4719 (N_4719,N_1372,N_888);
nor U4720 (N_4720,N_1172,N_2323);
and U4721 (N_4721,N_2058,N_1079);
nor U4722 (N_4722,N_801,N_1098);
and U4723 (N_4723,N_2391,N_2533);
or U4724 (N_4724,N_976,N_996);
or U4725 (N_4725,N_2560,N_2844);
and U4726 (N_4726,N_511,N_126);
xnor U4727 (N_4727,N_2990,N_1718);
and U4728 (N_4728,N_1174,N_2226);
and U4729 (N_4729,N_2448,N_1336);
nand U4730 (N_4730,N_1819,N_2297);
and U4731 (N_4731,N_2072,N_1442);
or U4732 (N_4732,N_1234,N_251);
or U4733 (N_4733,N_1034,N_1736);
and U4734 (N_4734,N_524,N_1450);
or U4735 (N_4735,N_56,N_1082);
and U4736 (N_4736,N_2630,N_1959);
nand U4737 (N_4737,N_399,N_2909);
and U4738 (N_4738,N_887,N_140);
and U4739 (N_4739,N_2101,N_2150);
nor U4740 (N_4740,N_529,N_656);
nor U4741 (N_4741,N_922,N_478);
nor U4742 (N_4742,N_1317,N_2307);
or U4743 (N_4743,N_2419,N_726);
and U4744 (N_4744,N_2999,N_590);
nand U4745 (N_4745,N_63,N_630);
nor U4746 (N_4746,N_2581,N_80);
nor U4747 (N_4747,N_2572,N_1757);
nand U4748 (N_4748,N_1624,N_629);
and U4749 (N_4749,N_160,N_540);
nor U4750 (N_4750,N_1557,N_2450);
or U4751 (N_4751,N_2131,N_824);
and U4752 (N_4752,N_2482,N_2943);
nor U4753 (N_4753,N_2662,N_1908);
nand U4754 (N_4754,N_485,N_1068);
nand U4755 (N_4755,N_1646,N_801);
nand U4756 (N_4756,N_1379,N_1666);
and U4757 (N_4757,N_2369,N_1610);
or U4758 (N_4758,N_639,N_2058);
nor U4759 (N_4759,N_200,N_2151);
nand U4760 (N_4760,N_869,N_2118);
nor U4761 (N_4761,N_1205,N_1473);
or U4762 (N_4762,N_2527,N_2939);
nor U4763 (N_4763,N_492,N_1108);
or U4764 (N_4764,N_403,N_1246);
and U4765 (N_4765,N_2806,N_2860);
nand U4766 (N_4766,N_951,N_2194);
nor U4767 (N_4767,N_1774,N_201);
or U4768 (N_4768,N_2940,N_1577);
nor U4769 (N_4769,N_1186,N_1187);
nand U4770 (N_4770,N_507,N_2792);
xor U4771 (N_4771,N_72,N_542);
nand U4772 (N_4772,N_2637,N_1208);
or U4773 (N_4773,N_1694,N_1368);
or U4774 (N_4774,N_1033,N_1106);
nor U4775 (N_4775,N_1702,N_2492);
nand U4776 (N_4776,N_131,N_1721);
or U4777 (N_4777,N_2692,N_1788);
nor U4778 (N_4778,N_1196,N_915);
or U4779 (N_4779,N_1659,N_2009);
nor U4780 (N_4780,N_1624,N_2186);
and U4781 (N_4781,N_2032,N_150);
or U4782 (N_4782,N_645,N_1681);
or U4783 (N_4783,N_541,N_1079);
and U4784 (N_4784,N_685,N_2766);
or U4785 (N_4785,N_1732,N_2487);
nand U4786 (N_4786,N_705,N_1500);
nor U4787 (N_4787,N_595,N_199);
nor U4788 (N_4788,N_1169,N_1229);
and U4789 (N_4789,N_497,N_1953);
and U4790 (N_4790,N_1903,N_2348);
and U4791 (N_4791,N_1127,N_1705);
nand U4792 (N_4792,N_1267,N_490);
nand U4793 (N_4793,N_1441,N_272);
or U4794 (N_4794,N_1062,N_1841);
nand U4795 (N_4795,N_2804,N_1136);
and U4796 (N_4796,N_977,N_1532);
or U4797 (N_4797,N_903,N_208);
nor U4798 (N_4798,N_2229,N_2827);
nand U4799 (N_4799,N_928,N_1488);
nand U4800 (N_4800,N_2350,N_2001);
and U4801 (N_4801,N_985,N_2425);
or U4802 (N_4802,N_224,N_2918);
or U4803 (N_4803,N_1850,N_1915);
nand U4804 (N_4804,N_2619,N_1732);
or U4805 (N_4805,N_1332,N_1926);
nor U4806 (N_4806,N_225,N_2879);
or U4807 (N_4807,N_250,N_2836);
nor U4808 (N_4808,N_1493,N_2834);
xor U4809 (N_4809,N_622,N_2274);
or U4810 (N_4810,N_2155,N_2206);
and U4811 (N_4811,N_2264,N_2209);
nor U4812 (N_4812,N_1167,N_351);
or U4813 (N_4813,N_1488,N_1249);
nor U4814 (N_4814,N_369,N_793);
or U4815 (N_4815,N_2796,N_1464);
nor U4816 (N_4816,N_871,N_2159);
nand U4817 (N_4817,N_1829,N_147);
nand U4818 (N_4818,N_105,N_1343);
nand U4819 (N_4819,N_1544,N_2509);
and U4820 (N_4820,N_2616,N_2502);
nand U4821 (N_4821,N_1389,N_2205);
nor U4822 (N_4822,N_261,N_212);
or U4823 (N_4823,N_434,N_1290);
and U4824 (N_4824,N_1223,N_2366);
or U4825 (N_4825,N_126,N_2485);
nand U4826 (N_4826,N_2906,N_1855);
nor U4827 (N_4827,N_1927,N_448);
or U4828 (N_4828,N_1128,N_2594);
nand U4829 (N_4829,N_255,N_1788);
or U4830 (N_4830,N_238,N_1224);
or U4831 (N_4831,N_619,N_36);
nand U4832 (N_4832,N_2777,N_2863);
nor U4833 (N_4833,N_668,N_2709);
nand U4834 (N_4834,N_2163,N_2191);
nand U4835 (N_4835,N_1820,N_2315);
nand U4836 (N_4836,N_1242,N_601);
nor U4837 (N_4837,N_397,N_1677);
nor U4838 (N_4838,N_1618,N_1678);
nor U4839 (N_4839,N_1220,N_1244);
or U4840 (N_4840,N_1000,N_2178);
nor U4841 (N_4841,N_1768,N_1156);
or U4842 (N_4842,N_2939,N_109);
or U4843 (N_4843,N_2083,N_1923);
nor U4844 (N_4844,N_2219,N_2131);
and U4845 (N_4845,N_2650,N_1815);
xor U4846 (N_4846,N_1957,N_1448);
and U4847 (N_4847,N_1563,N_478);
or U4848 (N_4848,N_2212,N_1029);
nand U4849 (N_4849,N_2354,N_1174);
nand U4850 (N_4850,N_2066,N_1463);
nand U4851 (N_4851,N_2548,N_2891);
nor U4852 (N_4852,N_122,N_1209);
and U4853 (N_4853,N_2788,N_329);
and U4854 (N_4854,N_1948,N_769);
nor U4855 (N_4855,N_2154,N_77);
or U4856 (N_4856,N_105,N_1786);
and U4857 (N_4857,N_17,N_1638);
nor U4858 (N_4858,N_318,N_1250);
nand U4859 (N_4859,N_2222,N_989);
nor U4860 (N_4860,N_1818,N_137);
or U4861 (N_4861,N_2507,N_2838);
xnor U4862 (N_4862,N_900,N_2242);
or U4863 (N_4863,N_352,N_2033);
nand U4864 (N_4864,N_2551,N_1035);
and U4865 (N_4865,N_1243,N_447);
nor U4866 (N_4866,N_2549,N_506);
and U4867 (N_4867,N_608,N_1960);
nand U4868 (N_4868,N_100,N_2175);
and U4869 (N_4869,N_336,N_220);
nand U4870 (N_4870,N_481,N_2802);
nor U4871 (N_4871,N_414,N_237);
nand U4872 (N_4872,N_304,N_823);
and U4873 (N_4873,N_964,N_1958);
or U4874 (N_4874,N_764,N_1610);
and U4875 (N_4875,N_1547,N_339);
nand U4876 (N_4876,N_1450,N_1342);
and U4877 (N_4877,N_993,N_699);
nand U4878 (N_4878,N_1790,N_2854);
and U4879 (N_4879,N_741,N_323);
nor U4880 (N_4880,N_2677,N_1875);
xor U4881 (N_4881,N_1972,N_109);
or U4882 (N_4882,N_1789,N_1603);
nor U4883 (N_4883,N_2204,N_2651);
and U4884 (N_4884,N_1170,N_1040);
nor U4885 (N_4885,N_2253,N_194);
nand U4886 (N_4886,N_2391,N_980);
nor U4887 (N_4887,N_52,N_1440);
nor U4888 (N_4888,N_1699,N_1652);
nor U4889 (N_4889,N_989,N_1855);
nor U4890 (N_4890,N_2568,N_1288);
or U4891 (N_4891,N_2088,N_1766);
nand U4892 (N_4892,N_1732,N_1571);
xor U4893 (N_4893,N_249,N_1915);
and U4894 (N_4894,N_2019,N_2595);
and U4895 (N_4895,N_1813,N_1064);
and U4896 (N_4896,N_676,N_237);
nand U4897 (N_4897,N_2876,N_161);
and U4898 (N_4898,N_962,N_2245);
and U4899 (N_4899,N_2964,N_416);
nor U4900 (N_4900,N_2146,N_414);
or U4901 (N_4901,N_16,N_1016);
or U4902 (N_4902,N_2570,N_2537);
and U4903 (N_4903,N_1565,N_2632);
or U4904 (N_4904,N_4,N_59);
or U4905 (N_4905,N_1100,N_2982);
and U4906 (N_4906,N_2682,N_2743);
and U4907 (N_4907,N_2516,N_2469);
and U4908 (N_4908,N_372,N_1353);
nor U4909 (N_4909,N_169,N_151);
or U4910 (N_4910,N_1423,N_2473);
and U4911 (N_4911,N_383,N_641);
or U4912 (N_4912,N_81,N_1977);
or U4913 (N_4913,N_2838,N_2307);
nand U4914 (N_4914,N_387,N_1738);
nor U4915 (N_4915,N_2488,N_2902);
xor U4916 (N_4916,N_2107,N_2067);
and U4917 (N_4917,N_2159,N_1856);
nand U4918 (N_4918,N_2306,N_331);
nand U4919 (N_4919,N_2085,N_1851);
and U4920 (N_4920,N_1077,N_759);
nor U4921 (N_4921,N_558,N_110);
or U4922 (N_4922,N_1182,N_995);
nand U4923 (N_4923,N_350,N_626);
nand U4924 (N_4924,N_1173,N_457);
or U4925 (N_4925,N_990,N_1275);
nor U4926 (N_4926,N_2620,N_931);
nand U4927 (N_4927,N_1365,N_744);
and U4928 (N_4928,N_2749,N_308);
and U4929 (N_4929,N_2351,N_1995);
nand U4930 (N_4930,N_2996,N_1265);
and U4931 (N_4931,N_698,N_200);
or U4932 (N_4932,N_2755,N_201);
or U4933 (N_4933,N_441,N_215);
or U4934 (N_4934,N_509,N_2502);
nand U4935 (N_4935,N_2284,N_2010);
nand U4936 (N_4936,N_310,N_2528);
xor U4937 (N_4937,N_813,N_2419);
nor U4938 (N_4938,N_408,N_1732);
nand U4939 (N_4939,N_264,N_1650);
and U4940 (N_4940,N_1962,N_2219);
nor U4941 (N_4941,N_2167,N_1512);
nand U4942 (N_4942,N_541,N_2035);
and U4943 (N_4943,N_1659,N_1958);
nand U4944 (N_4944,N_2715,N_2486);
nand U4945 (N_4945,N_776,N_426);
nand U4946 (N_4946,N_1811,N_2947);
or U4947 (N_4947,N_2344,N_2909);
nor U4948 (N_4948,N_2434,N_1066);
nor U4949 (N_4949,N_1511,N_2128);
nor U4950 (N_4950,N_1963,N_2337);
and U4951 (N_4951,N_1975,N_1254);
nor U4952 (N_4952,N_2262,N_2482);
or U4953 (N_4953,N_2708,N_1019);
and U4954 (N_4954,N_2945,N_2844);
nor U4955 (N_4955,N_2091,N_2812);
nor U4956 (N_4956,N_805,N_1041);
or U4957 (N_4957,N_660,N_348);
or U4958 (N_4958,N_173,N_1388);
and U4959 (N_4959,N_2303,N_2290);
nand U4960 (N_4960,N_1630,N_616);
nand U4961 (N_4961,N_834,N_971);
nand U4962 (N_4962,N_1237,N_272);
and U4963 (N_4963,N_1869,N_1756);
or U4964 (N_4964,N_2962,N_373);
and U4965 (N_4965,N_720,N_849);
nor U4966 (N_4966,N_2238,N_1543);
or U4967 (N_4967,N_1914,N_324);
or U4968 (N_4968,N_1487,N_938);
and U4969 (N_4969,N_2948,N_2700);
xnor U4970 (N_4970,N_2694,N_2090);
or U4971 (N_4971,N_1925,N_2911);
or U4972 (N_4972,N_2445,N_282);
or U4973 (N_4973,N_1278,N_2250);
nand U4974 (N_4974,N_419,N_1592);
or U4975 (N_4975,N_61,N_2584);
and U4976 (N_4976,N_231,N_2761);
and U4977 (N_4977,N_422,N_2291);
nor U4978 (N_4978,N_2019,N_2010);
nand U4979 (N_4979,N_1239,N_1828);
or U4980 (N_4980,N_1971,N_511);
nor U4981 (N_4981,N_1188,N_1714);
or U4982 (N_4982,N_223,N_2562);
nand U4983 (N_4983,N_516,N_311);
nor U4984 (N_4984,N_1503,N_2596);
nand U4985 (N_4985,N_2792,N_976);
and U4986 (N_4986,N_99,N_223);
and U4987 (N_4987,N_2763,N_2882);
nor U4988 (N_4988,N_2774,N_2494);
or U4989 (N_4989,N_2816,N_235);
or U4990 (N_4990,N_1847,N_1753);
and U4991 (N_4991,N_2943,N_234);
or U4992 (N_4992,N_2953,N_195);
and U4993 (N_4993,N_535,N_1399);
or U4994 (N_4994,N_2290,N_2813);
nor U4995 (N_4995,N_2656,N_1624);
and U4996 (N_4996,N_2494,N_1124);
nor U4997 (N_4997,N_1227,N_402);
nor U4998 (N_4998,N_1891,N_1958);
or U4999 (N_4999,N_1018,N_82);
nor U5000 (N_5000,N_1082,N_2406);
or U5001 (N_5001,N_2443,N_2827);
and U5002 (N_5002,N_2819,N_2269);
or U5003 (N_5003,N_2925,N_359);
and U5004 (N_5004,N_2995,N_206);
nor U5005 (N_5005,N_384,N_2261);
and U5006 (N_5006,N_2823,N_2140);
or U5007 (N_5007,N_2544,N_2409);
or U5008 (N_5008,N_2909,N_87);
nand U5009 (N_5009,N_1198,N_1203);
and U5010 (N_5010,N_691,N_2897);
nand U5011 (N_5011,N_2753,N_1290);
nor U5012 (N_5012,N_375,N_678);
nor U5013 (N_5013,N_2428,N_188);
or U5014 (N_5014,N_2959,N_2155);
nor U5015 (N_5015,N_2290,N_2201);
nand U5016 (N_5016,N_2153,N_1163);
nand U5017 (N_5017,N_2202,N_1619);
nor U5018 (N_5018,N_2091,N_70);
nor U5019 (N_5019,N_2966,N_2581);
and U5020 (N_5020,N_2961,N_500);
and U5021 (N_5021,N_2617,N_441);
nor U5022 (N_5022,N_2487,N_2063);
nor U5023 (N_5023,N_543,N_2675);
and U5024 (N_5024,N_468,N_433);
and U5025 (N_5025,N_2740,N_2327);
and U5026 (N_5026,N_2093,N_2225);
nand U5027 (N_5027,N_783,N_1208);
and U5028 (N_5028,N_537,N_768);
or U5029 (N_5029,N_75,N_568);
and U5030 (N_5030,N_325,N_680);
nor U5031 (N_5031,N_213,N_2942);
nor U5032 (N_5032,N_281,N_390);
nand U5033 (N_5033,N_2163,N_2868);
and U5034 (N_5034,N_1798,N_2096);
nand U5035 (N_5035,N_741,N_1613);
and U5036 (N_5036,N_895,N_569);
or U5037 (N_5037,N_1011,N_2533);
or U5038 (N_5038,N_2907,N_624);
and U5039 (N_5039,N_1301,N_1127);
nor U5040 (N_5040,N_2364,N_2370);
and U5041 (N_5041,N_1295,N_1738);
or U5042 (N_5042,N_2918,N_1266);
nand U5043 (N_5043,N_2479,N_377);
nand U5044 (N_5044,N_745,N_2981);
nand U5045 (N_5045,N_2337,N_79);
and U5046 (N_5046,N_1509,N_2760);
or U5047 (N_5047,N_2587,N_2299);
and U5048 (N_5048,N_646,N_2518);
nor U5049 (N_5049,N_1494,N_2797);
nand U5050 (N_5050,N_2355,N_1096);
nand U5051 (N_5051,N_879,N_1079);
nand U5052 (N_5052,N_1189,N_0);
and U5053 (N_5053,N_894,N_889);
nor U5054 (N_5054,N_1161,N_1801);
or U5055 (N_5055,N_421,N_1934);
nor U5056 (N_5056,N_277,N_2019);
or U5057 (N_5057,N_1001,N_2987);
nor U5058 (N_5058,N_2682,N_1484);
nand U5059 (N_5059,N_15,N_863);
and U5060 (N_5060,N_2263,N_915);
or U5061 (N_5061,N_1591,N_679);
nor U5062 (N_5062,N_1747,N_1448);
and U5063 (N_5063,N_1236,N_1400);
nor U5064 (N_5064,N_1171,N_721);
or U5065 (N_5065,N_1155,N_2986);
nand U5066 (N_5066,N_215,N_531);
and U5067 (N_5067,N_65,N_173);
or U5068 (N_5068,N_436,N_369);
and U5069 (N_5069,N_2844,N_258);
nor U5070 (N_5070,N_1312,N_296);
nand U5071 (N_5071,N_2419,N_537);
and U5072 (N_5072,N_413,N_1988);
nor U5073 (N_5073,N_1846,N_829);
or U5074 (N_5074,N_2123,N_2255);
or U5075 (N_5075,N_2913,N_555);
nor U5076 (N_5076,N_982,N_2914);
nor U5077 (N_5077,N_1600,N_1481);
and U5078 (N_5078,N_2365,N_1179);
nand U5079 (N_5079,N_2458,N_721);
or U5080 (N_5080,N_2787,N_2162);
and U5081 (N_5081,N_2024,N_2895);
and U5082 (N_5082,N_923,N_1715);
nor U5083 (N_5083,N_1481,N_2994);
nand U5084 (N_5084,N_1340,N_1515);
nor U5085 (N_5085,N_2761,N_266);
nor U5086 (N_5086,N_2639,N_575);
and U5087 (N_5087,N_692,N_1496);
or U5088 (N_5088,N_64,N_2379);
nor U5089 (N_5089,N_1856,N_2921);
and U5090 (N_5090,N_2055,N_1508);
nor U5091 (N_5091,N_1249,N_2612);
and U5092 (N_5092,N_973,N_1466);
nand U5093 (N_5093,N_2739,N_1493);
or U5094 (N_5094,N_2105,N_401);
nand U5095 (N_5095,N_2139,N_2468);
nand U5096 (N_5096,N_2741,N_2844);
nor U5097 (N_5097,N_1272,N_2407);
nor U5098 (N_5098,N_2365,N_1201);
nand U5099 (N_5099,N_1032,N_2523);
xnor U5100 (N_5100,N_2888,N_854);
and U5101 (N_5101,N_2279,N_1404);
and U5102 (N_5102,N_2324,N_991);
nor U5103 (N_5103,N_2208,N_2800);
or U5104 (N_5104,N_2820,N_2503);
or U5105 (N_5105,N_472,N_149);
nand U5106 (N_5106,N_2063,N_131);
and U5107 (N_5107,N_964,N_2291);
or U5108 (N_5108,N_1716,N_2978);
nand U5109 (N_5109,N_211,N_578);
nand U5110 (N_5110,N_11,N_2391);
nor U5111 (N_5111,N_989,N_2735);
or U5112 (N_5112,N_1285,N_2852);
or U5113 (N_5113,N_1747,N_1051);
or U5114 (N_5114,N_1595,N_297);
and U5115 (N_5115,N_2841,N_787);
or U5116 (N_5116,N_1344,N_367);
nor U5117 (N_5117,N_384,N_2764);
and U5118 (N_5118,N_70,N_1779);
or U5119 (N_5119,N_1447,N_896);
or U5120 (N_5120,N_1883,N_584);
nand U5121 (N_5121,N_212,N_393);
nand U5122 (N_5122,N_914,N_660);
nor U5123 (N_5123,N_2786,N_578);
nand U5124 (N_5124,N_336,N_2189);
nor U5125 (N_5125,N_2878,N_486);
nor U5126 (N_5126,N_2587,N_1774);
nor U5127 (N_5127,N_941,N_1870);
nand U5128 (N_5128,N_2674,N_2021);
and U5129 (N_5129,N_1458,N_1021);
or U5130 (N_5130,N_2074,N_2339);
or U5131 (N_5131,N_2913,N_1846);
nor U5132 (N_5132,N_2336,N_2959);
or U5133 (N_5133,N_2062,N_1830);
and U5134 (N_5134,N_1122,N_1681);
nand U5135 (N_5135,N_434,N_1496);
and U5136 (N_5136,N_238,N_414);
or U5137 (N_5137,N_860,N_209);
nor U5138 (N_5138,N_322,N_1301);
or U5139 (N_5139,N_421,N_2588);
xor U5140 (N_5140,N_980,N_433);
nand U5141 (N_5141,N_1994,N_2758);
or U5142 (N_5142,N_2205,N_64);
nand U5143 (N_5143,N_2782,N_190);
nand U5144 (N_5144,N_2564,N_1979);
nand U5145 (N_5145,N_1792,N_2596);
and U5146 (N_5146,N_2397,N_2307);
and U5147 (N_5147,N_1571,N_1115);
or U5148 (N_5148,N_1685,N_57);
nand U5149 (N_5149,N_477,N_1550);
nand U5150 (N_5150,N_637,N_1374);
nor U5151 (N_5151,N_1148,N_669);
nor U5152 (N_5152,N_2599,N_1922);
or U5153 (N_5153,N_1770,N_1961);
nor U5154 (N_5154,N_716,N_2648);
nor U5155 (N_5155,N_332,N_26);
or U5156 (N_5156,N_2872,N_2933);
nand U5157 (N_5157,N_1259,N_1090);
nand U5158 (N_5158,N_1491,N_765);
or U5159 (N_5159,N_1251,N_1965);
and U5160 (N_5160,N_1095,N_2755);
nand U5161 (N_5161,N_2314,N_2423);
xnor U5162 (N_5162,N_1845,N_1415);
nand U5163 (N_5163,N_881,N_1277);
and U5164 (N_5164,N_214,N_350);
and U5165 (N_5165,N_1101,N_158);
and U5166 (N_5166,N_627,N_143);
nor U5167 (N_5167,N_2878,N_2217);
or U5168 (N_5168,N_2331,N_2599);
nand U5169 (N_5169,N_1278,N_2653);
nand U5170 (N_5170,N_459,N_62);
and U5171 (N_5171,N_1561,N_218);
or U5172 (N_5172,N_282,N_1265);
and U5173 (N_5173,N_1876,N_614);
nor U5174 (N_5174,N_1522,N_1595);
or U5175 (N_5175,N_482,N_2332);
nor U5176 (N_5176,N_1340,N_41);
nor U5177 (N_5177,N_2023,N_505);
or U5178 (N_5178,N_2104,N_1797);
and U5179 (N_5179,N_2444,N_2515);
or U5180 (N_5180,N_2273,N_625);
or U5181 (N_5181,N_754,N_1809);
and U5182 (N_5182,N_2681,N_1779);
and U5183 (N_5183,N_1766,N_2098);
and U5184 (N_5184,N_2166,N_1361);
nor U5185 (N_5185,N_2327,N_521);
nand U5186 (N_5186,N_1281,N_2544);
nor U5187 (N_5187,N_776,N_543);
nor U5188 (N_5188,N_2883,N_509);
nand U5189 (N_5189,N_642,N_2515);
and U5190 (N_5190,N_1815,N_1834);
nand U5191 (N_5191,N_1930,N_900);
or U5192 (N_5192,N_828,N_2529);
or U5193 (N_5193,N_2059,N_1907);
nor U5194 (N_5194,N_1350,N_1354);
or U5195 (N_5195,N_784,N_1552);
nand U5196 (N_5196,N_539,N_1054);
and U5197 (N_5197,N_1070,N_2802);
nor U5198 (N_5198,N_582,N_1344);
or U5199 (N_5199,N_2201,N_529);
nor U5200 (N_5200,N_1662,N_976);
nand U5201 (N_5201,N_1333,N_2399);
nor U5202 (N_5202,N_290,N_1405);
nor U5203 (N_5203,N_1562,N_2599);
nand U5204 (N_5204,N_104,N_1124);
and U5205 (N_5205,N_2186,N_683);
and U5206 (N_5206,N_1505,N_978);
and U5207 (N_5207,N_1830,N_770);
nor U5208 (N_5208,N_1478,N_111);
nand U5209 (N_5209,N_2079,N_2251);
or U5210 (N_5210,N_1329,N_2310);
xnor U5211 (N_5211,N_2381,N_423);
and U5212 (N_5212,N_481,N_1579);
nand U5213 (N_5213,N_879,N_347);
or U5214 (N_5214,N_2193,N_1525);
and U5215 (N_5215,N_2761,N_2274);
nor U5216 (N_5216,N_800,N_529);
or U5217 (N_5217,N_942,N_2134);
and U5218 (N_5218,N_141,N_2605);
or U5219 (N_5219,N_999,N_781);
or U5220 (N_5220,N_2160,N_1623);
and U5221 (N_5221,N_889,N_977);
nand U5222 (N_5222,N_1994,N_1484);
nor U5223 (N_5223,N_1041,N_2242);
and U5224 (N_5224,N_2092,N_643);
or U5225 (N_5225,N_856,N_330);
or U5226 (N_5226,N_1518,N_1766);
and U5227 (N_5227,N_1825,N_752);
nand U5228 (N_5228,N_813,N_1049);
nand U5229 (N_5229,N_1636,N_25);
and U5230 (N_5230,N_243,N_1369);
or U5231 (N_5231,N_24,N_1615);
or U5232 (N_5232,N_1995,N_2007);
or U5233 (N_5233,N_1021,N_2020);
nand U5234 (N_5234,N_2370,N_421);
and U5235 (N_5235,N_2515,N_2504);
xor U5236 (N_5236,N_2897,N_2102);
nand U5237 (N_5237,N_1152,N_2834);
and U5238 (N_5238,N_1508,N_1);
nor U5239 (N_5239,N_1448,N_2320);
and U5240 (N_5240,N_2314,N_1531);
or U5241 (N_5241,N_392,N_114);
nor U5242 (N_5242,N_2603,N_2651);
nor U5243 (N_5243,N_1159,N_1852);
nor U5244 (N_5244,N_22,N_2865);
nor U5245 (N_5245,N_297,N_266);
nand U5246 (N_5246,N_2649,N_1643);
or U5247 (N_5247,N_2223,N_96);
and U5248 (N_5248,N_717,N_1173);
and U5249 (N_5249,N_2595,N_315);
and U5250 (N_5250,N_758,N_2414);
and U5251 (N_5251,N_318,N_316);
and U5252 (N_5252,N_640,N_2599);
or U5253 (N_5253,N_2208,N_1182);
nor U5254 (N_5254,N_2471,N_1309);
nand U5255 (N_5255,N_2110,N_1737);
nor U5256 (N_5256,N_973,N_2738);
nor U5257 (N_5257,N_524,N_187);
and U5258 (N_5258,N_2781,N_791);
nor U5259 (N_5259,N_2715,N_101);
or U5260 (N_5260,N_923,N_449);
and U5261 (N_5261,N_834,N_353);
or U5262 (N_5262,N_1793,N_619);
and U5263 (N_5263,N_2572,N_749);
nand U5264 (N_5264,N_262,N_1072);
or U5265 (N_5265,N_198,N_1954);
nand U5266 (N_5266,N_2152,N_2074);
nand U5267 (N_5267,N_1009,N_166);
nand U5268 (N_5268,N_2712,N_2657);
and U5269 (N_5269,N_1523,N_165);
or U5270 (N_5270,N_796,N_1869);
nor U5271 (N_5271,N_872,N_1544);
nor U5272 (N_5272,N_1633,N_1362);
nand U5273 (N_5273,N_933,N_1496);
or U5274 (N_5274,N_1034,N_619);
nand U5275 (N_5275,N_2587,N_1501);
nor U5276 (N_5276,N_1323,N_2594);
nand U5277 (N_5277,N_715,N_2580);
nor U5278 (N_5278,N_1067,N_1578);
nor U5279 (N_5279,N_2515,N_1458);
or U5280 (N_5280,N_2149,N_2926);
nand U5281 (N_5281,N_64,N_397);
nor U5282 (N_5282,N_2361,N_607);
nor U5283 (N_5283,N_1493,N_1307);
nand U5284 (N_5284,N_621,N_2351);
nand U5285 (N_5285,N_1273,N_632);
and U5286 (N_5286,N_2159,N_612);
or U5287 (N_5287,N_2540,N_1049);
or U5288 (N_5288,N_1546,N_641);
nand U5289 (N_5289,N_628,N_2305);
or U5290 (N_5290,N_1127,N_2016);
or U5291 (N_5291,N_2917,N_262);
or U5292 (N_5292,N_1642,N_393);
or U5293 (N_5293,N_590,N_1226);
and U5294 (N_5294,N_1248,N_676);
nor U5295 (N_5295,N_1524,N_1612);
nand U5296 (N_5296,N_2398,N_1578);
nand U5297 (N_5297,N_2518,N_2341);
or U5298 (N_5298,N_1392,N_710);
and U5299 (N_5299,N_1846,N_1138);
nor U5300 (N_5300,N_2086,N_1699);
or U5301 (N_5301,N_1321,N_218);
or U5302 (N_5302,N_2477,N_50);
and U5303 (N_5303,N_791,N_1245);
or U5304 (N_5304,N_1442,N_2985);
nand U5305 (N_5305,N_1688,N_2217);
nand U5306 (N_5306,N_2421,N_2713);
or U5307 (N_5307,N_2916,N_1452);
and U5308 (N_5308,N_1092,N_2903);
and U5309 (N_5309,N_1735,N_1452);
or U5310 (N_5310,N_2520,N_2987);
or U5311 (N_5311,N_3,N_165);
or U5312 (N_5312,N_1123,N_1286);
or U5313 (N_5313,N_2607,N_2850);
and U5314 (N_5314,N_373,N_319);
or U5315 (N_5315,N_541,N_70);
nand U5316 (N_5316,N_292,N_2298);
and U5317 (N_5317,N_950,N_2194);
nor U5318 (N_5318,N_2154,N_2612);
nand U5319 (N_5319,N_1151,N_1461);
nand U5320 (N_5320,N_1505,N_1552);
nand U5321 (N_5321,N_2072,N_2368);
and U5322 (N_5322,N_1111,N_344);
and U5323 (N_5323,N_2214,N_30);
or U5324 (N_5324,N_1752,N_1439);
nand U5325 (N_5325,N_152,N_2378);
nor U5326 (N_5326,N_2695,N_733);
and U5327 (N_5327,N_1451,N_2306);
and U5328 (N_5328,N_410,N_1426);
nand U5329 (N_5329,N_1053,N_548);
or U5330 (N_5330,N_1656,N_303);
nand U5331 (N_5331,N_277,N_2226);
nor U5332 (N_5332,N_1519,N_1828);
or U5333 (N_5333,N_1216,N_2675);
or U5334 (N_5334,N_498,N_2115);
nand U5335 (N_5335,N_649,N_2686);
or U5336 (N_5336,N_2461,N_1272);
nand U5337 (N_5337,N_1814,N_889);
or U5338 (N_5338,N_2034,N_1782);
nand U5339 (N_5339,N_629,N_1756);
and U5340 (N_5340,N_607,N_42);
or U5341 (N_5341,N_694,N_1552);
nor U5342 (N_5342,N_993,N_2244);
and U5343 (N_5343,N_1787,N_743);
and U5344 (N_5344,N_1452,N_1539);
and U5345 (N_5345,N_2790,N_2121);
nand U5346 (N_5346,N_933,N_892);
and U5347 (N_5347,N_175,N_955);
or U5348 (N_5348,N_1944,N_833);
nor U5349 (N_5349,N_1630,N_2153);
nor U5350 (N_5350,N_1414,N_769);
or U5351 (N_5351,N_813,N_2965);
nand U5352 (N_5352,N_2741,N_1422);
nor U5353 (N_5353,N_2279,N_2395);
and U5354 (N_5354,N_611,N_729);
and U5355 (N_5355,N_106,N_1554);
nand U5356 (N_5356,N_1234,N_287);
nor U5357 (N_5357,N_2114,N_2108);
nand U5358 (N_5358,N_2282,N_1595);
and U5359 (N_5359,N_1715,N_2090);
nor U5360 (N_5360,N_459,N_421);
nor U5361 (N_5361,N_2553,N_153);
and U5362 (N_5362,N_938,N_1862);
nand U5363 (N_5363,N_2550,N_330);
nand U5364 (N_5364,N_209,N_2156);
and U5365 (N_5365,N_945,N_387);
and U5366 (N_5366,N_2476,N_81);
or U5367 (N_5367,N_2779,N_1430);
and U5368 (N_5368,N_1118,N_2120);
nand U5369 (N_5369,N_449,N_1288);
nand U5370 (N_5370,N_1647,N_2232);
nor U5371 (N_5371,N_2295,N_2102);
and U5372 (N_5372,N_921,N_904);
nor U5373 (N_5373,N_2888,N_928);
nand U5374 (N_5374,N_1863,N_2001);
nand U5375 (N_5375,N_1647,N_2651);
nor U5376 (N_5376,N_1205,N_1374);
nor U5377 (N_5377,N_389,N_1513);
xor U5378 (N_5378,N_1808,N_212);
nand U5379 (N_5379,N_597,N_1939);
nor U5380 (N_5380,N_1240,N_700);
nand U5381 (N_5381,N_131,N_363);
nand U5382 (N_5382,N_1792,N_2931);
nand U5383 (N_5383,N_748,N_1693);
nand U5384 (N_5384,N_771,N_1708);
or U5385 (N_5385,N_1117,N_2192);
or U5386 (N_5386,N_108,N_1843);
nand U5387 (N_5387,N_2683,N_119);
or U5388 (N_5388,N_92,N_1258);
nand U5389 (N_5389,N_1861,N_659);
and U5390 (N_5390,N_2053,N_1217);
or U5391 (N_5391,N_2100,N_2775);
nand U5392 (N_5392,N_127,N_508);
nor U5393 (N_5393,N_2589,N_22);
nand U5394 (N_5394,N_1894,N_1281);
and U5395 (N_5395,N_1405,N_365);
nor U5396 (N_5396,N_1217,N_2489);
nor U5397 (N_5397,N_1950,N_1565);
nand U5398 (N_5398,N_213,N_2227);
nor U5399 (N_5399,N_996,N_2623);
and U5400 (N_5400,N_1578,N_1961);
or U5401 (N_5401,N_2625,N_1099);
or U5402 (N_5402,N_1699,N_2158);
nor U5403 (N_5403,N_566,N_2172);
and U5404 (N_5404,N_1886,N_2789);
or U5405 (N_5405,N_1292,N_2374);
or U5406 (N_5406,N_2890,N_1346);
nand U5407 (N_5407,N_184,N_2248);
and U5408 (N_5408,N_1974,N_1513);
nand U5409 (N_5409,N_891,N_1016);
and U5410 (N_5410,N_664,N_1414);
nand U5411 (N_5411,N_2016,N_1436);
or U5412 (N_5412,N_2827,N_1257);
or U5413 (N_5413,N_2788,N_223);
or U5414 (N_5414,N_1975,N_1746);
nor U5415 (N_5415,N_975,N_828);
or U5416 (N_5416,N_1173,N_164);
or U5417 (N_5417,N_2306,N_1783);
or U5418 (N_5418,N_2103,N_2969);
nand U5419 (N_5419,N_2757,N_1257);
nor U5420 (N_5420,N_2007,N_1508);
nor U5421 (N_5421,N_1582,N_1815);
or U5422 (N_5422,N_523,N_2465);
or U5423 (N_5423,N_2861,N_617);
nand U5424 (N_5424,N_458,N_2922);
or U5425 (N_5425,N_2590,N_922);
nand U5426 (N_5426,N_1432,N_280);
nor U5427 (N_5427,N_523,N_628);
or U5428 (N_5428,N_123,N_2692);
nor U5429 (N_5429,N_1317,N_2104);
and U5430 (N_5430,N_82,N_1217);
nor U5431 (N_5431,N_2432,N_86);
nand U5432 (N_5432,N_2918,N_2310);
and U5433 (N_5433,N_1245,N_2784);
nand U5434 (N_5434,N_769,N_2568);
nand U5435 (N_5435,N_2635,N_1209);
nor U5436 (N_5436,N_2290,N_2373);
or U5437 (N_5437,N_2970,N_1249);
and U5438 (N_5438,N_1814,N_2653);
or U5439 (N_5439,N_1178,N_237);
nor U5440 (N_5440,N_1140,N_659);
or U5441 (N_5441,N_1561,N_2242);
or U5442 (N_5442,N_2860,N_343);
and U5443 (N_5443,N_2190,N_1679);
nor U5444 (N_5444,N_314,N_1447);
nor U5445 (N_5445,N_632,N_2093);
and U5446 (N_5446,N_256,N_1385);
nand U5447 (N_5447,N_1684,N_2963);
and U5448 (N_5448,N_2556,N_2406);
nor U5449 (N_5449,N_161,N_306);
nand U5450 (N_5450,N_603,N_875);
nor U5451 (N_5451,N_54,N_1380);
nor U5452 (N_5452,N_1559,N_1644);
and U5453 (N_5453,N_322,N_2913);
or U5454 (N_5454,N_14,N_1592);
or U5455 (N_5455,N_2504,N_1979);
and U5456 (N_5456,N_2530,N_628);
or U5457 (N_5457,N_2601,N_929);
nand U5458 (N_5458,N_2807,N_2364);
nand U5459 (N_5459,N_1589,N_1959);
and U5460 (N_5460,N_1641,N_376);
and U5461 (N_5461,N_1613,N_1303);
nor U5462 (N_5462,N_1896,N_1811);
or U5463 (N_5463,N_1155,N_1960);
nor U5464 (N_5464,N_2122,N_1857);
or U5465 (N_5465,N_566,N_1245);
or U5466 (N_5466,N_1966,N_2245);
nor U5467 (N_5467,N_1939,N_1576);
nand U5468 (N_5468,N_2235,N_1549);
or U5469 (N_5469,N_307,N_2075);
nor U5470 (N_5470,N_809,N_2409);
nand U5471 (N_5471,N_1796,N_2978);
and U5472 (N_5472,N_519,N_28);
or U5473 (N_5473,N_805,N_966);
and U5474 (N_5474,N_447,N_1383);
or U5475 (N_5475,N_1739,N_1117);
nor U5476 (N_5476,N_182,N_177);
and U5477 (N_5477,N_994,N_1011);
or U5478 (N_5478,N_1040,N_2847);
nor U5479 (N_5479,N_992,N_1260);
or U5480 (N_5480,N_1805,N_1051);
and U5481 (N_5481,N_1006,N_2211);
and U5482 (N_5482,N_972,N_2825);
nand U5483 (N_5483,N_2986,N_1984);
nand U5484 (N_5484,N_1554,N_9);
nand U5485 (N_5485,N_1892,N_1765);
or U5486 (N_5486,N_1923,N_2501);
nand U5487 (N_5487,N_1285,N_981);
xnor U5488 (N_5488,N_2202,N_863);
nor U5489 (N_5489,N_978,N_2563);
nor U5490 (N_5490,N_2745,N_765);
nand U5491 (N_5491,N_1728,N_2907);
nand U5492 (N_5492,N_1118,N_2894);
and U5493 (N_5493,N_958,N_2343);
nor U5494 (N_5494,N_1208,N_283);
nand U5495 (N_5495,N_1596,N_1121);
and U5496 (N_5496,N_1496,N_195);
nor U5497 (N_5497,N_1159,N_1377);
or U5498 (N_5498,N_224,N_446);
and U5499 (N_5499,N_1738,N_813);
nor U5500 (N_5500,N_659,N_2536);
nand U5501 (N_5501,N_1878,N_2400);
and U5502 (N_5502,N_2102,N_2202);
and U5503 (N_5503,N_901,N_510);
and U5504 (N_5504,N_2574,N_2963);
nand U5505 (N_5505,N_1284,N_1336);
nor U5506 (N_5506,N_1805,N_1284);
nor U5507 (N_5507,N_468,N_1851);
nor U5508 (N_5508,N_2813,N_523);
and U5509 (N_5509,N_1823,N_2372);
nor U5510 (N_5510,N_1925,N_124);
and U5511 (N_5511,N_2634,N_1432);
nor U5512 (N_5512,N_1670,N_2666);
nand U5513 (N_5513,N_1675,N_2359);
nor U5514 (N_5514,N_721,N_2304);
and U5515 (N_5515,N_2861,N_374);
and U5516 (N_5516,N_2083,N_1587);
or U5517 (N_5517,N_459,N_1218);
nand U5518 (N_5518,N_1495,N_2995);
nand U5519 (N_5519,N_488,N_2485);
nand U5520 (N_5520,N_733,N_461);
nand U5521 (N_5521,N_1730,N_1949);
and U5522 (N_5522,N_2875,N_934);
nand U5523 (N_5523,N_224,N_1362);
nand U5524 (N_5524,N_1211,N_2918);
nand U5525 (N_5525,N_973,N_314);
and U5526 (N_5526,N_1461,N_2021);
and U5527 (N_5527,N_592,N_2554);
nand U5528 (N_5528,N_1798,N_494);
nor U5529 (N_5529,N_807,N_627);
nor U5530 (N_5530,N_1105,N_1888);
and U5531 (N_5531,N_1985,N_1579);
nor U5532 (N_5532,N_1341,N_742);
nand U5533 (N_5533,N_2343,N_1252);
and U5534 (N_5534,N_2798,N_1081);
nor U5535 (N_5535,N_1104,N_2717);
and U5536 (N_5536,N_2537,N_1362);
and U5537 (N_5537,N_2061,N_1772);
or U5538 (N_5538,N_848,N_2092);
nand U5539 (N_5539,N_926,N_56);
nor U5540 (N_5540,N_51,N_503);
or U5541 (N_5541,N_2267,N_548);
nand U5542 (N_5542,N_2423,N_2345);
and U5543 (N_5543,N_135,N_2156);
and U5544 (N_5544,N_2510,N_1384);
and U5545 (N_5545,N_50,N_2608);
and U5546 (N_5546,N_1124,N_1022);
nor U5547 (N_5547,N_980,N_595);
or U5548 (N_5548,N_2734,N_2796);
or U5549 (N_5549,N_2536,N_1527);
or U5550 (N_5550,N_2484,N_2360);
or U5551 (N_5551,N_541,N_2398);
xor U5552 (N_5552,N_1248,N_866);
or U5553 (N_5553,N_1011,N_1754);
or U5554 (N_5554,N_1393,N_2298);
and U5555 (N_5555,N_2843,N_2641);
nand U5556 (N_5556,N_234,N_1464);
nand U5557 (N_5557,N_803,N_2364);
and U5558 (N_5558,N_2605,N_2663);
nor U5559 (N_5559,N_1535,N_2879);
and U5560 (N_5560,N_1849,N_1717);
or U5561 (N_5561,N_998,N_2076);
nor U5562 (N_5562,N_613,N_1830);
or U5563 (N_5563,N_2303,N_489);
and U5564 (N_5564,N_2940,N_1685);
and U5565 (N_5565,N_1771,N_594);
or U5566 (N_5566,N_20,N_1460);
and U5567 (N_5567,N_2746,N_2760);
or U5568 (N_5568,N_1638,N_568);
and U5569 (N_5569,N_557,N_1218);
nor U5570 (N_5570,N_815,N_697);
or U5571 (N_5571,N_1454,N_190);
or U5572 (N_5572,N_2697,N_1485);
nor U5573 (N_5573,N_769,N_938);
xor U5574 (N_5574,N_1593,N_945);
nor U5575 (N_5575,N_550,N_690);
and U5576 (N_5576,N_2056,N_2315);
or U5577 (N_5577,N_787,N_1420);
or U5578 (N_5578,N_1598,N_1371);
and U5579 (N_5579,N_1789,N_1409);
and U5580 (N_5580,N_2852,N_1924);
or U5581 (N_5581,N_1119,N_1760);
and U5582 (N_5582,N_1725,N_767);
nor U5583 (N_5583,N_694,N_1840);
or U5584 (N_5584,N_776,N_1018);
nand U5585 (N_5585,N_2159,N_1727);
and U5586 (N_5586,N_1831,N_314);
or U5587 (N_5587,N_119,N_2999);
nand U5588 (N_5588,N_2597,N_2596);
nor U5589 (N_5589,N_569,N_1898);
or U5590 (N_5590,N_2071,N_2221);
nor U5591 (N_5591,N_1456,N_2566);
nand U5592 (N_5592,N_1268,N_2254);
nor U5593 (N_5593,N_2456,N_2626);
nand U5594 (N_5594,N_1199,N_1379);
or U5595 (N_5595,N_391,N_2823);
nor U5596 (N_5596,N_1468,N_1285);
and U5597 (N_5597,N_2078,N_1808);
and U5598 (N_5598,N_325,N_174);
nor U5599 (N_5599,N_401,N_930);
nor U5600 (N_5600,N_2652,N_2231);
nor U5601 (N_5601,N_1753,N_320);
nor U5602 (N_5602,N_1746,N_2187);
nand U5603 (N_5603,N_287,N_2125);
nor U5604 (N_5604,N_1161,N_2290);
nor U5605 (N_5605,N_671,N_2710);
and U5606 (N_5606,N_2370,N_1459);
or U5607 (N_5607,N_688,N_2588);
nand U5608 (N_5608,N_1147,N_1253);
and U5609 (N_5609,N_2271,N_2403);
and U5610 (N_5610,N_1317,N_2625);
nand U5611 (N_5611,N_2167,N_1311);
or U5612 (N_5612,N_1598,N_922);
and U5613 (N_5613,N_78,N_2231);
or U5614 (N_5614,N_1528,N_2079);
and U5615 (N_5615,N_1593,N_793);
nor U5616 (N_5616,N_1423,N_1210);
nor U5617 (N_5617,N_735,N_2974);
nor U5618 (N_5618,N_549,N_69);
nor U5619 (N_5619,N_746,N_794);
xor U5620 (N_5620,N_1844,N_2563);
nand U5621 (N_5621,N_2226,N_1210);
nand U5622 (N_5622,N_1130,N_881);
or U5623 (N_5623,N_118,N_430);
and U5624 (N_5624,N_364,N_0);
nand U5625 (N_5625,N_1408,N_2144);
or U5626 (N_5626,N_2429,N_886);
and U5627 (N_5627,N_691,N_1739);
or U5628 (N_5628,N_611,N_637);
and U5629 (N_5629,N_1462,N_2427);
nand U5630 (N_5630,N_816,N_2053);
or U5631 (N_5631,N_1987,N_2823);
or U5632 (N_5632,N_2236,N_590);
and U5633 (N_5633,N_674,N_2335);
and U5634 (N_5634,N_2531,N_1302);
nand U5635 (N_5635,N_1638,N_1192);
and U5636 (N_5636,N_1249,N_2541);
nor U5637 (N_5637,N_2091,N_1832);
or U5638 (N_5638,N_158,N_2011);
nor U5639 (N_5639,N_888,N_2550);
and U5640 (N_5640,N_2442,N_1726);
and U5641 (N_5641,N_2755,N_1713);
or U5642 (N_5642,N_2969,N_2273);
and U5643 (N_5643,N_2300,N_2162);
nor U5644 (N_5644,N_1710,N_1410);
nand U5645 (N_5645,N_2441,N_1164);
or U5646 (N_5646,N_250,N_1615);
and U5647 (N_5647,N_2943,N_1110);
nand U5648 (N_5648,N_830,N_1469);
or U5649 (N_5649,N_2270,N_2027);
nand U5650 (N_5650,N_805,N_2939);
or U5651 (N_5651,N_651,N_1015);
nand U5652 (N_5652,N_2405,N_2142);
nor U5653 (N_5653,N_455,N_1904);
and U5654 (N_5654,N_1005,N_2322);
or U5655 (N_5655,N_1143,N_463);
and U5656 (N_5656,N_2574,N_668);
or U5657 (N_5657,N_570,N_2765);
and U5658 (N_5658,N_1687,N_1594);
or U5659 (N_5659,N_2512,N_2063);
nor U5660 (N_5660,N_616,N_1136);
nor U5661 (N_5661,N_1474,N_2443);
nor U5662 (N_5662,N_2264,N_517);
xnor U5663 (N_5663,N_1490,N_2016);
or U5664 (N_5664,N_2961,N_549);
nand U5665 (N_5665,N_1964,N_2738);
nor U5666 (N_5666,N_1356,N_1264);
and U5667 (N_5667,N_1758,N_1889);
and U5668 (N_5668,N_202,N_2231);
nand U5669 (N_5669,N_2154,N_2861);
xor U5670 (N_5670,N_766,N_2314);
or U5671 (N_5671,N_2285,N_278);
nand U5672 (N_5672,N_183,N_800);
nand U5673 (N_5673,N_520,N_2682);
or U5674 (N_5674,N_1912,N_2355);
nor U5675 (N_5675,N_1182,N_927);
nand U5676 (N_5676,N_1462,N_2272);
or U5677 (N_5677,N_2502,N_1893);
nor U5678 (N_5678,N_1819,N_775);
or U5679 (N_5679,N_1016,N_347);
xnor U5680 (N_5680,N_2645,N_2912);
and U5681 (N_5681,N_2239,N_338);
nor U5682 (N_5682,N_2782,N_699);
nand U5683 (N_5683,N_2329,N_2514);
and U5684 (N_5684,N_806,N_1151);
nand U5685 (N_5685,N_1727,N_1486);
nand U5686 (N_5686,N_1015,N_2546);
and U5687 (N_5687,N_1474,N_1876);
and U5688 (N_5688,N_2623,N_840);
nor U5689 (N_5689,N_1069,N_1625);
or U5690 (N_5690,N_1177,N_925);
nor U5691 (N_5691,N_2852,N_1731);
nor U5692 (N_5692,N_1017,N_2583);
and U5693 (N_5693,N_365,N_790);
nor U5694 (N_5694,N_1604,N_2967);
or U5695 (N_5695,N_1594,N_2379);
nor U5696 (N_5696,N_1976,N_928);
nor U5697 (N_5697,N_455,N_1660);
and U5698 (N_5698,N_474,N_1986);
nor U5699 (N_5699,N_1266,N_1601);
and U5700 (N_5700,N_53,N_2809);
nor U5701 (N_5701,N_1134,N_2724);
nor U5702 (N_5702,N_2107,N_1326);
nor U5703 (N_5703,N_2289,N_610);
or U5704 (N_5704,N_2888,N_1897);
nand U5705 (N_5705,N_2101,N_2609);
or U5706 (N_5706,N_1400,N_1450);
nor U5707 (N_5707,N_63,N_1402);
or U5708 (N_5708,N_50,N_2166);
or U5709 (N_5709,N_2044,N_769);
and U5710 (N_5710,N_1705,N_2559);
or U5711 (N_5711,N_1762,N_1487);
nand U5712 (N_5712,N_2952,N_235);
and U5713 (N_5713,N_219,N_671);
nand U5714 (N_5714,N_2339,N_2090);
nand U5715 (N_5715,N_210,N_1770);
nor U5716 (N_5716,N_2661,N_2679);
or U5717 (N_5717,N_1864,N_306);
or U5718 (N_5718,N_1824,N_2940);
nand U5719 (N_5719,N_964,N_2240);
or U5720 (N_5720,N_637,N_2001);
nor U5721 (N_5721,N_2021,N_137);
nor U5722 (N_5722,N_285,N_435);
and U5723 (N_5723,N_2588,N_1329);
nand U5724 (N_5724,N_1264,N_2752);
or U5725 (N_5725,N_2078,N_912);
nand U5726 (N_5726,N_1891,N_1670);
nand U5727 (N_5727,N_998,N_2757);
or U5728 (N_5728,N_347,N_1896);
or U5729 (N_5729,N_2988,N_2099);
or U5730 (N_5730,N_704,N_1255);
nor U5731 (N_5731,N_1484,N_2809);
or U5732 (N_5732,N_2006,N_2883);
or U5733 (N_5733,N_1910,N_631);
nand U5734 (N_5734,N_2528,N_215);
nand U5735 (N_5735,N_850,N_1168);
or U5736 (N_5736,N_1502,N_169);
and U5737 (N_5737,N_2420,N_127);
and U5738 (N_5738,N_2456,N_1377);
nor U5739 (N_5739,N_496,N_1864);
nor U5740 (N_5740,N_184,N_976);
nand U5741 (N_5741,N_1956,N_2644);
nand U5742 (N_5742,N_1,N_759);
nand U5743 (N_5743,N_2929,N_2952);
or U5744 (N_5744,N_2397,N_644);
nand U5745 (N_5745,N_2203,N_1243);
and U5746 (N_5746,N_1951,N_1696);
nand U5747 (N_5747,N_1130,N_425);
nor U5748 (N_5748,N_353,N_1713);
nor U5749 (N_5749,N_824,N_498);
nand U5750 (N_5750,N_321,N_4);
and U5751 (N_5751,N_300,N_2907);
and U5752 (N_5752,N_2240,N_2888);
and U5753 (N_5753,N_74,N_1482);
or U5754 (N_5754,N_778,N_193);
nand U5755 (N_5755,N_2962,N_1057);
nor U5756 (N_5756,N_1599,N_2691);
or U5757 (N_5757,N_150,N_536);
and U5758 (N_5758,N_1629,N_2650);
and U5759 (N_5759,N_1227,N_632);
and U5760 (N_5760,N_2661,N_1586);
and U5761 (N_5761,N_2213,N_2198);
nor U5762 (N_5762,N_366,N_1408);
nand U5763 (N_5763,N_1343,N_966);
nand U5764 (N_5764,N_2141,N_2531);
nand U5765 (N_5765,N_916,N_60);
or U5766 (N_5766,N_2027,N_1245);
nor U5767 (N_5767,N_2194,N_755);
nand U5768 (N_5768,N_2868,N_2738);
and U5769 (N_5769,N_2865,N_1388);
and U5770 (N_5770,N_2177,N_538);
nand U5771 (N_5771,N_978,N_391);
nand U5772 (N_5772,N_3,N_379);
nor U5773 (N_5773,N_818,N_2097);
and U5774 (N_5774,N_959,N_944);
nor U5775 (N_5775,N_1614,N_842);
and U5776 (N_5776,N_2946,N_270);
nand U5777 (N_5777,N_687,N_2981);
nand U5778 (N_5778,N_1616,N_1633);
nand U5779 (N_5779,N_2208,N_2307);
xor U5780 (N_5780,N_1703,N_2703);
nor U5781 (N_5781,N_797,N_308);
nor U5782 (N_5782,N_1247,N_2306);
nand U5783 (N_5783,N_1875,N_340);
or U5784 (N_5784,N_297,N_2110);
or U5785 (N_5785,N_1769,N_2317);
nand U5786 (N_5786,N_2296,N_774);
nand U5787 (N_5787,N_2914,N_2428);
nor U5788 (N_5788,N_2932,N_387);
or U5789 (N_5789,N_678,N_394);
nand U5790 (N_5790,N_1836,N_1118);
or U5791 (N_5791,N_2915,N_912);
nor U5792 (N_5792,N_2694,N_909);
nand U5793 (N_5793,N_1164,N_2210);
nand U5794 (N_5794,N_2918,N_1400);
nand U5795 (N_5795,N_1999,N_805);
nand U5796 (N_5796,N_1107,N_1968);
xor U5797 (N_5797,N_1171,N_65);
nor U5798 (N_5798,N_2492,N_2401);
nor U5799 (N_5799,N_2380,N_1278);
nand U5800 (N_5800,N_2847,N_2044);
nor U5801 (N_5801,N_1476,N_1948);
and U5802 (N_5802,N_654,N_1434);
or U5803 (N_5803,N_1511,N_2315);
nor U5804 (N_5804,N_1823,N_1418);
nor U5805 (N_5805,N_1102,N_193);
and U5806 (N_5806,N_1170,N_533);
and U5807 (N_5807,N_1671,N_2304);
and U5808 (N_5808,N_1724,N_715);
and U5809 (N_5809,N_1045,N_739);
xnor U5810 (N_5810,N_2008,N_399);
nor U5811 (N_5811,N_1273,N_1570);
nand U5812 (N_5812,N_2300,N_1296);
nand U5813 (N_5813,N_2030,N_1869);
and U5814 (N_5814,N_1896,N_908);
nand U5815 (N_5815,N_412,N_286);
and U5816 (N_5816,N_1247,N_500);
xnor U5817 (N_5817,N_1468,N_485);
and U5818 (N_5818,N_176,N_2244);
and U5819 (N_5819,N_1254,N_1080);
or U5820 (N_5820,N_2909,N_2042);
and U5821 (N_5821,N_1238,N_1211);
and U5822 (N_5822,N_2929,N_1035);
or U5823 (N_5823,N_1335,N_803);
nand U5824 (N_5824,N_269,N_1284);
nand U5825 (N_5825,N_259,N_2133);
and U5826 (N_5826,N_629,N_1809);
and U5827 (N_5827,N_1725,N_485);
nor U5828 (N_5828,N_614,N_730);
nor U5829 (N_5829,N_1354,N_1683);
or U5830 (N_5830,N_1344,N_9);
and U5831 (N_5831,N_539,N_2014);
and U5832 (N_5832,N_2681,N_784);
nor U5833 (N_5833,N_1830,N_1683);
and U5834 (N_5834,N_1949,N_1383);
nand U5835 (N_5835,N_376,N_1027);
and U5836 (N_5836,N_2075,N_376);
nor U5837 (N_5837,N_2685,N_2921);
or U5838 (N_5838,N_523,N_1926);
and U5839 (N_5839,N_68,N_1646);
nand U5840 (N_5840,N_1241,N_635);
nor U5841 (N_5841,N_2662,N_1744);
or U5842 (N_5842,N_1675,N_1799);
or U5843 (N_5843,N_2465,N_1546);
nand U5844 (N_5844,N_1657,N_500);
and U5845 (N_5845,N_2416,N_2334);
nand U5846 (N_5846,N_2046,N_2986);
and U5847 (N_5847,N_2822,N_679);
nor U5848 (N_5848,N_2868,N_2887);
nand U5849 (N_5849,N_2906,N_2373);
xnor U5850 (N_5850,N_2789,N_608);
or U5851 (N_5851,N_2155,N_2260);
and U5852 (N_5852,N_482,N_636);
or U5853 (N_5853,N_752,N_2130);
and U5854 (N_5854,N_1765,N_2045);
nand U5855 (N_5855,N_2670,N_2372);
nand U5856 (N_5856,N_2167,N_150);
xnor U5857 (N_5857,N_690,N_2286);
nand U5858 (N_5858,N_298,N_2477);
or U5859 (N_5859,N_1101,N_294);
and U5860 (N_5860,N_1920,N_136);
or U5861 (N_5861,N_961,N_1311);
nand U5862 (N_5862,N_2965,N_1453);
nand U5863 (N_5863,N_2527,N_2214);
nor U5864 (N_5864,N_250,N_296);
and U5865 (N_5865,N_2885,N_200);
nand U5866 (N_5866,N_2892,N_423);
nand U5867 (N_5867,N_2970,N_2652);
or U5868 (N_5868,N_571,N_1918);
and U5869 (N_5869,N_697,N_942);
nand U5870 (N_5870,N_735,N_2320);
nor U5871 (N_5871,N_1317,N_461);
nand U5872 (N_5872,N_747,N_63);
nor U5873 (N_5873,N_1643,N_383);
nand U5874 (N_5874,N_48,N_2944);
nand U5875 (N_5875,N_2612,N_1413);
or U5876 (N_5876,N_1108,N_1819);
or U5877 (N_5877,N_1648,N_1267);
nand U5878 (N_5878,N_839,N_538);
nor U5879 (N_5879,N_2803,N_1856);
nand U5880 (N_5880,N_1789,N_867);
nor U5881 (N_5881,N_2364,N_1670);
nor U5882 (N_5882,N_1887,N_2665);
or U5883 (N_5883,N_1608,N_2623);
nor U5884 (N_5884,N_511,N_767);
nor U5885 (N_5885,N_2704,N_1707);
or U5886 (N_5886,N_1033,N_2695);
and U5887 (N_5887,N_835,N_1134);
and U5888 (N_5888,N_2645,N_1245);
nand U5889 (N_5889,N_1807,N_1373);
nand U5890 (N_5890,N_1604,N_2504);
or U5891 (N_5891,N_1561,N_1761);
and U5892 (N_5892,N_803,N_1353);
nand U5893 (N_5893,N_2349,N_936);
or U5894 (N_5894,N_1594,N_1880);
nor U5895 (N_5895,N_2740,N_1156);
nor U5896 (N_5896,N_2513,N_399);
nor U5897 (N_5897,N_1062,N_1610);
or U5898 (N_5898,N_1529,N_2124);
or U5899 (N_5899,N_1940,N_566);
nand U5900 (N_5900,N_131,N_507);
nand U5901 (N_5901,N_1131,N_1722);
nand U5902 (N_5902,N_162,N_1761);
nor U5903 (N_5903,N_1500,N_816);
and U5904 (N_5904,N_785,N_1358);
nor U5905 (N_5905,N_1885,N_2115);
and U5906 (N_5906,N_101,N_969);
and U5907 (N_5907,N_336,N_1636);
nand U5908 (N_5908,N_1945,N_2464);
or U5909 (N_5909,N_1912,N_462);
nand U5910 (N_5910,N_812,N_704);
nor U5911 (N_5911,N_592,N_156);
nor U5912 (N_5912,N_2090,N_361);
nand U5913 (N_5913,N_1639,N_2539);
nor U5914 (N_5914,N_68,N_837);
nand U5915 (N_5915,N_643,N_2538);
nand U5916 (N_5916,N_1668,N_118);
nand U5917 (N_5917,N_1764,N_186);
and U5918 (N_5918,N_2447,N_1329);
nor U5919 (N_5919,N_2043,N_1656);
or U5920 (N_5920,N_386,N_1946);
or U5921 (N_5921,N_2974,N_362);
xor U5922 (N_5922,N_1671,N_1298);
and U5923 (N_5923,N_847,N_1485);
and U5924 (N_5924,N_546,N_2627);
nand U5925 (N_5925,N_1846,N_845);
or U5926 (N_5926,N_143,N_1576);
or U5927 (N_5927,N_1227,N_2381);
nor U5928 (N_5928,N_2414,N_1615);
nor U5929 (N_5929,N_294,N_1201);
nand U5930 (N_5930,N_118,N_1699);
and U5931 (N_5931,N_2636,N_1095);
or U5932 (N_5932,N_1902,N_2991);
xnor U5933 (N_5933,N_2078,N_2393);
and U5934 (N_5934,N_1240,N_2890);
and U5935 (N_5935,N_474,N_2221);
nor U5936 (N_5936,N_963,N_390);
nor U5937 (N_5937,N_2523,N_2346);
nor U5938 (N_5938,N_2647,N_2056);
and U5939 (N_5939,N_1973,N_2121);
and U5940 (N_5940,N_2519,N_906);
and U5941 (N_5941,N_930,N_721);
nand U5942 (N_5942,N_2111,N_1697);
and U5943 (N_5943,N_2074,N_2010);
and U5944 (N_5944,N_2466,N_1436);
nand U5945 (N_5945,N_37,N_845);
and U5946 (N_5946,N_2474,N_1307);
and U5947 (N_5947,N_2936,N_199);
and U5948 (N_5948,N_2188,N_1898);
nand U5949 (N_5949,N_469,N_1745);
nand U5950 (N_5950,N_327,N_858);
nand U5951 (N_5951,N_779,N_1287);
nand U5952 (N_5952,N_2628,N_2530);
or U5953 (N_5953,N_1929,N_468);
or U5954 (N_5954,N_747,N_997);
nand U5955 (N_5955,N_1018,N_346);
xnor U5956 (N_5956,N_2380,N_1391);
and U5957 (N_5957,N_1312,N_765);
and U5958 (N_5958,N_1893,N_49);
nand U5959 (N_5959,N_1215,N_862);
nand U5960 (N_5960,N_2687,N_1336);
nand U5961 (N_5961,N_814,N_2812);
nand U5962 (N_5962,N_557,N_2280);
nor U5963 (N_5963,N_1366,N_11);
nand U5964 (N_5964,N_410,N_2555);
xor U5965 (N_5965,N_2159,N_613);
nor U5966 (N_5966,N_165,N_550);
and U5967 (N_5967,N_1979,N_1757);
nor U5968 (N_5968,N_1345,N_2624);
nor U5969 (N_5969,N_2136,N_181);
and U5970 (N_5970,N_1849,N_2842);
nor U5971 (N_5971,N_380,N_1156);
or U5972 (N_5972,N_2527,N_1059);
or U5973 (N_5973,N_563,N_845);
and U5974 (N_5974,N_918,N_1362);
nand U5975 (N_5975,N_2551,N_214);
nor U5976 (N_5976,N_960,N_2812);
and U5977 (N_5977,N_44,N_684);
and U5978 (N_5978,N_1487,N_1836);
xor U5979 (N_5979,N_2455,N_254);
or U5980 (N_5980,N_2057,N_1481);
or U5981 (N_5981,N_2467,N_2814);
nor U5982 (N_5982,N_2,N_386);
and U5983 (N_5983,N_412,N_2892);
and U5984 (N_5984,N_940,N_1639);
and U5985 (N_5985,N_865,N_209);
and U5986 (N_5986,N_1119,N_842);
nor U5987 (N_5987,N_2780,N_2437);
or U5988 (N_5988,N_254,N_2086);
or U5989 (N_5989,N_1683,N_2759);
and U5990 (N_5990,N_1734,N_51);
nand U5991 (N_5991,N_1244,N_11);
and U5992 (N_5992,N_2520,N_1859);
or U5993 (N_5993,N_1872,N_1364);
nand U5994 (N_5994,N_1886,N_1481);
and U5995 (N_5995,N_761,N_1393);
nand U5996 (N_5996,N_701,N_1642);
or U5997 (N_5997,N_2612,N_2719);
nand U5998 (N_5998,N_553,N_2091);
or U5999 (N_5999,N_1748,N_684);
and U6000 (N_6000,N_4135,N_3712);
nor U6001 (N_6001,N_3432,N_3940);
or U6002 (N_6002,N_5965,N_5555);
and U6003 (N_6003,N_3498,N_4675);
nor U6004 (N_6004,N_4127,N_5286);
and U6005 (N_6005,N_5293,N_4833);
nor U6006 (N_6006,N_5117,N_5536);
and U6007 (N_6007,N_5948,N_4424);
or U6008 (N_6008,N_4259,N_4768);
or U6009 (N_6009,N_3177,N_5349);
or U6010 (N_6010,N_4270,N_3874);
nand U6011 (N_6011,N_3417,N_3830);
or U6012 (N_6012,N_3872,N_5709);
and U6013 (N_6013,N_3152,N_3221);
nor U6014 (N_6014,N_5999,N_4050);
or U6015 (N_6015,N_4927,N_4951);
or U6016 (N_6016,N_3572,N_5572);
xor U6017 (N_6017,N_3604,N_5579);
nor U6018 (N_6018,N_4885,N_3916);
nand U6019 (N_6019,N_5667,N_3378);
or U6020 (N_6020,N_5204,N_3174);
nor U6021 (N_6021,N_5791,N_5362);
and U6022 (N_6022,N_3541,N_5081);
nand U6023 (N_6023,N_5495,N_5372);
or U6024 (N_6024,N_5937,N_4996);
nor U6025 (N_6025,N_4484,N_3521);
nand U6026 (N_6026,N_3476,N_4958);
nand U6027 (N_6027,N_4246,N_5818);
and U6028 (N_6028,N_4065,N_4546);
or U6029 (N_6029,N_4783,N_4745);
nor U6030 (N_6030,N_5784,N_5632);
nand U6031 (N_6031,N_4898,N_5766);
or U6032 (N_6032,N_5812,N_5001);
xnor U6033 (N_6033,N_3974,N_5714);
or U6034 (N_6034,N_4925,N_4504);
nor U6035 (N_6035,N_4180,N_4812);
or U6036 (N_6036,N_4487,N_3074);
nand U6037 (N_6037,N_5663,N_4528);
nor U6038 (N_6038,N_5570,N_4470);
nor U6039 (N_6039,N_4143,N_5509);
nand U6040 (N_6040,N_3021,N_5887);
nor U6041 (N_6041,N_3900,N_5181);
nor U6042 (N_6042,N_4580,N_3215);
nor U6043 (N_6043,N_3799,N_4434);
or U6044 (N_6044,N_5244,N_5689);
or U6045 (N_6045,N_3389,N_4374);
nand U6046 (N_6046,N_4632,N_4463);
nor U6047 (N_6047,N_4878,N_5401);
and U6048 (N_6048,N_5422,N_4491);
or U6049 (N_6049,N_4837,N_5185);
or U6050 (N_6050,N_5206,N_3016);
nor U6051 (N_6051,N_3017,N_4333);
nand U6052 (N_6052,N_5939,N_4058);
and U6053 (N_6053,N_3092,N_5606);
nand U6054 (N_6054,N_5108,N_5620);
nor U6055 (N_6055,N_4765,N_3956);
or U6056 (N_6056,N_5135,N_5953);
nand U6057 (N_6057,N_4365,N_5592);
or U6058 (N_6058,N_5674,N_5496);
and U6059 (N_6059,N_3402,N_5727);
nor U6060 (N_6060,N_5154,N_4617);
and U6061 (N_6061,N_4334,N_4339);
nand U6062 (N_6062,N_3136,N_5546);
or U6063 (N_6063,N_4027,N_3965);
nand U6064 (N_6064,N_5945,N_5829);
and U6065 (N_6065,N_5563,N_5972);
and U6066 (N_6066,N_3514,N_3774);
or U6067 (N_6067,N_4167,N_5212);
or U6068 (N_6068,N_5788,N_3587);
and U6069 (N_6069,N_4151,N_4586);
nand U6070 (N_6070,N_3489,N_4798);
and U6071 (N_6071,N_5000,N_4896);
and U6072 (N_6072,N_3471,N_3596);
xor U6073 (N_6073,N_5958,N_3153);
nand U6074 (N_6074,N_5919,N_4413);
or U6075 (N_6075,N_4467,N_3276);
nand U6076 (N_6076,N_4822,N_3796);
or U6077 (N_6077,N_3628,N_3800);
and U6078 (N_6078,N_3725,N_3537);
nand U6079 (N_6079,N_5210,N_3454);
and U6080 (N_6080,N_4698,N_3788);
nand U6081 (N_6081,N_4049,N_3146);
nor U6082 (N_6082,N_5540,N_5989);
nand U6083 (N_6083,N_5378,N_5090);
nand U6084 (N_6084,N_4303,N_5267);
nor U6085 (N_6085,N_5957,N_5601);
and U6086 (N_6086,N_3337,N_4733);
nor U6087 (N_6087,N_5180,N_4124);
nor U6088 (N_6088,N_5797,N_5234);
nor U6089 (N_6089,N_3223,N_3381);
and U6090 (N_6090,N_3166,N_4851);
nor U6091 (N_6091,N_4763,N_3551);
or U6092 (N_6092,N_5823,N_4918);
or U6093 (N_6093,N_3559,N_3191);
nand U6094 (N_6094,N_5415,N_5824);
nor U6095 (N_6095,N_4978,N_5035);
and U6096 (N_6096,N_5089,N_3444);
nor U6097 (N_6097,N_5578,N_3039);
or U6098 (N_6098,N_5595,N_4796);
and U6099 (N_6099,N_5188,N_3782);
nand U6100 (N_6100,N_5789,N_5653);
or U6101 (N_6101,N_5107,N_4842);
nor U6102 (N_6102,N_3430,N_3895);
nand U6103 (N_6103,N_5202,N_3346);
and U6104 (N_6104,N_5409,N_5011);
nor U6105 (N_6105,N_4808,N_4015);
nor U6106 (N_6106,N_3996,N_5715);
or U6107 (N_6107,N_3170,N_3375);
or U6108 (N_6108,N_5608,N_4541);
and U6109 (N_6109,N_3745,N_3845);
and U6110 (N_6110,N_3431,N_3114);
nand U6111 (N_6111,N_3682,N_4806);
nand U6112 (N_6112,N_4899,N_4486);
nor U6113 (N_6113,N_3778,N_5101);
and U6114 (N_6114,N_4905,N_4582);
or U6115 (N_6115,N_4844,N_4686);
xnor U6116 (N_6116,N_3014,N_5682);
nor U6117 (N_6117,N_5058,N_3440);
and U6118 (N_6118,N_4681,N_3200);
or U6119 (N_6119,N_3140,N_5319);
or U6120 (N_6120,N_5190,N_3742);
or U6121 (N_6121,N_3544,N_4692);
and U6122 (N_6122,N_5661,N_4678);
and U6123 (N_6123,N_4077,N_3717);
nor U6124 (N_6124,N_4335,N_4048);
or U6125 (N_6125,N_3127,N_3423);
nor U6126 (N_6126,N_5839,N_3159);
nand U6127 (N_6127,N_3202,N_4940);
and U6128 (N_6128,N_4710,N_4262);
or U6129 (N_6129,N_3864,N_4642);
and U6130 (N_6130,N_3770,N_4980);
or U6131 (N_6131,N_3930,N_5560);
nand U6132 (N_6132,N_3945,N_5765);
nand U6133 (N_6133,N_3964,N_5253);
nand U6134 (N_6134,N_4316,N_3789);
and U6135 (N_6135,N_5314,N_5738);
or U6136 (N_6136,N_5329,N_4082);
nor U6137 (N_6137,N_3100,N_5406);
nand U6138 (N_6138,N_5488,N_5126);
and U6139 (N_6139,N_3819,N_5106);
nand U6140 (N_6140,N_4519,N_3411);
nor U6141 (N_6141,N_4538,N_5449);
or U6142 (N_6142,N_4079,N_3213);
nor U6143 (N_6143,N_3069,N_5398);
nor U6144 (N_6144,N_3731,N_5491);
nand U6145 (N_6145,N_4574,N_3009);
nand U6146 (N_6146,N_5208,N_5451);
nand U6147 (N_6147,N_4596,N_5828);
nor U6148 (N_6148,N_5342,N_5301);
and U6149 (N_6149,N_4581,N_3102);
nand U6150 (N_6150,N_3515,N_5760);
nand U6151 (N_6151,N_5443,N_5984);
and U6152 (N_6152,N_3231,N_5732);
nand U6153 (N_6153,N_4070,N_5150);
and U6154 (N_6154,N_5221,N_4430);
or U6155 (N_6155,N_5985,N_3635);
nor U6156 (N_6156,N_3856,N_3970);
nand U6157 (N_6157,N_5635,N_3990);
or U6158 (N_6158,N_5790,N_5102);
and U6159 (N_6159,N_3442,N_4527);
nand U6160 (N_6160,N_3485,N_4740);
xnor U6161 (N_6161,N_3007,N_3410);
nand U6162 (N_6162,N_4092,N_3612);
nor U6163 (N_6163,N_4067,N_3034);
nor U6164 (N_6164,N_5162,N_3068);
and U6165 (N_6165,N_3364,N_5975);
nor U6166 (N_6166,N_4201,N_5844);
nor U6167 (N_6167,N_5328,N_3578);
nand U6168 (N_6168,N_4739,N_5508);
and U6169 (N_6169,N_3333,N_5430);
nor U6170 (N_6170,N_4173,N_4697);
nor U6171 (N_6171,N_5607,N_5571);
nor U6172 (N_6172,N_3086,N_5435);
nor U6173 (N_6173,N_4123,N_5144);
and U6174 (N_6174,N_3022,N_4320);
nand U6175 (N_6175,N_3481,N_4199);
xnor U6176 (N_6176,N_5631,N_4002);
nor U6177 (N_6177,N_5029,N_4182);
or U6178 (N_6178,N_3010,N_3666);
or U6179 (N_6179,N_3334,N_4962);
nand U6180 (N_6180,N_3362,N_3447);
nand U6181 (N_6181,N_5980,N_4174);
and U6182 (N_6182,N_3941,N_5821);
or U6183 (N_6183,N_4074,N_4263);
or U6184 (N_6184,N_5633,N_3827);
nor U6185 (N_6185,N_4052,N_4257);
nor U6186 (N_6186,N_4026,N_3403);
or U6187 (N_6187,N_4440,N_4863);
nand U6188 (N_6188,N_3101,N_3663);
nand U6189 (N_6189,N_4886,N_3873);
nor U6190 (N_6190,N_5273,N_5193);
and U6191 (N_6191,N_3668,N_5955);
nand U6192 (N_6192,N_4395,N_5820);
and U6193 (N_6193,N_4777,N_5442);
and U6194 (N_6194,N_4228,N_5318);
nor U6195 (N_6195,N_4832,N_5785);
or U6196 (N_6196,N_4737,N_4023);
nand U6197 (N_6197,N_4144,N_3253);
nor U6198 (N_6198,N_4616,N_5615);
or U6199 (N_6199,N_3434,N_3386);
nor U6200 (N_6200,N_5122,N_3160);
nor U6201 (N_6201,N_5929,N_5490);
nor U6202 (N_6202,N_3658,N_4985);
or U6203 (N_6203,N_5325,N_5163);
or U6204 (N_6204,N_5337,N_5211);
and U6205 (N_6205,N_4785,N_3449);
or U6206 (N_6206,N_5581,N_5994);
xor U6207 (N_6207,N_3083,N_5634);
nor U6208 (N_6208,N_4933,N_3684);
nand U6209 (N_6209,N_4959,N_5598);
nand U6210 (N_6210,N_5454,N_5708);
nor U6211 (N_6211,N_4560,N_3395);
and U6212 (N_6212,N_3525,N_3883);
nand U6213 (N_6213,N_5596,N_5426);
and U6214 (N_6214,N_4480,N_3311);
or U6215 (N_6215,N_5446,N_4350);
or U6216 (N_6216,N_4129,N_5165);
nor U6217 (N_6217,N_5854,N_3312);
or U6218 (N_6218,N_4846,N_3791);
or U6219 (N_6219,N_3670,N_3407);
nand U6220 (N_6220,N_4375,N_5280);
or U6221 (N_6221,N_5209,N_5220);
or U6222 (N_6222,N_4630,N_3749);
or U6223 (N_6223,N_5177,N_5137);
and U6224 (N_6224,N_5848,N_4555);
or U6225 (N_6225,N_5648,N_3734);
nand U6226 (N_6226,N_3997,N_4829);
or U6227 (N_6227,N_3833,N_4108);
nand U6228 (N_6228,N_4782,N_5018);
nor U6229 (N_6229,N_5014,N_4914);
nand U6230 (N_6230,N_5323,N_4405);
and U6231 (N_6231,N_4272,N_3835);
nand U6232 (N_6232,N_4593,N_4404);
and U6233 (N_6233,N_5877,N_5248);
nand U6234 (N_6234,N_3660,N_4443);
and U6235 (N_6235,N_3580,N_5237);
nand U6236 (N_6236,N_5541,N_3932);
or U6237 (N_6237,N_4598,N_3831);
and U6238 (N_6238,N_4707,N_5838);
nand U6239 (N_6239,N_4028,N_3131);
and U6240 (N_6240,N_4475,N_4030);
and U6241 (N_6241,N_3249,N_3917);
or U6242 (N_6242,N_4521,N_5590);
nor U6243 (N_6243,N_3351,N_5853);
or U6244 (N_6244,N_3278,N_4153);
nor U6245 (N_6245,N_3005,N_3821);
or U6246 (N_6246,N_3356,N_5679);
and U6247 (N_6247,N_5187,N_4068);
or U6248 (N_6248,N_4104,N_4993);
or U6249 (N_6249,N_3575,N_5941);
nor U6250 (N_6250,N_3980,N_5735);
nand U6251 (N_6251,N_4034,N_5299);
and U6252 (N_6252,N_3121,N_3700);
nand U6253 (N_6253,N_3920,N_3163);
or U6254 (N_6254,N_5695,N_5678);
nor U6255 (N_6255,N_5006,N_3622);
and U6256 (N_6256,N_4539,N_4848);
nand U6257 (N_6257,N_3469,N_5340);
or U6258 (N_6258,N_4523,N_5739);
or U6259 (N_6259,N_4076,N_4826);
or U6260 (N_6260,N_3500,N_3438);
nor U6261 (N_6261,N_5025,N_5503);
and U6262 (N_6262,N_4654,N_5140);
nor U6263 (N_6263,N_5704,N_4513);
or U6264 (N_6264,N_3882,N_4853);
nand U6265 (N_6265,N_5915,N_5285);
and U6266 (N_6266,N_3505,N_3348);
or U6267 (N_6267,N_5189,N_3557);
or U6268 (N_6268,N_5525,N_3610);
and U6269 (N_6269,N_4786,N_4159);
or U6270 (N_6270,N_4684,N_3093);
or U6271 (N_6271,N_4738,N_4543);
nor U6272 (N_6272,N_4234,N_4024);
or U6273 (N_6273,N_5060,N_3655);
nand U6274 (N_6274,N_3301,N_5353);
or U6275 (N_6275,N_4845,N_3230);
and U6276 (N_6276,N_4530,N_4166);
and U6277 (N_6277,N_5145,N_3621);
nor U6278 (N_6278,N_4811,N_3192);
and U6279 (N_6279,N_5021,N_5920);
nor U6280 (N_6280,N_3891,N_3598);
nand U6281 (N_6281,N_3556,N_4767);
nor U6282 (N_6282,N_4668,N_5124);
or U6283 (N_6283,N_5071,N_5279);
nand U6284 (N_6284,N_5537,N_4998);
nor U6285 (N_6285,N_3590,N_4236);
or U6286 (N_6286,N_4855,N_3972);
nor U6287 (N_6287,N_3106,N_3816);
and U6288 (N_6288,N_4330,N_3764);
or U6289 (N_6289,N_5054,N_4273);
or U6290 (N_6290,N_5557,N_5246);
nand U6291 (N_6291,N_4648,N_4468);
nand U6292 (N_6292,N_3851,N_5918);
or U6293 (N_6293,N_3099,N_5313);
or U6294 (N_6294,N_5688,N_5680);
nor U6295 (N_6295,N_4231,N_5917);
and U6296 (N_6296,N_3737,N_4305);
and U6297 (N_6297,N_5093,N_4906);
or U6298 (N_6298,N_4436,N_5482);
and U6299 (N_6299,N_5408,N_5448);
and U6300 (N_6300,N_3063,N_3360);
or U6301 (N_6301,N_5074,N_3907);
nor U6302 (N_6302,N_4396,N_4354);
nand U6303 (N_6303,N_4017,N_4761);
or U6304 (N_6304,N_3087,N_3052);
and U6305 (N_6305,N_5183,N_4992);
or U6306 (N_6306,N_4492,N_3549);
and U6307 (N_6307,N_5775,N_4132);
nor U6308 (N_6308,N_3728,N_5859);
nand U6309 (N_6309,N_5973,N_4526);
nand U6310 (N_6310,N_3340,N_5130);
and U6311 (N_6311,N_3280,N_3067);
and U6312 (N_6312,N_3524,N_5559);
nor U6313 (N_6313,N_3815,N_5758);
nor U6314 (N_6314,N_5665,N_5042);
or U6315 (N_6315,N_5959,N_4990);
or U6316 (N_6316,N_3397,N_3577);
nor U6317 (N_6317,N_3785,N_4847);
nand U6318 (N_6318,N_3429,N_5756);
and U6319 (N_6319,N_4974,N_5666);
or U6320 (N_6320,N_4329,N_3618);
or U6321 (N_6321,N_3164,N_3848);
and U6322 (N_6322,N_4731,N_5365);
nor U6323 (N_6323,N_4194,N_3415);
nand U6324 (N_6324,N_4912,N_4105);
nor U6325 (N_6325,N_5677,N_3295);
or U6326 (N_6326,N_5094,N_5773);
and U6327 (N_6327,N_5075,N_5764);
nand U6328 (N_6328,N_4016,N_5277);
or U6329 (N_6329,N_5305,N_4895);
nand U6330 (N_6330,N_4053,N_4340);
and U6331 (N_6331,N_3862,N_3228);
nor U6332 (N_6332,N_5876,N_3661);
or U6333 (N_6333,N_4455,N_4469);
nor U6334 (N_6334,N_4387,N_4169);
nand U6335 (N_6335,N_5338,N_4864);
or U6336 (N_6336,N_3188,N_4667);
or U6337 (N_6337,N_5461,N_3656);
nor U6338 (N_6338,N_5477,N_4266);
or U6339 (N_6339,N_3241,N_4061);
nor U6340 (N_6340,N_5425,N_5065);
nor U6341 (N_6341,N_5476,N_3025);
or U6342 (N_6342,N_5396,N_5683);
nand U6343 (N_6343,N_3341,N_3750);
and U6344 (N_6344,N_3269,N_5888);
and U6345 (N_6345,N_5669,N_3533);
and U6346 (N_6346,N_3171,N_3765);
nor U6347 (N_6347,N_5479,N_3755);
nand U6348 (N_6348,N_3975,N_4321);
and U6349 (N_6349,N_4422,N_5676);
nor U6350 (N_6350,N_5389,N_4827);
and U6351 (N_6351,N_3775,N_3463);
nor U6352 (N_6352,N_5229,N_4009);
xor U6353 (N_6353,N_4584,N_4131);
or U6354 (N_6354,N_5091,N_4022);
nand U6355 (N_6355,N_5597,N_4577);
or U6356 (N_6356,N_5049,N_3244);
nor U6357 (N_6357,N_4046,N_5961);
nand U6358 (N_6358,N_5291,N_5306);
and U6359 (N_6359,N_4602,N_4877);
nor U6360 (N_6360,N_4781,N_4306);
or U6361 (N_6361,N_4136,N_3828);
nor U6362 (N_6362,N_5174,N_4505);
and U6363 (N_6363,N_3178,N_5936);
nor U6364 (N_6364,N_5518,N_5630);
or U6365 (N_6365,N_3936,N_5110);
nor U6366 (N_6366,N_4545,N_3133);
and U6367 (N_6367,N_3446,N_5685);
and U6368 (N_6368,N_3421,N_3189);
and U6369 (N_6369,N_5528,N_3169);
nand U6370 (N_6370,N_5614,N_3124);
or U6371 (N_6371,N_5033,N_5825);
xnor U6372 (N_6372,N_4109,N_3150);
nand U6373 (N_6373,N_5830,N_5690);
or U6374 (N_6374,N_3287,N_4247);
and U6375 (N_6375,N_3075,N_3772);
nand U6376 (N_6376,N_4884,N_3272);
nand U6377 (N_6377,N_5740,N_3482);
nand U6378 (N_6378,N_4724,N_4639);
and U6379 (N_6379,N_4762,N_3018);
and U6380 (N_6380,N_4479,N_4566);
xnor U6381 (N_6381,N_3125,N_3232);
nor U6382 (N_6382,N_3927,N_3739);
or U6383 (N_6383,N_4036,N_4854);
nand U6384 (N_6384,N_3355,N_4702);
nor U6385 (N_6385,N_4482,N_5718);
or U6386 (N_6386,N_3490,N_3255);
nor U6387 (N_6387,N_3023,N_5628);
nor U6388 (N_6388,N_3605,N_5742);
nand U6389 (N_6389,N_4943,N_5658);
and U6390 (N_6390,N_4618,N_5966);
nand U6391 (N_6391,N_5483,N_5768);
nand U6392 (N_6392,N_5651,N_4571);
or U6393 (N_6393,N_5890,N_5886);
or U6394 (N_6394,N_3292,N_3766);
and U6395 (N_6395,N_4759,N_5127);
and U6396 (N_6396,N_4902,N_4881);
xor U6397 (N_6397,N_5971,N_3303);
and U6398 (N_6398,N_5321,N_4662);
nor U6399 (N_6399,N_3879,N_4032);
and U6400 (N_6400,N_5979,N_4597);
or U6401 (N_6401,N_4924,N_5645);
nor U6402 (N_6402,N_4267,N_3561);
or U6403 (N_6403,N_3894,N_5179);
and U6404 (N_6404,N_4919,N_3510);
and U6405 (N_6405,N_3723,N_4307);
or U6406 (N_6406,N_3155,N_4578);
xor U6407 (N_6407,N_4197,N_3090);
and U6408 (N_6408,N_3497,N_5410);
and U6409 (N_6409,N_4290,N_4410);
nand U6410 (N_6410,N_3646,N_5529);
nand U6411 (N_6411,N_5316,N_3871);
and U6412 (N_6412,N_5088,N_4154);
nor U6413 (N_6413,N_4145,N_4351);
and U6414 (N_6414,N_3844,N_4287);
or U6415 (N_6415,N_4331,N_3877);
nor U6416 (N_6416,N_4198,N_5250);
nor U6417 (N_6417,N_5473,N_3012);
nor U6418 (N_6418,N_3644,N_5346);
or U6419 (N_6419,N_5573,N_4458);
nor U6420 (N_6420,N_5474,N_3527);
and U6421 (N_6421,N_4368,N_3953);
and U6422 (N_6422,N_4400,N_4212);
nand U6423 (N_6423,N_5402,N_4549);
or U6424 (N_6424,N_4779,N_4152);
nor U6425 (N_6425,N_5170,N_3686);
nand U6426 (N_6426,N_3456,N_4726);
nand U6427 (N_6427,N_3371,N_4908);
nor U6428 (N_6428,N_5594,N_5885);
and U6429 (N_6429,N_3404,N_3047);
or U6430 (N_6430,N_5431,N_4947);
and U6431 (N_6431,N_3239,N_4117);
or U6432 (N_6432,N_3302,N_4183);
or U6433 (N_6433,N_5567,N_5743);
or U6434 (N_6434,N_3839,N_5687);
and U6435 (N_6435,N_4444,N_4086);
nor U6436 (N_6436,N_3809,N_4394);
or U6437 (N_6437,N_3522,N_3004);
nor U6438 (N_6438,N_4588,N_4298);
nor U6439 (N_6439,N_4789,N_3358);
nand U6440 (N_6440,N_5882,N_3671);
and U6441 (N_6441,N_4857,N_3992);
and U6442 (N_6442,N_4674,N_4483);
nor U6443 (N_6443,N_4465,N_5307);
nor U6444 (N_6444,N_4706,N_5550);
and U6445 (N_6445,N_3857,N_5935);
nand U6446 (N_6446,N_3715,N_3633);
nor U6447 (N_6447,N_4942,N_5502);
nand U6448 (N_6448,N_3433,N_4497);
nor U6449 (N_6449,N_5734,N_4606);
and U6450 (N_6450,N_3642,N_4012);
and U6451 (N_6451,N_5215,N_4242);
nor U6452 (N_6452,N_3252,N_3662);
nor U6453 (N_6453,N_5545,N_3049);
or U6454 (N_6454,N_5226,N_3795);
nand U6455 (N_6455,N_5519,N_5048);
nand U6456 (N_6456,N_3647,N_5281);
or U6457 (N_6457,N_4561,N_3754);
nand U6458 (N_6458,N_4670,N_5061);
and U6459 (N_6459,N_3254,N_4901);
and U6460 (N_6460,N_3842,N_3902);
and U6461 (N_6461,N_5752,N_4608);
or U6462 (N_6462,N_3070,N_5388);
nand U6463 (N_6463,N_4661,N_5681);
or U6464 (N_6464,N_5224,N_3973);
nand U6465 (N_6465,N_5111,N_5374);
and U6466 (N_6466,N_5288,N_4103);
or U6467 (N_6467,N_3690,N_3511);
nor U6468 (N_6468,N_3290,N_5118);
or U6469 (N_6469,N_5933,N_5112);
or U6470 (N_6470,N_3582,N_4031);
xor U6471 (N_6471,N_3692,N_5393);
or U6472 (N_6472,N_5390,N_5387);
and U6473 (N_6473,N_5171,N_5257);
nor U6474 (N_6474,N_5263,N_4817);
nand U6475 (N_6475,N_5650,N_4532);
nand U6476 (N_6476,N_3616,N_4386);
or U6477 (N_6477,N_5701,N_3986);
and U6478 (N_6478,N_4402,N_3983);
nor U6479 (N_6479,N_4338,N_4357);
nor U6480 (N_6480,N_4415,N_4148);
nand U6481 (N_6481,N_3840,N_5833);
or U6482 (N_6482,N_5960,N_3954);
nand U6483 (N_6483,N_5005,N_4534);
and U6484 (N_6484,N_3284,N_4872);
nor U6485 (N_6485,N_3260,N_3103);
and U6486 (N_6486,N_3190,N_4900);
or U6487 (N_6487,N_3571,N_3675);
nor U6488 (N_6488,N_3236,N_3905);
nor U6489 (N_6489,N_3137,N_5097);
nor U6490 (N_6490,N_3310,N_5618);
nand U6491 (N_6491,N_3735,N_3904);
or U6492 (N_6492,N_5897,N_4791);
nor U6493 (N_6493,N_4051,N_3787);
nor U6494 (N_6494,N_4909,N_3747);
and U6495 (N_6495,N_4965,N_5078);
and U6496 (N_6496,N_4130,N_5274);
nor U6497 (N_6497,N_3256,N_4713);
or U6498 (N_6498,N_3968,N_4510);
and U6499 (N_6499,N_3400,N_4435);
or U6500 (N_6500,N_3989,N_5691);
or U6501 (N_6501,N_4891,N_4647);
nand U6502 (N_6502,N_5535,N_4544);
and U6503 (N_6503,N_4213,N_5515);
nor U6504 (N_6504,N_4858,N_3299);
or U6505 (N_6505,N_4312,N_5024);
nand U6506 (N_6506,N_5022,N_3516);
nor U6507 (N_6507,N_5862,N_4818);
or U6508 (N_6508,N_4861,N_5672);
nand U6509 (N_6509,N_3792,N_4416);
or U6510 (N_6510,N_4917,N_4594);
and U6511 (N_6511,N_5298,N_3834);
nand U6512 (N_6512,N_3752,N_3377);
and U6513 (N_6513,N_5407,N_4114);
nand U6514 (N_6514,N_4230,N_3359);
and U6515 (N_6515,N_4520,N_3261);
and U6516 (N_6516,N_4188,N_5465);
nor U6517 (N_6517,N_3636,N_5400);
xor U6518 (N_6518,N_4776,N_5218);
or U6519 (N_6519,N_5798,N_4716);
or U6520 (N_6520,N_3592,N_4084);
nand U6521 (N_6521,N_5591,N_5433);
and U6522 (N_6522,N_3803,N_4205);
and U6523 (N_6523,N_4203,N_5087);
or U6524 (N_6524,N_3824,N_4669);
or U6525 (N_6525,N_5148,N_5901);
or U6526 (N_6526,N_3391,N_5511);
and U6527 (N_6527,N_5892,N_5439);
nor U6528 (N_6528,N_5282,N_5238);
and U6529 (N_6529,N_3654,N_5192);
or U6530 (N_6530,N_4454,N_4141);
and U6531 (N_6531,N_5312,N_4627);
and U6532 (N_6532,N_4437,N_5754);
or U6533 (N_6533,N_3467,N_4380);
or U6534 (N_6534,N_3625,N_3499);
or U6535 (N_6535,N_4433,N_5982);
and U6536 (N_6536,N_4446,N_5807);
or U6537 (N_6537,N_4836,N_4353);
nand U6538 (N_6538,N_5719,N_4268);
nor U6539 (N_6539,N_3643,N_3426);
or U6540 (N_6540,N_3638,N_4216);
and U6541 (N_6541,N_5796,N_4953);
and U6542 (N_6542,N_5549,N_3036);
and U6543 (N_6543,N_4873,N_4880);
nand U6544 (N_6544,N_5462,N_5946);
xor U6545 (N_6545,N_5684,N_3266);
nor U6546 (N_6546,N_4252,N_3242);
and U6547 (N_6547,N_5836,N_5532);
and U6548 (N_6548,N_5611,N_5134);
and U6549 (N_6549,N_4680,N_4072);
nor U6550 (N_6550,N_4831,N_4189);
nand U6551 (N_6551,N_3123,N_4223);
and U6552 (N_6552,N_3852,N_4042);
nor U6553 (N_6553,N_5456,N_4421);
and U6554 (N_6554,N_3088,N_3061);
nand U6555 (N_6555,N_4862,N_4770);
and U6556 (N_6556,N_5904,N_4494);
nand U6557 (N_6557,N_3172,N_5038);
or U6558 (N_6558,N_5548,N_5205);
and U6559 (N_6559,N_3144,N_3441);
and U6560 (N_6560,N_3229,N_5200);
nand U6561 (N_6561,N_5940,N_4461);
nand U6562 (N_6562,N_4773,N_5383);
nor U6563 (N_6563,N_5832,N_3318);
and U6564 (N_6564,N_3630,N_3929);
nand U6565 (N_6565,N_4349,N_3427);
and U6566 (N_6566,N_3680,N_4401);
or U6567 (N_6567,N_3767,N_5417);
and U6568 (N_6568,N_3637,N_5186);
or U6569 (N_6569,N_3797,N_4757);
nand U6570 (N_6570,N_5706,N_5334);
and U6571 (N_6571,N_5817,N_4645);
nor U6572 (N_6572,N_4575,N_5428);
nor U6573 (N_6573,N_4346,N_3027);
nor U6574 (N_6574,N_3769,N_3128);
nand U6575 (N_6575,N_3270,N_4619);
nor U6576 (N_6576,N_5032,N_3977);
or U6577 (N_6577,N_3032,N_5379);
nand U6578 (N_6578,N_4984,N_5543);
or U6579 (N_6579,N_4313,N_3387);
xnor U6580 (N_6580,N_4687,N_4816);
nor U6581 (N_6581,N_3711,N_4553);
and U6582 (N_6582,N_3494,N_5057);
and U6583 (N_6583,N_5753,N_5194);
nor U6584 (N_6584,N_3560,N_3187);
or U6585 (N_6585,N_4317,N_4643);
or U6586 (N_6586,N_4866,N_3705);
nor U6587 (N_6587,N_4677,N_4429);
nor U6588 (N_6588,N_3673,N_5745);
and U6589 (N_6589,N_5779,N_4176);
nand U6590 (N_6590,N_5156,N_3563);
nor U6591 (N_6591,N_5556,N_3573);
nand U6592 (N_6592,N_4038,N_5602);
nor U6593 (N_6593,N_4168,N_4477);
nor U6594 (N_6594,N_3345,N_4441);
and U6595 (N_6595,N_3217,N_4025);
and U6596 (N_6596,N_4366,N_3939);
or U6597 (N_6597,N_3714,N_4623);
nor U6598 (N_6598,N_3041,N_4033);
or U6599 (N_6599,N_4514,N_4903);
nand U6600 (N_6600,N_4550,N_4099);
nand U6601 (N_6601,N_4308,N_5031);
nand U6602 (N_6602,N_4653,N_4628);
nand U6603 (N_6603,N_3259,N_4381);
nand U6604 (N_6604,N_4403,N_3687);
or U6605 (N_6605,N_3376,N_3384);
nor U6606 (N_6606,N_4235,N_5816);
or U6607 (N_6607,N_5642,N_4088);
and U6608 (N_6608,N_5558,N_5243);
or U6609 (N_6609,N_4558,N_5309);
nor U6610 (N_6610,N_5644,N_4452);
nor U6611 (N_6611,N_4913,N_5582);
nand U6612 (N_6612,N_3222,N_3003);
nor U6613 (N_6613,N_5027,N_4202);
or U6614 (N_6614,N_4195,N_4932);
nand U6615 (N_6615,N_4080,N_5046);
and U6616 (N_6616,N_5991,N_3161);
nor U6617 (N_6617,N_5213,N_4251);
or U6618 (N_6618,N_4464,N_3509);
and U6619 (N_6619,N_5007,N_3205);
nor U6620 (N_6620,N_4910,N_4709);
nand U6621 (N_6621,N_3554,N_5143);
nor U6622 (N_6622,N_4283,N_4442);
nand U6623 (N_6623,N_5260,N_3282);
nand U6624 (N_6624,N_3555,N_3898);
or U6625 (N_6625,N_5988,N_4035);
nand U6626 (N_6626,N_5009,N_5343);
or U6627 (N_6627,N_4704,N_3777);
nor U6628 (N_6628,N_3491,N_3001);
and U6629 (N_6629,N_3059,N_4948);
or U6630 (N_6630,N_5178,N_4839);
xor U6631 (N_6631,N_4301,N_4809);
nor U6632 (N_6632,N_5245,N_5770);
or U6633 (N_6633,N_4241,N_5710);
xnor U6634 (N_6634,N_5802,N_5944);
nand U6635 (N_6635,N_3903,N_5840);
and U6636 (N_6636,N_5335,N_4841);
and U6637 (N_6637,N_4221,N_5066);
nand U6638 (N_6638,N_5405,N_3349);
nand U6639 (N_6639,N_3548,N_3042);
nand U6640 (N_6640,N_5157,N_3724);
nand U6641 (N_6641,N_3279,N_4986);
nand U6642 (N_6642,N_4473,N_4171);
or U6643 (N_6643,N_3506,N_4249);
nor U6644 (N_6644,N_3015,N_3323);
and U6645 (N_6645,N_3112,N_5172);
and U6646 (N_6646,N_3756,N_4218);
nand U6647 (N_6647,N_5331,N_5438);
and U6648 (N_6648,N_5819,N_3969);
or U6649 (N_6649,N_3118,N_4660);
nor U6650 (N_6650,N_5486,N_5616);
nand U6651 (N_6651,N_3428,N_4498);
nand U6652 (N_6652,N_5736,N_3165);
or U6653 (N_6653,N_3263,N_4794);
nor U6654 (N_6654,N_4744,N_4000);
or U6655 (N_6655,N_3854,N_4447);
nor U6656 (N_6656,N_5656,N_5911);
or U6657 (N_6657,N_3031,N_5705);
and U6658 (N_6658,N_3045,N_3392);
nor U6659 (N_6659,N_4659,N_5153);
nand U6660 (N_6660,N_3979,N_5969);
or U6661 (N_6661,N_4499,N_5943);
or U6662 (N_6662,N_3949,N_5921);
or U6663 (N_6663,N_5196,N_3810);
nand U6664 (N_6664,N_3987,N_4944);
nand U6665 (N_6665,N_5039,N_5303);
xnor U6666 (N_6666,N_4922,N_4609);
nor U6667 (N_6667,N_3496,N_3024);
nand U6668 (N_6668,N_4823,N_4690);
or U6669 (N_6669,N_4694,N_4325);
and U6670 (N_6670,N_3113,N_5534);
or U6671 (N_6671,N_4097,N_3285);
and U6672 (N_6672,N_3363,N_4299);
and U6673 (N_6673,N_5030,N_4258);
or U6674 (N_6674,N_4010,N_4592);
or U6675 (N_6675,N_4689,N_3425);
and U6676 (N_6676,N_5397,N_5175);
nand U6677 (N_6677,N_4208,N_3274);
and U6678 (N_6678,N_4233,N_3935);
and U6679 (N_6679,N_5239,N_5302);
nor U6680 (N_6680,N_5737,N_3327);
nand U6681 (N_6681,N_3855,N_5623);
nor U6682 (N_6682,N_5670,N_3218);
nand U6683 (N_6683,N_5772,N_5055);
nor U6684 (N_6684,N_5777,N_3892);
and U6685 (N_6685,N_5498,N_3072);
nor U6686 (N_6686,N_4559,N_3305);
xnor U6687 (N_6687,N_3841,N_4843);
and U6688 (N_6688,N_3703,N_4004);
and U6689 (N_6689,N_5427,N_5227);
nor U6690 (N_6690,N_3464,N_5881);
nor U6691 (N_6691,N_5925,N_3727);
nand U6692 (N_6692,N_5880,N_4466);
or U6693 (N_6693,N_5421,N_3508);
nor U6694 (N_6694,N_5506,N_3918);
or U6695 (N_6695,N_5721,N_4911);
and U6696 (N_6696,N_5809,N_4288);
nor U6697 (N_6697,N_3529,N_3488);
or U6698 (N_6698,N_4364,N_4390);
nand U6699 (N_6699,N_5808,N_3084);
or U6700 (N_6700,N_5468,N_4140);
and U6701 (N_6701,N_4705,N_5712);
nand U6702 (N_6702,N_3385,N_3098);
nor U6703 (N_6703,N_3419,N_4624);
and U6704 (N_6704,N_3503,N_4018);
or U6705 (N_6705,N_3773,N_3206);
nand U6706 (N_6706,N_5489,N_4797);
nand U6707 (N_6707,N_4314,N_3600);
or U6708 (N_6708,N_3458,N_4755);
nor U6709 (N_6709,N_5641,N_3958);
or U6710 (N_6710,N_3307,N_3388);
and U6711 (N_6711,N_5861,N_4968);
nor U6712 (N_6712,N_3688,N_4274);
or U6713 (N_6713,N_4883,N_4063);
nand U6714 (N_6714,N_4742,N_5585);
nand U6715 (N_6715,N_4815,N_3353);
nor U6716 (N_6716,N_5893,N_3736);
nand U6717 (N_6717,N_3568,N_3860);
or U6718 (N_6718,N_4859,N_3418);
nor U6719 (N_6719,N_5698,N_4576);
nor U6720 (N_6720,N_5017,N_4547);
and U6721 (N_6721,N_3967,N_3639);
nor U6722 (N_6722,N_3693,N_3293);
and U6723 (N_6723,N_5993,N_3151);
nor U6724 (N_6724,N_5128,N_3240);
and U6725 (N_6725,N_4098,N_4725);
and U6726 (N_6726,N_3317,N_5748);
nand U6727 (N_6727,N_5671,N_4193);
and U6728 (N_6728,N_5843,N_5133);
nor U6729 (N_6729,N_3976,N_4337);
nand U6730 (N_6730,N_4254,N_5849);
nor U6731 (N_6731,N_5330,N_4326);
or U6732 (N_6732,N_4296,N_4734);
xnor U6733 (N_6733,N_3350,N_3077);
nor U6734 (N_6734,N_3650,N_3814);
nor U6735 (N_6735,N_3320,N_5584);
or U6736 (N_6736,N_5173,N_3565);
nor U6737 (N_6737,N_4634,N_3479);
nand U6738 (N_6738,N_5716,N_5168);
nor U6739 (N_6739,N_4471,N_4923);
nand U6740 (N_6740,N_4711,N_4868);
nor U6741 (N_6741,N_4887,N_5242);
nor U6742 (N_6742,N_4569,N_4315);
or U6743 (N_6743,N_5787,N_4780);
and U6744 (N_6744,N_3910,N_4332);
nand U6745 (N_6745,N_5485,N_4345);
or U6746 (N_6746,N_3876,N_3550);
and U6747 (N_6747,N_4209,N_5095);
and U6748 (N_6748,N_4322,N_4834);
nor U6749 (N_6749,N_5553,N_4972);
nor U6750 (N_6750,N_4930,N_3858);
and U6751 (N_6751,N_3947,N_3271);
and U6752 (N_6752,N_3611,N_5799);
or U6753 (N_6753,N_3943,N_4860);
nor U6754 (N_6754,N_5504,N_4790);
and U6755 (N_6755,N_5040,N_4445);
nor U6756 (N_6756,N_4459,N_5310);
nand U6757 (N_6757,N_4453,N_3002);
nor U6758 (N_6758,N_4756,N_3056);
nor U6759 (N_6759,N_5416,N_5161);
or U6760 (N_6760,N_5668,N_4146);
nor U6761 (N_6761,N_5868,N_4120);
nor U6762 (N_6762,N_5922,N_4075);
or U6763 (N_6763,N_4535,N_3863);
or U6764 (N_6764,N_4775,N_3719);
nor U6765 (N_6765,N_4054,N_5588);
nor U6766 (N_6766,N_5894,N_5199);
nand U6767 (N_6767,N_5036,N_4253);
and U6768 (N_6768,N_5837,N_3547);
and U6769 (N_6769,N_5513,N_4937);
nand U6770 (N_6770,N_4936,N_5516);
or U6771 (N_6771,N_4294,N_4211);
nand U6772 (N_6772,N_3370,N_3694);
and U6773 (N_6773,N_4456,N_3435);
nand U6774 (N_6774,N_5441,N_5103);
or U6775 (N_6775,N_4754,N_3094);
nand U6776 (N_6776,N_5744,N_3546);
or U6777 (N_6777,N_4006,N_5453);
or U6778 (N_6778,N_3233,N_3536);
nand U6779 (N_6779,N_4629,N_3201);
or U6780 (N_6780,N_5564,N_3053);
and U6781 (N_6781,N_3322,N_3372);
nor U6782 (N_6782,N_5577,N_4055);
nor U6783 (N_6783,N_5345,N_4751);
and U6784 (N_6784,N_5382,N_4935);
or U6785 (N_6785,N_3768,N_3283);
and U6786 (N_6786,N_5121,N_4344);
or U6787 (N_6787,N_3297,N_4393);
and U6788 (N_6788,N_3944,N_5207);
nand U6789 (N_6789,N_5755,N_3881);
or U6790 (N_6790,N_3837,N_5255);
nor U6791 (N_6791,N_3665,N_3273);
and U6792 (N_6792,N_5891,N_4799);
or U6793 (N_6793,N_5654,N_5523);
nor U6794 (N_6794,N_3597,N_3523);
and U6795 (N_6795,N_5587,N_5741);
or U6796 (N_6796,N_3591,N_4496);
and U6797 (N_6797,N_3082,N_5864);
nand U6798 (N_6798,N_3566,N_5324);
nand U6799 (N_6799,N_4570,N_4931);
nor U6800 (N_6800,N_5804,N_5514);
and U6801 (N_6801,N_5652,N_3707);
nor U6802 (N_6802,N_4938,N_3710);
or U6803 (N_6803,N_4795,N_3176);
and U6804 (N_6804,N_3982,N_4342);
and U6805 (N_6805,N_3651,N_3950);
nand U6806 (N_6806,N_5947,N_3535);
and U6807 (N_6807,N_5729,N_3139);
or U6808 (N_6808,N_3994,N_3838);
and U6809 (N_6809,N_4388,N_5010);
nor U6810 (N_6810,N_3942,N_3382);
nand U6811 (N_6811,N_3532,N_5419);
nand U6812 (N_6812,N_3235,N_4425);
nor U6813 (N_6813,N_4769,N_5012);
or U6814 (N_6814,N_3478,N_5347);
nor U6815 (N_6815,N_3859,N_4341);
and U6816 (N_6816,N_4243,N_4838);
and U6817 (N_6817,N_3802,N_4150);
or U6818 (N_6818,N_4222,N_4852);
nor U6819 (N_6819,N_5463,N_3617);
and U6820 (N_6820,N_4073,N_4107);
nand U6821 (N_6821,N_3264,N_5327);
nor U6822 (N_6822,N_4650,N_5050);
nor U6823 (N_6823,N_5037,N_4728);
nand U6824 (N_6824,N_4495,N_3606);
nand U6825 (N_6825,N_4164,N_4760);
nor U6826 (N_6826,N_5236,N_3366);
or U6827 (N_6827,N_5909,N_5776);
and U6828 (N_6828,N_5903,N_5659);
nand U6829 (N_6829,N_4110,N_3607);
nor U6830 (N_6830,N_3495,N_5934);
or U6831 (N_6831,N_5505,N_3237);
or U6832 (N_6832,N_4814,N_4655);
and U6833 (N_6833,N_5080,N_3343);
or U6834 (N_6834,N_4157,N_5169);
and U6835 (N_6835,N_5300,N_3401);
xnor U6836 (N_6836,N_3294,N_4115);
and U6837 (N_6837,N_5045,N_5013);
or U6838 (N_6838,N_5530,N_4369);
or U6839 (N_6839,N_3619,N_3288);
or U6840 (N_6840,N_5831,N_5637);
nand U6841 (N_6841,N_3439,N_3659);
nand U6842 (N_6842,N_5411,N_4792);
or U6843 (N_6843,N_5230,N_4133);
nand U6844 (N_6844,N_5749,N_4890);
or U6845 (N_6845,N_3689,N_4995);
and U6846 (N_6846,N_5942,N_5850);
nand U6847 (N_6847,N_3048,N_5247);
nor U6848 (N_6848,N_4367,N_3695);
or U6849 (N_6849,N_4774,N_5160);
nor U6850 (N_6850,N_4476,N_4870);
nand U6851 (N_6851,N_5129,N_5501);
or U6852 (N_6852,N_3399,N_5912);
nor U6853 (N_6853,N_5520,N_3316);
nor U6854 (N_6854,N_5367,N_5954);
nand U6855 (N_6855,N_3373,N_4793);
and U6856 (N_6856,N_3985,N_5762);
nand U6857 (N_6857,N_4572,N_4044);
or U6858 (N_6858,N_5015,N_4610);
nand U6859 (N_6859,N_3971,N_4640);
nand U6860 (N_6860,N_3313,N_5198);
nor U6861 (N_6861,N_3595,N_5311);
nor U6862 (N_6862,N_4106,N_4971);
or U6863 (N_6863,N_4752,N_5377);
nand U6864 (N_6864,N_3887,N_5951);
or U6865 (N_6865,N_5475,N_3538);
nor U6866 (N_6866,N_3149,N_3286);
nor U6867 (N_6867,N_3216,N_3832);
nor U6868 (N_6868,N_4605,N_3332);
or U6869 (N_6869,N_3586,N_4502);
and U6870 (N_6870,N_5610,N_3609);
nor U6871 (N_6871,N_3908,N_4892);
nor U6872 (N_6872,N_3424,N_3296);
nand U6873 (N_6873,N_3208,N_3038);
and U6874 (N_6874,N_3798,N_3925);
nor U6875 (N_6875,N_5568,N_3450);
nor U6876 (N_6876,N_5141,N_4644);
or U6877 (N_6877,N_3472,N_3911);
and U6878 (N_6878,N_5003,N_3459);
and U6879 (N_6879,N_5413,N_3185);
and U6880 (N_6880,N_5970,N_3771);
nor U6881 (N_6881,N_3095,N_5368);
and U6882 (N_6882,N_4232,N_5987);
and U6883 (N_6883,N_3393,N_5023);
or U6884 (N_6884,N_4328,N_3129);
nand U6885 (N_6885,N_4389,N_5657);
nor U6886 (N_6886,N_5974,N_5096);
or U6887 (N_6887,N_5872,N_4607);
nand U6888 (N_6888,N_3051,N_5815);
or U6889 (N_6889,N_4727,N_5913);
or U6890 (N_6890,N_5484,N_4722);
nor U6891 (N_6891,N_4976,N_4184);
nand U6892 (N_6892,N_5292,N_4177);
or U6893 (N_6893,N_5526,N_5767);
and U6894 (N_6894,N_4481,N_4192);
nor U6895 (N_6895,N_3581,N_4210);
nand U6896 (N_6896,N_4611,N_3492);
nor U6897 (N_6897,N_4248,N_3921);
and U6898 (N_6898,N_3811,N_3126);
and U6899 (N_6899,N_4170,N_3585);
nor U6900 (N_6900,N_3452,N_4537);
or U6901 (N_6901,N_5916,N_3946);
nand U6902 (N_6902,N_4708,N_4419);
or U6903 (N_6903,N_4595,N_4635);
or U6904 (N_6904,N_5927,N_5539);
nor U6905 (N_6905,N_5662,N_5794);
and U6906 (N_6906,N_4256,N_3453);
nor U6907 (N_6907,N_4564,N_4186);
nor U6908 (N_6908,N_3209,N_4952);
nor U6909 (N_6909,N_3751,N_4991);
or U6910 (N_6910,N_5276,N_4090);
nand U6911 (N_6911,N_4255,N_5395);
or U6912 (N_6912,N_5521,N_3132);
or U6913 (N_6913,N_3652,N_4385);
or U6914 (N_6914,N_3594,N_3762);
or U6915 (N_6915,N_4007,N_4292);
or U6916 (N_6916,N_5810,N_5326);
nor U6917 (N_6917,N_3250,N_5928);
or U6918 (N_6918,N_4439,N_4688);
nor U6919 (N_6919,N_3955,N_5554);
nand U6920 (N_6920,N_5203,N_4059);
and U6921 (N_6921,N_3512,N_5976);
or U6922 (N_6922,N_5986,N_3262);
or U6923 (N_6923,N_4637,N_5026);
nand U6924 (N_6924,N_5696,N_3542);
or U6925 (N_6925,N_4700,N_3952);
nand U6926 (N_6926,N_4265,N_4348);
and U6927 (N_6927,N_3849,N_4703);
nand U6928 (N_6928,N_3267,N_5350);
and U6929 (N_6929,N_4291,N_4020);
and U6930 (N_6930,N_5341,N_4800);
or U6931 (N_6931,N_4748,N_4679);
or U6932 (N_6932,N_5452,N_3867);
and U6933 (N_6933,N_3698,N_5826);
or U6934 (N_6934,N_3822,N_3823);
or U6935 (N_6935,N_4215,N_4418);
nand U6936 (N_6936,N_5726,N_5697);
nand U6937 (N_6937,N_4718,N_5069);
nand U6938 (N_6938,N_4101,N_3044);
and U6939 (N_6939,N_5155,N_4565);
nor U6940 (N_6940,N_5278,N_3708);
nor U6941 (N_6941,N_5320,N_4163);
or U6942 (N_6942,N_5751,N_5494);
or U6943 (N_6943,N_4158,N_3981);
and U6944 (N_6944,N_5899,N_4701);
and U6945 (N_6945,N_3722,N_4967);
or U6946 (N_6946,N_3234,N_3567);
nand U6947 (N_6947,N_4869,N_5835);
nand U6948 (N_6948,N_3336,N_4112);
and U6949 (N_6949,N_3806,N_3394);
and U6950 (N_6950,N_3243,N_4142);
or U6951 (N_6951,N_3531,N_3258);
or U6952 (N_6952,N_5394,N_3706);
and U6953 (N_6953,N_4155,N_4652);
and U6954 (N_6954,N_5414,N_4856);
and U6955 (N_6955,N_3746,N_4651);
nand U6956 (N_6956,N_3043,N_5906);
and U6957 (N_6957,N_5159,N_4355);
nor U6958 (N_6958,N_4045,N_3520);
nor U6959 (N_6959,N_4438,N_3203);
or U6960 (N_6960,N_4975,N_3701);
nor U6961 (N_6961,N_3513,N_5317);
or U6962 (N_6962,N_4113,N_5344);
nand U6963 (N_6963,N_4462,N_5034);
and U6964 (N_6964,N_4840,N_4285);
and U6965 (N_6965,N_5322,N_3518);
nor U6966 (N_6966,N_4378,N_3627);
nor U6967 (N_6967,N_4005,N_5507);
nor U6968 (N_6968,N_5336,N_5240);
and U6969 (N_6969,N_3195,N_4309);
nand U6970 (N_6970,N_5841,N_4552);
and U6971 (N_6971,N_4787,N_3085);
or U6972 (N_6972,N_3078,N_3913);
nand U6973 (N_6973,N_3406,N_5875);
and U6974 (N_6974,N_5191,N_5251);
nor U6975 (N_6975,N_4362,N_5858);
nand U6976 (N_6976,N_5219,N_3147);
nand U6977 (N_6977,N_4835,N_5152);
and U6978 (N_6978,N_4490,N_4613);
or U6979 (N_6979,N_4493,N_3553);
nand U6980 (N_6980,N_5370,N_3380);
nor U6981 (N_6981,N_4488,N_3109);
nor U6982 (N_6982,N_3105,N_5801);
nor U6983 (N_6983,N_3653,N_3808);
nor U6984 (N_6984,N_3062,N_4172);
nand U6985 (N_6985,N_5763,N_3507);
nand U6986 (N_6986,N_5052,N_4250);
nor U6987 (N_6987,N_5105,N_4591);
and U6988 (N_6988,N_5098,N_4548);
or U6989 (N_6989,N_4563,N_5348);
and U6990 (N_6990,N_3623,N_3721);
or U6991 (N_6991,N_5480,N_4788);
or U6992 (N_6992,N_3926,N_5381);
and U6993 (N_6993,N_4179,N_4066);
nand U6994 (N_6994,N_4261,N_3897);
nand U6995 (N_6995,N_3909,N_5605);
or U6996 (N_6996,N_4293,N_3758);
nand U6997 (N_6997,N_4601,N_4524);
nand U6998 (N_6998,N_4408,N_3995);
nor U6999 (N_6999,N_3534,N_3257);
nand U7000 (N_7000,N_5923,N_4207);
nand U7001 (N_7001,N_3107,N_5847);
or U7002 (N_7002,N_3709,N_3504);
and U7003 (N_7003,N_4989,N_4003);
nor U7004 (N_7004,N_4448,N_4807);
nand U7005 (N_7005,N_4646,N_4121);
nor U7006 (N_7006,N_4715,N_3893);
nand U7007 (N_7007,N_4359,N_5512);
nor U7008 (N_7008,N_5624,N_5500);
or U7009 (N_7009,N_4206,N_4533);
and U7010 (N_7010,N_3526,N_3158);
xnor U7011 (N_7011,N_4663,N_5992);
xor U7012 (N_7012,N_3308,N_3246);
and U7013 (N_7013,N_5964,N_4507);
and U7014 (N_7014,N_5759,N_3519);
nand U7015 (N_7015,N_5233,N_5855);
and U7016 (N_7016,N_5871,N_5898);
nand U7017 (N_7017,N_5151,N_4522);
nor U7018 (N_7018,N_5938,N_3645);
nor U7019 (N_7019,N_4426,N_4100);
nor U7020 (N_7020,N_4508,N_3783);
nor U7021 (N_7021,N_3314,N_4275);
or U7022 (N_7022,N_3540,N_4356);
and U7023 (N_7023,N_3899,N_5047);
or U7024 (N_7024,N_4928,N_5360);
and U7025 (N_7025,N_4772,N_4138);
nor U7026 (N_7026,N_4134,N_3826);
and U7027 (N_7027,N_4460,N_3211);
and U7028 (N_7028,N_3924,N_3760);
or U7029 (N_7029,N_3720,N_4083);
or U7030 (N_7030,N_3928,N_4929);
nor U7031 (N_7031,N_4111,N_4397);
nor U7032 (N_7032,N_5547,N_5487);
nand U7033 (N_7033,N_5713,N_3820);
and U7034 (N_7034,N_3361,N_3028);
nand U7035 (N_7035,N_5852,N_3813);
nand U7036 (N_7036,N_5561,N_3776);
and U7037 (N_7037,N_3319,N_5392);
and U7038 (N_7038,N_4973,N_5296);
nor U7039 (N_7039,N_4040,N_3962);
and U7040 (N_7040,N_5099,N_3111);
nand U7041 (N_7041,N_4225,N_5391);
or U7042 (N_7042,N_4457,N_5355);
and U7043 (N_7043,N_3744,N_5182);
nor U7044 (N_7044,N_3878,N_4089);
or U7045 (N_7045,N_3574,N_5272);
and U7046 (N_7046,N_5997,N_3368);
nand U7047 (N_7047,N_3564,N_3588);
nor U7048 (N_7048,N_4226,N_3807);
nor U7049 (N_7049,N_4556,N_4376);
or U7050 (N_7050,N_3057,N_5522);
nand U7051 (N_7051,N_4318,N_3019);
or U7052 (N_7052,N_3468,N_4615);
nand U7053 (N_7053,N_5352,N_4324);
nand U7054 (N_7054,N_3248,N_3383);
and U7055 (N_7055,N_5481,N_4361);
or U7056 (N_7056,N_5692,N_4056);
nor U7057 (N_7057,N_5043,N_4904);
or U7058 (N_7058,N_5649,N_3412);
nor U7059 (N_7059,N_3696,N_3212);
or U7060 (N_7060,N_4746,N_5472);
nor U7061 (N_7061,N_4875,N_4162);
and U7062 (N_7062,N_3730,N_4021);
nand U7063 (N_7063,N_4411,N_5806);
nor U7064 (N_7064,N_4282,N_5412);
nor U7065 (N_7065,N_5583,N_5131);
or U7066 (N_7066,N_5067,N_3614);
or U7067 (N_7067,N_4149,N_4579);
nor U7068 (N_7068,N_3110,N_3919);
and U7069 (N_7069,N_3265,N_3961);
or U7070 (N_7070,N_3884,N_3761);
and U7071 (N_7071,N_5793,N_3681);
nor U7072 (N_7072,N_4427,N_5176);
or U7073 (N_7073,N_4062,N_4302);
or U7074 (N_7074,N_4828,N_5576);
or U7075 (N_7075,N_5464,N_5339);
or U7076 (N_7076,N_4178,N_4336);
and U7077 (N_7077,N_5447,N_3076);
nor U7078 (N_7078,N_4695,N_4360);
nand U7079 (N_7079,N_5846,N_3738);
nand U7080 (N_7080,N_4749,N_4525);
nor U7081 (N_7081,N_3569,N_3227);
nor U7082 (N_7082,N_5599,N_3699);
nand U7083 (N_7083,N_3309,N_3978);
or U7084 (N_7084,N_4758,N_5356);
nand U7085 (N_7085,N_3875,N_5609);
or U7086 (N_7086,N_5265,N_3963);
or U7087 (N_7087,N_4585,N_5424);
and U7088 (N_7088,N_3238,N_3182);
or U7089 (N_7089,N_4377,N_3759);
nand U7090 (N_7090,N_5883,N_3934);
nor U7091 (N_7091,N_5308,N_3781);
or U7092 (N_7092,N_5109,N_3347);
and U7093 (N_7093,N_4590,N_5429);
nor U7094 (N_7094,N_3801,N_3484);
nand U7095 (N_7095,N_5750,N_5932);
and U7096 (N_7096,N_3331,N_4961);
or U7097 (N_7097,N_5533,N_5724);
and U7098 (N_7098,N_5266,N_5586);
or U7099 (N_7099,N_5357,N_3896);
nand U7100 (N_7100,N_4604,N_3455);
nor U7101 (N_7101,N_4078,N_3142);
or U7102 (N_7102,N_5878,N_5907);
nand U7103 (N_7103,N_4229,N_4589);
nand U7104 (N_7104,N_5720,N_3579);
and U7105 (N_7105,N_5223,N_4803);
or U7106 (N_7106,N_5116,N_5467);
or U7107 (N_7107,N_5373,N_5983);
or U7108 (N_7108,N_3584,N_5445);
and U7109 (N_7109,N_5686,N_3888);
nand U7110 (N_7110,N_4165,N_3354);
and U7111 (N_7111,N_3743,N_5865);
or U7112 (N_7112,N_4988,N_3198);
or U7113 (N_7113,N_4039,N_4001);
nand U7114 (N_7114,N_3379,N_3960);
and U7115 (N_7115,N_3487,N_5811);
or U7116 (N_7116,N_5655,N_5699);
nand U7117 (N_7117,N_3138,N_5914);
and U7118 (N_7118,N_4432,N_5197);
or U7119 (N_7119,N_4699,N_3543);
nand U7120 (N_7120,N_3615,N_3013);
nand U7121 (N_7121,N_5019,N_5639);
xnor U7122 (N_7122,N_4057,N_4977);
or U7123 (N_7123,N_3869,N_5629);
nor U7124 (N_7124,N_5733,N_4047);
nand U7125 (N_7125,N_4540,N_3984);
nor U7126 (N_7126,N_5902,N_5115);
nor U7127 (N_7127,N_5104,N_3880);
and U7128 (N_7128,N_3486,N_5269);
or U7129 (N_7129,N_5717,N_4804);
nor U7130 (N_7130,N_3641,N_4196);
nand U7131 (N_7131,N_3726,N_5016);
or U7132 (N_7132,N_4573,N_4181);
and U7133 (N_7133,N_4542,N_5963);
nand U7134 (N_7134,N_5884,N_3938);
nor U7135 (N_7135,N_3020,N_5275);
nand U7136 (N_7136,N_3674,N_5926);
nor U7137 (N_7137,N_5792,N_5366);
and U7138 (N_7138,N_5142,N_5264);
or U7139 (N_7139,N_4363,N_4472);
and U7140 (N_7140,N_5351,N_3204);
nand U7141 (N_7141,N_5289,N_3130);
nor U7142 (N_7142,N_3154,N_3414);
nor U7143 (N_7143,N_4622,N_5497);
or U7144 (N_7144,N_3790,N_4894);
xor U7145 (N_7145,N_3931,N_4531);
nand U7146 (N_7146,N_5315,N_3207);
nand U7147 (N_7147,N_4175,N_3029);
nor U7148 (N_7148,N_5747,N_3865);
xor U7149 (N_7149,N_3325,N_3466);
and U7150 (N_7150,N_4916,N_4406);
nand U7151 (N_7151,N_3602,N_3245);
or U7152 (N_7152,N_4516,N_3732);
and U7153 (N_7153,N_3054,N_4214);
or U7154 (N_7154,N_4190,N_3805);
nor U7155 (N_7155,N_3613,N_5978);
and U7156 (N_7156,N_5723,N_4128);
nor U7157 (N_7157,N_4753,N_4311);
nor U7158 (N_7158,N_4719,N_3342);
or U7159 (N_7159,N_3008,N_3281);
nor U7160 (N_7160,N_3460,N_5458);
or U7161 (N_7161,N_5004,N_5949);
or U7162 (N_7162,N_3866,N_4732);
nor U7163 (N_7163,N_3631,N_4631);
or U7164 (N_7164,N_5643,N_3552);
and U7165 (N_7165,N_3558,N_4633);
and U7166 (N_7166,N_5722,N_4673);
and U7167 (N_7167,N_3037,N_3861);
nor U7168 (N_7168,N_4264,N_3214);
and U7169 (N_7169,N_4019,N_5694);
nor U7170 (N_7170,N_3416,N_4515);
nor U7171 (N_7171,N_5284,N_4289);
nor U7172 (N_7172,N_4509,N_3583);
or U7173 (N_7173,N_5725,N_4820);
nand U7174 (N_7174,N_5020,N_5638);
or U7175 (N_7175,N_3664,N_5761);
nand U7176 (N_7176,N_5385,N_5041);
or U7177 (N_7177,N_3870,N_3470);
or U7178 (N_7178,N_5700,N_5730);
and U7179 (N_7179,N_4501,N_3914);
and U7180 (N_7180,N_5910,N_3677);
or U7181 (N_7181,N_5231,N_4657);
nor U7182 (N_7182,N_4071,N_4879);
nor U7183 (N_7183,N_5551,N_3817);
nor U7184 (N_7184,N_4224,N_3398);
or U7185 (N_7185,N_5184,N_5249);
nor U7186 (N_7186,N_4500,N_3937);
or U7187 (N_7187,N_3648,N_3040);
nor U7188 (N_7188,N_4511,N_3374);
xnor U7189 (N_7189,N_3104,N_5085);
nor U7190 (N_7190,N_4244,N_5967);
and U7191 (N_7191,N_5998,N_4506);
nand U7192 (N_7192,N_4281,N_5056);
nand U7193 (N_7193,N_4778,N_3197);
or U7194 (N_7194,N_3829,N_5072);
or U7195 (N_7195,N_4137,N_5783);
nor U7196 (N_7196,N_5457,N_4747);
nor U7197 (N_7197,N_5466,N_3704);
or U7198 (N_7198,N_3780,N_4921);
xor U7199 (N_7199,N_4888,N_5908);
or U7200 (N_7200,N_5432,N_5499);
nand U7201 (N_7201,N_5418,N_4428);
or U7202 (N_7202,N_5510,N_3369);
or U7203 (N_7203,N_3634,N_4185);
or U7204 (N_7204,N_5380,N_4970);
nand U7205 (N_7205,N_3818,N_5166);
and U7206 (N_7206,N_5125,N_5860);
or U7207 (N_7207,N_5493,N_5603);
and U7208 (N_7208,N_4449,N_4160);
xor U7209 (N_7209,N_5062,N_4691);
and U7210 (N_7210,N_5369,N_3181);
or U7211 (N_7211,N_3367,N_4271);
nor U7212 (N_7212,N_4672,N_5222);
nor U7213 (N_7213,N_3741,N_3836);
nand U7214 (N_7214,N_4204,N_4554);
or U7215 (N_7215,N_4603,N_4300);
nor U7216 (N_7216,N_4717,N_5757);
or U7217 (N_7217,N_3786,N_3988);
and U7218 (N_7218,N_4279,N_4347);
nor U7219 (N_7219,N_4041,N_3672);
nor U7220 (N_7220,N_5580,N_4227);
nor U7221 (N_7221,N_3196,N_5214);
nand U7222 (N_7222,N_3275,N_3304);
and U7223 (N_7223,N_3991,N_3224);
or U7224 (N_7224,N_3624,N_3344);
nor U7225 (N_7225,N_4310,N_3060);
or U7226 (N_7226,N_4599,N_3409);
nor U7227 (N_7227,N_5354,N_4358);
and U7228 (N_7228,N_3640,N_4941);
and U7229 (N_7229,N_3948,N_4087);
nor U7230 (N_7230,N_5574,N_3676);
and U7231 (N_7231,N_5782,N_4304);
and U7232 (N_7232,N_4825,N_4801);
nand U7233 (N_7233,N_3784,N_5375);
or U7234 (N_7234,N_3156,N_5640);
and U7235 (N_7235,N_3089,N_4969);
nor U7236 (N_7236,N_4729,N_4399);
nand U7237 (N_7237,N_4714,N_3220);
nand U7238 (N_7238,N_4122,N_3779);
nand U7239 (N_7239,N_3493,N_3134);
or U7240 (N_7240,N_5444,N_3649);
or U7241 (N_7241,N_3993,N_4094);
and U7242 (N_7242,N_3599,N_4064);
nand U7243 (N_7243,N_5064,N_4297);
or U7244 (N_7244,N_5995,N_3175);
or U7245 (N_7245,N_5420,N_5235);
nand U7246 (N_7246,N_3168,N_4583);
or U7247 (N_7247,N_5673,N_3006);
nand U7248 (N_7248,N_4649,N_5879);
and U7249 (N_7249,N_3570,N_5827);
nor U7250 (N_7250,N_4187,N_4766);
or U7251 (N_7251,N_5621,N_3748);
nand U7252 (N_7252,N_3117,N_4983);
nand U7253 (N_7253,N_5647,N_3352);
nand U7254 (N_7254,N_5073,N_3324);
and U7255 (N_7255,N_4997,N_4409);
and U7256 (N_7256,N_5258,N_3853);
nor U7257 (N_7257,N_5403,N_4802);
xor U7258 (N_7258,N_4118,N_4963);
and U7259 (N_7259,N_5008,N_4116);
and U7260 (N_7260,N_5896,N_3315);
nand U7261 (N_7261,N_4407,N_4343);
nor U7262 (N_7262,N_5600,N_4934);
or U7263 (N_7263,N_5977,N_4156);
nor U7264 (N_7264,N_5851,N_4666);
nor U7265 (N_7265,N_5082,N_5569);
or U7266 (N_7266,N_3422,N_5100);
nand U7267 (N_7267,N_4518,N_3055);
and U7268 (N_7268,N_5931,N_4091);
and U7269 (N_7269,N_5814,N_4784);
nand U7270 (N_7270,N_5079,N_3167);
and U7271 (N_7271,N_4295,N_4621);
nor U7272 (N_7272,N_5361,N_4043);
and U7273 (N_7273,N_3268,N_5139);
and U7274 (N_7274,N_5386,N_5434);
or U7275 (N_7275,N_5527,N_3030);
and U7276 (N_7276,N_3143,N_5589);
nand U7277 (N_7277,N_5146,N_5304);
nor U7278 (N_7278,N_3657,N_4764);
or U7279 (N_7279,N_3413,N_3753);
nor U7280 (N_7280,N_4478,N_5711);
nor U7281 (N_7281,N_5962,N_3179);
or U7282 (N_7282,N_5290,N_5575);
or U7283 (N_7283,N_4641,N_3483);
nand U7284 (N_7284,N_3718,N_3886);
or U7285 (N_7285,N_3539,N_4813);
or U7286 (N_7286,N_5359,N_5195);
or U7287 (N_7287,N_3180,N_4920);
nor U7288 (N_7288,N_5552,N_4946);
nand U7289 (N_7289,N_3226,N_4161);
or U7290 (N_7290,N_3620,N_5132);
nor U7291 (N_7291,N_5201,N_3219);
nor U7292 (N_7292,N_3079,N_5332);
nand U7293 (N_7293,N_4238,N_3321);
nor U7294 (N_7294,N_4323,N_3306);
nor U7295 (N_7295,N_5542,N_5795);
nand U7296 (N_7296,N_3046,N_4371);
and U7297 (N_7297,N_3225,N_3457);
nand U7298 (N_7298,N_5083,N_4384);
nand U7299 (N_7299,N_4013,N_3702);
or U7300 (N_7300,N_5440,N_4536);
nor U7301 (N_7301,N_3679,N_5059);
nor U7302 (N_7302,N_5252,N_3298);
and U7303 (N_7303,N_4280,N_5857);
nand U7304 (N_7304,N_3289,N_3000);
or U7305 (N_7305,N_5950,N_5158);
xor U7306 (N_7306,N_5968,N_3576);
and U7307 (N_7307,N_5136,N_3716);
nand U7308 (N_7308,N_5952,N_4284);
and U7309 (N_7309,N_5086,N_4277);
and U7310 (N_7310,N_5470,N_3912);
nor U7311 (N_7311,N_5270,N_4420);
nor U7312 (N_7312,N_3697,N_3933);
nor U7313 (N_7313,N_4568,N_5460);
nand U7314 (N_7314,N_3906,N_5834);
nor U7315 (N_7315,N_4683,N_5077);
nor U7316 (N_7316,N_3066,N_4431);
and U7317 (N_7317,N_5805,N_3050);
and U7318 (N_7318,N_3448,N_3462);
and U7319 (N_7319,N_3589,N_4220);
and U7320 (N_7320,N_4503,N_3277);
or U7321 (N_7321,N_3115,N_4741);
and U7322 (N_7322,N_3183,N_3593);
nor U7323 (N_7323,N_3339,N_5437);
nand U7324 (N_7324,N_3465,N_3122);
nor U7325 (N_7325,N_3691,N_4567);
and U7326 (N_7326,N_5786,N_5728);
and U7327 (N_7327,N_5566,N_5225);
and U7328 (N_7328,N_4867,N_4352);
or U7329 (N_7329,N_3603,N_3847);
or U7330 (N_7330,N_3210,N_3064);
nand U7331 (N_7331,N_4200,N_4370);
nor U7332 (N_7332,N_4219,N_3885);
nor U7333 (N_7333,N_3011,N_5164);
nand U7334 (N_7334,N_4994,N_4874);
nand U7335 (N_7335,N_4907,N_5900);
and U7336 (N_7336,N_5636,N_4373);
or U7337 (N_7337,N_3890,N_4696);
nor U7338 (N_7338,N_3966,N_3793);
nand U7339 (N_7339,N_5256,N_5619);
nor U7340 (N_7340,N_5889,N_5450);
nor U7341 (N_7341,N_5262,N_4889);
nor U7342 (N_7342,N_4926,N_5813);
nor U7343 (N_7343,N_4893,N_4964);
or U7344 (N_7344,N_3713,N_3667);
nor U7345 (N_7345,N_3626,N_5531);
and U7346 (N_7346,N_3501,N_4423);
nor U7347 (N_7347,N_5114,N_5149);
and U7348 (N_7348,N_3081,N_5780);
nand U7349 (N_7349,N_5076,N_4096);
nor U7350 (N_7350,N_4417,N_3678);
and U7351 (N_7351,N_4191,N_5769);
and U7352 (N_7352,N_4955,N_4939);
and U7353 (N_7353,N_4237,N_3999);
and U7354 (N_7354,N_5956,N_3026);
and U7355 (N_7355,N_4981,N_3629);
nor U7356 (N_7356,N_5044,N_4450);
and U7357 (N_7357,N_3096,N_4830);
nand U7358 (N_7358,N_4723,N_4819);
nor U7359 (N_7359,N_4682,N_4865);
and U7360 (N_7360,N_5455,N_4636);
nand U7361 (N_7361,N_3477,N_4512);
nor U7362 (N_7362,N_3461,N_5371);
nor U7363 (N_7363,N_4600,N_3957);
and U7364 (N_7364,N_5297,N_5364);
or U7365 (N_7365,N_4260,N_5471);
and U7366 (N_7366,N_5294,N_5703);
nor U7367 (N_7367,N_4093,N_4736);
and U7368 (N_7368,N_5295,N_4095);
nand U7369 (N_7369,N_5562,N_5870);
nor U7370 (N_7370,N_5283,N_5120);
nand U7371 (N_7371,N_3408,N_4240);
or U7372 (N_7372,N_5612,N_4982);
and U7373 (N_7373,N_5856,N_5384);
nand U7374 (N_7374,N_3328,N_3108);
nor U7375 (N_7375,N_4489,N_5646);
xnor U7376 (N_7376,N_3601,N_3080);
nor U7377 (N_7377,N_5771,N_5622);
or U7378 (N_7378,N_3825,N_4949);
nand U7379 (N_7379,N_4276,N_4474);
or U7380 (N_7380,N_5866,N_3528);
nand U7381 (N_7381,N_4529,N_5800);
nand U7382 (N_7382,N_5874,N_3998);
xor U7383 (N_7383,N_3445,N_3502);
or U7384 (N_7384,N_5617,N_4245);
nor U7385 (N_7385,N_5626,N_4372);
nor U7386 (N_7386,N_3951,N_3148);
nor U7387 (N_7387,N_3437,N_4810);
nor U7388 (N_7388,N_4485,N_3475);
nor U7389 (N_7389,N_4897,N_5358);
nand U7390 (N_7390,N_4750,N_5254);
and U7391 (N_7391,N_5113,N_3120);
xor U7392 (N_7392,N_4805,N_3119);
xor U7393 (N_7393,N_3443,N_4720);
and U7394 (N_7394,N_5627,N_5228);
nor U7395 (N_7395,N_4956,N_5436);
nor U7396 (N_7396,N_4987,N_4379);
and U7397 (N_7397,N_5707,N_3794);
nand U7398 (N_7398,N_4712,N_3338);
or U7399 (N_7399,N_5625,N_4850);
nand U7400 (N_7400,N_4658,N_3763);
nand U7401 (N_7401,N_5063,N_4721);
or U7402 (N_7402,N_3451,N_3116);
and U7403 (N_7403,N_5996,N_5863);
nand U7404 (N_7404,N_3740,N_5675);
nand U7405 (N_7405,N_4125,N_5822);
or U7406 (N_7406,N_5905,N_3135);
nand U7407 (N_7407,N_5084,N_4743);
nand U7408 (N_7408,N_5930,N_5781);
nand U7409 (N_7409,N_3915,N_4008);
nand U7410 (N_7410,N_4391,N_5869);
and U7411 (N_7411,N_4412,N_3194);
nor U7412 (N_7412,N_5895,N_5664);
nand U7413 (N_7413,N_3632,N_3157);
and U7414 (N_7414,N_4821,N_4392);
nor U7415 (N_7415,N_3608,N_5478);
nor U7416 (N_7416,N_4954,N_4693);
nand U7417 (N_7417,N_3186,N_3480);
or U7418 (N_7418,N_3033,N_4037);
or U7419 (N_7419,N_5119,N_4612);
and U7420 (N_7420,N_4957,N_5924);
or U7421 (N_7421,N_4876,N_5660);
or U7422 (N_7422,N_3065,N_3517);
or U7423 (N_7423,N_3058,N_3329);
or U7424 (N_7424,N_3396,N_3073);
or U7425 (N_7425,N_4562,N_3901);
nor U7426 (N_7426,N_4665,N_5604);
nor U7427 (N_7427,N_5123,N_3850);
nor U7428 (N_7428,N_4966,N_4960);
or U7429 (N_7429,N_4664,N_4414);
or U7430 (N_7430,N_3247,N_4587);
xor U7431 (N_7431,N_5261,N_4638);
and U7432 (N_7432,N_4915,N_5241);
nand U7433 (N_7433,N_5845,N_4126);
and U7434 (N_7434,N_4319,N_4625);
nand U7435 (N_7435,N_3846,N_4147);
or U7436 (N_7436,N_3923,N_4945);
or U7437 (N_7437,N_5693,N_5028);
nor U7438 (N_7438,N_5232,N_3199);
or U7439 (N_7439,N_4069,N_5423);
nand U7440 (N_7440,N_3300,N_3843);
nand U7441 (N_7441,N_3365,N_5544);
nor U7442 (N_7442,N_3091,N_3405);
and U7443 (N_7443,N_4029,N_4849);
and U7444 (N_7444,N_5803,N_3683);
nor U7445 (N_7445,N_4085,N_5287);
or U7446 (N_7446,N_5981,N_5778);
or U7447 (N_7447,N_5842,N_4269);
and U7448 (N_7448,N_4081,N_3071);
or U7449 (N_7449,N_4383,N_4735);
nand U7450 (N_7450,N_5363,N_4327);
and U7451 (N_7451,N_4139,N_5524);
nor U7452 (N_7452,N_5731,N_5271);
nor U7453 (N_7453,N_4656,N_5147);
nand U7454 (N_7454,N_5002,N_3251);
nor U7455 (N_7455,N_5538,N_4979);
and U7456 (N_7456,N_4950,N_3530);
or U7457 (N_7457,N_4771,N_4999);
and U7458 (N_7458,N_3729,N_4671);
or U7459 (N_7459,N_3804,N_4382);
and U7460 (N_7460,N_4451,N_4557);
nand U7461 (N_7461,N_5259,N_5565);
nor U7462 (N_7462,N_5068,N_5070);
and U7463 (N_7463,N_4102,N_4882);
or U7464 (N_7464,N_3390,N_5376);
and U7465 (N_7465,N_3545,N_4014);
and U7466 (N_7466,N_4730,N_3420);
nand U7467 (N_7467,N_3757,N_5873);
nor U7468 (N_7468,N_3330,N_4824);
nand U7469 (N_7469,N_5613,N_4239);
nand U7470 (N_7470,N_3035,N_5774);
nand U7471 (N_7471,N_3473,N_4011);
and U7472 (N_7472,N_4119,N_3474);
or U7473 (N_7473,N_5459,N_3685);
or U7474 (N_7474,N_5867,N_4614);
and U7475 (N_7475,N_3889,N_3959);
and U7476 (N_7476,N_3162,N_3562);
and U7477 (N_7477,N_4517,N_3868);
nor U7478 (N_7478,N_4060,N_3669);
nand U7479 (N_7479,N_5492,N_4871);
nor U7480 (N_7480,N_3193,N_3812);
and U7481 (N_7481,N_4685,N_4551);
nand U7482 (N_7482,N_5593,N_5333);
and U7483 (N_7483,N_4620,N_3173);
and U7484 (N_7484,N_5702,N_5216);
and U7485 (N_7485,N_3141,N_4676);
nand U7486 (N_7486,N_5051,N_3733);
nor U7487 (N_7487,N_5517,N_3436);
and U7488 (N_7488,N_5399,N_3357);
or U7489 (N_7489,N_5990,N_5217);
and U7490 (N_7490,N_5469,N_3145);
and U7491 (N_7491,N_4626,N_4217);
nor U7492 (N_7492,N_4398,N_5092);
and U7493 (N_7493,N_3291,N_5268);
nor U7494 (N_7494,N_5746,N_3922);
and U7495 (N_7495,N_5404,N_3335);
nor U7496 (N_7496,N_3184,N_4278);
and U7497 (N_7497,N_5138,N_3326);
or U7498 (N_7498,N_5053,N_5167);
and U7499 (N_7499,N_4286,N_3097);
nor U7500 (N_7500,N_5203,N_3418);
and U7501 (N_7501,N_4665,N_4080);
and U7502 (N_7502,N_5944,N_4070);
or U7503 (N_7503,N_4353,N_3764);
nor U7504 (N_7504,N_3257,N_3549);
nand U7505 (N_7505,N_5657,N_5240);
nand U7506 (N_7506,N_4422,N_3705);
nand U7507 (N_7507,N_5996,N_3754);
nand U7508 (N_7508,N_3782,N_5925);
and U7509 (N_7509,N_5333,N_4280);
nand U7510 (N_7510,N_3102,N_4964);
and U7511 (N_7511,N_5621,N_4089);
nor U7512 (N_7512,N_4534,N_4028);
nand U7513 (N_7513,N_4525,N_5194);
nor U7514 (N_7514,N_4693,N_5805);
and U7515 (N_7515,N_3464,N_3240);
nand U7516 (N_7516,N_4023,N_5959);
and U7517 (N_7517,N_4600,N_3102);
nand U7518 (N_7518,N_5708,N_4159);
nand U7519 (N_7519,N_3083,N_5911);
nor U7520 (N_7520,N_5885,N_5535);
nor U7521 (N_7521,N_4845,N_5874);
nand U7522 (N_7522,N_4923,N_3766);
xor U7523 (N_7523,N_3534,N_5751);
or U7524 (N_7524,N_4047,N_4480);
and U7525 (N_7525,N_5759,N_3542);
and U7526 (N_7526,N_4311,N_3715);
or U7527 (N_7527,N_4800,N_3480);
or U7528 (N_7528,N_3746,N_3486);
and U7529 (N_7529,N_5433,N_4544);
nor U7530 (N_7530,N_5847,N_3261);
nand U7531 (N_7531,N_5077,N_3786);
or U7532 (N_7532,N_5395,N_3864);
nand U7533 (N_7533,N_4865,N_4846);
or U7534 (N_7534,N_5255,N_4076);
nor U7535 (N_7535,N_4186,N_4746);
nand U7536 (N_7536,N_4840,N_4973);
nor U7537 (N_7537,N_3487,N_4725);
nor U7538 (N_7538,N_4665,N_4198);
nor U7539 (N_7539,N_4850,N_5052);
nand U7540 (N_7540,N_3214,N_5620);
nor U7541 (N_7541,N_5640,N_3361);
and U7542 (N_7542,N_5709,N_3648);
or U7543 (N_7543,N_3602,N_3333);
nand U7544 (N_7544,N_4053,N_3478);
or U7545 (N_7545,N_3636,N_5038);
nand U7546 (N_7546,N_5237,N_4513);
and U7547 (N_7547,N_3074,N_4383);
or U7548 (N_7548,N_4691,N_3491);
nor U7549 (N_7549,N_3901,N_5167);
or U7550 (N_7550,N_3389,N_4340);
nor U7551 (N_7551,N_3015,N_5263);
nor U7552 (N_7552,N_5674,N_3242);
and U7553 (N_7553,N_4193,N_3985);
or U7554 (N_7554,N_5434,N_3161);
or U7555 (N_7555,N_3930,N_4187);
xnor U7556 (N_7556,N_5027,N_3042);
nand U7557 (N_7557,N_4191,N_3570);
or U7558 (N_7558,N_4219,N_4122);
nand U7559 (N_7559,N_4273,N_5041);
or U7560 (N_7560,N_3806,N_3161);
and U7561 (N_7561,N_3701,N_3563);
nand U7562 (N_7562,N_4322,N_3180);
nor U7563 (N_7563,N_3036,N_5431);
or U7564 (N_7564,N_3328,N_3780);
nand U7565 (N_7565,N_5538,N_5414);
nand U7566 (N_7566,N_5675,N_3211);
and U7567 (N_7567,N_5876,N_5368);
xor U7568 (N_7568,N_4823,N_5663);
nor U7569 (N_7569,N_5210,N_4082);
xnor U7570 (N_7570,N_5490,N_5306);
or U7571 (N_7571,N_4757,N_5217);
nor U7572 (N_7572,N_3052,N_4405);
or U7573 (N_7573,N_3068,N_4270);
and U7574 (N_7574,N_5886,N_3212);
nor U7575 (N_7575,N_4975,N_3798);
nand U7576 (N_7576,N_5867,N_5822);
nand U7577 (N_7577,N_3858,N_3714);
and U7578 (N_7578,N_3700,N_5297);
and U7579 (N_7579,N_3576,N_4705);
nor U7580 (N_7580,N_4942,N_5208);
and U7581 (N_7581,N_4127,N_4547);
nand U7582 (N_7582,N_3081,N_3793);
nand U7583 (N_7583,N_3009,N_4561);
nor U7584 (N_7584,N_3272,N_3691);
nand U7585 (N_7585,N_3124,N_5128);
nor U7586 (N_7586,N_4571,N_4224);
and U7587 (N_7587,N_4284,N_5143);
or U7588 (N_7588,N_5855,N_4183);
or U7589 (N_7589,N_4344,N_3802);
or U7590 (N_7590,N_5539,N_5633);
or U7591 (N_7591,N_5305,N_3265);
nand U7592 (N_7592,N_4352,N_4380);
nor U7593 (N_7593,N_4686,N_3925);
and U7594 (N_7594,N_5575,N_5880);
nor U7595 (N_7595,N_5961,N_5850);
nor U7596 (N_7596,N_5093,N_3584);
nand U7597 (N_7597,N_4460,N_3135);
xnor U7598 (N_7598,N_5315,N_4587);
nand U7599 (N_7599,N_4637,N_5451);
nand U7600 (N_7600,N_4066,N_4711);
or U7601 (N_7601,N_4140,N_3153);
nand U7602 (N_7602,N_4038,N_3320);
nor U7603 (N_7603,N_3331,N_3925);
and U7604 (N_7604,N_5785,N_5475);
and U7605 (N_7605,N_3219,N_5108);
and U7606 (N_7606,N_4420,N_3341);
and U7607 (N_7607,N_4037,N_4467);
nand U7608 (N_7608,N_5456,N_5998);
and U7609 (N_7609,N_4719,N_5503);
nor U7610 (N_7610,N_5114,N_3950);
and U7611 (N_7611,N_3202,N_3033);
nand U7612 (N_7612,N_5597,N_5977);
or U7613 (N_7613,N_3364,N_3427);
nor U7614 (N_7614,N_4279,N_5827);
or U7615 (N_7615,N_4880,N_5030);
nor U7616 (N_7616,N_5797,N_5482);
and U7617 (N_7617,N_5967,N_5048);
and U7618 (N_7618,N_3117,N_3230);
or U7619 (N_7619,N_4373,N_5981);
and U7620 (N_7620,N_5508,N_4854);
nand U7621 (N_7621,N_4775,N_3523);
or U7622 (N_7622,N_4863,N_5737);
or U7623 (N_7623,N_3590,N_5594);
or U7624 (N_7624,N_4692,N_5529);
nand U7625 (N_7625,N_5927,N_3112);
nand U7626 (N_7626,N_4517,N_5375);
nand U7627 (N_7627,N_3947,N_4781);
nor U7628 (N_7628,N_5003,N_4124);
nor U7629 (N_7629,N_5339,N_5427);
or U7630 (N_7630,N_4217,N_5079);
or U7631 (N_7631,N_3329,N_3826);
or U7632 (N_7632,N_4601,N_3354);
and U7633 (N_7633,N_3831,N_4301);
and U7634 (N_7634,N_5762,N_3929);
and U7635 (N_7635,N_5444,N_3839);
nand U7636 (N_7636,N_5029,N_3404);
nor U7637 (N_7637,N_4440,N_4989);
nor U7638 (N_7638,N_3514,N_4112);
nor U7639 (N_7639,N_3184,N_5713);
and U7640 (N_7640,N_4018,N_4729);
nor U7641 (N_7641,N_3453,N_3458);
nand U7642 (N_7642,N_5332,N_5385);
and U7643 (N_7643,N_5228,N_3015);
or U7644 (N_7644,N_5039,N_4433);
and U7645 (N_7645,N_5786,N_4114);
or U7646 (N_7646,N_3556,N_5750);
nor U7647 (N_7647,N_3882,N_3183);
or U7648 (N_7648,N_5073,N_4283);
nor U7649 (N_7649,N_4002,N_3119);
nand U7650 (N_7650,N_3626,N_3887);
nor U7651 (N_7651,N_4607,N_4537);
or U7652 (N_7652,N_4805,N_3840);
nor U7653 (N_7653,N_4280,N_5328);
or U7654 (N_7654,N_3928,N_3579);
nor U7655 (N_7655,N_5615,N_4324);
or U7656 (N_7656,N_4181,N_3624);
nor U7657 (N_7657,N_4014,N_5548);
nand U7658 (N_7658,N_5407,N_4023);
or U7659 (N_7659,N_3644,N_4431);
nand U7660 (N_7660,N_4809,N_4401);
nand U7661 (N_7661,N_4804,N_4132);
and U7662 (N_7662,N_3824,N_4045);
nor U7663 (N_7663,N_3277,N_3690);
nor U7664 (N_7664,N_4506,N_3890);
nand U7665 (N_7665,N_4141,N_4739);
nand U7666 (N_7666,N_5909,N_3761);
nand U7667 (N_7667,N_5651,N_3853);
nor U7668 (N_7668,N_4213,N_5171);
and U7669 (N_7669,N_5385,N_5583);
nand U7670 (N_7670,N_5208,N_3768);
and U7671 (N_7671,N_4818,N_5210);
nand U7672 (N_7672,N_4928,N_4398);
or U7673 (N_7673,N_4170,N_5254);
and U7674 (N_7674,N_5016,N_4133);
nand U7675 (N_7675,N_5070,N_3571);
nand U7676 (N_7676,N_5115,N_5717);
nand U7677 (N_7677,N_4514,N_3725);
or U7678 (N_7678,N_3271,N_3872);
or U7679 (N_7679,N_4124,N_4921);
nor U7680 (N_7680,N_4116,N_4864);
nor U7681 (N_7681,N_4693,N_4739);
nand U7682 (N_7682,N_5270,N_3186);
nor U7683 (N_7683,N_4212,N_3478);
and U7684 (N_7684,N_3063,N_3347);
nor U7685 (N_7685,N_3098,N_3925);
nor U7686 (N_7686,N_4774,N_3148);
and U7687 (N_7687,N_5806,N_4474);
or U7688 (N_7688,N_3385,N_3310);
nand U7689 (N_7689,N_4815,N_4153);
nand U7690 (N_7690,N_3516,N_4547);
and U7691 (N_7691,N_4412,N_4047);
or U7692 (N_7692,N_3149,N_3820);
or U7693 (N_7693,N_4442,N_4837);
nand U7694 (N_7694,N_5682,N_3893);
or U7695 (N_7695,N_3475,N_4760);
or U7696 (N_7696,N_5377,N_5737);
and U7697 (N_7697,N_3495,N_5512);
nand U7698 (N_7698,N_5967,N_4607);
nor U7699 (N_7699,N_3261,N_4662);
nor U7700 (N_7700,N_3898,N_3918);
nor U7701 (N_7701,N_5189,N_3974);
and U7702 (N_7702,N_5761,N_5837);
nand U7703 (N_7703,N_4656,N_3376);
nand U7704 (N_7704,N_3985,N_5593);
or U7705 (N_7705,N_4242,N_3456);
nand U7706 (N_7706,N_4212,N_5822);
nand U7707 (N_7707,N_3795,N_3544);
nor U7708 (N_7708,N_4094,N_5762);
or U7709 (N_7709,N_4943,N_4938);
nor U7710 (N_7710,N_5143,N_3877);
and U7711 (N_7711,N_4277,N_3345);
nor U7712 (N_7712,N_3297,N_4685);
nor U7713 (N_7713,N_5944,N_5938);
or U7714 (N_7714,N_4731,N_4903);
nand U7715 (N_7715,N_4258,N_5583);
nor U7716 (N_7716,N_5242,N_4147);
and U7717 (N_7717,N_5424,N_4535);
and U7718 (N_7718,N_5471,N_3818);
and U7719 (N_7719,N_3699,N_3886);
nor U7720 (N_7720,N_4387,N_3247);
or U7721 (N_7721,N_3466,N_3515);
xnor U7722 (N_7722,N_4290,N_3303);
or U7723 (N_7723,N_4127,N_4147);
xnor U7724 (N_7724,N_4814,N_5283);
nor U7725 (N_7725,N_4546,N_5766);
nand U7726 (N_7726,N_4843,N_3249);
nor U7727 (N_7727,N_3960,N_4058);
nor U7728 (N_7728,N_3295,N_3548);
and U7729 (N_7729,N_4625,N_3836);
or U7730 (N_7730,N_3555,N_3329);
and U7731 (N_7731,N_5548,N_5245);
nand U7732 (N_7732,N_5085,N_3253);
and U7733 (N_7733,N_3524,N_4037);
and U7734 (N_7734,N_5658,N_3374);
nor U7735 (N_7735,N_3291,N_4667);
or U7736 (N_7736,N_4835,N_3228);
or U7737 (N_7737,N_5426,N_5585);
or U7738 (N_7738,N_5629,N_4914);
and U7739 (N_7739,N_5903,N_3668);
nand U7740 (N_7740,N_4623,N_4522);
nand U7741 (N_7741,N_5656,N_4552);
nor U7742 (N_7742,N_5338,N_5744);
or U7743 (N_7743,N_5592,N_3647);
nand U7744 (N_7744,N_4995,N_3275);
and U7745 (N_7745,N_5292,N_3654);
and U7746 (N_7746,N_3395,N_4697);
nand U7747 (N_7747,N_4752,N_5301);
nand U7748 (N_7748,N_5504,N_5623);
and U7749 (N_7749,N_3543,N_4942);
nand U7750 (N_7750,N_3796,N_5685);
and U7751 (N_7751,N_5575,N_4487);
or U7752 (N_7752,N_3222,N_3549);
nand U7753 (N_7753,N_3213,N_4544);
or U7754 (N_7754,N_3446,N_3586);
or U7755 (N_7755,N_5924,N_3667);
nand U7756 (N_7756,N_3206,N_4106);
nor U7757 (N_7757,N_5924,N_3213);
and U7758 (N_7758,N_5925,N_4646);
nand U7759 (N_7759,N_5131,N_4301);
or U7760 (N_7760,N_3595,N_3940);
nor U7761 (N_7761,N_4294,N_4027);
or U7762 (N_7762,N_4450,N_3839);
nand U7763 (N_7763,N_4985,N_5568);
or U7764 (N_7764,N_5783,N_3769);
nand U7765 (N_7765,N_3005,N_5274);
or U7766 (N_7766,N_4086,N_5550);
and U7767 (N_7767,N_3909,N_5125);
and U7768 (N_7768,N_4370,N_4978);
nor U7769 (N_7769,N_4521,N_3992);
nand U7770 (N_7770,N_5459,N_3992);
or U7771 (N_7771,N_4473,N_5995);
nor U7772 (N_7772,N_5280,N_5444);
and U7773 (N_7773,N_5852,N_3200);
nor U7774 (N_7774,N_3019,N_5461);
nor U7775 (N_7775,N_5810,N_4023);
and U7776 (N_7776,N_4323,N_3810);
or U7777 (N_7777,N_5175,N_5833);
or U7778 (N_7778,N_3145,N_3532);
and U7779 (N_7779,N_4985,N_3036);
nand U7780 (N_7780,N_3864,N_5842);
nand U7781 (N_7781,N_4206,N_3961);
nor U7782 (N_7782,N_4327,N_4536);
nand U7783 (N_7783,N_5993,N_4271);
nand U7784 (N_7784,N_4302,N_5946);
nand U7785 (N_7785,N_3795,N_3438);
nor U7786 (N_7786,N_3122,N_4882);
or U7787 (N_7787,N_4982,N_5556);
nor U7788 (N_7788,N_5842,N_3929);
or U7789 (N_7789,N_3741,N_4426);
or U7790 (N_7790,N_5908,N_3575);
and U7791 (N_7791,N_5382,N_5902);
and U7792 (N_7792,N_5852,N_5192);
xnor U7793 (N_7793,N_5841,N_5435);
and U7794 (N_7794,N_3618,N_3284);
or U7795 (N_7795,N_4655,N_3170);
nor U7796 (N_7796,N_3360,N_5396);
and U7797 (N_7797,N_3405,N_5540);
or U7798 (N_7798,N_4059,N_4662);
nand U7799 (N_7799,N_5386,N_3791);
nand U7800 (N_7800,N_3040,N_3415);
and U7801 (N_7801,N_3008,N_5480);
nor U7802 (N_7802,N_5483,N_5688);
nand U7803 (N_7803,N_4300,N_3951);
nor U7804 (N_7804,N_3843,N_3820);
nand U7805 (N_7805,N_5453,N_4703);
and U7806 (N_7806,N_3406,N_3202);
or U7807 (N_7807,N_3827,N_3223);
nor U7808 (N_7808,N_4995,N_4858);
and U7809 (N_7809,N_3785,N_4245);
nor U7810 (N_7810,N_3029,N_4874);
nor U7811 (N_7811,N_4157,N_3775);
nor U7812 (N_7812,N_3761,N_5416);
and U7813 (N_7813,N_4629,N_5987);
or U7814 (N_7814,N_5767,N_3502);
nor U7815 (N_7815,N_3376,N_3161);
or U7816 (N_7816,N_4530,N_5499);
nand U7817 (N_7817,N_3005,N_5685);
or U7818 (N_7818,N_3224,N_3358);
nand U7819 (N_7819,N_4396,N_4378);
nand U7820 (N_7820,N_4001,N_3181);
and U7821 (N_7821,N_5091,N_4803);
or U7822 (N_7822,N_4139,N_4228);
nand U7823 (N_7823,N_5932,N_5702);
or U7824 (N_7824,N_4788,N_3279);
nor U7825 (N_7825,N_4490,N_4304);
or U7826 (N_7826,N_3925,N_3179);
nand U7827 (N_7827,N_5917,N_5157);
or U7828 (N_7828,N_5985,N_4109);
nor U7829 (N_7829,N_4008,N_5536);
nand U7830 (N_7830,N_5304,N_5801);
nand U7831 (N_7831,N_5387,N_4238);
nand U7832 (N_7832,N_4143,N_5453);
nand U7833 (N_7833,N_4563,N_3852);
or U7834 (N_7834,N_3391,N_3517);
nor U7835 (N_7835,N_4037,N_5293);
nor U7836 (N_7836,N_3061,N_3198);
and U7837 (N_7837,N_3157,N_3864);
nand U7838 (N_7838,N_5500,N_3903);
and U7839 (N_7839,N_4292,N_3882);
nand U7840 (N_7840,N_4247,N_5704);
or U7841 (N_7841,N_4427,N_5798);
nor U7842 (N_7842,N_5884,N_5485);
nor U7843 (N_7843,N_4423,N_5978);
nand U7844 (N_7844,N_4796,N_3666);
nor U7845 (N_7845,N_4566,N_3147);
nor U7846 (N_7846,N_4612,N_3852);
or U7847 (N_7847,N_4623,N_4552);
and U7848 (N_7848,N_5186,N_3719);
and U7849 (N_7849,N_4341,N_4336);
nor U7850 (N_7850,N_4773,N_5255);
or U7851 (N_7851,N_5428,N_3831);
nand U7852 (N_7852,N_5986,N_4370);
and U7853 (N_7853,N_5134,N_4272);
nand U7854 (N_7854,N_5225,N_4313);
and U7855 (N_7855,N_4222,N_3189);
or U7856 (N_7856,N_3256,N_3760);
nor U7857 (N_7857,N_5572,N_5643);
nand U7858 (N_7858,N_5983,N_4498);
nand U7859 (N_7859,N_3684,N_3189);
and U7860 (N_7860,N_4234,N_5050);
and U7861 (N_7861,N_5013,N_5282);
or U7862 (N_7862,N_4510,N_3307);
nor U7863 (N_7863,N_4851,N_4529);
nor U7864 (N_7864,N_3826,N_3125);
and U7865 (N_7865,N_4086,N_3357);
nand U7866 (N_7866,N_3426,N_3538);
nor U7867 (N_7867,N_3868,N_5689);
and U7868 (N_7868,N_5249,N_5880);
nor U7869 (N_7869,N_5024,N_4550);
and U7870 (N_7870,N_4689,N_3961);
or U7871 (N_7871,N_4861,N_5900);
nand U7872 (N_7872,N_5717,N_3222);
and U7873 (N_7873,N_5451,N_5121);
nand U7874 (N_7874,N_4538,N_5565);
xor U7875 (N_7875,N_5000,N_5633);
nor U7876 (N_7876,N_4632,N_3728);
and U7877 (N_7877,N_5979,N_5634);
and U7878 (N_7878,N_3757,N_3210);
and U7879 (N_7879,N_3997,N_5469);
xnor U7880 (N_7880,N_3605,N_5128);
nand U7881 (N_7881,N_5644,N_3000);
or U7882 (N_7882,N_3307,N_4811);
nor U7883 (N_7883,N_4135,N_5489);
or U7884 (N_7884,N_5997,N_3189);
nor U7885 (N_7885,N_4035,N_5623);
nand U7886 (N_7886,N_3265,N_3093);
or U7887 (N_7887,N_5993,N_5423);
and U7888 (N_7888,N_3399,N_3441);
and U7889 (N_7889,N_5516,N_4944);
or U7890 (N_7890,N_5375,N_3636);
nand U7891 (N_7891,N_4252,N_4683);
nand U7892 (N_7892,N_5726,N_3185);
or U7893 (N_7893,N_4805,N_4476);
nand U7894 (N_7894,N_5266,N_5860);
or U7895 (N_7895,N_5620,N_4876);
nand U7896 (N_7896,N_5159,N_5590);
nand U7897 (N_7897,N_4708,N_4655);
nand U7898 (N_7898,N_3924,N_3351);
xor U7899 (N_7899,N_3750,N_5371);
and U7900 (N_7900,N_5054,N_3301);
nand U7901 (N_7901,N_4861,N_4204);
nor U7902 (N_7902,N_4852,N_5023);
nand U7903 (N_7903,N_5220,N_5335);
or U7904 (N_7904,N_4754,N_4562);
and U7905 (N_7905,N_4934,N_5128);
or U7906 (N_7906,N_3546,N_5897);
and U7907 (N_7907,N_4684,N_5991);
and U7908 (N_7908,N_3547,N_3737);
nor U7909 (N_7909,N_5813,N_4639);
xor U7910 (N_7910,N_3425,N_4223);
or U7911 (N_7911,N_3848,N_3784);
and U7912 (N_7912,N_5690,N_5457);
nor U7913 (N_7913,N_3383,N_4810);
nand U7914 (N_7914,N_5551,N_3651);
or U7915 (N_7915,N_5656,N_3458);
nor U7916 (N_7916,N_5188,N_4448);
nand U7917 (N_7917,N_4710,N_4514);
nand U7918 (N_7918,N_4917,N_4726);
nand U7919 (N_7919,N_5386,N_3209);
or U7920 (N_7920,N_4873,N_4303);
xor U7921 (N_7921,N_4274,N_4085);
nor U7922 (N_7922,N_4125,N_3295);
nor U7923 (N_7923,N_5882,N_4049);
nor U7924 (N_7924,N_5810,N_5165);
and U7925 (N_7925,N_5507,N_5002);
and U7926 (N_7926,N_4659,N_4760);
or U7927 (N_7927,N_4853,N_5477);
nor U7928 (N_7928,N_5337,N_4820);
or U7929 (N_7929,N_4663,N_4903);
nor U7930 (N_7930,N_3824,N_3523);
or U7931 (N_7931,N_5027,N_3381);
and U7932 (N_7932,N_5810,N_3296);
nand U7933 (N_7933,N_5962,N_4366);
or U7934 (N_7934,N_4173,N_3593);
or U7935 (N_7935,N_4337,N_4060);
and U7936 (N_7936,N_5898,N_3160);
nand U7937 (N_7937,N_5000,N_5523);
or U7938 (N_7938,N_5303,N_5188);
or U7939 (N_7939,N_4173,N_3141);
nor U7940 (N_7940,N_4145,N_5585);
nand U7941 (N_7941,N_5191,N_4377);
or U7942 (N_7942,N_3827,N_4538);
nand U7943 (N_7943,N_3104,N_3102);
and U7944 (N_7944,N_5503,N_3723);
and U7945 (N_7945,N_4998,N_4746);
nand U7946 (N_7946,N_4830,N_4476);
or U7947 (N_7947,N_3448,N_3864);
or U7948 (N_7948,N_4708,N_4203);
or U7949 (N_7949,N_5518,N_5289);
and U7950 (N_7950,N_5140,N_3411);
nor U7951 (N_7951,N_4381,N_5202);
or U7952 (N_7952,N_3982,N_3834);
nand U7953 (N_7953,N_4379,N_4474);
nand U7954 (N_7954,N_5390,N_4655);
and U7955 (N_7955,N_5665,N_4085);
or U7956 (N_7956,N_5646,N_4218);
or U7957 (N_7957,N_5383,N_3299);
xnor U7958 (N_7958,N_4966,N_3098);
and U7959 (N_7959,N_3944,N_3917);
nand U7960 (N_7960,N_3519,N_3933);
nand U7961 (N_7961,N_4258,N_5125);
nor U7962 (N_7962,N_4053,N_4820);
or U7963 (N_7963,N_3880,N_3041);
nor U7964 (N_7964,N_5212,N_3489);
nor U7965 (N_7965,N_5316,N_4814);
nor U7966 (N_7966,N_3910,N_3035);
and U7967 (N_7967,N_3351,N_5823);
nor U7968 (N_7968,N_5977,N_5662);
or U7969 (N_7969,N_5722,N_4853);
and U7970 (N_7970,N_4787,N_4104);
or U7971 (N_7971,N_5107,N_5834);
and U7972 (N_7972,N_4027,N_5049);
or U7973 (N_7973,N_3393,N_4834);
nor U7974 (N_7974,N_5678,N_4624);
or U7975 (N_7975,N_4640,N_4259);
or U7976 (N_7976,N_4110,N_3363);
or U7977 (N_7977,N_4129,N_5640);
nor U7978 (N_7978,N_5111,N_5433);
nor U7979 (N_7979,N_3567,N_3404);
or U7980 (N_7980,N_3378,N_4775);
and U7981 (N_7981,N_3317,N_4620);
or U7982 (N_7982,N_3163,N_3330);
and U7983 (N_7983,N_3317,N_4846);
nor U7984 (N_7984,N_5596,N_4228);
nand U7985 (N_7985,N_4517,N_3513);
and U7986 (N_7986,N_4366,N_5010);
or U7987 (N_7987,N_5891,N_3926);
and U7988 (N_7988,N_4944,N_5440);
nand U7989 (N_7989,N_5942,N_5794);
nor U7990 (N_7990,N_4466,N_4257);
nand U7991 (N_7991,N_3706,N_3910);
nor U7992 (N_7992,N_4413,N_4698);
and U7993 (N_7993,N_4573,N_4706);
or U7994 (N_7994,N_3902,N_5896);
nor U7995 (N_7995,N_3094,N_5953);
nand U7996 (N_7996,N_3075,N_5858);
or U7997 (N_7997,N_4069,N_4670);
and U7998 (N_7998,N_3028,N_3734);
or U7999 (N_7999,N_3392,N_5503);
nor U8000 (N_8000,N_3854,N_3772);
nor U8001 (N_8001,N_4157,N_4620);
or U8002 (N_8002,N_5443,N_3163);
nor U8003 (N_8003,N_4268,N_4321);
and U8004 (N_8004,N_3205,N_3162);
and U8005 (N_8005,N_3569,N_3993);
nor U8006 (N_8006,N_4889,N_4453);
nand U8007 (N_8007,N_5019,N_5582);
nor U8008 (N_8008,N_3814,N_3478);
nand U8009 (N_8009,N_3968,N_3245);
nor U8010 (N_8010,N_5700,N_5151);
or U8011 (N_8011,N_4761,N_4725);
nor U8012 (N_8012,N_4430,N_5799);
xor U8013 (N_8013,N_3105,N_5029);
nor U8014 (N_8014,N_5196,N_3548);
and U8015 (N_8015,N_3046,N_3602);
nand U8016 (N_8016,N_4616,N_3408);
nand U8017 (N_8017,N_4126,N_4835);
and U8018 (N_8018,N_4642,N_5632);
and U8019 (N_8019,N_5454,N_4894);
or U8020 (N_8020,N_3263,N_5861);
and U8021 (N_8021,N_3785,N_5811);
or U8022 (N_8022,N_4969,N_5632);
or U8023 (N_8023,N_4450,N_5391);
and U8024 (N_8024,N_5208,N_4413);
and U8025 (N_8025,N_4413,N_5847);
and U8026 (N_8026,N_4134,N_3073);
nor U8027 (N_8027,N_3600,N_4459);
or U8028 (N_8028,N_3996,N_5884);
nand U8029 (N_8029,N_5167,N_5804);
or U8030 (N_8030,N_5474,N_4227);
or U8031 (N_8031,N_5462,N_4247);
nor U8032 (N_8032,N_4324,N_3605);
nand U8033 (N_8033,N_4549,N_5984);
or U8034 (N_8034,N_3677,N_4128);
and U8035 (N_8035,N_4364,N_3807);
and U8036 (N_8036,N_4497,N_5316);
or U8037 (N_8037,N_3846,N_4219);
or U8038 (N_8038,N_5586,N_4194);
nand U8039 (N_8039,N_4199,N_4472);
nor U8040 (N_8040,N_5180,N_4924);
or U8041 (N_8041,N_5287,N_4177);
or U8042 (N_8042,N_5109,N_5644);
xor U8043 (N_8043,N_4245,N_5796);
and U8044 (N_8044,N_3202,N_3646);
and U8045 (N_8045,N_3128,N_4614);
nor U8046 (N_8046,N_3153,N_5022);
or U8047 (N_8047,N_4462,N_4391);
nor U8048 (N_8048,N_3543,N_5748);
and U8049 (N_8049,N_4116,N_4179);
nor U8050 (N_8050,N_4262,N_4895);
nor U8051 (N_8051,N_3851,N_3817);
nor U8052 (N_8052,N_4530,N_4266);
nand U8053 (N_8053,N_4959,N_4597);
and U8054 (N_8054,N_5162,N_5221);
and U8055 (N_8055,N_4418,N_5466);
and U8056 (N_8056,N_5660,N_4123);
or U8057 (N_8057,N_3154,N_4502);
or U8058 (N_8058,N_3350,N_5666);
or U8059 (N_8059,N_5397,N_4258);
nor U8060 (N_8060,N_4368,N_3052);
or U8061 (N_8061,N_4450,N_3778);
or U8062 (N_8062,N_4605,N_3214);
or U8063 (N_8063,N_5596,N_4235);
and U8064 (N_8064,N_5490,N_4161);
nor U8065 (N_8065,N_3381,N_3968);
or U8066 (N_8066,N_3710,N_4855);
or U8067 (N_8067,N_3835,N_3224);
nor U8068 (N_8068,N_4097,N_5080);
and U8069 (N_8069,N_4232,N_4323);
and U8070 (N_8070,N_5454,N_3753);
nand U8071 (N_8071,N_4607,N_5937);
nand U8072 (N_8072,N_5794,N_4720);
nand U8073 (N_8073,N_4692,N_3033);
nand U8074 (N_8074,N_4377,N_5855);
and U8075 (N_8075,N_5832,N_3138);
nor U8076 (N_8076,N_5302,N_4126);
or U8077 (N_8077,N_4476,N_5767);
and U8078 (N_8078,N_4596,N_5043);
nor U8079 (N_8079,N_4936,N_5088);
nor U8080 (N_8080,N_5946,N_4389);
nand U8081 (N_8081,N_3507,N_4845);
nand U8082 (N_8082,N_4980,N_3984);
nand U8083 (N_8083,N_3286,N_5117);
or U8084 (N_8084,N_4103,N_5779);
nand U8085 (N_8085,N_3045,N_4142);
or U8086 (N_8086,N_5841,N_3586);
nor U8087 (N_8087,N_3621,N_3072);
and U8088 (N_8088,N_4815,N_5896);
nor U8089 (N_8089,N_4688,N_5316);
or U8090 (N_8090,N_3965,N_3641);
nand U8091 (N_8091,N_4223,N_3410);
or U8092 (N_8092,N_4442,N_3143);
nand U8093 (N_8093,N_5880,N_3913);
nand U8094 (N_8094,N_5166,N_3873);
and U8095 (N_8095,N_4605,N_3533);
nand U8096 (N_8096,N_5656,N_3305);
or U8097 (N_8097,N_3963,N_4802);
or U8098 (N_8098,N_5023,N_4679);
and U8099 (N_8099,N_4262,N_4513);
or U8100 (N_8100,N_5469,N_5716);
or U8101 (N_8101,N_5443,N_3819);
nand U8102 (N_8102,N_5833,N_5248);
and U8103 (N_8103,N_4426,N_3321);
and U8104 (N_8104,N_4531,N_4166);
or U8105 (N_8105,N_3116,N_4747);
or U8106 (N_8106,N_5292,N_4481);
nand U8107 (N_8107,N_5629,N_4298);
nand U8108 (N_8108,N_5606,N_3308);
and U8109 (N_8109,N_4426,N_5659);
nand U8110 (N_8110,N_4223,N_3587);
nor U8111 (N_8111,N_3610,N_5483);
or U8112 (N_8112,N_3838,N_4136);
or U8113 (N_8113,N_4732,N_4328);
nor U8114 (N_8114,N_3933,N_5784);
or U8115 (N_8115,N_4021,N_4103);
nand U8116 (N_8116,N_3742,N_4504);
nand U8117 (N_8117,N_4386,N_3641);
nor U8118 (N_8118,N_3127,N_5187);
nor U8119 (N_8119,N_5594,N_3695);
nor U8120 (N_8120,N_4599,N_3108);
nor U8121 (N_8121,N_5243,N_3211);
nand U8122 (N_8122,N_3721,N_3275);
nor U8123 (N_8123,N_3087,N_4606);
and U8124 (N_8124,N_4225,N_5284);
nor U8125 (N_8125,N_3072,N_3317);
nand U8126 (N_8126,N_5053,N_5741);
nand U8127 (N_8127,N_3063,N_5504);
and U8128 (N_8128,N_4066,N_4146);
nor U8129 (N_8129,N_5467,N_4248);
and U8130 (N_8130,N_3706,N_5987);
nand U8131 (N_8131,N_4328,N_3524);
nor U8132 (N_8132,N_4226,N_5094);
nor U8133 (N_8133,N_4805,N_5004);
or U8134 (N_8134,N_4360,N_4533);
nand U8135 (N_8135,N_3664,N_5158);
nand U8136 (N_8136,N_5380,N_4350);
nor U8137 (N_8137,N_4547,N_4612);
nand U8138 (N_8138,N_3872,N_3750);
or U8139 (N_8139,N_3947,N_5279);
nand U8140 (N_8140,N_5109,N_3830);
or U8141 (N_8141,N_4678,N_3438);
or U8142 (N_8142,N_5167,N_5471);
and U8143 (N_8143,N_4434,N_4780);
nand U8144 (N_8144,N_5895,N_4048);
and U8145 (N_8145,N_5092,N_4286);
and U8146 (N_8146,N_4091,N_3311);
nand U8147 (N_8147,N_4952,N_3258);
or U8148 (N_8148,N_4572,N_5124);
xnor U8149 (N_8149,N_3853,N_5616);
nand U8150 (N_8150,N_5780,N_5563);
nand U8151 (N_8151,N_5274,N_4928);
or U8152 (N_8152,N_3371,N_5942);
and U8153 (N_8153,N_4500,N_4363);
or U8154 (N_8154,N_3793,N_5061);
and U8155 (N_8155,N_4891,N_5375);
and U8156 (N_8156,N_4218,N_5618);
nand U8157 (N_8157,N_5483,N_5398);
nand U8158 (N_8158,N_3991,N_4433);
nand U8159 (N_8159,N_3740,N_4304);
and U8160 (N_8160,N_3260,N_4220);
nor U8161 (N_8161,N_4476,N_3342);
nand U8162 (N_8162,N_5818,N_4262);
nand U8163 (N_8163,N_4173,N_5385);
and U8164 (N_8164,N_4454,N_5031);
and U8165 (N_8165,N_5464,N_4783);
nand U8166 (N_8166,N_5895,N_3118);
nor U8167 (N_8167,N_5739,N_3648);
or U8168 (N_8168,N_5255,N_4770);
nand U8169 (N_8169,N_5674,N_3167);
nor U8170 (N_8170,N_5814,N_5678);
or U8171 (N_8171,N_4215,N_4053);
nand U8172 (N_8172,N_3983,N_5731);
or U8173 (N_8173,N_5532,N_3429);
and U8174 (N_8174,N_3533,N_3975);
nor U8175 (N_8175,N_3634,N_4961);
nor U8176 (N_8176,N_3562,N_5050);
or U8177 (N_8177,N_5473,N_4063);
nor U8178 (N_8178,N_5778,N_3717);
nand U8179 (N_8179,N_5246,N_5157);
and U8180 (N_8180,N_4180,N_3993);
nor U8181 (N_8181,N_5296,N_3414);
and U8182 (N_8182,N_5294,N_3848);
nand U8183 (N_8183,N_3477,N_5692);
or U8184 (N_8184,N_4609,N_5637);
nand U8185 (N_8185,N_3399,N_4214);
or U8186 (N_8186,N_3500,N_3518);
or U8187 (N_8187,N_4082,N_5825);
nand U8188 (N_8188,N_5996,N_3598);
and U8189 (N_8189,N_3300,N_5314);
nand U8190 (N_8190,N_3887,N_3970);
nand U8191 (N_8191,N_5499,N_3909);
nand U8192 (N_8192,N_4500,N_5265);
or U8193 (N_8193,N_5603,N_5971);
nand U8194 (N_8194,N_5150,N_3737);
and U8195 (N_8195,N_4606,N_5883);
and U8196 (N_8196,N_3697,N_4657);
or U8197 (N_8197,N_3953,N_5197);
nand U8198 (N_8198,N_5544,N_3340);
nor U8199 (N_8199,N_3004,N_3141);
nor U8200 (N_8200,N_3848,N_5793);
and U8201 (N_8201,N_4403,N_3057);
and U8202 (N_8202,N_4182,N_4822);
or U8203 (N_8203,N_5031,N_3515);
or U8204 (N_8204,N_3087,N_3037);
nand U8205 (N_8205,N_4773,N_3368);
nor U8206 (N_8206,N_4001,N_3045);
or U8207 (N_8207,N_4917,N_3116);
nor U8208 (N_8208,N_5420,N_5196);
nand U8209 (N_8209,N_5117,N_4012);
nand U8210 (N_8210,N_4472,N_5822);
nand U8211 (N_8211,N_4406,N_5929);
or U8212 (N_8212,N_4820,N_4513);
and U8213 (N_8213,N_5313,N_4487);
and U8214 (N_8214,N_3752,N_3620);
and U8215 (N_8215,N_5527,N_5997);
nor U8216 (N_8216,N_4779,N_3176);
and U8217 (N_8217,N_5636,N_3891);
nor U8218 (N_8218,N_5716,N_4566);
nor U8219 (N_8219,N_3629,N_5348);
or U8220 (N_8220,N_3666,N_4691);
and U8221 (N_8221,N_4247,N_4759);
and U8222 (N_8222,N_3942,N_4420);
nand U8223 (N_8223,N_4168,N_3338);
nor U8224 (N_8224,N_3509,N_5318);
or U8225 (N_8225,N_3317,N_3949);
or U8226 (N_8226,N_4195,N_3935);
and U8227 (N_8227,N_4516,N_4828);
nor U8228 (N_8228,N_3752,N_4466);
nand U8229 (N_8229,N_4948,N_5598);
nor U8230 (N_8230,N_5901,N_4432);
or U8231 (N_8231,N_5969,N_4419);
nor U8232 (N_8232,N_5249,N_3543);
and U8233 (N_8233,N_3498,N_5232);
or U8234 (N_8234,N_3702,N_3449);
nor U8235 (N_8235,N_5972,N_4981);
nor U8236 (N_8236,N_4839,N_4598);
or U8237 (N_8237,N_3221,N_5005);
or U8238 (N_8238,N_3586,N_4675);
nor U8239 (N_8239,N_5030,N_3625);
and U8240 (N_8240,N_5333,N_5121);
or U8241 (N_8241,N_5542,N_3735);
or U8242 (N_8242,N_3243,N_3013);
nand U8243 (N_8243,N_5118,N_3100);
and U8244 (N_8244,N_3974,N_4084);
nor U8245 (N_8245,N_5134,N_5163);
nor U8246 (N_8246,N_4540,N_3361);
or U8247 (N_8247,N_3609,N_3793);
or U8248 (N_8248,N_5380,N_3058);
nand U8249 (N_8249,N_3379,N_5059);
or U8250 (N_8250,N_3873,N_4055);
nor U8251 (N_8251,N_3320,N_5401);
nor U8252 (N_8252,N_5351,N_5881);
nor U8253 (N_8253,N_4497,N_4744);
and U8254 (N_8254,N_5228,N_5410);
and U8255 (N_8255,N_4695,N_4998);
nand U8256 (N_8256,N_3719,N_5100);
and U8257 (N_8257,N_3160,N_5114);
or U8258 (N_8258,N_5358,N_4645);
or U8259 (N_8259,N_4194,N_3381);
nor U8260 (N_8260,N_3854,N_5090);
nand U8261 (N_8261,N_3778,N_3985);
and U8262 (N_8262,N_3765,N_5332);
and U8263 (N_8263,N_3659,N_5765);
and U8264 (N_8264,N_4057,N_4490);
nor U8265 (N_8265,N_3593,N_5483);
nor U8266 (N_8266,N_4729,N_4187);
nor U8267 (N_8267,N_4241,N_3137);
or U8268 (N_8268,N_4594,N_4005);
nor U8269 (N_8269,N_5772,N_5250);
xnor U8270 (N_8270,N_5421,N_5533);
nand U8271 (N_8271,N_3137,N_4394);
or U8272 (N_8272,N_3725,N_5018);
and U8273 (N_8273,N_4248,N_3549);
nor U8274 (N_8274,N_5260,N_3169);
nor U8275 (N_8275,N_4250,N_4363);
and U8276 (N_8276,N_5018,N_4985);
nor U8277 (N_8277,N_3917,N_3271);
nor U8278 (N_8278,N_5443,N_3515);
xnor U8279 (N_8279,N_3087,N_4184);
or U8280 (N_8280,N_5701,N_3893);
nor U8281 (N_8281,N_4277,N_3375);
nand U8282 (N_8282,N_5242,N_4709);
and U8283 (N_8283,N_5101,N_5796);
nand U8284 (N_8284,N_4484,N_5584);
or U8285 (N_8285,N_5504,N_3271);
or U8286 (N_8286,N_4697,N_4463);
or U8287 (N_8287,N_5306,N_3470);
or U8288 (N_8288,N_5777,N_5539);
nor U8289 (N_8289,N_3156,N_5663);
and U8290 (N_8290,N_4396,N_4041);
or U8291 (N_8291,N_5518,N_4292);
or U8292 (N_8292,N_5287,N_3861);
or U8293 (N_8293,N_4746,N_3915);
or U8294 (N_8294,N_5290,N_4204);
nor U8295 (N_8295,N_5515,N_3053);
or U8296 (N_8296,N_3501,N_3268);
nand U8297 (N_8297,N_4966,N_4587);
or U8298 (N_8298,N_3235,N_4322);
nor U8299 (N_8299,N_4045,N_3515);
nand U8300 (N_8300,N_4811,N_4525);
and U8301 (N_8301,N_3296,N_3260);
and U8302 (N_8302,N_4716,N_4467);
nor U8303 (N_8303,N_3183,N_3389);
and U8304 (N_8304,N_5030,N_4834);
and U8305 (N_8305,N_3322,N_3737);
and U8306 (N_8306,N_5806,N_4163);
or U8307 (N_8307,N_4601,N_5510);
nand U8308 (N_8308,N_3172,N_4173);
and U8309 (N_8309,N_5866,N_5185);
nor U8310 (N_8310,N_3333,N_5362);
or U8311 (N_8311,N_4504,N_3935);
or U8312 (N_8312,N_4129,N_5934);
nor U8313 (N_8313,N_3456,N_4440);
and U8314 (N_8314,N_5877,N_4581);
or U8315 (N_8315,N_3930,N_4973);
and U8316 (N_8316,N_4921,N_4870);
xor U8317 (N_8317,N_3537,N_5865);
and U8318 (N_8318,N_5526,N_4521);
nand U8319 (N_8319,N_3796,N_4389);
or U8320 (N_8320,N_3359,N_5995);
nor U8321 (N_8321,N_5602,N_5111);
nand U8322 (N_8322,N_3913,N_4295);
and U8323 (N_8323,N_3830,N_3275);
xor U8324 (N_8324,N_3725,N_3043);
nor U8325 (N_8325,N_5568,N_3878);
nand U8326 (N_8326,N_4136,N_3087);
nand U8327 (N_8327,N_3858,N_3957);
nand U8328 (N_8328,N_3168,N_5139);
or U8329 (N_8329,N_3360,N_5052);
or U8330 (N_8330,N_5245,N_3554);
or U8331 (N_8331,N_4035,N_4973);
nor U8332 (N_8332,N_4357,N_4997);
or U8333 (N_8333,N_5437,N_4137);
nor U8334 (N_8334,N_4990,N_3934);
and U8335 (N_8335,N_3224,N_4098);
nor U8336 (N_8336,N_3092,N_4949);
or U8337 (N_8337,N_3637,N_5739);
and U8338 (N_8338,N_5278,N_5035);
and U8339 (N_8339,N_3483,N_3574);
and U8340 (N_8340,N_3331,N_5105);
nand U8341 (N_8341,N_4832,N_5749);
and U8342 (N_8342,N_4546,N_5832);
or U8343 (N_8343,N_4737,N_3027);
nor U8344 (N_8344,N_4085,N_4314);
nand U8345 (N_8345,N_4339,N_4882);
or U8346 (N_8346,N_5051,N_3661);
nor U8347 (N_8347,N_4406,N_3109);
nor U8348 (N_8348,N_4130,N_5817);
or U8349 (N_8349,N_3926,N_4336);
and U8350 (N_8350,N_3829,N_5096);
or U8351 (N_8351,N_5283,N_3949);
nor U8352 (N_8352,N_5104,N_4114);
nor U8353 (N_8353,N_5864,N_3273);
or U8354 (N_8354,N_3119,N_3143);
and U8355 (N_8355,N_5482,N_5396);
nand U8356 (N_8356,N_3042,N_5701);
nor U8357 (N_8357,N_3044,N_5674);
nor U8358 (N_8358,N_5400,N_3677);
or U8359 (N_8359,N_5712,N_3691);
nor U8360 (N_8360,N_3924,N_4703);
nand U8361 (N_8361,N_3228,N_4358);
nand U8362 (N_8362,N_5197,N_4450);
or U8363 (N_8363,N_3927,N_4001);
nand U8364 (N_8364,N_5614,N_3218);
nor U8365 (N_8365,N_5735,N_5278);
nand U8366 (N_8366,N_3902,N_4947);
nor U8367 (N_8367,N_4834,N_4035);
nor U8368 (N_8368,N_5805,N_4649);
and U8369 (N_8369,N_3862,N_3928);
nand U8370 (N_8370,N_5925,N_5143);
and U8371 (N_8371,N_5662,N_3981);
and U8372 (N_8372,N_5052,N_3936);
and U8373 (N_8373,N_5833,N_5106);
nor U8374 (N_8374,N_3007,N_4231);
nor U8375 (N_8375,N_5341,N_3248);
or U8376 (N_8376,N_4206,N_5802);
nand U8377 (N_8377,N_5804,N_5928);
and U8378 (N_8378,N_5683,N_4439);
nand U8379 (N_8379,N_3255,N_4424);
nor U8380 (N_8380,N_5229,N_4743);
or U8381 (N_8381,N_4196,N_5218);
or U8382 (N_8382,N_4171,N_4507);
nor U8383 (N_8383,N_3364,N_3378);
or U8384 (N_8384,N_4462,N_5170);
or U8385 (N_8385,N_4157,N_4729);
nand U8386 (N_8386,N_5866,N_5014);
and U8387 (N_8387,N_5421,N_3425);
nor U8388 (N_8388,N_4364,N_4830);
nand U8389 (N_8389,N_4421,N_5852);
nand U8390 (N_8390,N_4532,N_5043);
nor U8391 (N_8391,N_3294,N_5743);
or U8392 (N_8392,N_3951,N_4975);
nor U8393 (N_8393,N_5742,N_4037);
nand U8394 (N_8394,N_4434,N_5784);
nor U8395 (N_8395,N_5410,N_3404);
and U8396 (N_8396,N_4625,N_4282);
and U8397 (N_8397,N_3039,N_3177);
nand U8398 (N_8398,N_3643,N_3911);
nor U8399 (N_8399,N_4334,N_3986);
and U8400 (N_8400,N_4232,N_4744);
nand U8401 (N_8401,N_4958,N_3309);
and U8402 (N_8402,N_4291,N_5673);
and U8403 (N_8403,N_4484,N_4420);
nand U8404 (N_8404,N_3762,N_4236);
or U8405 (N_8405,N_5193,N_3239);
or U8406 (N_8406,N_5122,N_3142);
nor U8407 (N_8407,N_5470,N_3698);
and U8408 (N_8408,N_4797,N_3722);
and U8409 (N_8409,N_3431,N_4306);
xnor U8410 (N_8410,N_3858,N_3522);
nand U8411 (N_8411,N_5518,N_5443);
nor U8412 (N_8412,N_5526,N_3421);
nand U8413 (N_8413,N_3765,N_5488);
nand U8414 (N_8414,N_3553,N_3266);
and U8415 (N_8415,N_3029,N_3869);
nand U8416 (N_8416,N_4930,N_3006);
or U8417 (N_8417,N_5729,N_5513);
nand U8418 (N_8418,N_4373,N_5955);
and U8419 (N_8419,N_5615,N_4611);
or U8420 (N_8420,N_4677,N_3867);
or U8421 (N_8421,N_4761,N_4441);
or U8422 (N_8422,N_5338,N_4311);
nand U8423 (N_8423,N_4499,N_4569);
nand U8424 (N_8424,N_4757,N_4971);
nor U8425 (N_8425,N_5950,N_4982);
nor U8426 (N_8426,N_4759,N_5388);
or U8427 (N_8427,N_5439,N_5900);
nor U8428 (N_8428,N_4296,N_4694);
nor U8429 (N_8429,N_5078,N_5152);
nor U8430 (N_8430,N_4141,N_5476);
nor U8431 (N_8431,N_3599,N_5760);
or U8432 (N_8432,N_4635,N_3426);
and U8433 (N_8433,N_5620,N_3712);
nor U8434 (N_8434,N_4888,N_3372);
or U8435 (N_8435,N_5460,N_3465);
and U8436 (N_8436,N_4333,N_4555);
and U8437 (N_8437,N_3107,N_4316);
nand U8438 (N_8438,N_3805,N_5054);
nor U8439 (N_8439,N_5712,N_3533);
or U8440 (N_8440,N_4842,N_4202);
nand U8441 (N_8441,N_3676,N_3650);
nor U8442 (N_8442,N_4094,N_4173);
nand U8443 (N_8443,N_5976,N_4694);
or U8444 (N_8444,N_5551,N_5285);
and U8445 (N_8445,N_4375,N_3655);
nand U8446 (N_8446,N_4630,N_5801);
and U8447 (N_8447,N_5066,N_4523);
nor U8448 (N_8448,N_4563,N_3774);
and U8449 (N_8449,N_3420,N_4039);
or U8450 (N_8450,N_4990,N_5672);
and U8451 (N_8451,N_3465,N_4564);
nand U8452 (N_8452,N_4350,N_5997);
nor U8453 (N_8453,N_3449,N_3374);
nand U8454 (N_8454,N_4930,N_5225);
and U8455 (N_8455,N_4191,N_3954);
xor U8456 (N_8456,N_5851,N_3103);
nor U8457 (N_8457,N_3227,N_5199);
or U8458 (N_8458,N_4804,N_3823);
nand U8459 (N_8459,N_3778,N_4316);
and U8460 (N_8460,N_5692,N_4454);
nand U8461 (N_8461,N_4971,N_4931);
nor U8462 (N_8462,N_4623,N_5383);
nor U8463 (N_8463,N_5408,N_5597);
nand U8464 (N_8464,N_5537,N_5929);
and U8465 (N_8465,N_3028,N_5698);
nand U8466 (N_8466,N_5987,N_4061);
or U8467 (N_8467,N_4011,N_5681);
and U8468 (N_8468,N_3552,N_4034);
or U8469 (N_8469,N_3108,N_4071);
and U8470 (N_8470,N_4461,N_3993);
and U8471 (N_8471,N_4231,N_3614);
or U8472 (N_8472,N_5279,N_5567);
and U8473 (N_8473,N_4422,N_4808);
and U8474 (N_8474,N_4889,N_3086);
and U8475 (N_8475,N_5735,N_5437);
nor U8476 (N_8476,N_3589,N_3036);
or U8477 (N_8477,N_5640,N_3249);
and U8478 (N_8478,N_3541,N_3114);
nor U8479 (N_8479,N_3981,N_4948);
nor U8480 (N_8480,N_4895,N_3756);
or U8481 (N_8481,N_4598,N_4583);
or U8482 (N_8482,N_3271,N_4364);
and U8483 (N_8483,N_3023,N_4889);
nand U8484 (N_8484,N_3142,N_3603);
or U8485 (N_8485,N_3075,N_3140);
nand U8486 (N_8486,N_4353,N_3857);
and U8487 (N_8487,N_5743,N_3773);
nand U8488 (N_8488,N_5566,N_4545);
nand U8489 (N_8489,N_5870,N_4566);
and U8490 (N_8490,N_3311,N_3446);
or U8491 (N_8491,N_4897,N_4327);
nor U8492 (N_8492,N_3257,N_5128);
and U8493 (N_8493,N_3147,N_3619);
nor U8494 (N_8494,N_4283,N_3006);
or U8495 (N_8495,N_4296,N_3210);
or U8496 (N_8496,N_4594,N_3680);
nand U8497 (N_8497,N_3088,N_5866);
or U8498 (N_8498,N_3374,N_3277);
nand U8499 (N_8499,N_4340,N_4164);
nand U8500 (N_8500,N_3305,N_4852);
nor U8501 (N_8501,N_3963,N_3868);
and U8502 (N_8502,N_3617,N_5123);
nor U8503 (N_8503,N_4750,N_3753);
nand U8504 (N_8504,N_4874,N_4598);
and U8505 (N_8505,N_4459,N_5004);
or U8506 (N_8506,N_4899,N_3865);
nor U8507 (N_8507,N_3629,N_4245);
and U8508 (N_8508,N_5654,N_3450);
and U8509 (N_8509,N_3205,N_5710);
and U8510 (N_8510,N_5574,N_3620);
nor U8511 (N_8511,N_4578,N_3619);
nor U8512 (N_8512,N_4292,N_5219);
nand U8513 (N_8513,N_4055,N_5743);
and U8514 (N_8514,N_3174,N_5627);
xor U8515 (N_8515,N_5518,N_5989);
nand U8516 (N_8516,N_3105,N_3511);
nand U8517 (N_8517,N_5767,N_3338);
and U8518 (N_8518,N_4556,N_3261);
nor U8519 (N_8519,N_5890,N_4336);
nand U8520 (N_8520,N_5008,N_5420);
or U8521 (N_8521,N_3084,N_5090);
nand U8522 (N_8522,N_3701,N_3482);
or U8523 (N_8523,N_5490,N_4611);
xor U8524 (N_8524,N_3821,N_3830);
or U8525 (N_8525,N_5091,N_3883);
and U8526 (N_8526,N_4699,N_5177);
nand U8527 (N_8527,N_4982,N_5748);
nand U8528 (N_8528,N_4457,N_4439);
nand U8529 (N_8529,N_4925,N_5967);
and U8530 (N_8530,N_4118,N_5761);
and U8531 (N_8531,N_3848,N_4098);
nor U8532 (N_8532,N_3628,N_3816);
or U8533 (N_8533,N_4369,N_5307);
nor U8534 (N_8534,N_3840,N_4102);
nand U8535 (N_8535,N_4456,N_3848);
xnor U8536 (N_8536,N_4660,N_5915);
nand U8537 (N_8537,N_3599,N_5914);
nand U8538 (N_8538,N_3455,N_5278);
nor U8539 (N_8539,N_5574,N_3339);
and U8540 (N_8540,N_4495,N_3948);
or U8541 (N_8541,N_4471,N_4064);
and U8542 (N_8542,N_5681,N_4796);
nand U8543 (N_8543,N_3724,N_4895);
and U8544 (N_8544,N_5596,N_3325);
nand U8545 (N_8545,N_3844,N_4723);
and U8546 (N_8546,N_4906,N_4816);
nor U8547 (N_8547,N_3921,N_3753);
nor U8548 (N_8548,N_4975,N_3923);
or U8549 (N_8549,N_5988,N_5579);
nand U8550 (N_8550,N_5647,N_5090);
and U8551 (N_8551,N_3492,N_5807);
nor U8552 (N_8552,N_3877,N_5343);
or U8553 (N_8553,N_4264,N_4713);
and U8554 (N_8554,N_4218,N_4861);
nor U8555 (N_8555,N_4894,N_4189);
or U8556 (N_8556,N_5891,N_3640);
or U8557 (N_8557,N_4750,N_3673);
or U8558 (N_8558,N_4199,N_4285);
or U8559 (N_8559,N_5902,N_4642);
or U8560 (N_8560,N_3434,N_3158);
or U8561 (N_8561,N_3700,N_5616);
and U8562 (N_8562,N_3176,N_3186);
nor U8563 (N_8563,N_3462,N_3177);
and U8564 (N_8564,N_5131,N_5788);
or U8565 (N_8565,N_5216,N_4744);
nor U8566 (N_8566,N_3012,N_5260);
nand U8567 (N_8567,N_3638,N_5716);
nand U8568 (N_8568,N_5179,N_4480);
and U8569 (N_8569,N_4008,N_5406);
and U8570 (N_8570,N_5218,N_5896);
and U8571 (N_8571,N_3718,N_3471);
or U8572 (N_8572,N_5624,N_4470);
nand U8573 (N_8573,N_4981,N_3652);
and U8574 (N_8574,N_4326,N_3016);
nand U8575 (N_8575,N_3724,N_4188);
nand U8576 (N_8576,N_3476,N_3610);
and U8577 (N_8577,N_4700,N_3040);
nand U8578 (N_8578,N_4475,N_4908);
nand U8579 (N_8579,N_3887,N_3656);
nor U8580 (N_8580,N_3577,N_3293);
nor U8581 (N_8581,N_4041,N_4693);
or U8582 (N_8582,N_4901,N_3423);
or U8583 (N_8583,N_5730,N_3631);
nor U8584 (N_8584,N_3433,N_3145);
nand U8585 (N_8585,N_4189,N_4332);
nor U8586 (N_8586,N_4095,N_5787);
nor U8587 (N_8587,N_5046,N_5022);
nand U8588 (N_8588,N_4736,N_5305);
nand U8589 (N_8589,N_3124,N_4103);
nor U8590 (N_8590,N_4567,N_4841);
nand U8591 (N_8591,N_5597,N_3205);
and U8592 (N_8592,N_5463,N_5554);
and U8593 (N_8593,N_3874,N_3259);
nand U8594 (N_8594,N_5413,N_4603);
nand U8595 (N_8595,N_3841,N_5815);
nor U8596 (N_8596,N_3311,N_4152);
nand U8597 (N_8597,N_4208,N_4078);
or U8598 (N_8598,N_4894,N_5972);
or U8599 (N_8599,N_4590,N_5547);
nand U8600 (N_8600,N_4901,N_5172);
nand U8601 (N_8601,N_4430,N_4950);
and U8602 (N_8602,N_4295,N_4927);
or U8603 (N_8603,N_3451,N_5678);
nor U8604 (N_8604,N_5535,N_5939);
nor U8605 (N_8605,N_5011,N_5842);
nand U8606 (N_8606,N_3027,N_3362);
xnor U8607 (N_8607,N_4147,N_4265);
nand U8608 (N_8608,N_3627,N_4443);
nand U8609 (N_8609,N_3943,N_3864);
nor U8610 (N_8610,N_5807,N_3309);
or U8611 (N_8611,N_4527,N_4026);
nand U8612 (N_8612,N_5044,N_5322);
nor U8613 (N_8613,N_4196,N_4585);
and U8614 (N_8614,N_5257,N_3876);
nand U8615 (N_8615,N_4898,N_5444);
nor U8616 (N_8616,N_3420,N_4640);
and U8617 (N_8617,N_5996,N_4031);
nand U8618 (N_8618,N_4339,N_4140);
and U8619 (N_8619,N_4326,N_3918);
nor U8620 (N_8620,N_4322,N_5079);
and U8621 (N_8621,N_5180,N_5961);
or U8622 (N_8622,N_5211,N_3282);
nand U8623 (N_8623,N_5450,N_5801);
nor U8624 (N_8624,N_3800,N_3971);
nor U8625 (N_8625,N_5566,N_3097);
and U8626 (N_8626,N_4930,N_5384);
and U8627 (N_8627,N_5829,N_4581);
or U8628 (N_8628,N_5992,N_5163);
or U8629 (N_8629,N_5585,N_5203);
and U8630 (N_8630,N_5278,N_5457);
nor U8631 (N_8631,N_3982,N_4262);
nand U8632 (N_8632,N_4180,N_4963);
and U8633 (N_8633,N_5034,N_4470);
nand U8634 (N_8634,N_3257,N_4349);
or U8635 (N_8635,N_3099,N_5728);
and U8636 (N_8636,N_5516,N_4460);
or U8637 (N_8637,N_5457,N_3054);
or U8638 (N_8638,N_4933,N_3452);
nand U8639 (N_8639,N_3221,N_5980);
xnor U8640 (N_8640,N_5587,N_3944);
or U8641 (N_8641,N_5242,N_5456);
or U8642 (N_8642,N_5857,N_3488);
and U8643 (N_8643,N_5741,N_5730);
and U8644 (N_8644,N_4072,N_5110);
and U8645 (N_8645,N_5870,N_3455);
nor U8646 (N_8646,N_4389,N_5688);
nor U8647 (N_8647,N_3086,N_3934);
nor U8648 (N_8648,N_4598,N_3813);
and U8649 (N_8649,N_3097,N_5677);
and U8650 (N_8650,N_3083,N_3226);
xor U8651 (N_8651,N_3050,N_5102);
and U8652 (N_8652,N_5797,N_4276);
or U8653 (N_8653,N_4075,N_5617);
xor U8654 (N_8654,N_5744,N_4541);
nand U8655 (N_8655,N_3914,N_5501);
or U8656 (N_8656,N_5481,N_3675);
nor U8657 (N_8657,N_4092,N_3317);
or U8658 (N_8658,N_3481,N_3655);
and U8659 (N_8659,N_4853,N_3481);
nand U8660 (N_8660,N_4100,N_4902);
nor U8661 (N_8661,N_5933,N_4061);
nand U8662 (N_8662,N_5438,N_4701);
or U8663 (N_8663,N_4163,N_3969);
or U8664 (N_8664,N_3234,N_4857);
or U8665 (N_8665,N_5211,N_4428);
or U8666 (N_8666,N_5530,N_5967);
and U8667 (N_8667,N_4166,N_3467);
or U8668 (N_8668,N_3032,N_5047);
nor U8669 (N_8669,N_5508,N_5809);
nor U8670 (N_8670,N_3210,N_3284);
and U8671 (N_8671,N_5621,N_4361);
nor U8672 (N_8672,N_5125,N_5304);
and U8673 (N_8673,N_3560,N_5543);
nor U8674 (N_8674,N_3486,N_3094);
and U8675 (N_8675,N_3185,N_3845);
or U8676 (N_8676,N_5249,N_5038);
and U8677 (N_8677,N_5573,N_4989);
nand U8678 (N_8678,N_4450,N_3220);
and U8679 (N_8679,N_5991,N_4328);
and U8680 (N_8680,N_5368,N_5182);
and U8681 (N_8681,N_5633,N_3101);
nor U8682 (N_8682,N_4574,N_4450);
and U8683 (N_8683,N_5167,N_3064);
or U8684 (N_8684,N_4468,N_5225);
or U8685 (N_8685,N_5112,N_4382);
and U8686 (N_8686,N_3105,N_4797);
and U8687 (N_8687,N_4177,N_4325);
nand U8688 (N_8688,N_4251,N_4038);
and U8689 (N_8689,N_4131,N_3540);
and U8690 (N_8690,N_4609,N_5176);
nor U8691 (N_8691,N_3137,N_4926);
nor U8692 (N_8692,N_5889,N_5730);
nor U8693 (N_8693,N_3785,N_4033);
or U8694 (N_8694,N_4301,N_4611);
or U8695 (N_8695,N_3805,N_4229);
nor U8696 (N_8696,N_4956,N_3529);
and U8697 (N_8697,N_5481,N_5165);
or U8698 (N_8698,N_4483,N_4549);
nand U8699 (N_8699,N_5125,N_4983);
nor U8700 (N_8700,N_4808,N_3313);
nor U8701 (N_8701,N_5566,N_3137);
or U8702 (N_8702,N_3056,N_5561);
and U8703 (N_8703,N_3144,N_3234);
nor U8704 (N_8704,N_4349,N_3717);
nand U8705 (N_8705,N_4301,N_5816);
nor U8706 (N_8706,N_4504,N_3110);
nand U8707 (N_8707,N_3172,N_4760);
nor U8708 (N_8708,N_3372,N_5286);
nor U8709 (N_8709,N_5778,N_5757);
or U8710 (N_8710,N_4895,N_5291);
nor U8711 (N_8711,N_3601,N_3427);
nand U8712 (N_8712,N_4895,N_4947);
or U8713 (N_8713,N_4214,N_4682);
nand U8714 (N_8714,N_4143,N_5831);
nor U8715 (N_8715,N_5796,N_5045);
nand U8716 (N_8716,N_5145,N_5627);
and U8717 (N_8717,N_4397,N_4082);
nor U8718 (N_8718,N_3905,N_4786);
or U8719 (N_8719,N_4605,N_5533);
and U8720 (N_8720,N_4814,N_3222);
and U8721 (N_8721,N_5649,N_4444);
or U8722 (N_8722,N_4524,N_5288);
nor U8723 (N_8723,N_5443,N_3255);
or U8724 (N_8724,N_4630,N_4805);
or U8725 (N_8725,N_3210,N_5670);
and U8726 (N_8726,N_3269,N_5352);
nand U8727 (N_8727,N_4974,N_3421);
or U8728 (N_8728,N_5937,N_3329);
or U8729 (N_8729,N_5481,N_5980);
and U8730 (N_8730,N_3843,N_4059);
xnor U8731 (N_8731,N_4704,N_4664);
nand U8732 (N_8732,N_3691,N_4583);
or U8733 (N_8733,N_4470,N_3920);
nand U8734 (N_8734,N_3108,N_5861);
nor U8735 (N_8735,N_3182,N_5539);
nand U8736 (N_8736,N_3768,N_3288);
or U8737 (N_8737,N_5387,N_4637);
nor U8738 (N_8738,N_5359,N_3568);
nor U8739 (N_8739,N_3616,N_5650);
and U8740 (N_8740,N_4022,N_3845);
nor U8741 (N_8741,N_5598,N_5446);
nand U8742 (N_8742,N_3718,N_3046);
nand U8743 (N_8743,N_3299,N_4729);
or U8744 (N_8744,N_4638,N_3161);
or U8745 (N_8745,N_3554,N_4487);
nor U8746 (N_8746,N_5366,N_4318);
and U8747 (N_8747,N_4139,N_4733);
or U8748 (N_8748,N_4701,N_3036);
nand U8749 (N_8749,N_4132,N_3743);
nand U8750 (N_8750,N_3393,N_5932);
and U8751 (N_8751,N_5584,N_3162);
nor U8752 (N_8752,N_5256,N_3179);
nand U8753 (N_8753,N_3483,N_3217);
nor U8754 (N_8754,N_4455,N_3438);
or U8755 (N_8755,N_3492,N_5922);
and U8756 (N_8756,N_5253,N_5124);
nor U8757 (N_8757,N_3835,N_3248);
nor U8758 (N_8758,N_4430,N_3605);
nand U8759 (N_8759,N_5410,N_3108);
nand U8760 (N_8760,N_3577,N_3299);
or U8761 (N_8761,N_4903,N_4244);
or U8762 (N_8762,N_3912,N_4137);
and U8763 (N_8763,N_3662,N_5228);
or U8764 (N_8764,N_3913,N_4850);
nand U8765 (N_8765,N_4296,N_4254);
nand U8766 (N_8766,N_3723,N_3516);
or U8767 (N_8767,N_3898,N_5146);
and U8768 (N_8768,N_3392,N_3162);
and U8769 (N_8769,N_4816,N_5755);
nor U8770 (N_8770,N_5523,N_3527);
nor U8771 (N_8771,N_3959,N_3201);
or U8772 (N_8772,N_5894,N_3734);
and U8773 (N_8773,N_3164,N_3895);
nand U8774 (N_8774,N_3628,N_3194);
nand U8775 (N_8775,N_4504,N_4366);
and U8776 (N_8776,N_5848,N_5582);
nand U8777 (N_8777,N_3226,N_5997);
or U8778 (N_8778,N_5721,N_4433);
and U8779 (N_8779,N_4792,N_4814);
nand U8780 (N_8780,N_5648,N_4992);
or U8781 (N_8781,N_4986,N_3218);
nand U8782 (N_8782,N_3925,N_5881);
or U8783 (N_8783,N_3246,N_5742);
nor U8784 (N_8784,N_5022,N_4595);
and U8785 (N_8785,N_4858,N_4337);
nand U8786 (N_8786,N_3134,N_4498);
nor U8787 (N_8787,N_5854,N_3567);
nor U8788 (N_8788,N_4689,N_5066);
nand U8789 (N_8789,N_5541,N_5129);
xnor U8790 (N_8790,N_3931,N_4266);
nand U8791 (N_8791,N_3963,N_4348);
or U8792 (N_8792,N_5346,N_3840);
and U8793 (N_8793,N_5981,N_4612);
nor U8794 (N_8794,N_5704,N_4695);
nand U8795 (N_8795,N_5005,N_3037);
and U8796 (N_8796,N_3993,N_3622);
nor U8797 (N_8797,N_5356,N_5943);
nor U8798 (N_8798,N_5702,N_5112);
nand U8799 (N_8799,N_4628,N_5129);
nand U8800 (N_8800,N_3037,N_4572);
nand U8801 (N_8801,N_4568,N_4139);
and U8802 (N_8802,N_4384,N_5716);
and U8803 (N_8803,N_4353,N_3589);
nand U8804 (N_8804,N_5616,N_3429);
and U8805 (N_8805,N_4552,N_3013);
and U8806 (N_8806,N_5559,N_4851);
nor U8807 (N_8807,N_4781,N_3440);
nor U8808 (N_8808,N_4275,N_4580);
nor U8809 (N_8809,N_3673,N_3527);
and U8810 (N_8810,N_4490,N_5979);
nand U8811 (N_8811,N_4293,N_5132);
nor U8812 (N_8812,N_4300,N_4134);
and U8813 (N_8813,N_5082,N_3105);
nor U8814 (N_8814,N_5618,N_5848);
nand U8815 (N_8815,N_4385,N_5054);
or U8816 (N_8816,N_5524,N_4043);
nand U8817 (N_8817,N_5889,N_4417);
nand U8818 (N_8818,N_5272,N_4044);
xor U8819 (N_8819,N_5024,N_4038);
nand U8820 (N_8820,N_5479,N_3144);
and U8821 (N_8821,N_5881,N_3219);
nand U8822 (N_8822,N_3044,N_5321);
nand U8823 (N_8823,N_5049,N_4190);
nand U8824 (N_8824,N_3961,N_3363);
nand U8825 (N_8825,N_3355,N_3085);
nor U8826 (N_8826,N_4031,N_4340);
and U8827 (N_8827,N_5182,N_4488);
nand U8828 (N_8828,N_3139,N_5247);
and U8829 (N_8829,N_5036,N_5340);
or U8830 (N_8830,N_3570,N_4869);
nor U8831 (N_8831,N_4323,N_5432);
nor U8832 (N_8832,N_4610,N_4960);
nand U8833 (N_8833,N_4220,N_4179);
nand U8834 (N_8834,N_4798,N_5040);
nor U8835 (N_8835,N_4126,N_5582);
nand U8836 (N_8836,N_5670,N_4257);
or U8837 (N_8837,N_4381,N_4778);
or U8838 (N_8838,N_4561,N_4234);
and U8839 (N_8839,N_4430,N_3069);
xor U8840 (N_8840,N_5567,N_3123);
nor U8841 (N_8841,N_5394,N_3115);
nand U8842 (N_8842,N_5868,N_5543);
and U8843 (N_8843,N_3965,N_3025);
nor U8844 (N_8844,N_5780,N_4375);
nor U8845 (N_8845,N_4546,N_3449);
and U8846 (N_8846,N_4515,N_3869);
or U8847 (N_8847,N_5757,N_4564);
nor U8848 (N_8848,N_3076,N_3895);
nand U8849 (N_8849,N_3633,N_4291);
nor U8850 (N_8850,N_4585,N_5582);
nand U8851 (N_8851,N_5993,N_4119);
nand U8852 (N_8852,N_5522,N_3519);
and U8853 (N_8853,N_4814,N_5454);
and U8854 (N_8854,N_3346,N_5085);
or U8855 (N_8855,N_5171,N_5950);
nor U8856 (N_8856,N_3636,N_3856);
nor U8857 (N_8857,N_5405,N_3453);
nand U8858 (N_8858,N_4501,N_3965);
nor U8859 (N_8859,N_3868,N_3335);
nand U8860 (N_8860,N_4743,N_4899);
nand U8861 (N_8861,N_3820,N_4040);
nand U8862 (N_8862,N_4641,N_4417);
nand U8863 (N_8863,N_4463,N_5861);
nor U8864 (N_8864,N_3769,N_5859);
nor U8865 (N_8865,N_3043,N_5146);
nand U8866 (N_8866,N_3849,N_4346);
and U8867 (N_8867,N_3729,N_3085);
nand U8868 (N_8868,N_3143,N_5758);
nand U8869 (N_8869,N_5710,N_4931);
nor U8870 (N_8870,N_3606,N_5651);
nor U8871 (N_8871,N_3732,N_3979);
and U8872 (N_8872,N_4703,N_5470);
nor U8873 (N_8873,N_4420,N_3743);
and U8874 (N_8874,N_3978,N_5446);
and U8875 (N_8875,N_4756,N_4243);
or U8876 (N_8876,N_4657,N_4956);
nand U8877 (N_8877,N_3436,N_4548);
and U8878 (N_8878,N_5898,N_4957);
and U8879 (N_8879,N_4382,N_5770);
nor U8880 (N_8880,N_5637,N_5050);
nor U8881 (N_8881,N_3017,N_3427);
nor U8882 (N_8882,N_5353,N_3073);
nand U8883 (N_8883,N_4221,N_4370);
nand U8884 (N_8884,N_5558,N_3974);
or U8885 (N_8885,N_4991,N_5238);
or U8886 (N_8886,N_4277,N_4187);
nor U8887 (N_8887,N_3980,N_4386);
nand U8888 (N_8888,N_5757,N_5305);
nand U8889 (N_8889,N_5494,N_4659);
nand U8890 (N_8890,N_3101,N_3032);
or U8891 (N_8891,N_4089,N_5823);
nor U8892 (N_8892,N_4165,N_5325);
nand U8893 (N_8893,N_3017,N_4107);
nand U8894 (N_8894,N_5105,N_3464);
nand U8895 (N_8895,N_5247,N_3531);
or U8896 (N_8896,N_5619,N_4886);
nand U8897 (N_8897,N_3579,N_4165);
or U8898 (N_8898,N_5937,N_3319);
nand U8899 (N_8899,N_5665,N_5433);
nand U8900 (N_8900,N_3155,N_5077);
or U8901 (N_8901,N_4614,N_4634);
and U8902 (N_8902,N_3158,N_5922);
nor U8903 (N_8903,N_4828,N_4870);
nand U8904 (N_8904,N_4985,N_5828);
nand U8905 (N_8905,N_5967,N_4914);
nor U8906 (N_8906,N_4030,N_3802);
and U8907 (N_8907,N_3070,N_3636);
nor U8908 (N_8908,N_4475,N_4340);
and U8909 (N_8909,N_4779,N_3797);
nand U8910 (N_8910,N_4133,N_5392);
nor U8911 (N_8911,N_4432,N_4646);
and U8912 (N_8912,N_5370,N_4347);
nand U8913 (N_8913,N_3424,N_4481);
and U8914 (N_8914,N_3101,N_5059);
and U8915 (N_8915,N_5484,N_3934);
and U8916 (N_8916,N_4846,N_5404);
and U8917 (N_8917,N_4128,N_4872);
nand U8918 (N_8918,N_5351,N_4421);
and U8919 (N_8919,N_5521,N_5166);
nand U8920 (N_8920,N_5182,N_5163);
nor U8921 (N_8921,N_3764,N_3823);
nand U8922 (N_8922,N_4086,N_5205);
nand U8923 (N_8923,N_4139,N_4227);
nor U8924 (N_8924,N_4654,N_4046);
and U8925 (N_8925,N_4252,N_5184);
nand U8926 (N_8926,N_5517,N_4226);
or U8927 (N_8927,N_5032,N_3003);
nand U8928 (N_8928,N_3524,N_4465);
or U8929 (N_8929,N_3511,N_5710);
or U8930 (N_8930,N_3774,N_4472);
and U8931 (N_8931,N_4753,N_3689);
xnor U8932 (N_8932,N_4400,N_4216);
or U8933 (N_8933,N_4450,N_3169);
nand U8934 (N_8934,N_3740,N_4867);
and U8935 (N_8935,N_3221,N_3419);
xor U8936 (N_8936,N_5766,N_5325);
and U8937 (N_8937,N_5963,N_3073);
or U8938 (N_8938,N_4559,N_5239);
nor U8939 (N_8939,N_5091,N_3135);
nand U8940 (N_8940,N_5499,N_5392);
nor U8941 (N_8941,N_4221,N_5948);
and U8942 (N_8942,N_5815,N_5011);
nor U8943 (N_8943,N_3957,N_5238);
nand U8944 (N_8944,N_3271,N_3606);
and U8945 (N_8945,N_5419,N_5363);
nand U8946 (N_8946,N_5890,N_3993);
or U8947 (N_8947,N_5828,N_4507);
or U8948 (N_8948,N_5501,N_4364);
or U8949 (N_8949,N_3682,N_4014);
nor U8950 (N_8950,N_4603,N_3011);
nor U8951 (N_8951,N_4397,N_5877);
and U8952 (N_8952,N_5967,N_4968);
nand U8953 (N_8953,N_4834,N_3843);
nand U8954 (N_8954,N_5388,N_5259);
and U8955 (N_8955,N_5592,N_3047);
nand U8956 (N_8956,N_3163,N_5560);
and U8957 (N_8957,N_3094,N_3031);
nand U8958 (N_8958,N_3301,N_5769);
or U8959 (N_8959,N_3398,N_4681);
or U8960 (N_8960,N_3276,N_3825);
nand U8961 (N_8961,N_5661,N_5004);
and U8962 (N_8962,N_4298,N_4345);
and U8963 (N_8963,N_3072,N_3514);
nor U8964 (N_8964,N_3395,N_5821);
nor U8965 (N_8965,N_3966,N_4804);
nand U8966 (N_8966,N_4921,N_4138);
nor U8967 (N_8967,N_4682,N_5747);
nor U8968 (N_8968,N_4588,N_5797);
nor U8969 (N_8969,N_3129,N_3908);
nand U8970 (N_8970,N_4232,N_4238);
or U8971 (N_8971,N_4773,N_3851);
nand U8972 (N_8972,N_5875,N_4364);
nand U8973 (N_8973,N_4644,N_4179);
xnor U8974 (N_8974,N_3549,N_5351);
and U8975 (N_8975,N_4298,N_5016);
xnor U8976 (N_8976,N_3911,N_3662);
or U8977 (N_8977,N_5416,N_5758);
nor U8978 (N_8978,N_4934,N_5239);
or U8979 (N_8979,N_3038,N_5149);
and U8980 (N_8980,N_3761,N_5712);
and U8981 (N_8981,N_3726,N_3560);
nand U8982 (N_8982,N_5048,N_5114);
nor U8983 (N_8983,N_3021,N_4493);
nand U8984 (N_8984,N_5427,N_4199);
nor U8985 (N_8985,N_3612,N_5872);
and U8986 (N_8986,N_4917,N_5943);
or U8987 (N_8987,N_3538,N_3993);
nand U8988 (N_8988,N_3542,N_5209);
or U8989 (N_8989,N_5110,N_4506);
and U8990 (N_8990,N_3154,N_3067);
nand U8991 (N_8991,N_3869,N_3748);
nand U8992 (N_8992,N_4335,N_5828);
and U8993 (N_8993,N_3179,N_3041);
nand U8994 (N_8994,N_3445,N_4063);
and U8995 (N_8995,N_4251,N_4234);
nor U8996 (N_8996,N_3324,N_3179);
and U8997 (N_8997,N_3423,N_5610);
nand U8998 (N_8998,N_4120,N_5631);
and U8999 (N_8999,N_4695,N_4591);
and U9000 (N_9000,N_6074,N_6449);
or U9001 (N_9001,N_8638,N_6833);
or U9002 (N_9002,N_6171,N_8322);
nor U9003 (N_9003,N_8391,N_7755);
nand U9004 (N_9004,N_7784,N_7385);
nor U9005 (N_9005,N_8127,N_6462);
and U9006 (N_9006,N_6821,N_6489);
nor U9007 (N_9007,N_8728,N_7192);
nor U9008 (N_9008,N_6593,N_6009);
nor U9009 (N_9009,N_6406,N_7248);
nor U9010 (N_9010,N_6674,N_6215);
or U9011 (N_9011,N_8982,N_8546);
nor U9012 (N_9012,N_7509,N_7383);
nand U9013 (N_9013,N_8251,N_6638);
nand U9014 (N_9014,N_6338,N_6668);
nor U9015 (N_9015,N_6071,N_8755);
and U9016 (N_9016,N_6120,N_7963);
or U9017 (N_9017,N_7149,N_8571);
and U9018 (N_9018,N_8059,N_8511);
or U9019 (N_9019,N_8049,N_6032);
nand U9020 (N_9020,N_7614,N_6095);
or U9021 (N_9021,N_7982,N_8459);
and U9022 (N_9022,N_6587,N_6892);
nor U9023 (N_9023,N_6970,N_7098);
nor U9024 (N_9024,N_6619,N_6244);
nand U9025 (N_9025,N_6793,N_6503);
and U9026 (N_9026,N_6553,N_8815);
nor U9027 (N_9027,N_7018,N_6877);
and U9028 (N_9028,N_8502,N_7631);
xnor U9029 (N_9029,N_8592,N_7618);
nor U9030 (N_9030,N_6866,N_7245);
nor U9031 (N_9031,N_6394,N_8804);
or U9032 (N_9032,N_6349,N_6600);
nand U9033 (N_9033,N_7589,N_7605);
nor U9034 (N_9034,N_6034,N_7947);
xor U9035 (N_9035,N_8715,N_7859);
or U9036 (N_9036,N_6015,N_7325);
nor U9037 (N_9037,N_7587,N_6166);
or U9038 (N_9038,N_8359,N_7062);
xor U9039 (N_9039,N_8560,N_7709);
and U9040 (N_9040,N_8368,N_6792);
and U9041 (N_9041,N_6673,N_7979);
nor U9042 (N_9042,N_7918,N_8138);
nand U9043 (N_9043,N_6969,N_8435);
nand U9044 (N_9044,N_7370,N_7592);
and U9045 (N_9045,N_8051,N_8438);
and U9046 (N_9046,N_8526,N_7850);
nor U9047 (N_9047,N_8772,N_8885);
and U9048 (N_9048,N_7070,N_8031);
or U9049 (N_9049,N_7422,N_6057);
nand U9050 (N_9050,N_7120,N_6750);
nand U9051 (N_9051,N_6301,N_8298);
nor U9052 (N_9052,N_6158,N_7684);
or U9053 (N_9053,N_8266,N_7968);
nor U9054 (N_9054,N_8242,N_8426);
nor U9055 (N_9055,N_8413,N_6966);
or U9056 (N_9056,N_8588,N_6791);
xnor U9057 (N_9057,N_7505,N_7643);
nand U9058 (N_9058,N_7522,N_8597);
nand U9059 (N_9059,N_7271,N_6558);
or U9060 (N_9060,N_7392,N_8479);
nand U9061 (N_9061,N_6569,N_7057);
nor U9062 (N_9062,N_8997,N_7000);
or U9063 (N_9063,N_7717,N_8768);
and U9064 (N_9064,N_7626,N_6498);
or U9065 (N_9065,N_7822,N_7699);
and U9066 (N_9066,N_8725,N_6919);
nor U9067 (N_9067,N_6096,N_6081);
nor U9068 (N_9068,N_8183,N_6716);
or U9069 (N_9069,N_6367,N_8732);
nor U9070 (N_9070,N_7294,N_8122);
and U9071 (N_9071,N_7519,N_6997);
nand U9072 (N_9072,N_6828,N_8893);
and U9073 (N_9073,N_6205,N_6423);
xnor U9074 (N_9074,N_6521,N_7367);
or U9075 (N_9075,N_8551,N_8157);
and U9076 (N_9076,N_7609,N_8965);
and U9077 (N_9077,N_8939,N_6139);
and U9078 (N_9078,N_6764,N_7082);
nor U9079 (N_9079,N_8108,N_6108);
nor U9080 (N_9080,N_6143,N_8954);
nand U9081 (N_9081,N_7576,N_7697);
or U9082 (N_9082,N_8678,N_6141);
and U9083 (N_9083,N_6512,N_8996);
nor U9084 (N_9084,N_7913,N_8080);
nor U9085 (N_9085,N_6159,N_7242);
xnor U9086 (N_9086,N_6537,N_8581);
nor U9087 (N_9087,N_7443,N_8495);
nor U9088 (N_9088,N_6613,N_6805);
or U9089 (N_9089,N_7147,N_6956);
nand U9090 (N_9090,N_6777,N_7845);
nor U9091 (N_9091,N_7164,N_7286);
nor U9092 (N_9092,N_6534,N_6149);
nor U9093 (N_9093,N_7063,N_6766);
or U9094 (N_9094,N_7529,N_6293);
nor U9095 (N_9095,N_7226,N_7312);
nand U9096 (N_9096,N_8473,N_8855);
nand U9097 (N_9097,N_8660,N_6295);
or U9098 (N_9098,N_6785,N_8057);
or U9099 (N_9099,N_8883,N_7518);
and U9100 (N_9100,N_6984,N_8914);
nand U9101 (N_9101,N_6263,N_8096);
or U9102 (N_9102,N_7711,N_7467);
nor U9103 (N_9103,N_8602,N_7438);
or U9104 (N_9104,N_6098,N_7897);
nand U9105 (N_9105,N_7673,N_8116);
nor U9106 (N_9106,N_6645,N_8789);
nand U9107 (N_9107,N_7616,N_7334);
xnor U9108 (N_9108,N_8330,N_6599);
nor U9109 (N_9109,N_7788,N_6637);
and U9110 (N_9110,N_8155,N_8380);
or U9111 (N_9111,N_8625,N_7282);
nor U9112 (N_9112,N_6376,N_8288);
or U9113 (N_9113,N_7702,N_7409);
nand U9114 (N_9114,N_6331,N_8751);
nand U9115 (N_9115,N_8469,N_7310);
and U9116 (N_9116,N_6632,N_8184);
or U9117 (N_9117,N_7730,N_7005);
nand U9118 (N_9118,N_6216,N_6085);
nor U9119 (N_9119,N_7515,N_6588);
nor U9120 (N_9120,N_7229,N_8877);
nand U9121 (N_9121,N_6891,N_6902);
and U9122 (N_9122,N_7278,N_7813);
xnor U9123 (N_9123,N_6398,N_7588);
nand U9124 (N_9124,N_6383,N_6621);
nand U9125 (N_9125,N_7314,N_7181);
or U9126 (N_9126,N_8753,N_6905);
and U9127 (N_9127,N_8670,N_7414);
or U9128 (N_9128,N_8820,N_8448);
nand U9129 (N_9129,N_7346,N_8270);
nand U9130 (N_9130,N_8975,N_6439);
nor U9131 (N_9131,N_7578,N_8962);
and U9132 (N_9132,N_6304,N_7376);
or U9133 (N_9133,N_7874,N_6958);
nand U9134 (N_9134,N_8112,N_6385);
or U9135 (N_9135,N_7397,N_7797);
and U9136 (N_9136,N_8240,N_7944);
and U9137 (N_9137,N_7139,N_6242);
and U9138 (N_9138,N_8527,N_7061);
nand U9139 (N_9139,N_8609,N_7764);
or U9140 (N_9140,N_7273,N_8023);
and U9141 (N_9141,N_8803,N_8689);
or U9142 (N_9142,N_8523,N_7115);
and U9143 (N_9143,N_7929,N_8197);
and U9144 (N_9144,N_7465,N_7773);
and U9145 (N_9145,N_6035,N_8770);
and U9146 (N_9146,N_7761,N_7378);
and U9147 (N_9147,N_8690,N_7633);
nand U9148 (N_9148,N_7598,N_8009);
and U9149 (N_9149,N_8462,N_7805);
nor U9150 (N_9150,N_6745,N_8243);
nand U9151 (N_9151,N_8465,N_6411);
nand U9152 (N_9152,N_7332,N_8538);
or U9153 (N_9153,N_7321,N_7583);
nand U9154 (N_9154,N_7958,N_7928);
or U9155 (N_9155,N_6430,N_7856);
and U9156 (N_9156,N_8757,N_8830);
and U9157 (N_9157,N_6758,N_7050);
xnor U9158 (N_9158,N_7710,N_8907);
or U9159 (N_9159,N_6709,N_7683);
or U9160 (N_9160,N_6723,N_6202);
nand U9161 (N_9161,N_6756,N_8904);
or U9162 (N_9162,N_7669,N_8507);
nor U9163 (N_9163,N_6072,N_8860);
nand U9164 (N_9164,N_8695,N_7153);
and U9165 (N_9165,N_8151,N_6451);
nand U9166 (N_9166,N_7379,N_8159);
nor U9167 (N_9167,N_6843,N_8759);
nand U9168 (N_9168,N_6841,N_8515);
and U9169 (N_9169,N_6461,N_8875);
or U9170 (N_9170,N_8482,N_8084);
or U9171 (N_9171,N_7328,N_6618);
nand U9172 (N_9172,N_7503,N_7652);
nand U9173 (N_9173,N_8774,N_6237);
nor U9174 (N_9174,N_6675,N_6965);
and U9175 (N_9175,N_6884,N_7624);
and U9176 (N_9176,N_8230,N_6351);
nand U9177 (N_9177,N_6812,N_8760);
nor U9178 (N_9178,N_7645,N_7860);
and U9179 (N_9179,N_8795,N_8248);
xor U9180 (N_9180,N_7969,N_6784);
and U9181 (N_9181,N_6872,N_6604);
nand U9182 (N_9182,N_8231,N_6657);
or U9183 (N_9183,N_6934,N_7794);
nand U9184 (N_9184,N_7218,N_6715);
and U9185 (N_9185,N_6686,N_7069);
xnor U9186 (N_9186,N_8852,N_6084);
and U9187 (N_9187,N_8345,N_7081);
or U9188 (N_9188,N_7851,N_7439);
nand U9189 (N_9189,N_7582,N_6525);
or U9190 (N_9190,N_6809,N_7787);
and U9191 (N_9191,N_6146,N_8333);
nor U9192 (N_9192,N_7132,N_6772);
nor U9193 (N_9193,N_8843,N_6518);
or U9194 (N_9194,N_6730,N_7146);
and U9195 (N_9195,N_8662,N_6798);
nand U9196 (N_9196,N_8436,N_6420);
and U9197 (N_9197,N_6527,N_8898);
nand U9198 (N_9198,N_8086,N_7125);
or U9199 (N_9199,N_7203,N_8525);
nand U9200 (N_9200,N_7361,N_7572);
or U9201 (N_9201,N_6614,N_8844);
nand U9202 (N_9202,N_6670,N_6991);
and U9203 (N_9203,N_8208,N_7932);
nor U9204 (N_9204,N_7469,N_8015);
nor U9205 (N_9205,N_8134,N_6818);
and U9206 (N_9206,N_6950,N_7237);
nand U9207 (N_9207,N_8748,N_7573);
xnor U9208 (N_9208,N_7309,N_8309);
or U9209 (N_9209,N_8563,N_6387);
nor U9210 (N_9210,N_6200,N_6029);
nor U9211 (N_9211,N_6561,N_6460);
or U9212 (N_9212,N_7627,N_8763);
nor U9213 (N_9213,N_6729,N_7528);
or U9214 (N_9214,N_6168,N_8220);
nand U9215 (N_9215,N_8120,N_7388);
and U9216 (N_9216,N_7756,N_7009);
nand U9217 (N_9217,N_6667,N_6836);
nor U9218 (N_9218,N_6397,N_8617);
nand U9219 (N_9219,N_6033,N_8033);
or U9220 (N_9220,N_6820,N_8456);
or U9221 (N_9221,N_6539,N_6025);
and U9222 (N_9222,N_8600,N_7954);
or U9223 (N_9223,N_6664,N_8857);
nor U9224 (N_9224,N_6261,N_8547);
or U9225 (N_9225,N_8932,N_7844);
nand U9226 (N_9226,N_6834,N_7360);
nor U9227 (N_9227,N_8257,N_6265);
and U9228 (N_9228,N_6290,N_7010);
nand U9229 (N_9229,N_6916,N_8468);
or U9230 (N_9230,N_7180,N_7306);
nand U9231 (N_9231,N_7548,N_8191);
nand U9232 (N_9232,N_7060,N_6307);
or U9233 (N_9233,N_8392,N_7092);
nand U9234 (N_9234,N_8655,N_6232);
or U9235 (N_9235,N_8668,N_7274);
nor U9236 (N_9236,N_6344,N_6038);
nor U9237 (N_9237,N_8953,N_7540);
or U9238 (N_9238,N_8708,N_8776);
and U9239 (N_9239,N_7289,N_6363);
or U9240 (N_9240,N_6191,N_7891);
or U9241 (N_9241,N_7987,N_7925);
nor U9242 (N_9242,N_8420,N_7076);
and U9243 (N_9243,N_8219,N_8692);
or U9244 (N_9244,N_7819,N_6783);
and U9245 (N_9245,N_7601,N_6324);
nand U9246 (N_9246,N_7671,N_7089);
or U9247 (N_9247,N_7163,N_6907);
nor U9248 (N_9248,N_6125,N_6375);
nor U9249 (N_9249,N_7110,N_8299);
xnor U9250 (N_9250,N_7570,N_6343);
or U9251 (N_9251,N_7389,N_7425);
and U9252 (N_9252,N_8428,N_6332);
nor U9253 (N_9253,N_6138,N_6094);
nor U9254 (N_9254,N_8529,N_7738);
nand U9255 (N_9255,N_8048,N_8360);
nand U9256 (N_9256,N_6762,N_8376);
nand U9257 (N_9257,N_8401,N_7489);
and U9258 (N_9258,N_7099,N_6887);
or U9259 (N_9259,N_7140,N_7073);
nor U9260 (N_9260,N_7222,N_8362);
nor U9261 (N_9261,N_6277,N_8816);
nor U9262 (N_9262,N_6540,N_8902);
and U9263 (N_9263,N_8577,N_7508);
nand U9264 (N_9264,N_7701,N_8210);
and U9265 (N_9265,N_7604,N_7637);
nand U9266 (N_9266,N_8200,N_6157);
and U9267 (N_9267,N_8653,N_7001);
and U9268 (N_9268,N_8659,N_6359);
and U9269 (N_9269,N_8147,N_6677);
or U9270 (N_9270,N_8038,N_6366);
and U9271 (N_9271,N_8794,N_6628);
or U9272 (N_9272,N_8273,N_8342);
nand U9273 (N_9273,N_6052,N_8195);
nand U9274 (N_9274,N_7243,N_7571);
nor U9275 (N_9275,N_7088,N_7101);
and U9276 (N_9276,N_7384,N_6752);
nand U9277 (N_9277,N_7718,N_7511);
or U9278 (N_9278,N_8223,N_7326);
and U9279 (N_9279,N_8859,N_8111);
nand U9280 (N_9280,N_6271,N_6152);
and U9281 (N_9281,N_6704,N_6162);
or U9282 (N_9282,N_6878,N_8260);
and U9283 (N_9283,N_7833,N_8556);
nor U9284 (N_9284,N_8161,N_7715);
nor U9285 (N_9285,N_6725,N_6601);
or U9286 (N_9286,N_8204,N_7246);
or U9287 (N_9287,N_7525,N_7586);
and U9288 (N_9288,N_7569,N_7602);
and U9289 (N_9289,N_7330,N_8036);
or U9290 (N_9290,N_7757,N_7214);
and U9291 (N_9291,N_8186,N_6584);
or U9292 (N_9292,N_8979,N_8865);
nor U9293 (N_9293,N_8265,N_7369);
nor U9294 (N_9294,N_8381,N_6814);
nor U9295 (N_9295,N_7364,N_7220);
or U9296 (N_9296,N_7216,N_8306);
nor U9297 (N_9297,N_8218,N_6708);
and U9298 (N_9298,N_8056,N_7816);
or U9299 (N_9299,N_8909,N_7014);
and U9300 (N_9300,N_7554,N_8641);
or U9301 (N_9301,N_7279,N_8619);
nor U9302 (N_9302,N_6165,N_7667);
and U9303 (N_9303,N_8156,N_6838);
or U9304 (N_9304,N_7723,N_8199);
nand U9305 (N_9305,N_7191,N_6135);
and U9306 (N_9306,N_8267,N_6867);
nand U9307 (N_9307,N_6083,N_7473);
and U9308 (N_9308,N_7906,N_7724);
or U9309 (N_9309,N_6633,N_6296);
and U9310 (N_9310,N_6482,N_7536);
or U9311 (N_9311,N_7961,N_6594);
nor U9312 (N_9312,N_7353,N_6949);
nor U9313 (N_9313,N_8178,N_6233);
and U9314 (N_9314,N_8943,N_6697);
or U9315 (N_9315,N_6921,N_7029);
and U9316 (N_9316,N_8371,N_7974);
nor U9317 (N_9317,N_7753,N_7148);
or U9318 (N_9318,N_6655,N_7762);
nor U9319 (N_9319,N_7510,N_7656);
nor U9320 (N_9320,N_6678,N_8312);
nand U9321 (N_9321,N_8882,N_8945);
and U9322 (N_9322,N_8058,N_8269);
nor U9323 (N_9323,N_6235,N_6079);
or U9324 (N_9324,N_6473,N_7750);
nor U9325 (N_9325,N_8007,N_8226);
nand U9326 (N_9326,N_7240,N_7707);
or U9327 (N_9327,N_6030,N_7333);
nand U9328 (N_9328,N_7786,N_6370);
nor U9329 (N_9329,N_8378,N_8082);
and U9330 (N_9330,N_8478,N_6974);
or U9331 (N_9331,N_6505,N_6371);
and U9332 (N_9332,N_7054,N_6199);
nor U9333 (N_9333,N_6087,N_8864);
nand U9334 (N_9334,N_6517,N_8951);
or U9335 (N_9335,N_6542,N_8940);
and U9336 (N_9336,N_6182,N_6802);
nor U9337 (N_9337,N_8418,N_8193);
and U9338 (N_9338,N_6622,N_6778);
nand U9339 (N_9339,N_7043,N_8704);
or U9340 (N_9340,N_7032,N_6231);
nor U9341 (N_9341,N_6024,N_6495);
nor U9342 (N_9342,N_7477,N_6070);
nand U9343 (N_9343,N_8919,N_7183);
and U9344 (N_9344,N_7682,N_7990);
or U9345 (N_9345,N_8450,N_7698);
or U9346 (N_9346,N_6787,N_6687);
nor U9347 (N_9347,N_8969,N_7112);
and U9348 (N_9348,N_6133,N_7597);
or U9349 (N_9349,N_8106,N_8908);
or U9350 (N_9350,N_8044,N_7623);
or U9351 (N_9351,N_8358,N_6454);
or U9352 (N_9352,N_6544,N_6946);
nor U9353 (N_9353,N_8061,N_8315);
or U9354 (N_9354,N_7027,N_8812);
and U9355 (N_9355,N_8966,N_8881);
and U9356 (N_9356,N_8363,N_8314);
nor U9357 (N_9357,N_8476,N_6190);
nand U9358 (N_9358,N_7461,N_6858);
and U9359 (N_9359,N_7094,N_8093);
nand U9360 (N_9360,N_7559,N_6894);
and U9361 (N_9361,N_7065,N_6873);
nor U9362 (N_9362,N_6514,N_8915);
nand U9363 (N_9363,N_8873,N_7517);
or U9364 (N_9364,N_6502,N_7311);
nand U9365 (N_9365,N_8524,N_6167);
nand U9366 (N_9366,N_7350,N_6917);
and U9367 (N_9367,N_6480,N_6719);
nand U9368 (N_9368,N_8397,N_7765);
nor U9369 (N_9369,N_6585,N_6443);
nor U9370 (N_9370,N_6695,N_8618);
nand U9371 (N_9371,N_6744,N_6666);
or U9372 (N_9372,N_8762,N_8206);
nor U9373 (N_9373,N_6499,N_8612);
and U9374 (N_9374,N_7319,N_7790);
xor U9375 (N_9375,N_6876,N_7662);
or U9376 (N_9376,N_6901,N_6530);
nor U9377 (N_9377,N_8452,N_6257);
or U9378 (N_9378,N_8006,N_6767);
nor U9379 (N_9379,N_8451,N_6132);
nor U9380 (N_9380,N_6546,N_7173);
or U9381 (N_9381,N_7830,N_8797);
nand U9382 (N_9382,N_6204,N_8846);
nand U9383 (N_9383,N_8946,N_7038);
nor U9384 (N_9384,N_6640,N_7351);
nor U9385 (N_9385,N_7408,N_8025);
or U9386 (N_9386,N_8172,N_8721);
nor U9387 (N_9387,N_6849,N_7455);
nand U9388 (N_9388,N_7087,N_8531);
nor U9389 (N_9389,N_8717,N_8549);
nor U9390 (N_9390,N_8090,N_8694);
nand U9391 (N_9391,N_7871,N_8425);
nor U9392 (N_9392,N_8722,N_8483);
nand U9393 (N_9393,N_7541,N_6911);
nand U9394 (N_9394,N_6826,N_7903);
and U9395 (N_9395,N_7551,N_7391);
nand U9396 (N_9396,N_8500,N_6951);
and U9397 (N_9397,N_7375,N_7459);
nor U9398 (N_9398,N_7064,N_6283);
nand U9399 (N_9399,N_7211,N_6000);
and U9400 (N_9400,N_7747,N_8575);
nor U9401 (N_9401,N_7934,N_6415);
nor U9402 (N_9402,N_7372,N_8377);
or U9403 (N_9403,N_8424,N_8505);
nand U9404 (N_9404,N_8880,N_8684);
or U9405 (N_9405,N_7013,N_7468);
nand U9406 (N_9406,N_8598,N_6662);
and U9407 (N_9407,N_6591,N_8836);
nand U9408 (N_9408,N_6732,N_7972);
xnor U9409 (N_9409,N_8075,N_8020);
and U9410 (N_9410,N_7782,N_8289);
and U9411 (N_9411,N_7911,N_7412);
nand U9412 (N_9412,N_8104,N_6427);
and U9413 (N_9413,N_6998,N_6580);
and U9414 (N_9414,N_7653,N_8842);
and U9415 (N_9415,N_7262,N_7728);
and U9416 (N_9416,N_6513,N_8792);
and U9417 (N_9417,N_7909,N_7985);
and U9418 (N_9418,N_7654,N_7268);
and U9419 (N_9419,N_7686,N_8921);
nand U9420 (N_9420,N_6273,N_6131);
or U9421 (N_9421,N_8393,N_6472);
nor U9422 (N_9422,N_6679,N_8540);
and U9423 (N_9423,N_7866,N_6047);
nand U9424 (N_9424,N_7336,N_8756);
and U9425 (N_9425,N_6317,N_7177);
nand U9426 (N_9426,N_6925,N_7655);
nand U9427 (N_9427,N_7742,N_8109);
and U9428 (N_9428,N_8083,N_6360);
nor U9429 (N_9429,N_6747,N_8594);
nor U9430 (N_9430,N_6623,N_7665);
nand U9431 (N_9431,N_7155,N_6795);
nand U9432 (N_9432,N_8201,N_7386);
or U9433 (N_9433,N_7758,N_7949);
or U9434 (N_9434,N_8286,N_8978);
nor U9435 (N_9435,N_7436,N_8984);
nor U9436 (N_9436,N_6845,N_6455);
or U9437 (N_9437,N_6247,N_8487);
and U9438 (N_9438,N_8329,N_6882);
or U9439 (N_9439,N_7971,N_6631);
or U9440 (N_9440,N_8743,N_6501);
or U9441 (N_9441,N_6642,N_6508);
nand U9442 (N_9442,N_7953,N_7564);
or U9443 (N_9443,N_7066,N_8620);
nand U9444 (N_9444,N_7496,N_8014);
nand U9445 (N_9445,N_8045,N_7740);
and U9446 (N_9446,N_7324,N_7495);
and U9447 (N_9447,N_8073,N_6804);
or U9448 (N_9448,N_8354,N_6090);
xnor U9449 (N_9449,N_6605,N_8861);
or U9450 (N_9450,N_6676,N_6571);
and U9451 (N_9451,N_8422,N_7848);
nand U9452 (N_9452,N_6330,N_8629);
nand U9453 (N_9453,N_6021,N_7283);
nand U9454 (N_9454,N_8383,N_8955);
or U9455 (N_9455,N_6869,N_6938);
and U9456 (N_9456,N_8234,N_8076);
nor U9457 (N_9457,N_6971,N_8528);
or U9458 (N_9458,N_7205,N_7121);
and U9459 (N_9459,N_6401,N_8236);
or U9460 (N_9460,N_7938,N_7122);
or U9461 (N_9461,N_7767,N_6796);
or U9462 (N_9462,N_8307,N_8666);
nand U9463 (N_9463,N_6835,N_6661);
nand U9464 (N_9464,N_7834,N_6746);
nand U9465 (N_9465,N_6189,N_6660);
or U9466 (N_9466,N_7781,N_8189);
nand U9467 (N_9467,N_6178,N_7359);
or U9468 (N_9468,N_8202,N_7644);
or U9469 (N_9469,N_7343,N_6980);
nor U9470 (N_9470,N_7272,N_6961);
or U9471 (N_9471,N_8334,N_6595);
nand U9472 (N_9472,N_7206,N_6365);
nand U9473 (N_9473,N_8222,N_8651);
or U9474 (N_9474,N_6890,N_6348);
nand U9475 (N_9475,N_6909,N_8353);
nand U9476 (N_9476,N_7416,N_8675);
nand U9477 (N_9477,N_8746,N_8323);
or U9478 (N_9478,N_6065,N_7354);
or U9479 (N_9479,N_8379,N_6102);
nor U9480 (N_9480,N_8841,N_7269);
or U9481 (N_9481,N_6560,N_6963);
nand U9482 (N_9482,N_8734,N_7558);
or U9483 (N_9483,N_6759,N_8336);
nand U9484 (N_9484,N_6755,N_6912);
or U9485 (N_9485,N_7424,N_7453);
and U9486 (N_9486,N_8968,N_7862);
nand U9487 (N_9487,N_8512,N_8870);
or U9488 (N_9488,N_6976,N_6054);
nor U9489 (N_9489,N_7713,N_8827);
and U9490 (N_9490,N_7941,N_6811);
or U9491 (N_9491,N_7745,N_8936);
nor U9492 (N_9492,N_7055,N_7997);
nand U9493 (N_9493,N_8355,N_8608);
or U9494 (N_9494,N_8471,N_7708);
or U9495 (N_9495,N_8832,N_7224);
nor U9496 (N_9496,N_7568,N_7280);
nor U9497 (N_9497,N_6983,N_8989);
nand U9498 (N_9498,N_7084,N_8102);
nand U9499 (N_9499,N_6382,N_6148);
nor U9500 (N_9500,N_8510,N_8647);
nand U9501 (N_9501,N_8649,N_8390);
or U9502 (N_9502,N_7366,N_6388);
and U9503 (N_9503,N_7429,N_8153);
nor U9504 (N_9504,N_6346,N_7256);
xor U9505 (N_9505,N_8894,N_7666);
or U9506 (N_9506,N_7821,N_6774);
nand U9507 (N_9507,N_6711,N_8822);
nor U9508 (N_9508,N_6176,N_7401);
and U9509 (N_9509,N_8285,N_6305);
nor U9510 (N_9510,N_8055,N_6868);
nand U9511 (N_9511,N_6886,N_6404);
nor U9512 (N_9512,N_8372,N_6727);
nand U9513 (N_9513,N_6652,N_6684);
or U9514 (N_9514,N_6776,N_7887);
or U9515 (N_9515,N_6438,N_7560);
or U9516 (N_9516,N_7421,N_6328);
or U9517 (N_9517,N_8233,N_7824);
and U9518 (N_9518,N_6060,N_7893);
nand U9519 (N_9519,N_7402,N_8958);
nor U9520 (N_9520,N_8252,N_8905);
xnor U9521 (N_9521,N_7940,N_8673);
nor U9522 (N_9522,N_8778,N_7892);
nor U9523 (N_9523,N_8064,N_6769);
nand U9524 (N_9524,N_7817,N_6292);
and U9525 (N_9525,N_8806,N_8933);
and U9526 (N_9526,N_6369,N_6266);
or U9527 (N_9527,N_6109,N_8530);
or U9528 (N_9528,N_7689,N_8077);
nand U9529 (N_9529,N_7865,N_6405);
nor U9530 (N_9530,N_8925,N_8942);
nand U9531 (N_9531,N_6110,N_8947);
nand U9532 (N_9532,N_6364,N_7323);
or U9533 (N_9533,N_8247,N_6078);
and U9534 (N_9534,N_7877,N_6497);
nand U9535 (N_9535,N_8466,N_7802);
and U9536 (N_9536,N_8626,N_7020);
nand U9537 (N_9537,N_7512,N_7107);
or U9538 (N_9538,N_7239,N_7899);
nor U9539 (N_9539,N_8114,N_7329);
nand U9540 (N_9540,N_8570,N_6915);
nand U9541 (N_9541,N_6634,N_8458);
xor U9542 (N_9542,N_6442,N_6853);
nor U9543 (N_9543,N_6140,N_6245);
nand U9544 (N_9544,N_7233,N_6770);
nor U9545 (N_9545,N_7640,N_8838);
and U9546 (N_9546,N_8475,N_6700);
and U9547 (N_9547,N_6506,N_6753);
or U9548 (N_9548,N_8735,N_6724);
nor U9549 (N_9549,N_6436,N_8654);
nor U9550 (N_9550,N_8423,N_8727);
or U9551 (N_9551,N_8665,N_6280);
nor U9552 (N_9552,N_8493,N_7025);
or U9553 (N_9553,N_8047,N_7493);
nand U9554 (N_9554,N_6865,N_7810);
and U9555 (N_9555,N_7863,N_6113);
nand U9556 (N_9556,N_7317,N_6471);
or U9557 (N_9557,N_8386,N_7658);
and U9558 (N_9558,N_8534,N_7868);
nand U9559 (N_9559,N_8308,N_6465);
and U9560 (N_9560,N_6568,N_8327);
and U9561 (N_9561,N_8485,N_6922);
or U9562 (N_9562,N_8863,N_7625);
nor U9563 (N_9563,N_6183,N_7235);
nand U9564 (N_9564,N_8878,N_8118);
or U9565 (N_9565,N_6748,N_7244);
nand U9566 (N_9566,N_6448,N_6197);
or U9567 (N_9567,N_7413,N_7657);
or U9568 (N_9568,N_6590,N_8325);
or U9569 (N_9569,N_7427,N_8646);
and U9570 (N_9570,N_8621,N_7685);
or U9571 (N_9571,N_7676,N_8399);
and U9572 (N_9572,N_7450,N_6248);
nor U9573 (N_9573,N_8280,N_6392);
nand U9574 (N_9574,N_6421,N_8516);
nor U9575 (N_9575,N_7942,N_6358);
or U9576 (N_9576,N_8113,N_6194);
or U9577 (N_9577,N_8593,N_7875);
nand U9578 (N_9578,N_8761,N_8564);
and U9579 (N_9579,N_6260,N_7035);
or U9580 (N_9580,N_7721,N_8677);
or U9581 (N_9581,N_7002,N_8823);
nand U9582 (N_9582,N_6903,N_6617);
nand U9583 (N_9583,N_7172,N_8352);
or U9584 (N_9584,N_8918,N_7145);
or U9585 (N_9585,N_6011,N_8070);
nand U9586 (N_9586,N_7056,N_8011);
nand U9587 (N_9587,N_7046,N_6829);
or U9588 (N_9588,N_6425,N_8998);
or U9589 (N_9589,N_6088,N_7746);
nor U9590 (N_9590,N_7635,N_6957);
nand U9591 (N_9591,N_7894,N_8503);
and U9592 (N_9592,N_7921,N_8499);
and U9593 (N_9593,N_8171,N_8484);
and U9594 (N_9594,N_8065,N_7607);
or U9595 (N_9595,N_8067,N_7965);
or U9596 (N_9596,N_8636,N_6386);
nand U9597 (N_9597,N_7475,N_8656);
nor U9598 (N_9598,N_7952,N_8085);
nand U9599 (N_9599,N_8930,N_7642);
nor U9600 (N_9600,N_7499,N_7567);
or U9601 (N_9601,N_6302,N_6781);
or U9602 (N_9602,N_6066,N_8562);
or U9603 (N_9603,N_6467,N_6322);
or U9604 (N_9604,N_6020,N_6738);
or U9605 (N_9605,N_8414,N_6410);
nor U9606 (N_9606,N_6847,N_8896);
nor U9607 (N_9607,N_8514,N_6797);
nor U9608 (N_9608,N_7629,N_8099);
nor U9609 (N_9609,N_7458,N_8364);
and U9610 (N_9610,N_8052,N_7776);
nand U9611 (N_9611,N_6046,N_8163);
nor U9612 (N_9612,N_7639,N_6988);
nor U9613 (N_9613,N_6111,N_7189);
or U9614 (N_9614,N_7792,N_8010);
and U9615 (N_9615,N_7371,N_7498);
nor U9616 (N_9616,N_6393,N_7338);
or U9617 (N_9617,N_6967,N_8098);
and U9618 (N_9618,N_7159,N_7470);
or U9619 (N_9619,N_7879,N_6996);
nor U9620 (N_9620,N_8141,N_8634);
and U9621 (N_9621,N_6063,N_8054);
and U9622 (N_9622,N_8501,N_6663);
and U9623 (N_9623,N_6474,N_8884);
nor U9624 (N_9624,N_8000,N_8847);
nand U9625 (N_9625,N_6062,N_8680);
or U9626 (N_9626,N_8635,N_6531);
or U9627 (N_9627,N_7476,N_7610);
and U9628 (N_9628,N_6819,N_7542);
and U9629 (N_9629,N_7889,N_7335);
nor U9630 (N_9630,N_6940,N_6572);
or U9631 (N_9631,N_6879,N_6630);
nor U9632 (N_9632,N_6142,N_6037);
xor U9633 (N_9633,N_6105,N_7307);
nor U9634 (N_9634,N_8985,N_8209);
and U9635 (N_9635,N_7188,N_6672);
nor U9636 (N_9636,N_7133,N_8375);
or U9637 (N_9637,N_6702,N_8693);
nor U9638 (N_9638,N_8739,N_6538);
and U9639 (N_9639,N_8439,N_8582);
nor U9640 (N_9640,N_7275,N_6626);
nor U9641 (N_9641,N_8143,N_6717);
and U9642 (N_9642,N_7768,N_7741);
or U9643 (N_9643,N_7590,N_8624);
and U9644 (N_9644,N_7404,N_6788);
and U9645 (N_9645,N_6377,N_8971);
and U9646 (N_9646,N_8706,N_7044);
and U9647 (N_9647,N_6962,N_8357);
nor U9648 (N_9648,N_7300,N_7727);
nand U9649 (N_9649,N_7134,N_6414);
nand U9650 (N_9650,N_8078,N_8028);
and U9651 (N_9651,N_6432,N_8311);
and U9652 (N_9652,N_6577,N_6089);
and U9653 (N_9653,N_6075,N_7019);
nand U9654 (N_9654,N_8796,N_7530);
and U9655 (N_9655,N_7980,N_7053);
nand U9656 (N_9656,N_8402,N_8198);
and U9657 (N_9657,N_8576,N_8276);
and U9658 (N_9658,N_7483,N_8851);
nor U9659 (N_9659,N_7426,N_7022);
or U9660 (N_9660,N_7759,N_7960);
nand U9661 (N_9661,N_6234,N_8264);
nor U9662 (N_9662,N_6318,N_7632);
nand U9663 (N_9663,N_6192,N_7305);
or U9664 (N_9664,N_6281,N_7197);
nor U9665 (N_9665,N_7532,N_6986);
nand U9666 (N_9666,N_7118,N_7136);
nor U9667 (N_9667,N_8906,N_7111);
or U9668 (N_9668,N_8369,N_7600);
or U9669 (N_9669,N_8291,N_7538);
or U9670 (N_9670,N_7234,N_6127);
nor U9671 (N_9671,N_7168,N_7479);
and U9672 (N_9672,N_6813,N_8173);
or U9673 (N_9673,N_7823,N_8601);
nor U9674 (N_9674,N_6519,N_7585);
or U9675 (N_9675,N_6270,N_7349);
nor U9676 (N_9676,N_8453,N_7930);
nand U9677 (N_9677,N_8454,N_7456);
nor U9678 (N_9678,N_6920,N_6228);
nand U9679 (N_9679,N_8658,N_6264);
or U9680 (N_9680,N_6221,N_8382);
nor U9681 (N_9681,N_8633,N_6705);
or U9682 (N_9682,N_6646,N_8021);
nand U9683 (N_9683,N_6665,N_8868);
and U9684 (N_9684,N_7783,N_6130);
xnor U9685 (N_9685,N_6064,N_8750);
or U9686 (N_9686,N_8818,N_8974);
and U9687 (N_9687,N_6718,N_6579);
nor U9688 (N_9688,N_6464,N_7497);
and U9689 (N_9689,N_6452,N_6567);
or U9690 (N_9690,N_7199,N_8977);
nand U9691 (N_9691,N_6582,N_7668);
and U9692 (N_9692,N_6217,N_6557);
or U9693 (N_9693,N_8229,N_6391);
nand U9694 (N_9694,N_8980,N_7919);
nand U9695 (N_9695,N_7647,N_6556);
nor U9696 (N_9696,N_6353,N_8331);
and U9697 (N_9697,N_6609,N_7190);
nand U9698 (N_9698,N_7574,N_8741);
nand U9699 (N_9699,N_6300,N_8922);
or U9700 (N_9700,N_7085,N_8506);
or U9701 (N_9701,N_7051,N_7341);
nor U9702 (N_9702,N_8272,N_7119);
nor U9703 (N_9703,N_7288,N_7471);
and U9704 (N_9704,N_7238,N_6516);
and U9705 (N_9705,N_7520,N_8071);
and U9706 (N_9706,N_8132,N_6453);
nand U9707 (N_9707,N_8972,N_7799);
and U9708 (N_9708,N_7620,N_7608);
nor U9709 (N_9709,N_7846,N_7484);
nor U9710 (N_9710,N_6990,N_7945);
and U9711 (N_9711,N_7651,N_7796);
and U9712 (N_9712,N_8472,N_8623);
nor U9713 (N_9713,N_6463,N_7179);
nand U9714 (N_9714,N_6698,N_6941);
nand U9715 (N_9715,N_8548,N_8888);
nand U9716 (N_9716,N_6104,N_7621);
nand U9717 (N_9717,N_7225,N_6629);
nor U9718 (N_9718,N_8956,N_8644);
and U9719 (N_9719,N_6888,N_8912);
and U9720 (N_9720,N_7622,N_7261);
or U9721 (N_9721,N_6285,N_7864);
nor U9722 (N_9722,N_8139,N_7544);
or U9723 (N_9723,N_8321,N_6839);
nand U9724 (N_9724,N_8742,N_6541);
nor U9725 (N_9725,N_8565,N_6968);
nor U9726 (N_9726,N_6459,N_6028);
or U9727 (N_9727,N_6824,N_8411);
and U9728 (N_9728,N_6710,N_8738);
and U9729 (N_9729,N_8995,N_6413);
or U9730 (N_9730,N_7599,N_8688);
or U9731 (N_9731,N_6275,N_8959);
nor U9732 (N_9732,N_8164,N_6799);
or U9733 (N_9733,N_7247,N_6241);
nor U9734 (N_9734,N_6859,N_6603);
nor U9735 (N_9735,N_8879,N_7808);
or U9736 (N_9736,N_8853,N_8994);
nand U9737 (N_9737,N_6213,N_7725);
and U9738 (N_9738,N_6615,N_6620);
nor U9739 (N_9739,N_6050,N_7048);
nand U9740 (N_9740,N_8012,N_8615);
and U9741 (N_9741,N_7144,N_7124);
nand U9742 (N_9742,N_6022,N_6483);
nor U9743 (N_9743,N_8347,N_7795);
nand U9744 (N_9744,N_8920,N_7184);
or U9745 (N_9745,N_7252,N_6830);
nand U9746 (N_9746,N_7052,N_6575);
and U9747 (N_9747,N_8926,N_8555);
nand U9748 (N_9748,N_6786,N_6350);
nor U9749 (N_9749,N_6933,N_7837);
and U9750 (N_9750,N_7302,N_6608);
nor U9751 (N_9751,N_6760,N_6053);
nand U9752 (N_9752,N_6975,N_7948);
and U9753 (N_9753,N_7803,N_7719);
nand U9754 (N_9754,N_7417,N_6596);
and U9755 (N_9755,N_7074,N_8340);
or U9756 (N_9756,N_6279,N_6379);
nand U9757 (N_9757,N_8042,N_7908);
nor U9758 (N_9758,N_8319,N_7998);
or U9759 (N_9759,N_7991,N_8101);
and U9760 (N_9760,N_6931,N_6316);
or U9761 (N_9761,N_6691,N_7313);
nor U9762 (N_9762,N_8697,N_7555);
and U9763 (N_9763,N_6832,N_7935);
nor U9764 (N_9764,N_7843,N_6932);
nor U9765 (N_9765,N_8990,N_6278);
nor U9766 (N_9766,N_8814,N_6566);
nor U9767 (N_9767,N_8295,N_8324);
nor U9768 (N_9768,N_8709,N_6509);
and U9769 (N_9769,N_6198,N_7357);
nor U9770 (N_9770,N_6681,N_6536);
or U9771 (N_9771,N_6736,N_6254);
nor U9772 (N_9772,N_6252,N_6606);
and U9773 (N_9773,N_8829,N_7912);
or U9774 (N_9774,N_6511,N_7502);
nand U9775 (N_9775,N_7674,N_7345);
nand U9776 (N_9776,N_6688,N_7752);
or U9777 (N_9777,N_7594,N_8606);
nor U9778 (N_9778,N_8934,N_7126);
nand U9779 (N_9779,N_7196,N_6694);
or U9780 (N_9780,N_7690,N_7348);
nand U9781 (N_9781,N_7575,N_7299);
nand U9782 (N_9782,N_8287,N_8737);
nand U9783 (N_9783,N_7959,N_6689);
nor U9784 (N_9784,N_7251,N_7358);
nor U9785 (N_9785,N_6230,N_8250);
or U9786 (N_9786,N_7318,N_6073);
nor U9787 (N_9787,N_6400,N_6186);
nor U9788 (N_9788,N_8440,N_6340);
nor U9789 (N_9789,N_6311,N_6040);
nor U9790 (N_9790,N_8825,N_8177);
and U9791 (N_9791,N_6308,N_6150);
and U9792 (N_9792,N_6635,N_7630);
or U9793 (N_9793,N_7331,N_8981);
and U9794 (N_9794,N_8019,N_7423);
or U9795 (N_9795,N_6129,N_8497);
or U9796 (N_9796,N_7996,N_8253);
and U9797 (N_9797,N_8712,N_6426);
nand U9798 (N_9798,N_6999,N_8350);
nor U9799 (N_9799,N_6654,N_8237);
and U9800 (N_9800,N_7263,N_8003);
nor U9801 (N_9801,N_7798,N_6528);
nand U9802 (N_9802,N_7664,N_8088);
nand U9803 (N_9803,N_7793,N_6486);
or U9804 (N_9804,N_8572,N_7854);
and U9805 (N_9805,N_8518,N_7552);
nor U9806 (N_9806,N_8463,N_7394);
and U9807 (N_9807,N_6611,N_6936);
nor U9808 (N_9808,N_7705,N_8871);
and U9809 (N_9809,N_8388,N_6701);
or U9810 (N_9810,N_6122,N_8938);
nor U9811 (N_9811,N_6487,N_7104);
and U9812 (N_9812,N_7650,N_8258);
and U9813 (N_9813,N_7936,N_7403);
nand U9814 (N_9814,N_6973,N_6721);
and U9815 (N_9815,N_6180,N_7437);
nand U9816 (N_9816,N_8674,N_8805);
nand U9817 (N_9817,N_8719,N_7420);
nor U9818 (N_9818,N_7754,N_8136);
nand U9819 (N_9819,N_6533,N_7562);
and U9820 (N_9820,N_8987,N_7154);
nand U9821 (N_9821,N_8405,N_7841);
or U9822 (N_9822,N_8119,N_7749);
nor U9823 (N_9823,N_8941,N_6552);
nand U9824 (N_9824,N_8935,N_6352);
and U9825 (N_9825,N_6058,N_7150);
nand U9826 (N_9826,N_7549,N_7999);
or U9827 (N_9827,N_6355,N_6602);
or U9828 (N_9828,N_8215,N_7986);
nor U9829 (N_9829,N_7223,N_7611);
nor U9830 (N_9830,N_7736,N_7442);
nand U9831 (N_9831,N_7152,N_6128);
nand U9832 (N_9832,N_8457,N_7964);
or U9833 (N_9833,N_8261,N_7165);
nor U9834 (N_9834,N_8773,N_8005);
xor U9835 (N_9835,N_7907,N_7812);
nand U9836 (N_9836,N_6526,N_6779);
nand U9837 (N_9837,N_8008,N_6312);
and U9838 (N_9838,N_6156,N_7204);
or U9839 (N_9839,N_7169,N_8211);
and U9840 (N_9840,N_8304,N_7086);
nand U9841 (N_9841,N_7726,N_6207);
or U9842 (N_9842,N_7071,N_7955);
nand U9843 (N_9843,N_8239,N_7956);
or U9844 (N_9844,N_6173,N_6771);
or U9845 (N_9845,N_8389,N_6116);
and U9846 (N_9846,N_8771,N_7151);
nand U9847 (N_9847,N_6831,N_7660);
and U9848 (N_9848,N_7737,N_8683);
or U9849 (N_9849,N_8707,N_8800);
nor U9850 (N_9850,N_8283,N_7902);
nor U9851 (N_9851,N_7208,N_6690);
nor U9852 (N_9852,N_7221,N_7537);
or U9853 (N_9853,N_7857,N_7373);
and U9854 (N_9854,N_6942,N_8026);
xnor U9855 (N_9855,N_8320,N_7451);
nand U9856 (N_9856,N_8179,N_6522);
or U9857 (N_9857,N_8895,N_7933);
nor U9858 (N_9858,N_7596,N_8802);
or U9859 (N_9859,N_6712,N_7462);
or U9860 (N_9860,N_6403,N_7791);
and U9861 (N_9861,N_7067,N_7504);
nor U9862 (N_9862,N_6906,N_8491);
nand U9863 (N_9863,N_8246,N_7962);
nor U9864 (N_9864,N_7751,N_7779);
nand U9865 (N_9865,N_8676,N_6042);
or U9866 (N_9866,N_6856,N_8889);
nor U9867 (N_9867,N_8671,N_6782);
nand U9868 (N_9868,N_8245,N_8274);
nor U9869 (N_9869,N_7265,N_8837);
nand U9870 (N_9870,N_6396,N_7617);
or U9871 (N_9871,N_6825,N_8664);
and U9872 (N_9872,N_6017,N_7083);
and U9873 (N_9873,N_6555,N_8244);
nand U9874 (N_9874,N_6044,N_8282);
nor U9875 (N_9875,N_7143,N_8290);
nand U9876 (N_9876,N_7603,N_6943);
nor U9877 (N_9877,N_8869,N_6315);
nand U9878 (N_9878,N_7881,N_7849);
nor U9879 (N_9879,N_7415,N_7157);
and U9880 (N_9880,N_8607,N_6954);
nor U9881 (N_9881,N_6240,N_8259);
nand U9882 (N_9882,N_8188,N_7876);
and U9883 (N_9883,N_7185,N_7951);
and U9884 (N_9884,N_6549,N_6155);
and U9885 (N_9885,N_8887,N_6447);
and U9886 (N_9886,N_8024,N_6291);
nor U9887 (N_9887,N_6456,N_8344);
or U9888 (N_9888,N_8160,N_8650);
or U9889 (N_9889,N_7011,N_6172);
and U9890 (N_9890,N_7636,N_8744);
and U9891 (N_9891,N_8911,N_8262);
or U9892 (N_9892,N_6987,N_7693);
nand U9893 (N_9893,N_7516,N_6256);
nand U9894 (N_9894,N_8780,N_8190);
nand U9895 (N_9895,N_6177,N_8890);
or U9896 (N_9896,N_6193,N_8303);
or U9897 (N_9897,N_8480,N_8856);
nand U9898 (N_9898,N_7628,N_6218);
and U9899 (N_9899,N_6395,N_8544);
or U9900 (N_9900,N_7615,N_6842);
or U9901 (N_9901,N_6860,N_8481);
nor U9902 (N_9902,N_6823,N_7448);
or U9903 (N_9903,N_6504,N_6754);
or U9904 (N_9904,N_8097,N_8924);
nor U9905 (N_9905,N_7418,N_6806);
nor U9906 (N_9906,N_6201,N_8589);
nor U9907 (N_9907,N_6854,N_6412);
or U9908 (N_9908,N_7920,N_7563);
or U9909 (N_9909,N_7284,N_7463);
nand U9910 (N_9910,N_8637,N_8498);
and U9911 (N_9911,N_8539,N_6515);
nand U9912 (N_9912,N_6713,N_8221);
or U9913 (N_9913,N_8613,N_7474);
nand U9914 (N_9914,N_6012,N_6523);
or U9915 (N_9915,N_8819,N_7780);
nor U9916 (N_9916,N_8667,N_6647);
and U9917 (N_9917,N_7973,N_6124);
nand U9918 (N_9918,N_6069,N_6239);
or U9919 (N_9919,N_8241,N_7826);
or U9920 (N_9920,N_7281,N_6313);
nand U9921 (N_9921,N_8168,N_8567);
xor U9922 (N_9922,N_8228,N_6895);
nor U9923 (N_9923,N_7840,N_7296);
or U9924 (N_9924,N_8949,N_6563);
and U9925 (N_9925,N_8691,N_8128);
or U9926 (N_9926,N_6117,N_8710);
nor U9927 (N_9927,N_8910,N_7452);
or U9928 (N_9928,N_8037,N_7646);
or U9929 (N_9929,N_7444,N_8632);
nand U9930 (N_9930,N_8872,N_7026);
and U9931 (N_9931,N_7801,N_7105);
or U9932 (N_9932,N_7241,N_7387);
nand U9933 (N_9933,N_6203,N_7356);
or U9934 (N_9934,N_7141,N_8212);
and U9935 (N_9935,N_6993,N_6810);
or U9936 (N_9936,N_6573,N_7079);
or U9937 (N_9937,N_6303,N_6319);
or U9938 (N_9938,N_6068,N_6045);
nand U9939 (N_9939,N_7093,N_8752);
nor U9940 (N_9940,N_7774,N_7487);
or U9941 (N_9941,N_7533,N_8135);
or U9942 (N_9942,N_8779,N_7228);
and U9943 (N_9943,N_8950,N_7253);
or U9944 (N_9944,N_7007,N_6524);
nor U9945 (N_9945,N_6294,N_8700);
nand U9946 (N_9946,N_6817,N_8488);
or U9947 (N_9947,N_8016,N_8541);
and U9948 (N_9948,N_6112,N_8022);
nand U9949 (N_9949,N_8574,N_7488);
and U9950 (N_9950,N_7075,N_7017);
nand U9951 (N_9951,N_6535,N_8256);
nand U9952 (N_9952,N_8145,N_6852);
or U9953 (N_9953,N_6749,N_6327);
nor U9954 (N_9954,N_8578,N_8278);
nor U9955 (N_9955,N_6885,N_8227);
or U9956 (N_9956,N_6669,N_7946);
or U9957 (N_9957,N_6883,N_8758);
nand U9958 (N_9958,N_8899,N_8509);
nand U9959 (N_9959,N_7820,N_6003);
and U9960 (N_9960,N_6236,N_8370);
or U9961 (N_9961,N_8409,N_7303);
nand U9962 (N_9962,N_7524,N_8519);
nand U9963 (N_9963,N_7731,N_8142);
and U9964 (N_9964,N_8035,N_8992);
nor U9965 (N_9965,N_7293,N_7440);
nand U9966 (N_9966,N_6179,N_7853);
and U9967 (N_9967,N_8986,N_8374);
nand U9968 (N_9968,N_7814,N_7342);
or U9969 (N_9969,N_6742,N_6431);
or U9970 (N_9970,N_6336,N_7123);
nor U9971 (N_9971,N_7399,N_8777);
nand U9972 (N_9972,N_7036,N_6390);
nand U9973 (N_9973,N_8412,N_6918);
nor U9974 (N_9974,N_7485,N_7700);
nand U9975 (N_9975,N_7267,N_7835);
and U9976 (N_9976,N_7434,N_6298);
nor U9977 (N_9977,N_7984,N_6434);
or U9978 (N_9978,N_7748,N_7285);
nor U9979 (N_9979,N_7838,N_8685);
nor U9980 (N_9980,N_7695,N_7127);
nand U9981 (N_9981,N_8648,N_7789);
nand U9982 (N_9982,N_7449,N_6147);
nor U9983 (N_9983,N_6589,N_8126);
nor U9984 (N_9984,N_7445,N_6607);
or U9985 (N_9985,N_6051,N_7547);
nor U9986 (N_9986,N_6761,N_7040);
or U9987 (N_9987,N_7100,N_7481);
and U9988 (N_9988,N_7250,N_6908);
or U9989 (N_9989,N_8533,N_8470);
nand U9990 (N_9990,N_7068,N_6592);
or U9991 (N_9991,N_6297,N_6658);
nand U9992 (N_9992,N_8596,N_7187);
nor U9993 (N_9993,N_7212,N_7593);
xor U9994 (N_9994,N_7478,N_6496);
and U9995 (N_9995,N_7156,N_7297);
or U9996 (N_9996,N_8365,N_7352);
and U9997 (N_9997,N_6284,N_6481);
nand U9998 (N_9998,N_7039,N_8069);
or U9999 (N_9999,N_7855,N_6653);
or U10000 (N_10000,N_7649,N_7916);
nor U10001 (N_10001,N_7454,N_6576);
or U10002 (N_10002,N_6636,N_6100);
nand U10003 (N_10003,N_6381,N_7322);
nand U10004 (N_10004,N_6944,N_8595);
nor U10005 (N_10005,N_6337,N_8062);
and U10006 (N_10006,N_6299,N_8404);
and U10007 (N_10007,N_8148,N_6259);
and U10008 (N_10008,N_6226,N_6018);
and U10009 (N_10009,N_7460,N_6001);
and U10010 (N_10010,N_7883,N_6310);
or U10011 (N_10011,N_7613,N_6227);
nor U10012 (N_10012,N_8729,N_7320);
nand U10013 (N_10013,N_7291,N_7988);
or U10014 (N_10014,N_8999,N_6016);
nor U10015 (N_10015,N_8810,N_6048);
nand U10016 (N_10016,N_6077,N_8316);
nor U10017 (N_10017,N_6402,N_8296);
nand U10018 (N_10018,N_8263,N_8973);
and U10019 (N_10019,N_6238,N_8271);
nor U10020 (N_10020,N_8929,N_8769);
nand U10021 (N_10021,N_6977,N_8279);
and U10022 (N_10022,N_7207,N_8103);
and U10023 (N_10023,N_6651,N_6743);
nor U10024 (N_10024,N_8723,N_6320);
or U10025 (N_10025,N_6570,N_7008);
nand U10026 (N_10026,N_8801,N_7521);
or U10027 (N_10027,N_7390,N_6650);
nand U10028 (N_10028,N_6004,N_6007);
nor U10029 (N_10029,N_7004,N_7825);
nand U10030 (N_10030,N_7258,N_7130);
nor U10031 (N_10031,N_7937,N_6494);
or U10032 (N_10032,N_7096,N_6790);
nand U10033 (N_10033,N_6361,N_6253);
nand U10034 (N_10034,N_8745,N_8294);
nor U10035 (N_10035,N_7117,N_7870);
nor U10036 (N_10036,N_7393,N_6080);
xor U10037 (N_10037,N_6106,N_8284);
nor U10038 (N_10038,N_7045,N_8736);
nor U10039 (N_10039,N_6101,N_6408);
nand U10040 (N_10040,N_8149,N_6864);
nand U10041 (N_10041,N_7257,N_6446);
and U10042 (N_10042,N_6722,N_7677);
or U10043 (N_10043,N_6445,N_6510);
nor U10044 (N_10044,N_6175,N_8703);
nor U10045 (N_10045,N_6031,N_7772);
nor U10046 (N_10046,N_6092,N_8892);
or U10047 (N_10047,N_8639,N_8661);
or U10048 (N_10048,N_7744,N_7992);
nand U10049 (N_10049,N_7023,N_6728);
nand U10050 (N_10050,N_7049,N_7901);
or U10051 (N_10051,N_6267,N_8952);
nor U10052 (N_10052,N_7514,N_8799);
nor U10053 (N_10053,N_6696,N_7301);
and U10054 (N_10054,N_7255,N_7565);
or U10055 (N_10055,N_7419,N_6529);
nor U10056 (N_10056,N_8764,N_6682);
xor U10057 (N_10057,N_8900,N_8492);
or U10058 (N_10058,N_7337,N_8897);
and U10059 (N_10059,N_7230,N_7435);
and U10060 (N_10060,N_6643,N_6107);
or U10061 (N_10061,N_8150,N_6741);
nand U10062 (N_10062,N_7162,N_8027);
or U10063 (N_10063,N_6897,N_7174);
and U10064 (N_10064,N_8441,N_6659);
nor U10065 (N_10065,N_7720,N_6126);
and U10066 (N_10066,N_7398,N_7202);
nand U10067 (N_10067,N_8477,N_8913);
xor U10068 (N_10068,N_8559,N_8867);
nor U10069 (N_10069,N_6904,N_8105);
or U10070 (N_10070,N_7171,N_8782);
nor U10071 (N_10071,N_6417,N_6641);
or U10072 (N_10072,N_8034,N_8642);
nor U10073 (N_10073,N_6952,N_7818);
nor U10074 (N_10074,N_6181,N_6583);
nor U10075 (N_10075,N_8181,N_7975);
nor U10076 (N_10076,N_6484,N_8419);
nand U10077 (N_10077,N_6734,N_8726);
nand U10078 (N_10078,N_8050,N_7106);
and U10079 (N_10079,N_8766,N_6160);
and U10080 (N_10080,N_8927,N_6008);
nor U10081 (N_10081,N_6212,N_6578);
or U10082 (N_10082,N_7663,N_6161);
nand U10083 (N_10083,N_8845,N_8591);
and U10084 (N_10084,N_6889,N_6979);
nand U10085 (N_10085,N_8385,N_7006);
nand U10086 (N_10086,N_8603,N_6656);
and U10087 (N_10087,N_7766,N_6211);
nor U10088 (N_10088,N_7178,N_7446);
nor U10089 (N_10089,N_8964,N_8249);
and U10090 (N_10090,N_6726,N_6082);
or U10091 (N_10091,N_8948,N_7861);
or U10092 (N_10092,N_7591,N_7734);
and U10093 (N_10093,N_6775,N_6061);
or U10094 (N_10094,N_8580,N_6076);
nand U10095 (N_10095,N_6219,N_6306);
and U10096 (N_10096,N_7777,N_6978);
or U10097 (N_10097,N_7904,N_7103);
nand U10098 (N_10098,N_6773,N_8686);
and U10099 (N_10099,N_7213,N_7910);
nor U10100 (N_10100,N_6170,N_7577);
or U10101 (N_10101,N_8254,N_8698);
or U10102 (N_10102,N_6923,N_6648);
and U10103 (N_10103,N_6268,N_6612);
nor U10104 (N_10104,N_8554,N_6815);
and U10105 (N_10105,N_8702,N_8095);
or U10106 (N_10106,N_7831,N_8281);
and U10107 (N_10107,N_8550,N_8124);
or U10108 (N_10108,N_8348,N_8599);
nand U10109 (N_10109,N_6624,N_7595);
and U10110 (N_10110,N_7109,N_7031);
and U10111 (N_10111,N_7080,N_6163);
nor U10112 (N_10112,N_8217,N_6435);
and U10113 (N_10113,N_8991,N_6325);
and U10114 (N_10114,N_7847,N_6893);
or U10115 (N_10115,N_8657,N_8558);
nor U10116 (N_10116,N_6992,N_8793);
nor U10117 (N_10117,N_7539,N_6041);
nand U10118 (N_10118,N_8586,N_7970);
or U10119 (N_10119,N_6955,N_7905);
nor U10120 (N_10120,N_8410,N_8131);
or U10121 (N_10121,N_7193,N_8687);
and U10122 (N_10122,N_8313,N_7634);
nand U10123 (N_10123,N_8373,N_8584);
nand U10124 (N_10124,N_8429,N_7059);
nor U10125 (N_10125,N_8367,N_6610);
nor U10126 (N_10126,N_8361,N_6372);
nand U10127 (N_10127,N_6939,N_8317);
or U10128 (N_10128,N_8813,N_7692);
nor U10129 (N_10129,N_7612,N_7231);
or U10130 (N_10130,N_6409,N_8396);
nor U10131 (N_10131,N_6597,N_6627);
or U10132 (N_10132,N_6803,N_8002);
nand U10133 (N_10133,N_8573,N_7377);
or U10134 (N_10134,N_8196,N_6816);
or U10135 (N_10135,N_7917,N_6309);
nand U10136 (N_10136,N_7976,N_7374);
or U10137 (N_10137,N_8194,N_6444);
or U10138 (N_10138,N_8614,N_7923);
or U10139 (N_10139,N_6768,N_8765);
and U10140 (N_10140,N_8960,N_8679);
and U10141 (N_10141,N_7884,N_7722);
nor U10142 (N_10142,N_8041,N_7832);
nor U10143 (N_10143,N_7995,N_7195);
nor U10144 (N_10144,N_7433,N_8089);
nand U10145 (N_10145,N_8886,N_7347);
nand U10146 (N_10146,N_7116,N_6206);
or U10147 (N_10147,N_7828,N_6468);
nand U10148 (N_10148,N_6995,N_7943);
or U10149 (N_10149,N_7785,N_8115);
or U10150 (N_10150,N_6134,N_7546);
and U10151 (N_10151,N_8643,N_6565);
nand U10152 (N_10152,N_7507,N_8213);
nor U10153 (N_10153,N_7950,N_8807);
nand U10154 (N_10154,N_6255,N_8310);
and U10155 (N_10155,N_6027,N_6707);
nand U10156 (N_10156,N_7012,N_8579);
nand U10157 (N_10157,N_6953,N_6994);
nor U10158 (N_10158,N_7362,N_6005);
or U10159 (N_10159,N_8730,N_6964);
and U10160 (N_10160,N_7771,N_8826);
nor U10161 (N_10161,N_7543,N_8696);
nor U10162 (N_10162,N_8681,N_7581);
nand U10163 (N_10163,N_8724,N_6930);
nor U10164 (N_10164,N_7880,N_7775);
nor U10165 (N_10165,N_6598,N_6214);
nor U10166 (N_10166,N_7492,N_6735);
and U10167 (N_10167,N_6625,N_8455);
nor U10168 (N_10168,N_6959,N_8790);
nand U10169 (N_10169,N_8917,N_8277);
or U10170 (N_10170,N_8754,N_6794);
nand U10171 (N_10171,N_6422,N_7236);
nand U10172 (N_10172,N_7194,N_8187);
and U10173 (N_10173,N_6581,N_7827);
nand U10174 (N_10174,N_7978,N_8824);
nor U10175 (N_10175,N_6276,N_6861);
nor U10176 (N_10176,N_8740,N_7158);
nand U10177 (N_10177,N_7382,N_7270);
nand U10178 (N_10178,N_8783,N_8214);
or U10179 (N_10179,N_8916,N_6384);
and U10180 (N_10180,N_8961,N_7531);
and U10181 (N_10181,N_8834,N_8092);
or U10182 (N_10182,N_6288,N_8169);
or U10183 (N_10183,N_6475,N_7535);
and U10184 (N_10184,N_8421,N_6185);
and U10185 (N_10185,N_8716,N_8165);
nor U10186 (N_10186,N_6209,N_6851);
nand U10187 (N_10187,N_7114,N_7807);
nor U10188 (N_10188,N_6989,N_7015);
nand U10189 (N_10189,N_8175,N_8039);
and U10190 (N_10190,N_8901,N_6137);
nand U10191 (N_10191,N_8107,N_6972);
nand U10192 (N_10192,N_7315,N_6418);
nand U10193 (N_10193,N_7078,N_8255);
or U10194 (N_10194,N_8787,N_6269);
and U10195 (N_10195,N_6478,N_6685);
and U10196 (N_10196,N_6055,N_7340);
or U10197 (N_10197,N_6416,N_8628);
or U10198 (N_10198,N_8604,N_8017);
nand U10199 (N_10199,N_7021,N_8630);
nor U10200 (N_10200,N_6321,N_6224);
nand U10201 (N_10201,N_8416,N_8032);
nand U10202 (N_10202,N_6195,N_8535);
nor U10203 (N_10203,N_6220,N_7457);
nor U10204 (N_10204,N_7410,N_8443);
nand U10205 (N_10205,N_6801,N_6900);
or U10206 (N_10206,N_8944,N_6036);
or U10207 (N_10207,N_8063,N_7482);
nand U10208 (N_10208,N_8583,N_7743);
or U10209 (N_10209,N_6928,N_7900);
nor U10210 (N_10210,N_7994,N_6091);
or U10211 (N_10211,N_8682,N_6354);
or U10212 (N_10212,N_8705,N_7142);
or U10213 (N_10213,N_6948,N_6863);
or U10214 (N_10214,N_6844,N_6739);
and U10215 (N_10215,N_8817,N_7809);
nor U10216 (N_10216,N_6692,N_7210);
nor U10217 (N_10217,N_8522,N_6981);
nand U10218 (N_10218,N_7977,N_8091);
nor U10219 (N_10219,N_6457,N_8349);
and U10220 (N_10220,N_7466,N_8384);
nand U10221 (N_10221,N_7778,N_6870);
nor U10222 (N_10222,N_8081,N_7381);
and U10223 (N_10223,N_7500,N_7491);
or U10224 (N_10224,N_6789,N_6857);
and U10225 (N_10225,N_8590,N_8339);
nand U10226 (N_10226,N_7028,N_7201);
nand U10227 (N_10227,N_7566,N_6274);
and U10228 (N_10228,N_7714,N_8338);
nand U10229 (N_10229,N_7447,N_8747);
nand U10230 (N_10230,N_7327,N_8963);
and U10231 (N_10231,N_8434,N_7395);
nor U10232 (N_10232,N_7287,N_6368);
nor U10233 (N_10233,N_8068,N_7703);
and U10234 (N_10234,N_7896,N_6424);
nand U10235 (N_10235,N_8967,N_7659);
and U10236 (N_10236,N_6429,N_7030);
nor U10237 (N_10237,N_6272,N_8394);
and U10238 (N_10238,N_7580,N_8616);
nor U10239 (N_10239,N_7885,N_7513);
and U10240 (N_10240,N_6550,N_8431);
and U10241 (N_10241,N_8216,N_6019);
or U10242 (N_10242,N_8125,N_7735);
nand U10243 (N_10243,N_8442,N_6477);
or U10244 (N_10244,N_7526,N_8508);
and U10245 (N_10245,N_6362,N_6229);
nand U10246 (N_10246,N_7895,N_6574);
nor U10247 (N_10247,N_7927,N_8521);
or U10248 (N_10248,N_7523,N_7441);
and U10249 (N_10249,N_6683,N_7003);
or U10250 (N_10250,N_6982,N_7219);
and U10251 (N_10251,N_7553,N_7561);
or U10252 (N_10252,N_6026,N_7687);
nand U10253 (N_10253,N_6765,N_8566);
or U10254 (N_10254,N_6243,N_7129);
nor U10255 (N_10255,N_8144,N_8335);
and U10256 (N_10256,N_7672,N_7712);
nand U10257 (N_10257,N_8874,N_6714);
and U10258 (N_10258,N_8627,N_6559);
or U10259 (N_10259,N_7209,N_8170);
and U10260 (N_10260,N_6757,N_8833);
nand U10261 (N_10261,N_6002,N_8970);
or U10262 (N_10262,N_7732,N_8123);
or U10263 (N_10263,N_6006,N_7556);
and U10264 (N_10264,N_7339,N_7113);
or U10265 (N_10265,N_7681,N_7648);
nand U10266 (N_10266,N_8207,N_7989);
or U10267 (N_10267,N_8713,N_8798);
and U10268 (N_10268,N_7706,N_7939);
nor U10269 (N_10269,N_7733,N_6154);
nor U10270 (N_10270,N_6225,N_6151);
nor U10271 (N_10271,N_7873,N_8400);
nand U10272 (N_10272,N_8040,N_6169);
nor U10273 (N_10273,N_7135,N_7890);
and U10274 (N_10274,N_6086,N_7276);
and U10275 (N_10275,N_6945,N_8403);
or U10276 (N_10276,N_7534,N_7170);
and U10277 (N_10277,N_6543,N_6374);
nand U10278 (N_10278,N_6067,N_8490);
or U10279 (N_10279,N_6562,N_8937);
and U10280 (N_10280,N_8043,N_8862);
nand U10281 (N_10281,N_8720,N_6440);
or U10282 (N_10282,N_6144,N_8622);
nand U10283 (N_10283,N_7494,N_7619);
nand U10284 (N_10284,N_7678,N_8356);
nor U10285 (N_10285,N_6326,N_7363);
nor U10286 (N_10286,N_6389,N_6874);
xor U10287 (N_10287,N_7926,N_8517);
and U10288 (N_10288,N_6323,N_7166);
or U10289 (N_10289,N_7344,N_7739);
nor U10290 (N_10290,N_7254,N_6118);
and U10291 (N_10291,N_8866,N_6947);
nor U10292 (N_10292,N_8652,N_8060);
and U10293 (N_10293,N_8133,N_6013);
nand U10294 (N_10294,N_7606,N_8552);
nand U10295 (N_10295,N_6314,N_6097);
or U10296 (N_10296,N_8714,N_6329);
xor U10297 (N_10297,N_6476,N_6532);
or U10298 (N_10298,N_8326,N_6545);
or U10299 (N_10299,N_6250,N_8532);
or U10300 (N_10300,N_6049,N_7464);
or U10301 (N_10301,N_8203,N_8030);
nand U10302 (N_10302,N_6935,N_6380);
nor U10303 (N_10303,N_7292,N_6282);
nand U10304 (N_10304,N_7882,N_7033);
nand U10305 (N_10305,N_6039,N_8631);
and U10306 (N_10306,N_7922,N_8415);
nand U10307 (N_10307,N_7806,N_6450);
nor U10308 (N_10308,N_6913,N_6010);
or U10309 (N_10309,N_6924,N_8293);
xnor U10310 (N_10310,N_8891,N_8167);
or U10311 (N_10311,N_7217,N_8074);
nor U10312 (N_10312,N_8784,N_6649);
nor U10313 (N_10313,N_7760,N_6357);
nor U10314 (N_10314,N_8520,N_7957);
or U10315 (N_10315,N_8332,N_8100);
or U10316 (N_10316,N_6807,N_8225);
or U10317 (N_10317,N_6059,N_6554);
nor U10318 (N_10318,N_6910,N_7430);
or U10319 (N_10319,N_7914,N_8976);
nor U10320 (N_10320,N_8146,N_8406);
or U10321 (N_10321,N_8858,N_6119);
or U10322 (N_10322,N_8407,N_6929);
nand U10323 (N_10323,N_7227,N_8072);
or U10324 (N_10324,N_7811,N_7878);
nand U10325 (N_10325,N_6703,N_8781);
nor U10326 (N_10326,N_8398,N_8983);
nor U10327 (N_10327,N_6564,N_7872);
nor U10328 (N_10328,N_8494,N_7898);
nor U10329 (N_10329,N_8557,N_6153);
nor U10330 (N_10330,N_8542,N_6470);
and U10331 (N_10331,N_7501,N_6114);
and U10332 (N_10332,N_6896,N_8749);
and U10333 (N_10333,N_6174,N_7308);
nor U10334 (N_10334,N_7016,N_6493);
nand U10335 (N_10335,N_7131,N_6469);
and U10336 (N_10336,N_8174,N_7260);
nand U10337 (N_10337,N_7090,N_8545);
nor U10338 (N_10338,N_7966,N_8447);
nand U10339 (N_10339,N_6871,N_7967);
nor U10340 (N_10340,N_7557,N_6551);
and U10341 (N_10341,N_7993,N_7411);
and U10342 (N_10342,N_8094,N_8504);
and U10343 (N_10343,N_7680,N_6099);
nand U10344 (N_10344,N_8300,N_8162);
or U10345 (N_10345,N_7675,N_6356);
or U10346 (N_10346,N_6927,N_6222);
nor U10347 (N_10347,N_8087,N_7858);
and U10348 (N_10348,N_7091,N_8232);
nor U10349 (N_10349,N_7431,N_6043);
nand U10350 (N_10350,N_8110,N_6639);
and U10351 (N_10351,N_8854,N_6208);
and U10352 (N_10352,N_8731,N_8536);
and U10353 (N_10353,N_6491,N_6246);
xor U10354 (N_10354,N_6441,N_6616);
or U10355 (N_10355,N_8699,N_7694);
nand U10356 (N_10356,N_8788,N_6258);
nor U10357 (N_10357,N_6780,N_8301);
nor U10358 (N_10358,N_8786,N_6333);
and U10359 (N_10359,N_6093,N_8432);
and U10360 (N_10360,N_7829,N_8701);
or U10361 (N_10361,N_6880,N_6680);
or U10362 (N_10362,N_7215,N_6740);
or U10363 (N_10363,N_8328,N_7037);
nand U10364 (N_10364,N_6196,N_8663);
nor U10365 (N_10365,N_7800,N_8467);
nand U10366 (N_10366,N_7716,N_7641);
and U10367 (N_10367,N_8835,N_6763);
nand U10368 (N_10368,N_7550,N_8117);
or U10369 (N_10369,N_7983,N_6937);
nor U10370 (N_10370,N_6500,N_6737);
or U10371 (N_10371,N_7304,N_8569);
or U10372 (N_10372,N_6720,N_6699);
nor U10373 (N_10373,N_7232,N_8839);
or U10374 (N_10374,N_8645,N_6850);
nand U10375 (N_10375,N_7490,N_8464);
or U10376 (N_10376,N_7175,N_8733);
nor U10377 (N_10377,N_6262,N_6407);
or U10378 (N_10378,N_8341,N_7047);
nand U10379 (N_10379,N_7924,N_6466);
nor U10380 (N_10380,N_6399,N_8553);
or U10381 (N_10381,N_8931,N_8013);
nand U10382 (N_10382,N_6458,N_6249);
or U10383 (N_10383,N_6881,N_7506);
nand U10384 (N_10384,N_6115,N_6808);
nand U10385 (N_10385,N_7400,N_8154);
nand U10386 (N_10386,N_7182,N_6862);
nor U10387 (N_10387,N_8001,N_7679);
or U10388 (N_10388,N_6671,N_7042);
and U10389 (N_10389,N_6827,N_6023);
nand U10390 (N_10390,N_7931,N_8205);
and U10391 (N_10391,N_6014,N_7024);
or U10392 (N_10392,N_8568,N_7432);
or U10393 (N_10393,N_8605,N_7888);
or U10394 (N_10394,N_6123,N_7058);
nand U10395 (N_10395,N_7249,N_8587);
nor U10396 (N_10396,N_8268,N_8182);
and U10397 (N_10397,N_8238,N_8297);
or U10398 (N_10398,N_7034,N_7097);
nor U10399 (N_10399,N_6145,N_6056);
and U10400 (N_10400,N_7167,N_7295);
or U10401 (N_10401,N_6223,N_8437);
nor U10402 (N_10402,N_8537,N_8140);
and U10403 (N_10403,N_6373,N_6837);
and U10404 (N_10404,N_7160,N_7486);
and U10405 (N_10405,N_8079,N_8445);
nand U10406 (N_10406,N_8387,N_7259);
or U10407 (N_10407,N_8408,N_8346);
nand U10408 (N_10408,N_7277,N_6855);
or U10409 (N_10409,N_8808,N_8446);
nor U10410 (N_10410,N_7770,N_8137);
and U10411 (N_10411,N_7661,N_8928);
nand U10412 (N_10412,N_7842,N_8474);
or U10413 (N_10413,N_6479,N_6164);
nor U10414 (N_10414,N_6187,N_8235);
nor U10415 (N_10415,N_6985,N_8849);
and U10416 (N_10416,N_7688,N_8343);
nand U10417 (N_10417,N_7290,N_6914);
nor U10418 (N_10418,N_7298,N_7316);
or U10419 (N_10419,N_7108,N_8489);
or U10420 (N_10420,N_6800,N_7867);
or U10421 (N_10421,N_8821,N_8718);
nand U10422 (N_10422,N_7804,N_7137);
and U10423 (N_10423,N_8430,N_8185);
and U10424 (N_10424,N_8337,N_8513);
nor U10425 (N_10425,N_6341,N_8417);
nand U10426 (N_10426,N_7176,N_8460);
nand U10427 (N_10427,N_8669,N_6184);
nand U10428 (N_10428,N_8444,N_6706);
or U10429 (N_10429,N_8988,N_8292);
nor U10430 (N_10430,N_8993,N_8004);
and U10431 (N_10431,N_7696,N_6751);
nand U10432 (N_10432,N_8640,N_6840);
nand U10433 (N_10433,N_7869,N_8611);
and U10434 (N_10434,N_8767,N_7545);
or U10435 (N_10435,N_6335,N_8923);
nor U10436 (N_10436,N_7161,N_6492);
or U10437 (N_10437,N_7407,N_7365);
or U10438 (N_10438,N_6848,N_8192);
nand U10439 (N_10439,N_8809,N_6490);
or U10440 (N_10440,N_7198,N_7691);
or U10441 (N_10441,N_8876,N_8366);
or U10442 (N_10442,N_6548,N_7704);
nand U10443 (N_10443,N_8351,N_7041);
nor U10444 (N_10444,N_8158,N_8711);
nand U10445 (N_10445,N_8585,N_6488);
and U10446 (N_10446,N_8433,N_6644);
and U10447 (N_10447,N_6251,N_7102);
nor U10448 (N_10448,N_7670,N_6121);
or U10449 (N_10449,N_7915,N_8129);
nor U10450 (N_10450,N_8775,N_6899);
or U10451 (N_10451,N_6507,N_7428);
nor U10452 (N_10452,N_7480,N_8840);
or U10453 (N_10453,N_8496,N_6287);
or U10454 (N_10454,N_8811,N_7396);
and U10455 (N_10455,N_6586,N_7095);
or U10456 (N_10456,N_8828,N_8180);
and U10457 (N_10457,N_8224,N_8672);
or U10458 (N_10458,N_8053,N_6693);
nand U10459 (N_10459,N_7186,N_8066);
and U10460 (N_10460,N_7584,N_7128);
nand U10461 (N_10461,N_7264,N_7981);
and U10462 (N_10462,N_8046,N_8395);
nand U10463 (N_10463,N_6520,N_6875);
and U10464 (N_10464,N_7852,N_6347);
and U10465 (N_10465,N_8427,N_8610);
nor U10466 (N_10466,N_6898,N_6822);
or U10467 (N_10467,N_8903,N_8791);
nor U10468 (N_10468,N_8166,N_6419);
nor U10469 (N_10469,N_8152,N_8461);
or U10470 (N_10470,N_7200,N_8018);
nand U10471 (N_10471,N_6136,N_8130);
or U10472 (N_10472,N_6345,N_7072);
or U10473 (N_10473,N_6210,N_8176);
nand U10474 (N_10474,N_6289,N_7579);
or U10475 (N_10475,N_6547,N_8486);
and U10476 (N_10476,N_8029,N_8785);
nor U10477 (N_10477,N_7405,N_7527);
nand U10478 (N_10478,N_7077,N_7815);
or U10479 (N_10479,N_6485,N_6926);
or U10480 (N_10480,N_7355,N_8561);
nand U10481 (N_10481,N_8449,N_6339);
nand U10482 (N_10482,N_7763,N_6731);
nor U10483 (N_10483,N_7472,N_7886);
nor U10484 (N_10484,N_6188,N_8121);
nand U10485 (N_10485,N_8831,N_7769);
nor U10486 (N_10486,N_6960,N_7836);
nand U10487 (N_10487,N_6433,N_6437);
xor U10488 (N_10488,N_7839,N_8275);
nand U10489 (N_10489,N_8318,N_8543);
and U10490 (N_10490,N_6846,N_6103);
or U10491 (N_10491,N_8848,N_6286);
and U10492 (N_10492,N_6342,N_8850);
nor U10493 (N_10493,N_7729,N_6334);
or U10494 (N_10494,N_7138,N_7266);
and U10495 (N_10495,N_8305,N_6733);
nor U10496 (N_10496,N_7406,N_7638);
and U10497 (N_10497,N_8957,N_6378);
or U10498 (N_10498,N_8302,N_6428);
nor U10499 (N_10499,N_7368,N_7380);
nand U10500 (N_10500,N_6215,N_7603);
nor U10501 (N_10501,N_8410,N_6359);
nor U10502 (N_10502,N_8928,N_7477);
nand U10503 (N_10503,N_7653,N_8291);
or U10504 (N_10504,N_7781,N_7353);
nor U10505 (N_10505,N_8220,N_7951);
or U10506 (N_10506,N_8390,N_8278);
nand U10507 (N_10507,N_7215,N_6673);
nand U10508 (N_10508,N_7951,N_6032);
nor U10509 (N_10509,N_7285,N_7079);
nand U10510 (N_10510,N_8094,N_6782);
nor U10511 (N_10511,N_7917,N_6819);
nor U10512 (N_10512,N_7601,N_6185);
or U10513 (N_10513,N_6564,N_7132);
and U10514 (N_10514,N_8115,N_8047);
or U10515 (N_10515,N_8643,N_8313);
nor U10516 (N_10516,N_6329,N_7438);
nand U10517 (N_10517,N_8094,N_6440);
nor U10518 (N_10518,N_7219,N_8581);
or U10519 (N_10519,N_6030,N_7231);
nand U10520 (N_10520,N_8994,N_6327);
nor U10521 (N_10521,N_7577,N_7924);
nor U10522 (N_10522,N_7960,N_7487);
or U10523 (N_10523,N_6957,N_7830);
nand U10524 (N_10524,N_8410,N_7662);
or U10525 (N_10525,N_6189,N_6444);
and U10526 (N_10526,N_6037,N_6451);
and U10527 (N_10527,N_7296,N_8449);
and U10528 (N_10528,N_8532,N_6964);
or U10529 (N_10529,N_6951,N_7138);
nor U10530 (N_10530,N_6477,N_7493);
nor U10531 (N_10531,N_8090,N_7825);
or U10532 (N_10532,N_7397,N_7290);
nor U10533 (N_10533,N_6350,N_8241);
and U10534 (N_10534,N_8150,N_6035);
or U10535 (N_10535,N_6752,N_6857);
and U10536 (N_10536,N_8408,N_7226);
or U10537 (N_10537,N_6567,N_6246);
and U10538 (N_10538,N_8896,N_7244);
or U10539 (N_10539,N_8809,N_6440);
and U10540 (N_10540,N_7032,N_8931);
nor U10541 (N_10541,N_8899,N_7725);
nand U10542 (N_10542,N_6851,N_6032);
and U10543 (N_10543,N_6624,N_7492);
nand U10544 (N_10544,N_8127,N_7898);
nor U10545 (N_10545,N_6376,N_6713);
nand U10546 (N_10546,N_8996,N_6891);
nand U10547 (N_10547,N_6873,N_7775);
nor U10548 (N_10548,N_7106,N_6588);
and U10549 (N_10549,N_7966,N_6337);
nor U10550 (N_10550,N_6477,N_7788);
or U10551 (N_10551,N_7258,N_6535);
nor U10552 (N_10552,N_7175,N_8470);
nand U10553 (N_10553,N_6126,N_8095);
xnor U10554 (N_10554,N_7595,N_6415);
nand U10555 (N_10555,N_8580,N_8309);
and U10556 (N_10556,N_8715,N_7726);
and U10557 (N_10557,N_6910,N_6629);
and U10558 (N_10558,N_8592,N_7524);
nor U10559 (N_10559,N_7356,N_6636);
nor U10560 (N_10560,N_7254,N_6621);
or U10561 (N_10561,N_7927,N_8404);
nand U10562 (N_10562,N_8704,N_7247);
nand U10563 (N_10563,N_8150,N_7211);
nand U10564 (N_10564,N_8300,N_6455);
nor U10565 (N_10565,N_6015,N_6302);
and U10566 (N_10566,N_6942,N_7470);
and U10567 (N_10567,N_8329,N_7679);
nand U10568 (N_10568,N_6822,N_7180);
nor U10569 (N_10569,N_7080,N_8781);
nand U10570 (N_10570,N_7491,N_7056);
or U10571 (N_10571,N_7999,N_8704);
nand U10572 (N_10572,N_8502,N_8690);
or U10573 (N_10573,N_8568,N_7764);
nor U10574 (N_10574,N_8594,N_8161);
nand U10575 (N_10575,N_7785,N_7609);
and U10576 (N_10576,N_8862,N_7213);
and U10577 (N_10577,N_7976,N_6477);
and U10578 (N_10578,N_8494,N_6568);
nand U10579 (N_10579,N_6475,N_6758);
nand U10580 (N_10580,N_8920,N_6622);
nand U10581 (N_10581,N_6347,N_7244);
nor U10582 (N_10582,N_7544,N_6522);
nor U10583 (N_10583,N_6544,N_7362);
nor U10584 (N_10584,N_7486,N_6447);
nand U10585 (N_10585,N_7625,N_7196);
nand U10586 (N_10586,N_7151,N_8634);
and U10587 (N_10587,N_7854,N_8546);
or U10588 (N_10588,N_6614,N_7700);
and U10589 (N_10589,N_7374,N_8138);
nor U10590 (N_10590,N_7189,N_6621);
nand U10591 (N_10591,N_7927,N_6069);
and U10592 (N_10592,N_7591,N_8687);
nand U10593 (N_10593,N_8716,N_8975);
and U10594 (N_10594,N_6532,N_7394);
and U10595 (N_10595,N_6985,N_6321);
nand U10596 (N_10596,N_6733,N_6908);
or U10597 (N_10597,N_6758,N_8826);
nor U10598 (N_10598,N_7849,N_7892);
and U10599 (N_10599,N_8058,N_8018);
or U10600 (N_10600,N_6722,N_8005);
nor U10601 (N_10601,N_7601,N_6887);
nor U10602 (N_10602,N_8773,N_6615);
nand U10603 (N_10603,N_7433,N_6521);
nand U10604 (N_10604,N_8633,N_8806);
and U10605 (N_10605,N_6157,N_8802);
or U10606 (N_10606,N_6345,N_8729);
or U10607 (N_10607,N_6724,N_7892);
and U10608 (N_10608,N_6274,N_7289);
or U10609 (N_10609,N_7140,N_8448);
and U10610 (N_10610,N_7877,N_8130);
or U10611 (N_10611,N_8087,N_8428);
nor U10612 (N_10612,N_8765,N_7017);
or U10613 (N_10613,N_7002,N_6056);
nor U10614 (N_10614,N_7997,N_7572);
nand U10615 (N_10615,N_7335,N_8259);
and U10616 (N_10616,N_6780,N_8663);
nor U10617 (N_10617,N_6737,N_8052);
nor U10618 (N_10618,N_7590,N_6521);
nand U10619 (N_10619,N_8261,N_7619);
or U10620 (N_10620,N_6034,N_6739);
nand U10621 (N_10621,N_8476,N_8041);
and U10622 (N_10622,N_8219,N_6833);
nor U10623 (N_10623,N_8050,N_7685);
and U10624 (N_10624,N_7007,N_8601);
xor U10625 (N_10625,N_8694,N_6893);
nor U10626 (N_10626,N_6766,N_6655);
nor U10627 (N_10627,N_7440,N_8023);
nand U10628 (N_10628,N_8557,N_6568);
and U10629 (N_10629,N_7902,N_7707);
and U10630 (N_10630,N_7287,N_6812);
and U10631 (N_10631,N_6634,N_8032);
nor U10632 (N_10632,N_8337,N_8653);
nand U10633 (N_10633,N_8279,N_8113);
and U10634 (N_10634,N_6181,N_6045);
nand U10635 (N_10635,N_7301,N_8749);
nand U10636 (N_10636,N_7762,N_6697);
nand U10637 (N_10637,N_6077,N_6513);
or U10638 (N_10638,N_8482,N_8254);
nor U10639 (N_10639,N_7449,N_7897);
or U10640 (N_10640,N_8241,N_7590);
nor U10641 (N_10641,N_7295,N_8487);
nand U10642 (N_10642,N_7849,N_6208);
nand U10643 (N_10643,N_7074,N_7017);
or U10644 (N_10644,N_7800,N_7236);
nand U10645 (N_10645,N_8000,N_7856);
or U10646 (N_10646,N_8379,N_7772);
nor U10647 (N_10647,N_7295,N_8473);
nand U10648 (N_10648,N_6274,N_6816);
nor U10649 (N_10649,N_6618,N_8015);
nand U10650 (N_10650,N_8181,N_7303);
and U10651 (N_10651,N_7422,N_8522);
nor U10652 (N_10652,N_6862,N_7022);
and U10653 (N_10653,N_8486,N_7488);
nor U10654 (N_10654,N_8034,N_6482);
and U10655 (N_10655,N_8118,N_8967);
nor U10656 (N_10656,N_6886,N_8500);
nor U10657 (N_10657,N_6317,N_8361);
nand U10658 (N_10658,N_8703,N_7725);
nand U10659 (N_10659,N_6205,N_7526);
or U10660 (N_10660,N_7552,N_8290);
nand U10661 (N_10661,N_8829,N_7073);
nand U10662 (N_10662,N_8124,N_6122);
nor U10663 (N_10663,N_8152,N_8037);
and U10664 (N_10664,N_8213,N_7583);
and U10665 (N_10665,N_7065,N_6308);
or U10666 (N_10666,N_7237,N_7181);
nand U10667 (N_10667,N_6649,N_6819);
nand U10668 (N_10668,N_7680,N_6725);
and U10669 (N_10669,N_7864,N_8139);
or U10670 (N_10670,N_6869,N_8536);
or U10671 (N_10671,N_6425,N_8145);
nand U10672 (N_10672,N_6417,N_6066);
nand U10673 (N_10673,N_7318,N_8975);
or U10674 (N_10674,N_6048,N_7109);
and U10675 (N_10675,N_8346,N_6137);
and U10676 (N_10676,N_8539,N_7827);
nor U10677 (N_10677,N_8151,N_7153);
and U10678 (N_10678,N_6360,N_8628);
and U10679 (N_10679,N_6023,N_7725);
or U10680 (N_10680,N_7574,N_8038);
or U10681 (N_10681,N_8424,N_7761);
nor U10682 (N_10682,N_6088,N_6671);
and U10683 (N_10683,N_7949,N_6688);
nor U10684 (N_10684,N_6690,N_7892);
and U10685 (N_10685,N_7589,N_6804);
nand U10686 (N_10686,N_8680,N_6741);
nor U10687 (N_10687,N_7501,N_6373);
and U10688 (N_10688,N_7808,N_7039);
and U10689 (N_10689,N_7188,N_8234);
nor U10690 (N_10690,N_6254,N_8755);
or U10691 (N_10691,N_8763,N_8171);
and U10692 (N_10692,N_6931,N_7306);
or U10693 (N_10693,N_7482,N_6647);
nor U10694 (N_10694,N_6930,N_7308);
and U10695 (N_10695,N_7681,N_8094);
nor U10696 (N_10696,N_8156,N_6891);
or U10697 (N_10697,N_7166,N_6307);
and U10698 (N_10698,N_6732,N_8431);
nand U10699 (N_10699,N_8545,N_8816);
nand U10700 (N_10700,N_7324,N_8196);
xor U10701 (N_10701,N_8357,N_8787);
or U10702 (N_10702,N_7007,N_8775);
or U10703 (N_10703,N_8275,N_7848);
nor U10704 (N_10704,N_6383,N_7108);
nor U10705 (N_10705,N_8734,N_6571);
and U10706 (N_10706,N_8469,N_6649);
nand U10707 (N_10707,N_6650,N_7880);
nand U10708 (N_10708,N_7950,N_7151);
or U10709 (N_10709,N_6632,N_7868);
or U10710 (N_10710,N_7095,N_7388);
or U10711 (N_10711,N_8399,N_7411);
and U10712 (N_10712,N_7905,N_6390);
or U10713 (N_10713,N_7624,N_8736);
or U10714 (N_10714,N_8082,N_7204);
and U10715 (N_10715,N_6942,N_8572);
and U10716 (N_10716,N_8774,N_8956);
or U10717 (N_10717,N_6529,N_7686);
nor U10718 (N_10718,N_8672,N_6730);
and U10719 (N_10719,N_8439,N_8318);
nand U10720 (N_10720,N_6004,N_8811);
or U10721 (N_10721,N_7531,N_6577);
and U10722 (N_10722,N_7564,N_8546);
or U10723 (N_10723,N_7738,N_8224);
nor U10724 (N_10724,N_7777,N_7909);
nor U10725 (N_10725,N_7530,N_6315);
and U10726 (N_10726,N_7584,N_6206);
or U10727 (N_10727,N_7521,N_8597);
nand U10728 (N_10728,N_8640,N_7963);
nor U10729 (N_10729,N_6227,N_8181);
nand U10730 (N_10730,N_8144,N_7917);
nor U10731 (N_10731,N_7492,N_6769);
or U10732 (N_10732,N_6639,N_8131);
nand U10733 (N_10733,N_7558,N_8551);
or U10734 (N_10734,N_8291,N_6932);
nor U10735 (N_10735,N_7337,N_6707);
or U10736 (N_10736,N_8987,N_7875);
nor U10737 (N_10737,N_7613,N_7516);
and U10738 (N_10738,N_7951,N_6473);
or U10739 (N_10739,N_8270,N_7381);
or U10740 (N_10740,N_6555,N_7978);
or U10741 (N_10741,N_8505,N_7255);
nand U10742 (N_10742,N_8338,N_6774);
nor U10743 (N_10743,N_7637,N_7506);
and U10744 (N_10744,N_8383,N_8172);
and U10745 (N_10745,N_6925,N_7897);
and U10746 (N_10746,N_8302,N_7346);
or U10747 (N_10747,N_6958,N_6593);
nor U10748 (N_10748,N_6183,N_6533);
nor U10749 (N_10749,N_6938,N_7498);
or U10750 (N_10750,N_8148,N_8133);
and U10751 (N_10751,N_6022,N_8099);
nand U10752 (N_10752,N_6016,N_6417);
nand U10753 (N_10753,N_6588,N_6794);
nor U10754 (N_10754,N_8095,N_6793);
and U10755 (N_10755,N_8504,N_6791);
or U10756 (N_10756,N_6487,N_6080);
nand U10757 (N_10757,N_7998,N_6521);
nand U10758 (N_10758,N_6635,N_8655);
and U10759 (N_10759,N_7217,N_6878);
nand U10760 (N_10760,N_6742,N_6901);
or U10761 (N_10761,N_6167,N_7480);
nand U10762 (N_10762,N_7616,N_8565);
nand U10763 (N_10763,N_8013,N_6579);
or U10764 (N_10764,N_8076,N_7991);
and U10765 (N_10765,N_6707,N_6424);
or U10766 (N_10766,N_6499,N_6444);
nand U10767 (N_10767,N_7029,N_8005);
and U10768 (N_10768,N_7530,N_8346);
and U10769 (N_10769,N_7618,N_6439);
or U10770 (N_10770,N_8389,N_8426);
or U10771 (N_10771,N_8324,N_7930);
nor U10772 (N_10772,N_7517,N_7599);
or U10773 (N_10773,N_7908,N_7856);
or U10774 (N_10774,N_7010,N_8344);
nor U10775 (N_10775,N_6044,N_8946);
or U10776 (N_10776,N_7357,N_7863);
or U10777 (N_10777,N_8930,N_8724);
xnor U10778 (N_10778,N_7168,N_6692);
nand U10779 (N_10779,N_6130,N_7649);
nand U10780 (N_10780,N_6867,N_8050);
and U10781 (N_10781,N_6407,N_7145);
or U10782 (N_10782,N_8175,N_6786);
or U10783 (N_10783,N_8238,N_8367);
and U10784 (N_10784,N_7769,N_6060);
nand U10785 (N_10785,N_6271,N_8912);
nor U10786 (N_10786,N_6457,N_7308);
or U10787 (N_10787,N_8088,N_7123);
nor U10788 (N_10788,N_8754,N_6531);
nor U10789 (N_10789,N_7858,N_8795);
nand U10790 (N_10790,N_6021,N_6349);
nor U10791 (N_10791,N_7500,N_7436);
nor U10792 (N_10792,N_7991,N_7285);
and U10793 (N_10793,N_7415,N_8707);
nand U10794 (N_10794,N_8155,N_8044);
and U10795 (N_10795,N_6598,N_7147);
nor U10796 (N_10796,N_8418,N_8562);
and U10797 (N_10797,N_8541,N_6902);
nor U10798 (N_10798,N_6637,N_6392);
and U10799 (N_10799,N_8498,N_6606);
and U10800 (N_10800,N_7555,N_6987);
nand U10801 (N_10801,N_8900,N_6058);
nand U10802 (N_10802,N_6949,N_8324);
and U10803 (N_10803,N_7654,N_7513);
nand U10804 (N_10804,N_8051,N_8434);
nand U10805 (N_10805,N_8558,N_7830);
nor U10806 (N_10806,N_7106,N_6811);
nand U10807 (N_10807,N_6840,N_7113);
nand U10808 (N_10808,N_7533,N_6607);
or U10809 (N_10809,N_6375,N_7357);
nor U10810 (N_10810,N_7327,N_8729);
nor U10811 (N_10811,N_7020,N_7438);
nor U10812 (N_10812,N_7838,N_6137);
nand U10813 (N_10813,N_8535,N_7441);
and U10814 (N_10814,N_7451,N_8467);
nand U10815 (N_10815,N_8799,N_7511);
xor U10816 (N_10816,N_7780,N_6527);
nor U10817 (N_10817,N_8836,N_6919);
and U10818 (N_10818,N_7910,N_7578);
nand U10819 (N_10819,N_7525,N_8308);
nor U10820 (N_10820,N_6180,N_8009);
nor U10821 (N_10821,N_8305,N_6177);
nand U10822 (N_10822,N_8617,N_8770);
or U10823 (N_10823,N_7594,N_8558);
or U10824 (N_10824,N_7223,N_7165);
nand U10825 (N_10825,N_8024,N_8577);
nor U10826 (N_10826,N_8618,N_7778);
and U10827 (N_10827,N_8375,N_6101);
or U10828 (N_10828,N_7012,N_6313);
nand U10829 (N_10829,N_6624,N_6335);
or U10830 (N_10830,N_6904,N_7509);
nor U10831 (N_10831,N_7081,N_8838);
nand U10832 (N_10832,N_8345,N_8654);
xor U10833 (N_10833,N_7339,N_6705);
nand U10834 (N_10834,N_8217,N_7919);
and U10835 (N_10835,N_6286,N_8248);
and U10836 (N_10836,N_7508,N_8904);
or U10837 (N_10837,N_6681,N_7933);
or U10838 (N_10838,N_6048,N_6145);
nor U10839 (N_10839,N_7588,N_6251);
nand U10840 (N_10840,N_7226,N_6925);
and U10841 (N_10841,N_8525,N_8033);
and U10842 (N_10842,N_8931,N_7273);
and U10843 (N_10843,N_7539,N_8154);
or U10844 (N_10844,N_7603,N_7199);
nand U10845 (N_10845,N_8207,N_7800);
nor U10846 (N_10846,N_6675,N_8103);
nand U10847 (N_10847,N_8712,N_6918);
nand U10848 (N_10848,N_8476,N_7776);
and U10849 (N_10849,N_7583,N_7813);
nor U10850 (N_10850,N_6988,N_8227);
nor U10851 (N_10851,N_7812,N_8796);
and U10852 (N_10852,N_7110,N_7005);
and U10853 (N_10853,N_7437,N_6169);
or U10854 (N_10854,N_6512,N_7105);
or U10855 (N_10855,N_6955,N_8393);
nor U10856 (N_10856,N_8042,N_7346);
nor U10857 (N_10857,N_7256,N_6771);
nor U10858 (N_10858,N_6281,N_6302);
or U10859 (N_10859,N_7517,N_8729);
or U10860 (N_10860,N_7302,N_8555);
nand U10861 (N_10861,N_7848,N_6012);
or U10862 (N_10862,N_7315,N_7002);
nand U10863 (N_10863,N_8915,N_7156);
nand U10864 (N_10864,N_7837,N_8828);
nand U10865 (N_10865,N_8868,N_7219);
or U10866 (N_10866,N_6900,N_6755);
nand U10867 (N_10867,N_6038,N_8827);
and U10868 (N_10868,N_8367,N_6524);
or U10869 (N_10869,N_8717,N_7908);
xnor U10870 (N_10870,N_8438,N_7435);
or U10871 (N_10871,N_7907,N_6662);
or U10872 (N_10872,N_7318,N_8845);
or U10873 (N_10873,N_7067,N_7833);
xnor U10874 (N_10874,N_8035,N_6728);
nand U10875 (N_10875,N_8148,N_6518);
nand U10876 (N_10876,N_6779,N_7031);
nor U10877 (N_10877,N_7361,N_8663);
and U10878 (N_10878,N_6731,N_8405);
nor U10879 (N_10879,N_8941,N_7609);
or U10880 (N_10880,N_7611,N_6657);
or U10881 (N_10881,N_6655,N_6761);
and U10882 (N_10882,N_7042,N_8782);
nor U10883 (N_10883,N_7335,N_7272);
and U10884 (N_10884,N_6529,N_7311);
and U10885 (N_10885,N_7434,N_8555);
nand U10886 (N_10886,N_8822,N_7818);
nand U10887 (N_10887,N_7434,N_6095);
nor U10888 (N_10888,N_8448,N_7078);
or U10889 (N_10889,N_7338,N_7834);
nor U10890 (N_10890,N_7598,N_8844);
and U10891 (N_10891,N_6676,N_6503);
nand U10892 (N_10892,N_8102,N_8929);
and U10893 (N_10893,N_6282,N_6758);
xor U10894 (N_10894,N_6404,N_6472);
and U10895 (N_10895,N_6605,N_8109);
or U10896 (N_10896,N_7441,N_7398);
and U10897 (N_10897,N_6695,N_7078);
or U10898 (N_10898,N_6028,N_7317);
nor U10899 (N_10899,N_6996,N_8286);
nand U10900 (N_10900,N_7767,N_6510);
nand U10901 (N_10901,N_6511,N_6400);
or U10902 (N_10902,N_6005,N_6552);
or U10903 (N_10903,N_7465,N_8684);
or U10904 (N_10904,N_8959,N_8416);
nor U10905 (N_10905,N_8614,N_6376);
or U10906 (N_10906,N_6162,N_8586);
and U10907 (N_10907,N_7791,N_6020);
or U10908 (N_10908,N_8409,N_6566);
nor U10909 (N_10909,N_8942,N_8670);
and U10910 (N_10910,N_8654,N_6042);
nor U10911 (N_10911,N_6902,N_8790);
nor U10912 (N_10912,N_8423,N_8293);
nand U10913 (N_10913,N_8781,N_7889);
nor U10914 (N_10914,N_6132,N_7413);
nand U10915 (N_10915,N_6243,N_7166);
and U10916 (N_10916,N_7404,N_6992);
and U10917 (N_10917,N_7258,N_6130);
and U10918 (N_10918,N_6055,N_6816);
nor U10919 (N_10919,N_7662,N_8706);
nor U10920 (N_10920,N_6970,N_8263);
nand U10921 (N_10921,N_6195,N_8146);
and U10922 (N_10922,N_8773,N_7992);
or U10923 (N_10923,N_6785,N_6889);
and U10924 (N_10924,N_7544,N_7397);
and U10925 (N_10925,N_8546,N_7625);
nand U10926 (N_10926,N_7431,N_7617);
nand U10927 (N_10927,N_6666,N_7601);
nand U10928 (N_10928,N_6602,N_7872);
and U10929 (N_10929,N_7817,N_7783);
nor U10930 (N_10930,N_6874,N_7964);
or U10931 (N_10931,N_6627,N_6832);
and U10932 (N_10932,N_6515,N_6607);
nand U10933 (N_10933,N_6068,N_6762);
and U10934 (N_10934,N_6404,N_8573);
and U10935 (N_10935,N_6916,N_8768);
nand U10936 (N_10936,N_8398,N_6508);
and U10937 (N_10937,N_7064,N_7548);
nand U10938 (N_10938,N_6352,N_7260);
and U10939 (N_10939,N_7349,N_6265);
xor U10940 (N_10940,N_8175,N_8406);
nor U10941 (N_10941,N_6050,N_8616);
and U10942 (N_10942,N_7909,N_7049);
nand U10943 (N_10943,N_8006,N_6505);
nand U10944 (N_10944,N_8642,N_8216);
and U10945 (N_10945,N_8694,N_6734);
nor U10946 (N_10946,N_8559,N_8404);
and U10947 (N_10947,N_7480,N_7299);
nand U10948 (N_10948,N_6243,N_8605);
and U10949 (N_10949,N_7141,N_8657);
or U10950 (N_10950,N_7384,N_6544);
and U10951 (N_10951,N_8847,N_6028);
nor U10952 (N_10952,N_8191,N_7915);
or U10953 (N_10953,N_7736,N_7720);
nor U10954 (N_10954,N_8791,N_8986);
nand U10955 (N_10955,N_6536,N_6916);
and U10956 (N_10956,N_8624,N_7897);
nand U10957 (N_10957,N_6211,N_7589);
and U10958 (N_10958,N_6554,N_7934);
and U10959 (N_10959,N_7280,N_7150);
and U10960 (N_10960,N_8467,N_8683);
nand U10961 (N_10961,N_6719,N_6841);
nand U10962 (N_10962,N_6271,N_7286);
or U10963 (N_10963,N_6373,N_6421);
and U10964 (N_10964,N_6311,N_6186);
or U10965 (N_10965,N_6126,N_6846);
and U10966 (N_10966,N_7925,N_6832);
nor U10967 (N_10967,N_8172,N_7611);
nand U10968 (N_10968,N_7305,N_8784);
and U10969 (N_10969,N_7129,N_8219);
or U10970 (N_10970,N_6345,N_7585);
nand U10971 (N_10971,N_8562,N_6904);
nor U10972 (N_10972,N_8896,N_7967);
and U10973 (N_10973,N_6431,N_6962);
nand U10974 (N_10974,N_6210,N_6458);
or U10975 (N_10975,N_8178,N_6236);
nand U10976 (N_10976,N_8232,N_7752);
nand U10977 (N_10977,N_6893,N_6452);
or U10978 (N_10978,N_8074,N_7664);
nand U10979 (N_10979,N_6639,N_6122);
and U10980 (N_10980,N_8031,N_8528);
nor U10981 (N_10981,N_8878,N_8500);
or U10982 (N_10982,N_7466,N_8593);
or U10983 (N_10983,N_6516,N_8827);
nand U10984 (N_10984,N_6334,N_6122);
nand U10985 (N_10985,N_6619,N_7047);
nor U10986 (N_10986,N_6261,N_7855);
and U10987 (N_10987,N_8691,N_8187);
nor U10988 (N_10988,N_8700,N_8716);
and U10989 (N_10989,N_6342,N_7358);
nand U10990 (N_10990,N_8993,N_6598);
and U10991 (N_10991,N_8162,N_6328);
or U10992 (N_10992,N_8046,N_8020);
nor U10993 (N_10993,N_7955,N_8098);
or U10994 (N_10994,N_6066,N_6845);
nor U10995 (N_10995,N_6504,N_7783);
or U10996 (N_10996,N_6580,N_8773);
nand U10997 (N_10997,N_8261,N_6085);
or U10998 (N_10998,N_8190,N_6723);
or U10999 (N_10999,N_8504,N_8305);
and U11000 (N_11000,N_8013,N_6537);
nor U11001 (N_11001,N_7063,N_8107);
nand U11002 (N_11002,N_6529,N_6103);
nand U11003 (N_11003,N_6338,N_8959);
nand U11004 (N_11004,N_8968,N_7147);
xnor U11005 (N_11005,N_6477,N_8910);
nand U11006 (N_11006,N_6598,N_7528);
and U11007 (N_11007,N_8270,N_7616);
or U11008 (N_11008,N_6027,N_7563);
nor U11009 (N_11009,N_6882,N_7999);
and U11010 (N_11010,N_6739,N_7965);
nand U11011 (N_11011,N_8602,N_8574);
nor U11012 (N_11012,N_7396,N_6739);
or U11013 (N_11013,N_6620,N_6618);
or U11014 (N_11014,N_8047,N_8851);
nand U11015 (N_11015,N_7403,N_6738);
or U11016 (N_11016,N_7493,N_8256);
and U11017 (N_11017,N_7475,N_6060);
nand U11018 (N_11018,N_7111,N_6504);
and U11019 (N_11019,N_8441,N_7909);
and U11020 (N_11020,N_6879,N_6764);
or U11021 (N_11021,N_8157,N_6001);
and U11022 (N_11022,N_8300,N_8372);
and U11023 (N_11023,N_6284,N_7924);
or U11024 (N_11024,N_6846,N_8308);
or U11025 (N_11025,N_8483,N_7428);
nand U11026 (N_11026,N_7107,N_7088);
and U11027 (N_11027,N_8531,N_6134);
and U11028 (N_11028,N_7524,N_8183);
nand U11029 (N_11029,N_6525,N_8167);
or U11030 (N_11030,N_6132,N_8086);
nand U11031 (N_11031,N_8467,N_7889);
nand U11032 (N_11032,N_8843,N_6877);
nand U11033 (N_11033,N_7926,N_7210);
nand U11034 (N_11034,N_8879,N_7117);
and U11035 (N_11035,N_8457,N_7000);
nand U11036 (N_11036,N_8281,N_7590);
nor U11037 (N_11037,N_7802,N_6761);
nand U11038 (N_11038,N_6103,N_7564);
nor U11039 (N_11039,N_6082,N_7098);
or U11040 (N_11040,N_6596,N_8234);
and U11041 (N_11041,N_7363,N_7606);
nand U11042 (N_11042,N_7321,N_7863);
nor U11043 (N_11043,N_8782,N_8231);
and U11044 (N_11044,N_7910,N_6499);
or U11045 (N_11045,N_8763,N_8211);
nor U11046 (N_11046,N_7997,N_6514);
xor U11047 (N_11047,N_6920,N_7051);
and U11048 (N_11048,N_6997,N_8320);
or U11049 (N_11049,N_6669,N_8431);
nor U11050 (N_11050,N_6593,N_8107);
or U11051 (N_11051,N_7116,N_7024);
and U11052 (N_11052,N_6356,N_6604);
nand U11053 (N_11053,N_8988,N_7798);
nor U11054 (N_11054,N_7019,N_7490);
nor U11055 (N_11055,N_7508,N_6254);
nand U11056 (N_11056,N_8149,N_6540);
and U11057 (N_11057,N_8955,N_7834);
and U11058 (N_11058,N_6597,N_8627);
nor U11059 (N_11059,N_8358,N_7582);
or U11060 (N_11060,N_6346,N_6770);
nand U11061 (N_11061,N_7527,N_8526);
nand U11062 (N_11062,N_7434,N_7367);
nor U11063 (N_11063,N_6184,N_7608);
and U11064 (N_11064,N_6731,N_7083);
and U11065 (N_11065,N_8844,N_7603);
nand U11066 (N_11066,N_8182,N_7865);
and U11067 (N_11067,N_8370,N_8032);
nor U11068 (N_11068,N_7544,N_8143);
or U11069 (N_11069,N_8835,N_6672);
nor U11070 (N_11070,N_7138,N_7513);
nand U11071 (N_11071,N_6256,N_7212);
and U11072 (N_11072,N_8605,N_7542);
or U11073 (N_11073,N_7662,N_6747);
or U11074 (N_11074,N_7909,N_6559);
nor U11075 (N_11075,N_6651,N_7023);
nand U11076 (N_11076,N_7876,N_7489);
nand U11077 (N_11077,N_7946,N_7731);
nor U11078 (N_11078,N_8903,N_8921);
nand U11079 (N_11079,N_6608,N_8396);
nand U11080 (N_11080,N_7154,N_7037);
nand U11081 (N_11081,N_7537,N_7649);
and U11082 (N_11082,N_7560,N_7992);
nand U11083 (N_11083,N_7100,N_8895);
nor U11084 (N_11084,N_6915,N_7408);
or U11085 (N_11085,N_7264,N_7293);
and U11086 (N_11086,N_8451,N_7933);
and U11087 (N_11087,N_8103,N_6703);
nor U11088 (N_11088,N_6620,N_7154);
nor U11089 (N_11089,N_7728,N_8068);
nand U11090 (N_11090,N_7663,N_6832);
and U11091 (N_11091,N_7959,N_8546);
or U11092 (N_11092,N_7341,N_8726);
or U11093 (N_11093,N_8774,N_8402);
and U11094 (N_11094,N_6241,N_8326);
nor U11095 (N_11095,N_6740,N_8303);
nor U11096 (N_11096,N_8714,N_7101);
nand U11097 (N_11097,N_6927,N_7084);
nor U11098 (N_11098,N_6614,N_6944);
nand U11099 (N_11099,N_8702,N_7113);
nand U11100 (N_11100,N_6108,N_8362);
nand U11101 (N_11101,N_7792,N_6883);
nor U11102 (N_11102,N_6985,N_6922);
nor U11103 (N_11103,N_7267,N_8299);
and U11104 (N_11104,N_6870,N_8597);
or U11105 (N_11105,N_7450,N_8881);
xor U11106 (N_11106,N_7499,N_8077);
nor U11107 (N_11107,N_7892,N_6586);
nand U11108 (N_11108,N_6219,N_6799);
or U11109 (N_11109,N_7097,N_6674);
or U11110 (N_11110,N_7833,N_7402);
nor U11111 (N_11111,N_8965,N_7776);
or U11112 (N_11112,N_6185,N_7289);
nor U11113 (N_11113,N_8028,N_6514);
or U11114 (N_11114,N_7565,N_8834);
and U11115 (N_11115,N_8273,N_6812);
nand U11116 (N_11116,N_7635,N_6637);
nor U11117 (N_11117,N_7014,N_8434);
or U11118 (N_11118,N_8411,N_8690);
and U11119 (N_11119,N_8095,N_8306);
or U11120 (N_11120,N_6206,N_6177);
or U11121 (N_11121,N_7525,N_6677);
or U11122 (N_11122,N_8836,N_7158);
or U11123 (N_11123,N_6607,N_8702);
or U11124 (N_11124,N_6784,N_7323);
or U11125 (N_11125,N_7257,N_8045);
or U11126 (N_11126,N_6544,N_8735);
or U11127 (N_11127,N_7591,N_7420);
nor U11128 (N_11128,N_6729,N_7936);
or U11129 (N_11129,N_8702,N_7821);
and U11130 (N_11130,N_8138,N_7278);
or U11131 (N_11131,N_6580,N_8854);
nand U11132 (N_11132,N_8653,N_6637);
nand U11133 (N_11133,N_7834,N_7315);
nor U11134 (N_11134,N_7499,N_7945);
nand U11135 (N_11135,N_7446,N_6216);
nand U11136 (N_11136,N_6101,N_7337);
nor U11137 (N_11137,N_6551,N_8530);
and U11138 (N_11138,N_6895,N_8316);
nand U11139 (N_11139,N_8599,N_6363);
nand U11140 (N_11140,N_6684,N_6802);
and U11141 (N_11141,N_6586,N_7886);
and U11142 (N_11142,N_8049,N_7452);
or U11143 (N_11143,N_6465,N_7448);
nor U11144 (N_11144,N_6739,N_8257);
xnor U11145 (N_11145,N_8434,N_6003);
and U11146 (N_11146,N_8425,N_6697);
and U11147 (N_11147,N_7026,N_7002);
nand U11148 (N_11148,N_6594,N_6266);
nand U11149 (N_11149,N_8981,N_8169);
nand U11150 (N_11150,N_6595,N_7553);
or U11151 (N_11151,N_6463,N_7990);
nor U11152 (N_11152,N_8235,N_6952);
and U11153 (N_11153,N_8183,N_6511);
or U11154 (N_11154,N_8868,N_6697);
or U11155 (N_11155,N_6969,N_7402);
or U11156 (N_11156,N_6375,N_8870);
and U11157 (N_11157,N_6855,N_6218);
and U11158 (N_11158,N_6368,N_6902);
and U11159 (N_11159,N_8883,N_6211);
nor U11160 (N_11160,N_7531,N_6164);
nand U11161 (N_11161,N_6909,N_6857);
nand U11162 (N_11162,N_8195,N_8052);
and U11163 (N_11163,N_8519,N_8788);
and U11164 (N_11164,N_6387,N_6356);
or U11165 (N_11165,N_7412,N_8520);
nor U11166 (N_11166,N_7848,N_8690);
nand U11167 (N_11167,N_6776,N_6252);
and U11168 (N_11168,N_6732,N_7307);
and U11169 (N_11169,N_6901,N_7547);
nor U11170 (N_11170,N_6681,N_6729);
nand U11171 (N_11171,N_6364,N_6775);
and U11172 (N_11172,N_8305,N_6132);
nand U11173 (N_11173,N_8655,N_7147);
nor U11174 (N_11174,N_7241,N_7589);
nor U11175 (N_11175,N_6378,N_6281);
or U11176 (N_11176,N_6970,N_8308);
nor U11177 (N_11177,N_7904,N_8302);
or U11178 (N_11178,N_7717,N_6644);
nand U11179 (N_11179,N_8087,N_6861);
nand U11180 (N_11180,N_8930,N_6091);
or U11181 (N_11181,N_6806,N_7087);
nand U11182 (N_11182,N_7949,N_8256);
nor U11183 (N_11183,N_7055,N_6915);
and U11184 (N_11184,N_8097,N_6516);
nand U11185 (N_11185,N_7892,N_6266);
nand U11186 (N_11186,N_6496,N_8441);
nor U11187 (N_11187,N_7640,N_8410);
or U11188 (N_11188,N_8299,N_7126);
and U11189 (N_11189,N_8016,N_7710);
nor U11190 (N_11190,N_6497,N_6485);
nand U11191 (N_11191,N_6120,N_8812);
nor U11192 (N_11192,N_8995,N_8090);
or U11193 (N_11193,N_8541,N_7228);
nor U11194 (N_11194,N_8481,N_6059);
nor U11195 (N_11195,N_8304,N_7597);
or U11196 (N_11196,N_8804,N_6493);
and U11197 (N_11197,N_6617,N_8583);
nand U11198 (N_11198,N_6630,N_7787);
and U11199 (N_11199,N_8054,N_7728);
or U11200 (N_11200,N_7081,N_8192);
or U11201 (N_11201,N_6511,N_8515);
or U11202 (N_11202,N_8537,N_6984);
or U11203 (N_11203,N_6245,N_6130);
and U11204 (N_11204,N_7853,N_8765);
nand U11205 (N_11205,N_6635,N_6380);
nor U11206 (N_11206,N_8053,N_8404);
nor U11207 (N_11207,N_7002,N_6904);
nand U11208 (N_11208,N_8154,N_8446);
nor U11209 (N_11209,N_7192,N_8443);
and U11210 (N_11210,N_6565,N_8930);
and U11211 (N_11211,N_8599,N_6108);
or U11212 (N_11212,N_6622,N_6020);
and U11213 (N_11213,N_7653,N_8371);
nand U11214 (N_11214,N_7608,N_8546);
and U11215 (N_11215,N_7323,N_8411);
and U11216 (N_11216,N_6432,N_7924);
or U11217 (N_11217,N_8319,N_6567);
and U11218 (N_11218,N_6738,N_7246);
nor U11219 (N_11219,N_6077,N_8541);
and U11220 (N_11220,N_7062,N_6951);
and U11221 (N_11221,N_7922,N_7950);
or U11222 (N_11222,N_8952,N_7261);
and U11223 (N_11223,N_7675,N_7852);
or U11224 (N_11224,N_8159,N_6535);
and U11225 (N_11225,N_7325,N_6889);
nand U11226 (N_11226,N_7489,N_6225);
nor U11227 (N_11227,N_8717,N_8364);
or U11228 (N_11228,N_7300,N_8432);
nor U11229 (N_11229,N_8080,N_6236);
and U11230 (N_11230,N_7336,N_6709);
or U11231 (N_11231,N_8144,N_6533);
nand U11232 (N_11232,N_7402,N_7522);
nor U11233 (N_11233,N_6180,N_8061);
or U11234 (N_11234,N_7213,N_8598);
nand U11235 (N_11235,N_7048,N_7314);
and U11236 (N_11236,N_7331,N_6465);
nand U11237 (N_11237,N_8672,N_8102);
and U11238 (N_11238,N_7489,N_8786);
nor U11239 (N_11239,N_8345,N_7279);
or U11240 (N_11240,N_7026,N_8781);
nand U11241 (N_11241,N_6079,N_8226);
nor U11242 (N_11242,N_8668,N_6308);
or U11243 (N_11243,N_6875,N_7113);
or U11244 (N_11244,N_7379,N_8389);
nand U11245 (N_11245,N_8409,N_6149);
or U11246 (N_11246,N_7497,N_6987);
and U11247 (N_11247,N_6040,N_6651);
or U11248 (N_11248,N_6070,N_7662);
nor U11249 (N_11249,N_7655,N_8694);
nand U11250 (N_11250,N_7373,N_7789);
nor U11251 (N_11251,N_8883,N_6759);
and U11252 (N_11252,N_6255,N_6007);
nor U11253 (N_11253,N_6714,N_6465);
or U11254 (N_11254,N_7629,N_8417);
nand U11255 (N_11255,N_6446,N_7098);
and U11256 (N_11256,N_8045,N_8719);
and U11257 (N_11257,N_7541,N_7116);
or U11258 (N_11258,N_6844,N_8164);
nand U11259 (N_11259,N_6508,N_8883);
and U11260 (N_11260,N_8634,N_6105);
and U11261 (N_11261,N_7632,N_8382);
nor U11262 (N_11262,N_7057,N_7794);
or U11263 (N_11263,N_8099,N_6267);
nand U11264 (N_11264,N_8501,N_8942);
or U11265 (N_11265,N_8610,N_6340);
nand U11266 (N_11266,N_7419,N_6632);
and U11267 (N_11267,N_7341,N_7471);
or U11268 (N_11268,N_6311,N_8661);
and U11269 (N_11269,N_6449,N_6274);
and U11270 (N_11270,N_7837,N_8319);
nand U11271 (N_11271,N_6292,N_7487);
and U11272 (N_11272,N_7495,N_7638);
nor U11273 (N_11273,N_6099,N_8121);
nor U11274 (N_11274,N_7928,N_7275);
and U11275 (N_11275,N_7110,N_7773);
nor U11276 (N_11276,N_6442,N_6938);
nor U11277 (N_11277,N_7647,N_6431);
or U11278 (N_11278,N_8372,N_7204);
nand U11279 (N_11279,N_7941,N_7015);
nor U11280 (N_11280,N_7867,N_8242);
nor U11281 (N_11281,N_6053,N_7153);
and U11282 (N_11282,N_7644,N_8087);
nand U11283 (N_11283,N_6891,N_8053);
and U11284 (N_11284,N_6865,N_8977);
nand U11285 (N_11285,N_7133,N_7195);
or U11286 (N_11286,N_7496,N_6758);
or U11287 (N_11287,N_8637,N_7050);
nor U11288 (N_11288,N_8435,N_7300);
nor U11289 (N_11289,N_8165,N_8188);
nand U11290 (N_11290,N_7899,N_6546);
or U11291 (N_11291,N_7482,N_6405);
nor U11292 (N_11292,N_6552,N_6321);
nand U11293 (N_11293,N_8633,N_7441);
or U11294 (N_11294,N_8991,N_7526);
nor U11295 (N_11295,N_8040,N_6365);
and U11296 (N_11296,N_7725,N_6780);
nand U11297 (N_11297,N_8645,N_7369);
nand U11298 (N_11298,N_8192,N_7216);
and U11299 (N_11299,N_6287,N_7650);
or U11300 (N_11300,N_6746,N_8453);
and U11301 (N_11301,N_7679,N_6229);
or U11302 (N_11302,N_6847,N_7409);
or U11303 (N_11303,N_6796,N_8430);
nor U11304 (N_11304,N_6591,N_8558);
or U11305 (N_11305,N_6824,N_6602);
nand U11306 (N_11306,N_7361,N_6105);
and U11307 (N_11307,N_6891,N_8507);
nand U11308 (N_11308,N_8132,N_6294);
and U11309 (N_11309,N_7354,N_7444);
and U11310 (N_11310,N_6920,N_8240);
nor U11311 (N_11311,N_8679,N_6659);
or U11312 (N_11312,N_8443,N_6615);
nand U11313 (N_11313,N_8436,N_6950);
nor U11314 (N_11314,N_7062,N_7742);
xor U11315 (N_11315,N_6386,N_8272);
and U11316 (N_11316,N_7204,N_6561);
nor U11317 (N_11317,N_7342,N_8111);
nor U11318 (N_11318,N_8111,N_6908);
nor U11319 (N_11319,N_6660,N_7067);
or U11320 (N_11320,N_8284,N_6401);
nand U11321 (N_11321,N_8956,N_8204);
and U11322 (N_11322,N_6290,N_7162);
and U11323 (N_11323,N_8495,N_8663);
or U11324 (N_11324,N_8135,N_8000);
nor U11325 (N_11325,N_6548,N_6293);
nor U11326 (N_11326,N_7649,N_7643);
nand U11327 (N_11327,N_7250,N_6348);
nor U11328 (N_11328,N_6058,N_6825);
and U11329 (N_11329,N_6221,N_6420);
nor U11330 (N_11330,N_8625,N_8781);
nand U11331 (N_11331,N_6649,N_6014);
and U11332 (N_11332,N_7473,N_8689);
or U11333 (N_11333,N_8789,N_7967);
nor U11334 (N_11334,N_6293,N_6752);
nor U11335 (N_11335,N_7159,N_8495);
nand U11336 (N_11336,N_8780,N_6861);
or U11337 (N_11337,N_7375,N_6843);
or U11338 (N_11338,N_6339,N_6010);
or U11339 (N_11339,N_7466,N_8221);
and U11340 (N_11340,N_6542,N_8163);
and U11341 (N_11341,N_7479,N_8701);
or U11342 (N_11342,N_6715,N_6472);
or U11343 (N_11343,N_6817,N_7245);
nor U11344 (N_11344,N_7059,N_6972);
nand U11345 (N_11345,N_6089,N_8130);
or U11346 (N_11346,N_8653,N_8592);
nand U11347 (N_11347,N_6615,N_8249);
nor U11348 (N_11348,N_7327,N_8133);
nand U11349 (N_11349,N_6130,N_6577);
nand U11350 (N_11350,N_6948,N_6340);
nand U11351 (N_11351,N_8143,N_7776);
or U11352 (N_11352,N_8392,N_8327);
or U11353 (N_11353,N_6507,N_7323);
and U11354 (N_11354,N_7133,N_7664);
or U11355 (N_11355,N_6558,N_7679);
nor U11356 (N_11356,N_7615,N_8899);
and U11357 (N_11357,N_8589,N_6627);
nor U11358 (N_11358,N_6134,N_8458);
nand U11359 (N_11359,N_8067,N_8837);
nand U11360 (N_11360,N_6189,N_6296);
and U11361 (N_11361,N_8387,N_6465);
nand U11362 (N_11362,N_6657,N_7939);
and U11363 (N_11363,N_7992,N_6250);
nand U11364 (N_11364,N_8397,N_6607);
nand U11365 (N_11365,N_8046,N_7665);
nand U11366 (N_11366,N_8580,N_6767);
or U11367 (N_11367,N_7976,N_7226);
or U11368 (N_11368,N_6550,N_8848);
or U11369 (N_11369,N_7423,N_7386);
and U11370 (N_11370,N_6652,N_7083);
nor U11371 (N_11371,N_6132,N_8481);
nor U11372 (N_11372,N_7538,N_8544);
nor U11373 (N_11373,N_8351,N_7751);
or U11374 (N_11374,N_8897,N_7907);
nor U11375 (N_11375,N_6022,N_8419);
nand U11376 (N_11376,N_7926,N_7757);
nor U11377 (N_11377,N_7250,N_6452);
nand U11378 (N_11378,N_6498,N_8395);
xnor U11379 (N_11379,N_8694,N_8597);
and U11380 (N_11380,N_8078,N_8248);
and U11381 (N_11381,N_8280,N_6517);
or U11382 (N_11382,N_6982,N_8544);
or U11383 (N_11383,N_8709,N_6969);
or U11384 (N_11384,N_7499,N_6703);
and U11385 (N_11385,N_8080,N_8286);
and U11386 (N_11386,N_7425,N_6402);
nand U11387 (N_11387,N_6445,N_8303);
xnor U11388 (N_11388,N_6687,N_8911);
nand U11389 (N_11389,N_8204,N_7749);
and U11390 (N_11390,N_8009,N_8353);
and U11391 (N_11391,N_8636,N_6983);
nor U11392 (N_11392,N_6449,N_7151);
or U11393 (N_11393,N_8336,N_8657);
nor U11394 (N_11394,N_8046,N_6111);
or U11395 (N_11395,N_6782,N_8708);
and U11396 (N_11396,N_7064,N_8429);
or U11397 (N_11397,N_6971,N_8739);
nor U11398 (N_11398,N_7141,N_7842);
and U11399 (N_11399,N_7794,N_6169);
or U11400 (N_11400,N_7082,N_7560);
nor U11401 (N_11401,N_7794,N_6510);
and U11402 (N_11402,N_8263,N_6843);
or U11403 (N_11403,N_7638,N_6001);
nor U11404 (N_11404,N_8400,N_7272);
nor U11405 (N_11405,N_7335,N_7447);
or U11406 (N_11406,N_6785,N_7453);
nand U11407 (N_11407,N_6173,N_8664);
nand U11408 (N_11408,N_8855,N_6426);
nand U11409 (N_11409,N_7765,N_8586);
and U11410 (N_11410,N_6978,N_7892);
and U11411 (N_11411,N_7418,N_8685);
nand U11412 (N_11412,N_6203,N_6111);
or U11413 (N_11413,N_8052,N_8341);
nand U11414 (N_11414,N_8295,N_6762);
and U11415 (N_11415,N_7114,N_8908);
nand U11416 (N_11416,N_8910,N_8827);
and U11417 (N_11417,N_7757,N_7065);
and U11418 (N_11418,N_7828,N_7343);
or U11419 (N_11419,N_7238,N_6996);
and U11420 (N_11420,N_8914,N_8167);
or U11421 (N_11421,N_7035,N_7736);
nor U11422 (N_11422,N_7371,N_8392);
nand U11423 (N_11423,N_6542,N_7766);
or U11424 (N_11424,N_6222,N_7094);
and U11425 (N_11425,N_8454,N_7804);
nand U11426 (N_11426,N_7174,N_7709);
nand U11427 (N_11427,N_8339,N_7668);
nand U11428 (N_11428,N_8087,N_7733);
or U11429 (N_11429,N_6865,N_6924);
nand U11430 (N_11430,N_8596,N_6118);
and U11431 (N_11431,N_7163,N_7176);
or U11432 (N_11432,N_8079,N_8944);
nand U11433 (N_11433,N_8123,N_6755);
and U11434 (N_11434,N_8213,N_7108);
nand U11435 (N_11435,N_8764,N_7371);
or U11436 (N_11436,N_7177,N_6032);
or U11437 (N_11437,N_8928,N_7319);
nor U11438 (N_11438,N_8784,N_7495);
and U11439 (N_11439,N_8660,N_6259);
or U11440 (N_11440,N_6858,N_7153);
nor U11441 (N_11441,N_7244,N_8224);
nor U11442 (N_11442,N_7702,N_6401);
nand U11443 (N_11443,N_6845,N_6046);
and U11444 (N_11444,N_7370,N_8250);
and U11445 (N_11445,N_6463,N_7366);
nor U11446 (N_11446,N_8989,N_7052);
or U11447 (N_11447,N_8994,N_8178);
and U11448 (N_11448,N_8688,N_6959);
or U11449 (N_11449,N_8200,N_7011);
and U11450 (N_11450,N_6802,N_7236);
nand U11451 (N_11451,N_7854,N_7133);
nor U11452 (N_11452,N_6170,N_8954);
nand U11453 (N_11453,N_7605,N_7990);
or U11454 (N_11454,N_8830,N_6883);
and U11455 (N_11455,N_7456,N_7910);
nand U11456 (N_11456,N_8047,N_7158);
or U11457 (N_11457,N_6674,N_6656);
xnor U11458 (N_11458,N_7165,N_7415);
nand U11459 (N_11459,N_7400,N_6996);
nor U11460 (N_11460,N_8675,N_7098);
nor U11461 (N_11461,N_6442,N_7524);
nor U11462 (N_11462,N_8083,N_8627);
and U11463 (N_11463,N_7206,N_7185);
xnor U11464 (N_11464,N_6764,N_7592);
nand U11465 (N_11465,N_8990,N_8356);
nor U11466 (N_11466,N_8285,N_7730);
or U11467 (N_11467,N_8778,N_8701);
nor U11468 (N_11468,N_6401,N_7007);
and U11469 (N_11469,N_6831,N_6051);
nor U11470 (N_11470,N_6835,N_7741);
nand U11471 (N_11471,N_8332,N_6482);
nor U11472 (N_11472,N_7063,N_8734);
nor U11473 (N_11473,N_7950,N_6767);
and U11474 (N_11474,N_7975,N_8242);
or U11475 (N_11475,N_7039,N_7140);
nor U11476 (N_11476,N_7364,N_6406);
and U11477 (N_11477,N_6653,N_7221);
and U11478 (N_11478,N_8564,N_8630);
nand U11479 (N_11479,N_7945,N_6371);
or U11480 (N_11480,N_8100,N_8179);
nor U11481 (N_11481,N_8822,N_6762);
and U11482 (N_11482,N_6437,N_6842);
nand U11483 (N_11483,N_7129,N_7389);
nand U11484 (N_11484,N_6390,N_6128);
nand U11485 (N_11485,N_8299,N_8339);
and U11486 (N_11486,N_7803,N_6169);
or U11487 (N_11487,N_6401,N_8343);
or U11488 (N_11488,N_7870,N_6042);
or U11489 (N_11489,N_7947,N_7967);
xnor U11490 (N_11490,N_6053,N_7901);
nor U11491 (N_11491,N_8069,N_7770);
nor U11492 (N_11492,N_7756,N_7066);
and U11493 (N_11493,N_6862,N_6649);
nand U11494 (N_11494,N_6286,N_8319);
or U11495 (N_11495,N_6470,N_7025);
and U11496 (N_11496,N_8817,N_8836);
and U11497 (N_11497,N_6417,N_6614);
nor U11498 (N_11498,N_8640,N_7561);
nand U11499 (N_11499,N_7292,N_6909);
nor U11500 (N_11500,N_6135,N_6200);
nor U11501 (N_11501,N_7498,N_8137);
nand U11502 (N_11502,N_8393,N_7655);
or U11503 (N_11503,N_6889,N_8145);
nor U11504 (N_11504,N_7524,N_8869);
and U11505 (N_11505,N_7570,N_8112);
nand U11506 (N_11506,N_7025,N_6723);
and U11507 (N_11507,N_8365,N_6233);
or U11508 (N_11508,N_8800,N_8669);
nand U11509 (N_11509,N_6860,N_8193);
and U11510 (N_11510,N_6413,N_8182);
and U11511 (N_11511,N_7756,N_8057);
nor U11512 (N_11512,N_6529,N_8390);
nor U11513 (N_11513,N_7956,N_6298);
nor U11514 (N_11514,N_8857,N_6016);
and U11515 (N_11515,N_6141,N_6636);
nand U11516 (N_11516,N_6861,N_8145);
nand U11517 (N_11517,N_7143,N_7878);
nand U11518 (N_11518,N_7499,N_7820);
nand U11519 (N_11519,N_8655,N_6552);
nor U11520 (N_11520,N_6010,N_8902);
or U11521 (N_11521,N_7275,N_6537);
nand U11522 (N_11522,N_8778,N_7070);
nand U11523 (N_11523,N_7526,N_7528);
nor U11524 (N_11524,N_7788,N_6049);
nand U11525 (N_11525,N_8041,N_7010);
nand U11526 (N_11526,N_8450,N_8447);
nor U11527 (N_11527,N_8095,N_7818);
nor U11528 (N_11528,N_7953,N_7064);
or U11529 (N_11529,N_8202,N_6695);
and U11530 (N_11530,N_8677,N_7230);
or U11531 (N_11531,N_6560,N_7095);
nor U11532 (N_11532,N_8688,N_7565);
and U11533 (N_11533,N_7129,N_8111);
and U11534 (N_11534,N_7127,N_6438);
nand U11535 (N_11535,N_7135,N_8975);
and U11536 (N_11536,N_8816,N_7463);
or U11537 (N_11537,N_8216,N_8694);
nor U11538 (N_11538,N_7329,N_6535);
nor U11539 (N_11539,N_8469,N_6983);
nand U11540 (N_11540,N_6915,N_6555);
or U11541 (N_11541,N_7992,N_7486);
or U11542 (N_11542,N_7010,N_7466);
or U11543 (N_11543,N_7364,N_7283);
or U11544 (N_11544,N_8625,N_6407);
nor U11545 (N_11545,N_6248,N_7262);
nand U11546 (N_11546,N_6281,N_8826);
nor U11547 (N_11547,N_7238,N_8818);
nand U11548 (N_11548,N_8817,N_7344);
nor U11549 (N_11549,N_6574,N_7854);
or U11550 (N_11550,N_8225,N_7510);
and U11551 (N_11551,N_7954,N_7090);
or U11552 (N_11552,N_8838,N_6426);
or U11553 (N_11553,N_6072,N_8816);
or U11554 (N_11554,N_6704,N_8227);
nand U11555 (N_11555,N_7236,N_6098);
or U11556 (N_11556,N_8678,N_7353);
nand U11557 (N_11557,N_7723,N_6876);
nor U11558 (N_11558,N_8573,N_8633);
and U11559 (N_11559,N_8329,N_7268);
nor U11560 (N_11560,N_7639,N_6926);
nand U11561 (N_11561,N_8961,N_6990);
or U11562 (N_11562,N_6529,N_7759);
nor U11563 (N_11563,N_6486,N_6829);
nor U11564 (N_11564,N_6789,N_6258);
and U11565 (N_11565,N_8060,N_6647);
nand U11566 (N_11566,N_6310,N_7521);
nand U11567 (N_11567,N_7041,N_8585);
nor U11568 (N_11568,N_8337,N_7006);
nand U11569 (N_11569,N_6770,N_8887);
or U11570 (N_11570,N_8611,N_6360);
or U11571 (N_11571,N_8833,N_6438);
xnor U11572 (N_11572,N_6672,N_7254);
nor U11573 (N_11573,N_8736,N_8868);
and U11574 (N_11574,N_7570,N_7239);
and U11575 (N_11575,N_7237,N_8946);
or U11576 (N_11576,N_6949,N_7912);
or U11577 (N_11577,N_7560,N_7933);
nor U11578 (N_11578,N_7776,N_7566);
and U11579 (N_11579,N_6296,N_8027);
and U11580 (N_11580,N_8972,N_6364);
nor U11581 (N_11581,N_7926,N_8554);
or U11582 (N_11582,N_7298,N_8273);
or U11583 (N_11583,N_8823,N_8054);
and U11584 (N_11584,N_8599,N_7206);
nor U11585 (N_11585,N_8242,N_6048);
or U11586 (N_11586,N_6488,N_7368);
nand U11587 (N_11587,N_6027,N_8774);
nor U11588 (N_11588,N_7448,N_7087);
or U11589 (N_11589,N_7754,N_7457);
xnor U11590 (N_11590,N_6755,N_6063);
and U11591 (N_11591,N_8688,N_8490);
and U11592 (N_11592,N_8607,N_8458);
nand U11593 (N_11593,N_6380,N_7328);
and U11594 (N_11594,N_6962,N_8602);
nand U11595 (N_11595,N_7565,N_7881);
or U11596 (N_11596,N_7194,N_6922);
nor U11597 (N_11597,N_7976,N_7283);
nand U11598 (N_11598,N_7608,N_7292);
or U11599 (N_11599,N_8852,N_7503);
and U11600 (N_11600,N_7705,N_6457);
or U11601 (N_11601,N_6545,N_6879);
nor U11602 (N_11602,N_7783,N_8295);
or U11603 (N_11603,N_7394,N_6271);
nand U11604 (N_11604,N_8146,N_7012);
and U11605 (N_11605,N_6279,N_6503);
and U11606 (N_11606,N_8080,N_6131);
or U11607 (N_11607,N_8774,N_6387);
nor U11608 (N_11608,N_7631,N_8764);
nand U11609 (N_11609,N_7922,N_6673);
nor U11610 (N_11610,N_7049,N_7852);
nand U11611 (N_11611,N_6892,N_7807);
nand U11612 (N_11612,N_6407,N_8183);
nand U11613 (N_11613,N_7543,N_6703);
nor U11614 (N_11614,N_6212,N_6386);
nand U11615 (N_11615,N_7775,N_6258);
nor U11616 (N_11616,N_7156,N_7175);
or U11617 (N_11617,N_6862,N_6973);
or U11618 (N_11618,N_6190,N_6207);
nand U11619 (N_11619,N_7765,N_8360);
nor U11620 (N_11620,N_6600,N_7281);
or U11621 (N_11621,N_7718,N_6262);
nand U11622 (N_11622,N_6757,N_8357);
and U11623 (N_11623,N_6449,N_7903);
nand U11624 (N_11624,N_6684,N_8416);
nor U11625 (N_11625,N_6409,N_7320);
nor U11626 (N_11626,N_6499,N_6751);
nand U11627 (N_11627,N_6838,N_6678);
and U11628 (N_11628,N_6651,N_8949);
nor U11629 (N_11629,N_8324,N_7495);
nand U11630 (N_11630,N_8478,N_7535);
and U11631 (N_11631,N_8822,N_8485);
and U11632 (N_11632,N_8010,N_7621);
nor U11633 (N_11633,N_7372,N_7681);
or U11634 (N_11634,N_6345,N_7434);
nand U11635 (N_11635,N_7274,N_8074);
nand U11636 (N_11636,N_6506,N_8057);
nand U11637 (N_11637,N_8977,N_8547);
nor U11638 (N_11638,N_6237,N_6408);
nor U11639 (N_11639,N_7870,N_8952);
and U11640 (N_11640,N_8226,N_8280);
or U11641 (N_11641,N_7530,N_8410);
and U11642 (N_11642,N_6007,N_6477);
nor U11643 (N_11643,N_6962,N_8503);
or U11644 (N_11644,N_8868,N_6813);
xor U11645 (N_11645,N_7752,N_7614);
and U11646 (N_11646,N_8627,N_7515);
nor U11647 (N_11647,N_7130,N_6328);
nand U11648 (N_11648,N_8290,N_7976);
and U11649 (N_11649,N_8342,N_8174);
or U11650 (N_11650,N_7976,N_6288);
and U11651 (N_11651,N_6812,N_8311);
or U11652 (N_11652,N_6034,N_6267);
and U11653 (N_11653,N_8608,N_7000);
nand U11654 (N_11654,N_8347,N_7063);
nor U11655 (N_11655,N_7968,N_7878);
or U11656 (N_11656,N_8132,N_7906);
nor U11657 (N_11657,N_8895,N_6657);
and U11658 (N_11658,N_6117,N_7845);
nand U11659 (N_11659,N_6253,N_7300);
or U11660 (N_11660,N_7826,N_6201);
nand U11661 (N_11661,N_6403,N_6643);
nand U11662 (N_11662,N_7202,N_8415);
nand U11663 (N_11663,N_6511,N_8008);
xor U11664 (N_11664,N_6396,N_7105);
or U11665 (N_11665,N_6336,N_6582);
and U11666 (N_11666,N_7788,N_6835);
or U11667 (N_11667,N_7435,N_8687);
nand U11668 (N_11668,N_6703,N_8142);
or U11669 (N_11669,N_6153,N_6429);
or U11670 (N_11670,N_6396,N_8421);
nor U11671 (N_11671,N_7459,N_7483);
and U11672 (N_11672,N_7660,N_6280);
xor U11673 (N_11673,N_6437,N_7463);
nand U11674 (N_11674,N_6056,N_6859);
and U11675 (N_11675,N_8844,N_6355);
and U11676 (N_11676,N_6667,N_6110);
or U11677 (N_11677,N_7712,N_6071);
and U11678 (N_11678,N_6560,N_8537);
or U11679 (N_11679,N_7847,N_6499);
nand U11680 (N_11680,N_6995,N_8006);
and U11681 (N_11681,N_8855,N_8030);
nor U11682 (N_11682,N_7105,N_6571);
or U11683 (N_11683,N_6298,N_6462);
and U11684 (N_11684,N_7216,N_6585);
or U11685 (N_11685,N_6453,N_6634);
and U11686 (N_11686,N_7352,N_8566);
or U11687 (N_11687,N_6001,N_8243);
or U11688 (N_11688,N_6076,N_6719);
and U11689 (N_11689,N_8110,N_7043);
or U11690 (N_11690,N_8279,N_8223);
nor U11691 (N_11691,N_6810,N_7422);
or U11692 (N_11692,N_7482,N_7157);
nand U11693 (N_11693,N_6532,N_7002);
nor U11694 (N_11694,N_6494,N_8040);
and U11695 (N_11695,N_7529,N_7934);
or U11696 (N_11696,N_7456,N_7540);
xor U11697 (N_11697,N_6186,N_8932);
nor U11698 (N_11698,N_8478,N_6268);
or U11699 (N_11699,N_8978,N_6576);
nand U11700 (N_11700,N_7768,N_6004);
and U11701 (N_11701,N_6688,N_7925);
or U11702 (N_11702,N_6861,N_8700);
nor U11703 (N_11703,N_6693,N_6501);
nor U11704 (N_11704,N_8850,N_6132);
or U11705 (N_11705,N_6339,N_6323);
nor U11706 (N_11706,N_8686,N_8536);
or U11707 (N_11707,N_8359,N_6348);
xor U11708 (N_11708,N_7349,N_8258);
or U11709 (N_11709,N_6626,N_8798);
and U11710 (N_11710,N_7731,N_6918);
nand U11711 (N_11711,N_8595,N_7860);
or U11712 (N_11712,N_6278,N_8744);
nand U11713 (N_11713,N_6531,N_8740);
and U11714 (N_11714,N_6589,N_8957);
nor U11715 (N_11715,N_8910,N_6571);
nor U11716 (N_11716,N_7791,N_7582);
or U11717 (N_11717,N_7164,N_7789);
or U11718 (N_11718,N_7891,N_7948);
nor U11719 (N_11719,N_8477,N_7186);
and U11720 (N_11720,N_7361,N_8240);
and U11721 (N_11721,N_6384,N_8004);
nor U11722 (N_11722,N_6228,N_7331);
nor U11723 (N_11723,N_8242,N_7006);
and U11724 (N_11724,N_6242,N_8532);
or U11725 (N_11725,N_6236,N_7821);
and U11726 (N_11726,N_7013,N_6784);
nand U11727 (N_11727,N_6989,N_8493);
nand U11728 (N_11728,N_8259,N_7929);
nand U11729 (N_11729,N_6795,N_8517);
nand U11730 (N_11730,N_7686,N_8704);
nand U11731 (N_11731,N_6781,N_7960);
and U11732 (N_11732,N_8226,N_6677);
nand U11733 (N_11733,N_6203,N_6544);
xnor U11734 (N_11734,N_6649,N_6172);
and U11735 (N_11735,N_6935,N_7681);
nor U11736 (N_11736,N_7116,N_6896);
or U11737 (N_11737,N_7591,N_6850);
and U11738 (N_11738,N_7492,N_6565);
nor U11739 (N_11739,N_8118,N_8677);
nand U11740 (N_11740,N_7497,N_7593);
nor U11741 (N_11741,N_8032,N_8319);
and U11742 (N_11742,N_7947,N_6157);
or U11743 (N_11743,N_6430,N_7192);
xnor U11744 (N_11744,N_6506,N_6578);
or U11745 (N_11745,N_8187,N_8337);
nand U11746 (N_11746,N_8909,N_7018);
and U11747 (N_11747,N_7159,N_8605);
nand U11748 (N_11748,N_6903,N_6291);
or U11749 (N_11749,N_8999,N_6978);
or U11750 (N_11750,N_8635,N_8294);
nor U11751 (N_11751,N_7189,N_6548);
or U11752 (N_11752,N_6762,N_6876);
and U11753 (N_11753,N_7242,N_6535);
nor U11754 (N_11754,N_8117,N_6996);
or U11755 (N_11755,N_7221,N_8752);
and U11756 (N_11756,N_8668,N_8671);
and U11757 (N_11757,N_6457,N_8354);
or U11758 (N_11758,N_6284,N_6048);
nor U11759 (N_11759,N_6090,N_6073);
nor U11760 (N_11760,N_6464,N_8212);
and U11761 (N_11761,N_8304,N_7646);
and U11762 (N_11762,N_7493,N_6590);
or U11763 (N_11763,N_8280,N_8485);
or U11764 (N_11764,N_7359,N_7029);
nor U11765 (N_11765,N_6399,N_6901);
and U11766 (N_11766,N_7808,N_8869);
nor U11767 (N_11767,N_8683,N_7958);
nor U11768 (N_11768,N_8671,N_6699);
and U11769 (N_11769,N_8653,N_7378);
nor U11770 (N_11770,N_8077,N_7941);
nor U11771 (N_11771,N_7544,N_8675);
and U11772 (N_11772,N_7551,N_8906);
or U11773 (N_11773,N_6761,N_6841);
or U11774 (N_11774,N_7151,N_6208);
and U11775 (N_11775,N_6819,N_6029);
and U11776 (N_11776,N_7679,N_7194);
nand U11777 (N_11777,N_8046,N_8786);
or U11778 (N_11778,N_8970,N_8639);
and U11779 (N_11779,N_7245,N_7971);
and U11780 (N_11780,N_7779,N_6901);
or U11781 (N_11781,N_7097,N_6885);
or U11782 (N_11782,N_7656,N_7807);
and U11783 (N_11783,N_7719,N_6196);
nand U11784 (N_11784,N_8311,N_8533);
nor U11785 (N_11785,N_8754,N_8692);
nor U11786 (N_11786,N_8741,N_6010);
xnor U11787 (N_11787,N_6026,N_6310);
nor U11788 (N_11788,N_7047,N_6962);
and U11789 (N_11789,N_6185,N_8712);
or U11790 (N_11790,N_7969,N_8562);
and U11791 (N_11791,N_7974,N_8926);
and U11792 (N_11792,N_8888,N_8880);
and U11793 (N_11793,N_7244,N_6725);
xor U11794 (N_11794,N_6267,N_8787);
and U11795 (N_11795,N_8419,N_7277);
or U11796 (N_11796,N_6846,N_6169);
or U11797 (N_11797,N_6067,N_7340);
and U11798 (N_11798,N_7456,N_8231);
and U11799 (N_11799,N_6633,N_8320);
nand U11800 (N_11800,N_7712,N_6630);
nand U11801 (N_11801,N_7763,N_6159);
xnor U11802 (N_11802,N_7062,N_7246);
and U11803 (N_11803,N_8826,N_7697);
nor U11804 (N_11804,N_6489,N_7191);
nor U11805 (N_11805,N_6809,N_7041);
or U11806 (N_11806,N_6975,N_7462);
and U11807 (N_11807,N_8957,N_6006);
and U11808 (N_11808,N_7069,N_7845);
and U11809 (N_11809,N_7552,N_6390);
or U11810 (N_11810,N_8862,N_8036);
or U11811 (N_11811,N_7695,N_6883);
nand U11812 (N_11812,N_8462,N_8658);
nand U11813 (N_11813,N_8604,N_6049);
nor U11814 (N_11814,N_6476,N_8939);
nor U11815 (N_11815,N_7107,N_6957);
and U11816 (N_11816,N_7829,N_8630);
and U11817 (N_11817,N_6621,N_8913);
or U11818 (N_11818,N_6792,N_8746);
and U11819 (N_11819,N_7502,N_7550);
xor U11820 (N_11820,N_6046,N_8280);
and U11821 (N_11821,N_7956,N_8643);
nor U11822 (N_11822,N_7738,N_6301);
nand U11823 (N_11823,N_8335,N_7399);
or U11824 (N_11824,N_6992,N_8049);
or U11825 (N_11825,N_8369,N_8476);
nor U11826 (N_11826,N_6513,N_7278);
nor U11827 (N_11827,N_8644,N_8163);
nand U11828 (N_11828,N_8309,N_6061);
nor U11829 (N_11829,N_6083,N_8637);
nor U11830 (N_11830,N_6025,N_6495);
nor U11831 (N_11831,N_8141,N_6768);
nand U11832 (N_11832,N_6290,N_7062);
nor U11833 (N_11833,N_7435,N_7633);
nand U11834 (N_11834,N_8750,N_6737);
nor U11835 (N_11835,N_8509,N_8365);
or U11836 (N_11836,N_7203,N_8541);
nor U11837 (N_11837,N_8054,N_6728);
and U11838 (N_11838,N_6307,N_7674);
or U11839 (N_11839,N_8907,N_7865);
and U11840 (N_11840,N_6221,N_8741);
and U11841 (N_11841,N_7937,N_6673);
nand U11842 (N_11842,N_8167,N_6812);
and U11843 (N_11843,N_7556,N_6358);
or U11844 (N_11844,N_7595,N_7235);
and U11845 (N_11845,N_8473,N_6511);
or U11846 (N_11846,N_7481,N_6192);
nand U11847 (N_11847,N_6521,N_7636);
and U11848 (N_11848,N_7842,N_6162);
and U11849 (N_11849,N_7263,N_8734);
and U11850 (N_11850,N_6712,N_6506);
nand U11851 (N_11851,N_8268,N_8556);
and U11852 (N_11852,N_7810,N_8586);
and U11853 (N_11853,N_8971,N_7667);
nor U11854 (N_11854,N_6382,N_8519);
nand U11855 (N_11855,N_8742,N_7057);
nor U11856 (N_11856,N_8039,N_6381);
nor U11857 (N_11857,N_6789,N_6795);
nor U11858 (N_11858,N_7460,N_7334);
nand U11859 (N_11859,N_7525,N_8068);
or U11860 (N_11860,N_7569,N_6354);
nand U11861 (N_11861,N_6164,N_8758);
or U11862 (N_11862,N_7812,N_7911);
nand U11863 (N_11863,N_8306,N_6058);
and U11864 (N_11864,N_8305,N_8099);
nand U11865 (N_11865,N_6932,N_6760);
nand U11866 (N_11866,N_6952,N_7085);
nand U11867 (N_11867,N_7202,N_7152);
nand U11868 (N_11868,N_8471,N_6896);
nor U11869 (N_11869,N_8210,N_7955);
xor U11870 (N_11870,N_8879,N_7011);
nand U11871 (N_11871,N_8348,N_7597);
and U11872 (N_11872,N_7316,N_7799);
and U11873 (N_11873,N_6497,N_8302);
nand U11874 (N_11874,N_7506,N_7991);
or U11875 (N_11875,N_8655,N_8133);
nand U11876 (N_11876,N_6328,N_6073);
nor U11877 (N_11877,N_8175,N_6594);
or U11878 (N_11878,N_6366,N_6615);
nand U11879 (N_11879,N_8002,N_7372);
or U11880 (N_11880,N_7325,N_8308);
nor U11881 (N_11881,N_6412,N_7422);
nand U11882 (N_11882,N_7538,N_6872);
or U11883 (N_11883,N_8562,N_6773);
nor U11884 (N_11884,N_7510,N_8349);
or U11885 (N_11885,N_7983,N_7006);
nand U11886 (N_11886,N_8570,N_8493);
or U11887 (N_11887,N_7424,N_8662);
and U11888 (N_11888,N_8482,N_6724);
and U11889 (N_11889,N_6093,N_8466);
or U11890 (N_11890,N_8725,N_7463);
nand U11891 (N_11891,N_8437,N_6184);
and U11892 (N_11892,N_6192,N_7928);
nor U11893 (N_11893,N_7394,N_8592);
nor U11894 (N_11894,N_7732,N_7997);
and U11895 (N_11895,N_8631,N_8444);
or U11896 (N_11896,N_7221,N_7057);
nor U11897 (N_11897,N_8173,N_6223);
nand U11898 (N_11898,N_6619,N_7003);
nand U11899 (N_11899,N_7614,N_6075);
nand U11900 (N_11900,N_7307,N_6866);
and U11901 (N_11901,N_7084,N_8458);
nand U11902 (N_11902,N_8422,N_6923);
and U11903 (N_11903,N_6508,N_6141);
or U11904 (N_11904,N_8869,N_8457);
and U11905 (N_11905,N_6487,N_8860);
nand U11906 (N_11906,N_8061,N_8636);
and U11907 (N_11907,N_6083,N_6432);
nand U11908 (N_11908,N_8818,N_6840);
or U11909 (N_11909,N_7106,N_7377);
xnor U11910 (N_11910,N_6293,N_6007);
xnor U11911 (N_11911,N_7519,N_7994);
and U11912 (N_11912,N_7565,N_6332);
nand U11913 (N_11913,N_7855,N_7156);
or U11914 (N_11914,N_8470,N_7861);
and U11915 (N_11915,N_6052,N_8477);
xnor U11916 (N_11916,N_7360,N_7692);
and U11917 (N_11917,N_7046,N_7536);
nor U11918 (N_11918,N_8282,N_8638);
nand U11919 (N_11919,N_7221,N_7997);
or U11920 (N_11920,N_8279,N_8609);
and U11921 (N_11921,N_7482,N_7168);
nand U11922 (N_11922,N_6001,N_6906);
nor U11923 (N_11923,N_6401,N_6974);
nor U11924 (N_11924,N_8273,N_6226);
nor U11925 (N_11925,N_7440,N_7684);
nor U11926 (N_11926,N_8416,N_8260);
and U11927 (N_11927,N_8769,N_6618);
nand U11928 (N_11928,N_8688,N_8634);
or U11929 (N_11929,N_7394,N_7781);
nor U11930 (N_11930,N_7467,N_6980);
and U11931 (N_11931,N_7976,N_7609);
or U11932 (N_11932,N_8099,N_7711);
nand U11933 (N_11933,N_8163,N_6241);
nor U11934 (N_11934,N_6475,N_6219);
or U11935 (N_11935,N_6541,N_7646);
or U11936 (N_11936,N_6682,N_6537);
and U11937 (N_11937,N_8566,N_6584);
nor U11938 (N_11938,N_6665,N_6236);
nand U11939 (N_11939,N_6805,N_8854);
nor U11940 (N_11940,N_7860,N_6870);
nor U11941 (N_11941,N_7129,N_6241);
nand U11942 (N_11942,N_6938,N_8529);
and U11943 (N_11943,N_6052,N_7738);
or U11944 (N_11944,N_8516,N_7250);
nand U11945 (N_11945,N_8861,N_8925);
nand U11946 (N_11946,N_6855,N_8157);
or U11947 (N_11947,N_6588,N_8673);
and U11948 (N_11948,N_8607,N_6563);
and U11949 (N_11949,N_7690,N_7077);
or U11950 (N_11950,N_7206,N_7168);
nor U11951 (N_11951,N_6703,N_6967);
or U11952 (N_11952,N_6124,N_8412);
and U11953 (N_11953,N_8433,N_7643);
nor U11954 (N_11954,N_7590,N_8308);
or U11955 (N_11955,N_8410,N_8201);
or U11956 (N_11956,N_7308,N_6761);
and U11957 (N_11957,N_7936,N_7944);
and U11958 (N_11958,N_6446,N_6716);
nor U11959 (N_11959,N_7275,N_7343);
or U11960 (N_11960,N_8894,N_8746);
nand U11961 (N_11961,N_6233,N_6035);
or U11962 (N_11962,N_7561,N_8966);
and U11963 (N_11963,N_7409,N_6517);
nor U11964 (N_11964,N_7966,N_8710);
xnor U11965 (N_11965,N_7525,N_7697);
nor U11966 (N_11966,N_6614,N_8561);
nor U11967 (N_11967,N_7252,N_7643);
nor U11968 (N_11968,N_6216,N_6987);
nand U11969 (N_11969,N_7959,N_8768);
and U11970 (N_11970,N_6030,N_7720);
and U11971 (N_11971,N_6542,N_7193);
and U11972 (N_11972,N_7704,N_6888);
or U11973 (N_11973,N_6496,N_8216);
or U11974 (N_11974,N_6990,N_7012);
nand U11975 (N_11975,N_6903,N_8297);
nor U11976 (N_11976,N_6590,N_7150);
nor U11977 (N_11977,N_6679,N_7117);
and U11978 (N_11978,N_6815,N_6567);
nand U11979 (N_11979,N_7958,N_8574);
or U11980 (N_11980,N_6380,N_6834);
and U11981 (N_11981,N_6980,N_7721);
and U11982 (N_11982,N_7449,N_6771);
or U11983 (N_11983,N_7333,N_8858);
nor U11984 (N_11984,N_7730,N_8282);
nand U11985 (N_11985,N_6498,N_7207);
or U11986 (N_11986,N_6441,N_8527);
nor U11987 (N_11987,N_8196,N_6898);
nor U11988 (N_11988,N_8826,N_6669);
nor U11989 (N_11989,N_8034,N_8592);
nor U11990 (N_11990,N_8954,N_8678);
or U11991 (N_11991,N_6525,N_7100);
nand U11992 (N_11992,N_6206,N_6933);
nor U11993 (N_11993,N_6951,N_6530);
nand U11994 (N_11994,N_7559,N_7476);
nand U11995 (N_11995,N_6467,N_8777);
or U11996 (N_11996,N_8050,N_7009);
nor U11997 (N_11997,N_8075,N_8973);
nor U11998 (N_11998,N_7806,N_8425);
nand U11999 (N_11999,N_6674,N_6595);
nor U12000 (N_12000,N_9530,N_9893);
nand U12001 (N_12001,N_11146,N_11773);
or U12002 (N_12002,N_10714,N_9401);
or U12003 (N_12003,N_10870,N_10263);
or U12004 (N_12004,N_9286,N_11030);
nand U12005 (N_12005,N_11778,N_10594);
or U12006 (N_12006,N_10636,N_11798);
or U12007 (N_12007,N_11581,N_11749);
nand U12008 (N_12008,N_11683,N_9880);
nor U12009 (N_12009,N_11110,N_9715);
nand U12010 (N_12010,N_11973,N_9967);
or U12011 (N_12011,N_9537,N_10847);
and U12012 (N_12012,N_10293,N_10166);
nand U12013 (N_12013,N_9483,N_10030);
nor U12014 (N_12014,N_11547,N_11682);
and U12015 (N_12015,N_9691,N_10027);
and U12016 (N_12016,N_10015,N_10734);
nand U12017 (N_12017,N_11212,N_10444);
or U12018 (N_12018,N_10508,N_11584);
or U12019 (N_12019,N_11236,N_9885);
nand U12020 (N_12020,N_10695,N_11366);
nor U12021 (N_12021,N_9550,N_10253);
nor U12022 (N_12022,N_10958,N_10597);
nand U12023 (N_12023,N_10850,N_11566);
nor U12024 (N_12024,N_11887,N_10001);
or U12025 (N_12025,N_11324,N_9037);
nand U12026 (N_12026,N_10837,N_11823);
or U12027 (N_12027,N_9130,N_11949);
and U12028 (N_12028,N_11830,N_11619);
nand U12029 (N_12029,N_10688,N_9134);
nand U12030 (N_12030,N_9342,N_9190);
nor U12031 (N_12031,N_11289,N_10407);
nor U12032 (N_12032,N_11158,N_9036);
nand U12033 (N_12033,N_9090,N_11608);
nand U12034 (N_12034,N_10338,N_9437);
and U12035 (N_12035,N_9093,N_9380);
or U12036 (N_12036,N_11684,N_10925);
or U12037 (N_12037,N_10484,N_11803);
or U12038 (N_12038,N_10894,N_10178);
nand U12039 (N_12039,N_11609,N_10254);
nand U12040 (N_12040,N_9433,N_11101);
nand U12041 (N_12041,N_9317,N_9923);
nand U12042 (N_12042,N_11771,N_9259);
nor U12043 (N_12043,N_9235,N_11863);
nor U12044 (N_12044,N_11148,N_11415);
or U12045 (N_12045,N_10219,N_10247);
or U12046 (N_12046,N_11482,N_11718);
nand U12047 (N_12047,N_10327,N_11859);
nor U12048 (N_12048,N_11067,N_11042);
nand U12049 (N_12049,N_9770,N_11210);
or U12050 (N_12050,N_11019,N_9646);
or U12051 (N_12051,N_9170,N_11669);
nand U12052 (N_12052,N_10693,N_9898);
and U12053 (N_12053,N_11967,N_10056);
nand U12054 (N_12054,N_9132,N_10857);
or U12055 (N_12055,N_10835,N_10377);
or U12056 (N_12056,N_11305,N_9331);
or U12057 (N_12057,N_10421,N_10304);
or U12058 (N_12058,N_11636,N_10501);
or U12059 (N_12059,N_11387,N_10188);
nor U12060 (N_12060,N_10707,N_11027);
nand U12061 (N_12061,N_10141,N_9091);
or U12062 (N_12062,N_10262,N_11736);
nor U12063 (N_12063,N_10897,N_10665);
nor U12064 (N_12064,N_11745,N_9397);
nor U12065 (N_12065,N_9551,N_10766);
or U12066 (N_12066,N_11977,N_11392);
and U12067 (N_12067,N_10483,N_10034);
xor U12068 (N_12068,N_9907,N_11638);
nand U12069 (N_12069,N_11672,N_11201);
or U12070 (N_12070,N_9320,N_9527);
nor U12071 (N_12071,N_9487,N_11449);
nand U12072 (N_12072,N_10481,N_9221);
nor U12073 (N_12073,N_10186,N_10995);
nor U12074 (N_12074,N_9582,N_11132);
and U12075 (N_12075,N_10982,N_11821);
and U12076 (N_12076,N_9446,N_11685);
and U12077 (N_12077,N_9447,N_9694);
nand U12078 (N_12078,N_11913,N_11023);
nor U12079 (N_12079,N_10562,N_9304);
or U12080 (N_12080,N_11364,N_11417);
or U12081 (N_12081,N_10558,N_10643);
or U12082 (N_12082,N_11556,N_10456);
and U12083 (N_12083,N_11633,N_10703);
nand U12084 (N_12084,N_11807,N_11353);
and U12085 (N_12085,N_9746,N_11492);
nand U12086 (N_12086,N_11532,N_9709);
or U12087 (N_12087,N_11781,N_10265);
nor U12088 (N_12088,N_9948,N_11907);
nand U12089 (N_12089,N_11138,N_9965);
nand U12090 (N_12090,N_10374,N_10035);
nor U12091 (N_12091,N_10316,N_11969);
and U12092 (N_12092,N_10639,N_10742);
nor U12093 (N_12093,N_11994,N_11620);
nand U12094 (N_12094,N_10286,N_10940);
nor U12095 (N_12095,N_11281,N_11167);
and U12096 (N_12096,N_11530,N_9863);
nand U12097 (N_12097,N_9059,N_9457);
nor U12098 (N_12098,N_10725,N_10081);
nor U12099 (N_12099,N_11508,N_10041);
nor U12100 (N_12100,N_11463,N_10086);
or U12101 (N_12101,N_10302,N_9816);
nand U12102 (N_12102,N_9847,N_10774);
and U12103 (N_12103,N_11577,N_10069);
xor U12104 (N_12104,N_10129,N_10278);
or U12105 (N_12105,N_11119,N_11618);
or U12106 (N_12106,N_9281,N_11561);
nor U12107 (N_12107,N_9147,N_11077);
nor U12108 (N_12108,N_9957,N_10517);
nor U12109 (N_12109,N_9300,N_11627);
nand U12110 (N_12110,N_9249,N_11924);
nand U12111 (N_12111,N_9776,N_11342);
or U12112 (N_12112,N_10846,N_11501);
and U12113 (N_12113,N_10037,N_9149);
and U12114 (N_12114,N_9063,N_9443);
nor U12115 (N_12115,N_11088,N_9505);
nor U12116 (N_12116,N_10529,N_11036);
and U12117 (N_12117,N_10719,N_11135);
nand U12118 (N_12118,N_9414,N_11017);
nor U12119 (N_12119,N_9857,N_11432);
or U12120 (N_12120,N_9563,N_10807);
nor U12121 (N_12121,N_10965,N_10053);
nand U12122 (N_12122,N_11563,N_11471);
nor U12123 (N_12123,N_11287,N_10343);
and U12124 (N_12124,N_11918,N_10108);
and U12125 (N_12125,N_9566,N_11813);
nor U12126 (N_12126,N_11710,N_9502);
or U12127 (N_12127,N_11767,N_10770);
nor U12128 (N_12128,N_10794,N_10854);
and U12129 (N_12129,N_11900,N_10782);
or U12130 (N_12130,N_10899,N_9222);
nand U12131 (N_12131,N_10157,N_9970);
or U12132 (N_12132,N_11445,N_10922);
and U12133 (N_12133,N_9705,N_9061);
and U12134 (N_12134,N_11586,N_10303);
nor U12135 (N_12135,N_10942,N_11106);
nor U12136 (N_12136,N_11843,N_9291);
or U12137 (N_12137,N_11565,N_11022);
and U12138 (N_12138,N_9617,N_10195);
nand U12139 (N_12139,N_9516,N_11122);
and U12140 (N_12140,N_9879,N_10627);
nand U12141 (N_12141,N_9593,N_11762);
and U12142 (N_12142,N_9892,N_10171);
or U12143 (N_12143,N_11705,N_9372);
nand U12144 (N_12144,N_11011,N_10049);
nand U12145 (N_12145,N_9804,N_9402);
or U12146 (N_12146,N_9318,N_10152);
nand U12147 (N_12147,N_10551,N_11457);
nor U12148 (N_12148,N_10866,N_11065);
and U12149 (N_12149,N_9600,N_11856);
and U12150 (N_12150,N_10324,N_10826);
or U12151 (N_12151,N_9116,N_11297);
and U12152 (N_12152,N_11384,N_11742);
nand U12153 (N_12153,N_11372,N_11630);
or U12154 (N_12154,N_10469,N_9205);
nor U12155 (N_12155,N_11646,N_9018);
nand U12156 (N_12156,N_11689,N_9913);
nor U12157 (N_12157,N_10104,N_9854);
or U12158 (N_12158,N_9655,N_9634);
and U12159 (N_12159,N_11734,N_11634);
or U12160 (N_12160,N_11242,N_11075);
or U12161 (N_12161,N_9615,N_11976);
nand U12162 (N_12162,N_9980,N_10347);
nor U12163 (N_12163,N_11336,N_9189);
nor U12164 (N_12164,N_11920,N_11335);
or U12165 (N_12165,N_10706,N_11162);
and U12166 (N_12166,N_11279,N_9111);
nor U12167 (N_12167,N_10080,N_10518);
and U12168 (N_12168,N_10934,N_10282);
or U12169 (N_12169,N_11737,N_10388);
and U12170 (N_12170,N_11664,N_11564);
nand U12171 (N_12171,N_11776,N_11025);
or U12172 (N_12172,N_11044,N_9420);
and U12173 (N_12173,N_9821,N_11395);
nor U12174 (N_12174,N_9417,N_10477);
nand U12175 (N_12175,N_10118,N_9576);
nor U12176 (N_12176,N_11483,N_9667);
or U12177 (N_12177,N_10221,N_9981);
nand U12178 (N_12178,N_11985,N_10582);
nand U12179 (N_12179,N_10193,N_9412);
nand U12180 (N_12180,N_11637,N_9031);
nand U12181 (N_12181,N_9444,N_9491);
and U12182 (N_12182,N_11677,N_11730);
nand U12183 (N_12183,N_10084,N_11422);
nor U12184 (N_12184,N_10635,N_9522);
or U12185 (N_12185,N_9390,N_9805);
nor U12186 (N_12186,N_10196,N_11408);
nand U12187 (N_12187,N_10888,N_10771);
or U12188 (N_12188,N_10073,N_11264);
nand U12189 (N_12189,N_11667,N_10482);
or U12190 (N_12190,N_11639,N_9951);
nand U12191 (N_12191,N_11394,N_9668);
or U12192 (N_12192,N_9202,N_10829);
nor U12193 (N_12193,N_9324,N_10592);
or U12194 (N_12194,N_11173,N_9993);
or U12195 (N_12195,N_9405,N_10154);
nor U12196 (N_12196,N_10756,N_10179);
or U12197 (N_12197,N_9197,N_9440);
or U12198 (N_12198,N_9148,N_11622);
or U12199 (N_12199,N_10266,N_11296);
and U12200 (N_12200,N_10396,N_10307);
or U12201 (N_12201,N_9922,N_10968);
and U12202 (N_12202,N_10137,N_9125);
and U12203 (N_12203,N_11702,N_11783);
xnor U12204 (N_12204,N_11413,N_9734);
or U12205 (N_12205,N_10754,N_11943);
nand U12206 (N_12206,N_10395,N_10608);
or U12207 (N_12207,N_11754,N_10452);
and U12208 (N_12208,N_11020,N_10046);
nor U12209 (N_12209,N_11465,N_9374);
nand U12210 (N_12210,N_9688,N_9445);
or U12211 (N_12211,N_9478,N_9313);
nand U12212 (N_12212,N_9573,N_9706);
or U12213 (N_12213,N_11176,N_11551);
or U12214 (N_12214,N_11200,N_9039);
and U12215 (N_12215,N_9302,N_11916);
or U12216 (N_12216,N_11219,N_9939);
nand U12217 (N_12217,N_10723,N_10811);
nor U12218 (N_12218,N_9439,N_11590);
or U12219 (N_12219,N_10117,N_11248);
nor U12220 (N_12220,N_9200,N_11321);
nor U12221 (N_12221,N_11359,N_10532);
and U12222 (N_12222,N_10543,N_9619);
nand U12223 (N_12223,N_11751,N_10406);
nor U12224 (N_12224,N_9650,N_10561);
nand U12225 (N_12225,N_9652,N_9643);
and U12226 (N_12226,N_10270,N_10735);
nor U12227 (N_12227,N_11116,N_11363);
and U12228 (N_12228,N_9739,N_11621);
and U12229 (N_12229,N_11750,N_11085);
and U12230 (N_12230,N_9921,N_9424);
and U12231 (N_12231,N_10649,N_9784);
and U12232 (N_12232,N_11837,N_11653);
nand U12233 (N_12233,N_10954,N_11740);
nand U12234 (N_12234,N_11720,N_10533);
nand U12235 (N_12235,N_9775,N_11066);
nand U12236 (N_12236,N_10353,N_9261);
or U12237 (N_12237,N_10061,N_10333);
and U12238 (N_12238,N_10748,N_9081);
and U12239 (N_12239,N_10684,N_10675);
nand U12240 (N_12240,N_11955,N_9565);
or U12241 (N_12241,N_10528,N_9299);
or U12242 (N_12242,N_9729,N_9486);
nand U12243 (N_12243,N_9112,N_10566);
nor U12244 (N_12244,N_9097,N_10641);
nand U12245 (N_12245,N_11727,N_11427);
nor U12246 (N_12246,N_10202,N_9428);
nand U12247 (N_12247,N_9518,N_9160);
nor U12248 (N_12248,N_11999,N_10047);
and U12249 (N_12249,N_10309,N_9323);
nor U12250 (N_12250,N_10223,N_10652);
or U12251 (N_12251,N_10726,N_10973);
and U12252 (N_12252,N_9224,N_11486);
nor U12253 (N_12253,N_9823,N_11129);
nand U12254 (N_12254,N_10586,N_10085);
and U12255 (N_12255,N_10985,N_9388);
and U12256 (N_12256,N_11842,N_10509);
and U12257 (N_12257,N_9226,N_10859);
and U12258 (N_12258,N_9779,N_11991);
or U12259 (N_12259,N_11487,N_11145);
nor U12260 (N_12260,N_10245,N_10392);
nand U12261 (N_12261,N_9984,N_11052);
nor U12262 (N_12262,N_9864,N_10553);
and U12263 (N_12263,N_11056,N_9525);
nor U12264 (N_12264,N_11000,N_10383);
or U12265 (N_12265,N_10852,N_9436);
nand U12266 (N_12266,N_9630,N_10148);
nand U12267 (N_12267,N_11546,N_10230);
nand U12268 (N_12268,N_10342,N_10306);
and U12269 (N_12269,N_10050,N_11930);
or U12270 (N_12270,N_11139,N_10775);
or U12271 (N_12271,N_11081,N_11261);
and U12272 (N_12272,N_10401,N_10783);
and U12273 (N_12273,N_9698,N_9968);
nor U12274 (N_12274,N_10746,N_11704);
nor U12275 (N_12275,N_9943,N_9215);
or U12276 (N_12276,N_9768,N_10984);
and U12277 (N_12277,N_10929,N_9560);
or U12278 (N_12278,N_9684,N_9819);
and U12279 (N_12279,N_11191,N_9931);
or U12280 (N_12280,N_9099,N_10651);
nor U12281 (N_12281,N_10698,N_10970);
or U12282 (N_12282,N_9852,N_11280);
and U12283 (N_12283,N_9273,N_10580);
nor U12284 (N_12284,N_10348,N_9271);
nor U12285 (N_12285,N_10346,N_11941);
nor U12286 (N_12286,N_11935,N_11759);
or U12287 (N_12287,N_10902,N_10900);
or U12288 (N_12288,N_9946,N_11974);
or U12289 (N_12289,N_10339,N_10840);
and U12290 (N_12290,N_9631,N_10587);
and U12291 (N_12291,N_10439,N_9407);
nor U12292 (N_12292,N_9531,N_10631);
nand U12293 (N_12293,N_10883,N_11123);
nand U12294 (N_12294,N_10419,N_9987);
or U12295 (N_12295,N_10550,N_9870);
nand U12296 (N_12296,N_10564,N_11390);
or U12297 (N_12297,N_10412,N_10619);
and U12298 (N_12298,N_9151,N_11500);
nand U12299 (N_12299,N_9911,N_10087);
nor U12300 (N_12300,N_11361,N_10674);
or U12301 (N_12301,N_9541,N_11034);
nand U12302 (N_12302,N_9868,N_10459);
nand U12303 (N_12303,N_11520,N_9935);
nor U12304 (N_12304,N_11589,N_10806);
and U12305 (N_12305,N_11499,N_9076);
nand U12306 (N_12306,N_10938,N_10424);
and U12307 (N_12307,N_11478,N_10535);
or U12308 (N_12308,N_9367,N_9512);
nand U12309 (N_12309,N_11403,N_11093);
or U12310 (N_12310,N_10426,N_9985);
nand U12311 (N_12311,N_11801,N_11005);
nor U12312 (N_12312,N_9697,N_9395);
or U12313 (N_12313,N_10417,N_9442);
or U12314 (N_12314,N_10858,N_9422);
and U12315 (N_12315,N_9726,N_9660);
nor U12316 (N_12316,N_9358,N_9232);
nand U12317 (N_12317,N_9592,N_11882);
nand U12318 (N_12318,N_11569,N_11354);
or U12319 (N_12319,N_11018,N_10497);
nor U12320 (N_12320,N_11657,N_11035);
and U12321 (N_12321,N_10058,N_10364);
or U12322 (N_12322,N_10602,N_9381);
nand U12323 (N_12323,N_9473,N_10089);
nor U12324 (N_12324,N_10875,N_10299);
nand U12325 (N_12325,N_10464,N_10743);
nand U12326 (N_12326,N_9789,N_10345);
and U12327 (N_12327,N_9553,N_9554);
nand U12328 (N_12328,N_9168,N_10096);
nand U12329 (N_12329,N_9877,N_10176);
nor U12330 (N_12330,N_9398,N_11833);
and U12331 (N_12331,N_9699,N_11814);
nand U12332 (N_12332,N_11865,N_11687);
or U12333 (N_12333,N_10493,N_9196);
nor U12334 (N_12334,N_9394,N_9046);
nor U12335 (N_12335,N_11143,N_9693);
and U12336 (N_12336,N_11883,N_9211);
and U12337 (N_12337,N_11755,N_9426);
or U12338 (N_12338,N_9558,N_10352);
or U12339 (N_12339,N_9166,N_10335);
nand U12340 (N_12340,N_10006,N_9359);
nand U12341 (N_12341,N_10787,N_11678);
and U12342 (N_12342,N_10716,N_9139);
nor U12343 (N_12343,N_11697,N_11448);
nor U12344 (N_12344,N_10704,N_10921);
nand U12345 (N_12345,N_10959,N_11835);
nand U12346 (N_12346,N_10884,N_11374);
nand U12347 (N_12347,N_10963,N_10721);
and U12348 (N_12348,N_9572,N_9741);
and U12349 (N_12349,N_10045,N_10622);
and U12350 (N_12350,N_10790,N_9027);
or U12351 (N_12351,N_11185,N_9484);
nand U12352 (N_12352,N_9192,N_11344);
nor U12353 (N_12353,N_9343,N_11871);
xor U12354 (N_12354,N_9774,N_11451);
nand U12355 (N_12355,N_11049,N_9389);
nor U12356 (N_12356,N_9887,N_9703);
nand U12357 (N_12357,N_10511,N_11700);
nor U12358 (N_12358,N_11831,N_9665);
nor U12359 (N_12359,N_9078,N_11908);
and U12360 (N_12360,N_10372,N_11905);
or U12361 (N_12361,N_10733,N_9795);
or U12362 (N_12362,N_9647,N_11369);
nor U12363 (N_12363,N_11679,N_10163);
nand U12364 (N_12364,N_10492,N_11961);
and U12365 (N_12365,N_11719,N_10393);
or U12366 (N_12366,N_9810,N_10005);
nor U12367 (N_12367,N_9322,N_11131);
nand U12368 (N_12368,N_11885,N_9843);
nand U12369 (N_12369,N_11378,N_11975);
or U12370 (N_12370,N_9024,N_11199);
nand U12371 (N_12371,N_11029,N_10066);
and U12372 (N_12372,N_10632,N_11168);
and U12373 (N_12373,N_11788,N_11558);
nor U12374 (N_12374,N_11197,N_10927);
or U12375 (N_12375,N_11959,N_11543);
or U12376 (N_12376,N_9602,N_9798);
or U12377 (N_12377,N_10634,N_9051);
nand U12378 (N_12378,N_11238,N_9754);
nor U12379 (N_12379,N_10368,N_11611);
and U12380 (N_12380,N_9788,N_11873);
and U12381 (N_12381,N_9140,N_10106);
and U12382 (N_12382,N_11136,N_10548);
and U12383 (N_12383,N_11707,N_9785);
and U12384 (N_12384,N_9825,N_11090);
or U12385 (N_12385,N_9986,N_9861);
and U12386 (N_12386,N_9000,N_10074);
nor U12387 (N_12387,N_10397,N_9158);
and U12388 (N_12388,N_11466,N_11229);
nand U12389 (N_12389,N_9777,N_9945);
nor U12390 (N_12390,N_10809,N_11834);
nand U12391 (N_12391,N_9504,N_10885);
or U12392 (N_12392,N_9562,N_9396);
and U12393 (N_12393,N_11698,N_9839);
nor U12394 (N_12394,N_9293,N_10654);
or U12395 (N_12395,N_9674,N_9828);
nand U12396 (N_12396,N_9385,N_9966);
and U12397 (N_12397,N_11869,N_10758);
or U12398 (N_12398,N_9365,N_11244);
nand U12399 (N_12399,N_11157,N_10391);
or U12400 (N_12400,N_11895,N_11911);
or U12401 (N_12401,N_11937,N_9142);
or U12402 (N_12402,N_9599,N_11993);
nand U12403 (N_12403,N_10088,N_9737);
or U12404 (N_12404,N_9283,N_10190);
nand U12405 (N_12405,N_11899,N_9418);
nand U12406 (N_12406,N_10461,N_9506);
or U12407 (N_12407,N_9707,N_9579);
and U12408 (N_12408,N_9383,N_9071);
and U12409 (N_12409,N_11626,N_11925);
or U12410 (N_12410,N_9203,N_11944);
nand U12411 (N_12411,N_9416,N_11805);
or U12412 (N_12412,N_9964,N_9217);
and U12413 (N_12413,N_9791,N_10994);
nor U12414 (N_12414,N_11385,N_11064);
or U12415 (N_12415,N_11681,N_10070);
or U12416 (N_12416,N_10191,N_11701);
nor U12417 (N_12417,N_10662,N_10798);
nor U12418 (N_12418,N_10004,N_10312);
and U12419 (N_12419,N_10795,N_9766);
nor U12420 (N_12420,N_11610,N_11105);
or U12421 (N_12421,N_10199,N_11291);
and U12422 (N_12422,N_11998,N_9057);
and U12423 (N_12423,N_9613,N_11819);
or U12424 (N_12424,N_11855,N_11827);
or U12425 (N_12425,N_11560,N_9616);
nor U12426 (N_12426,N_9186,N_11523);
nor U12427 (N_12427,N_10325,N_10712);
and U12428 (N_12428,N_11596,N_11473);
nand U12429 (N_12429,N_11256,N_10438);
nand U12430 (N_12430,N_11995,N_11850);
nand U12431 (N_12431,N_11437,N_10336);
nor U12432 (N_12432,N_11922,N_10863);
and U12433 (N_12433,N_9356,N_9812);
nand U12434 (N_12434,N_10246,N_10673);
nand U12435 (N_12435,N_9678,N_9845);
nor U12436 (N_12436,N_10642,N_11957);
and U12437 (N_12437,N_10822,N_10495);
or U12438 (N_12438,N_11832,N_11927);
and U12439 (N_12439,N_9888,N_9364);
or U12440 (N_12440,N_9666,N_11992);
and U12441 (N_12441,N_11534,N_10120);
and U12442 (N_12442,N_11808,N_11194);
or U12443 (N_12443,N_11779,N_9903);
and U12444 (N_12444,N_10600,N_11772);
and U12445 (N_12445,N_11493,N_9858);
or U12446 (N_12446,N_10728,N_9201);
nor U12447 (N_12447,N_9242,N_10488);
nor U12448 (N_12448,N_11470,N_10572);
nand U12449 (N_12449,N_10057,N_11480);
nor U12450 (N_12450,N_10741,N_9464);
nor U12451 (N_12451,N_11728,N_9761);
or U12452 (N_12452,N_10877,N_10554);
or U12453 (N_12453,N_10827,N_11529);
and U12454 (N_12454,N_10930,N_9471);
nand U12455 (N_12455,N_11195,N_9480);
and U12456 (N_12456,N_11447,N_11016);
nor U12457 (N_12457,N_10121,N_10454);
nor U12458 (N_12458,N_11325,N_10192);
and U12459 (N_12459,N_11076,N_11858);
or U12460 (N_12460,N_11915,N_10321);
or U12461 (N_12461,N_11602,N_11268);
nor U12462 (N_12462,N_9080,N_11355);
and U12463 (N_12463,N_10623,N_9883);
and U12464 (N_12464,N_11892,N_10433);
nand U12465 (N_12465,N_9441,N_10480);
nor U12466 (N_12466,N_11345,N_10209);
and U12467 (N_12467,N_9559,N_9288);
nor U12468 (N_12468,N_10563,N_10217);
nor U12469 (N_12469,N_11756,N_9329);
or U12470 (N_12470,N_11582,N_11316);
and U12471 (N_12471,N_9757,N_9497);
nor U12472 (N_12472,N_11625,N_9386);
nand U12473 (N_12473,N_11134,N_11362);
and U12474 (N_12474,N_9783,N_9360);
or U12475 (N_12475,N_9833,N_11786);
and U12476 (N_12476,N_11950,N_11285);
and U12477 (N_12477,N_10479,N_11425);
nor U12478 (N_12478,N_9079,N_11598);
nor U12479 (N_12479,N_9749,N_10538);
nand U12480 (N_12480,N_10128,N_11929);
and U12481 (N_12481,N_9008,N_9207);
nand U12482 (N_12482,N_10686,N_11294);
and U12483 (N_12483,N_11398,N_10935);
nand U12484 (N_12484,N_9521,N_10633);
nand U12485 (N_12485,N_9640,N_9580);
nor U12486 (N_12486,N_11358,N_10910);
nand U12487 (N_12487,N_11531,N_10720);
and U12488 (N_12488,N_9824,N_10378);
nand U12489 (N_12489,N_9252,N_10996);
nand U12490 (N_12490,N_11045,N_10140);
nand U12491 (N_12491,N_11746,N_11507);
and U12492 (N_12492,N_10376,N_9260);
nand U12493 (N_12493,N_10909,N_9278);
nor U12494 (N_12494,N_11028,N_10976);
and U12495 (N_12495,N_11796,N_10546);
or U12496 (N_12496,N_10932,N_11102);
or U12497 (N_12497,N_9419,N_9346);
and U12498 (N_12498,N_9756,N_9875);
or U12499 (N_12499,N_11635,N_11806);
nand U12500 (N_12500,N_9157,N_10616);
nand U12501 (N_12501,N_11450,N_9725);
or U12502 (N_12502,N_9614,N_9673);
and U12503 (N_12503,N_10201,N_11690);
or U12504 (N_12504,N_10646,N_9287);
nor U12505 (N_12505,N_10441,N_10919);
nand U12506 (N_12506,N_11711,N_10229);
nor U12507 (N_12507,N_11379,N_10625);
or U12508 (N_12508,N_11232,N_10340);
or U12509 (N_12509,N_11249,N_10276);
and U12510 (N_12510,N_10845,N_9781);
nand U12511 (N_12511,N_9626,N_9924);
nand U12512 (N_12512,N_11643,N_11062);
and U12513 (N_12513,N_11193,N_11645);
nor U12514 (N_12514,N_9241,N_9228);
and U12515 (N_12515,N_11443,N_10802);
and U12516 (N_12516,N_11152,N_10914);
nor U12517 (N_12517,N_9223,N_10975);
and U12518 (N_12518,N_10314,N_10269);
nand U12519 (N_12519,N_9545,N_11380);
or U12520 (N_12520,N_10960,N_10585);
nand U12521 (N_12521,N_10000,N_11576);
and U12522 (N_12522,N_10135,N_10411);
nand U12523 (N_12523,N_10853,N_10234);
or U12524 (N_12524,N_9431,N_11524);
nor U12525 (N_12525,N_9896,N_9762);
nand U12526 (N_12526,N_11713,N_10872);
nand U12527 (N_12527,N_9255,N_11938);
nor U12528 (N_12528,N_9639,N_9889);
nor U12529 (N_12529,N_9182,N_11241);
and U12530 (N_12530,N_10273,N_11880);
nand U12531 (N_12531,N_11562,N_11488);
and U12532 (N_12532,N_10887,N_11087);
or U12533 (N_12533,N_10218,N_11477);
and U12534 (N_12534,N_9826,N_11775);
or U12535 (N_12535,N_10659,N_11726);
nor U12536 (N_12536,N_10896,N_10164);
and U12537 (N_12537,N_11259,N_9696);
nand U12538 (N_12538,N_10801,N_11187);
nor U12539 (N_12539,N_11037,N_10628);
and U12540 (N_12540,N_9335,N_11795);
or U12541 (N_12541,N_10011,N_9989);
nor U12542 (N_12542,N_11793,N_11648);
nand U12543 (N_12543,N_9369,N_11980);
and U12544 (N_12544,N_9654,N_10653);
or U12545 (N_12545,N_11420,N_11410);
nor U12546 (N_12546,N_11226,N_9129);
or U12547 (N_12547,N_9865,N_9662);
nor U12548 (N_12548,N_9060,N_9423);
or U12549 (N_12549,N_11245,N_11300);
or U12550 (N_12550,N_11641,N_9107);
and U12551 (N_12551,N_11897,N_9792);
nand U12552 (N_12552,N_9786,N_9371);
and U12553 (N_12553,N_11503,N_9927);
nand U12554 (N_12554,N_9169,N_9495);
and U12555 (N_12555,N_11770,N_11051);
xor U12556 (N_12556,N_10620,N_11227);
nor U12557 (N_12557,N_11346,N_9680);
nand U12558 (N_12558,N_11108,N_10261);
and U12559 (N_12559,N_9354,N_10116);
and U12560 (N_12560,N_10028,N_9137);
or U12561 (N_12561,N_9043,N_11587);
nor U12562 (N_12562,N_11881,N_10796);
and U12563 (N_12563,N_11026,N_10060);
and U12564 (N_12564,N_9178,N_10889);
nor U12565 (N_12565,N_9032,N_10008);
nand U12566 (N_12566,N_11223,N_9701);
nor U12567 (N_12567,N_9738,N_11706);
nor U12568 (N_12568,N_11349,N_11290);
or U12569 (N_12569,N_11515,N_11252);
nor U12570 (N_12570,N_10904,N_9982);
nand U12571 (N_12571,N_11603,N_9998);
and U12572 (N_12572,N_10769,N_10055);
nand U12573 (N_12573,N_9585,N_9303);
and U12574 (N_12574,N_10486,N_11903);
and U12575 (N_12575,N_11774,N_10664);
nor U12576 (N_12576,N_9351,N_11549);
xor U12577 (N_12577,N_9977,N_9919);
nor U12578 (N_12578,N_10506,N_11299);
and U12579 (N_12579,N_9733,N_10054);
nor U12580 (N_12580,N_11069,N_9154);
or U12581 (N_12581,N_11860,N_10002);
nor U12582 (N_12582,N_10332,N_10494);
nor U12583 (N_12583,N_10228,N_9244);
nand U12584 (N_12584,N_11965,N_10986);
nand U12585 (N_12585,N_11120,N_9049);
nor U12586 (N_12586,N_10966,N_9878);
nor U12587 (N_12587,N_11475,N_9295);
nand U12588 (N_12588,N_9044,N_11867);
or U12589 (N_12589,N_9641,N_11725);
and U12590 (N_12590,N_9347,N_11777);
and U12591 (N_12591,N_10891,N_10090);
nand U12592 (N_12592,N_10779,N_11172);
nand U12593 (N_12593,N_11295,N_11878);
nand U12594 (N_12594,N_9003,N_10151);
or U12595 (N_12595,N_10834,N_11815);
nand U12596 (N_12596,N_10717,N_9535);
or U12597 (N_12597,N_10422,N_10009);
nand U12598 (N_12598,N_11092,N_11401);
and U12599 (N_12599,N_11262,N_11192);
or U12600 (N_12600,N_10830,N_11014);
and U12601 (N_12601,N_9298,N_9571);
or U12602 (N_12602,N_10231,N_11919);
and U12603 (N_12603,N_9934,N_10258);
and U12604 (N_12604,N_11166,N_11512);
nand U12605 (N_12605,N_9568,N_9163);
and U12606 (N_12606,N_10350,N_11953);
nor U12607 (N_12607,N_11811,N_11840);
or U12608 (N_12608,N_11658,N_11968);
or U12609 (N_12609,N_11298,N_11591);
nand U12610 (N_12610,N_10267,N_11495);
or U12611 (N_12611,N_10415,N_10715);
and U12612 (N_12612,N_9642,N_11411);
nand U12613 (N_12613,N_10026,N_10124);
nand U12614 (N_12614,N_11141,N_10638);
or U12615 (N_12615,N_9475,N_11033);
and U12616 (N_12616,N_11375,N_9933);
nor U12617 (N_12617,N_9465,N_9276);
nor U12618 (N_12618,N_10222,N_9013);
or U12619 (N_12619,N_11002,N_9704);
or U12620 (N_12620,N_9509,N_10204);
nand U12621 (N_12621,N_10530,N_11054);
nor U12622 (N_12622,N_10432,N_10578);
and U12623 (N_12623,N_9671,N_9117);
and U12624 (N_12624,N_9605,N_10611);
and U12625 (N_12625,N_11951,N_11253);
or U12626 (N_12626,N_11659,N_10989);
and U12627 (N_12627,N_9025,N_10109);
nand U12628 (N_12628,N_10337,N_9866);
nand U12629 (N_12629,N_9460,N_10077);
nand U12630 (N_12630,N_10420,N_9002);
or U12631 (N_12631,N_11491,N_10161);
nand U12632 (N_12632,N_10599,N_11570);
nand U12633 (N_12633,N_11693,N_9476);
nor U12634 (N_12634,N_11496,N_10819);
nand U12635 (N_12635,N_10418,N_9790);
or U12636 (N_12636,N_11370,N_10851);
nor U12637 (N_12637,N_9123,N_10521);
nand U12638 (N_12638,N_9748,N_10820);
or U12639 (N_12639,N_10663,N_9020);
and U12640 (N_12640,N_11371,N_9014);
and U12641 (N_12641,N_11872,N_10123);
and U12642 (N_12642,N_9477,N_9456);
nor U12643 (N_12643,N_9362,N_10937);
and U12644 (N_12644,N_11594,N_10355);
and U12645 (N_12645,N_9803,N_11382);
or U12646 (N_12646,N_9627,N_10012);
nand U12647 (N_12647,N_9899,N_10040);
and U12648 (N_12648,N_9102,N_10203);
nand U12649 (N_12649,N_11928,N_9095);
nand U12650 (N_12650,N_11548,N_9556);
nand U12651 (N_12651,N_10113,N_9454);
nor U12652 (N_12652,N_10573,N_11671);
or U12653 (N_12653,N_11651,N_11984);
nand U12654 (N_12654,N_11274,N_10042);
and U12655 (N_12655,N_10472,N_9234);
nand U12656 (N_12656,N_11079,N_9840);
nand U12657 (N_12657,N_11997,N_9004);
nand U12658 (N_12658,N_11130,N_9960);
nand U12659 (N_12659,N_11309,N_11113);
nand U12660 (N_12660,N_9213,N_9088);
nor U12661 (N_12661,N_9162,N_10579);
or U12662 (N_12662,N_9867,N_11539);
or U12663 (N_12663,N_11053,N_11171);
or U12664 (N_12664,N_10526,N_9622);
and U12665 (N_12665,N_10291,N_10251);
nor U12666 (N_12666,N_9153,N_9595);
nor U12667 (N_12667,N_11647,N_11251);
nand U12668 (N_12668,N_11761,N_10864);
or U12669 (N_12669,N_10658,N_11469);
nor U12670 (N_12670,N_10075,N_11196);
and U12671 (N_12671,N_11159,N_11163);
nor U12672 (N_12672,N_10833,N_11306);
nand U12673 (N_12673,N_11861,N_10365);
or U12674 (N_12674,N_10825,N_11024);
nand U12675 (N_12675,N_10577,N_10560);
or U12676 (N_12676,N_9056,N_9246);
or U12677 (N_12677,N_10895,N_9474);
nand U12678 (N_12678,N_10294,N_11235);
nor U12679 (N_12679,N_9941,N_11712);
xnor U12680 (N_12680,N_9929,N_11100);
and U12681 (N_12681,N_11839,N_11246);
or U12682 (N_12682,N_11160,N_10784);
nor U12683 (N_12683,N_9104,N_9458);
nand U12684 (N_12684,N_11981,N_11217);
nand U12685 (N_12685,N_9567,N_9316);
nand U12686 (N_12686,N_11179,N_11099);
or U12687 (N_12687,N_9068,N_10358);
nand U12688 (N_12688,N_9969,N_9555);
nor U12689 (N_12689,N_11642,N_10951);
nand U12690 (N_12690,N_11341,N_9523);
nand U12691 (N_12691,N_10861,N_10657);
and U12692 (N_12692,N_11960,N_9597);
nor U12693 (N_12693,N_10216,N_10855);
and U12694 (N_12694,N_11818,N_11164);
nor U12695 (N_12695,N_10869,N_9047);
nand U12696 (N_12696,N_11624,N_11886);
or U12697 (N_12697,N_9620,N_9481);
or U12698 (N_12698,N_9237,N_10277);
nand U12699 (N_12699,N_10512,N_9740);
nand U12700 (N_12700,N_9070,N_9758);
nor U12701 (N_12701,N_10435,N_11841);
nor U12702 (N_12702,N_10797,N_11810);
and U12703 (N_12703,N_10757,N_11061);
and U12704 (N_12704,N_9220,N_10936);
nor U12705 (N_12705,N_11744,N_9494);
and U12706 (N_12706,N_10752,N_11074);
nand U12707 (N_12707,N_11111,N_10115);
nor U12708 (N_12708,N_9838,N_9349);
or U12709 (N_12709,N_9256,N_10048);
and U12710 (N_12710,N_11434,N_9400);
nand U12711 (N_12711,N_11741,N_9711);
nor U12712 (N_12712,N_9198,N_11180);
nor U12713 (N_12713,N_10067,N_11096);
nand U12714 (N_12714,N_11351,N_11812);
xnor U12715 (N_12715,N_11303,N_11334);
or U12716 (N_12716,N_10540,N_9308);
nand U12717 (N_12717,N_11041,N_10250);
nor U12718 (N_12718,N_11320,N_11497);
nor U12719 (N_12719,N_10524,N_9664);
or U12720 (N_12720,N_10575,N_11008);
nor U12721 (N_12721,N_10403,N_9006);
and U12722 (N_12722,N_11484,N_10740);
and U12723 (N_12723,N_10102,N_9656);
nor U12724 (N_12724,N_11825,N_10789);
nor U12725 (N_12725,N_10175,N_10205);
and U12726 (N_12726,N_11824,N_11304);
xnor U12727 (N_12727,N_9856,N_9488);
nand U12728 (N_12728,N_11494,N_9219);
and U12729 (N_12729,N_10371,N_11763);
nor U12730 (N_12730,N_10330,N_10626);
nor U12731 (N_12731,N_10100,N_10173);
nor U12732 (N_12732,N_10737,N_10878);
and U12733 (N_12733,N_10295,N_10727);
and U12734 (N_12734,N_9282,N_11010);
or U12735 (N_12735,N_9230,N_11012);
and U12736 (N_12736,N_10677,N_11050);
nor U12737 (N_12737,N_11675,N_10134);
nor U12738 (N_12738,N_9963,N_11605);
or U12739 (N_12739,N_10823,N_11912);
nor U12740 (N_12740,N_10142,N_11038);
nor U12741 (N_12741,N_9310,N_10781);
and U12742 (N_12742,N_10541,N_11456);
or U12743 (N_12743,N_10021,N_11430);
nand U12744 (N_12744,N_9434,N_11352);
nand U12745 (N_12745,N_10792,N_9608);
nor U12746 (N_12746,N_11902,N_11789);
and U12747 (N_12747,N_9542,N_9370);
or U12748 (N_12748,N_11233,N_9411);
or U12749 (N_12749,N_9764,N_9884);
nor U12750 (N_12750,N_10948,N_11691);
xor U12751 (N_12751,N_9583,N_10198);
nor U12752 (N_12752,N_9301,N_9325);
or U12753 (N_12753,N_10977,N_10394);
and U12754 (N_12754,N_9247,N_10760);
or U12755 (N_12755,N_11822,N_9493);
nor U12756 (N_12756,N_9152,N_10308);
nand U12757 (N_12757,N_9482,N_10923);
and U12758 (N_12758,N_10373,N_9820);
or U12759 (N_12759,N_10590,N_10023);
nand U12760 (N_12760,N_11007,N_9953);
nand U12761 (N_12761,N_10763,N_11936);
and U12762 (N_12762,N_11505,N_9735);
nor U12763 (N_12763,N_9610,N_11239);
and U12764 (N_12764,N_9468,N_9409);
nand U12765 (N_12765,N_9384,N_9227);
nor U12766 (N_12766,N_9971,N_10928);
nor U12767 (N_12767,N_9687,N_10409);
and U12768 (N_12768,N_11339,N_9589);
nor U12769 (N_12769,N_10044,N_10200);
and U12770 (N_12770,N_11293,N_10793);
and U12771 (N_12771,N_9285,N_9517);
nor U12772 (N_12772,N_10924,N_9485);
and U12773 (N_12773,N_10458,N_10804);
or U12774 (N_12774,N_9188,N_10437);
nand U12775 (N_12775,N_9780,N_9120);
nand U12776 (N_12776,N_9114,N_10099);
or U12777 (N_12777,N_10010,N_9159);
nand U12778 (N_12778,N_10886,N_10860);
or U12779 (N_12779,N_10762,N_9808);
or U12780 (N_12780,N_9724,N_10785);
or U12781 (N_12781,N_10232,N_9108);
nand U12782 (N_12782,N_10465,N_11519);
and U12783 (N_12783,N_9728,N_11149);
nor U12784 (N_12784,N_10534,N_10591);
and U12785 (N_12785,N_10275,N_11844);
or U12786 (N_12786,N_11003,N_10767);
and U12787 (N_12787,N_10359,N_9806);
nor U12788 (N_12788,N_10356,N_9011);
nand U12789 (N_12789,N_10156,N_10531);
and U12790 (N_12790,N_10856,N_10547);
nand U12791 (N_12791,N_9685,N_11461);
nor U12792 (N_12792,N_9363,N_10696);
nor U12793 (N_12793,N_11424,N_10516);
nor U12794 (N_12794,N_9624,N_9990);
or U12795 (N_12795,N_10062,N_11753);
nand U12796 (N_12796,N_11875,N_9799);
nor U12797 (N_12797,N_9053,N_11588);
and U12798 (N_12798,N_9837,N_9466);
and U12799 (N_12799,N_11593,N_9250);
or U12800 (N_12800,N_10640,N_11521);
nand U12801 (N_12801,N_9603,N_10843);
nor U12802 (N_12802,N_11567,N_9961);
and U12803 (N_12803,N_9330,N_11031);
or U12804 (N_12804,N_11552,N_9793);
or U12805 (N_12805,N_11663,N_11506);
or U12806 (N_12806,N_9333,N_9700);
nor U12807 (N_12807,N_10969,N_11866);
and U12808 (N_12808,N_11169,N_11383);
nor U12809 (N_12809,N_10943,N_10739);
nor U12810 (N_12810,N_9510,N_11578);
nand U12811 (N_12811,N_10366,N_9399);
or U12812 (N_12812,N_9164,N_10815);
and U12813 (N_12813,N_10849,N_11544);
and U12814 (N_12814,N_10159,N_9874);
or U12815 (N_12815,N_11435,N_10593);
nor U12816 (N_12816,N_11939,N_11743);
nand U12817 (N_12817,N_9978,N_10617);
or U12818 (N_12818,N_11006,N_11406);
nor U12819 (N_12819,N_9538,N_9127);
and U12820 (N_12820,N_9366,N_9378);
nor U12821 (N_12821,N_9916,N_11948);
nor U12822 (N_12822,N_9101,N_11302);
xnor U12823 (N_12823,N_10672,N_11849);
nand U12824 (N_12824,N_10722,N_10603);
and U12825 (N_12825,N_11055,N_9578);
nor U12826 (N_12826,N_11071,N_9809);
nand U12827 (N_12827,N_9753,N_11439);
nor U12828 (N_12828,N_11933,N_11386);
nand U12829 (N_12829,N_9822,N_10298);
and U12830 (N_12830,N_10882,N_11277);
nand U12831 (N_12831,N_10842,N_11686);
nand U12832 (N_12832,N_9064,N_10387);
nand U12833 (N_12833,N_10281,N_9853);
or U12834 (N_12834,N_9144,N_9459);
nor U12835 (N_12835,N_10105,N_10127);
nor U12836 (N_12836,N_9782,N_10428);
and U12837 (N_12837,N_9936,N_10318);
nor U12838 (N_12838,N_9587,N_9606);
and U12839 (N_12839,N_10430,N_9683);
nand U12840 (N_12840,N_9297,N_11739);
or U12841 (N_12841,N_10736,N_9479);
nor U12842 (N_12842,N_10903,N_11688);
nor U12843 (N_12843,N_10685,N_11926);
nor U12844 (N_12844,N_9677,N_10700);
and U12845 (N_12845,N_11270,N_9055);
nor U12846 (N_12846,N_9850,N_10519);
or U12847 (N_12847,N_10300,N_11988);
or U12848 (N_12848,N_9187,N_11893);
nand U12849 (N_12849,N_9126,N_9596);
or U12850 (N_12850,N_10279,N_10369);
nand U12851 (N_12851,N_11932,N_9882);
nand U12852 (N_12852,N_10146,N_11575);
and U12853 (N_12853,N_9185,N_9262);
nand U12854 (N_12854,N_11715,N_10227);
and U12855 (N_12855,N_10466,N_9972);
nor U12856 (N_12856,N_10865,N_10003);
or U12857 (N_12857,N_10939,N_10559);
nand U12858 (N_12858,N_10920,N_9269);
nor U12859 (N_12859,N_9797,N_11722);
nand U12860 (N_12860,N_11237,N_11124);
or U12861 (N_12861,N_9723,N_11094);
nor U12862 (N_12862,N_10950,N_10280);
xor U12863 (N_12863,N_11396,N_10505);
nor U12864 (N_12864,N_9672,N_9584);
nand U12865 (N_12865,N_10893,N_9636);
nand U12866 (N_12866,N_10210,N_10445);
and U12867 (N_12867,N_9042,N_11444);
or U12868 (N_12868,N_9326,N_11190);
nand U12869 (N_12869,N_10816,N_10778);
nand U12870 (N_12870,N_10810,N_9873);
nand U12871 (N_12871,N_9901,N_10381);
or U12872 (N_12872,N_11360,N_10103);
and U12873 (N_12873,N_10147,N_11467);
nand U12874 (N_12874,N_11868,N_11428);
nand U12875 (N_12875,N_9996,N_9225);
nand U12876 (N_12876,N_9341,N_10661);
nand U12877 (N_12877,N_9925,N_10522);
nor U12878 (N_12878,N_9072,N_10478);
or U12879 (N_12879,N_11032,N_9932);
or U12880 (N_12880,N_9462,N_9334);
nor U12881 (N_12881,N_11258,N_9659);
nor U12882 (N_12882,N_11694,N_10898);
or U12883 (N_12883,N_9501,N_11782);
and U12884 (N_12884,N_10667,N_9938);
nand U12885 (N_12885,N_9802,N_9712);
or U12886 (N_12886,N_11768,N_11322);
and U12887 (N_12887,N_10918,N_11059);
nand U12888 (N_12888,N_10971,N_10581);
nor U12889 (N_12889,N_9258,N_9470);
nand U12890 (N_12890,N_11267,N_11545);
nand U12891 (N_12891,N_10694,N_9912);
nand U12892 (N_12892,N_10018,N_11266);
nand U12893 (N_12893,N_9312,N_9609);
nand U12894 (N_12894,N_9212,N_9176);
and U12895 (N_12895,N_11662,N_10093);
nor U12896 (N_12896,N_11522,N_9801);
or U12897 (N_12897,N_11283,N_11107);
and U12898 (N_12898,N_11282,N_9827);
nand U12899 (N_12899,N_10130,N_10655);
nor U12900 (N_12900,N_9814,N_11760);
nand U12901 (N_12901,N_11126,N_10022);
or U12902 (N_12902,N_10025,N_9204);
or U12903 (N_12903,N_9150,N_10818);
or U12904 (N_12904,N_11889,N_11314);
or U12905 (N_12905,N_11525,N_10031);
nand U12906 (N_12906,N_10375,N_10749);
or U12907 (N_12907,N_10125,N_11799);
and U12908 (N_12908,N_9859,N_10690);
and U12909 (N_12909,N_10776,N_11784);
and U12910 (N_12910,N_10380,N_9094);
nor U12911 (N_12911,N_10515,N_9005);
nor U12912 (N_12912,N_10791,N_10941);
nand U12913 (N_12913,N_11198,N_9974);
nand U12914 (N_12914,N_10570,N_11464);
nor U12915 (N_12915,N_9377,N_9175);
nand U12916 (N_12916,N_11250,N_10607);
nor U12917 (N_12917,N_9344,N_9604);
nand U12918 (N_12918,N_11923,N_9534);
or U12919 (N_12919,N_11133,N_10212);
and U12920 (N_12920,N_10676,N_10064);
nor U12921 (N_12921,N_11877,N_9180);
or U12922 (N_12922,N_10448,N_11389);
nor U12923 (N_12923,N_9448,N_11084);
and U12924 (N_12924,N_9086,N_11884);
or U12925 (N_12925,N_9930,N_11436);
nand U12926 (N_12926,N_11215,N_11404);
nand U12927 (N_12927,N_10901,N_10399);
nor U12928 (N_12928,N_9309,N_10370);
and U12929 (N_12929,N_11391,N_11629);
nand U12930 (N_12930,N_10386,N_10718);
and U12931 (N_12931,N_11864,N_10467);
nor U12932 (N_12932,N_9040,N_9266);
nor U12933 (N_12933,N_10197,N_9894);
and U12934 (N_12934,N_9955,N_9280);
or U12935 (N_12935,N_11340,N_9009);
and U12936 (N_12936,N_10908,N_9747);
nand U12937 (N_12937,N_9765,N_9500);
and U12938 (N_12938,N_9695,N_10136);
or U12939 (N_12939,N_9248,N_10926);
nor U12940 (N_12940,N_11732,N_11934);
or U12941 (N_12941,N_9956,N_9908);
nand U12942 (N_12942,N_11947,N_9612);
nand U12943 (N_12943,N_9778,N_11747);
nand U12944 (N_12944,N_11231,N_11442);
and U12945 (N_12945,N_10185,N_9472);
nor U12946 (N_12946,N_11650,N_11541);
or U12947 (N_12947,N_11607,N_9897);
or U12948 (N_12948,N_11091,N_9021);
nand U12949 (N_12949,N_10078,N_9292);
and U12950 (N_12950,N_11516,N_11426);
and U12951 (N_12951,N_11585,N_10398);
nand U12952 (N_12952,N_11117,N_11292);
nand U12953 (N_12953,N_11537,N_10331);
nor U12954 (N_12954,N_11550,N_9975);
nor U12955 (N_12955,N_10692,N_11431);
nor U12956 (N_12956,N_9962,N_11203);
or U12957 (N_12957,N_11703,N_9744);
nand U12958 (N_12958,N_9339,N_11848);
nor U12959 (N_12959,N_10036,N_9918);
and U12960 (N_12960,N_11940,N_10257);
nor U12961 (N_12961,N_10384,N_9979);
nand U12962 (N_12962,N_10389,N_10537);
nand U12963 (N_12963,N_9769,N_9074);
nor U12964 (N_12964,N_11553,N_10838);
or U12965 (N_12965,N_11368,N_11373);
nor U12966 (N_12966,N_9529,N_11121);
nand U12967 (N_12967,N_9862,N_11357);
nor U12968 (N_12968,N_10032,N_10944);
nand U12969 (N_12969,N_9272,N_9601);
or U12970 (N_12970,N_9498,N_9382);
or U12971 (N_12971,N_9052,N_9143);
nand U12972 (N_12972,N_10786,N_11790);
nand U12973 (N_12973,N_10979,N_11527);
nand U12974 (N_12974,N_10007,N_9909);
and U12975 (N_12975,N_11791,N_9546);
nand U12976 (N_12976,N_9621,N_11716);
or U12977 (N_12977,N_9118,N_11182);
or U12978 (N_12978,N_9679,N_9937);
and U12979 (N_12979,N_9638,N_11367);
nand U12980 (N_12980,N_11758,N_11538);
and U12981 (N_12981,N_11468,N_11004);
nand U12982 (N_12982,N_10596,N_9670);
nor U12983 (N_12983,N_10239,N_9959);
nand U12984 (N_12984,N_11901,N_9430);
or U12985 (N_12985,N_10504,N_10423);
or U12986 (N_12986,N_9172,N_10983);
or U12987 (N_12987,N_9928,N_10604);
and U12988 (N_12988,N_9736,N_10033);
nand U12989 (N_12989,N_11278,N_11612);
nor U12990 (N_12990,N_9109,N_11479);
or U12991 (N_12991,N_11013,N_10567);
and U12992 (N_12992,N_9284,N_9607);
or U12993 (N_12993,N_10313,N_11535);
and U12994 (N_12994,N_9179,N_11189);
nor U12995 (N_12995,N_9415,N_11906);
nand U12996 (N_12996,N_11952,N_9944);
nand U12997 (N_12997,N_9075,N_11388);
nand U12998 (N_12998,N_10241,N_11186);
or U12999 (N_12999,N_9570,N_9676);
nand U13000 (N_13000,N_11504,N_10824);
nor U13001 (N_13001,N_10408,N_9876);
nand U13002 (N_13002,N_9438,N_10689);
nand U13003 (N_13003,N_9361,N_11616);
and U13004 (N_13004,N_9328,N_11904);
nand U13005 (N_13005,N_11764,N_10367);
or U13006 (N_13006,N_9719,N_11979);
or U13007 (N_13007,N_10172,N_11896);
or U13008 (N_13008,N_9264,N_10385);
and U13009 (N_13009,N_10065,N_11942);
nor U13010 (N_13010,N_10446,N_10867);
and U13011 (N_13011,N_10630,N_9702);
or U13012 (N_13012,N_9832,N_9054);
nor U13013 (N_13013,N_10773,N_11717);
nand U13014 (N_13014,N_10949,N_10126);
or U13015 (N_13015,N_10240,N_11459);
nor U13016 (N_13016,N_9564,N_11205);
or U13017 (N_13017,N_11271,N_9450);
nand U13018 (N_13018,N_9540,N_9727);
nor U13019 (N_13019,N_9306,N_10363);
nand U13020 (N_13020,N_10145,N_10536);
and U13021 (N_13021,N_9763,N_9526);
nand U13022 (N_13022,N_9016,N_11082);
nor U13023 (N_13023,N_9658,N_11319);
nor U13024 (N_13024,N_9455,N_9069);
or U13025 (N_13025,N_10569,N_11601);
nor U13026 (N_13026,N_10256,N_9586);
or U13027 (N_13027,N_9767,N_11511);
nor U13028 (N_13028,N_9548,N_10890);
nand U13029 (N_13029,N_9026,N_10059);
nand U13030 (N_13030,N_10132,N_11481);
nor U13031 (N_13031,N_9842,N_10549);
or U13032 (N_13032,N_11318,N_11785);
and U13033 (N_13033,N_10682,N_11476);
nor U13034 (N_13034,N_9257,N_11510);
and U13035 (N_13035,N_11230,N_9240);
nor U13036 (N_13036,N_9073,N_11654);
nand U13037 (N_13037,N_10656,N_11222);
nand U13038 (N_13038,N_10098,N_9557);
nand U13039 (N_13039,N_11579,N_11151);
and U13040 (N_13040,N_10143,N_10139);
and U13041 (N_13041,N_9087,N_9653);
nor U13042 (N_13042,N_9871,N_9633);
nand U13043 (N_13043,N_9713,N_11649);
nand U13044 (N_13044,N_9716,N_11177);
nor U13045 (N_13045,N_10647,N_10244);
nand U13046 (N_13046,N_10555,N_9124);
nor U13047 (N_13047,N_10039,N_9023);
nor U13048 (N_13048,N_11438,N_11221);
nor U13049 (N_13049,N_10068,N_10588);
nor U13050 (N_13050,N_10525,N_11247);
or U13051 (N_13051,N_9637,N_11870);
and U13052 (N_13052,N_9760,N_10072);
xnor U13053 (N_13053,N_10666,N_10076);
nor U13054 (N_13054,N_11891,N_9155);
and U13055 (N_13055,N_9618,N_11332);
or U13056 (N_13056,N_10029,N_10731);
and U13057 (N_13057,N_11308,N_9844);
nand U13058 (N_13058,N_11307,N_9817);
nand U13059 (N_13059,N_9575,N_10848);
nor U13060 (N_13060,N_9904,N_10917);
or U13061 (N_13061,N_10317,N_9432);
and U13062 (N_13062,N_11655,N_10836);
nand U13063 (N_13063,N_9229,N_10315);
or U13064 (N_13064,N_10450,N_11640);
or U13065 (N_13065,N_10668,N_10708);
and U13066 (N_13066,N_11156,N_11845);
nand U13067 (N_13067,N_11412,N_10705);
nand U13068 (N_13068,N_9588,N_11536);
nor U13069 (N_13069,N_9406,N_11632);
and U13070 (N_13070,N_10730,N_9332);
and U13071 (N_13071,N_11829,N_11518);
nand U13072 (N_13072,N_10207,N_9983);
or U13073 (N_13073,N_11862,N_11931);
and U13074 (N_13074,N_9033,N_9690);
or U13075 (N_13075,N_11125,N_10813);
and U13076 (N_13076,N_10083,N_10710);
nand U13077 (N_13077,N_9835,N_10933);
or U13078 (N_13078,N_10168,N_10955);
nand U13079 (N_13079,N_9449,N_10014);
nor U13080 (N_13080,N_9350,N_10557);
or U13081 (N_13081,N_11001,N_10138);
nand U13082 (N_13082,N_11597,N_11676);
or U13083 (N_13083,N_9467,N_9796);
nor U13084 (N_13084,N_9632,N_9759);
nor U13085 (N_13085,N_9836,N_9999);
nor U13086 (N_13086,N_10987,N_11218);
nand U13087 (N_13087,N_9569,N_11458);
or U13088 (N_13088,N_11954,N_11216);
nor U13089 (N_13089,N_9019,N_11255);
nor U13090 (N_13090,N_11528,N_11154);
nor U13091 (N_13091,N_11086,N_9135);
nor U13092 (N_13092,N_9954,N_10320);
or U13093 (N_13093,N_9254,N_9869);
nor U13094 (N_13094,N_9421,N_9590);
and U13095 (N_13095,N_10468,N_9581);
or U13096 (N_13096,N_9920,N_9772);
nor U13097 (N_13097,N_11400,N_10750);
nor U13098 (N_13098,N_9336,N_10539);
and U13099 (N_13099,N_9539,N_10814);
or U13100 (N_13100,N_9552,N_10576);
nor U13101 (N_13101,N_9851,N_10598);
or U13102 (N_13102,N_11617,N_11098);
or U13103 (N_13103,N_10584,N_11879);
or U13104 (N_13104,N_10334,N_9121);
nor U13105 (N_13105,N_11571,N_11898);
nor U13106 (N_13106,N_9519,N_9030);
nand U13107 (N_13107,N_9514,N_11721);
or U13108 (N_13108,N_10964,N_10500);
and U13109 (N_13109,N_11070,N_10297);
and U13110 (N_13110,N_11946,N_9574);
and U13111 (N_13111,N_10443,N_9136);
nand U13112 (N_13112,N_10507,N_9131);
and U13113 (N_13113,N_11542,N_9233);
nor U13114 (N_13114,N_11170,N_11276);
nand U13115 (N_13115,N_9028,N_9663);
nor U13116 (N_13116,N_10980,N_11440);
or U13117 (N_13117,N_11735,N_10020);
or U13118 (N_13118,N_9895,N_10357);
and U13119 (N_13119,N_10208,N_11804);
nand U13120 (N_13120,N_10788,N_11257);
and U13121 (N_13121,N_11724,N_10618);
nand U13122 (N_13122,N_10911,N_10612);
nand U13123 (N_13123,N_11797,N_10476);
or U13124 (N_13124,N_10874,N_10390);
or U13125 (N_13125,N_9800,N_10181);
or U13126 (N_13126,N_11820,N_9900);
or U13127 (N_13127,N_9742,N_10052);
or U13128 (N_13128,N_11140,N_9958);
nand U13129 (N_13129,N_9392,N_9238);
or U13130 (N_13130,N_11462,N_10711);
and U13131 (N_13131,N_9315,N_9181);
and U13132 (N_13132,N_10967,N_10473);
nor U13133 (N_13133,N_10931,N_11989);
nand U13134 (N_13134,N_11987,N_11220);
nor U13135 (N_13135,N_10713,N_11572);
or U13136 (N_13136,N_11260,N_10510);
nor U13137 (N_13137,N_10947,N_11595);
and U13138 (N_13138,N_9881,N_9110);
and U13139 (N_13139,N_10660,N_9165);
or U13140 (N_13140,N_11207,N_10431);
nand U13141 (N_13141,N_10905,N_10162);
nor U13142 (N_13142,N_10496,N_10709);
or U13143 (N_13143,N_9177,N_9997);
and U13144 (N_13144,N_9314,N_11063);
nand U13145 (N_13145,N_11381,N_9045);
nor U13146 (N_13146,N_11917,N_11574);
nand U13147 (N_13147,N_11058,N_10999);
or U13148 (N_13148,N_11365,N_11606);
nor U13149 (N_13149,N_11043,N_9089);
nand U13150 (N_13150,N_10961,N_11661);
xnor U13151 (N_13151,N_11128,N_11009);
and U13152 (N_13152,N_9947,N_11311);
and U13153 (N_13153,N_11921,N_9327);
and U13154 (N_13154,N_10097,N_9007);
and U13155 (N_13155,N_11329,N_9231);
or U13156 (N_13156,N_11513,N_11853);
nor U13157 (N_13157,N_11982,N_11174);
nand U13158 (N_13158,N_10153,N_9098);
nor U13159 (N_13159,N_11708,N_10990);
nand U13160 (N_13160,N_9594,N_10761);
nor U13161 (N_13161,N_9345,N_9290);
and U13162 (N_13162,N_9085,N_9988);
xnor U13163 (N_13163,N_11614,N_11656);
or U13164 (N_13164,N_11097,N_10416);
nor U13165 (N_13165,N_11165,N_9661);
nand U13166 (N_13166,N_10956,N_9771);
and U13167 (N_13167,N_10226,N_9425);
or U13168 (N_13168,N_11996,N_9243);
and U13169 (N_13169,N_10323,N_9387);
or U13170 (N_13170,N_10800,N_9489);
nor U13171 (N_13171,N_11852,N_9103);
nor U13172 (N_13172,N_9084,N_9161);
and U13173 (N_13173,N_10079,N_9174);
nor U13174 (N_13174,N_10679,N_9105);
or U13175 (N_13175,N_9195,N_10906);
nand U13176 (N_13176,N_11613,N_11874);
nand U13177 (N_13177,N_11828,N_10523);
nor U13178 (N_13178,N_9373,N_11208);
or U13179 (N_13179,N_10962,N_11514);
or U13180 (N_13180,N_9682,N_10839);
and U13181 (N_13181,N_11666,N_11670);
or U13182 (N_13182,N_10946,N_9492);
or U13183 (N_13183,N_10092,N_11668);
and U13184 (N_13184,N_10017,N_9113);
nor U13185 (N_13185,N_10155,N_9834);
and U13186 (N_13186,N_10747,N_11972);
or U13187 (N_13187,N_10268,N_10238);
nor U13188 (N_13188,N_11665,N_11147);
or U13189 (N_13189,N_9058,N_10974);
and U13190 (N_13190,N_10264,N_11213);
nor U13191 (N_13191,N_9270,N_10913);
nor U13192 (N_13192,N_11554,N_10289);
or U13193 (N_13193,N_9718,N_11254);
and U13194 (N_13194,N_10169,N_10527);
and U13195 (N_13195,N_11714,N_10215);
and U13196 (N_13196,N_9692,N_9976);
or U13197 (N_13197,N_10645,N_9628);
nand U13198 (N_13198,N_11472,N_11847);
and U13199 (N_13199,N_9649,N_10290);
nand U13200 (N_13200,N_9171,N_11214);
nor U13201 (N_13201,N_10755,N_9890);
nand U13202 (N_13202,N_9503,N_11399);
nand U13203 (N_13203,N_10379,N_10470);
or U13204 (N_13204,N_9686,N_9206);
nand U13205 (N_13205,N_10972,N_9435);
nand U13206 (N_13206,N_9066,N_9651);
or U13207 (N_13207,N_11978,N_9730);
nor U13208 (N_13208,N_11265,N_9041);
or U13209 (N_13209,N_10595,N_9183);
nand U13210 (N_13210,N_9274,N_10871);
nor U13211 (N_13211,N_11517,N_11826);
and U13212 (N_13212,N_10831,N_10485);
or U13213 (N_13213,N_9942,N_9267);
nor U13214 (N_13214,N_10436,N_11418);
nor U13215 (N_13215,N_11330,N_10650);
nand U13216 (N_13216,N_11460,N_9048);
and U13217 (N_13217,N_10978,N_11015);
nor U13218 (N_13218,N_11419,N_9511);
nor U13219 (N_13219,N_11089,N_10271);
and U13220 (N_13220,N_9829,N_11115);
and U13221 (N_13221,N_10764,N_10879);
nand U13222 (N_13222,N_9379,N_10475);
and U13223 (N_13223,N_11240,N_11809);
nor U13224 (N_13224,N_10114,N_9549);
nor U13225 (N_13225,N_10150,N_9408);
nor U13226 (N_13226,N_11183,N_11313);
or U13227 (N_13227,N_11206,N_11243);
and U13228 (N_13228,N_11315,N_9915);
or U13229 (N_13229,N_11263,N_10844);
nor U13230 (N_13230,N_10019,N_9917);
nand U13231 (N_13231,N_9083,N_9635);
and U13232 (N_13232,N_10637,N_9122);
nand U13233 (N_13233,N_11072,N_9138);
or U13234 (N_13234,N_10425,N_11509);
nor U13235 (N_13235,N_10624,N_10158);
nand U13236 (N_13236,N_9167,N_10410);
nand U13237 (N_13237,N_10213,N_10174);
nand U13238 (N_13238,N_9029,N_11914);
nor U13239 (N_13239,N_10220,N_10702);
or U13240 (N_13240,N_11644,N_11748);
xor U13241 (N_13241,N_9994,N_9750);
and U13242 (N_13242,N_10991,N_10669);
or U13243 (N_13243,N_10699,N_10413);
or U13244 (N_13244,N_10724,N_9353);
nand U13245 (N_13245,N_11945,N_10988);
nand U13246 (N_13246,N_10131,N_9452);
or U13247 (N_13247,N_9133,N_11409);
or U13248 (N_13248,N_10382,N_9543);
nor U13249 (N_13249,N_10402,N_9340);
and U13250 (N_13250,N_10349,N_10091);
nand U13251 (N_13251,N_10344,N_11970);
or U13252 (N_13252,N_9268,N_10680);
nor U13253 (N_13253,N_11350,N_11846);
nand U13254 (N_13254,N_10447,N_11854);
nand U13255 (N_13255,N_9721,N_9461);
and U13256 (N_13256,N_11211,N_10236);
nor U13257 (N_13257,N_10916,N_9950);
nor U13258 (N_13258,N_9731,N_10803);
xnor U13259 (N_13259,N_11048,N_11331);
and U13260 (N_13260,N_9860,N_11348);
nor U13261 (N_13261,N_10119,N_9846);
nand U13262 (N_13262,N_11323,N_11455);
nand U13263 (N_13263,N_10177,N_10404);
or U13264 (N_13264,N_10687,N_9106);
nor U13265 (N_13265,N_10681,N_9239);
or U13266 (N_13266,N_11894,N_9886);
or U13267 (N_13267,N_9499,N_10489);
or U13268 (N_13268,N_9532,N_9311);
nor U13269 (N_13269,N_11080,N_11792);
nor U13270 (N_13270,N_11709,N_11184);
or U13271 (N_13271,N_10427,N_11769);
xor U13272 (N_13272,N_11397,N_10287);
nor U13273 (N_13273,N_10499,N_10149);
nor U13274 (N_13274,N_11273,N_10460);
nand U13275 (N_13275,N_9391,N_9732);
and U13276 (N_13276,N_9815,N_9001);
or U13277 (N_13277,N_10945,N_11555);
or U13278 (N_13278,N_10170,N_11699);
nor U13279 (N_13279,N_11416,N_9156);
nand U13280 (N_13280,N_10360,N_9128);
nor U13281 (N_13281,N_9751,N_10233);
and U13282 (N_13282,N_10471,N_10288);
or U13283 (N_13283,N_9902,N_11228);
and U13284 (N_13284,N_10862,N_11800);
and U13285 (N_13285,N_11990,N_9669);
and U13286 (N_13286,N_11446,N_10248);
nor U13287 (N_13287,N_9245,N_10463);
or U13288 (N_13288,N_11333,N_9807);
nand U13289 (N_13289,N_11729,N_9348);
nor U13290 (N_13290,N_10112,N_11474);
nor U13291 (N_13291,N_9265,N_9469);
nand U13292 (N_13292,N_10670,N_10552);
and U13293 (N_13293,N_11673,N_10183);
nor U13294 (N_13294,N_10629,N_10111);
nor U13295 (N_13295,N_9413,N_10571);
nor U13296 (N_13296,N_11114,N_9236);
or U13297 (N_13297,N_9355,N_11326);
nand U13298 (N_13298,N_11338,N_11490);
nor U13299 (N_13299,N_11407,N_9752);
nand U13300 (N_13300,N_11502,N_10644);
or U13301 (N_13301,N_9184,N_10957);
nor U13302 (N_13302,N_9119,N_11405);
nand U13303 (N_13303,N_11802,N_11986);
nor U13304 (N_13304,N_10613,N_10296);
nand U13305 (N_13305,N_9745,N_10678);
or U13306 (N_13306,N_9952,N_9352);
or U13307 (N_13307,N_9034,N_10283);
nor U13308 (N_13308,N_11312,N_10284);
nor U13309 (N_13309,N_10165,N_10542);
nand U13310 (N_13310,N_10556,N_10881);
nand U13311 (N_13311,N_10992,N_10180);
and U13312 (N_13312,N_11137,N_11142);
or U13313 (N_13313,N_10043,N_9289);
and U13314 (N_13314,N_9012,N_10328);
nor U13315 (N_13315,N_11286,N_11269);
and U13316 (N_13316,N_10615,N_10738);
nor U13317 (N_13317,N_10583,N_9644);
nor U13318 (N_13318,N_10235,N_11202);
or U13319 (N_13319,N_11723,N_9191);
nand U13320 (N_13320,N_10341,N_11794);
and U13321 (N_13321,N_9818,N_10574);
and U13322 (N_13322,N_9507,N_10400);
nor U13323 (N_13323,N_9393,N_10329);
nand U13324 (N_13324,N_11526,N_11150);
nand U13325 (N_13325,N_9193,N_10513);
or U13326 (N_13326,N_11966,N_11816);
and U13327 (N_13327,N_9949,N_10122);
nor U13328 (N_13328,N_10745,N_10133);
nor U13329 (N_13329,N_11175,N_10082);
nand U13330 (N_13330,N_10821,N_10568);
and U13331 (N_13331,N_10144,N_10753);
or U13332 (N_13332,N_9251,N_11583);
nand U13333 (N_13333,N_11680,N_11592);
nand U13334 (N_13334,N_9813,N_10491);
and U13335 (N_13335,N_11393,N_10799);
and U13336 (N_13336,N_10759,N_10777);
nor U13337 (N_13337,N_9940,N_9038);
nor U13338 (N_13338,N_10434,N_11733);
or U13339 (N_13339,N_11838,N_10405);
nand U13340 (N_13340,N_9305,N_10817);
nand U13341 (N_13341,N_10351,N_9010);
or U13342 (N_13342,N_10187,N_9717);
nand U13343 (N_13343,N_9490,N_11817);
or U13344 (N_13344,N_11234,N_9625);
nor U13345 (N_13345,N_11310,N_11836);
and U13346 (N_13346,N_11078,N_11127);
or U13347 (N_13347,N_10765,N_10211);
nor U13348 (N_13348,N_9429,N_11731);
xor U13349 (N_13349,N_10981,N_10319);
nand U13350 (N_13350,N_10880,N_11095);
and U13351 (N_13351,N_9906,N_10605);
and U13352 (N_13352,N_9277,N_11956);
nor U13353 (N_13353,N_11765,N_10255);
and U13354 (N_13354,N_9536,N_10095);
or U13355 (N_13355,N_9321,N_10016);
and U13356 (N_13356,N_10997,N_10260);
nand U13357 (N_13357,N_11414,N_10892);
nor U13358 (N_13358,N_9794,N_9216);
and U13359 (N_13359,N_9453,N_11047);
or U13360 (N_13360,N_9914,N_11103);
or U13361 (N_13361,N_11083,N_9710);
or U13362 (N_13362,N_9720,N_9722);
or U13363 (N_13363,N_10601,N_10876);
and U13364 (N_13364,N_11343,N_11423);
and U13365 (N_13365,N_9831,N_9035);
nand U13366 (N_13366,N_10160,N_9368);
nor U13367 (N_13367,N_11631,N_11962);
and U13368 (N_13368,N_10301,N_10184);
and U13369 (N_13369,N_11652,N_9337);
or U13370 (N_13370,N_9743,N_11060);
nand U13371 (N_13371,N_9849,N_9145);
nand U13372 (N_13372,N_10683,N_9992);
nand U13373 (N_13373,N_11696,N_10520);
nand U13374 (N_13374,N_9279,N_11604);
nor U13375 (N_13375,N_10024,N_9689);
nand U13376 (N_13376,N_11780,N_10110);
nand U13377 (N_13377,N_10545,N_9926);
nor U13378 (N_13378,N_11204,N_10252);
and U13379 (N_13379,N_9755,N_10832);
nor U13380 (N_13380,N_9905,N_10744);
nand U13381 (N_13381,N_10224,N_11225);
nor U13382 (N_13382,N_10182,N_10214);
and U13383 (N_13383,N_11890,N_9067);
nand U13384 (N_13384,N_9194,N_9623);
and U13385 (N_13385,N_10621,N_11557);
or U13386 (N_13386,N_11040,N_11224);
nor U13387 (N_13387,N_11454,N_11559);
nor U13388 (N_13388,N_9062,N_11317);
nor U13389 (N_13389,N_10691,N_10589);
nand U13390 (N_13390,N_10311,N_11766);
or U13391 (N_13391,N_11109,N_10502);
or U13392 (N_13392,N_10952,N_10609);
and U13393 (N_13393,N_10462,N_11738);
nand U13394 (N_13394,N_11498,N_10751);
nor U13395 (N_13395,N_9210,N_9319);
nor U13396 (N_13396,N_11347,N_9910);
and U13397 (N_13397,N_11489,N_9547);
or U13398 (N_13398,N_9995,N_11275);
and U13399 (N_13399,N_9077,N_10455);
nor U13400 (N_13400,N_9065,N_11046);
and U13401 (N_13401,N_10243,N_9357);
or U13402 (N_13402,N_10449,N_9714);
or U13403 (N_13403,N_11337,N_9427);
and U13404 (N_13404,N_10051,N_9528);
nor U13405 (N_13405,N_10453,N_9830);
nor U13406 (N_13406,N_10189,N_9022);
or U13407 (N_13407,N_11963,N_11695);
xor U13408 (N_13408,N_10474,N_10729);
xor U13409 (N_13409,N_11453,N_10812);
nor U13410 (N_13410,N_11328,N_10487);
or U13411 (N_13411,N_11876,N_9648);
nand U13412 (N_13412,N_9991,N_10868);
nand U13413 (N_13413,N_10701,N_9520);
and U13414 (N_13414,N_10953,N_10998);
and U13415 (N_13415,N_11327,N_9403);
nor U13416 (N_13416,N_11615,N_11144);
nor U13417 (N_13417,N_10873,N_9017);
nand U13418 (N_13418,N_11971,N_11039);
nor U13419 (N_13419,N_11857,N_11188);
or U13420 (N_13420,N_11377,N_11692);
nand U13421 (N_13421,N_10206,N_9513);
nand U13422 (N_13422,N_11181,N_10094);
and U13423 (N_13423,N_10772,N_11573);
nor U13424 (N_13424,N_9561,N_10322);
nand U13425 (N_13425,N_10828,N_11073);
and U13426 (N_13426,N_11057,N_9681);
or U13427 (N_13427,N_11155,N_11402);
or U13428 (N_13428,N_9375,N_10071);
and U13429 (N_13429,N_9100,N_9294);
and U13430 (N_13430,N_9811,N_9296);
or U13431 (N_13431,N_9253,N_9629);
nand U13432 (N_13432,N_9082,N_9708);
nor U13433 (N_13433,N_10915,N_10732);
nand U13434 (N_13434,N_9841,N_9657);
nor U13435 (N_13435,N_11599,N_9404);
and U13436 (N_13436,N_11153,N_10610);
or U13437 (N_13437,N_10310,N_10671);
and U13438 (N_13438,N_9214,N_9218);
nor U13439 (N_13439,N_10780,N_9872);
nor U13440 (N_13440,N_9591,N_10063);
nor U13441 (N_13441,N_9209,N_10768);
nand U13442 (N_13442,N_10285,N_10907);
nor U13443 (N_13443,N_11112,N_11660);
or U13444 (N_13444,N_10451,N_9598);
and U13445 (N_13445,N_10305,N_10274);
and U13446 (N_13446,N_11284,N_10242);
nor U13447 (N_13447,N_9973,N_9015);
nand U13448 (N_13448,N_11118,N_10697);
nor U13449 (N_13449,N_11533,N_10272);
nand U13450 (N_13450,N_10013,N_11272);
nor U13451 (N_13451,N_10440,N_9092);
and U13452 (N_13452,N_9463,N_9533);
nor U13453 (N_13453,N_9275,N_9577);
and U13454 (N_13454,N_10194,N_9338);
or U13455 (N_13455,N_9855,N_10565);
nor U13456 (N_13456,N_9787,N_10354);
and U13457 (N_13457,N_10841,N_9496);
or U13458 (N_13458,N_11376,N_11429);
or U13459 (N_13459,N_11580,N_10805);
or U13460 (N_13460,N_9208,N_10414);
nand U13461 (N_13461,N_10326,N_11356);
and U13462 (N_13462,N_10225,N_11752);
nand U13463 (N_13463,N_9773,N_11787);
xor U13464 (N_13464,N_10514,N_10442);
nor U13465 (N_13465,N_10993,N_11485);
xnor U13466 (N_13466,N_10101,N_10167);
nor U13467 (N_13467,N_9050,N_10292);
nor U13468 (N_13468,N_10038,N_10606);
nor U13469 (N_13469,N_9263,N_11161);
or U13470 (N_13470,N_10429,N_10912);
nand U13471 (N_13471,N_11757,N_10457);
and U13472 (N_13472,N_11888,N_11964);
or U13473 (N_13473,N_10259,N_11623);
nand U13474 (N_13474,N_11851,N_9675);
or U13475 (N_13475,N_10490,N_11452);
nor U13476 (N_13476,N_11983,N_11600);
and U13477 (N_13477,N_9115,N_9096);
or U13478 (N_13478,N_11568,N_11910);
nor U13479 (N_13479,N_9173,N_11958);
nand U13480 (N_13480,N_11674,N_11021);
or U13481 (N_13481,N_9410,N_10361);
nand U13482 (N_13482,N_10498,N_9146);
nor U13483 (N_13483,N_11909,N_9508);
nor U13484 (N_13484,N_10249,N_10614);
or U13485 (N_13485,N_9611,N_10648);
nor U13486 (N_13486,N_11441,N_10107);
or U13487 (N_13487,N_11433,N_9515);
nand U13488 (N_13488,N_11421,N_11301);
nand U13489 (N_13489,N_9891,N_10544);
or U13490 (N_13490,N_9451,N_9307);
and U13491 (N_13491,N_11628,N_9848);
nand U13492 (N_13492,N_10503,N_11209);
nand U13493 (N_13493,N_9544,N_9199);
nor U13494 (N_13494,N_10808,N_9141);
nand U13495 (N_13495,N_10237,N_9645);
nand U13496 (N_13496,N_11178,N_10362);
or U13497 (N_13497,N_9524,N_11288);
and U13498 (N_13498,N_11540,N_11068);
or U13499 (N_13499,N_11104,N_9376);
or U13500 (N_13500,N_9591,N_9570);
nor U13501 (N_13501,N_11217,N_11851);
and U13502 (N_13502,N_11223,N_9074);
nand U13503 (N_13503,N_11925,N_11320);
and U13504 (N_13504,N_11637,N_11478);
nor U13505 (N_13505,N_9178,N_11951);
or U13506 (N_13506,N_11115,N_11153);
and U13507 (N_13507,N_11204,N_10542);
nand U13508 (N_13508,N_10890,N_11865);
nand U13509 (N_13509,N_11815,N_9238);
nor U13510 (N_13510,N_11913,N_10247);
and U13511 (N_13511,N_9361,N_9472);
and U13512 (N_13512,N_9915,N_10304);
nor U13513 (N_13513,N_11299,N_11307);
nand U13514 (N_13514,N_10786,N_11594);
or U13515 (N_13515,N_11177,N_9834);
or U13516 (N_13516,N_9379,N_10654);
and U13517 (N_13517,N_11034,N_9107);
or U13518 (N_13518,N_9645,N_10491);
nand U13519 (N_13519,N_11541,N_11269);
and U13520 (N_13520,N_11802,N_11485);
and U13521 (N_13521,N_10448,N_11579);
nand U13522 (N_13522,N_10336,N_11823);
nor U13523 (N_13523,N_11971,N_10860);
nand U13524 (N_13524,N_10256,N_10925);
nor U13525 (N_13525,N_10809,N_9816);
and U13526 (N_13526,N_10850,N_10348);
nand U13527 (N_13527,N_10216,N_10247);
nor U13528 (N_13528,N_11923,N_9144);
or U13529 (N_13529,N_9503,N_10436);
nand U13530 (N_13530,N_9253,N_9037);
nand U13531 (N_13531,N_11776,N_9961);
nand U13532 (N_13532,N_10107,N_11370);
and U13533 (N_13533,N_9860,N_10320);
and U13534 (N_13534,N_11131,N_10314);
and U13535 (N_13535,N_9732,N_10287);
or U13536 (N_13536,N_10948,N_11565);
nand U13537 (N_13537,N_9801,N_9302);
and U13538 (N_13538,N_11565,N_10920);
or U13539 (N_13539,N_9599,N_9579);
and U13540 (N_13540,N_11072,N_10016);
nand U13541 (N_13541,N_11284,N_10771);
and U13542 (N_13542,N_9892,N_11901);
nand U13543 (N_13543,N_10098,N_9263);
and U13544 (N_13544,N_11782,N_11277);
or U13545 (N_13545,N_10340,N_10856);
nand U13546 (N_13546,N_10592,N_10325);
nor U13547 (N_13547,N_9163,N_9087);
nand U13548 (N_13548,N_11847,N_11263);
nor U13549 (N_13549,N_10024,N_9329);
nor U13550 (N_13550,N_9150,N_10950);
or U13551 (N_13551,N_10516,N_11939);
and U13552 (N_13552,N_9139,N_11984);
nand U13553 (N_13553,N_10328,N_11210);
nor U13554 (N_13554,N_10946,N_9255);
nand U13555 (N_13555,N_11144,N_11488);
nor U13556 (N_13556,N_9053,N_10065);
or U13557 (N_13557,N_10721,N_10688);
nor U13558 (N_13558,N_11255,N_10808);
nand U13559 (N_13559,N_10241,N_9341);
or U13560 (N_13560,N_9389,N_11274);
nor U13561 (N_13561,N_9196,N_9753);
nand U13562 (N_13562,N_10725,N_10097);
or U13563 (N_13563,N_11412,N_11752);
and U13564 (N_13564,N_9130,N_9044);
nand U13565 (N_13565,N_11386,N_10323);
nand U13566 (N_13566,N_9395,N_10626);
and U13567 (N_13567,N_10684,N_10067);
nand U13568 (N_13568,N_9036,N_9679);
and U13569 (N_13569,N_11666,N_11482);
nor U13570 (N_13570,N_10507,N_11337);
and U13571 (N_13571,N_10219,N_9962);
nor U13572 (N_13572,N_10991,N_9425);
or U13573 (N_13573,N_10367,N_9187);
or U13574 (N_13574,N_9087,N_11575);
or U13575 (N_13575,N_9468,N_9806);
nor U13576 (N_13576,N_11472,N_10670);
nor U13577 (N_13577,N_10487,N_11089);
or U13578 (N_13578,N_11068,N_9651);
or U13579 (N_13579,N_10208,N_10808);
nand U13580 (N_13580,N_9088,N_9776);
and U13581 (N_13581,N_10975,N_11610);
xor U13582 (N_13582,N_10092,N_11581);
or U13583 (N_13583,N_9480,N_10298);
nor U13584 (N_13584,N_10849,N_10561);
nor U13585 (N_13585,N_10164,N_9925);
nand U13586 (N_13586,N_10716,N_9948);
and U13587 (N_13587,N_10610,N_10533);
nand U13588 (N_13588,N_9858,N_11749);
or U13589 (N_13589,N_9330,N_10856);
and U13590 (N_13590,N_9741,N_9611);
nor U13591 (N_13591,N_11807,N_10215);
nor U13592 (N_13592,N_10916,N_11127);
nor U13593 (N_13593,N_11163,N_9103);
or U13594 (N_13594,N_9238,N_9380);
or U13595 (N_13595,N_11199,N_10591);
nand U13596 (N_13596,N_11207,N_10928);
or U13597 (N_13597,N_11491,N_10993);
nor U13598 (N_13598,N_11690,N_10061);
and U13599 (N_13599,N_9074,N_9472);
nand U13600 (N_13600,N_9166,N_9993);
and U13601 (N_13601,N_9604,N_9448);
nand U13602 (N_13602,N_10117,N_9400);
or U13603 (N_13603,N_9329,N_10061);
or U13604 (N_13604,N_10895,N_11064);
and U13605 (N_13605,N_10113,N_9941);
nand U13606 (N_13606,N_11937,N_11417);
xnor U13607 (N_13607,N_10796,N_10140);
nand U13608 (N_13608,N_10893,N_9075);
nand U13609 (N_13609,N_9747,N_9289);
nor U13610 (N_13610,N_9985,N_10451);
and U13611 (N_13611,N_10484,N_9722);
and U13612 (N_13612,N_11374,N_10106);
nor U13613 (N_13613,N_9815,N_10484);
or U13614 (N_13614,N_9835,N_9427);
nor U13615 (N_13615,N_9444,N_9175);
nor U13616 (N_13616,N_11125,N_11395);
or U13617 (N_13617,N_11223,N_10334);
or U13618 (N_13618,N_10253,N_10213);
or U13619 (N_13619,N_10207,N_9605);
nand U13620 (N_13620,N_9449,N_11608);
nor U13621 (N_13621,N_11784,N_11672);
nand U13622 (N_13622,N_10520,N_9655);
and U13623 (N_13623,N_10455,N_9025);
nand U13624 (N_13624,N_11533,N_9546);
nand U13625 (N_13625,N_11473,N_11661);
and U13626 (N_13626,N_9613,N_10226);
nand U13627 (N_13627,N_10040,N_9016);
nor U13628 (N_13628,N_9862,N_10762);
and U13629 (N_13629,N_9799,N_11274);
and U13630 (N_13630,N_9069,N_9271);
nor U13631 (N_13631,N_9783,N_9615);
nor U13632 (N_13632,N_10742,N_11620);
nand U13633 (N_13633,N_10917,N_9469);
nand U13634 (N_13634,N_11665,N_9315);
or U13635 (N_13635,N_10238,N_10774);
nor U13636 (N_13636,N_10285,N_10182);
and U13637 (N_13637,N_10642,N_10151);
nor U13638 (N_13638,N_11259,N_9465);
nand U13639 (N_13639,N_11173,N_10772);
nand U13640 (N_13640,N_10585,N_9600);
nor U13641 (N_13641,N_10151,N_9688);
nor U13642 (N_13642,N_11269,N_11623);
and U13643 (N_13643,N_11573,N_9449);
and U13644 (N_13644,N_9830,N_10463);
nand U13645 (N_13645,N_9740,N_11313);
nand U13646 (N_13646,N_9177,N_9150);
nand U13647 (N_13647,N_10742,N_10761);
nor U13648 (N_13648,N_9907,N_11341);
or U13649 (N_13649,N_9086,N_9835);
and U13650 (N_13650,N_10445,N_11193);
or U13651 (N_13651,N_11164,N_10806);
or U13652 (N_13652,N_9652,N_10227);
and U13653 (N_13653,N_9755,N_9809);
or U13654 (N_13654,N_9054,N_10736);
nor U13655 (N_13655,N_9595,N_10970);
and U13656 (N_13656,N_10781,N_10198);
and U13657 (N_13657,N_10414,N_11207);
nand U13658 (N_13658,N_9409,N_10381);
nor U13659 (N_13659,N_11125,N_10459);
or U13660 (N_13660,N_11370,N_11928);
and U13661 (N_13661,N_9645,N_10499);
nand U13662 (N_13662,N_9170,N_10685);
or U13663 (N_13663,N_11963,N_10981);
or U13664 (N_13664,N_9817,N_10454);
and U13665 (N_13665,N_10464,N_11505);
or U13666 (N_13666,N_9488,N_11799);
or U13667 (N_13667,N_11421,N_11859);
xnor U13668 (N_13668,N_11047,N_9938);
nor U13669 (N_13669,N_11809,N_9945);
and U13670 (N_13670,N_11934,N_9287);
nor U13671 (N_13671,N_11895,N_10887);
or U13672 (N_13672,N_10872,N_10288);
nor U13673 (N_13673,N_10702,N_9128);
nand U13674 (N_13674,N_10551,N_10614);
or U13675 (N_13675,N_9593,N_10930);
or U13676 (N_13676,N_11961,N_9855);
nor U13677 (N_13677,N_9586,N_9788);
and U13678 (N_13678,N_10130,N_11022);
and U13679 (N_13679,N_9833,N_10943);
or U13680 (N_13680,N_10198,N_10490);
or U13681 (N_13681,N_9450,N_11049);
nor U13682 (N_13682,N_10905,N_9856);
or U13683 (N_13683,N_9057,N_9125);
nand U13684 (N_13684,N_9330,N_11899);
or U13685 (N_13685,N_9813,N_11983);
and U13686 (N_13686,N_11402,N_11844);
and U13687 (N_13687,N_10822,N_9510);
nor U13688 (N_13688,N_9518,N_9752);
nand U13689 (N_13689,N_10367,N_11887);
and U13690 (N_13690,N_10958,N_9424);
nor U13691 (N_13691,N_9264,N_9447);
nand U13692 (N_13692,N_11004,N_10483);
nand U13693 (N_13693,N_10813,N_9574);
or U13694 (N_13694,N_10236,N_9003);
and U13695 (N_13695,N_10638,N_9254);
nand U13696 (N_13696,N_11743,N_10697);
xnor U13697 (N_13697,N_10634,N_10684);
or U13698 (N_13698,N_9779,N_10164);
and U13699 (N_13699,N_10293,N_10319);
and U13700 (N_13700,N_11699,N_11301);
and U13701 (N_13701,N_10986,N_11115);
or U13702 (N_13702,N_11724,N_10489);
or U13703 (N_13703,N_11187,N_10312);
nand U13704 (N_13704,N_9403,N_9189);
and U13705 (N_13705,N_11501,N_10641);
or U13706 (N_13706,N_11184,N_10304);
nand U13707 (N_13707,N_11119,N_11606);
nor U13708 (N_13708,N_11880,N_10990);
nand U13709 (N_13709,N_11515,N_11659);
and U13710 (N_13710,N_10498,N_10927);
or U13711 (N_13711,N_10306,N_10529);
or U13712 (N_13712,N_9414,N_9112);
nor U13713 (N_13713,N_11041,N_9788);
nand U13714 (N_13714,N_9647,N_9272);
nand U13715 (N_13715,N_10589,N_11826);
or U13716 (N_13716,N_11443,N_10614);
nor U13717 (N_13717,N_10090,N_9488);
nand U13718 (N_13718,N_9339,N_10588);
or U13719 (N_13719,N_11047,N_11028);
nand U13720 (N_13720,N_11051,N_11002);
and U13721 (N_13721,N_11800,N_11462);
and U13722 (N_13722,N_11740,N_11491);
nand U13723 (N_13723,N_10712,N_9698);
nand U13724 (N_13724,N_11951,N_9021);
nand U13725 (N_13725,N_11812,N_11852);
nor U13726 (N_13726,N_9765,N_9767);
or U13727 (N_13727,N_10605,N_10657);
or U13728 (N_13728,N_9288,N_9813);
nor U13729 (N_13729,N_11182,N_9313);
or U13730 (N_13730,N_9102,N_11303);
nand U13731 (N_13731,N_9081,N_9128);
nor U13732 (N_13732,N_9769,N_11287);
and U13733 (N_13733,N_10057,N_9850);
nor U13734 (N_13734,N_11671,N_10309);
and U13735 (N_13735,N_11734,N_11443);
and U13736 (N_13736,N_11880,N_10443);
and U13737 (N_13737,N_11635,N_10867);
nand U13738 (N_13738,N_9840,N_11240);
and U13739 (N_13739,N_10014,N_10983);
nor U13740 (N_13740,N_9992,N_11612);
nor U13741 (N_13741,N_10895,N_9317);
or U13742 (N_13742,N_11099,N_11843);
nor U13743 (N_13743,N_11092,N_11136);
and U13744 (N_13744,N_9578,N_9706);
nor U13745 (N_13745,N_9300,N_10453);
and U13746 (N_13746,N_10493,N_10333);
nand U13747 (N_13747,N_11148,N_9448);
and U13748 (N_13748,N_9721,N_11341);
and U13749 (N_13749,N_10095,N_10550);
or U13750 (N_13750,N_10975,N_10141);
nand U13751 (N_13751,N_11805,N_11037);
nand U13752 (N_13752,N_10091,N_11172);
nor U13753 (N_13753,N_11011,N_10935);
or U13754 (N_13754,N_11651,N_10772);
and U13755 (N_13755,N_10665,N_10531);
and U13756 (N_13756,N_10254,N_9496);
and U13757 (N_13757,N_9089,N_11878);
nor U13758 (N_13758,N_10225,N_11278);
or U13759 (N_13759,N_9356,N_9832);
nor U13760 (N_13760,N_11264,N_9449);
nor U13761 (N_13761,N_11811,N_11779);
or U13762 (N_13762,N_11488,N_10087);
and U13763 (N_13763,N_11354,N_10439);
and U13764 (N_13764,N_11570,N_11609);
nor U13765 (N_13765,N_11747,N_10448);
nor U13766 (N_13766,N_10928,N_10572);
nor U13767 (N_13767,N_9864,N_10726);
nand U13768 (N_13768,N_11748,N_9524);
nor U13769 (N_13769,N_11444,N_11424);
nor U13770 (N_13770,N_10798,N_9581);
and U13771 (N_13771,N_10498,N_11736);
and U13772 (N_13772,N_10038,N_9326);
or U13773 (N_13773,N_11313,N_9236);
and U13774 (N_13774,N_10515,N_10671);
and U13775 (N_13775,N_11100,N_9235);
and U13776 (N_13776,N_10596,N_9618);
and U13777 (N_13777,N_10942,N_9402);
or U13778 (N_13778,N_10353,N_9958);
nand U13779 (N_13779,N_11045,N_11320);
nor U13780 (N_13780,N_10052,N_10138);
nand U13781 (N_13781,N_9041,N_11032);
or U13782 (N_13782,N_11088,N_11081);
or U13783 (N_13783,N_9521,N_9483);
nand U13784 (N_13784,N_11879,N_10636);
and U13785 (N_13785,N_10675,N_9141);
nand U13786 (N_13786,N_10842,N_10979);
or U13787 (N_13787,N_9638,N_9307);
and U13788 (N_13788,N_10727,N_9980);
and U13789 (N_13789,N_9737,N_11224);
nor U13790 (N_13790,N_11303,N_9599);
or U13791 (N_13791,N_9753,N_11019);
xor U13792 (N_13792,N_9614,N_11230);
and U13793 (N_13793,N_9387,N_10017);
or U13794 (N_13794,N_9032,N_11254);
or U13795 (N_13795,N_9606,N_11560);
or U13796 (N_13796,N_10325,N_11384);
nor U13797 (N_13797,N_10538,N_9200);
or U13798 (N_13798,N_9008,N_10883);
nor U13799 (N_13799,N_9104,N_10171);
nand U13800 (N_13800,N_11911,N_9892);
nor U13801 (N_13801,N_11914,N_10161);
or U13802 (N_13802,N_10260,N_9004);
or U13803 (N_13803,N_10372,N_10060);
or U13804 (N_13804,N_9292,N_11293);
nor U13805 (N_13805,N_9229,N_11691);
and U13806 (N_13806,N_10658,N_10936);
nand U13807 (N_13807,N_11820,N_11074);
nor U13808 (N_13808,N_11875,N_10794);
nor U13809 (N_13809,N_11313,N_10483);
nand U13810 (N_13810,N_11253,N_10607);
or U13811 (N_13811,N_10918,N_9841);
nor U13812 (N_13812,N_10527,N_11796);
nor U13813 (N_13813,N_9524,N_10403);
or U13814 (N_13814,N_10474,N_9759);
nand U13815 (N_13815,N_10901,N_10022);
nor U13816 (N_13816,N_9100,N_11367);
nor U13817 (N_13817,N_9344,N_10270);
and U13818 (N_13818,N_10106,N_9679);
and U13819 (N_13819,N_11276,N_10850);
nand U13820 (N_13820,N_11863,N_11698);
nor U13821 (N_13821,N_9383,N_11027);
or U13822 (N_13822,N_9627,N_11737);
nor U13823 (N_13823,N_9825,N_11151);
nor U13824 (N_13824,N_10959,N_11419);
or U13825 (N_13825,N_11032,N_10061);
nand U13826 (N_13826,N_11115,N_11055);
nand U13827 (N_13827,N_10495,N_11487);
or U13828 (N_13828,N_9375,N_9269);
or U13829 (N_13829,N_9163,N_11520);
and U13830 (N_13830,N_11155,N_10653);
nor U13831 (N_13831,N_9236,N_9414);
and U13832 (N_13832,N_9299,N_11363);
nand U13833 (N_13833,N_10306,N_11183);
or U13834 (N_13834,N_11695,N_10499);
nor U13835 (N_13835,N_9902,N_9497);
or U13836 (N_13836,N_10506,N_9339);
nor U13837 (N_13837,N_9394,N_9988);
nor U13838 (N_13838,N_9638,N_9979);
nand U13839 (N_13839,N_9300,N_11985);
nor U13840 (N_13840,N_10713,N_11349);
nor U13841 (N_13841,N_10168,N_9032);
nand U13842 (N_13842,N_10080,N_11358);
nor U13843 (N_13843,N_9864,N_11007);
nand U13844 (N_13844,N_10116,N_9562);
nor U13845 (N_13845,N_11821,N_10440);
nand U13846 (N_13846,N_11957,N_11573);
xor U13847 (N_13847,N_10988,N_10133);
nor U13848 (N_13848,N_10249,N_10103);
and U13849 (N_13849,N_10615,N_11735);
nor U13850 (N_13850,N_9652,N_11950);
nand U13851 (N_13851,N_10518,N_10909);
nor U13852 (N_13852,N_9376,N_11180);
or U13853 (N_13853,N_9318,N_9098);
or U13854 (N_13854,N_11407,N_9348);
and U13855 (N_13855,N_9470,N_9610);
nand U13856 (N_13856,N_9793,N_11980);
and U13857 (N_13857,N_9120,N_9118);
nand U13858 (N_13858,N_10790,N_11097);
nand U13859 (N_13859,N_11265,N_11323);
or U13860 (N_13860,N_11323,N_11920);
and U13861 (N_13861,N_11509,N_11817);
or U13862 (N_13862,N_10822,N_11569);
nor U13863 (N_13863,N_11139,N_9303);
nor U13864 (N_13864,N_9313,N_9735);
nand U13865 (N_13865,N_9119,N_9484);
nor U13866 (N_13866,N_9881,N_11461);
or U13867 (N_13867,N_11621,N_11398);
nor U13868 (N_13868,N_10341,N_11670);
and U13869 (N_13869,N_10815,N_9693);
nand U13870 (N_13870,N_9472,N_9693);
nand U13871 (N_13871,N_11818,N_10558);
nor U13872 (N_13872,N_10322,N_11830);
or U13873 (N_13873,N_11373,N_10393);
nor U13874 (N_13874,N_9681,N_11822);
nand U13875 (N_13875,N_10474,N_11967);
nand U13876 (N_13876,N_9106,N_11017);
and U13877 (N_13877,N_9874,N_10407);
nor U13878 (N_13878,N_11532,N_10674);
nand U13879 (N_13879,N_10141,N_10285);
nor U13880 (N_13880,N_10687,N_10217);
and U13881 (N_13881,N_9594,N_9936);
or U13882 (N_13882,N_10311,N_9782);
and U13883 (N_13883,N_11873,N_11408);
or U13884 (N_13884,N_10842,N_11083);
and U13885 (N_13885,N_9276,N_11089);
and U13886 (N_13886,N_11917,N_10638);
nor U13887 (N_13887,N_10406,N_9714);
or U13888 (N_13888,N_9108,N_11056);
nand U13889 (N_13889,N_11664,N_11942);
nand U13890 (N_13890,N_11424,N_11340);
nor U13891 (N_13891,N_11901,N_9464);
nor U13892 (N_13892,N_9897,N_9065);
nor U13893 (N_13893,N_10569,N_10682);
nand U13894 (N_13894,N_9198,N_10451);
nand U13895 (N_13895,N_10620,N_10694);
or U13896 (N_13896,N_10270,N_9350);
nand U13897 (N_13897,N_9849,N_9084);
nor U13898 (N_13898,N_11049,N_10638);
and U13899 (N_13899,N_11464,N_9415);
and U13900 (N_13900,N_10052,N_11231);
nand U13901 (N_13901,N_9304,N_10384);
nor U13902 (N_13902,N_9182,N_11369);
and U13903 (N_13903,N_10525,N_11486);
or U13904 (N_13904,N_11863,N_10901);
and U13905 (N_13905,N_11924,N_9869);
nand U13906 (N_13906,N_9807,N_11630);
nor U13907 (N_13907,N_10655,N_11073);
xor U13908 (N_13908,N_10381,N_11074);
nor U13909 (N_13909,N_10443,N_9759);
nor U13910 (N_13910,N_10673,N_9308);
nand U13911 (N_13911,N_11399,N_11212);
and U13912 (N_13912,N_10511,N_10057);
or U13913 (N_13913,N_11473,N_9333);
xnor U13914 (N_13914,N_11359,N_10325);
nand U13915 (N_13915,N_9459,N_10468);
nor U13916 (N_13916,N_11512,N_10365);
nand U13917 (N_13917,N_11874,N_11721);
nand U13918 (N_13918,N_9323,N_11394);
nor U13919 (N_13919,N_11627,N_11881);
nor U13920 (N_13920,N_9623,N_11435);
nor U13921 (N_13921,N_9932,N_11296);
nand U13922 (N_13922,N_11451,N_9673);
nand U13923 (N_13923,N_9514,N_9999);
nor U13924 (N_13924,N_10026,N_11630);
and U13925 (N_13925,N_10172,N_11310);
and U13926 (N_13926,N_9586,N_11697);
nor U13927 (N_13927,N_10655,N_10754);
nor U13928 (N_13928,N_9290,N_10251);
and U13929 (N_13929,N_9551,N_10541);
nand U13930 (N_13930,N_10535,N_9770);
nand U13931 (N_13931,N_10354,N_11154);
nor U13932 (N_13932,N_10238,N_9269);
and U13933 (N_13933,N_11641,N_10648);
nor U13934 (N_13934,N_11463,N_9335);
and U13935 (N_13935,N_9937,N_9946);
nand U13936 (N_13936,N_9296,N_9624);
nor U13937 (N_13937,N_11804,N_10648);
nand U13938 (N_13938,N_11105,N_9257);
nor U13939 (N_13939,N_9357,N_11413);
nor U13940 (N_13940,N_11610,N_10971);
and U13941 (N_13941,N_11230,N_11728);
or U13942 (N_13942,N_10535,N_11028);
nor U13943 (N_13943,N_9925,N_10820);
or U13944 (N_13944,N_10979,N_11658);
nor U13945 (N_13945,N_11943,N_9414);
or U13946 (N_13946,N_9926,N_9277);
nor U13947 (N_13947,N_9708,N_11622);
or U13948 (N_13948,N_10278,N_11557);
or U13949 (N_13949,N_9556,N_11186);
nor U13950 (N_13950,N_9532,N_9265);
nand U13951 (N_13951,N_9679,N_10202);
or U13952 (N_13952,N_11571,N_10547);
or U13953 (N_13953,N_9155,N_10412);
or U13954 (N_13954,N_9291,N_9405);
and U13955 (N_13955,N_11003,N_11656);
nor U13956 (N_13956,N_10021,N_9937);
nand U13957 (N_13957,N_9641,N_10382);
or U13958 (N_13958,N_11559,N_9114);
nand U13959 (N_13959,N_10376,N_11144);
nor U13960 (N_13960,N_10631,N_9446);
or U13961 (N_13961,N_9644,N_11929);
and U13962 (N_13962,N_10574,N_11048);
and U13963 (N_13963,N_9730,N_10427);
nor U13964 (N_13964,N_11843,N_10136);
nor U13965 (N_13965,N_11676,N_10675);
and U13966 (N_13966,N_11098,N_9291);
nor U13967 (N_13967,N_10262,N_10041);
nand U13968 (N_13968,N_10500,N_11202);
and U13969 (N_13969,N_10763,N_9424);
or U13970 (N_13970,N_9024,N_11746);
nor U13971 (N_13971,N_11070,N_11241);
nand U13972 (N_13972,N_9932,N_9774);
and U13973 (N_13973,N_10400,N_11251);
and U13974 (N_13974,N_9098,N_11125);
nor U13975 (N_13975,N_9028,N_11237);
and U13976 (N_13976,N_9853,N_10472);
or U13977 (N_13977,N_9171,N_9501);
or U13978 (N_13978,N_9564,N_11947);
or U13979 (N_13979,N_11756,N_11023);
or U13980 (N_13980,N_10487,N_10684);
or U13981 (N_13981,N_10582,N_11421);
nand U13982 (N_13982,N_11654,N_11542);
and U13983 (N_13983,N_10612,N_10754);
nor U13984 (N_13984,N_10024,N_9007);
and U13985 (N_13985,N_11574,N_9661);
nor U13986 (N_13986,N_10265,N_11067);
and U13987 (N_13987,N_9707,N_9050);
nor U13988 (N_13988,N_11363,N_9329);
nor U13989 (N_13989,N_9830,N_10685);
or U13990 (N_13990,N_11824,N_9658);
or U13991 (N_13991,N_9409,N_9279);
and U13992 (N_13992,N_10027,N_11418);
and U13993 (N_13993,N_11922,N_10713);
or U13994 (N_13994,N_9168,N_9824);
nor U13995 (N_13995,N_11538,N_9945);
or U13996 (N_13996,N_10395,N_10425);
or U13997 (N_13997,N_9632,N_11724);
nand U13998 (N_13998,N_10101,N_10381);
and U13999 (N_13999,N_10636,N_9672);
or U14000 (N_14000,N_11935,N_10287);
nand U14001 (N_14001,N_9447,N_9349);
xnor U14002 (N_14002,N_9046,N_11516);
nand U14003 (N_14003,N_9850,N_9290);
nor U14004 (N_14004,N_9178,N_9882);
and U14005 (N_14005,N_11713,N_9022);
nand U14006 (N_14006,N_10668,N_9782);
or U14007 (N_14007,N_9318,N_11344);
nor U14008 (N_14008,N_9855,N_9520);
nand U14009 (N_14009,N_10523,N_11817);
nor U14010 (N_14010,N_9486,N_9159);
and U14011 (N_14011,N_11214,N_9042);
nor U14012 (N_14012,N_9590,N_11110);
or U14013 (N_14013,N_11936,N_11481);
nor U14014 (N_14014,N_9414,N_10516);
and U14015 (N_14015,N_10437,N_10775);
nor U14016 (N_14016,N_10236,N_11182);
nor U14017 (N_14017,N_9275,N_11774);
or U14018 (N_14018,N_10189,N_11895);
nor U14019 (N_14019,N_11170,N_11424);
nand U14020 (N_14020,N_10450,N_10439);
and U14021 (N_14021,N_11767,N_10204);
nor U14022 (N_14022,N_10881,N_11342);
or U14023 (N_14023,N_9994,N_11500);
and U14024 (N_14024,N_9762,N_9977);
and U14025 (N_14025,N_11051,N_11749);
or U14026 (N_14026,N_9853,N_10682);
or U14027 (N_14027,N_11229,N_10210);
or U14028 (N_14028,N_11605,N_11279);
and U14029 (N_14029,N_10123,N_9597);
nand U14030 (N_14030,N_11710,N_11317);
and U14031 (N_14031,N_10293,N_9031);
and U14032 (N_14032,N_9029,N_10376);
or U14033 (N_14033,N_11363,N_9189);
and U14034 (N_14034,N_11705,N_10099);
and U14035 (N_14035,N_10667,N_10501);
and U14036 (N_14036,N_10536,N_11729);
or U14037 (N_14037,N_9207,N_11253);
or U14038 (N_14038,N_10106,N_11554);
nor U14039 (N_14039,N_9813,N_9679);
nand U14040 (N_14040,N_9445,N_9630);
nor U14041 (N_14041,N_10832,N_11217);
and U14042 (N_14042,N_9654,N_11735);
or U14043 (N_14043,N_10118,N_11810);
and U14044 (N_14044,N_9221,N_10405);
and U14045 (N_14045,N_11842,N_11836);
and U14046 (N_14046,N_10651,N_11286);
or U14047 (N_14047,N_11706,N_9240);
or U14048 (N_14048,N_11617,N_9555);
and U14049 (N_14049,N_11359,N_9327);
nor U14050 (N_14050,N_11126,N_10975);
and U14051 (N_14051,N_9538,N_9126);
or U14052 (N_14052,N_11626,N_11573);
nand U14053 (N_14053,N_9596,N_9146);
nand U14054 (N_14054,N_10718,N_10851);
or U14055 (N_14055,N_10053,N_10538);
nor U14056 (N_14056,N_11222,N_10963);
or U14057 (N_14057,N_11231,N_10442);
nand U14058 (N_14058,N_9519,N_9548);
nor U14059 (N_14059,N_10835,N_10861);
or U14060 (N_14060,N_9575,N_10273);
nor U14061 (N_14061,N_9305,N_11786);
nor U14062 (N_14062,N_11865,N_11976);
nand U14063 (N_14063,N_9647,N_9056);
nand U14064 (N_14064,N_11387,N_11722);
or U14065 (N_14065,N_9217,N_9482);
and U14066 (N_14066,N_9337,N_11928);
nor U14067 (N_14067,N_10267,N_10434);
or U14068 (N_14068,N_10562,N_11102);
nand U14069 (N_14069,N_9907,N_10922);
or U14070 (N_14070,N_9014,N_10997);
nand U14071 (N_14071,N_11790,N_10648);
and U14072 (N_14072,N_11181,N_11574);
nand U14073 (N_14073,N_11921,N_11872);
nor U14074 (N_14074,N_11319,N_9174);
nor U14075 (N_14075,N_10177,N_11435);
nand U14076 (N_14076,N_9417,N_10529);
or U14077 (N_14077,N_10431,N_9679);
nor U14078 (N_14078,N_11024,N_11796);
or U14079 (N_14079,N_11479,N_10474);
and U14080 (N_14080,N_11199,N_10112);
nand U14081 (N_14081,N_9768,N_10604);
or U14082 (N_14082,N_11527,N_11258);
or U14083 (N_14083,N_10802,N_9017);
nor U14084 (N_14084,N_11273,N_9214);
or U14085 (N_14085,N_9754,N_9127);
nand U14086 (N_14086,N_10373,N_9131);
and U14087 (N_14087,N_11865,N_10327);
and U14088 (N_14088,N_10548,N_10929);
or U14089 (N_14089,N_10916,N_11236);
and U14090 (N_14090,N_9602,N_10136);
nor U14091 (N_14091,N_9386,N_9429);
or U14092 (N_14092,N_9571,N_10814);
and U14093 (N_14093,N_10737,N_11595);
nor U14094 (N_14094,N_9091,N_9301);
or U14095 (N_14095,N_10659,N_10266);
nor U14096 (N_14096,N_11553,N_11060);
nor U14097 (N_14097,N_9961,N_10275);
or U14098 (N_14098,N_9431,N_10609);
and U14099 (N_14099,N_9261,N_10298);
nand U14100 (N_14100,N_10219,N_10164);
nand U14101 (N_14101,N_10561,N_11111);
xor U14102 (N_14102,N_11400,N_11647);
nand U14103 (N_14103,N_10529,N_10485);
and U14104 (N_14104,N_10421,N_10363);
and U14105 (N_14105,N_10807,N_9950);
and U14106 (N_14106,N_10655,N_10411);
and U14107 (N_14107,N_11518,N_11188);
or U14108 (N_14108,N_10376,N_11235);
and U14109 (N_14109,N_11587,N_9468);
or U14110 (N_14110,N_9614,N_10980);
and U14111 (N_14111,N_10526,N_11038);
or U14112 (N_14112,N_11258,N_10874);
nand U14113 (N_14113,N_11535,N_10460);
nor U14114 (N_14114,N_9878,N_10651);
nor U14115 (N_14115,N_11039,N_9366);
nand U14116 (N_14116,N_11470,N_11083);
or U14117 (N_14117,N_11928,N_10108);
or U14118 (N_14118,N_11671,N_9867);
nand U14119 (N_14119,N_11962,N_11784);
or U14120 (N_14120,N_11211,N_10333);
or U14121 (N_14121,N_10624,N_11782);
nor U14122 (N_14122,N_10950,N_10251);
nand U14123 (N_14123,N_9709,N_11555);
or U14124 (N_14124,N_9420,N_11203);
or U14125 (N_14125,N_9462,N_9514);
nand U14126 (N_14126,N_10702,N_10960);
nor U14127 (N_14127,N_9381,N_9307);
and U14128 (N_14128,N_10907,N_9406);
and U14129 (N_14129,N_11445,N_10058);
nand U14130 (N_14130,N_11240,N_10300);
or U14131 (N_14131,N_9441,N_9432);
xnor U14132 (N_14132,N_11697,N_11971);
nor U14133 (N_14133,N_10367,N_11270);
nand U14134 (N_14134,N_9483,N_10474);
and U14135 (N_14135,N_9085,N_10042);
or U14136 (N_14136,N_10981,N_10404);
nor U14137 (N_14137,N_10989,N_9608);
nor U14138 (N_14138,N_10881,N_10760);
nor U14139 (N_14139,N_9203,N_10953);
or U14140 (N_14140,N_9667,N_10307);
nor U14141 (N_14141,N_9772,N_10604);
or U14142 (N_14142,N_10218,N_11188);
nand U14143 (N_14143,N_9662,N_9989);
and U14144 (N_14144,N_11835,N_9676);
nor U14145 (N_14145,N_11966,N_10183);
nand U14146 (N_14146,N_9127,N_10508);
nor U14147 (N_14147,N_10153,N_9874);
and U14148 (N_14148,N_11512,N_10509);
nor U14149 (N_14149,N_9238,N_10794);
or U14150 (N_14150,N_11526,N_10454);
or U14151 (N_14151,N_11701,N_10129);
and U14152 (N_14152,N_9382,N_9618);
nand U14153 (N_14153,N_9868,N_9130);
nor U14154 (N_14154,N_10474,N_11749);
and U14155 (N_14155,N_11308,N_11391);
and U14156 (N_14156,N_11850,N_10737);
and U14157 (N_14157,N_10791,N_11606);
nand U14158 (N_14158,N_11655,N_9054);
or U14159 (N_14159,N_9015,N_9235);
nor U14160 (N_14160,N_11144,N_9902);
or U14161 (N_14161,N_10921,N_9051);
nor U14162 (N_14162,N_11137,N_9699);
and U14163 (N_14163,N_10811,N_9567);
and U14164 (N_14164,N_10078,N_11272);
or U14165 (N_14165,N_11061,N_10033);
and U14166 (N_14166,N_11290,N_9227);
and U14167 (N_14167,N_10988,N_10680);
nand U14168 (N_14168,N_9798,N_11850);
nand U14169 (N_14169,N_9550,N_11370);
nor U14170 (N_14170,N_10126,N_9170);
nand U14171 (N_14171,N_10453,N_9069);
nand U14172 (N_14172,N_10357,N_11318);
nor U14173 (N_14173,N_10476,N_10478);
nor U14174 (N_14174,N_10489,N_11320);
nor U14175 (N_14175,N_10303,N_11223);
nor U14176 (N_14176,N_11316,N_11142);
nand U14177 (N_14177,N_10169,N_9187);
nor U14178 (N_14178,N_11399,N_11711);
nand U14179 (N_14179,N_9458,N_10281);
nor U14180 (N_14180,N_10131,N_10342);
nor U14181 (N_14181,N_11692,N_9541);
nor U14182 (N_14182,N_10049,N_10715);
or U14183 (N_14183,N_11780,N_10259);
nor U14184 (N_14184,N_9909,N_10716);
nor U14185 (N_14185,N_9263,N_10558);
or U14186 (N_14186,N_9630,N_9028);
or U14187 (N_14187,N_11860,N_10587);
nand U14188 (N_14188,N_9062,N_10640);
nor U14189 (N_14189,N_10852,N_10389);
nor U14190 (N_14190,N_11441,N_10020);
nand U14191 (N_14191,N_9344,N_11185);
nor U14192 (N_14192,N_10249,N_10824);
nand U14193 (N_14193,N_11858,N_10048);
and U14194 (N_14194,N_10086,N_9101);
and U14195 (N_14195,N_9561,N_10248);
and U14196 (N_14196,N_10205,N_9979);
nor U14197 (N_14197,N_9968,N_11941);
nor U14198 (N_14198,N_10923,N_10595);
or U14199 (N_14199,N_10188,N_11425);
and U14200 (N_14200,N_10646,N_9737);
nor U14201 (N_14201,N_9158,N_9624);
and U14202 (N_14202,N_10535,N_9564);
or U14203 (N_14203,N_11480,N_10048);
xor U14204 (N_14204,N_9373,N_9199);
nand U14205 (N_14205,N_10694,N_11173);
nand U14206 (N_14206,N_10375,N_11382);
nand U14207 (N_14207,N_9450,N_10509);
nand U14208 (N_14208,N_11483,N_11998);
and U14209 (N_14209,N_11395,N_9357);
or U14210 (N_14210,N_9968,N_11400);
nor U14211 (N_14211,N_9264,N_11141);
or U14212 (N_14212,N_9504,N_9961);
and U14213 (N_14213,N_10191,N_9287);
nor U14214 (N_14214,N_11905,N_9812);
nand U14215 (N_14215,N_11070,N_11377);
or U14216 (N_14216,N_10086,N_9557);
or U14217 (N_14217,N_9867,N_9150);
or U14218 (N_14218,N_9993,N_9456);
and U14219 (N_14219,N_10287,N_10977);
or U14220 (N_14220,N_11256,N_9967);
nor U14221 (N_14221,N_11481,N_10007);
nor U14222 (N_14222,N_11699,N_9794);
nor U14223 (N_14223,N_10513,N_11830);
nor U14224 (N_14224,N_11192,N_10666);
and U14225 (N_14225,N_11227,N_10822);
nand U14226 (N_14226,N_10310,N_11722);
nand U14227 (N_14227,N_10247,N_10402);
nor U14228 (N_14228,N_9368,N_10720);
nor U14229 (N_14229,N_11406,N_10512);
and U14230 (N_14230,N_10104,N_11160);
and U14231 (N_14231,N_11831,N_11265);
xor U14232 (N_14232,N_9799,N_9563);
nor U14233 (N_14233,N_9362,N_10134);
or U14234 (N_14234,N_11484,N_11636);
and U14235 (N_14235,N_10725,N_11870);
nor U14236 (N_14236,N_10196,N_11031);
nand U14237 (N_14237,N_10335,N_10060);
or U14238 (N_14238,N_9087,N_9093);
nor U14239 (N_14239,N_11608,N_9785);
nand U14240 (N_14240,N_11521,N_9181);
nor U14241 (N_14241,N_10470,N_10364);
nand U14242 (N_14242,N_9108,N_11613);
nor U14243 (N_14243,N_11591,N_11963);
or U14244 (N_14244,N_11406,N_11670);
or U14245 (N_14245,N_10470,N_9867);
or U14246 (N_14246,N_10888,N_11311);
nand U14247 (N_14247,N_11288,N_10836);
nand U14248 (N_14248,N_9433,N_10438);
nand U14249 (N_14249,N_10563,N_9627);
nand U14250 (N_14250,N_9214,N_10871);
and U14251 (N_14251,N_10846,N_10057);
and U14252 (N_14252,N_11244,N_10194);
and U14253 (N_14253,N_11964,N_11443);
and U14254 (N_14254,N_9755,N_10467);
nor U14255 (N_14255,N_9966,N_9977);
nor U14256 (N_14256,N_10000,N_9720);
nand U14257 (N_14257,N_10502,N_10938);
or U14258 (N_14258,N_9893,N_10295);
or U14259 (N_14259,N_10976,N_11422);
or U14260 (N_14260,N_11626,N_9910);
and U14261 (N_14261,N_10202,N_10773);
nand U14262 (N_14262,N_9256,N_9654);
and U14263 (N_14263,N_10151,N_11613);
or U14264 (N_14264,N_9623,N_10744);
or U14265 (N_14265,N_11992,N_9063);
or U14266 (N_14266,N_10378,N_11020);
nand U14267 (N_14267,N_10339,N_11869);
or U14268 (N_14268,N_10436,N_9355);
and U14269 (N_14269,N_10797,N_9332);
nor U14270 (N_14270,N_11325,N_11598);
nor U14271 (N_14271,N_11900,N_10659);
nor U14272 (N_14272,N_10073,N_11822);
nand U14273 (N_14273,N_9378,N_9861);
nor U14274 (N_14274,N_9252,N_9775);
nor U14275 (N_14275,N_9926,N_9273);
and U14276 (N_14276,N_11720,N_9269);
nor U14277 (N_14277,N_9815,N_11325);
nor U14278 (N_14278,N_10059,N_11421);
nand U14279 (N_14279,N_9045,N_11240);
nand U14280 (N_14280,N_10953,N_9879);
nor U14281 (N_14281,N_9767,N_10566);
or U14282 (N_14282,N_11405,N_10652);
nor U14283 (N_14283,N_9294,N_9659);
nand U14284 (N_14284,N_11705,N_10357);
or U14285 (N_14285,N_9515,N_11152);
and U14286 (N_14286,N_10983,N_11421);
nor U14287 (N_14287,N_10875,N_9308);
nand U14288 (N_14288,N_9143,N_10642);
nor U14289 (N_14289,N_11534,N_10049);
nand U14290 (N_14290,N_11276,N_10385);
and U14291 (N_14291,N_11424,N_10895);
nand U14292 (N_14292,N_10248,N_9444);
or U14293 (N_14293,N_10424,N_11101);
nor U14294 (N_14294,N_9272,N_10648);
nand U14295 (N_14295,N_11409,N_9377);
and U14296 (N_14296,N_11672,N_9496);
and U14297 (N_14297,N_9491,N_11145);
or U14298 (N_14298,N_10417,N_9381);
nor U14299 (N_14299,N_9627,N_9573);
nor U14300 (N_14300,N_10553,N_9339);
nand U14301 (N_14301,N_10484,N_9775);
nor U14302 (N_14302,N_9381,N_9526);
nor U14303 (N_14303,N_9611,N_10736);
and U14304 (N_14304,N_10697,N_10488);
or U14305 (N_14305,N_10810,N_9045);
nand U14306 (N_14306,N_9585,N_11026);
nand U14307 (N_14307,N_10445,N_9572);
nor U14308 (N_14308,N_10762,N_9890);
and U14309 (N_14309,N_9475,N_11252);
xnor U14310 (N_14310,N_9440,N_10067);
nor U14311 (N_14311,N_10519,N_10134);
nand U14312 (N_14312,N_11477,N_10885);
or U14313 (N_14313,N_9854,N_10585);
nor U14314 (N_14314,N_10207,N_10107);
and U14315 (N_14315,N_9378,N_11131);
and U14316 (N_14316,N_11446,N_11289);
nand U14317 (N_14317,N_9027,N_10243);
nor U14318 (N_14318,N_11475,N_10835);
nand U14319 (N_14319,N_10503,N_11756);
nand U14320 (N_14320,N_10636,N_11413);
nand U14321 (N_14321,N_9121,N_9038);
nand U14322 (N_14322,N_9231,N_9563);
nand U14323 (N_14323,N_9015,N_9890);
xor U14324 (N_14324,N_9641,N_11900);
nand U14325 (N_14325,N_10005,N_10956);
nand U14326 (N_14326,N_11192,N_9959);
and U14327 (N_14327,N_10760,N_9982);
and U14328 (N_14328,N_9891,N_9713);
nand U14329 (N_14329,N_11478,N_10948);
or U14330 (N_14330,N_10972,N_10845);
nand U14331 (N_14331,N_11924,N_10396);
nor U14332 (N_14332,N_9364,N_10802);
and U14333 (N_14333,N_10174,N_10833);
and U14334 (N_14334,N_11675,N_9573);
xor U14335 (N_14335,N_10902,N_11266);
nor U14336 (N_14336,N_9945,N_11397);
or U14337 (N_14337,N_11361,N_11745);
nor U14338 (N_14338,N_9616,N_11983);
nor U14339 (N_14339,N_11125,N_10619);
nand U14340 (N_14340,N_11092,N_11847);
or U14341 (N_14341,N_9345,N_9080);
and U14342 (N_14342,N_10002,N_11821);
nor U14343 (N_14343,N_11430,N_11232);
nand U14344 (N_14344,N_10444,N_9143);
nand U14345 (N_14345,N_11377,N_9967);
nand U14346 (N_14346,N_9410,N_11668);
or U14347 (N_14347,N_9949,N_11984);
nor U14348 (N_14348,N_10179,N_10523);
or U14349 (N_14349,N_10835,N_10648);
and U14350 (N_14350,N_10133,N_10840);
and U14351 (N_14351,N_10792,N_11075);
nand U14352 (N_14352,N_9829,N_9740);
or U14353 (N_14353,N_10806,N_9672);
nand U14354 (N_14354,N_9687,N_11016);
and U14355 (N_14355,N_11835,N_11164);
or U14356 (N_14356,N_9802,N_9282);
and U14357 (N_14357,N_9666,N_10118);
nand U14358 (N_14358,N_11759,N_9401);
nor U14359 (N_14359,N_9537,N_9033);
or U14360 (N_14360,N_9939,N_10214);
and U14361 (N_14361,N_11207,N_11897);
nand U14362 (N_14362,N_9761,N_9588);
nor U14363 (N_14363,N_9851,N_10471);
nand U14364 (N_14364,N_11986,N_9263);
nor U14365 (N_14365,N_10139,N_9290);
nand U14366 (N_14366,N_9006,N_11677);
nor U14367 (N_14367,N_11280,N_9310);
and U14368 (N_14368,N_9953,N_10808);
and U14369 (N_14369,N_9267,N_9589);
nor U14370 (N_14370,N_11285,N_11286);
nor U14371 (N_14371,N_9675,N_11141);
or U14372 (N_14372,N_9864,N_11500);
nand U14373 (N_14373,N_10690,N_9755);
nand U14374 (N_14374,N_11814,N_9661);
nand U14375 (N_14375,N_9089,N_9740);
nand U14376 (N_14376,N_11300,N_11512);
nor U14377 (N_14377,N_10167,N_10131);
and U14378 (N_14378,N_10852,N_10819);
or U14379 (N_14379,N_10847,N_9815);
nand U14380 (N_14380,N_11725,N_9214);
or U14381 (N_14381,N_10094,N_11886);
nor U14382 (N_14382,N_11419,N_11354);
xor U14383 (N_14383,N_11990,N_11456);
nand U14384 (N_14384,N_11772,N_9724);
and U14385 (N_14385,N_11743,N_9970);
and U14386 (N_14386,N_9219,N_10563);
or U14387 (N_14387,N_9300,N_10581);
nand U14388 (N_14388,N_11847,N_10432);
nor U14389 (N_14389,N_10949,N_9144);
or U14390 (N_14390,N_11151,N_11102);
or U14391 (N_14391,N_10867,N_10360);
and U14392 (N_14392,N_10478,N_9658);
nor U14393 (N_14393,N_11704,N_9693);
nor U14394 (N_14394,N_11204,N_11711);
nor U14395 (N_14395,N_9438,N_11611);
nor U14396 (N_14396,N_10632,N_11074);
nor U14397 (N_14397,N_11267,N_9576);
or U14398 (N_14398,N_10178,N_10046);
or U14399 (N_14399,N_9827,N_10514);
nor U14400 (N_14400,N_10407,N_11961);
nand U14401 (N_14401,N_9603,N_11797);
or U14402 (N_14402,N_11172,N_10442);
nor U14403 (N_14403,N_11502,N_10065);
nor U14404 (N_14404,N_9332,N_10450);
xnor U14405 (N_14405,N_10951,N_10253);
or U14406 (N_14406,N_10159,N_11695);
or U14407 (N_14407,N_10123,N_11225);
nor U14408 (N_14408,N_10865,N_11488);
nand U14409 (N_14409,N_9820,N_9520);
or U14410 (N_14410,N_9169,N_11827);
nor U14411 (N_14411,N_9041,N_10727);
nand U14412 (N_14412,N_9253,N_11708);
nand U14413 (N_14413,N_9406,N_10393);
or U14414 (N_14414,N_9113,N_11178);
or U14415 (N_14415,N_10859,N_9967);
nor U14416 (N_14416,N_9792,N_9560);
nor U14417 (N_14417,N_9748,N_11257);
nand U14418 (N_14418,N_10930,N_9927);
or U14419 (N_14419,N_11134,N_10767);
xor U14420 (N_14420,N_11399,N_10216);
nor U14421 (N_14421,N_9839,N_9302);
or U14422 (N_14422,N_11486,N_9577);
nand U14423 (N_14423,N_9770,N_10256);
nand U14424 (N_14424,N_9632,N_9192);
nand U14425 (N_14425,N_9602,N_11185);
or U14426 (N_14426,N_9746,N_11488);
nor U14427 (N_14427,N_9311,N_9046);
nand U14428 (N_14428,N_9538,N_11128);
or U14429 (N_14429,N_9901,N_9142);
nor U14430 (N_14430,N_9136,N_11722);
nand U14431 (N_14431,N_11675,N_11567);
or U14432 (N_14432,N_10251,N_9564);
or U14433 (N_14433,N_9630,N_11635);
nor U14434 (N_14434,N_11582,N_11061);
nor U14435 (N_14435,N_10913,N_11989);
and U14436 (N_14436,N_11027,N_11133);
nor U14437 (N_14437,N_10157,N_10998);
nor U14438 (N_14438,N_9106,N_9228);
nor U14439 (N_14439,N_10648,N_9782);
or U14440 (N_14440,N_9760,N_9198);
nor U14441 (N_14441,N_9108,N_10295);
or U14442 (N_14442,N_11595,N_11525);
nor U14443 (N_14443,N_9195,N_11082);
or U14444 (N_14444,N_11935,N_9049);
or U14445 (N_14445,N_9638,N_11226);
nor U14446 (N_14446,N_9033,N_10713);
and U14447 (N_14447,N_9434,N_10270);
nand U14448 (N_14448,N_9499,N_10437);
nor U14449 (N_14449,N_10381,N_11677);
and U14450 (N_14450,N_11154,N_10959);
or U14451 (N_14451,N_9514,N_10959);
nand U14452 (N_14452,N_11067,N_11829);
or U14453 (N_14453,N_10229,N_11740);
nor U14454 (N_14454,N_9426,N_9006);
nor U14455 (N_14455,N_10555,N_9803);
or U14456 (N_14456,N_11840,N_9612);
nand U14457 (N_14457,N_11919,N_11858);
nand U14458 (N_14458,N_10084,N_11153);
or U14459 (N_14459,N_11439,N_9219);
nor U14460 (N_14460,N_11161,N_9163);
nor U14461 (N_14461,N_10365,N_10399);
or U14462 (N_14462,N_9530,N_11764);
nand U14463 (N_14463,N_9881,N_11579);
nor U14464 (N_14464,N_11339,N_10583);
or U14465 (N_14465,N_9408,N_9626);
nand U14466 (N_14466,N_9687,N_10805);
nor U14467 (N_14467,N_10101,N_11044);
nor U14468 (N_14468,N_11104,N_10682);
or U14469 (N_14469,N_9688,N_10682);
and U14470 (N_14470,N_10892,N_9700);
nand U14471 (N_14471,N_11028,N_10027);
nor U14472 (N_14472,N_10498,N_10281);
nor U14473 (N_14473,N_10643,N_11245);
or U14474 (N_14474,N_9593,N_9525);
nor U14475 (N_14475,N_10528,N_11308);
nor U14476 (N_14476,N_9580,N_10935);
or U14477 (N_14477,N_9953,N_10765);
nor U14478 (N_14478,N_9093,N_9685);
nand U14479 (N_14479,N_10517,N_9930);
nand U14480 (N_14480,N_9561,N_9505);
nor U14481 (N_14481,N_11502,N_9501);
xor U14482 (N_14482,N_11493,N_10070);
nor U14483 (N_14483,N_10901,N_10310);
and U14484 (N_14484,N_10268,N_9661);
and U14485 (N_14485,N_10127,N_10832);
or U14486 (N_14486,N_9693,N_11883);
nand U14487 (N_14487,N_11464,N_9665);
or U14488 (N_14488,N_10727,N_10994);
and U14489 (N_14489,N_11563,N_11992);
nor U14490 (N_14490,N_9273,N_11743);
or U14491 (N_14491,N_9179,N_9208);
nand U14492 (N_14492,N_10015,N_11376);
or U14493 (N_14493,N_9864,N_10195);
or U14494 (N_14494,N_10910,N_10415);
and U14495 (N_14495,N_11111,N_9479);
or U14496 (N_14496,N_10974,N_10325);
or U14497 (N_14497,N_11387,N_9508);
nor U14498 (N_14498,N_10583,N_9021);
nor U14499 (N_14499,N_9597,N_11165);
nand U14500 (N_14500,N_9606,N_11984);
or U14501 (N_14501,N_11068,N_9492);
nand U14502 (N_14502,N_9194,N_11023);
nor U14503 (N_14503,N_10678,N_10444);
or U14504 (N_14504,N_10686,N_11653);
nor U14505 (N_14505,N_10068,N_9890);
or U14506 (N_14506,N_9047,N_9049);
or U14507 (N_14507,N_10471,N_9601);
and U14508 (N_14508,N_10153,N_9859);
or U14509 (N_14509,N_9724,N_9692);
nor U14510 (N_14510,N_10644,N_10522);
or U14511 (N_14511,N_10451,N_9120);
and U14512 (N_14512,N_9575,N_10639);
or U14513 (N_14513,N_9166,N_11750);
and U14514 (N_14514,N_9589,N_9041);
or U14515 (N_14515,N_10368,N_11603);
nor U14516 (N_14516,N_11972,N_10945);
nor U14517 (N_14517,N_9431,N_9311);
or U14518 (N_14518,N_9614,N_11666);
and U14519 (N_14519,N_9503,N_9904);
or U14520 (N_14520,N_11635,N_9274);
nand U14521 (N_14521,N_9143,N_9994);
nand U14522 (N_14522,N_11401,N_10730);
and U14523 (N_14523,N_9230,N_10398);
nor U14524 (N_14524,N_10136,N_9133);
nor U14525 (N_14525,N_11792,N_10575);
nor U14526 (N_14526,N_10241,N_9470);
nand U14527 (N_14527,N_9924,N_10380);
nor U14528 (N_14528,N_11320,N_9479);
nor U14529 (N_14529,N_10198,N_10531);
and U14530 (N_14530,N_10743,N_10217);
or U14531 (N_14531,N_9163,N_11999);
or U14532 (N_14532,N_9001,N_10646);
or U14533 (N_14533,N_11927,N_10459);
nor U14534 (N_14534,N_9568,N_10244);
nand U14535 (N_14535,N_11800,N_11913);
or U14536 (N_14536,N_10808,N_9546);
and U14537 (N_14537,N_9516,N_10660);
or U14538 (N_14538,N_10758,N_11734);
nor U14539 (N_14539,N_9001,N_10747);
nor U14540 (N_14540,N_9663,N_9084);
or U14541 (N_14541,N_10767,N_9713);
or U14542 (N_14542,N_9771,N_11594);
and U14543 (N_14543,N_9951,N_10513);
nor U14544 (N_14544,N_10112,N_10517);
nor U14545 (N_14545,N_9834,N_9074);
nor U14546 (N_14546,N_9814,N_10920);
nor U14547 (N_14547,N_10809,N_11470);
and U14548 (N_14548,N_11997,N_9255);
and U14549 (N_14549,N_9915,N_11422);
and U14550 (N_14550,N_10448,N_10304);
nand U14551 (N_14551,N_9248,N_9962);
and U14552 (N_14552,N_9028,N_11356);
nor U14553 (N_14553,N_11623,N_10482);
nor U14554 (N_14554,N_9419,N_10395);
or U14555 (N_14555,N_11239,N_10192);
nand U14556 (N_14556,N_10816,N_9056);
or U14557 (N_14557,N_11600,N_9016);
and U14558 (N_14558,N_11401,N_10627);
or U14559 (N_14559,N_10861,N_9973);
and U14560 (N_14560,N_9823,N_10616);
nand U14561 (N_14561,N_10247,N_10664);
and U14562 (N_14562,N_10522,N_10253);
or U14563 (N_14563,N_9903,N_11327);
nand U14564 (N_14564,N_11424,N_11625);
nor U14565 (N_14565,N_10936,N_11779);
nor U14566 (N_14566,N_11524,N_10874);
and U14567 (N_14567,N_11504,N_11142);
nand U14568 (N_14568,N_10921,N_10323);
or U14569 (N_14569,N_9219,N_11641);
or U14570 (N_14570,N_11544,N_11732);
nor U14571 (N_14571,N_11199,N_10106);
or U14572 (N_14572,N_11367,N_9411);
or U14573 (N_14573,N_9918,N_10287);
or U14574 (N_14574,N_9695,N_10486);
or U14575 (N_14575,N_11714,N_10297);
nor U14576 (N_14576,N_10884,N_10028);
nand U14577 (N_14577,N_11365,N_10909);
nand U14578 (N_14578,N_11646,N_11343);
or U14579 (N_14579,N_9621,N_9044);
nor U14580 (N_14580,N_11235,N_11030);
or U14581 (N_14581,N_10316,N_10897);
and U14582 (N_14582,N_9378,N_11819);
and U14583 (N_14583,N_9660,N_9250);
nand U14584 (N_14584,N_9323,N_9290);
and U14585 (N_14585,N_11757,N_11435);
nor U14586 (N_14586,N_11139,N_10457);
nand U14587 (N_14587,N_9972,N_11144);
and U14588 (N_14588,N_9314,N_11591);
or U14589 (N_14589,N_11923,N_10799);
and U14590 (N_14590,N_11495,N_9443);
nor U14591 (N_14591,N_10850,N_9139);
nand U14592 (N_14592,N_11588,N_10770);
nor U14593 (N_14593,N_10920,N_9719);
nor U14594 (N_14594,N_9012,N_9075);
nor U14595 (N_14595,N_10824,N_9128);
nand U14596 (N_14596,N_11048,N_10385);
and U14597 (N_14597,N_9707,N_11134);
xnor U14598 (N_14598,N_9222,N_11732);
nand U14599 (N_14599,N_10257,N_11326);
or U14600 (N_14600,N_10805,N_10966);
nor U14601 (N_14601,N_11780,N_9884);
or U14602 (N_14602,N_9101,N_9421);
and U14603 (N_14603,N_10351,N_9880);
or U14604 (N_14604,N_11640,N_10454);
and U14605 (N_14605,N_10250,N_9747);
nor U14606 (N_14606,N_11023,N_10922);
nor U14607 (N_14607,N_9061,N_11253);
or U14608 (N_14608,N_11998,N_11349);
nand U14609 (N_14609,N_10233,N_9592);
nand U14610 (N_14610,N_10369,N_10550);
nor U14611 (N_14611,N_9797,N_10073);
nor U14612 (N_14612,N_9547,N_11154);
nand U14613 (N_14613,N_11010,N_11675);
nor U14614 (N_14614,N_11323,N_11573);
nand U14615 (N_14615,N_11043,N_11150);
or U14616 (N_14616,N_11700,N_9778);
nand U14617 (N_14617,N_10127,N_9099);
nand U14618 (N_14618,N_10824,N_9126);
and U14619 (N_14619,N_11633,N_10280);
and U14620 (N_14620,N_9239,N_11113);
or U14621 (N_14621,N_9420,N_11452);
and U14622 (N_14622,N_11699,N_9650);
or U14623 (N_14623,N_11472,N_9359);
and U14624 (N_14624,N_10124,N_11440);
nor U14625 (N_14625,N_11081,N_11134);
nor U14626 (N_14626,N_11688,N_10873);
nor U14627 (N_14627,N_10574,N_10251);
nand U14628 (N_14628,N_9389,N_11957);
nor U14629 (N_14629,N_11667,N_9461);
and U14630 (N_14630,N_9969,N_11002);
nand U14631 (N_14631,N_10570,N_9076);
nor U14632 (N_14632,N_11790,N_11946);
nand U14633 (N_14633,N_9443,N_11302);
and U14634 (N_14634,N_9020,N_10602);
nand U14635 (N_14635,N_11280,N_10542);
nor U14636 (N_14636,N_10754,N_11235);
or U14637 (N_14637,N_9903,N_9622);
or U14638 (N_14638,N_10387,N_9495);
or U14639 (N_14639,N_9925,N_11193);
nor U14640 (N_14640,N_9027,N_10973);
nor U14641 (N_14641,N_10504,N_11084);
nand U14642 (N_14642,N_11553,N_10865);
or U14643 (N_14643,N_11210,N_9206);
or U14644 (N_14644,N_10805,N_11700);
or U14645 (N_14645,N_9870,N_11817);
nand U14646 (N_14646,N_10859,N_11192);
or U14647 (N_14647,N_10377,N_10467);
and U14648 (N_14648,N_11466,N_10085);
nand U14649 (N_14649,N_11301,N_10102);
and U14650 (N_14650,N_11555,N_11233);
or U14651 (N_14651,N_11457,N_10079);
nor U14652 (N_14652,N_9877,N_10658);
and U14653 (N_14653,N_11041,N_10035);
nor U14654 (N_14654,N_11174,N_10654);
or U14655 (N_14655,N_11623,N_10880);
or U14656 (N_14656,N_10806,N_11944);
nor U14657 (N_14657,N_11973,N_11425);
and U14658 (N_14658,N_9710,N_11664);
nor U14659 (N_14659,N_10654,N_10316);
nand U14660 (N_14660,N_11633,N_11441);
and U14661 (N_14661,N_11494,N_11495);
or U14662 (N_14662,N_9368,N_9797);
nand U14663 (N_14663,N_11033,N_9830);
nand U14664 (N_14664,N_11137,N_10398);
and U14665 (N_14665,N_11751,N_10847);
nand U14666 (N_14666,N_9495,N_10966);
nor U14667 (N_14667,N_10600,N_11900);
or U14668 (N_14668,N_9021,N_10059);
and U14669 (N_14669,N_10732,N_11143);
nor U14670 (N_14670,N_10893,N_10189);
nand U14671 (N_14671,N_9703,N_10875);
nor U14672 (N_14672,N_10796,N_9913);
nor U14673 (N_14673,N_9221,N_11560);
nand U14674 (N_14674,N_9629,N_11165);
nand U14675 (N_14675,N_9878,N_10266);
nor U14676 (N_14676,N_11009,N_11277);
and U14677 (N_14677,N_9354,N_11537);
nor U14678 (N_14678,N_11625,N_9232);
and U14679 (N_14679,N_10465,N_9716);
nor U14680 (N_14680,N_11304,N_10580);
or U14681 (N_14681,N_9355,N_9769);
nand U14682 (N_14682,N_11117,N_10263);
or U14683 (N_14683,N_11660,N_11433);
or U14684 (N_14684,N_9265,N_11733);
or U14685 (N_14685,N_9806,N_11346);
nand U14686 (N_14686,N_9284,N_9235);
or U14687 (N_14687,N_10925,N_9104);
or U14688 (N_14688,N_10780,N_10436);
and U14689 (N_14689,N_10773,N_11497);
and U14690 (N_14690,N_11436,N_11161);
and U14691 (N_14691,N_11769,N_10166);
nand U14692 (N_14692,N_9855,N_9941);
and U14693 (N_14693,N_11006,N_11890);
nand U14694 (N_14694,N_10456,N_10927);
and U14695 (N_14695,N_9375,N_9896);
nand U14696 (N_14696,N_10797,N_9518);
nand U14697 (N_14697,N_9822,N_11442);
nor U14698 (N_14698,N_9037,N_9031);
or U14699 (N_14699,N_9830,N_11422);
nand U14700 (N_14700,N_10751,N_9748);
nor U14701 (N_14701,N_10282,N_11417);
nor U14702 (N_14702,N_9032,N_10508);
nor U14703 (N_14703,N_11050,N_10536);
or U14704 (N_14704,N_10385,N_10527);
or U14705 (N_14705,N_11933,N_11567);
or U14706 (N_14706,N_10894,N_9062);
nand U14707 (N_14707,N_9025,N_11186);
and U14708 (N_14708,N_10410,N_10759);
and U14709 (N_14709,N_9455,N_11058);
nor U14710 (N_14710,N_9837,N_10010);
or U14711 (N_14711,N_11631,N_10814);
nand U14712 (N_14712,N_9091,N_10003);
and U14713 (N_14713,N_9126,N_9733);
nor U14714 (N_14714,N_9436,N_10711);
and U14715 (N_14715,N_11258,N_9370);
nor U14716 (N_14716,N_10462,N_9618);
xnor U14717 (N_14717,N_9062,N_10673);
and U14718 (N_14718,N_9853,N_11101);
nor U14719 (N_14719,N_11932,N_10174);
and U14720 (N_14720,N_10204,N_9139);
and U14721 (N_14721,N_9874,N_10567);
nand U14722 (N_14722,N_10900,N_11805);
nand U14723 (N_14723,N_11412,N_10044);
nor U14724 (N_14724,N_11877,N_9638);
or U14725 (N_14725,N_11706,N_10091);
nand U14726 (N_14726,N_9772,N_10610);
and U14727 (N_14727,N_9237,N_10295);
nand U14728 (N_14728,N_9715,N_10096);
and U14729 (N_14729,N_10293,N_9501);
nand U14730 (N_14730,N_9702,N_11030);
nor U14731 (N_14731,N_9386,N_11866);
xnor U14732 (N_14732,N_11929,N_9796);
and U14733 (N_14733,N_10308,N_11758);
or U14734 (N_14734,N_11322,N_9864);
and U14735 (N_14735,N_11824,N_9168);
and U14736 (N_14736,N_9998,N_9716);
nand U14737 (N_14737,N_11777,N_9219);
or U14738 (N_14738,N_11116,N_10280);
nor U14739 (N_14739,N_11262,N_9024);
or U14740 (N_14740,N_10186,N_9766);
or U14741 (N_14741,N_11829,N_11299);
or U14742 (N_14742,N_9859,N_11998);
nor U14743 (N_14743,N_10968,N_11731);
or U14744 (N_14744,N_11662,N_10685);
and U14745 (N_14745,N_11928,N_10687);
or U14746 (N_14746,N_9468,N_11746);
nand U14747 (N_14747,N_10485,N_11940);
or U14748 (N_14748,N_10534,N_9606);
or U14749 (N_14749,N_11236,N_9603);
nand U14750 (N_14750,N_9332,N_9324);
and U14751 (N_14751,N_10922,N_9921);
nand U14752 (N_14752,N_9124,N_11082);
nor U14753 (N_14753,N_10513,N_11475);
or U14754 (N_14754,N_9721,N_10987);
nor U14755 (N_14755,N_11116,N_10194);
and U14756 (N_14756,N_9579,N_10658);
or U14757 (N_14757,N_9406,N_10655);
nand U14758 (N_14758,N_9799,N_11595);
nor U14759 (N_14759,N_10211,N_10238);
or U14760 (N_14760,N_10833,N_9898);
and U14761 (N_14761,N_9955,N_9743);
and U14762 (N_14762,N_9983,N_9809);
nand U14763 (N_14763,N_10753,N_10868);
nand U14764 (N_14764,N_10417,N_9430);
or U14765 (N_14765,N_11901,N_10048);
and U14766 (N_14766,N_10248,N_9396);
nand U14767 (N_14767,N_11034,N_11905);
nor U14768 (N_14768,N_10201,N_11415);
xor U14769 (N_14769,N_9546,N_9991);
and U14770 (N_14770,N_10375,N_10301);
and U14771 (N_14771,N_9139,N_9229);
and U14772 (N_14772,N_10546,N_10552);
and U14773 (N_14773,N_9773,N_9357);
nor U14774 (N_14774,N_10763,N_9685);
and U14775 (N_14775,N_11815,N_10884);
or U14776 (N_14776,N_10488,N_11688);
and U14777 (N_14777,N_11793,N_10360);
or U14778 (N_14778,N_10498,N_11969);
or U14779 (N_14779,N_9902,N_9106);
nand U14780 (N_14780,N_9936,N_10804);
or U14781 (N_14781,N_11140,N_11119);
or U14782 (N_14782,N_11189,N_11003);
nor U14783 (N_14783,N_10271,N_9573);
nor U14784 (N_14784,N_10416,N_10038);
or U14785 (N_14785,N_9406,N_9384);
nor U14786 (N_14786,N_10767,N_9317);
and U14787 (N_14787,N_9317,N_11643);
or U14788 (N_14788,N_9880,N_9678);
nor U14789 (N_14789,N_10358,N_10301);
or U14790 (N_14790,N_11784,N_11503);
nor U14791 (N_14791,N_10595,N_10256);
or U14792 (N_14792,N_11823,N_11032);
nor U14793 (N_14793,N_9711,N_11878);
nor U14794 (N_14794,N_9903,N_9390);
nand U14795 (N_14795,N_11555,N_9016);
nand U14796 (N_14796,N_11246,N_9288);
and U14797 (N_14797,N_11350,N_9539);
or U14798 (N_14798,N_10142,N_11101);
and U14799 (N_14799,N_10051,N_9653);
nand U14800 (N_14800,N_10704,N_11735);
or U14801 (N_14801,N_10640,N_10668);
nand U14802 (N_14802,N_11312,N_9557);
nor U14803 (N_14803,N_9137,N_10328);
nor U14804 (N_14804,N_10695,N_11081);
and U14805 (N_14805,N_10994,N_11826);
nor U14806 (N_14806,N_9689,N_11402);
or U14807 (N_14807,N_9867,N_10709);
nand U14808 (N_14808,N_10032,N_10623);
nor U14809 (N_14809,N_9041,N_10585);
or U14810 (N_14810,N_11065,N_9077);
and U14811 (N_14811,N_11622,N_10444);
or U14812 (N_14812,N_11194,N_9697);
nor U14813 (N_14813,N_9867,N_11249);
nand U14814 (N_14814,N_10051,N_11155);
and U14815 (N_14815,N_11781,N_9333);
or U14816 (N_14816,N_11522,N_11312);
or U14817 (N_14817,N_11325,N_9189);
or U14818 (N_14818,N_11809,N_11844);
nand U14819 (N_14819,N_10313,N_9909);
or U14820 (N_14820,N_9719,N_11748);
and U14821 (N_14821,N_10340,N_9279);
nor U14822 (N_14822,N_9160,N_10903);
nor U14823 (N_14823,N_11414,N_9710);
or U14824 (N_14824,N_9921,N_9226);
or U14825 (N_14825,N_11406,N_9728);
and U14826 (N_14826,N_9508,N_10809);
nand U14827 (N_14827,N_11317,N_9952);
nor U14828 (N_14828,N_11411,N_11133);
nor U14829 (N_14829,N_11418,N_10756);
or U14830 (N_14830,N_9070,N_10304);
or U14831 (N_14831,N_10097,N_11519);
and U14832 (N_14832,N_10486,N_9030);
nor U14833 (N_14833,N_9931,N_9342);
or U14834 (N_14834,N_10272,N_10069);
nor U14835 (N_14835,N_11065,N_11671);
and U14836 (N_14836,N_10984,N_10528);
and U14837 (N_14837,N_11767,N_9413);
nand U14838 (N_14838,N_10148,N_9828);
and U14839 (N_14839,N_11269,N_10359);
or U14840 (N_14840,N_9160,N_11161);
or U14841 (N_14841,N_11793,N_10661);
and U14842 (N_14842,N_9677,N_10363);
nand U14843 (N_14843,N_10519,N_9755);
and U14844 (N_14844,N_11218,N_10377);
or U14845 (N_14845,N_11086,N_10861);
or U14846 (N_14846,N_9268,N_9607);
nor U14847 (N_14847,N_11115,N_9694);
nand U14848 (N_14848,N_11122,N_9737);
nand U14849 (N_14849,N_11138,N_10717);
or U14850 (N_14850,N_10343,N_10676);
nand U14851 (N_14851,N_9672,N_10177);
or U14852 (N_14852,N_9755,N_9638);
and U14853 (N_14853,N_11229,N_11401);
nor U14854 (N_14854,N_9096,N_11522);
nor U14855 (N_14855,N_9370,N_11115);
or U14856 (N_14856,N_9030,N_10094);
or U14857 (N_14857,N_10423,N_11251);
nand U14858 (N_14858,N_9266,N_10811);
nand U14859 (N_14859,N_11130,N_11648);
nand U14860 (N_14860,N_11632,N_11672);
and U14861 (N_14861,N_9278,N_11437);
and U14862 (N_14862,N_10351,N_10474);
or U14863 (N_14863,N_10467,N_9945);
nand U14864 (N_14864,N_11112,N_11335);
or U14865 (N_14865,N_9543,N_9330);
nand U14866 (N_14866,N_9761,N_10780);
nand U14867 (N_14867,N_10584,N_9317);
nand U14868 (N_14868,N_11099,N_10543);
or U14869 (N_14869,N_9045,N_11723);
nand U14870 (N_14870,N_10478,N_11637);
or U14871 (N_14871,N_10842,N_10050);
nand U14872 (N_14872,N_11155,N_11115);
and U14873 (N_14873,N_11850,N_9034);
or U14874 (N_14874,N_11866,N_11768);
and U14875 (N_14875,N_11676,N_9310);
or U14876 (N_14876,N_10410,N_11598);
nand U14877 (N_14877,N_11675,N_11510);
or U14878 (N_14878,N_10763,N_9080);
nor U14879 (N_14879,N_11205,N_10568);
nor U14880 (N_14880,N_10187,N_10111);
nand U14881 (N_14881,N_11806,N_10343);
and U14882 (N_14882,N_9681,N_11168);
nor U14883 (N_14883,N_11608,N_9378);
nor U14884 (N_14884,N_9223,N_11709);
nand U14885 (N_14885,N_11911,N_11104);
nand U14886 (N_14886,N_11187,N_9636);
nor U14887 (N_14887,N_9833,N_11212);
nand U14888 (N_14888,N_11478,N_9296);
nor U14889 (N_14889,N_11414,N_11551);
or U14890 (N_14890,N_11032,N_11077);
and U14891 (N_14891,N_9052,N_10474);
nand U14892 (N_14892,N_9911,N_11954);
nand U14893 (N_14893,N_11852,N_11153);
nand U14894 (N_14894,N_11090,N_11939);
or U14895 (N_14895,N_9785,N_10301);
and U14896 (N_14896,N_11517,N_9518);
and U14897 (N_14897,N_9710,N_10842);
and U14898 (N_14898,N_9084,N_10803);
nand U14899 (N_14899,N_10773,N_11986);
nand U14900 (N_14900,N_10823,N_9457);
and U14901 (N_14901,N_10482,N_9799);
nor U14902 (N_14902,N_11960,N_11481);
nor U14903 (N_14903,N_9897,N_9872);
nand U14904 (N_14904,N_10957,N_10126);
or U14905 (N_14905,N_9945,N_10255);
nor U14906 (N_14906,N_10487,N_9456);
or U14907 (N_14907,N_11691,N_10825);
nor U14908 (N_14908,N_11613,N_11907);
nor U14909 (N_14909,N_10081,N_10977);
and U14910 (N_14910,N_11371,N_11600);
nor U14911 (N_14911,N_11533,N_11996);
or U14912 (N_14912,N_9552,N_9319);
nor U14913 (N_14913,N_11309,N_10176);
nor U14914 (N_14914,N_9633,N_9049);
or U14915 (N_14915,N_9056,N_9545);
or U14916 (N_14916,N_11145,N_9576);
nor U14917 (N_14917,N_9337,N_9720);
and U14918 (N_14918,N_11913,N_9327);
and U14919 (N_14919,N_9141,N_9226);
nand U14920 (N_14920,N_11087,N_10498);
nor U14921 (N_14921,N_9169,N_11956);
nor U14922 (N_14922,N_9290,N_11056);
and U14923 (N_14923,N_10559,N_10409);
nor U14924 (N_14924,N_10645,N_11532);
and U14925 (N_14925,N_9764,N_11351);
nand U14926 (N_14926,N_10296,N_11929);
and U14927 (N_14927,N_11670,N_11731);
or U14928 (N_14928,N_9247,N_9902);
and U14929 (N_14929,N_10149,N_10849);
nor U14930 (N_14930,N_10662,N_11888);
or U14931 (N_14931,N_11380,N_10336);
and U14932 (N_14932,N_11936,N_10978);
or U14933 (N_14933,N_9328,N_11953);
nand U14934 (N_14934,N_11871,N_9710);
and U14935 (N_14935,N_10283,N_9205);
nor U14936 (N_14936,N_10802,N_10172);
nand U14937 (N_14937,N_11458,N_9568);
nor U14938 (N_14938,N_9825,N_11626);
nand U14939 (N_14939,N_9252,N_11164);
nand U14940 (N_14940,N_9820,N_9937);
nor U14941 (N_14941,N_10668,N_9788);
and U14942 (N_14942,N_10051,N_9721);
or U14943 (N_14943,N_9339,N_10006);
nand U14944 (N_14944,N_11511,N_11683);
nor U14945 (N_14945,N_10221,N_11222);
or U14946 (N_14946,N_10676,N_10484);
nand U14947 (N_14947,N_10080,N_10748);
nor U14948 (N_14948,N_11899,N_11657);
or U14949 (N_14949,N_10935,N_11275);
nand U14950 (N_14950,N_11279,N_9256);
nand U14951 (N_14951,N_10170,N_9128);
nor U14952 (N_14952,N_11866,N_11996);
and U14953 (N_14953,N_10378,N_11725);
and U14954 (N_14954,N_11407,N_10881);
and U14955 (N_14955,N_9913,N_9655);
nor U14956 (N_14956,N_11728,N_10753);
nor U14957 (N_14957,N_10683,N_10577);
nand U14958 (N_14958,N_11585,N_10890);
and U14959 (N_14959,N_11980,N_11685);
nor U14960 (N_14960,N_10832,N_10112);
or U14961 (N_14961,N_9675,N_9950);
or U14962 (N_14962,N_10615,N_10508);
or U14963 (N_14963,N_10043,N_11051);
nand U14964 (N_14964,N_10517,N_11227);
nand U14965 (N_14965,N_10416,N_10396);
and U14966 (N_14966,N_11598,N_9841);
nand U14967 (N_14967,N_11163,N_9160);
and U14968 (N_14968,N_11583,N_10376);
and U14969 (N_14969,N_10885,N_10554);
nand U14970 (N_14970,N_11996,N_9174);
nor U14971 (N_14971,N_11822,N_10906);
nand U14972 (N_14972,N_10875,N_9357);
nor U14973 (N_14973,N_9702,N_10247);
and U14974 (N_14974,N_10678,N_11289);
xor U14975 (N_14975,N_9445,N_9146);
nand U14976 (N_14976,N_11701,N_11822);
nand U14977 (N_14977,N_10502,N_11188);
nand U14978 (N_14978,N_10170,N_10529);
nor U14979 (N_14979,N_9583,N_10215);
nand U14980 (N_14980,N_9201,N_9825);
nor U14981 (N_14981,N_9540,N_11549);
nand U14982 (N_14982,N_10249,N_9992);
nand U14983 (N_14983,N_9724,N_9387);
or U14984 (N_14984,N_10231,N_10837);
and U14985 (N_14985,N_9388,N_9227);
nand U14986 (N_14986,N_11545,N_11910);
nand U14987 (N_14987,N_11880,N_11889);
nor U14988 (N_14988,N_9727,N_10333);
or U14989 (N_14989,N_11632,N_11826);
nor U14990 (N_14990,N_11593,N_9246);
nor U14991 (N_14991,N_9122,N_10225);
nand U14992 (N_14992,N_11546,N_9845);
and U14993 (N_14993,N_11200,N_10385);
nand U14994 (N_14994,N_10328,N_10724);
nor U14995 (N_14995,N_9977,N_11928);
and U14996 (N_14996,N_10531,N_10736);
or U14997 (N_14997,N_9556,N_9202);
nand U14998 (N_14998,N_10292,N_10183);
xor U14999 (N_14999,N_9367,N_9535);
nand UO_0 (O_0,N_14291,N_13043);
nand UO_1 (O_1,N_13186,N_13784);
nor UO_2 (O_2,N_12609,N_14423);
and UO_3 (O_3,N_12183,N_13926);
and UO_4 (O_4,N_13316,N_13975);
nand UO_5 (O_5,N_14607,N_12330);
nor UO_6 (O_6,N_13729,N_13830);
nand UO_7 (O_7,N_12418,N_13852);
nand UO_8 (O_8,N_12594,N_14337);
nand UO_9 (O_9,N_12904,N_14404);
nand UO_10 (O_10,N_13237,N_13315);
nor UO_11 (O_11,N_14642,N_12605);
nand UO_12 (O_12,N_14233,N_12930);
and UO_13 (O_13,N_14018,N_12027);
or UO_14 (O_14,N_12675,N_13628);
or UO_15 (O_15,N_14668,N_12948);
nor UO_16 (O_16,N_14096,N_14646);
nor UO_17 (O_17,N_13670,N_14293);
or UO_18 (O_18,N_12516,N_14990);
or UO_19 (O_19,N_12499,N_13905);
nor UO_20 (O_20,N_14399,N_14497);
or UO_21 (O_21,N_13909,N_12747);
and UO_22 (O_22,N_14521,N_12789);
or UO_23 (O_23,N_14620,N_12051);
or UO_24 (O_24,N_14093,N_14139);
and UO_25 (O_25,N_12462,N_13003);
nand UO_26 (O_26,N_14266,N_14199);
nor UO_27 (O_27,N_14057,N_14530);
nand UO_28 (O_28,N_12742,N_12206);
or UO_29 (O_29,N_14379,N_14185);
nand UO_30 (O_30,N_14572,N_13528);
nand UO_31 (O_31,N_14363,N_14887);
nand UO_32 (O_32,N_13219,N_12372);
xnor UO_33 (O_33,N_13626,N_14056);
nor UO_34 (O_34,N_13236,N_14837);
or UO_35 (O_35,N_14581,N_12097);
or UO_36 (O_36,N_13199,N_13195);
nor UO_37 (O_37,N_12883,N_14566);
or UO_38 (O_38,N_13532,N_13733);
nor UO_39 (O_39,N_14709,N_14638);
and UO_40 (O_40,N_12967,N_13846);
and UO_41 (O_41,N_12293,N_13781);
nor UO_42 (O_42,N_13211,N_12996);
or UO_43 (O_43,N_13115,N_13412);
nor UO_44 (O_44,N_12313,N_14147);
nand UO_45 (O_45,N_12705,N_14600);
nand UO_46 (O_46,N_14737,N_14470);
nor UO_47 (O_47,N_14747,N_13568);
nor UO_48 (O_48,N_14987,N_14697);
and UO_49 (O_49,N_12893,N_12068);
and UO_50 (O_50,N_13821,N_14844);
nor UO_51 (O_51,N_13375,N_14224);
nor UO_52 (O_52,N_12799,N_14691);
nor UO_53 (O_53,N_12038,N_13740);
or UO_54 (O_54,N_14252,N_13664);
and UO_55 (O_55,N_14834,N_13441);
or UO_56 (O_56,N_13997,N_13650);
or UO_57 (O_57,N_14241,N_12739);
and UO_58 (O_58,N_13840,N_13228);
or UO_59 (O_59,N_12238,N_12307);
nand UO_60 (O_60,N_12392,N_12656);
nor UO_61 (O_61,N_12718,N_13659);
and UO_62 (O_62,N_12899,N_14878);
or UO_63 (O_63,N_12055,N_13036);
nand UO_64 (O_64,N_14124,N_12316);
and UO_65 (O_65,N_14755,N_12683);
or UO_66 (O_66,N_13053,N_13411);
nand UO_67 (O_67,N_12821,N_12783);
nor UO_68 (O_68,N_14659,N_12182);
nor UO_69 (O_69,N_13968,N_12442);
and UO_70 (O_70,N_14223,N_12896);
nor UO_71 (O_71,N_12792,N_13941);
nand UO_72 (O_72,N_13871,N_12842);
and UO_73 (O_73,N_14068,N_12597);
or UO_74 (O_74,N_12255,N_13390);
or UO_75 (O_75,N_12518,N_12550);
nor UO_76 (O_76,N_13421,N_12922);
nand UO_77 (O_77,N_14695,N_13566);
and UO_78 (O_78,N_14564,N_14806);
nand UO_79 (O_79,N_12318,N_12651);
or UO_80 (O_80,N_13489,N_12449);
nand UO_81 (O_81,N_12757,N_13482);
or UO_82 (O_82,N_13067,N_13317);
and UO_83 (O_83,N_12288,N_12588);
and UO_84 (O_84,N_13320,N_13266);
and UO_85 (O_85,N_14970,N_12104);
nor UO_86 (O_86,N_14963,N_13303);
and UO_87 (O_87,N_12787,N_13092);
and UO_88 (O_88,N_13560,N_12401);
or UO_89 (O_89,N_12990,N_12088);
nand UO_90 (O_90,N_14140,N_13319);
nor UO_91 (O_91,N_14822,N_13343);
nand UO_92 (O_92,N_12827,N_13354);
nand UO_93 (O_93,N_13527,N_13251);
and UO_94 (O_94,N_12014,N_12947);
nand UO_95 (O_95,N_12579,N_12431);
or UO_96 (O_96,N_12059,N_14354);
and UO_97 (O_97,N_14075,N_13582);
or UO_98 (O_98,N_12774,N_14098);
and UO_99 (O_99,N_13774,N_13042);
and UO_100 (O_100,N_14122,N_12213);
or UO_101 (O_101,N_14089,N_12737);
nor UO_102 (O_102,N_12666,N_14084);
nand UO_103 (O_103,N_12634,N_14651);
or UO_104 (O_104,N_13791,N_13785);
and UO_105 (O_105,N_13338,N_12872);
or UO_106 (O_106,N_13983,N_14571);
nand UO_107 (O_107,N_12423,N_13451);
nand UO_108 (O_108,N_13171,N_13614);
or UO_109 (O_109,N_13282,N_12141);
or UO_110 (O_110,N_13253,N_13299);
nand UO_111 (O_111,N_14920,N_12758);
nand UO_112 (O_112,N_14393,N_12830);
nor UO_113 (O_113,N_12101,N_12025);
nor UO_114 (O_114,N_14242,N_14469);
and UO_115 (O_115,N_12212,N_12080);
nand UO_116 (O_116,N_13134,N_12252);
or UO_117 (O_117,N_12366,N_13698);
nand UO_118 (O_118,N_13807,N_12409);
xnor UO_119 (O_119,N_13818,N_14263);
nor UO_120 (O_120,N_12573,N_14001);
or UO_121 (O_121,N_14891,N_13839);
nand UO_122 (O_122,N_14474,N_13351);
or UO_123 (O_123,N_14429,N_12469);
nor UO_124 (O_124,N_14149,N_13748);
nand UO_125 (O_125,N_12009,N_12087);
or UO_126 (O_126,N_14687,N_13082);
or UO_127 (O_127,N_13561,N_14246);
or UO_128 (O_128,N_13672,N_12982);
or UO_129 (O_129,N_13433,N_12636);
and UO_130 (O_130,N_14849,N_14126);
nor UO_131 (O_131,N_13537,N_13629);
nor UO_132 (O_132,N_13386,N_12233);
or UO_133 (O_133,N_13610,N_12730);
and UO_134 (O_134,N_14013,N_14681);
nor UO_135 (O_135,N_13161,N_12696);
and UO_136 (O_136,N_14117,N_12997);
nor UO_137 (O_137,N_13529,N_14708);
or UO_138 (O_138,N_14678,N_14721);
and UO_139 (O_139,N_13979,N_12297);
or UO_140 (O_140,N_12549,N_14996);
or UO_141 (O_141,N_14824,N_12970);
or UO_142 (O_142,N_13165,N_13724);
nor UO_143 (O_143,N_12750,N_12617);
nor UO_144 (O_144,N_12091,N_12034);
nand UO_145 (O_145,N_12833,N_14957);
or UO_146 (O_146,N_14475,N_13126);
or UO_147 (O_147,N_14658,N_14842);
or UO_148 (O_148,N_14087,N_12711);
nor UO_149 (O_149,N_12196,N_14498);
and UO_150 (O_150,N_14345,N_14739);
nor UO_151 (O_151,N_13802,N_12993);
and UO_152 (O_152,N_14751,N_12593);
nand UO_153 (O_153,N_13458,N_12801);
or UO_154 (O_154,N_12586,N_13328);
nand UO_155 (O_155,N_12358,N_12150);
or UO_156 (O_156,N_13372,N_13661);
or UO_157 (O_157,N_13795,N_13046);
and UO_158 (O_158,N_13246,N_13542);
nand UO_159 (O_159,N_14509,N_13565);
or UO_160 (O_160,N_13240,N_13304);
nand UO_161 (O_161,N_14713,N_12164);
and UO_162 (O_162,N_14921,N_12260);
nor UO_163 (O_163,N_12199,N_13068);
nand UO_164 (O_164,N_13974,N_14900);
nor UO_165 (O_165,N_14437,N_13244);
nor UO_166 (O_166,N_13217,N_13947);
nand UO_167 (O_167,N_14042,N_13706);
nor UO_168 (O_168,N_13008,N_14489);
nor UO_169 (O_169,N_14249,N_13765);
and UO_170 (O_170,N_14361,N_12959);
and UO_171 (O_171,N_13292,N_14298);
nand UO_172 (O_172,N_14176,N_14194);
and UO_173 (O_173,N_12826,N_13462);
nand UO_174 (O_174,N_13914,N_13048);
nand UO_175 (O_175,N_14508,N_14501);
nor UO_176 (O_176,N_13581,N_12795);
nor UO_177 (O_177,N_14245,N_13584);
nor UO_178 (O_178,N_14238,N_12684);
nand UO_179 (O_179,N_12048,N_13612);
or UO_180 (O_180,N_12393,N_13178);
and UO_181 (O_181,N_12067,N_13409);
nor UO_182 (O_182,N_14861,N_13310);
nor UO_183 (O_183,N_13533,N_12314);
and UO_184 (O_184,N_12995,N_13488);
nand UO_185 (O_185,N_13984,N_13596);
nand UO_186 (O_186,N_12460,N_12941);
nand UO_187 (O_187,N_12385,N_12489);
nand UO_188 (O_188,N_13723,N_12224);
nor UO_189 (O_189,N_13295,N_14698);
nor UO_190 (O_190,N_13191,N_12601);
nor UO_191 (O_191,N_14729,N_14253);
nand UO_192 (O_192,N_13583,N_13058);
nand UO_193 (O_193,N_12823,N_12585);
nand UO_194 (O_194,N_14071,N_12357);
nor UO_195 (O_195,N_13604,N_12003);
nor UO_196 (O_196,N_12679,N_13794);
and UO_197 (O_197,N_14874,N_14503);
or UO_198 (O_198,N_13929,N_13097);
and UO_199 (O_199,N_12762,N_14652);
nor UO_200 (O_200,N_13373,N_12610);
nor UO_201 (O_201,N_12669,N_13619);
or UO_202 (O_202,N_12955,N_14738);
or UO_203 (O_203,N_12875,N_12805);
or UO_204 (O_204,N_12292,N_14434);
nand UO_205 (O_205,N_12111,N_13241);
and UO_206 (O_206,N_14209,N_12698);
or UO_207 (O_207,N_14618,N_13452);
and UO_208 (O_208,N_12845,N_13496);
nand UO_209 (O_209,N_14592,N_14511);
or UO_210 (O_210,N_12444,N_12323);
nand UO_211 (O_211,N_12294,N_13197);
and UO_212 (O_212,N_13668,N_12603);
nor UO_213 (O_213,N_14555,N_14030);
nand UO_214 (O_214,N_13049,N_12116);
nor UO_215 (O_215,N_13232,N_13051);
and UO_216 (O_216,N_12640,N_13358);
nor UO_217 (O_217,N_14240,N_14810);
nand UO_218 (O_218,N_12380,N_13579);
nand UO_219 (O_219,N_12804,N_14981);
nor UO_220 (O_220,N_13878,N_12638);
or UO_221 (O_221,N_14567,N_12176);
nor UO_222 (O_222,N_13213,N_12708);
or UO_223 (O_223,N_14527,N_13759);
or UO_224 (O_224,N_12608,N_13311);
nor UO_225 (O_225,N_12022,N_14621);
nand UO_226 (O_226,N_12514,N_12886);
nand UO_227 (O_227,N_13953,N_13880);
nand UO_228 (O_228,N_14959,N_12012);
nand UO_229 (O_229,N_13558,N_14825);
nand UO_230 (O_230,N_12258,N_14364);
and UO_231 (O_231,N_12935,N_12151);
or UO_232 (O_232,N_13167,N_13940);
and UO_233 (O_233,N_14519,N_12250);
nand UO_234 (O_234,N_12342,N_13757);
nand UO_235 (O_235,N_13066,N_14730);
or UO_236 (O_236,N_13907,N_13312);
nand UO_237 (O_237,N_14984,N_13737);
or UO_238 (O_238,N_12533,N_13635);
xnor UO_239 (O_239,N_12735,N_13599);
nand UO_240 (O_240,N_14287,N_14529);
nand UO_241 (O_241,N_12999,N_13927);
or UO_242 (O_242,N_13897,N_14127);
or UO_243 (O_243,N_13032,N_13817);
nor UO_244 (O_244,N_13687,N_14107);
or UO_245 (O_245,N_13615,N_14988);
nand UO_246 (O_246,N_13022,N_14026);
and UO_247 (O_247,N_13270,N_12340);
nand UO_248 (O_248,N_12631,N_12060);
nand UO_249 (O_249,N_13603,N_13469);
nor UO_250 (O_250,N_13720,N_14282);
nand UO_251 (O_251,N_14804,N_12349);
nor UO_252 (O_252,N_14675,N_14673);
nor UO_253 (O_253,N_12869,N_14760);
and UO_254 (O_254,N_12225,N_14095);
nor UO_255 (O_255,N_12822,N_14259);
nand UO_256 (O_256,N_14841,N_13291);
nand UO_257 (O_257,N_13392,N_14630);
xor UO_258 (O_258,N_12596,N_12156);
or UO_259 (O_259,N_12074,N_14701);
and UO_260 (O_260,N_13350,N_12987);
or UO_261 (O_261,N_14785,N_14303);
nand UO_262 (O_262,N_12543,N_14882);
or UO_263 (O_263,N_12979,N_12374);
nor UO_264 (O_264,N_12132,N_13047);
nand UO_265 (O_265,N_13353,N_13778);
nand UO_266 (O_266,N_12071,N_14307);
and UO_267 (O_267,N_12271,N_13401);
or UO_268 (O_268,N_12991,N_14575);
and UO_269 (O_269,N_12818,N_12037);
and UO_270 (O_270,N_12179,N_13288);
nor UO_271 (O_271,N_12910,N_13284);
or UO_272 (O_272,N_14328,N_13007);
nand UO_273 (O_273,N_13344,N_14348);
or UO_274 (O_274,N_14192,N_14174);
nor UO_275 (O_275,N_12298,N_12047);
and UO_276 (O_276,N_14860,N_13478);
or UO_277 (O_277,N_13406,N_12824);
nand UO_278 (O_278,N_12919,N_12720);
nor UO_279 (O_279,N_12016,N_13324);
or UO_280 (O_280,N_12744,N_12944);
nor UO_281 (O_281,N_14934,N_14022);
and UO_282 (O_282,N_13507,N_13297);
or UO_283 (O_283,N_14945,N_14088);
nor UO_284 (O_284,N_13473,N_13223);
and UO_285 (O_285,N_14905,N_12455);
nand UO_286 (O_286,N_13497,N_12646);
and UO_287 (O_287,N_13182,N_14831);
nor UO_288 (O_288,N_13864,N_14868);
and UO_289 (O_289,N_14960,N_12688);
and UO_290 (O_290,N_12337,N_14008);
nand UO_291 (O_291,N_12054,N_13648);
or UO_292 (O_292,N_12246,N_14565);
nand UO_293 (O_293,N_12558,N_13509);
xor UO_294 (O_294,N_13300,N_12254);
or UO_295 (O_295,N_12198,N_14157);
and UO_296 (O_296,N_13959,N_13019);
xnor UO_297 (O_297,N_12650,N_13836);
nor UO_298 (O_298,N_12599,N_12344);
and UO_299 (O_299,N_14230,N_13775);
nand UO_300 (O_300,N_12419,N_14991);
or UO_301 (O_301,N_14388,N_12494);
and UO_302 (O_302,N_12479,N_14256);
nand UO_303 (O_303,N_13040,N_14932);
nand UO_304 (O_304,N_13313,N_14597);
nor UO_305 (O_305,N_14270,N_12839);
nand UO_306 (O_306,N_14405,N_13922);
and UO_307 (O_307,N_14189,N_14829);
nand UO_308 (O_308,N_13826,N_14702);
nor UO_309 (O_309,N_14789,N_13281);
nand UO_310 (O_310,N_13415,N_14438);
and UO_311 (O_311,N_13318,N_14373);
nor UO_312 (O_312,N_12129,N_12001);
nor UO_313 (O_313,N_14232,N_14294);
nor UO_314 (O_314,N_13556,N_14772);
nand UO_315 (O_315,N_14243,N_13783);
nand UO_316 (O_316,N_14525,N_12226);
and UO_317 (O_317,N_13238,N_13541);
nand UO_318 (O_318,N_14975,N_13021);
nand UO_319 (O_319,N_14228,N_12445);
nand UO_320 (O_320,N_14439,N_13719);
nor UO_321 (O_321,N_14599,N_14601);
nor UO_322 (O_322,N_12881,N_14129);
and UO_323 (O_323,N_14025,N_14258);
nor UO_324 (O_324,N_14412,N_12362);
nor UO_325 (O_325,N_13824,N_12786);
and UO_326 (O_326,N_14944,N_14911);
nor UO_327 (O_327,N_14936,N_14915);
and UO_328 (O_328,N_12642,N_12763);
or UO_329 (O_329,N_12951,N_12148);
and UO_330 (O_330,N_12776,N_12185);
and UO_331 (O_331,N_13632,N_14705);
nor UO_332 (O_332,N_13866,N_12147);
or UO_333 (O_333,N_14541,N_14244);
nand UO_334 (O_334,N_14531,N_14451);
nor UO_335 (O_335,N_12474,N_13276);
nor UO_336 (O_336,N_14856,N_14338);
nor UO_337 (O_337,N_13924,N_14455);
xor UO_338 (O_338,N_13133,N_13704);
nor UO_339 (O_339,N_12194,N_12332);
nor UO_340 (O_340,N_14366,N_14289);
nand UO_341 (O_341,N_14622,N_13884);
nor UO_342 (O_342,N_14716,N_13277);
or UO_343 (O_343,N_13339,N_12595);
nor UO_344 (O_344,N_12771,N_14648);
or UO_345 (O_345,N_14769,N_13766);
nand UO_346 (O_346,N_13860,N_12190);
nand UO_347 (O_347,N_14200,N_12808);
nor UO_348 (O_348,N_14778,N_14910);
or UO_349 (O_349,N_13695,N_13993);
nand UO_350 (O_350,N_13002,N_12565);
nor UO_351 (O_351,N_12230,N_12440);
nor UO_352 (O_352,N_12811,N_13814);
or UO_353 (O_353,N_12261,N_12598);
or UO_354 (O_354,N_14329,N_13728);
nand UO_355 (O_355,N_14711,N_14972);
nand UO_356 (O_356,N_14748,N_14576);
nor UO_357 (O_357,N_13459,N_14392);
nand UO_358 (O_358,N_13586,N_12645);
and UO_359 (O_359,N_14735,N_12201);
and UO_360 (O_360,N_13293,N_14496);
and UO_361 (O_361,N_14391,N_14593);
or UO_362 (O_362,N_14781,N_13662);
nor UO_363 (O_363,N_12251,N_14595);
nor UO_364 (O_364,N_13999,N_13378);
or UO_365 (O_365,N_12906,N_12633);
and UO_366 (O_366,N_12365,N_14523);
nand UO_367 (O_367,N_12039,N_12623);
nor UO_368 (O_368,N_14826,N_12784);
and UO_369 (O_369,N_13268,N_14236);
nand UO_370 (O_370,N_12884,N_14649);
or UO_371 (O_371,N_14226,N_12106);
nand UO_372 (O_372,N_12352,N_14492);
nand UO_373 (O_373,N_12653,N_12473);
nand UO_374 (O_374,N_13861,N_12490);
and UO_375 (O_375,N_14173,N_14467);
and UO_376 (O_376,N_12882,N_12963);
and UO_377 (O_377,N_13853,N_13831);
and UO_378 (O_378,N_14250,N_13847);
nand UO_379 (O_379,N_12343,N_12350);
xor UO_380 (O_380,N_13099,N_13259);
nor UO_381 (O_381,N_12501,N_14331);
nand UO_382 (O_382,N_13511,N_12277);
nand UO_383 (O_383,N_13395,N_13083);
and UO_384 (O_384,N_13901,N_14038);
nor UO_385 (O_385,N_14867,N_14623);
nand UO_386 (O_386,N_13660,N_14798);
nand UO_387 (O_387,N_14273,N_12079);
nor UO_388 (O_388,N_13536,N_12351);
or UO_389 (O_389,N_14103,N_14833);
and UO_390 (O_390,N_14546,N_14993);
nor UO_391 (O_391,N_13889,N_12364);
or UO_392 (O_392,N_14815,N_12527);
and UO_393 (O_393,N_14073,N_14894);
or UO_394 (O_394,N_13547,N_12746);
xor UO_395 (O_395,N_13617,N_12211);
and UO_396 (O_396,N_14502,N_12897);
nor UO_397 (O_397,N_14692,N_14375);
nor UO_398 (O_398,N_12706,N_12866);
nand UO_399 (O_399,N_14603,N_12940);
nor UO_400 (O_400,N_14097,N_13689);
nor UO_401 (O_401,N_13075,N_14888);
nor UO_402 (O_402,N_14105,N_13873);
or UO_403 (O_403,N_12764,N_13333);
nand UO_404 (O_404,N_12145,N_13813);
or UO_405 (O_405,N_13913,N_13346);
nand UO_406 (O_406,N_13652,N_14752);
and UO_407 (O_407,N_12552,N_12123);
nor UO_408 (O_408,N_13883,N_14195);
nor UO_409 (O_409,N_12689,N_12761);
nand UO_410 (O_410,N_12387,N_12045);
nand UO_411 (O_411,N_13389,N_14432);
nand UO_412 (O_412,N_12992,N_13340);
or UO_413 (O_413,N_13772,N_13621);
nor UO_414 (O_414,N_12551,N_12876);
nand UO_415 (O_415,N_12028,N_14415);
nor UO_416 (O_416,N_14536,N_13329);
or UO_417 (O_417,N_14578,N_12269);
and UO_418 (O_418,N_13519,N_13812);
nor UO_419 (O_419,N_13911,N_13858);
and UO_420 (O_420,N_14543,N_14854);
and UO_421 (O_421,N_13750,N_14418);
nand UO_422 (O_422,N_13693,N_13206);
or UO_423 (O_423,N_13247,N_13214);
or UO_424 (O_424,N_13606,N_14344);
nor UO_425 (O_425,N_13535,N_12015);
nor UO_426 (O_426,N_14980,N_12933);
or UO_427 (O_427,N_12478,N_14665);
and UO_428 (O_428,N_13990,N_12870);
or UO_429 (O_429,N_14956,N_14931);
or UO_430 (O_430,N_14614,N_14974);
nor UO_431 (O_431,N_13111,N_13801);
or UO_432 (O_432,N_12895,N_14004);
and UO_433 (O_433,N_13675,N_12484);
or UO_434 (O_434,N_14385,N_14398);
nor UO_435 (O_435,N_13903,N_13827);
nand UO_436 (O_436,N_14694,N_12539);
nor UO_437 (O_437,N_14362,N_12495);
nor UO_438 (O_438,N_13559,N_13444);
or UO_439 (O_439,N_13498,N_14167);
nand UO_440 (O_440,N_14821,N_13327);
nor UO_441 (O_441,N_12138,N_14720);
or UO_442 (O_442,N_12265,N_14091);
and UO_443 (O_443,N_14717,N_12917);
or UO_444 (O_444,N_12980,N_13256);
or UO_445 (O_445,N_13424,N_14351);
or UO_446 (O_446,N_12532,N_13505);
and UO_447 (O_447,N_12788,N_13280);
and UO_448 (O_448,N_12729,N_12195);
nor UO_449 (O_449,N_14895,N_14274);
nand UO_450 (O_450,N_13054,N_14955);
nand UO_451 (O_451,N_12981,N_14285);
nand UO_452 (O_452,N_13138,N_12432);
or UO_453 (O_453,N_13856,N_12434);
nor UO_454 (O_454,N_12453,N_12278);
and UO_455 (O_455,N_12538,N_13707);
nand UO_456 (O_456,N_14201,N_13263);
or UO_457 (O_457,N_13257,N_12812);
nor UO_458 (O_458,N_14283,N_13136);
nand UO_459 (O_459,N_13001,N_14413);
and UO_460 (O_460,N_13520,N_14181);
or UO_461 (O_461,N_12984,N_14484);
nor UO_462 (O_462,N_12457,N_14872);
or UO_463 (O_463,N_14594,N_12791);
nand UO_464 (O_464,N_12960,N_13077);
nand UO_465 (O_465,N_14703,N_13789);
and UO_466 (O_466,N_13419,N_13116);
and UO_467 (O_467,N_12107,N_14645);
nand UO_468 (O_468,N_12328,N_12128);
or UO_469 (O_469,N_12751,N_14280);
nor UO_470 (O_470,N_12333,N_13718);
and UO_471 (O_471,N_12630,N_14464);
nor UO_472 (O_472,N_13934,N_12639);
or UO_473 (O_473,N_13466,N_14141);
xor UO_474 (O_474,N_12856,N_13899);
nand UO_475 (O_475,N_12607,N_12486);
and UO_476 (O_476,N_12506,N_12019);
and UO_477 (O_477,N_12621,N_14357);
and UO_478 (O_478,N_14033,N_12384);
and UO_479 (O_479,N_12282,N_14335);
or UO_480 (O_480,N_13657,N_14014);
or UO_481 (O_481,N_14902,N_13551);
nor UO_482 (O_482,N_12065,N_13651);
or UO_483 (O_483,N_13222,N_12086);
and UO_484 (O_484,N_13027,N_14965);
nand UO_485 (O_485,N_13731,N_12591);
nand UO_486 (O_486,N_13502,N_14465);
nor UO_487 (O_487,N_14884,N_12503);
or UO_488 (O_488,N_14780,N_13755);
or UO_489 (O_489,N_12069,N_12697);
nor UO_490 (O_490,N_14390,N_14537);
nor UO_491 (O_491,N_14397,N_13763);
and UO_492 (O_492,N_14402,N_13637);
nor UO_493 (O_493,N_13751,N_13404);
nor UO_494 (O_494,N_13286,N_14770);
or UO_495 (O_495,N_14473,N_14689);
or UO_496 (O_496,N_14165,N_14319);
nor UO_497 (O_497,N_14669,N_12912);
nand UO_498 (O_498,N_13376,N_13101);
nand UO_499 (O_499,N_12908,N_14846);
or UO_500 (O_500,N_14542,N_13538);
and UO_501 (O_501,N_12388,N_14381);
nand UO_502 (O_502,N_13643,N_14545);
nand UO_503 (O_503,N_13923,N_13302);
and UO_504 (O_504,N_14143,N_12662);
nor UO_505 (O_505,N_12006,N_13309);
and UO_506 (O_506,N_13210,N_12043);
nor UO_507 (O_507,N_13198,N_14039);
or UO_508 (O_508,N_14672,N_12546);
or UO_509 (O_509,N_13932,N_14172);
nor UO_510 (O_510,N_14290,N_14229);
and UO_511 (O_511,N_13620,N_13904);
and UO_512 (O_512,N_14933,N_14156);
or UO_513 (O_513,N_12174,N_12722);
or UO_514 (O_514,N_13655,N_13301);
xnor UO_515 (O_515,N_13521,N_12512);
or UO_516 (O_516,N_13699,N_14995);
or UO_517 (O_517,N_13164,N_12461);
nor UO_518 (O_518,N_13103,N_12341);
or UO_519 (O_519,N_14724,N_13855);
and UO_520 (O_520,N_12447,N_12652);
nor UO_521 (O_521,N_14719,N_13936);
or UO_522 (O_522,N_12077,N_12188);
nor UO_523 (O_523,N_14763,N_14297);
xnor UO_524 (O_524,N_12248,N_12215);
nand UO_525 (O_525,N_14491,N_13017);
or UO_526 (O_526,N_14162,N_13330);
nor UO_527 (O_527,N_14355,N_12618);
and UO_528 (O_528,N_13796,N_12778);
nand UO_529 (O_529,N_12200,N_13605);
or UO_530 (O_530,N_12485,N_12862);
and UO_531 (O_531,N_13271,N_13961);
or UO_532 (O_532,N_14512,N_14548);
nand UO_533 (O_533,N_12702,N_14712);
and UO_534 (O_534,N_12438,N_14268);
nor UO_535 (O_535,N_12070,N_12810);
and UO_536 (O_536,N_14637,N_14485);
nand UO_537 (O_537,N_14740,N_13758);
nor UO_538 (O_538,N_13290,N_12901);
and UO_539 (O_539,N_13227,N_14370);
and UO_540 (O_540,N_13102,N_14389);
and UO_541 (O_541,N_13705,N_14938);
and UO_542 (O_542,N_13769,N_13684);
or UO_543 (O_543,N_12042,N_12399);
nor UO_544 (O_544,N_13091,N_14903);
and UO_545 (O_545,N_12670,N_13512);
or UO_546 (O_546,N_13753,N_13726);
and UO_547 (O_547,N_12853,N_14560);
and UO_548 (O_548,N_14916,N_12865);
nand UO_549 (O_549,N_13475,N_14327);
nand UO_550 (O_550,N_14146,N_12172);
nor UO_551 (O_551,N_14985,N_13806);
nor UO_552 (O_552,N_12429,N_12394);
or UO_553 (O_553,N_12407,N_12681);
nor UO_554 (O_554,N_14066,N_13188);
or UO_555 (O_555,N_12050,N_13712);
or UO_556 (O_556,N_13996,N_13965);
nand UO_557 (O_557,N_14119,N_14914);
or UO_558 (O_558,N_12975,N_14336);
and UO_559 (O_559,N_12322,N_12846);
and UO_560 (O_560,N_12961,N_14326);
nor UO_561 (O_561,N_12504,N_14550);
nand UO_562 (O_562,N_14617,N_13157);
or UO_563 (O_563,N_14520,N_14788);
xnor UO_564 (O_564,N_12584,N_12428);
nand UO_565 (O_565,N_14365,N_13006);
nor UO_566 (O_566,N_12189,N_12241);
nor UO_567 (O_567,N_14160,N_14288);
nand UO_568 (O_568,N_12436,N_13886);
and UO_569 (O_569,N_13166,N_14812);
and UO_570 (O_570,N_13308,N_14264);
nand UO_571 (O_571,N_14941,N_13641);
nor UO_572 (O_572,N_13449,N_13744);
nor UO_573 (O_573,N_14483,N_12085);
nor UO_574 (O_574,N_12184,N_14396);
nand UO_575 (O_575,N_12770,N_14532);
or UO_576 (O_576,N_14976,N_14655);
or UO_577 (O_577,N_14472,N_13084);
nand UO_578 (O_578,N_13638,N_13669);
nor UO_579 (O_579,N_13235,N_14002);
xnor UO_580 (O_580,N_12105,N_13437);
and UO_581 (O_581,N_12998,N_12140);
or UO_582 (O_582,N_14518,N_14374);
and UO_583 (O_583,N_13964,N_12040);
nor UO_584 (O_584,N_13803,N_12965);
or UO_585 (O_585,N_14376,N_13180);
nor UO_586 (O_586,N_14947,N_13665);
and UO_587 (O_587,N_14634,N_12094);
nand UO_588 (O_588,N_12687,N_12379);
xor UO_589 (O_589,N_13939,N_14794);
or UO_590 (O_590,N_13747,N_13967);
nand UO_591 (O_591,N_14481,N_12157);
or UO_592 (O_592,N_13642,N_14445);
and UO_593 (O_593,N_14009,N_14609);
nand UO_594 (O_594,N_12554,N_13109);
nand UO_595 (O_595,N_13591,N_12170);
and UO_596 (O_596,N_14145,N_13039);
and UO_597 (O_597,N_14494,N_14431);
nor UO_598 (O_598,N_12658,N_12168);
nand UO_599 (O_599,N_12719,N_12918);
nor UO_600 (O_600,N_14216,N_13100);
or UO_601 (O_601,N_14734,N_12715);
nor UO_602 (O_602,N_13374,N_12044);
and UO_603 (O_603,N_14078,N_14113);
nand UO_604 (O_604,N_12663,N_14086);
or UO_605 (O_605,N_14862,N_14704);
nand UO_606 (O_606,N_12117,N_12120);
nor UO_607 (O_607,N_12854,N_12075);
nand UO_608 (O_608,N_14925,N_12325);
and UO_609 (O_609,N_14631,N_14011);
nand UO_610 (O_610,N_14857,N_12767);
or UO_611 (O_611,N_13095,N_12813);
nand UO_612 (O_612,N_14880,N_14969);
nand UO_613 (O_613,N_14128,N_14851);
xor UO_614 (O_614,N_13954,N_13548);
and UO_615 (O_615,N_14881,N_12682);
and UO_616 (O_616,N_12754,N_12338);
nor UO_617 (O_617,N_12216,N_12809);
or UO_618 (O_618,N_14171,N_14644);
and UO_619 (O_619,N_13985,N_12738);
nand UO_620 (O_620,N_14382,N_14024);
and UO_621 (O_621,N_13207,N_12165);
nand UO_622 (O_622,N_12131,N_12637);
nor UO_623 (O_623,N_13773,N_13052);
or UO_624 (O_624,N_13543,N_12417);
and UO_625 (O_625,N_13274,N_14504);
and UO_626 (O_626,N_14021,N_13143);
or UO_627 (O_627,N_12446,N_13436);
or UO_628 (O_628,N_13177,N_14114);
or UO_629 (O_629,N_12249,N_13739);
nor UO_630 (O_630,N_14424,N_12815);
and UO_631 (O_631,N_14308,N_12759);
nor UO_632 (O_632,N_14696,N_14436);
or UO_633 (O_633,N_14387,N_13486);
nor UO_634 (O_634,N_14892,N_12525);
nand UO_635 (O_635,N_13667,N_14378);
nand UO_636 (O_636,N_13239,N_13920);
nor UO_637 (O_637,N_12056,N_13978);
nand UO_638 (O_638,N_14453,N_13129);
and UO_639 (O_639,N_13141,N_12741);
or UO_640 (O_640,N_12266,N_14380);
and UO_641 (O_641,N_13782,N_14507);
and UO_642 (O_642,N_14653,N_13196);
nand UO_643 (O_643,N_13673,N_13948);
nor UO_644 (O_644,N_13434,N_13185);
nor UO_645 (O_645,N_13044,N_12871);
nand UO_646 (O_646,N_14526,N_13423);
or UO_647 (O_647,N_14049,N_14707);
nand UO_648 (O_648,N_12716,N_12841);
nor UO_649 (O_649,N_14108,N_12320);
or UO_650 (O_650,N_13624,N_14219);
or UO_651 (O_651,N_13992,N_14725);
nand UO_652 (O_652,N_14099,N_14315);
nor UO_653 (O_653,N_14569,N_13666);
and UO_654 (O_654,N_12740,N_12286);
nor UO_655 (O_655,N_12890,N_12018);
or UO_656 (O_656,N_14299,N_14175);
and UO_657 (O_657,N_12611,N_14795);
or UO_658 (O_658,N_14346,N_13094);
nand UO_659 (O_659,N_13476,N_12709);
nor UO_660 (O_660,N_14449,N_13159);
and UO_661 (O_661,N_12613,N_12122);
or UO_662 (O_662,N_13862,N_12529);
nand UO_663 (O_663,N_12030,N_12777);
nor UO_664 (O_664,N_14403,N_14510);
or UO_665 (O_665,N_12988,N_14460);
nand UO_666 (O_666,N_12644,N_14235);
and UO_667 (O_667,N_13676,N_12564);
or UO_668 (O_668,N_12578,N_14870);
nor UO_669 (O_669,N_14773,N_12699);
or UO_670 (O_670,N_13004,N_13369);
and UO_671 (O_671,N_12210,N_14919);
and UO_672 (O_672,N_14598,N_13962);
nand UO_673 (O_673,N_14163,N_13587);
nand UO_674 (O_674,N_12589,N_14488);
nor UO_675 (O_675,N_12580,N_12142);
nor UO_676 (O_676,N_14211,N_13949);
or UO_677 (O_677,N_12280,N_14768);
and UO_678 (O_678,N_12727,N_12467);
and UO_679 (O_679,N_14203,N_14746);
and UO_680 (O_680,N_13825,N_13589);
or UO_681 (O_681,N_12377,N_14476);
nand UO_682 (O_682,N_13531,N_12002);
nor UO_683 (O_683,N_12615,N_12221);
and UO_684 (O_684,N_12240,N_14456);
nand UO_685 (O_685,N_12456,N_13105);
nand UO_686 (O_686,N_12517,N_12084);
or UO_687 (O_687,N_12262,N_13254);
or UO_688 (O_688,N_12451,N_13245);
or UO_689 (O_689,N_13041,N_14908);
nand UO_690 (O_690,N_12559,N_14120);
or UO_691 (O_691,N_13492,N_14836);
nand UO_692 (O_692,N_14367,N_14222);
xor UO_693 (O_693,N_13011,N_14558);
nand UO_694 (O_694,N_13446,N_12302);
nor UO_695 (O_695,N_13816,N_14893);
nor UO_696 (O_696,N_12962,N_12507);
nand UO_697 (O_697,N_12903,N_14349);
nand UO_698 (O_698,N_13050,N_14577);
nand UO_699 (O_699,N_12555,N_14670);
nor UO_700 (O_700,N_14757,N_13916);
nand UO_701 (O_701,N_13690,N_14845);
or UO_702 (O_702,N_12424,N_12569);
and UO_703 (O_703,N_13215,N_14817);
nor UO_704 (O_704,N_14419,N_13854);
nand UO_705 (O_705,N_13152,N_12731);
or UO_706 (O_706,N_13460,N_12062);
and UO_707 (O_707,N_13574,N_13357);
nand UO_708 (O_708,N_14863,N_14359);
and UO_709 (O_709,N_14462,N_12725);
nor UO_710 (O_710,N_14736,N_12234);
nor UO_711 (O_711,N_13877,N_12259);
and UO_712 (O_712,N_12861,N_13155);
and UO_713 (O_713,N_12649,N_13870);
and UO_714 (O_714,N_12500,N_12847);
nor UO_715 (O_715,N_13627,N_14205);
nor UO_716 (O_716,N_13345,N_14448);
or UO_717 (O_717,N_12655,N_12969);
nor UO_718 (O_718,N_14440,N_12972);
or UO_719 (O_719,N_12287,N_14796);
nand UO_720 (O_720,N_14685,N_12781);
nor UO_721 (O_721,N_14950,N_12152);
and UO_722 (O_722,N_13224,N_14753);
or UO_723 (O_723,N_12547,N_12437);
nor UO_724 (O_724,N_13279,N_14131);
nand UO_725 (O_725,N_12817,N_13117);
xnor UO_726 (O_726,N_13893,N_13364);
or UO_727 (O_727,N_12193,N_14077);
or UO_728 (O_728,N_12521,N_13994);
and UO_729 (O_729,N_14411,N_13685);
nand UO_730 (O_730,N_12680,N_12118);
nand UO_731 (O_731,N_12700,N_13427);
or UO_732 (O_732,N_14761,N_14262);
nand UO_733 (O_733,N_12868,N_14277);
and UO_734 (O_734,N_13777,N_13562);
nor UO_735 (O_735,N_14304,N_12335);
or UO_736 (O_736,N_14662,N_14486);
or UO_737 (O_737,N_12950,N_14050);
nand UO_738 (O_738,N_14316,N_12239);
or UO_739 (O_739,N_13012,N_13593);
or UO_740 (O_740,N_13780,N_12939);
nand UO_741 (O_741,N_14109,N_12492);
or UO_742 (O_742,N_13991,N_13760);
and UO_743 (O_743,N_13578,N_13336);
or UO_744 (O_744,N_12391,N_13952);
or UO_745 (O_745,N_12304,N_13575);
nand UO_746 (O_746,N_14613,N_14776);
nand UO_747 (O_747,N_14158,N_12619);
nor UO_748 (O_748,N_12674,N_12158);
or UO_749 (O_749,N_14556,N_13514);
nor UO_750 (O_750,N_14534,N_13534);
or UO_751 (O_751,N_14153,N_14994);
or UO_752 (O_752,N_14272,N_13859);
and UO_753 (O_753,N_12756,N_13225);
nor UO_754 (O_754,N_14198,N_12511);
and UO_755 (O_755,N_14540,N_13074);
nor UO_756 (O_756,N_12296,N_12907);
nor UO_757 (O_757,N_13325,N_14535);
and UO_758 (O_758,N_14633,N_13874);
nand UO_759 (O_759,N_12202,N_14466);
nor UO_760 (O_760,N_12124,N_13554);
nor UO_761 (O_761,N_12284,N_14356);
and UO_762 (O_762,N_12072,N_13031);
nand UO_763 (O_763,N_14027,N_13062);
or UO_764 (O_764,N_12488,N_14046);
or UO_765 (O_765,N_13298,N_14859);
nand UO_766 (O_766,N_13352,N_12782);
and UO_767 (O_767,N_12408,N_14275);
and UO_768 (O_768,N_13849,N_12496);
nor UO_769 (O_769,N_14311,N_14977);
or UO_770 (O_770,N_14783,N_12100);
or UO_771 (O_771,N_13289,N_12435);
nor UO_772 (O_772,N_13108,N_14801);
nor UO_773 (O_773,N_12191,N_14048);
and UO_774 (O_774,N_14883,N_12885);
nand UO_775 (O_775,N_14321,N_13815);
nor UO_776 (O_776,N_13037,N_13416);
nand UO_777 (O_777,N_13089,N_13956);
nand UO_778 (O_778,N_12834,N_13153);
and UO_779 (O_779,N_12994,N_13644);
and UO_780 (O_780,N_14479,N_12929);
and UO_781 (O_781,N_14010,N_12838);
or UO_782 (O_782,N_14023,N_12548);
or UO_783 (O_783,N_12368,N_14168);
and UO_784 (O_784,N_12976,N_13697);
or UO_785 (O_785,N_13071,N_12576);
and UO_786 (O_786,N_13065,N_13518);
or UO_787 (O_787,N_12796,N_13016);
nand UO_788 (O_788,N_12814,N_14745);
and UO_789 (O_789,N_14208,N_13283);
or UO_790 (O_790,N_12181,N_14410);
nor UO_791 (O_791,N_13443,N_13220);
and UO_792 (O_792,N_12966,N_12160);
nand UO_793 (O_793,N_12732,N_13957);
or UO_794 (O_794,N_12923,N_12482);
nor UO_795 (O_795,N_12932,N_12163);
nor UO_796 (O_796,N_13829,N_14939);
and UO_797 (O_797,N_12583,N_12888);
or UO_798 (O_798,N_13176,N_13762);
nor UO_799 (O_799,N_12849,N_12857);
nand UO_800 (O_800,N_14639,N_14879);
nand UO_801 (O_801,N_12095,N_12369);
or UO_802 (O_802,N_13808,N_12289);
or UO_803 (O_803,N_14586,N_14251);
and UO_804 (O_804,N_14179,N_13761);
nand UO_805 (O_805,N_12441,N_12542);
and UO_806 (O_806,N_12471,N_14610);
nand UO_807 (O_807,N_13725,N_13341);
and UO_808 (O_808,N_12053,N_12513);
or UO_809 (O_809,N_12820,N_12528);
nor UO_810 (O_810,N_14583,N_12458);
nor UO_811 (O_811,N_14762,N_12276);
and UO_812 (O_812,N_12285,N_12530);
or UO_813 (O_813,N_14314,N_13921);
and UO_814 (O_814,N_14573,N_14408);
nor UO_815 (O_815,N_13976,N_14400);
or UO_816 (O_816,N_13170,N_13025);
and UO_817 (O_817,N_14930,N_12892);
nor UO_818 (O_818,N_13151,N_12665);
and UO_819 (O_819,N_12667,N_12673);
or UO_820 (O_820,N_12121,N_14953);
nand UO_821 (O_821,N_13033,N_14420);
or UO_822 (O_822,N_13879,N_13499);
and UO_823 (O_823,N_14615,N_13145);
and UO_824 (O_824,N_14342,N_13491);
nor UO_825 (O_825,N_12021,N_14818);
xnor UO_826 (O_826,N_14929,N_12167);
or UO_827 (O_827,N_12779,N_13680);
nand UO_828 (O_828,N_14196,N_14898);
nand UO_829 (O_829,N_12078,N_14343);
and UO_830 (O_830,N_14587,N_13630);
and UO_831 (O_831,N_13118,N_14588);
and UO_832 (O_832,N_14371,N_12879);
or UO_833 (O_833,N_13070,N_14395);
and UO_834 (O_834,N_14718,N_14043);
nor UO_835 (O_835,N_12398,N_13229);
nand UO_836 (O_836,N_13918,N_13634);
and UO_837 (O_837,N_14051,N_13209);
nand UO_838 (O_838,N_14480,N_14722);
or UO_839 (O_839,N_13233,N_13367);
nor UO_840 (O_840,N_12481,N_14055);
nand UO_841 (O_841,N_14619,N_12171);
or UO_842 (O_842,N_13377,N_12553);
or UO_843 (O_843,N_13881,N_14549);
and UO_844 (O_844,N_13487,N_12524);
nor UO_845 (O_845,N_12242,N_13592);
nor UO_846 (O_846,N_14997,N_14212);
nand UO_847 (O_847,N_12468,N_12616);
xnor UO_848 (O_848,N_14452,N_14820);
or UO_849 (O_849,N_13294,N_13756);
nand UO_850 (O_850,N_13394,N_12819);
nor UO_851 (O_851,N_14877,N_13851);
nor UO_852 (O_852,N_14276,N_13980);
and UO_853 (O_853,N_12402,N_12773);
or UO_854 (O_854,N_14983,N_14132);
nand UO_855 (O_855,N_12267,N_14838);
nor UO_856 (O_856,N_13832,N_12497);
and UO_857 (O_857,N_14559,N_12076);
nor UO_858 (O_858,N_12851,N_12137);
or UO_859 (O_859,N_13064,N_13549);
nand UO_860 (O_860,N_13602,N_14368);
or UO_861 (O_861,N_13580,N_14813);
nand UO_862 (O_862,N_13397,N_14797);
and UO_863 (O_863,N_14425,N_14267);
nor UO_864 (O_864,N_13163,N_13450);
nor UO_865 (O_865,N_14731,N_14333);
and UO_866 (O_866,N_13252,N_14517);
nand UO_867 (O_867,N_12274,N_13950);
nand UO_868 (O_868,N_13080,N_13714);
or UO_869 (O_869,N_12925,N_12427);
or UO_870 (O_870,N_14741,N_12470);
and UO_871 (O_871,N_13843,N_14803);
or UO_872 (O_872,N_14570,N_12413);
and UO_873 (O_873,N_12383,N_12253);
nand UO_874 (O_874,N_13844,N_13243);
and UO_875 (O_875,N_14394,N_14835);
nor UO_876 (O_876,N_12291,N_13696);
or UO_877 (O_877,N_12301,N_14028);
nor UO_878 (O_878,N_14214,N_13149);
and UO_879 (O_879,N_13622,N_12326);
and UO_880 (O_880,N_14775,N_14909);
or UO_881 (O_881,N_13658,N_13716);
and UO_882 (O_882,N_12334,N_13023);
and UO_883 (O_883,N_13850,N_12775);
or UO_884 (O_884,N_13144,N_13745);
nand UO_885 (O_885,N_13332,N_13798);
and UO_886 (O_886,N_12008,N_13121);
nor UO_887 (O_887,N_12728,N_13470);
nand UO_888 (O_888,N_12880,N_13013);
nand UO_889 (O_889,N_13570,N_12480);
nand UO_890 (O_890,N_12541,N_14166);
nand UO_891 (O_891,N_12209,N_14544);
or UO_892 (O_892,N_13876,N_12159);
or UO_893 (O_893,N_13504,N_14040);
nand UO_894 (O_894,N_12832,N_12723);
or UO_895 (O_895,N_12245,N_13799);
or UO_896 (O_896,N_12375,N_14123);
nand UO_897 (O_897,N_13454,N_14279);
or UO_898 (O_898,N_13713,N_13998);
nand UO_899 (O_899,N_13355,N_14310);
nor UO_900 (O_900,N_14052,N_13865);
nor UO_901 (O_901,N_12629,N_14562);
nor UO_902 (O_902,N_14210,N_12166);
and UO_903 (O_903,N_12303,N_13722);
nor UO_904 (O_904,N_14515,N_12920);
or UO_905 (O_905,N_13275,N_14538);
nand UO_906 (O_906,N_12389,N_13130);
or UO_907 (O_907,N_12113,N_14799);
or UO_908 (O_908,N_14218,N_14585);
nor UO_909 (O_909,N_14062,N_14072);
or UO_910 (O_910,N_14732,N_14255);
or UO_911 (O_911,N_14482,N_13123);
or UO_912 (O_912,N_14092,N_12958);
and UO_913 (O_913,N_13793,N_13925);
and UO_914 (O_914,N_12873,N_12604);
or UO_915 (O_915,N_14948,N_13337);
nor UO_916 (O_916,N_12222,N_14221);
nor UO_917 (O_917,N_13408,N_14154);
nand UO_918 (O_918,N_13752,N_12887);
nor UO_919 (O_919,N_12931,N_14656);
and UO_920 (O_920,N_14847,N_14461);
and UO_921 (O_921,N_12625,N_14101);
nand UO_922 (O_922,N_14104,N_12378);
nand UO_923 (O_923,N_12308,N_13741);
nor UO_924 (O_924,N_12400,N_12557);
and UO_925 (O_925,N_13088,N_12096);
nand UO_926 (O_926,N_12704,N_14115);
and UO_927 (O_927,N_13218,N_13371);
or UO_928 (O_928,N_14913,N_12035);
nand UO_929 (O_929,N_12946,N_12476);
nand UO_930 (O_930,N_12425,N_14848);
nor UO_931 (O_931,N_12703,N_13407);
and UO_932 (O_932,N_14727,N_13841);
and UO_933 (O_933,N_12648,N_13835);
nand UO_934 (O_934,N_13383,N_14155);
nor UO_935 (O_935,N_14875,N_14539);
and UO_936 (O_936,N_13833,N_14422);
nor UO_937 (O_937,N_14766,N_14800);
and UO_938 (O_938,N_12421,N_13601);
and UO_939 (O_939,N_13933,N_13483);
and UO_940 (O_940,N_14135,N_14992);
or UO_941 (O_941,N_13837,N_12024);
or UO_942 (O_942,N_14943,N_13147);
and UO_943 (O_943,N_13467,N_12523);
and UO_944 (O_944,N_12347,N_13937);
nand UO_945 (O_945,N_12562,N_14901);
nand UO_946 (O_946,N_13391,N_12797);
nand UO_947 (O_947,N_14907,N_13399);
and UO_948 (O_948,N_13400,N_14034);
or UO_949 (O_949,N_14952,N_14605);
or UO_950 (O_950,N_13788,N_14180);
nand UO_951 (O_951,N_12273,N_12894);
nand UO_952 (O_952,N_14922,N_12414);
nand UO_953 (O_953,N_13205,N_13649);
nor UO_954 (O_954,N_12915,N_14495);
nor UO_955 (O_955,N_13438,N_14676);
or UO_956 (O_956,N_12229,N_14430);
or UO_957 (O_957,N_12721,N_14271);
nor UO_958 (O_958,N_12386,N_13010);
or UO_959 (O_959,N_13474,N_13702);
nand UO_960 (O_960,N_13131,N_12668);
nor UO_961 (O_961,N_13828,N_12843);
or UO_962 (O_962,N_14791,N_12133);
nand UO_963 (O_963,N_12766,N_12733);
nor UO_964 (O_964,N_12785,N_13258);
nor UO_965 (O_965,N_12371,N_12036);
nand UO_966 (O_966,N_14446,N_14624);
nor UO_967 (O_967,N_12459,N_12264);
or UO_968 (O_968,N_14186,N_13035);
or UO_969 (O_969,N_12205,N_14524);
nor UO_970 (O_970,N_13432,N_13314);
or UO_971 (O_971,N_13955,N_14102);
and UO_972 (O_972,N_12217,N_12772);
or UO_973 (O_973,N_13973,N_13063);
nand UO_974 (O_974,N_14743,N_14823);
nor UO_975 (O_975,N_13683,N_12831);
nand UO_976 (O_976,N_12493,N_14871);
nand UO_977 (O_977,N_12321,N_13285);
and UO_978 (O_978,N_12487,N_14627);
and UO_979 (O_979,N_13595,N_14961);
or UO_980 (O_980,N_12848,N_14130);
nor UO_981 (O_981,N_14300,N_13892);
or UO_982 (O_982,N_14758,N_13429);
or UO_983 (O_983,N_14679,N_14330);
nand UO_984 (O_984,N_14671,N_12571);
or UO_985 (O_985,N_14635,N_13264);
nand UO_986 (O_986,N_14169,N_14674);
nor UO_987 (O_987,N_12033,N_12592);
and UO_988 (O_988,N_12657,N_13366);
nor UO_989 (O_989,N_12672,N_14471);
nor UO_990 (O_990,N_13168,N_14632);
or UO_991 (O_991,N_14301,N_13515);
nor UO_992 (O_992,N_12695,N_13958);
nor UO_993 (O_993,N_12878,N_12187);
and UO_994 (O_994,N_13611,N_12753);
and UO_995 (O_995,N_12112,N_13347);
nand UO_996 (O_996,N_12390,N_12952);
and UO_997 (O_997,N_14159,N_13732);
nand UO_998 (O_998,N_14574,N_14151);
nand UO_999 (O_999,N_13365,N_13078);
or UO_1000 (O_1000,N_12108,N_13935);
nand UO_1001 (O_1001,N_13405,N_13173);
or UO_1002 (O_1002,N_14989,N_14080);
or UO_1003 (O_1003,N_12005,N_12143);
nand UO_1004 (O_1004,N_13735,N_14964);
nor UO_1005 (O_1005,N_12426,N_14188);
nand UO_1006 (O_1006,N_13425,N_14064);
nand UO_1007 (O_1007,N_14663,N_12173);
nand UO_1008 (O_1008,N_14830,N_12017);
and UO_1009 (O_1009,N_13148,N_13154);
nor UO_1010 (O_1010,N_12945,N_13413);
xnor UO_1011 (O_1011,N_14885,N_14458);
nor UO_1012 (O_1012,N_14966,N_14416);
nand UO_1013 (O_1013,N_13484,N_12577);
or UO_1014 (O_1014,N_12130,N_14407);
or UO_1015 (O_1015,N_12175,N_13607);
or UO_1016 (O_1016,N_14463,N_12283);
or UO_1017 (O_1017,N_13321,N_12852);
or UO_1018 (O_1018,N_13770,N_13800);
or UO_1019 (O_1019,N_13384,N_12909);
nand UO_1020 (O_1020,N_13081,N_12309);
or UO_1021 (O_1021,N_12204,N_12066);
nand UO_1022 (O_1022,N_14962,N_13387);
nor UO_1023 (O_1023,N_14190,N_13189);
or UO_1024 (O_1024,N_12243,N_13646);
or UO_1025 (O_1025,N_14063,N_13059);
and UO_1026 (O_1026,N_12049,N_14478);
and UO_1027 (O_1027,N_14756,N_12860);
nand UO_1028 (O_1028,N_14771,N_12928);
and UO_1029 (O_1029,N_13125,N_12614);
nand UO_1030 (O_1030,N_12073,N_14206);
or UO_1031 (O_1031,N_14350,N_14369);
nand UO_1032 (O_1032,N_14468,N_14690);
or UO_1033 (O_1033,N_13863,N_14207);
nand UO_1034 (O_1034,N_12023,N_13573);
nor UO_1035 (O_1035,N_12235,N_13616);
nor UO_1036 (O_1036,N_14832,N_12227);
and UO_1037 (O_1037,N_12448,N_12346);
nor UO_1038 (O_1038,N_13442,N_13448);
or UO_1039 (O_1039,N_14254,N_13085);
or UO_1040 (O_1040,N_13823,N_14889);
and UO_1041 (O_1041,N_14383,N_13420);
nand UO_1042 (O_1042,N_13805,N_13296);
nand UO_1043 (O_1043,N_12263,N_13820);
nor UO_1044 (O_1044,N_14191,N_12465);
nand UO_1045 (O_1045,N_12115,N_14060);
nor UO_1046 (O_1046,N_14417,N_13963);
and UO_1047 (O_1047,N_14053,N_12063);
or UO_1048 (O_1048,N_13456,N_14958);
nand UO_1049 (O_1049,N_14234,N_14926);
nor UO_1050 (O_1050,N_14706,N_14591);
and UO_1051 (O_1051,N_13230,N_12061);
or UO_1052 (O_1052,N_12228,N_12010);
nand UO_1053 (O_1053,N_12582,N_13786);
or UO_1054 (O_1054,N_12305,N_12971);
nand UO_1055 (O_1055,N_13677,N_14553);
nor UO_1056 (O_1056,N_14144,N_13872);
nand UO_1057 (O_1057,N_12641,N_13857);
nor UO_1058 (O_1058,N_12464,N_14454);
or UO_1059 (O_1059,N_13787,N_12415);
or UO_1060 (O_1060,N_12125,N_12178);
nor UO_1061 (O_1061,N_13912,N_14579);
nor UO_1062 (O_1062,N_13045,N_14657);
nor UO_1063 (O_1063,N_12864,N_13600);
or UO_1064 (O_1064,N_13945,N_13526);
and UO_1065 (O_1065,N_14505,N_14116);
nor UO_1066 (O_1066,N_14443,N_13494);
nand UO_1067 (O_1067,N_14265,N_14421);
xnor UO_1068 (O_1068,N_14324,N_12606);
and UO_1069 (O_1069,N_13226,N_14121);
nand UO_1070 (O_1070,N_13221,N_13588);
nor UO_1071 (O_1071,N_14554,N_14935);
nor UO_1072 (O_1072,N_13653,N_14584);
and UO_1073 (O_1073,N_13307,N_14516);
nor UO_1074 (O_1074,N_14611,N_14260);
or UO_1075 (O_1075,N_12396,N_12691);
and UO_1076 (O_1076,N_12581,N_12701);
nor UO_1077 (O_1077,N_13393,N_13370);
and UO_1078 (O_1078,N_13172,N_14876);
and UO_1079 (O_1079,N_13447,N_14138);
nand UO_1080 (O_1080,N_13431,N_13692);
and UO_1081 (O_1081,N_12026,N_13234);
or UO_1082 (O_1082,N_13960,N_14360);
or UO_1083 (O_1083,N_12443,N_13190);
and UO_1084 (O_1084,N_13160,N_14499);
nand UO_1085 (O_1085,N_13417,N_13072);
and UO_1086 (O_1086,N_14641,N_12602);
nand UO_1087 (O_1087,N_12590,N_13598);
and UO_1088 (O_1088,N_14759,N_13717);
or UO_1089 (O_1089,N_13530,N_13771);
or UO_1090 (O_1090,N_13550,N_13972);
nand UO_1091 (O_1091,N_13201,N_13261);
nor UO_1092 (O_1092,N_14853,N_14261);
nor UO_1093 (O_1093,N_13132,N_14069);
nand UO_1094 (O_1094,N_13380,N_12556);
and UO_1095 (O_1095,N_12973,N_12726);
and UO_1096 (O_1096,N_14090,N_13938);
and UO_1097 (O_1097,N_14257,N_13545);
and UO_1098 (O_1098,N_12136,N_13845);
nor UO_1099 (O_1099,N_12643,N_13981);
nand UO_1100 (O_1100,N_12272,N_13200);
nand UO_1101 (O_1101,N_14000,N_14414);
or UO_1102 (O_1102,N_14015,N_12844);
nor UO_1103 (O_1103,N_14320,N_14710);
nor UO_1104 (O_1104,N_13754,N_13465);
or UO_1105 (O_1105,N_14094,N_13540);
or UO_1106 (O_1106,N_13572,N_13267);
and UO_1107 (O_1107,N_12677,N_13890);
nand UO_1108 (O_1108,N_13426,N_12237);
or UO_1109 (O_1109,N_12498,N_14792);
and UO_1110 (O_1110,N_12452,N_13457);
and UO_1111 (O_1111,N_14054,N_12219);
and UO_1112 (O_1112,N_13098,N_12509);
and UO_1113 (O_1113,N_13398,N_12483);
and UO_1114 (O_1114,N_12093,N_14082);
nor UO_1115 (O_1115,N_13506,N_13942);
and UO_1116 (O_1116,N_13738,N_12411);
nor UO_1117 (O_1117,N_13636,N_12900);
or UO_1118 (O_1118,N_14334,N_12620);
nand UO_1119 (O_1119,N_14680,N_13678);
and UO_1120 (O_1120,N_12545,N_14079);
nand UO_1121 (O_1121,N_14557,N_12752);
or UO_1122 (O_1122,N_14604,N_12508);
or UO_1123 (O_1123,N_12802,N_12502);
and UO_1124 (O_1124,N_12046,N_12755);
and UO_1125 (O_1125,N_13721,N_14640);
and UO_1126 (O_1126,N_13867,N_14513);
or UO_1127 (O_1127,N_13428,N_13977);
and UO_1128 (O_1128,N_12937,N_12433);
nand UO_1129 (O_1129,N_13174,N_14852);
or UO_1130 (O_1130,N_12647,N_12382);
nand UO_1131 (O_1131,N_12710,N_14865);
or UO_1132 (O_1132,N_12736,N_12835);
or UO_1133 (O_1133,N_13014,N_12926);
nand UO_1134 (O_1134,N_14608,N_13110);
nor UO_1135 (O_1135,N_12134,N_12600);
and UO_1136 (O_1136,N_12090,N_12404);
or UO_1137 (O_1137,N_13272,N_13477);
or UO_1138 (O_1138,N_12299,N_12466);
nor UO_1139 (O_1139,N_13422,N_14808);
nor UO_1140 (O_1140,N_14332,N_13359);
nor UO_1141 (O_1141,N_14928,N_12454);
nor UO_1142 (O_1142,N_13323,N_12570);
or UO_1143 (O_1143,N_12098,N_13362);
and UO_1144 (O_1144,N_12439,N_14384);
and UO_1145 (O_1145,N_12257,N_14693);
and UO_1146 (O_1146,N_12220,N_14003);
and UO_1147 (O_1147,N_12968,N_14193);
or UO_1148 (O_1148,N_12671,N_14596);
nor UO_1149 (O_1149,N_14231,N_13403);
or UO_1150 (O_1150,N_12956,N_12676);
nor UO_1151 (O_1151,N_12177,N_13804);
nand UO_1152 (O_1152,N_13435,N_12154);
and UO_1153 (O_1153,N_14045,N_14715);
nor UO_1154 (O_1154,N_14827,N_13896);
nand UO_1155 (O_1155,N_14643,N_14552);
or UO_1156 (O_1156,N_14580,N_12692);
and UO_1157 (O_1157,N_14500,N_14522);
and UO_1158 (O_1158,N_12373,N_13445);
and UO_1159 (O_1159,N_12825,N_13119);
nor UO_1160 (O_1160,N_12403,N_14312);
or UO_1161 (O_1161,N_14754,N_14946);
nor UO_1162 (O_1162,N_13891,N_12567);
and UO_1163 (O_1163,N_12381,N_13503);
or UO_1164 (O_1164,N_14085,N_14372);
nor UO_1165 (O_1165,N_13334,N_14866);
nor UO_1166 (O_1166,N_12139,N_13982);
or UO_1167 (O_1167,N_14873,N_14306);
nor UO_1168 (O_1168,N_14787,N_12745);
or UO_1169 (O_1169,N_12780,N_14248);
xnor UO_1170 (O_1170,N_14677,N_12110);
and UO_1171 (O_1171,N_12370,N_12126);
and UO_1172 (O_1172,N_13248,N_14917);
or UO_1173 (O_1173,N_14217,N_14007);
and UO_1174 (O_1174,N_13156,N_13674);
and UO_1175 (O_1175,N_14971,N_12627);
nor UO_1176 (O_1176,N_12798,N_13790);
nand UO_1177 (O_1177,N_14629,N_12300);
nor UO_1178 (O_1178,N_12510,N_12540);
nor UO_1179 (O_1179,N_13711,N_12336);
nand UO_1180 (O_1180,N_13005,N_14041);
nor UO_1181 (O_1181,N_12013,N_12806);
or UO_1182 (O_1182,N_13767,N_12660);
nand UO_1183 (O_1183,N_13142,N_14184);
nand UO_1184 (O_1184,N_13571,N_13701);
nand UO_1185 (O_1185,N_12339,N_12109);
or UO_1186 (O_1186,N_12208,N_14777);
nand UO_1187 (O_1187,N_14409,N_14979);
nand UO_1188 (O_1188,N_12155,N_13269);
nor UO_1189 (O_1189,N_13966,N_12064);
or UO_1190 (O_1190,N_14111,N_12686);
and UO_1191 (O_1191,N_12161,N_12913);
nor UO_1192 (O_1192,N_14699,N_14493);
nand UO_1193 (O_1193,N_13730,N_13875);
or UO_1194 (O_1194,N_14840,N_14213);
and UO_1195 (O_1195,N_14178,N_14106);
or UO_1196 (O_1196,N_12007,N_14582);
nor UO_1197 (O_1197,N_12089,N_12353);
nand UO_1198 (O_1198,N_13439,N_14386);
nand UO_1199 (O_1199,N_13495,N_13631);
nand UO_1200 (O_1200,N_12561,N_13609);
nor UO_1201 (O_1201,N_14220,N_14177);
or UO_1202 (O_1202,N_12840,N_14110);
nand UO_1203 (O_1203,N_14949,N_12936);
nand UO_1204 (O_1204,N_13242,N_14202);
or UO_1205 (O_1205,N_13086,N_12410);
nor UO_1206 (O_1206,N_13951,N_12769);
nor UO_1207 (O_1207,N_13613,N_12661);
or UO_1208 (O_1208,N_13326,N_12693);
nor UO_1209 (O_1209,N_12626,N_14793);
or UO_1210 (O_1210,N_12324,N_13989);
and UO_1211 (O_1211,N_14435,N_12360);
and UO_1212 (O_1212,N_14433,N_13746);
or UO_1213 (O_1213,N_12985,N_14309);
nor UO_1214 (O_1214,N_13150,N_14726);
and UO_1215 (O_1215,N_14428,N_13349);
or UO_1216 (O_1216,N_13525,N_12954);
and UO_1217 (O_1217,N_14118,N_13187);
nor UO_1218 (O_1218,N_13749,N_12119);
or UO_1219 (O_1219,N_12587,N_13385);
or UO_1220 (O_1220,N_12114,N_14317);
nor UO_1221 (O_1221,N_12032,N_14547);
nor UO_1222 (O_1222,N_12828,N_14967);
or UO_1223 (O_1223,N_12491,N_14864);
and UO_1224 (O_1224,N_13917,N_14197);
or UO_1225 (O_1225,N_14136,N_14032);
nor UO_1226 (O_1226,N_13900,N_12144);
or UO_1227 (O_1227,N_12977,N_14951);
nand UO_1228 (O_1228,N_12236,N_14019);
nor UO_1229 (O_1229,N_12331,N_13710);
nand UO_1230 (O_1230,N_14125,N_12397);
or UO_1231 (O_1231,N_14764,N_13278);
or UO_1232 (O_1232,N_12355,N_14247);
and UO_1233 (O_1233,N_13908,N_13910);
nand UO_1234 (O_1234,N_12420,N_12162);
nand UO_1235 (O_1235,N_14765,N_14899);
nor UO_1236 (O_1236,N_12534,N_14204);
nand UO_1237 (O_1237,N_13472,N_12477);
and UO_1238 (O_1238,N_12694,N_14982);
and UO_1239 (O_1239,N_12103,N_13479);
nor UO_1240 (O_1240,N_12463,N_14923);
nor UO_1241 (O_1241,N_12102,N_12748);
nor UO_1242 (O_1242,N_14016,N_13087);
or UO_1243 (O_1243,N_12311,N_13030);
and UO_1244 (O_1244,N_13943,N_14742);
xor UO_1245 (O_1245,N_13453,N_13096);
nand UO_1246 (O_1246,N_14814,N_13842);
nor UO_1247 (O_1247,N_14686,N_13093);
nand UO_1248 (O_1248,N_12836,N_14281);
nor UO_1249 (O_1249,N_12628,N_12354);
and UO_1250 (O_1250,N_12829,N_13553);
or UO_1251 (O_1251,N_14029,N_12083);
nand UO_1252 (O_1252,N_14661,N_13524);
or UO_1253 (O_1253,N_14020,N_12566);
or UO_1254 (O_1254,N_14684,N_13564);
and UO_1255 (O_1255,N_14714,N_14031);
nand UO_1256 (O_1256,N_12816,N_14150);
nand UO_1257 (O_1257,N_13682,N_13124);
nand UO_1258 (O_1258,N_13034,N_12041);
or UO_1259 (O_1259,N_13029,N_13181);
and UO_1260 (O_1260,N_12560,N_12029);
xor UO_1261 (O_1261,N_13810,N_13585);
or UO_1262 (O_1262,N_12612,N_13122);
nor UO_1263 (O_1263,N_13204,N_12270);
nand UO_1264 (O_1264,N_12714,N_12268);
or UO_1265 (O_1265,N_12632,N_14318);
nor UO_1266 (O_1266,N_13396,N_14626);
or UO_1267 (O_1267,N_14660,N_14890);
nand UO_1268 (O_1268,N_13510,N_14161);
and UO_1269 (O_1269,N_14450,N_13694);
and UO_1270 (O_1270,N_13517,N_14790);
nand UO_1271 (O_1271,N_12348,N_13885);
nand UO_1272 (O_1272,N_13887,N_14061);
nor UO_1273 (O_1273,N_13727,N_13995);
and UO_1274 (O_1274,N_14286,N_12800);
or UO_1275 (O_1275,N_14927,N_14506);
nand UO_1276 (O_1276,N_14401,N_12149);
nand UO_1277 (O_1277,N_12522,N_12180);
or UO_1278 (O_1278,N_13691,N_13112);
nand UO_1279 (O_1279,N_13608,N_12911);
nand UO_1280 (O_1280,N_14805,N_13838);
nor UO_1281 (O_1281,N_13306,N_13169);
or UO_1282 (O_1282,N_14081,N_13523);
and UO_1283 (O_1283,N_12450,N_13061);
or UO_1284 (O_1284,N_12275,N_13175);
or UO_1285 (O_1285,N_12057,N_12743);
and UO_1286 (O_1286,N_13944,N_13715);
nor UO_1287 (O_1287,N_14869,N_13379);
nor UO_1288 (O_1288,N_13597,N_14352);
nor UO_1289 (O_1289,N_13262,N_13797);
and UO_1290 (O_1290,N_12863,N_13625);
and UO_1291 (O_1291,N_14816,N_14442);
nand UO_1292 (O_1292,N_13516,N_14278);
nor UO_1293 (O_1293,N_13203,N_13418);
nand UO_1294 (O_1294,N_14855,N_13928);
nand UO_1295 (O_1295,N_14444,N_14973);
nand UO_1296 (O_1296,N_12356,N_14666);
nor UO_1297 (O_1297,N_13986,N_14134);
and UO_1298 (O_1298,N_14148,N_14700);
or UO_1299 (O_1299,N_13577,N_12867);
and UO_1300 (O_1300,N_14296,N_12807);
or UO_1301 (O_1301,N_14323,N_12927);
or UO_1302 (O_1302,N_12654,N_13544);
or UO_1303 (O_1303,N_13388,N_14358);
nand UO_1304 (O_1304,N_14767,N_13906);
and UO_1305 (O_1305,N_13569,N_12395);
nor UO_1306 (O_1306,N_14843,N_14076);
and UO_1307 (O_1307,N_13895,N_12678);
nand UO_1308 (O_1308,N_13331,N_12953);
and UO_1309 (O_1309,N_14047,N_12563);
nand UO_1310 (O_1310,N_14377,N_13656);
nor UO_1311 (O_1311,N_13193,N_13137);
and UO_1312 (O_1312,N_14811,N_12310);
nand UO_1313 (O_1313,N_13090,N_13402);
or UO_1314 (O_1314,N_13055,N_12515);
or UO_1315 (O_1315,N_12281,N_13834);
nand UO_1316 (O_1316,N_13869,N_14100);
nor UO_1317 (O_1317,N_14563,N_12207);
or UO_1318 (O_1318,N_12058,N_13127);
nor UO_1319 (O_1319,N_14682,N_12475);
and UO_1320 (O_1320,N_12760,N_12232);
nor UO_1321 (O_1321,N_12327,N_12905);
nand UO_1322 (O_1322,N_12902,N_13681);
and UO_1323 (O_1323,N_12472,N_12989);
nor UO_1324 (O_1324,N_12315,N_14170);
and UO_1325 (O_1325,N_12889,N_12231);
nand UO_1326 (O_1326,N_12664,N_12519);
or UO_1327 (O_1327,N_13356,N_12574);
and UO_1328 (O_1328,N_14036,N_13618);
nor UO_1329 (O_1329,N_14602,N_14897);
or UO_1330 (O_1330,N_12244,N_13743);
nor UO_1331 (O_1331,N_13481,N_12290);
or UO_1332 (O_1332,N_13335,N_12544);
nand UO_1333 (O_1333,N_13106,N_13522);
nand UO_1334 (O_1334,N_14058,N_14237);
and UO_1335 (O_1335,N_14490,N_12135);
and UO_1336 (O_1336,N_14183,N_12568);
and UO_1337 (O_1337,N_12943,N_14239);
and UO_1338 (O_1338,N_13764,N_13184);
nand UO_1339 (O_1339,N_13736,N_13255);
nor UO_1340 (O_1340,N_12921,N_13819);
and UO_1341 (O_1341,N_12319,N_13038);
nand UO_1342 (O_1342,N_14683,N_14353);
or UO_1343 (O_1343,N_12877,N_13742);
and UO_1344 (O_1344,N_14858,N_13647);
or UO_1345 (O_1345,N_14606,N_14650);
and UO_1346 (O_1346,N_13490,N_13557);
nand UO_1347 (O_1347,N_14937,N_12412);
and UO_1348 (O_1348,N_14284,N_14628);
and UO_1349 (O_1349,N_14017,N_13216);
nand UO_1350 (O_1350,N_13183,N_12531);
and UO_1351 (O_1351,N_13654,N_14005);
and UO_1352 (O_1352,N_13158,N_13688);
nand UO_1353 (O_1353,N_13894,N_13464);
nor UO_1354 (O_1354,N_12011,N_14142);
nand UO_1355 (O_1355,N_13430,N_13440);
or UO_1356 (O_1356,N_12859,N_14427);
nor UO_1357 (O_1357,N_13988,N_13679);
and UO_1358 (O_1358,N_13703,N_12974);
nor UO_1359 (O_1359,N_12197,N_12713);
and UO_1360 (O_1360,N_13056,N_12430);
nand UO_1361 (O_1361,N_14074,N_14786);
or UO_1362 (O_1362,N_13015,N_12092);
nand UO_1363 (O_1363,N_14782,N_13020);
and UO_1364 (O_1364,N_13135,N_12898);
nor UO_1365 (O_1365,N_13987,N_13576);
and UO_1366 (O_1366,N_12924,N_13888);
nand UO_1367 (O_1367,N_13930,N_12855);
xor UO_1368 (O_1368,N_13363,N_14133);
nand UO_1369 (O_1369,N_13563,N_14802);
nand UO_1370 (O_1370,N_12405,N_14528);
and UO_1371 (O_1371,N_12376,N_12526);
nor UO_1372 (O_1372,N_12192,N_14728);
nor UO_1373 (O_1373,N_12214,N_13026);
or UO_1374 (O_1374,N_14182,N_14037);
or UO_1375 (O_1375,N_13455,N_14839);
nor UO_1376 (O_1376,N_12000,N_13009);
and UO_1377 (O_1377,N_14477,N_14339);
and UO_1378 (O_1378,N_12983,N_13500);
nor UO_1379 (O_1379,N_14065,N_14886);
and UO_1380 (O_1380,N_14688,N_13969);
and UO_1381 (O_1381,N_14809,N_14744);
nand UO_1382 (O_1382,N_14940,N_14012);
and UO_1383 (O_1383,N_12978,N_14551);
nand UO_1384 (O_1384,N_12367,N_14654);
nor UO_1385 (O_1385,N_12850,N_13463);
xnor UO_1386 (O_1386,N_13468,N_14906);
nand UO_1387 (O_1387,N_13000,N_13931);
nand UO_1388 (O_1388,N_13114,N_14589);
xor UO_1389 (O_1389,N_14779,N_14292);
nor UO_1390 (O_1390,N_14325,N_12505);
nand UO_1391 (O_1391,N_13208,N_14302);
or UO_1392 (O_1392,N_14340,N_13113);
nand UO_1393 (O_1393,N_12099,N_13671);
or UO_1394 (O_1394,N_14313,N_13822);
and UO_1395 (O_1395,N_14426,N_12858);
and UO_1396 (O_1396,N_14059,N_13179);
or UO_1397 (O_1397,N_13868,N_14784);
nand UO_1398 (O_1398,N_13645,N_13639);
and UO_1399 (O_1399,N_14225,N_14616);
or UO_1400 (O_1400,N_12964,N_12986);
nor UO_1401 (O_1401,N_12279,N_14667);
nand UO_1402 (O_1402,N_13128,N_12004);
nor UO_1403 (O_1403,N_12127,N_13265);
nor UO_1404 (O_1404,N_14561,N_14647);
and UO_1405 (O_1405,N_13640,N_12203);
nand UO_1406 (O_1406,N_12690,N_14850);
nor UO_1407 (O_1407,N_14164,N_13461);
and UO_1408 (O_1408,N_12803,N_12712);
and UO_1409 (O_1409,N_12717,N_12707);
or UO_1410 (O_1410,N_13073,N_14954);
or UO_1411 (O_1411,N_14942,N_13898);
or UO_1412 (O_1412,N_12052,N_12406);
or UO_1413 (O_1413,N_12934,N_13882);
nor UO_1414 (O_1414,N_13140,N_13057);
and UO_1415 (O_1415,N_14487,N_14918);
nand UO_1416 (O_1416,N_13700,N_14998);
nand UO_1417 (O_1417,N_14533,N_14568);
and UO_1418 (O_1418,N_14067,N_13539);
and UO_1419 (O_1419,N_14035,N_12768);
nand UO_1420 (O_1420,N_13555,N_14441);
xnor UO_1421 (O_1421,N_14112,N_14447);
or UO_1422 (O_1422,N_12685,N_12329);
or UO_1423 (O_1423,N_12146,N_12520);
or UO_1424 (O_1424,N_12256,N_12536);
or UO_1425 (O_1425,N_14406,N_12635);
nor UO_1426 (O_1426,N_13069,N_13273);
and UO_1427 (O_1427,N_13250,N_14807);
nand UO_1428 (O_1428,N_13480,N_14625);
nor UO_1429 (O_1429,N_14459,N_14733);
and UO_1430 (O_1430,N_13686,N_13471);
nor UO_1431 (O_1431,N_13508,N_12218);
or UO_1432 (O_1432,N_13594,N_13546);
nor UO_1433 (O_1433,N_12942,N_13776);
or UO_1434 (O_1434,N_12938,N_12874);
or UO_1435 (O_1435,N_13120,N_14986);
nand UO_1436 (O_1436,N_13361,N_13368);
nor UO_1437 (O_1437,N_12082,N_13485);
or UO_1438 (O_1438,N_13382,N_12031);
or UO_1439 (O_1439,N_13946,N_12622);
nand UO_1440 (O_1440,N_12575,N_13018);
nand UO_1441 (O_1441,N_13360,N_12957);
and UO_1442 (O_1442,N_14612,N_12535);
nor UO_1443 (O_1443,N_14269,N_13348);
and UO_1444 (O_1444,N_12363,N_13971);
nor UO_1445 (O_1445,N_13779,N_13848);
or UO_1446 (O_1446,N_13501,N_13146);
nor UO_1447 (O_1447,N_13079,N_13231);
nand UO_1448 (O_1448,N_14457,N_14904);
nor UO_1449 (O_1449,N_14295,N_12537);
nand UO_1450 (O_1450,N_13552,N_14227);
and UO_1451 (O_1451,N_12749,N_13919);
or UO_1452 (O_1452,N_12295,N_12793);
nor UO_1453 (O_1453,N_13811,N_14187);
nand UO_1454 (O_1454,N_14322,N_13768);
nor UO_1455 (O_1455,N_14305,N_14347);
nand UO_1456 (O_1456,N_14774,N_13107);
or UO_1457 (O_1457,N_12949,N_14152);
or UO_1458 (O_1458,N_13809,N_13792);
nand UO_1459 (O_1459,N_14723,N_12247);
and UO_1460 (O_1460,N_13709,N_13493);
xnor UO_1461 (O_1461,N_13567,N_13287);
nor UO_1462 (O_1462,N_13513,N_14896);
and UO_1463 (O_1463,N_13410,N_12794);
and UO_1464 (O_1464,N_14590,N_12416);
nor UO_1465 (O_1465,N_14819,N_13322);
nor UO_1466 (O_1466,N_12624,N_14749);
and UO_1467 (O_1467,N_12359,N_13708);
nand UO_1468 (O_1468,N_14828,N_14664);
nor UO_1469 (O_1469,N_12765,N_13104);
nor UO_1470 (O_1470,N_14341,N_13902);
and UO_1471 (O_1471,N_14924,N_13192);
nand UO_1472 (O_1472,N_12312,N_13414);
nand UO_1473 (O_1473,N_12361,N_14750);
and UO_1474 (O_1474,N_12734,N_12724);
or UO_1475 (O_1475,N_13139,N_14070);
nor UO_1476 (O_1476,N_13024,N_12081);
and UO_1477 (O_1477,N_14044,N_13342);
or UO_1478 (O_1478,N_12345,N_12306);
or UO_1479 (O_1479,N_13260,N_14999);
or UO_1480 (O_1480,N_12223,N_12422);
and UO_1481 (O_1481,N_14137,N_14636);
nand UO_1482 (O_1482,N_12837,N_12572);
or UO_1483 (O_1483,N_12659,N_12914);
and UO_1484 (O_1484,N_13381,N_12790);
nand UO_1485 (O_1485,N_13915,N_12186);
or UO_1486 (O_1486,N_14912,N_13590);
or UO_1487 (O_1487,N_13663,N_13202);
nor UO_1488 (O_1488,N_13162,N_14514);
nand UO_1489 (O_1489,N_13076,N_12020);
and UO_1490 (O_1490,N_14978,N_12153);
nor UO_1491 (O_1491,N_12891,N_13028);
or UO_1492 (O_1492,N_14968,N_13060);
nor UO_1493 (O_1493,N_13249,N_12317);
or UO_1494 (O_1494,N_13623,N_14083);
nand UO_1495 (O_1495,N_12916,N_13633);
or UO_1496 (O_1496,N_13212,N_13970);
nor UO_1497 (O_1497,N_13734,N_14215);
nor UO_1498 (O_1498,N_14006,N_13194);
xnor UO_1499 (O_1499,N_13305,N_12169);
or UO_1500 (O_1500,N_12905,N_12398);
and UO_1501 (O_1501,N_14081,N_12710);
nand UO_1502 (O_1502,N_14547,N_14358);
xnor UO_1503 (O_1503,N_14206,N_13059);
nor UO_1504 (O_1504,N_12353,N_12854);
nor UO_1505 (O_1505,N_12610,N_13393);
or UO_1506 (O_1506,N_13899,N_13606);
nand UO_1507 (O_1507,N_14421,N_13339);
or UO_1508 (O_1508,N_12618,N_14843);
nand UO_1509 (O_1509,N_13901,N_12215);
nand UO_1510 (O_1510,N_12213,N_13199);
nand UO_1511 (O_1511,N_12931,N_13672);
nor UO_1512 (O_1512,N_13514,N_12043);
and UO_1513 (O_1513,N_14719,N_12247);
nand UO_1514 (O_1514,N_14213,N_13076);
nor UO_1515 (O_1515,N_13817,N_13763);
or UO_1516 (O_1516,N_13391,N_14656);
and UO_1517 (O_1517,N_14176,N_12616);
nand UO_1518 (O_1518,N_12960,N_13634);
nand UO_1519 (O_1519,N_12194,N_12387);
nor UO_1520 (O_1520,N_12775,N_12615);
nand UO_1521 (O_1521,N_13034,N_14788);
or UO_1522 (O_1522,N_12708,N_13040);
and UO_1523 (O_1523,N_13218,N_12065);
nor UO_1524 (O_1524,N_13564,N_14799);
or UO_1525 (O_1525,N_12647,N_13637);
and UO_1526 (O_1526,N_12003,N_14565);
nor UO_1527 (O_1527,N_13327,N_14978);
nor UO_1528 (O_1528,N_14360,N_12576);
and UO_1529 (O_1529,N_12104,N_14058);
and UO_1530 (O_1530,N_13552,N_12262);
and UO_1531 (O_1531,N_13725,N_13161);
nor UO_1532 (O_1532,N_14924,N_14159);
and UO_1533 (O_1533,N_13609,N_13453);
nand UO_1534 (O_1534,N_12268,N_12224);
nand UO_1535 (O_1535,N_14607,N_12333);
or UO_1536 (O_1536,N_13104,N_12329);
nand UO_1537 (O_1537,N_12293,N_14994);
nand UO_1538 (O_1538,N_14544,N_14453);
nor UO_1539 (O_1539,N_13732,N_14903);
and UO_1540 (O_1540,N_14210,N_12543);
and UO_1541 (O_1541,N_13386,N_12072);
and UO_1542 (O_1542,N_13406,N_14506);
nor UO_1543 (O_1543,N_12520,N_13365);
or UO_1544 (O_1544,N_12246,N_12266);
or UO_1545 (O_1545,N_14061,N_14845);
and UO_1546 (O_1546,N_12681,N_13989);
nor UO_1547 (O_1547,N_12849,N_14056);
and UO_1548 (O_1548,N_14817,N_14532);
or UO_1549 (O_1549,N_12375,N_14825);
nand UO_1550 (O_1550,N_12191,N_12906);
nor UO_1551 (O_1551,N_14304,N_13829);
nand UO_1552 (O_1552,N_13162,N_12104);
or UO_1553 (O_1553,N_12572,N_14312);
nand UO_1554 (O_1554,N_14835,N_14615);
and UO_1555 (O_1555,N_14052,N_12465);
nand UO_1556 (O_1556,N_13129,N_14652);
nand UO_1557 (O_1557,N_13086,N_13125);
and UO_1558 (O_1558,N_12135,N_14227);
and UO_1559 (O_1559,N_12521,N_13802);
nor UO_1560 (O_1560,N_12671,N_14461);
or UO_1561 (O_1561,N_14104,N_14902);
and UO_1562 (O_1562,N_13539,N_13403);
nand UO_1563 (O_1563,N_14280,N_14694);
or UO_1564 (O_1564,N_12660,N_13657);
nand UO_1565 (O_1565,N_12008,N_14835);
and UO_1566 (O_1566,N_12796,N_12697);
and UO_1567 (O_1567,N_13267,N_14999);
nor UO_1568 (O_1568,N_12358,N_14639);
or UO_1569 (O_1569,N_14950,N_14436);
and UO_1570 (O_1570,N_14281,N_14190);
nand UO_1571 (O_1571,N_12747,N_13439);
and UO_1572 (O_1572,N_14761,N_13489);
or UO_1573 (O_1573,N_12123,N_13544);
nor UO_1574 (O_1574,N_13343,N_12651);
and UO_1575 (O_1575,N_13972,N_13886);
nor UO_1576 (O_1576,N_14212,N_14431);
or UO_1577 (O_1577,N_12559,N_14622);
nand UO_1578 (O_1578,N_12652,N_12434);
and UO_1579 (O_1579,N_13184,N_13100);
and UO_1580 (O_1580,N_14522,N_12127);
nor UO_1581 (O_1581,N_14223,N_12941);
nand UO_1582 (O_1582,N_13389,N_14105);
nand UO_1583 (O_1583,N_12928,N_12778);
or UO_1584 (O_1584,N_12087,N_13668);
and UO_1585 (O_1585,N_12484,N_13382);
and UO_1586 (O_1586,N_13123,N_14869);
or UO_1587 (O_1587,N_13470,N_12578);
nand UO_1588 (O_1588,N_13620,N_14709);
nand UO_1589 (O_1589,N_14236,N_14426);
and UO_1590 (O_1590,N_13212,N_14844);
or UO_1591 (O_1591,N_12050,N_13179);
or UO_1592 (O_1592,N_12912,N_13876);
and UO_1593 (O_1593,N_13440,N_14734);
nand UO_1594 (O_1594,N_13692,N_12000);
nor UO_1595 (O_1595,N_13341,N_12285);
nand UO_1596 (O_1596,N_14006,N_12250);
or UO_1597 (O_1597,N_14545,N_14208);
and UO_1598 (O_1598,N_13636,N_13867);
or UO_1599 (O_1599,N_13970,N_14229);
or UO_1600 (O_1600,N_12700,N_14438);
nand UO_1601 (O_1601,N_13770,N_14692);
nand UO_1602 (O_1602,N_13276,N_13544);
and UO_1603 (O_1603,N_13660,N_13939);
and UO_1604 (O_1604,N_12614,N_14011);
or UO_1605 (O_1605,N_13796,N_14136);
nor UO_1606 (O_1606,N_12370,N_12468);
or UO_1607 (O_1607,N_14643,N_14784);
and UO_1608 (O_1608,N_14427,N_14349);
nor UO_1609 (O_1609,N_13838,N_14083);
or UO_1610 (O_1610,N_13857,N_12500);
nor UO_1611 (O_1611,N_12444,N_13826);
nand UO_1612 (O_1612,N_12203,N_12116);
or UO_1613 (O_1613,N_13054,N_12829);
and UO_1614 (O_1614,N_12523,N_14302);
nor UO_1615 (O_1615,N_12320,N_13904);
and UO_1616 (O_1616,N_12349,N_13165);
and UO_1617 (O_1617,N_12178,N_12209);
nand UO_1618 (O_1618,N_13396,N_14148);
nand UO_1619 (O_1619,N_12436,N_14525);
nand UO_1620 (O_1620,N_12254,N_14986);
nand UO_1621 (O_1621,N_14536,N_13755);
and UO_1622 (O_1622,N_12793,N_13718);
nor UO_1623 (O_1623,N_12595,N_12807);
nand UO_1624 (O_1624,N_13121,N_14274);
nand UO_1625 (O_1625,N_13836,N_12171);
or UO_1626 (O_1626,N_13993,N_14944);
nor UO_1627 (O_1627,N_12110,N_12030);
and UO_1628 (O_1628,N_14576,N_14218);
or UO_1629 (O_1629,N_14228,N_14514);
or UO_1630 (O_1630,N_13421,N_13345);
and UO_1631 (O_1631,N_12684,N_13479);
nor UO_1632 (O_1632,N_13709,N_14388);
or UO_1633 (O_1633,N_14794,N_14597);
nand UO_1634 (O_1634,N_14612,N_13378);
nand UO_1635 (O_1635,N_14528,N_12407);
and UO_1636 (O_1636,N_13488,N_14507);
or UO_1637 (O_1637,N_13119,N_14488);
nand UO_1638 (O_1638,N_14328,N_14718);
and UO_1639 (O_1639,N_13605,N_13425);
nor UO_1640 (O_1640,N_14659,N_14053);
nor UO_1641 (O_1641,N_13632,N_14905);
and UO_1642 (O_1642,N_13543,N_13934);
nand UO_1643 (O_1643,N_12771,N_13854);
or UO_1644 (O_1644,N_12289,N_13354);
nand UO_1645 (O_1645,N_14250,N_13330);
nand UO_1646 (O_1646,N_12910,N_14069);
and UO_1647 (O_1647,N_12135,N_12635);
nor UO_1648 (O_1648,N_12828,N_12192);
nand UO_1649 (O_1649,N_13932,N_13074);
nor UO_1650 (O_1650,N_14489,N_14077);
nand UO_1651 (O_1651,N_14234,N_14123);
nor UO_1652 (O_1652,N_12677,N_12044);
nor UO_1653 (O_1653,N_12726,N_12691);
and UO_1654 (O_1654,N_13865,N_14394);
or UO_1655 (O_1655,N_13537,N_12225);
and UO_1656 (O_1656,N_12909,N_12968);
nand UO_1657 (O_1657,N_12066,N_13373);
or UO_1658 (O_1658,N_14237,N_13070);
and UO_1659 (O_1659,N_14418,N_14975);
or UO_1660 (O_1660,N_14125,N_12924);
or UO_1661 (O_1661,N_12230,N_14556);
nor UO_1662 (O_1662,N_14386,N_14556);
nor UO_1663 (O_1663,N_13727,N_13556);
nand UO_1664 (O_1664,N_13835,N_13967);
or UO_1665 (O_1665,N_12409,N_12066);
or UO_1666 (O_1666,N_12541,N_14211);
or UO_1667 (O_1667,N_14069,N_12410);
or UO_1668 (O_1668,N_14643,N_12574);
nand UO_1669 (O_1669,N_14838,N_12268);
and UO_1670 (O_1670,N_14174,N_12520);
or UO_1671 (O_1671,N_13503,N_14304);
and UO_1672 (O_1672,N_14730,N_12729);
or UO_1673 (O_1673,N_13679,N_14014);
and UO_1674 (O_1674,N_12365,N_13664);
nor UO_1675 (O_1675,N_13735,N_12547);
nor UO_1676 (O_1676,N_12226,N_12511);
or UO_1677 (O_1677,N_13208,N_14835);
nor UO_1678 (O_1678,N_13754,N_13351);
or UO_1679 (O_1679,N_14181,N_13890);
nand UO_1680 (O_1680,N_13290,N_14660);
and UO_1681 (O_1681,N_13996,N_14250);
nand UO_1682 (O_1682,N_13807,N_14709);
nand UO_1683 (O_1683,N_12818,N_13485);
nand UO_1684 (O_1684,N_13688,N_13654);
and UO_1685 (O_1685,N_14654,N_13779);
xnor UO_1686 (O_1686,N_14760,N_13162);
nor UO_1687 (O_1687,N_13361,N_12232);
and UO_1688 (O_1688,N_13915,N_14110);
nor UO_1689 (O_1689,N_13495,N_12345);
and UO_1690 (O_1690,N_14303,N_12673);
xnor UO_1691 (O_1691,N_13130,N_13705);
nor UO_1692 (O_1692,N_12355,N_13143);
and UO_1693 (O_1693,N_14384,N_14631);
and UO_1694 (O_1694,N_13639,N_13586);
xnor UO_1695 (O_1695,N_12401,N_13847);
nor UO_1696 (O_1696,N_13445,N_13318);
nand UO_1697 (O_1697,N_13911,N_14032);
nor UO_1698 (O_1698,N_12083,N_12021);
nand UO_1699 (O_1699,N_13240,N_14307);
nand UO_1700 (O_1700,N_14841,N_13380);
or UO_1701 (O_1701,N_12213,N_14550);
and UO_1702 (O_1702,N_14748,N_12254);
nand UO_1703 (O_1703,N_13664,N_14844);
nand UO_1704 (O_1704,N_14945,N_12946);
or UO_1705 (O_1705,N_12428,N_14135);
or UO_1706 (O_1706,N_13588,N_14144);
nor UO_1707 (O_1707,N_12629,N_13651);
nor UO_1708 (O_1708,N_14981,N_12888);
and UO_1709 (O_1709,N_14767,N_14869);
nand UO_1710 (O_1710,N_12045,N_13577);
or UO_1711 (O_1711,N_13509,N_14021);
and UO_1712 (O_1712,N_14901,N_14137);
nand UO_1713 (O_1713,N_12773,N_14227);
and UO_1714 (O_1714,N_12664,N_14769);
or UO_1715 (O_1715,N_12480,N_14728);
nor UO_1716 (O_1716,N_12930,N_13356);
nand UO_1717 (O_1717,N_12030,N_12759);
nor UO_1718 (O_1718,N_12950,N_12165);
or UO_1719 (O_1719,N_13169,N_13397);
nor UO_1720 (O_1720,N_13781,N_12965);
and UO_1721 (O_1721,N_13034,N_14929);
and UO_1722 (O_1722,N_12546,N_14858);
and UO_1723 (O_1723,N_14385,N_14920);
nor UO_1724 (O_1724,N_12884,N_12123);
and UO_1725 (O_1725,N_14615,N_13387);
nor UO_1726 (O_1726,N_14793,N_13944);
and UO_1727 (O_1727,N_14184,N_13172);
nor UO_1728 (O_1728,N_12543,N_14830);
and UO_1729 (O_1729,N_14691,N_14002);
or UO_1730 (O_1730,N_14250,N_14135);
or UO_1731 (O_1731,N_13254,N_12389);
and UO_1732 (O_1732,N_12256,N_13505);
or UO_1733 (O_1733,N_14570,N_13387);
or UO_1734 (O_1734,N_12943,N_14141);
and UO_1735 (O_1735,N_14548,N_14006);
and UO_1736 (O_1736,N_12906,N_14001);
or UO_1737 (O_1737,N_13511,N_14430);
nand UO_1738 (O_1738,N_13156,N_12988);
nor UO_1739 (O_1739,N_12878,N_12369);
or UO_1740 (O_1740,N_12217,N_13804);
and UO_1741 (O_1741,N_13244,N_12610);
nand UO_1742 (O_1742,N_12856,N_14165);
xnor UO_1743 (O_1743,N_14420,N_12488);
nor UO_1744 (O_1744,N_14766,N_12499);
and UO_1745 (O_1745,N_13515,N_14062);
nand UO_1746 (O_1746,N_14924,N_13990);
nor UO_1747 (O_1747,N_14313,N_12824);
or UO_1748 (O_1748,N_12592,N_14503);
nand UO_1749 (O_1749,N_14619,N_12142);
or UO_1750 (O_1750,N_14686,N_13145);
and UO_1751 (O_1751,N_12301,N_14785);
nand UO_1752 (O_1752,N_14938,N_13974);
nor UO_1753 (O_1753,N_14307,N_14267);
or UO_1754 (O_1754,N_13835,N_12342);
nand UO_1755 (O_1755,N_12334,N_13347);
and UO_1756 (O_1756,N_13956,N_12115);
nor UO_1757 (O_1757,N_13166,N_12610);
and UO_1758 (O_1758,N_13873,N_14840);
nand UO_1759 (O_1759,N_13265,N_14823);
nand UO_1760 (O_1760,N_12317,N_12248);
nor UO_1761 (O_1761,N_12303,N_12688);
and UO_1762 (O_1762,N_14652,N_12808);
or UO_1763 (O_1763,N_14789,N_14502);
nand UO_1764 (O_1764,N_14849,N_14608);
nor UO_1765 (O_1765,N_13879,N_14195);
nor UO_1766 (O_1766,N_14768,N_12575);
and UO_1767 (O_1767,N_12505,N_14915);
or UO_1768 (O_1768,N_14082,N_13376);
nor UO_1769 (O_1769,N_12678,N_13819);
nor UO_1770 (O_1770,N_12654,N_13032);
nand UO_1771 (O_1771,N_13820,N_13305);
nand UO_1772 (O_1772,N_14187,N_12710);
nor UO_1773 (O_1773,N_12224,N_12094);
and UO_1774 (O_1774,N_12277,N_13521);
and UO_1775 (O_1775,N_13370,N_13639);
nor UO_1776 (O_1776,N_13510,N_13418);
nor UO_1777 (O_1777,N_13551,N_12953);
nand UO_1778 (O_1778,N_14334,N_12886);
and UO_1779 (O_1779,N_14565,N_12196);
or UO_1780 (O_1780,N_13648,N_12841);
nor UO_1781 (O_1781,N_13661,N_14397);
and UO_1782 (O_1782,N_14638,N_12900);
nor UO_1783 (O_1783,N_12194,N_14596);
nor UO_1784 (O_1784,N_14068,N_14526);
nor UO_1785 (O_1785,N_12854,N_12585);
nor UO_1786 (O_1786,N_14258,N_12565);
nor UO_1787 (O_1787,N_14106,N_14328);
and UO_1788 (O_1788,N_14952,N_13983);
and UO_1789 (O_1789,N_13651,N_12167);
nand UO_1790 (O_1790,N_13598,N_12862);
nand UO_1791 (O_1791,N_14707,N_12283);
and UO_1792 (O_1792,N_14984,N_12532);
or UO_1793 (O_1793,N_12450,N_13026);
and UO_1794 (O_1794,N_12712,N_14303);
and UO_1795 (O_1795,N_13283,N_13940);
and UO_1796 (O_1796,N_14519,N_12969);
nor UO_1797 (O_1797,N_13477,N_14730);
or UO_1798 (O_1798,N_13646,N_12758);
nand UO_1799 (O_1799,N_14664,N_12453);
or UO_1800 (O_1800,N_13209,N_14022);
and UO_1801 (O_1801,N_12841,N_14766);
or UO_1802 (O_1802,N_12786,N_12393);
or UO_1803 (O_1803,N_13883,N_12321);
and UO_1804 (O_1804,N_12063,N_12854);
or UO_1805 (O_1805,N_14561,N_14158);
nand UO_1806 (O_1806,N_14298,N_14414);
nor UO_1807 (O_1807,N_12117,N_14168);
and UO_1808 (O_1808,N_13347,N_13991);
nor UO_1809 (O_1809,N_12542,N_13032);
nor UO_1810 (O_1810,N_14000,N_13277);
and UO_1811 (O_1811,N_14616,N_12003);
or UO_1812 (O_1812,N_14566,N_14048);
nand UO_1813 (O_1813,N_14983,N_12491);
and UO_1814 (O_1814,N_13923,N_12471);
or UO_1815 (O_1815,N_14499,N_13595);
nand UO_1816 (O_1816,N_13698,N_12872);
and UO_1817 (O_1817,N_12398,N_14471);
or UO_1818 (O_1818,N_12673,N_12326);
or UO_1819 (O_1819,N_14648,N_13787);
and UO_1820 (O_1820,N_14464,N_13569);
and UO_1821 (O_1821,N_14265,N_13895);
and UO_1822 (O_1822,N_13166,N_14855);
or UO_1823 (O_1823,N_14611,N_13865);
nor UO_1824 (O_1824,N_13005,N_14230);
nor UO_1825 (O_1825,N_12727,N_14846);
nor UO_1826 (O_1826,N_12343,N_14599);
nand UO_1827 (O_1827,N_13546,N_12659);
nand UO_1828 (O_1828,N_14801,N_14646);
or UO_1829 (O_1829,N_13142,N_14591);
nor UO_1830 (O_1830,N_14424,N_14826);
nand UO_1831 (O_1831,N_13463,N_12014);
and UO_1832 (O_1832,N_13326,N_12178);
nand UO_1833 (O_1833,N_13657,N_14661);
and UO_1834 (O_1834,N_12852,N_14376);
nor UO_1835 (O_1835,N_12611,N_14667);
nor UO_1836 (O_1836,N_13508,N_12908);
and UO_1837 (O_1837,N_14159,N_14045);
and UO_1838 (O_1838,N_14051,N_12972);
nor UO_1839 (O_1839,N_14880,N_14905);
or UO_1840 (O_1840,N_14634,N_13219);
and UO_1841 (O_1841,N_14568,N_13268);
nand UO_1842 (O_1842,N_14346,N_13981);
and UO_1843 (O_1843,N_14422,N_13288);
nand UO_1844 (O_1844,N_12461,N_14300);
nor UO_1845 (O_1845,N_14295,N_12792);
nor UO_1846 (O_1846,N_13740,N_12710);
and UO_1847 (O_1847,N_14428,N_14299);
nor UO_1848 (O_1848,N_12302,N_14203);
nor UO_1849 (O_1849,N_13406,N_12781);
or UO_1850 (O_1850,N_12642,N_14901);
nand UO_1851 (O_1851,N_13185,N_13111);
or UO_1852 (O_1852,N_12013,N_13704);
nor UO_1853 (O_1853,N_13101,N_13925);
nor UO_1854 (O_1854,N_14071,N_14915);
nand UO_1855 (O_1855,N_14972,N_12224);
nor UO_1856 (O_1856,N_12840,N_12167);
nor UO_1857 (O_1857,N_14333,N_12220);
nor UO_1858 (O_1858,N_13317,N_14142);
nand UO_1859 (O_1859,N_12195,N_12636);
or UO_1860 (O_1860,N_14482,N_14080);
nor UO_1861 (O_1861,N_13196,N_12550);
and UO_1862 (O_1862,N_12477,N_12048);
nor UO_1863 (O_1863,N_13001,N_14560);
nand UO_1864 (O_1864,N_13430,N_14321);
and UO_1865 (O_1865,N_12669,N_13121);
nand UO_1866 (O_1866,N_13186,N_13321);
or UO_1867 (O_1867,N_14811,N_12213);
and UO_1868 (O_1868,N_14193,N_14644);
or UO_1869 (O_1869,N_13640,N_12582);
nand UO_1870 (O_1870,N_13259,N_13797);
nand UO_1871 (O_1871,N_14759,N_12018);
nand UO_1872 (O_1872,N_14784,N_12066);
nor UO_1873 (O_1873,N_14437,N_13767);
nor UO_1874 (O_1874,N_12892,N_13463);
nor UO_1875 (O_1875,N_13138,N_12692);
and UO_1876 (O_1876,N_14749,N_13268);
or UO_1877 (O_1877,N_13818,N_13722);
nor UO_1878 (O_1878,N_12551,N_12564);
and UO_1879 (O_1879,N_13657,N_12256);
or UO_1880 (O_1880,N_12591,N_13533);
or UO_1881 (O_1881,N_13986,N_12859);
and UO_1882 (O_1882,N_14370,N_14567);
xnor UO_1883 (O_1883,N_14017,N_13632);
and UO_1884 (O_1884,N_14052,N_13112);
and UO_1885 (O_1885,N_14873,N_13683);
nor UO_1886 (O_1886,N_12821,N_12430);
nand UO_1887 (O_1887,N_12527,N_14625);
nand UO_1888 (O_1888,N_13433,N_12665);
nand UO_1889 (O_1889,N_13000,N_14568);
or UO_1890 (O_1890,N_14671,N_13068);
and UO_1891 (O_1891,N_12809,N_14693);
nand UO_1892 (O_1892,N_12603,N_14709);
or UO_1893 (O_1893,N_13693,N_13348);
and UO_1894 (O_1894,N_13916,N_12297);
nand UO_1895 (O_1895,N_14326,N_13386);
nor UO_1896 (O_1896,N_12124,N_13364);
nor UO_1897 (O_1897,N_13350,N_14577);
nand UO_1898 (O_1898,N_12947,N_12547);
or UO_1899 (O_1899,N_13602,N_14567);
nor UO_1900 (O_1900,N_14344,N_13210);
nand UO_1901 (O_1901,N_14264,N_13013);
or UO_1902 (O_1902,N_12091,N_12255);
and UO_1903 (O_1903,N_12258,N_14547);
nor UO_1904 (O_1904,N_12554,N_14135);
and UO_1905 (O_1905,N_14834,N_14136);
nand UO_1906 (O_1906,N_14966,N_13499);
or UO_1907 (O_1907,N_14960,N_12315);
nor UO_1908 (O_1908,N_12366,N_14825);
or UO_1909 (O_1909,N_14462,N_13449);
or UO_1910 (O_1910,N_14683,N_14918);
nor UO_1911 (O_1911,N_13413,N_14358);
or UO_1912 (O_1912,N_13289,N_12620);
or UO_1913 (O_1913,N_12234,N_13495);
nor UO_1914 (O_1914,N_13083,N_13756);
and UO_1915 (O_1915,N_14739,N_12259);
or UO_1916 (O_1916,N_14925,N_13092);
nor UO_1917 (O_1917,N_13763,N_14763);
and UO_1918 (O_1918,N_12268,N_13445);
nor UO_1919 (O_1919,N_12425,N_13336);
and UO_1920 (O_1920,N_12306,N_13123);
or UO_1921 (O_1921,N_14953,N_14385);
nor UO_1922 (O_1922,N_13872,N_12907);
nor UO_1923 (O_1923,N_13146,N_12494);
or UO_1924 (O_1924,N_13033,N_12629);
nor UO_1925 (O_1925,N_14371,N_12854);
or UO_1926 (O_1926,N_12243,N_13234);
nor UO_1927 (O_1927,N_13811,N_12407);
nor UO_1928 (O_1928,N_14972,N_12924);
and UO_1929 (O_1929,N_14873,N_12264);
and UO_1930 (O_1930,N_13511,N_13401);
and UO_1931 (O_1931,N_13869,N_14755);
or UO_1932 (O_1932,N_13939,N_14378);
and UO_1933 (O_1933,N_13551,N_13629);
or UO_1934 (O_1934,N_12474,N_14673);
nand UO_1935 (O_1935,N_12655,N_14363);
nor UO_1936 (O_1936,N_12262,N_13706);
nor UO_1937 (O_1937,N_14719,N_13885);
nand UO_1938 (O_1938,N_13791,N_12032);
and UO_1939 (O_1939,N_12903,N_13234);
nor UO_1940 (O_1940,N_13184,N_14222);
and UO_1941 (O_1941,N_13777,N_14134);
nand UO_1942 (O_1942,N_14965,N_13082);
nor UO_1943 (O_1943,N_12287,N_12577);
and UO_1944 (O_1944,N_12894,N_12056);
or UO_1945 (O_1945,N_12748,N_13381);
nand UO_1946 (O_1946,N_12877,N_13537);
nand UO_1947 (O_1947,N_13967,N_12344);
nand UO_1948 (O_1948,N_12282,N_14409);
or UO_1949 (O_1949,N_14566,N_12802);
or UO_1950 (O_1950,N_13239,N_12156);
or UO_1951 (O_1951,N_12137,N_14275);
nor UO_1952 (O_1952,N_14330,N_13216);
or UO_1953 (O_1953,N_13400,N_14797);
and UO_1954 (O_1954,N_13974,N_14884);
or UO_1955 (O_1955,N_14207,N_14762);
nor UO_1956 (O_1956,N_14774,N_13056);
and UO_1957 (O_1957,N_13490,N_13739);
nand UO_1958 (O_1958,N_12058,N_14614);
nand UO_1959 (O_1959,N_13951,N_12623);
or UO_1960 (O_1960,N_14140,N_14696);
nand UO_1961 (O_1961,N_14968,N_13194);
nand UO_1962 (O_1962,N_14495,N_13307);
and UO_1963 (O_1963,N_13243,N_14476);
or UO_1964 (O_1964,N_12796,N_13704);
and UO_1965 (O_1965,N_14150,N_13332);
nor UO_1966 (O_1966,N_13969,N_13164);
and UO_1967 (O_1967,N_12589,N_13205);
nand UO_1968 (O_1968,N_13306,N_14844);
nor UO_1969 (O_1969,N_12767,N_13271);
nand UO_1970 (O_1970,N_12782,N_12057);
nor UO_1971 (O_1971,N_14040,N_12142);
and UO_1972 (O_1972,N_12007,N_14869);
or UO_1973 (O_1973,N_12552,N_14842);
nand UO_1974 (O_1974,N_13660,N_13667);
nand UO_1975 (O_1975,N_13977,N_12998);
and UO_1976 (O_1976,N_13189,N_12570);
nor UO_1977 (O_1977,N_12589,N_13540);
or UO_1978 (O_1978,N_12968,N_12546);
nand UO_1979 (O_1979,N_13778,N_14712);
nor UO_1980 (O_1980,N_12915,N_12665);
nand UO_1981 (O_1981,N_14023,N_12295);
or UO_1982 (O_1982,N_13035,N_12628);
and UO_1983 (O_1983,N_12508,N_14261);
and UO_1984 (O_1984,N_14223,N_14427);
and UO_1985 (O_1985,N_12664,N_14010);
nand UO_1986 (O_1986,N_12448,N_12196);
nor UO_1987 (O_1987,N_14732,N_12650);
nor UO_1988 (O_1988,N_14515,N_13023);
nand UO_1989 (O_1989,N_12754,N_14050);
nor UO_1990 (O_1990,N_12522,N_12563);
or UO_1991 (O_1991,N_14325,N_13105);
nor UO_1992 (O_1992,N_12529,N_13919);
nor UO_1993 (O_1993,N_14075,N_12152);
or UO_1994 (O_1994,N_12461,N_14676);
or UO_1995 (O_1995,N_14451,N_13729);
nand UO_1996 (O_1996,N_14840,N_12390);
and UO_1997 (O_1997,N_12977,N_14392);
and UO_1998 (O_1998,N_12713,N_13743);
nand UO_1999 (O_1999,N_14489,N_14776);
endmodule