module basic_500_3000_500_15_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_382,In_466);
and U1 (N_1,In_53,In_164);
nand U2 (N_2,In_273,In_486);
nor U3 (N_3,In_219,In_94);
or U4 (N_4,In_327,In_258);
nand U5 (N_5,In_121,In_422);
or U6 (N_6,In_122,In_3);
nor U7 (N_7,In_112,In_481);
and U8 (N_8,In_6,In_139);
nand U9 (N_9,In_189,In_363);
nand U10 (N_10,In_170,In_418);
nand U11 (N_11,In_476,In_407);
nand U12 (N_12,In_414,In_470);
or U13 (N_13,In_140,In_410);
and U14 (N_14,In_288,In_337);
nand U15 (N_15,In_372,In_235);
nand U16 (N_16,In_149,In_256);
xor U17 (N_17,In_1,In_283);
or U18 (N_18,In_161,In_428);
xor U19 (N_19,In_40,In_480);
nor U20 (N_20,In_276,In_157);
nor U21 (N_21,In_234,In_8);
and U22 (N_22,In_326,In_30);
or U23 (N_23,In_24,In_240);
xnor U24 (N_24,In_393,In_242);
xnor U25 (N_25,In_330,In_250);
nor U26 (N_26,In_284,In_346);
and U27 (N_27,In_493,In_33);
nor U28 (N_28,In_150,In_181);
nand U29 (N_29,In_387,In_299);
xnor U30 (N_30,In_453,In_148);
nor U31 (N_31,In_119,In_357);
and U32 (N_32,In_311,In_308);
and U33 (N_33,In_394,In_82);
nor U34 (N_34,In_39,In_179);
or U35 (N_35,In_177,In_430);
or U36 (N_36,In_472,In_19);
and U37 (N_37,In_4,In_59);
and U38 (N_38,In_236,In_305);
and U39 (N_39,In_404,In_265);
nand U40 (N_40,In_79,In_75);
and U41 (N_41,In_268,In_351);
xnor U42 (N_42,In_309,In_100);
or U43 (N_43,In_67,In_335);
nor U44 (N_44,In_98,In_319);
or U45 (N_45,In_312,In_445);
nand U46 (N_46,In_201,In_241);
or U47 (N_47,In_347,In_383);
nand U48 (N_48,In_434,In_130);
nor U49 (N_49,In_277,In_211);
nand U50 (N_50,In_377,In_341);
or U51 (N_51,In_446,In_187);
or U52 (N_52,In_498,In_190);
nor U53 (N_53,In_314,In_172);
and U54 (N_54,In_62,In_29);
nor U55 (N_55,In_208,In_448);
or U56 (N_56,In_301,In_171);
nor U57 (N_57,In_93,In_415);
and U58 (N_58,In_144,In_15);
or U59 (N_59,In_424,In_416);
and U60 (N_60,In_426,In_478);
xor U61 (N_61,In_120,In_359);
or U62 (N_62,In_460,In_12);
or U63 (N_63,In_35,In_266);
or U64 (N_64,In_125,In_248);
or U65 (N_65,In_74,In_361);
or U66 (N_66,In_197,In_70);
xor U67 (N_67,In_151,In_117);
nor U68 (N_68,In_88,In_21);
and U69 (N_69,In_267,In_465);
nand U70 (N_70,In_290,In_207);
and U71 (N_71,In_95,In_343);
nor U72 (N_72,In_46,In_63);
nor U73 (N_73,In_31,In_222);
and U74 (N_74,In_160,In_254);
nor U75 (N_75,In_229,In_73);
or U76 (N_76,In_362,In_396);
xnor U77 (N_77,In_375,In_405);
nand U78 (N_78,In_442,In_44);
nand U79 (N_79,In_7,In_247);
and U80 (N_80,In_191,In_60);
nor U81 (N_81,In_497,In_370);
nor U82 (N_82,In_444,In_141);
nand U83 (N_83,In_175,In_402);
nor U84 (N_84,In_477,In_84);
nand U85 (N_85,In_441,In_25);
or U86 (N_86,In_452,In_420);
or U87 (N_87,In_80,In_193);
nand U88 (N_88,In_376,In_495);
nor U89 (N_89,In_168,In_432);
or U90 (N_90,In_230,In_295);
nand U91 (N_91,In_218,In_342);
or U92 (N_92,In_65,In_163);
or U93 (N_93,In_102,In_281);
and U94 (N_94,In_491,In_315);
and U95 (N_95,In_439,In_304);
nand U96 (N_96,In_51,In_123);
nand U97 (N_97,In_440,In_239);
or U98 (N_98,In_228,In_313);
nor U99 (N_99,In_317,In_352);
and U100 (N_100,In_492,In_490);
or U101 (N_101,In_106,In_0);
and U102 (N_102,In_473,In_61);
and U103 (N_103,In_64,In_488);
nand U104 (N_104,In_105,In_300);
and U105 (N_105,In_464,In_145);
nor U106 (N_106,In_159,In_41);
and U107 (N_107,In_209,In_328);
nand U108 (N_108,In_435,In_354);
and U109 (N_109,In_329,In_479);
or U110 (N_110,In_110,In_255);
nor U111 (N_111,In_221,In_340);
nor U112 (N_112,In_185,In_483);
xor U113 (N_113,In_499,In_243);
and U114 (N_114,In_156,In_38);
nor U115 (N_115,In_433,In_78);
nand U116 (N_116,In_323,In_214);
or U117 (N_117,In_485,In_43);
nor U118 (N_118,In_338,In_48);
nand U119 (N_119,In_167,In_182);
nand U120 (N_120,In_374,In_114);
nand U121 (N_121,In_431,In_42);
nor U122 (N_122,In_96,In_97);
nand U123 (N_123,In_350,In_457);
and U124 (N_124,In_303,In_274);
nand U125 (N_125,In_14,In_467);
and U126 (N_126,In_259,In_23);
and U127 (N_127,In_132,In_129);
nand U128 (N_128,In_320,In_220);
and U129 (N_129,In_245,In_13);
or U130 (N_130,In_26,In_166);
xor U131 (N_131,In_463,In_390);
nand U132 (N_132,In_366,In_389);
or U133 (N_133,In_395,In_400);
nand U134 (N_134,In_293,In_22);
and U135 (N_135,In_56,In_127);
and U136 (N_136,In_28,In_456);
and U137 (N_137,In_417,In_469);
or U138 (N_138,In_118,In_461);
nor U139 (N_139,In_286,In_291);
nor U140 (N_140,In_468,In_198);
nand U141 (N_141,In_232,In_162);
nand U142 (N_142,In_487,In_55);
and U143 (N_143,In_365,In_378);
nand U144 (N_144,In_421,In_412);
and U145 (N_145,In_392,In_364);
and U146 (N_146,In_462,In_47);
nand U147 (N_147,In_257,In_380);
and U148 (N_148,In_484,In_113);
and U149 (N_149,In_302,In_386);
and U150 (N_150,In_194,In_333);
nor U151 (N_151,In_325,In_134);
or U152 (N_152,In_17,In_213);
and U153 (N_153,In_180,In_454);
nand U154 (N_154,In_272,In_173);
or U155 (N_155,In_262,In_89);
nor U156 (N_156,In_107,In_379);
nor U157 (N_157,In_388,In_360);
and U158 (N_158,In_356,In_178);
nand U159 (N_159,In_270,In_436);
or U160 (N_160,In_494,In_344);
or U161 (N_161,In_251,In_158);
nand U162 (N_162,In_438,In_451);
nor U163 (N_163,In_349,In_289);
or U164 (N_164,In_152,In_353);
or U165 (N_165,In_136,In_409);
or U166 (N_166,In_91,In_244);
and U167 (N_167,In_104,In_449);
xnor U168 (N_168,In_336,In_116);
or U169 (N_169,In_5,In_216);
xnor U170 (N_170,In_332,In_367);
nor U171 (N_171,In_58,In_369);
and U172 (N_172,In_36,In_307);
or U173 (N_173,In_85,In_403);
xnor U174 (N_174,In_408,In_135);
nand U175 (N_175,In_126,In_310);
nand U176 (N_176,In_482,In_18);
and U177 (N_177,In_225,In_32);
and U178 (N_178,In_423,In_271);
or U179 (N_179,In_206,In_72);
nand U180 (N_180,In_165,In_186);
xor U181 (N_181,In_210,In_54);
xnor U182 (N_182,In_458,In_2);
nand U183 (N_183,In_397,In_419);
and U184 (N_184,In_90,In_294);
nor U185 (N_185,In_298,In_237);
nand U186 (N_186,In_16,In_52);
or U187 (N_187,In_77,In_204);
nand U188 (N_188,In_406,In_45);
and U189 (N_189,In_224,In_183);
or U190 (N_190,In_143,In_188);
nor U191 (N_191,In_306,In_109);
or U192 (N_192,In_174,In_108);
and U193 (N_193,In_195,In_348);
nand U194 (N_194,In_324,In_83);
nand U195 (N_195,In_101,In_249);
nand U196 (N_196,In_287,In_50);
nor U197 (N_197,In_411,In_81);
nand U198 (N_198,In_69,In_279);
xnor U199 (N_199,In_450,In_202);
nand U200 (N_200,In_292,N_108);
nor U201 (N_201,N_85,In_429);
nor U202 (N_202,N_72,In_384);
or U203 (N_203,N_53,In_223);
or U204 (N_204,In_138,N_97);
or U205 (N_205,In_37,N_79);
nor U206 (N_206,N_35,N_188);
or U207 (N_207,In_212,N_127);
nand U208 (N_208,N_187,N_33);
xnor U209 (N_209,N_115,N_95);
and U210 (N_210,N_51,N_167);
or U211 (N_211,In_282,N_26);
and U212 (N_212,N_184,In_401);
nor U213 (N_213,N_34,In_142);
or U214 (N_214,In_280,In_128);
or U215 (N_215,N_68,N_157);
nand U216 (N_216,N_25,N_37);
or U217 (N_217,In_345,N_142);
nor U218 (N_218,N_164,N_10);
and U219 (N_219,In_355,N_102);
or U220 (N_220,N_156,N_165);
nand U221 (N_221,In_238,In_381);
nor U222 (N_222,N_160,In_316);
and U223 (N_223,In_425,N_112);
nand U224 (N_224,N_4,N_135);
and U225 (N_225,In_111,N_128);
and U226 (N_226,N_86,In_200);
xnor U227 (N_227,N_137,N_19);
nand U228 (N_228,In_398,N_11);
and U229 (N_229,N_21,In_260);
or U230 (N_230,N_44,N_100);
or U231 (N_231,N_153,In_358);
nor U232 (N_232,In_455,N_91);
xor U233 (N_233,N_22,N_123);
and U234 (N_234,N_71,N_186);
nand U235 (N_235,N_129,In_153);
nor U236 (N_236,N_40,N_138);
nor U237 (N_237,N_89,In_137);
or U238 (N_238,N_136,In_391);
or U239 (N_239,N_50,N_32);
xnor U240 (N_240,N_119,N_190);
or U241 (N_241,In_34,N_45);
nor U242 (N_242,N_49,In_76);
and U243 (N_243,N_3,N_81);
nor U244 (N_244,N_75,N_146);
or U245 (N_245,N_158,N_57);
and U246 (N_246,N_9,In_318);
xor U247 (N_247,N_192,N_126);
xor U248 (N_248,N_24,N_87);
nand U249 (N_249,In_399,N_139);
and U250 (N_250,N_197,N_17);
nor U251 (N_251,N_177,In_133);
nand U252 (N_252,N_194,N_134);
nand U253 (N_253,N_103,In_71);
xor U254 (N_254,In_154,N_29);
or U255 (N_255,N_198,In_475);
or U256 (N_256,In_169,In_131);
and U257 (N_257,In_474,In_443);
nor U258 (N_258,In_115,N_124);
and U259 (N_259,N_59,In_246);
xnor U260 (N_260,N_18,N_98);
nand U261 (N_261,In_471,N_38);
nand U262 (N_262,N_196,N_155);
xor U263 (N_263,In_146,N_64);
nor U264 (N_264,In_233,N_8);
nand U265 (N_265,N_181,In_215);
nand U266 (N_266,In_322,In_275);
and U267 (N_267,N_141,N_195);
and U268 (N_268,N_27,N_47);
and U269 (N_269,In_489,N_163);
nand U270 (N_270,In_68,In_87);
nand U271 (N_271,N_73,N_122);
nand U272 (N_272,N_109,N_111);
nor U273 (N_273,N_16,In_296);
xor U274 (N_274,N_193,N_179);
and U275 (N_275,N_7,In_331);
nand U276 (N_276,In_263,N_46);
nor U277 (N_277,N_14,N_133);
or U278 (N_278,N_125,In_227);
and U279 (N_279,N_99,In_253);
nor U280 (N_280,N_23,N_183);
and U281 (N_281,In_192,N_28);
or U282 (N_282,N_131,N_105);
nor U283 (N_283,In_203,In_205);
nand U284 (N_284,N_6,N_92);
xor U285 (N_285,N_159,N_117);
or U286 (N_286,N_149,N_185);
nand U287 (N_287,In_385,In_103);
nand U288 (N_288,N_175,N_101);
nand U289 (N_289,N_80,In_496);
nand U290 (N_290,N_106,In_437);
nor U291 (N_291,N_143,N_60);
nor U292 (N_292,N_42,N_116);
nand U293 (N_293,In_147,In_368);
nor U294 (N_294,In_196,N_171);
xnor U295 (N_295,N_173,N_121);
nand U296 (N_296,N_74,N_66);
nand U297 (N_297,N_144,In_226);
nor U298 (N_298,N_36,N_88);
nand U299 (N_299,N_77,N_118);
nand U300 (N_300,N_172,N_189);
nand U301 (N_301,N_162,N_2);
nor U302 (N_302,N_148,N_78);
xnor U303 (N_303,In_278,N_20);
and U304 (N_304,N_120,In_99);
or U305 (N_305,In_459,In_66);
xnor U306 (N_306,In_413,N_147);
and U307 (N_307,In_269,In_27);
nand U308 (N_308,In_231,N_31);
nand U309 (N_309,N_166,N_170);
nand U310 (N_310,In_447,N_113);
or U311 (N_311,N_154,N_130);
or U312 (N_312,In_217,N_12);
and U313 (N_313,N_84,N_94);
nand U314 (N_314,N_182,N_58);
nand U315 (N_315,N_69,N_83);
nand U316 (N_316,N_43,In_252);
and U317 (N_317,N_96,N_5);
nand U318 (N_318,N_178,N_140);
and U319 (N_319,N_76,N_180);
xnor U320 (N_320,In_321,In_285);
and U321 (N_321,N_176,N_55);
xor U322 (N_322,N_132,N_150);
nor U323 (N_323,N_41,In_92);
xor U324 (N_324,N_168,N_82);
nor U325 (N_325,In_334,In_261);
or U326 (N_326,N_1,N_39);
or U327 (N_327,N_107,In_49);
nand U328 (N_328,In_124,N_48);
and U329 (N_329,N_0,In_199);
xnor U330 (N_330,N_30,N_145);
or U331 (N_331,N_54,N_151);
and U332 (N_332,N_114,N_104);
nand U333 (N_333,N_56,N_174);
xor U334 (N_334,N_161,N_93);
xor U335 (N_335,In_86,N_61);
nor U336 (N_336,N_169,In_10);
nand U337 (N_337,N_191,N_13);
nor U338 (N_338,In_155,In_373);
and U339 (N_339,N_65,N_63);
or U340 (N_340,In_371,N_90);
or U341 (N_341,N_15,In_264);
xnor U342 (N_342,In_20,In_176);
and U343 (N_343,In_11,In_9);
and U344 (N_344,In_427,N_62);
nor U345 (N_345,N_199,In_339);
nor U346 (N_346,N_110,N_52);
nor U347 (N_347,In_184,N_152);
or U348 (N_348,In_57,In_297);
or U349 (N_349,N_70,N_67);
nor U350 (N_350,N_159,N_49);
nor U351 (N_351,N_35,N_37);
and U352 (N_352,N_138,N_75);
and U353 (N_353,In_20,N_132);
nand U354 (N_354,N_4,In_413);
nand U355 (N_355,N_8,N_66);
or U356 (N_356,N_106,N_23);
nand U357 (N_357,N_87,N_14);
or U358 (N_358,N_110,N_16);
nand U359 (N_359,In_296,N_160);
nand U360 (N_360,N_129,N_179);
nor U361 (N_361,N_149,N_24);
nand U362 (N_362,N_5,In_133);
or U363 (N_363,N_31,N_57);
nor U364 (N_364,N_66,N_155);
nand U365 (N_365,N_94,N_133);
and U366 (N_366,N_89,N_178);
and U367 (N_367,N_67,In_264);
or U368 (N_368,N_169,N_172);
or U369 (N_369,N_145,N_57);
nand U370 (N_370,In_147,In_459);
nand U371 (N_371,N_168,In_200);
nor U372 (N_372,In_263,In_169);
nor U373 (N_373,N_14,In_399);
and U374 (N_374,N_65,N_34);
and U375 (N_375,N_48,N_35);
xor U376 (N_376,N_132,N_82);
and U377 (N_377,N_185,N_15);
nand U378 (N_378,In_231,N_86);
or U379 (N_379,N_148,N_47);
nor U380 (N_380,N_96,N_180);
nor U381 (N_381,N_68,N_39);
nand U382 (N_382,N_161,N_97);
or U383 (N_383,N_102,N_179);
nor U384 (N_384,In_233,In_205);
and U385 (N_385,N_133,N_167);
nand U386 (N_386,In_321,N_15);
nand U387 (N_387,N_1,In_142);
nand U388 (N_388,N_158,N_128);
and U389 (N_389,In_261,N_85);
nand U390 (N_390,N_81,In_443);
nor U391 (N_391,In_199,In_331);
nor U392 (N_392,N_166,N_71);
and U393 (N_393,N_187,N_101);
nand U394 (N_394,N_44,N_190);
nand U395 (N_395,N_4,N_174);
or U396 (N_396,In_49,In_443);
nor U397 (N_397,N_62,N_78);
nor U398 (N_398,N_105,N_0);
or U399 (N_399,N_147,In_391);
nor U400 (N_400,N_259,N_292);
and U401 (N_401,N_294,N_213);
xor U402 (N_402,N_381,N_327);
and U403 (N_403,N_280,N_312);
xnor U404 (N_404,N_313,N_206);
nand U405 (N_405,N_257,N_375);
nand U406 (N_406,N_270,N_242);
or U407 (N_407,N_384,N_247);
or U408 (N_408,N_216,N_231);
xnor U409 (N_409,N_374,N_237);
or U410 (N_410,N_303,N_387);
or U411 (N_411,N_388,N_396);
or U412 (N_412,N_367,N_202);
nor U413 (N_413,N_272,N_398);
xor U414 (N_414,N_220,N_291);
or U415 (N_415,N_266,N_253);
and U416 (N_416,N_382,N_289);
or U417 (N_417,N_263,N_347);
nor U418 (N_418,N_329,N_271);
or U419 (N_419,N_325,N_223);
nor U420 (N_420,N_261,N_395);
nand U421 (N_421,N_331,N_243);
nand U422 (N_422,N_345,N_298);
xor U423 (N_423,N_355,N_283);
and U424 (N_424,N_248,N_228);
nor U425 (N_425,N_262,N_309);
nor U426 (N_426,N_344,N_318);
nor U427 (N_427,N_336,N_288);
and U428 (N_428,N_350,N_208);
or U429 (N_429,N_249,N_377);
nand U430 (N_430,N_364,N_360);
and U431 (N_431,N_362,N_332);
xor U432 (N_432,N_239,N_225);
nand U433 (N_433,N_222,N_235);
or U434 (N_434,N_392,N_293);
and U435 (N_435,N_229,N_307);
and U436 (N_436,N_393,N_348);
or U437 (N_437,N_258,N_201);
and U438 (N_438,N_390,N_300);
xnor U439 (N_439,N_264,N_366);
and U440 (N_440,N_308,N_246);
and U441 (N_441,N_323,N_321);
or U442 (N_442,N_207,N_351);
nand U443 (N_443,N_317,N_214);
and U444 (N_444,N_273,N_359);
and U445 (N_445,N_341,N_328);
and U446 (N_446,N_363,N_279);
or U447 (N_447,N_334,N_338);
or U448 (N_448,N_267,N_333);
or U449 (N_449,N_352,N_212);
xor U450 (N_450,N_397,N_250);
and U451 (N_451,N_337,N_282);
and U452 (N_452,N_343,N_200);
nor U453 (N_453,N_301,N_302);
or U454 (N_454,N_357,N_369);
nor U455 (N_455,N_217,N_315);
xor U456 (N_456,N_277,N_233);
or U457 (N_457,N_358,N_304);
xor U458 (N_458,N_278,N_286);
xor U459 (N_459,N_274,N_296);
or U460 (N_460,N_346,N_215);
and U461 (N_461,N_339,N_379);
nand U462 (N_462,N_340,N_254);
nor U463 (N_463,N_276,N_324);
nand U464 (N_464,N_373,N_319);
and U465 (N_465,N_256,N_252);
and U466 (N_466,N_349,N_383);
nor U467 (N_467,N_285,N_275);
or U468 (N_468,N_224,N_240);
nand U469 (N_469,N_342,N_260);
and U470 (N_470,N_205,N_320);
xor U471 (N_471,N_389,N_211);
nand U472 (N_472,N_376,N_269);
nand U473 (N_473,N_361,N_297);
and U474 (N_474,N_368,N_219);
nand U475 (N_475,N_265,N_290);
or U476 (N_476,N_230,N_232);
and U477 (N_477,N_221,N_365);
xor U478 (N_478,N_314,N_326);
and U479 (N_479,N_203,N_305);
nand U480 (N_480,N_255,N_226);
and U481 (N_481,N_399,N_284);
or U482 (N_482,N_372,N_281);
nor U483 (N_483,N_204,N_391);
xor U484 (N_484,N_316,N_353);
nand U485 (N_485,N_311,N_218);
nor U486 (N_486,N_371,N_380);
and U487 (N_487,N_306,N_287);
and U488 (N_488,N_378,N_210);
or U489 (N_489,N_251,N_394);
nand U490 (N_490,N_299,N_241);
and U491 (N_491,N_322,N_385);
xnor U492 (N_492,N_245,N_370);
nand U493 (N_493,N_227,N_268);
xor U494 (N_494,N_354,N_386);
xor U495 (N_495,N_234,N_356);
nor U496 (N_496,N_209,N_236);
and U497 (N_497,N_330,N_238);
or U498 (N_498,N_244,N_295);
nand U499 (N_499,N_335,N_310);
nand U500 (N_500,N_348,N_212);
xnor U501 (N_501,N_222,N_266);
or U502 (N_502,N_327,N_293);
nor U503 (N_503,N_276,N_370);
nor U504 (N_504,N_213,N_367);
nor U505 (N_505,N_228,N_354);
nand U506 (N_506,N_385,N_347);
or U507 (N_507,N_306,N_352);
and U508 (N_508,N_247,N_260);
nand U509 (N_509,N_278,N_208);
nand U510 (N_510,N_332,N_219);
or U511 (N_511,N_237,N_345);
nor U512 (N_512,N_204,N_239);
nor U513 (N_513,N_375,N_275);
nand U514 (N_514,N_251,N_302);
xor U515 (N_515,N_397,N_337);
xor U516 (N_516,N_275,N_297);
or U517 (N_517,N_312,N_326);
and U518 (N_518,N_382,N_201);
or U519 (N_519,N_221,N_346);
and U520 (N_520,N_217,N_208);
and U521 (N_521,N_342,N_298);
nand U522 (N_522,N_396,N_260);
nand U523 (N_523,N_311,N_210);
or U524 (N_524,N_321,N_246);
nand U525 (N_525,N_365,N_375);
nand U526 (N_526,N_339,N_229);
nand U527 (N_527,N_224,N_222);
and U528 (N_528,N_368,N_390);
nand U529 (N_529,N_302,N_271);
nand U530 (N_530,N_305,N_362);
nor U531 (N_531,N_395,N_382);
and U532 (N_532,N_363,N_271);
and U533 (N_533,N_235,N_293);
xnor U534 (N_534,N_286,N_213);
xor U535 (N_535,N_395,N_356);
and U536 (N_536,N_279,N_243);
nand U537 (N_537,N_256,N_248);
nor U538 (N_538,N_309,N_295);
or U539 (N_539,N_310,N_208);
nor U540 (N_540,N_377,N_375);
nand U541 (N_541,N_265,N_345);
or U542 (N_542,N_220,N_300);
nand U543 (N_543,N_248,N_324);
or U544 (N_544,N_337,N_213);
xnor U545 (N_545,N_392,N_350);
nor U546 (N_546,N_359,N_228);
nor U547 (N_547,N_241,N_356);
nor U548 (N_548,N_243,N_318);
or U549 (N_549,N_381,N_203);
or U550 (N_550,N_349,N_348);
xnor U551 (N_551,N_234,N_327);
nand U552 (N_552,N_329,N_370);
nand U553 (N_553,N_340,N_202);
or U554 (N_554,N_202,N_378);
or U555 (N_555,N_263,N_326);
nand U556 (N_556,N_367,N_302);
or U557 (N_557,N_264,N_234);
nand U558 (N_558,N_290,N_281);
nor U559 (N_559,N_242,N_210);
nand U560 (N_560,N_265,N_248);
and U561 (N_561,N_244,N_301);
or U562 (N_562,N_254,N_337);
nor U563 (N_563,N_325,N_244);
nor U564 (N_564,N_232,N_366);
and U565 (N_565,N_248,N_253);
or U566 (N_566,N_237,N_325);
nand U567 (N_567,N_321,N_299);
or U568 (N_568,N_301,N_352);
xor U569 (N_569,N_239,N_251);
xor U570 (N_570,N_217,N_316);
xnor U571 (N_571,N_355,N_259);
and U572 (N_572,N_359,N_254);
nor U573 (N_573,N_365,N_207);
or U574 (N_574,N_333,N_332);
or U575 (N_575,N_316,N_336);
nand U576 (N_576,N_275,N_254);
or U577 (N_577,N_373,N_336);
xnor U578 (N_578,N_353,N_277);
nand U579 (N_579,N_249,N_229);
nand U580 (N_580,N_366,N_369);
xnor U581 (N_581,N_290,N_345);
and U582 (N_582,N_270,N_389);
nor U583 (N_583,N_378,N_268);
or U584 (N_584,N_251,N_321);
or U585 (N_585,N_245,N_391);
nand U586 (N_586,N_397,N_365);
nor U587 (N_587,N_229,N_395);
nor U588 (N_588,N_329,N_209);
and U589 (N_589,N_380,N_311);
and U590 (N_590,N_364,N_226);
or U591 (N_591,N_231,N_322);
nand U592 (N_592,N_342,N_303);
or U593 (N_593,N_285,N_335);
or U594 (N_594,N_340,N_292);
xnor U595 (N_595,N_247,N_241);
or U596 (N_596,N_339,N_221);
nand U597 (N_597,N_301,N_280);
xor U598 (N_598,N_343,N_264);
nor U599 (N_599,N_227,N_319);
or U600 (N_600,N_571,N_589);
nand U601 (N_601,N_528,N_419);
and U602 (N_602,N_524,N_514);
xor U603 (N_603,N_443,N_557);
nor U604 (N_604,N_574,N_453);
nor U605 (N_605,N_521,N_568);
nor U606 (N_606,N_486,N_551);
nor U607 (N_607,N_469,N_534);
nand U608 (N_608,N_479,N_455);
nor U609 (N_609,N_492,N_467);
nor U610 (N_610,N_559,N_457);
nor U611 (N_611,N_517,N_530);
nor U612 (N_612,N_561,N_598);
xor U613 (N_613,N_539,N_411);
nand U614 (N_614,N_442,N_424);
nand U615 (N_615,N_407,N_405);
nand U616 (N_616,N_560,N_511);
nor U617 (N_617,N_505,N_416);
and U618 (N_618,N_520,N_435);
nand U619 (N_619,N_414,N_577);
nor U620 (N_620,N_579,N_410);
xor U621 (N_621,N_592,N_531);
and U622 (N_622,N_474,N_438);
or U623 (N_623,N_464,N_554);
and U624 (N_624,N_460,N_458);
or U625 (N_625,N_433,N_509);
nand U626 (N_626,N_562,N_471);
or U627 (N_627,N_498,N_441);
or U628 (N_628,N_515,N_555);
nand U629 (N_629,N_450,N_549);
xor U630 (N_630,N_428,N_525);
or U631 (N_631,N_522,N_501);
nand U632 (N_632,N_432,N_495);
nand U633 (N_633,N_552,N_484);
or U634 (N_634,N_526,N_550);
nor U635 (N_635,N_545,N_527);
nor U636 (N_636,N_566,N_586);
nor U637 (N_637,N_544,N_445);
and U638 (N_638,N_439,N_436);
nor U639 (N_639,N_459,N_476);
or U640 (N_640,N_487,N_535);
nand U641 (N_641,N_409,N_415);
or U642 (N_642,N_567,N_485);
nand U643 (N_643,N_444,N_556);
nand U644 (N_644,N_516,N_538);
nor U645 (N_645,N_596,N_582);
xnor U646 (N_646,N_512,N_456);
or U647 (N_647,N_451,N_565);
and U648 (N_648,N_494,N_518);
nor U649 (N_649,N_401,N_519);
xor U650 (N_650,N_472,N_437);
or U651 (N_651,N_402,N_461);
or U652 (N_652,N_507,N_490);
and U653 (N_653,N_434,N_426);
nor U654 (N_654,N_597,N_452);
nor U655 (N_655,N_481,N_413);
or U656 (N_656,N_580,N_446);
or U657 (N_657,N_475,N_403);
or U658 (N_658,N_422,N_595);
or U659 (N_659,N_513,N_548);
nand U660 (N_660,N_536,N_529);
and U661 (N_661,N_404,N_569);
nand U662 (N_662,N_547,N_496);
nand U663 (N_663,N_502,N_504);
or U664 (N_664,N_425,N_599);
and U665 (N_665,N_482,N_546);
and U666 (N_666,N_454,N_553);
nand U667 (N_667,N_543,N_506);
and U668 (N_668,N_523,N_491);
and U669 (N_669,N_537,N_508);
and U670 (N_670,N_584,N_563);
xor U671 (N_671,N_418,N_542);
xnor U672 (N_672,N_423,N_590);
nand U673 (N_673,N_421,N_427);
or U674 (N_674,N_540,N_499);
or U675 (N_675,N_478,N_408);
nor U676 (N_676,N_429,N_587);
nor U677 (N_677,N_466,N_468);
nor U678 (N_678,N_477,N_572);
nand U679 (N_679,N_575,N_570);
and U680 (N_680,N_510,N_583);
and U681 (N_681,N_480,N_489);
nor U682 (N_682,N_449,N_497);
nand U683 (N_683,N_417,N_493);
or U684 (N_684,N_591,N_412);
or U685 (N_685,N_420,N_448);
nand U686 (N_686,N_576,N_581);
nor U687 (N_687,N_483,N_406);
and U688 (N_688,N_430,N_573);
nor U689 (N_689,N_541,N_578);
or U690 (N_690,N_558,N_440);
and U691 (N_691,N_473,N_532);
nor U692 (N_692,N_533,N_431);
and U693 (N_693,N_447,N_500);
nor U694 (N_694,N_400,N_470);
and U695 (N_695,N_503,N_593);
nand U696 (N_696,N_462,N_588);
nor U697 (N_697,N_594,N_488);
or U698 (N_698,N_465,N_463);
or U699 (N_699,N_564,N_585);
and U700 (N_700,N_482,N_426);
or U701 (N_701,N_455,N_405);
or U702 (N_702,N_450,N_460);
xnor U703 (N_703,N_513,N_545);
nand U704 (N_704,N_404,N_553);
nand U705 (N_705,N_496,N_413);
and U706 (N_706,N_433,N_542);
nor U707 (N_707,N_477,N_475);
nor U708 (N_708,N_463,N_521);
nand U709 (N_709,N_504,N_509);
and U710 (N_710,N_531,N_417);
or U711 (N_711,N_426,N_491);
xnor U712 (N_712,N_534,N_438);
or U713 (N_713,N_400,N_441);
or U714 (N_714,N_594,N_430);
and U715 (N_715,N_487,N_441);
nand U716 (N_716,N_431,N_433);
or U717 (N_717,N_446,N_437);
nand U718 (N_718,N_500,N_544);
nand U719 (N_719,N_446,N_411);
nor U720 (N_720,N_406,N_420);
or U721 (N_721,N_564,N_546);
nand U722 (N_722,N_584,N_509);
and U723 (N_723,N_578,N_471);
nand U724 (N_724,N_562,N_536);
nor U725 (N_725,N_554,N_451);
or U726 (N_726,N_412,N_507);
or U727 (N_727,N_505,N_549);
or U728 (N_728,N_428,N_575);
nor U729 (N_729,N_543,N_487);
and U730 (N_730,N_455,N_410);
and U731 (N_731,N_595,N_488);
or U732 (N_732,N_405,N_449);
and U733 (N_733,N_550,N_453);
or U734 (N_734,N_591,N_527);
nand U735 (N_735,N_523,N_462);
nand U736 (N_736,N_407,N_404);
or U737 (N_737,N_486,N_501);
nand U738 (N_738,N_403,N_507);
nor U739 (N_739,N_587,N_417);
nand U740 (N_740,N_574,N_478);
or U741 (N_741,N_453,N_590);
xor U742 (N_742,N_404,N_585);
nand U743 (N_743,N_524,N_530);
nand U744 (N_744,N_550,N_417);
nor U745 (N_745,N_537,N_488);
and U746 (N_746,N_418,N_584);
nor U747 (N_747,N_541,N_519);
nor U748 (N_748,N_577,N_410);
or U749 (N_749,N_452,N_427);
and U750 (N_750,N_547,N_430);
nor U751 (N_751,N_448,N_557);
and U752 (N_752,N_465,N_492);
nand U753 (N_753,N_440,N_406);
and U754 (N_754,N_448,N_414);
nand U755 (N_755,N_507,N_515);
nand U756 (N_756,N_444,N_501);
and U757 (N_757,N_441,N_472);
nand U758 (N_758,N_492,N_545);
nand U759 (N_759,N_559,N_585);
nand U760 (N_760,N_567,N_449);
nand U761 (N_761,N_463,N_496);
or U762 (N_762,N_595,N_586);
xor U763 (N_763,N_489,N_419);
xnor U764 (N_764,N_411,N_428);
and U765 (N_765,N_412,N_575);
nand U766 (N_766,N_543,N_554);
xnor U767 (N_767,N_498,N_453);
nor U768 (N_768,N_502,N_554);
nand U769 (N_769,N_585,N_529);
or U770 (N_770,N_455,N_548);
nor U771 (N_771,N_433,N_401);
xnor U772 (N_772,N_436,N_528);
and U773 (N_773,N_480,N_477);
nor U774 (N_774,N_402,N_400);
xor U775 (N_775,N_449,N_453);
nand U776 (N_776,N_496,N_472);
nor U777 (N_777,N_410,N_548);
nor U778 (N_778,N_544,N_444);
xnor U779 (N_779,N_518,N_592);
or U780 (N_780,N_518,N_405);
nor U781 (N_781,N_518,N_462);
nor U782 (N_782,N_583,N_588);
or U783 (N_783,N_581,N_502);
and U784 (N_784,N_596,N_541);
or U785 (N_785,N_550,N_565);
nand U786 (N_786,N_512,N_432);
nand U787 (N_787,N_450,N_420);
nand U788 (N_788,N_547,N_442);
and U789 (N_789,N_541,N_567);
nor U790 (N_790,N_471,N_510);
and U791 (N_791,N_536,N_555);
or U792 (N_792,N_434,N_481);
nand U793 (N_793,N_499,N_491);
or U794 (N_794,N_564,N_434);
xor U795 (N_795,N_509,N_488);
or U796 (N_796,N_595,N_558);
nor U797 (N_797,N_494,N_509);
nor U798 (N_798,N_553,N_546);
and U799 (N_799,N_576,N_504);
nand U800 (N_800,N_602,N_738);
or U801 (N_801,N_732,N_664);
or U802 (N_802,N_723,N_780);
and U803 (N_803,N_693,N_613);
nor U804 (N_804,N_646,N_735);
nand U805 (N_805,N_609,N_641);
nor U806 (N_806,N_757,N_619);
xor U807 (N_807,N_783,N_616);
and U808 (N_808,N_617,N_736);
or U809 (N_809,N_796,N_600);
and U810 (N_810,N_795,N_663);
or U811 (N_811,N_784,N_715);
nor U812 (N_812,N_702,N_709);
and U813 (N_813,N_742,N_699);
and U814 (N_814,N_744,N_650);
nor U815 (N_815,N_769,N_770);
or U816 (N_816,N_799,N_618);
nor U817 (N_817,N_666,N_791);
nand U818 (N_818,N_767,N_772);
nor U819 (N_819,N_730,N_703);
xor U820 (N_820,N_675,N_763);
nand U821 (N_821,N_648,N_759);
nand U822 (N_822,N_665,N_718);
xnor U823 (N_823,N_751,N_671);
and U824 (N_824,N_745,N_739);
and U825 (N_825,N_667,N_606);
or U826 (N_826,N_798,N_610);
nor U827 (N_827,N_797,N_728);
nand U828 (N_828,N_614,N_668);
xor U829 (N_829,N_725,N_704);
or U830 (N_830,N_627,N_684);
or U831 (N_831,N_719,N_706);
and U832 (N_832,N_773,N_607);
and U833 (N_833,N_603,N_793);
nor U834 (N_834,N_722,N_752);
nor U835 (N_835,N_724,N_669);
or U836 (N_836,N_695,N_747);
nand U837 (N_837,N_774,N_781);
nand U838 (N_838,N_792,N_685);
nand U839 (N_839,N_676,N_740);
nand U840 (N_840,N_622,N_635);
and U841 (N_841,N_655,N_626);
nor U842 (N_842,N_657,N_687);
and U843 (N_843,N_653,N_758);
nor U844 (N_844,N_660,N_630);
xnor U845 (N_845,N_775,N_678);
nor U846 (N_846,N_682,N_612);
and U847 (N_847,N_681,N_726);
nand U848 (N_848,N_672,N_636);
nor U849 (N_849,N_778,N_605);
nor U850 (N_850,N_696,N_639);
and U851 (N_851,N_679,N_746);
and U852 (N_852,N_727,N_674);
or U853 (N_853,N_683,N_748);
nand U854 (N_854,N_688,N_608);
and U855 (N_855,N_689,N_633);
nand U856 (N_856,N_638,N_777);
and U857 (N_857,N_753,N_714);
nand U858 (N_858,N_720,N_700);
nor U859 (N_859,N_756,N_661);
and U860 (N_860,N_680,N_787);
and U861 (N_861,N_686,N_768);
xor U862 (N_862,N_737,N_765);
nor U863 (N_863,N_734,N_654);
nor U864 (N_864,N_697,N_766);
nand U865 (N_865,N_621,N_623);
nor U866 (N_866,N_649,N_733);
nor U867 (N_867,N_764,N_652);
nor U868 (N_868,N_761,N_624);
xnor U869 (N_869,N_629,N_631);
nor U870 (N_870,N_640,N_637);
and U871 (N_871,N_749,N_755);
or U872 (N_872,N_786,N_673);
or U873 (N_873,N_785,N_771);
and U874 (N_874,N_632,N_754);
xor U875 (N_875,N_794,N_711);
or U876 (N_876,N_628,N_788);
nand U877 (N_877,N_743,N_691);
and U878 (N_878,N_779,N_615);
nand U879 (N_879,N_760,N_662);
nand U880 (N_880,N_634,N_731);
and U881 (N_881,N_611,N_790);
nand U882 (N_882,N_651,N_712);
and U883 (N_883,N_625,N_677);
and U884 (N_884,N_647,N_644);
nand U885 (N_885,N_601,N_789);
and U886 (N_886,N_716,N_645);
and U887 (N_887,N_659,N_698);
nand U888 (N_888,N_762,N_729);
or U889 (N_889,N_620,N_656);
or U890 (N_890,N_705,N_708);
nor U891 (N_891,N_694,N_707);
nor U892 (N_892,N_776,N_643);
and U893 (N_893,N_692,N_710);
or U894 (N_894,N_782,N_604);
and U895 (N_895,N_717,N_713);
nand U896 (N_896,N_670,N_750);
or U897 (N_897,N_701,N_741);
nand U898 (N_898,N_658,N_690);
nor U899 (N_899,N_721,N_642);
and U900 (N_900,N_633,N_680);
and U901 (N_901,N_778,N_752);
and U902 (N_902,N_638,N_793);
nand U903 (N_903,N_798,N_726);
xor U904 (N_904,N_778,N_729);
nor U905 (N_905,N_764,N_785);
nor U906 (N_906,N_644,N_688);
nand U907 (N_907,N_623,N_787);
and U908 (N_908,N_712,N_746);
or U909 (N_909,N_604,N_708);
and U910 (N_910,N_619,N_716);
nand U911 (N_911,N_755,N_605);
nor U912 (N_912,N_782,N_658);
and U913 (N_913,N_720,N_702);
and U914 (N_914,N_664,N_743);
or U915 (N_915,N_778,N_725);
nor U916 (N_916,N_770,N_755);
or U917 (N_917,N_602,N_778);
and U918 (N_918,N_736,N_780);
nand U919 (N_919,N_776,N_634);
or U920 (N_920,N_674,N_751);
or U921 (N_921,N_637,N_711);
nand U922 (N_922,N_693,N_602);
and U923 (N_923,N_677,N_731);
nand U924 (N_924,N_677,N_661);
and U925 (N_925,N_634,N_605);
and U926 (N_926,N_778,N_755);
nand U927 (N_927,N_693,N_691);
nor U928 (N_928,N_712,N_794);
or U929 (N_929,N_780,N_731);
nor U930 (N_930,N_622,N_790);
nor U931 (N_931,N_798,N_785);
nor U932 (N_932,N_723,N_639);
nor U933 (N_933,N_718,N_694);
nand U934 (N_934,N_718,N_755);
or U935 (N_935,N_782,N_620);
xnor U936 (N_936,N_711,N_656);
or U937 (N_937,N_640,N_735);
nor U938 (N_938,N_796,N_706);
xnor U939 (N_939,N_736,N_666);
nand U940 (N_940,N_690,N_630);
nor U941 (N_941,N_786,N_674);
xor U942 (N_942,N_619,N_685);
and U943 (N_943,N_690,N_659);
and U944 (N_944,N_747,N_773);
or U945 (N_945,N_731,N_698);
nor U946 (N_946,N_664,N_620);
nand U947 (N_947,N_686,N_703);
and U948 (N_948,N_608,N_627);
nor U949 (N_949,N_646,N_768);
nor U950 (N_950,N_799,N_681);
nor U951 (N_951,N_706,N_623);
and U952 (N_952,N_613,N_793);
nand U953 (N_953,N_666,N_679);
nand U954 (N_954,N_696,N_626);
nor U955 (N_955,N_633,N_642);
nand U956 (N_956,N_769,N_685);
and U957 (N_957,N_697,N_643);
nor U958 (N_958,N_781,N_645);
nand U959 (N_959,N_649,N_663);
and U960 (N_960,N_661,N_666);
nor U961 (N_961,N_716,N_630);
and U962 (N_962,N_715,N_730);
nor U963 (N_963,N_758,N_705);
nand U964 (N_964,N_755,N_722);
or U965 (N_965,N_764,N_757);
nand U966 (N_966,N_794,N_725);
nand U967 (N_967,N_621,N_730);
nand U968 (N_968,N_633,N_792);
nor U969 (N_969,N_734,N_685);
nor U970 (N_970,N_621,N_681);
nor U971 (N_971,N_655,N_605);
nand U972 (N_972,N_669,N_722);
nand U973 (N_973,N_778,N_662);
xor U974 (N_974,N_760,N_777);
nand U975 (N_975,N_615,N_603);
nand U976 (N_976,N_795,N_781);
xnor U977 (N_977,N_629,N_662);
and U978 (N_978,N_717,N_652);
nor U979 (N_979,N_699,N_730);
and U980 (N_980,N_762,N_645);
nor U981 (N_981,N_716,N_725);
and U982 (N_982,N_760,N_684);
nand U983 (N_983,N_623,N_748);
nand U984 (N_984,N_786,N_639);
nor U985 (N_985,N_678,N_691);
and U986 (N_986,N_777,N_617);
and U987 (N_987,N_791,N_717);
nor U988 (N_988,N_711,N_680);
nand U989 (N_989,N_746,N_748);
and U990 (N_990,N_723,N_647);
nor U991 (N_991,N_683,N_706);
and U992 (N_992,N_782,N_680);
nand U993 (N_993,N_768,N_760);
and U994 (N_994,N_786,N_687);
nor U995 (N_995,N_699,N_799);
nand U996 (N_996,N_694,N_656);
nand U997 (N_997,N_798,N_658);
nand U998 (N_998,N_770,N_723);
xnor U999 (N_999,N_796,N_749);
nor U1000 (N_1000,N_856,N_987);
or U1001 (N_1001,N_909,N_818);
and U1002 (N_1002,N_966,N_915);
nand U1003 (N_1003,N_908,N_984);
or U1004 (N_1004,N_939,N_976);
nor U1005 (N_1005,N_916,N_910);
or U1006 (N_1006,N_982,N_907);
nor U1007 (N_1007,N_924,N_957);
or U1008 (N_1008,N_835,N_829);
xor U1009 (N_1009,N_843,N_825);
nor U1010 (N_1010,N_828,N_935);
xnor U1011 (N_1011,N_881,N_880);
nand U1012 (N_1012,N_855,N_864);
and U1013 (N_1013,N_967,N_807);
or U1014 (N_1014,N_955,N_969);
nor U1015 (N_1015,N_882,N_922);
or U1016 (N_1016,N_863,N_917);
xnor U1017 (N_1017,N_903,N_857);
and U1018 (N_1018,N_932,N_951);
nor U1019 (N_1019,N_943,N_879);
nor U1020 (N_1020,N_896,N_914);
and U1021 (N_1021,N_933,N_980);
and U1022 (N_1022,N_859,N_898);
nor U1023 (N_1023,N_901,N_848);
nand U1024 (N_1024,N_956,N_990);
nand U1025 (N_1025,N_838,N_962);
nor U1026 (N_1026,N_808,N_826);
nor U1027 (N_1027,N_862,N_851);
and U1028 (N_1028,N_830,N_891);
nand U1029 (N_1029,N_888,N_930);
xnor U1030 (N_1030,N_964,N_853);
nor U1031 (N_1031,N_865,N_994);
or U1032 (N_1032,N_997,N_906);
nand U1033 (N_1033,N_827,N_806);
nand U1034 (N_1034,N_961,N_945);
and U1035 (N_1035,N_833,N_873);
or U1036 (N_1036,N_870,N_940);
nor U1037 (N_1037,N_817,N_953);
nand U1038 (N_1038,N_998,N_886);
or U1039 (N_1039,N_876,N_878);
nand U1040 (N_1040,N_804,N_902);
nor U1041 (N_1041,N_931,N_900);
and U1042 (N_1042,N_970,N_959);
nor U1043 (N_1043,N_812,N_847);
xor U1044 (N_1044,N_822,N_958);
nor U1045 (N_1045,N_963,N_872);
and U1046 (N_1046,N_913,N_960);
nor U1047 (N_1047,N_954,N_831);
and U1048 (N_1048,N_911,N_801);
and U1049 (N_1049,N_884,N_895);
nand U1050 (N_1050,N_810,N_978);
and U1051 (N_1051,N_837,N_839);
and U1052 (N_1052,N_854,N_946);
or U1053 (N_1053,N_813,N_952);
nand U1054 (N_1054,N_821,N_925);
nand U1055 (N_1055,N_824,N_819);
or U1056 (N_1056,N_868,N_849);
nor U1057 (N_1057,N_928,N_905);
and U1058 (N_1058,N_832,N_988);
and U1059 (N_1059,N_918,N_845);
or U1060 (N_1060,N_803,N_942);
nor U1061 (N_1061,N_815,N_965);
nand U1062 (N_1062,N_986,N_866);
nor U1063 (N_1063,N_974,N_887);
nand U1064 (N_1064,N_938,N_941);
nand U1065 (N_1065,N_948,N_893);
or U1066 (N_1066,N_936,N_811);
nor U1067 (N_1067,N_972,N_877);
nor U1068 (N_1068,N_890,N_885);
nand U1069 (N_1069,N_937,N_858);
nand U1070 (N_1070,N_844,N_814);
nand U1071 (N_1071,N_971,N_934);
xor U1072 (N_1072,N_991,N_983);
nor U1073 (N_1073,N_929,N_949);
nand U1074 (N_1074,N_993,N_944);
nor U1075 (N_1075,N_985,N_850);
nand U1076 (N_1076,N_897,N_892);
xor U1077 (N_1077,N_950,N_973);
and U1078 (N_1078,N_999,N_823);
nor U1079 (N_1079,N_889,N_947);
and U1080 (N_1080,N_996,N_883);
and U1081 (N_1081,N_920,N_805);
nor U1082 (N_1082,N_979,N_968);
xor U1083 (N_1083,N_904,N_975);
and U1084 (N_1084,N_921,N_981);
and U1085 (N_1085,N_995,N_800);
nor U1086 (N_1086,N_894,N_869);
nand U1087 (N_1087,N_802,N_834);
nor U1088 (N_1088,N_867,N_977);
or U1089 (N_1089,N_899,N_923);
xnor U1090 (N_1090,N_816,N_820);
nand U1091 (N_1091,N_841,N_926);
or U1092 (N_1092,N_860,N_836);
nand U1093 (N_1093,N_861,N_927);
nor U1094 (N_1094,N_874,N_842);
nor U1095 (N_1095,N_809,N_871);
nor U1096 (N_1096,N_912,N_852);
or U1097 (N_1097,N_989,N_919);
or U1098 (N_1098,N_992,N_840);
and U1099 (N_1099,N_846,N_875);
and U1100 (N_1100,N_904,N_963);
nand U1101 (N_1101,N_893,N_917);
or U1102 (N_1102,N_808,N_863);
nor U1103 (N_1103,N_878,N_868);
nand U1104 (N_1104,N_955,N_868);
nor U1105 (N_1105,N_990,N_998);
and U1106 (N_1106,N_819,N_932);
and U1107 (N_1107,N_957,N_955);
nand U1108 (N_1108,N_962,N_980);
nor U1109 (N_1109,N_865,N_853);
or U1110 (N_1110,N_828,N_912);
xnor U1111 (N_1111,N_830,N_814);
nand U1112 (N_1112,N_878,N_993);
or U1113 (N_1113,N_957,N_917);
and U1114 (N_1114,N_923,N_865);
or U1115 (N_1115,N_821,N_967);
nor U1116 (N_1116,N_828,N_976);
nor U1117 (N_1117,N_907,N_911);
nand U1118 (N_1118,N_859,N_936);
and U1119 (N_1119,N_925,N_977);
and U1120 (N_1120,N_942,N_902);
nand U1121 (N_1121,N_899,N_871);
nor U1122 (N_1122,N_905,N_922);
and U1123 (N_1123,N_920,N_934);
nor U1124 (N_1124,N_977,N_909);
nand U1125 (N_1125,N_952,N_862);
or U1126 (N_1126,N_850,N_957);
and U1127 (N_1127,N_887,N_827);
nand U1128 (N_1128,N_860,N_926);
or U1129 (N_1129,N_885,N_981);
nand U1130 (N_1130,N_938,N_922);
nor U1131 (N_1131,N_897,N_993);
nor U1132 (N_1132,N_906,N_888);
and U1133 (N_1133,N_986,N_989);
nor U1134 (N_1134,N_982,N_875);
and U1135 (N_1135,N_949,N_801);
nand U1136 (N_1136,N_844,N_822);
and U1137 (N_1137,N_992,N_943);
and U1138 (N_1138,N_859,N_999);
or U1139 (N_1139,N_809,N_968);
nor U1140 (N_1140,N_992,N_910);
and U1141 (N_1141,N_940,N_923);
xnor U1142 (N_1142,N_958,N_903);
and U1143 (N_1143,N_812,N_916);
xnor U1144 (N_1144,N_969,N_837);
and U1145 (N_1145,N_987,N_943);
or U1146 (N_1146,N_864,N_874);
or U1147 (N_1147,N_876,N_902);
nor U1148 (N_1148,N_946,N_807);
nand U1149 (N_1149,N_905,N_871);
and U1150 (N_1150,N_974,N_854);
or U1151 (N_1151,N_966,N_899);
nor U1152 (N_1152,N_880,N_876);
xor U1153 (N_1153,N_806,N_903);
nand U1154 (N_1154,N_838,N_806);
or U1155 (N_1155,N_995,N_953);
nor U1156 (N_1156,N_924,N_958);
and U1157 (N_1157,N_936,N_984);
xnor U1158 (N_1158,N_851,N_899);
nand U1159 (N_1159,N_873,N_903);
and U1160 (N_1160,N_985,N_919);
nand U1161 (N_1161,N_860,N_846);
xnor U1162 (N_1162,N_817,N_939);
nand U1163 (N_1163,N_973,N_958);
xor U1164 (N_1164,N_902,N_971);
nand U1165 (N_1165,N_809,N_911);
xor U1166 (N_1166,N_891,N_899);
xor U1167 (N_1167,N_852,N_954);
or U1168 (N_1168,N_867,N_801);
nand U1169 (N_1169,N_975,N_933);
and U1170 (N_1170,N_924,N_976);
or U1171 (N_1171,N_867,N_855);
nor U1172 (N_1172,N_809,N_910);
xnor U1173 (N_1173,N_842,N_888);
nand U1174 (N_1174,N_860,N_925);
nor U1175 (N_1175,N_853,N_866);
and U1176 (N_1176,N_861,N_894);
nor U1177 (N_1177,N_948,N_932);
nand U1178 (N_1178,N_831,N_944);
or U1179 (N_1179,N_907,N_868);
nor U1180 (N_1180,N_948,N_973);
nor U1181 (N_1181,N_826,N_804);
nor U1182 (N_1182,N_975,N_819);
nand U1183 (N_1183,N_839,N_990);
and U1184 (N_1184,N_868,N_920);
xnor U1185 (N_1185,N_878,N_952);
nand U1186 (N_1186,N_919,N_835);
and U1187 (N_1187,N_833,N_986);
and U1188 (N_1188,N_935,N_937);
nor U1189 (N_1189,N_878,N_812);
nor U1190 (N_1190,N_893,N_811);
or U1191 (N_1191,N_882,N_997);
or U1192 (N_1192,N_821,N_874);
or U1193 (N_1193,N_883,N_804);
and U1194 (N_1194,N_816,N_879);
nor U1195 (N_1195,N_945,N_833);
and U1196 (N_1196,N_993,N_828);
and U1197 (N_1197,N_976,N_983);
and U1198 (N_1198,N_927,N_964);
or U1199 (N_1199,N_959,N_872);
nand U1200 (N_1200,N_1055,N_1050);
nand U1201 (N_1201,N_1181,N_1195);
nor U1202 (N_1202,N_1089,N_1149);
nand U1203 (N_1203,N_1000,N_1018);
nand U1204 (N_1204,N_1069,N_1124);
xnor U1205 (N_1205,N_1038,N_1015);
or U1206 (N_1206,N_1155,N_1125);
nor U1207 (N_1207,N_1040,N_1074);
and U1208 (N_1208,N_1105,N_1183);
or U1209 (N_1209,N_1029,N_1177);
nand U1210 (N_1210,N_1192,N_1167);
xnor U1211 (N_1211,N_1141,N_1056);
and U1212 (N_1212,N_1073,N_1019);
xnor U1213 (N_1213,N_1198,N_1086);
and U1214 (N_1214,N_1006,N_1174);
nor U1215 (N_1215,N_1163,N_1152);
nand U1216 (N_1216,N_1091,N_1165);
and U1217 (N_1217,N_1159,N_1042);
nor U1218 (N_1218,N_1139,N_1103);
nor U1219 (N_1219,N_1184,N_1083);
nor U1220 (N_1220,N_1122,N_1017);
or U1221 (N_1221,N_1087,N_1063);
and U1222 (N_1222,N_1013,N_1156);
nor U1223 (N_1223,N_1128,N_1021);
or U1224 (N_1224,N_1153,N_1037);
xnor U1225 (N_1225,N_1016,N_1150);
or U1226 (N_1226,N_1060,N_1136);
nor U1227 (N_1227,N_1095,N_1022);
nand U1228 (N_1228,N_1147,N_1170);
xnor U1229 (N_1229,N_1144,N_1048);
nor U1230 (N_1230,N_1140,N_1098);
and U1231 (N_1231,N_1020,N_1109);
nand U1232 (N_1232,N_1187,N_1067);
nor U1233 (N_1233,N_1070,N_1065);
or U1234 (N_1234,N_1045,N_1185);
and U1235 (N_1235,N_1032,N_1189);
or U1236 (N_1236,N_1179,N_1161);
xnor U1237 (N_1237,N_1151,N_1142);
or U1238 (N_1238,N_1009,N_1080);
nand U1239 (N_1239,N_1078,N_1160);
and U1240 (N_1240,N_1137,N_1110);
nand U1241 (N_1241,N_1010,N_1085);
nor U1242 (N_1242,N_1154,N_1053);
xnor U1243 (N_1243,N_1082,N_1025);
nor U1244 (N_1244,N_1043,N_1166);
and U1245 (N_1245,N_1123,N_1148);
or U1246 (N_1246,N_1001,N_1191);
nor U1247 (N_1247,N_1024,N_1115);
nor U1248 (N_1248,N_1090,N_1143);
nor U1249 (N_1249,N_1075,N_1002);
or U1250 (N_1250,N_1196,N_1097);
nor U1251 (N_1251,N_1041,N_1106);
and U1252 (N_1252,N_1004,N_1146);
and U1253 (N_1253,N_1113,N_1101);
xor U1254 (N_1254,N_1118,N_1039);
nand U1255 (N_1255,N_1164,N_1133);
and U1256 (N_1256,N_1061,N_1180);
xor U1257 (N_1257,N_1188,N_1028);
or U1258 (N_1258,N_1052,N_1047);
nand U1259 (N_1259,N_1138,N_1173);
and U1260 (N_1260,N_1054,N_1175);
xnor U1261 (N_1261,N_1072,N_1057);
and U1262 (N_1262,N_1107,N_1007);
nand U1263 (N_1263,N_1099,N_1176);
xor U1264 (N_1264,N_1172,N_1114);
or U1265 (N_1265,N_1135,N_1102);
and U1266 (N_1266,N_1116,N_1117);
and U1267 (N_1267,N_1044,N_1079);
and U1268 (N_1268,N_1076,N_1131);
nand U1269 (N_1269,N_1158,N_1049);
nand U1270 (N_1270,N_1100,N_1186);
and U1271 (N_1271,N_1077,N_1129);
or U1272 (N_1272,N_1157,N_1197);
and U1273 (N_1273,N_1026,N_1121);
nand U1274 (N_1274,N_1168,N_1036);
xor U1275 (N_1275,N_1126,N_1093);
nand U1276 (N_1276,N_1092,N_1062);
or U1277 (N_1277,N_1199,N_1023);
nor U1278 (N_1278,N_1108,N_1120);
nand U1279 (N_1279,N_1068,N_1003);
and U1280 (N_1280,N_1011,N_1132);
nor U1281 (N_1281,N_1030,N_1169);
nor U1282 (N_1282,N_1190,N_1031);
and U1283 (N_1283,N_1008,N_1071);
and U1284 (N_1284,N_1005,N_1058);
nand U1285 (N_1285,N_1193,N_1134);
nor U1286 (N_1286,N_1084,N_1096);
nor U1287 (N_1287,N_1111,N_1104);
xnor U1288 (N_1288,N_1059,N_1127);
nand U1289 (N_1289,N_1094,N_1051);
or U1290 (N_1290,N_1119,N_1033);
xnor U1291 (N_1291,N_1012,N_1027);
nor U1292 (N_1292,N_1035,N_1171);
nand U1293 (N_1293,N_1088,N_1112);
or U1294 (N_1294,N_1034,N_1130);
xnor U1295 (N_1295,N_1162,N_1046);
or U1296 (N_1296,N_1178,N_1081);
nor U1297 (N_1297,N_1145,N_1064);
nor U1298 (N_1298,N_1194,N_1182);
and U1299 (N_1299,N_1066,N_1014);
xor U1300 (N_1300,N_1090,N_1109);
xnor U1301 (N_1301,N_1116,N_1187);
nand U1302 (N_1302,N_1099,N_1051);
nand U1303 (N_1303,N_1101,N_1039);
and U1304 (N_1304,N_1085,N_1025);
nor U1305 (N_1305,N_1142,N_1164);
or U1306 (N_1306,N_1088,N_1001);
and U1307 (N_1307,N_1001,N_1029);
or U1308 (N_1308,N_1098,N_1105);
nand U1309 (N_1309,N_1059,N_1092);
or U1310 (N_1310,N_1087,N_1061);
or U1311 (N_1311,N_1007,N_1178);
and U1312 (N_1312,N_1108,N_1054);
or U1313 (N_1313,N_1063,N_1016);
or U1314 (N_1314,N_1067,N_1130);
xor U1315 (N_1315,N_1139,N_1191);
or U1316 (N_1316,N_1020,N_1116);
nor U1317 (N_1317,N_1133,N_1064);
and U1318 (N_1318,N_1115,N_1105);
nor U1319 (N_1319,N_1113,N_1094);
nor U1320 (N_1320,N_1124,N_1072);
xor U1321 (N_1321,N_1058,N_1002);
nand U1322 (N_1322,N_1056,N_1050);
nor U1323 (N_1323,N_1155,N_1147);
nand U1324 (N_1324,N_1088,N_1012);
nor U1325 (N_1325,N_1051,N_1075);
nor U1326 (N_1326,N_1199,N_1156);
xor U1327 (N_1327,N_1055,N_1152);
or U1328 (N_1328,N_1029,N_1084);
nand U1329 (N_1329,N_1147,N_1027);
nand U1330 (N_1330,N_1018,N_1139);
or U1331 (N_1331,N_1169,N_1111);
nand U1332 (N_1332,N_1157,N_1116);
xnor U1333 (N_1333,N_1077,N_1052);
nor U1334 (N_1334,N_1147,N_1003);
and U1335 (N_1335,N_1101,N_1137);
nand U1336 (N_1336,N_1183,N_1153);
nor U1337 (N_1337,N_1064,N_1053);
nand U1338 (N_1338,N_1003,N_1043);
and U1339 (N_1339,N_1127,N_1130);
nand U1340 (N_1340,N_1100,N_1141);
nand U1341 (N_1341,N_1187,N_1142);
nand U1342 (N_1342,N_1161,N_1166);
nor U1343 (N_1343,N_1062,N_1125);
nand U1344 (N_1344,N_1103,N_1077);
nor U1345 (N_1345,N_1170,N_1036);
or U1346 (N_1346,N_1050,N_1103);
nor U1347 (N_1347,N_1093,N_1027);
or U1348 (N_1348,N_1011,N_1022);
nor U1349 (N_1349,N_1153,N_1027);
nor U1350 (N_1350,N_1128,N_1006);
or U1351 (N_1351,N_1076,N_1129);
and U1352 (N_1352,N_1168,N_1189);
nor U1353 (N_1353,N_1195,N_1042);
nor U1354 (N_1354,N_1026,N_1161);
or U1355 (N_1355,N_1065,N_1002);
or U1356 (N_1356,N_1050,N_1098);
nor U1357 (N_1357,N_1147,N_1097);
nand U1358 (N_1358,N_1041,N_1145);
and U1359 (N_1359,N_1177,N_1158);
nor U1360 (N_1360,N_1052,N_1196);
nand U1361 (N_1361,N_1020,N_1067);
and U1362 (N_1362,N_1123,N_1099);
or U1363 (N_1363,N_1083,N_1149);
and U1364 (N_1364,N_1084,N_1185);
and U1365 (N_1365,N_1053,N_1144);
and U1366 (N_1366,N_1122,N_1049);
and U1367 (N_1367,N_1080,N_1100);
xor U1368 (N_1368,N_1160,N_1147);
nor U1369 (N_1369,N_1011,N_1104);
and U1370 (N_1370,N_1149,N_1026);
nand U1371 (N_1371,N_1027,N_1133);
nor U1372 (N_1372,N_1129,N_1045);
or U1373 (N_1373,N_1053,N_1158);
nand U1374 (N_1374,N_1052,N_1182);
xnor U1375 (N_1375,N_1008,N_1002);
nor U1376 (N_1376,N_1035,N_1148);
or U1377 (N_1377,N_1138,N_1139);
nand U1378 (N_1378,N_1042,N_1150);
nor U1379 (N_1379,N_1199,N_1086);
nand U1380 (N_1380,N_1180,N_1006);
nor U1381 (N_1381,N_1045,N_1197);
nand U1382 (N_1382,N_1092,N_1033);
and U1383 (N_1383,N_1076,N_1088);
or U1384 (N_1384,N_1104,N_1091);
nand U1385 (N_1385,N_1161,N_1128);
and U1386 (N_1386,N_1120,N_1028);
and U1387 (N_1387,N_1088,N_1146);
nor U1388 (N_1388,N_1106,N_1023);
nor U1389 (N_1389,N_1069,N_1136);
or U1390 (N_1390,N_1056,N_1187);
and U1391 (N_1391,N_1058,N_1050);
nor U1392 (N_1392,N_1181,N_1136);
nor U1393 (N_1393,N_1183,N_1127);
or U1394 (N_1394,N_1138,N_1035);
or U1395 (N_1395,N_1099,N_1080);
nand U1396 (N_1396,N_1158,N_1006);
nor U1397 (N_1397,N_1069,N_1153);
nor U1398 (N_1398,N_1086,N_1165);
and U1399 (N_1399,N_1071,N_1114);
nor U1400 (N_1400,N_1325,N_1296);
nor U1401 (N_1401,N_1205,N_1336);
nor U1402 (N_1402,N_1349,N_1230);
and U1403 (N_1403,N_1292,N_1289);
and U1404 (N_1404,N_1209,N_1321);
and U1405 (N_1405,N_1278,N_1342);
nand U1406 (N_1406,N_1246,N_1316);
nand U1407 (N_1407,N_1203,N_1333);
and U1408 (N_1408,N_1396,N_1263);
xor U1409 (N_1409,N_1388,N_1304);
nand U1410 (N_1410,N_1368,N_1354);
or U1411 (N_1411,N_1298,N_1262);
and U1412 (N_1412,N_1233,N_1254);
and U1413 (N_1413,N_1227,N_1282);
and U1414 (N_1414,N_1270,N_1358);
nand U1415 (N_1415,N_1366,N_1361);
and U1416 (N_1416,N_1343,N_1319);
and U1417 (N_1417,N_1335,N_1323);
and U1418 (N_1418,N_1272,N_1211);
nand U1419 (N_1419,N_1344,N_1390);
nand U1420 (N_1420,N_1302,N_1332);
nand U1421 (N_1421,N_1357,N_1317);
nand U1422 (N_1422,N_1347,N_1339);
nor U1423 (N_1423,N_1311,N_1310);
or U1424 (N_1424,N_1277,N_1338);
or U1425 (N_1425,N_1394,N_1223);
or U1426 (N_1426,N_1309,N_1228);
nand U1427 (N_1427,N_1322,N_1269);
or U1428 (N_1428,N_1220,N_1330);
nand U1429 (N_1429,N_1375,N_1285);
or U1430 (N_1430,N_1256,N_1283);
or U1431 (N_1431,N_1363,N_1294);
nand U1432 (N_1432,N_1379,N_1329);
or U1433 (N_1433,N_1260,N_1244);
and U1434 (N_1434,N_1251,N_1257);
or U1435 (N_1435,N_1208,N_1236);
nor U1436 (N_1436,N_1359,N_1350);
nor U1437 (N_1437,N_1393,N_1318);
and U1438 (N_1438,N_1364,N_1307);
or U1439 (N_1439,N_1266,N_1265);
xnor U1440 (N_1440,N_1217,N_1314);
nand U1441 (N_1441,N_1267,N_1389);
xnor U1442 (N_1442,N_1235,N_1242);
xor U1443 (N_1443,N_1232,N_1219);
or U1444 (N_1444,N_1258,N_1261);
nand U1445 (N_1445,N_1312,N_1229);
nand U1446 (N_1446,N_1273,N_1351);
and U1447 (N_1447,N_1313,N_1345);
and U1448 (N_1448,N_1303,N_1249);
or U1449 (N_1449,N_1215,N_1372);
nand U1450 (N_1450,N_1238,N_1290);
nand U1451 (N_1451,N_1240,N_1327);
or U1452 (N_1452,N_1207,N_1381);
nand U1453 (N_1453,N_1218,N_1337);
and U1454 (N_1454,N_1370,N_1324);
nand U1455 (N_1455,N_1280,N_1356);
or U1456 (N_1456,N_1221,N_1248);
and U1457 (N_1457,N_1247,N_1222);
nand U1458 (N_1458,N_1271,N_1206);
or U1459 (N_1459,N_1213,N_1281);
nand U1460 (N_1460,N_1276,N_1395);
nor U1461 (N_1461,N_1387,N_1397);
or U1462 (N_1462,N_1200,N_1340);
and U1463 (N_1463,N_1214,N_1376);
or U1464 (N_1464,N_1224,N_1378);
or U1465 (N_1465,N_1299,N_1315);
and U1466 (N_1466,N_1386,N_1239);
nand U1467 (N_1467,N_1286,N_1301);
nand U1468 (N_1468,N_1353,N_1331);
and U1469 (N_1469,N_1320,N_1399);
nor U1470 (N_1470,N_1392,N_1385);
nor U1471 (N_1471,N_1268,N_1279);
and U1472 (N_1472,N_1346,N_1245);
xor U1473 (N_1473,N_1371,N_1360);
or U1474 (N_1474,N_1306,N_1328);
and U1475 (N_1475,N_1326,N_1398);
nor U1476 (N_1476,N_1380,N_1295);
or U1477 (N_1477,N_1210,N_1300);
xnor U1478 (N_1478,N_1264,N_1255);
nor U1479 (N_1479,N_1391,N_1341);
nor U1480 (N_1480,N_1369,N_1382);
nor U1481 (N_1481,N_1237,N_1383);
xnor U1482 (N_1482,N_1202,N_1259);
nor U1483 (N_1483,N_1204,N_1365);
nor U1484 (N_1484,N_1216,N_1367);
nor U1485 (N_1485,N_1201,N_1291);
xnor U1486 (N_1486,N_1212,N_1274);
and U1487 (N_1487,N_1305,N_1297);
nor U1488 (N_1488,N_1287,N_1377);
nor U1489 (N_1489,N_1231,N_1384);
nor U1490 (N_1490,N_1253,N_1250);
or U1491 (N_1491,N_1288,N_1308);
nand U1492 (N_1492,N_1348,N_1226);
nand U1493 (N_1493,N_1243,N_1334);
nor U1494 (N_1494,N_1252,N_1362);
nand U1495 (N_1495,N_1373,N_1355);
nor U1496 (N_1496,N_1284,N_1225);
or U1497 (N_1497,N_1293,N_1241);
nor U1498 (N_1498,N_1275,N_1374);
nor U1499 (N_1499,N_1234,N_1352);
and U1500 (N_1500,N_1379,N_1303);
or U1501 (N_1501,N_1278,N_1204);
or U1502 (N_1502,N_1252,N_1221);
xnor U1503 (N_1503,N_1288,N_1323);
xor U1504 (N_1504,N_1214,N_1347);
nor U1505 (N_1505,N_1337,N_1254);
xor U1506 (N_1506,N_1327,N_1350);
nor U1507 (N_1507,N_1378,N_1231);
or U1508 (N_1508,N_1235,N_1315);
or U1509 (N_1509,N_1382,N_1322);
nor U1510 (N_1510,N_1283,N_1202);
nor U1511 (N_1511,N_1235,N_1345);
xor U1512 (N_1512,N_1337,N_1234);
and U1513 (N_1513,N_1318,N_1246);
and U1514 (N_1514,N_1209,N_1385);
xnor U1515 (N_1515,N_1270,N_1246);
and U1516 (N_1516,N_1291,N_1324);
and U1517 (N_1517,N_1396,N_1367);
or U1518 (N_1518,N_1395,N_1348);
nor U1519 (N_1519,N_1375,N_1210);
or U1520 (N_1520,N_1384,N_1269);
or U1521 (N_1521,N_1249,N_1287);
and U1522 (N_1522,N_1271,N_1323);
and U1523 (N_1523,N_1258,N_1349);
nand U1524 (N_1524,N_1354,N_1329);
nor U1525 (N_1525,N_1261,N_1220);
nor U1526 (N_1526,N_1322,N_1295);
nand U1527 (N_1527,N_1392,N_1300);
nand U1528 (N_1528,N_1351,N_1260);
and U1529 (N_1529,N_1320,N_1234);
nor U1530 (N_1530,N_1267,N_1224);
nor U1531 (N_1531,N_1204,N_1251);
or U1532 (N_1532,N_1251,N_1302);
or U1533 (N_1533,N_1329,N_1216);
xnor U1534 (N_1534,N_1237,N_1285);
or U1535 (N_1535,N_1351,N_1358);
and U1536 (N_1536,N_1320,N_1308);
nand U1537 (N_1537,N_1248,N_1391);
and U1538 (N_1538,N_1291,N_1295);
nand U1539 (N_1539,N_1336,N_1202);
nand U1540 (N_1540,N_1341,N_1250);
or U1541 (N_1541,N_1241,N_1335);
nand U1542 (N_1542,N_1395,N_1386);
and U1543 (N_1543,N_1390,N_1208);
or U1544 (N_1544,N_1327,N_1311);
or U1545 (N_1545,N_1255,N_1327);
nand U1546 (N_1546,N_1262,N_1283);
xnor U1547 (N_1547,N_1319,N_1239);
and U1548 (N_1548,N_1324,N_1335);
nor U1549 (N_1549,N_1261,N_1222);
or U1550 (N_1550,N_1389,N_1320);
xnor U1551 (N_1551,N_1269,N_1291);
or U1552 (N_1552,N_1225,N_1305);
nor U1553 (N_1553,N_1352,N_1318);
and U1554 (N_1554,N_1378,N_1360);
nor U1555 (N_1555,N_1239,N_1279);
and U1556 (N_1556,N_1269,N_1275);
or U1557 (N_1557,N_1234,N_1339);
nor U1558 (N_1558,N_1392,N_1233);
and U1559 (N_1559,N_1300,N_1274);
and U1560 (N_1560,N_1208,N_1231);
xnor U1561 (N_1561,N_1390,N_1233);
nand U1562 (N_1562,N_1385,N_1273);
nand U1563 (N_1563,N_1252,N_1266);
xor U1564 (N_1564,N_1292,N_1247);
and U1565 (N_1565,N_1394,N_1219);
xnor U1566 (N_1566,N_1222,N_1277);
and U1567 (N_1567,N_1332,N_1357);
or U1568 (N_1568,N_1265,N_1336);
or U1569 (N_1569,N_1380,N_1272);
nor U1570 (N_1570,N_1366,N_1339);
nand U1571 (N_1571,N_1351,N_1241);
nand U1572 (N_1572,N_1206,N_1310);
or U1573 (N_1573,N_1393,N_1308);
xnor U1574 (N_1574,N_1312,N_1302);
xor U1575 (N_1575,N_1331,N_1393);
or U1576 (N_1576,N_1361,N_1398);
xor U1577 (N_1577,N_1239,N_1281);
xnor U1578 (N_1578,N_1312,N_1319);
nand U1579 (N_1579,N_1202,N_1385);
and U1580 (N_1580,N_1307,N_1244);
and U1581 (N_1581,N_1224,N_1262);
or U1582 (N_1582,N_1266,N_1393);
nand U1583 (N_1583,N_1204,N_1240);
nand U1584 (N_1584,N_1323,N_1359);
and U1585 (N_1585,N_1321,N_1203);
or U1586 (N_1586,N_1315,N_1202);
and U1587 (N_1587,N_1201,N_1208);
nand U1588 (N_1588,N_1356,N_1315);
or U1589 (N_1589,N_1326,N_1277);
and U1590 (N_1590,N_1207,N_1225);
nand U1591 (N_1591,N_1389,N_1258);
nand U1592 (N_1592,N_1295,N_1367);
nor U1593 (N_1593,N_1378,N_1239);
and U1594 (N_1594,N_1268,N_1211);
and U1595 (N_1595,N_1293,N_1309);
and U1596 (N_1596,N_1387,N_1355);
nand U1597 (N_1597,N_1209,N_1223);
nor U1598 (N_1598,N_1274,N_1208);
and U1599 (N_1599,N_1305,N_1294);
or U1600 (N_1600,N_1457,N_1567);
nor U1601 (N_1601,N_1566,N_1517);
nand U1602 (N_1602,N_1415,N_1558);
and U1603 (N_1603,N_1447,N_1445);
xnor U1604 (N_1604,N_1568,N_1531);
nor U1605 (N_1605,N_1475,N_1489);
and U1606 (N_1606,N_1564,N_1538);
nand U1607 (N_1607,N_1551,N_1408);
xor U1608 (N_1608,N_1527,N_1453);
nor U1609 (N_1609,N_1591,N_1500);
or U1610 (N_1610,N_1565,N_1523);
nand U1611 (N_1611,N_1425,N_1449);
nor U1612 (N_1612,N_1407,N_1465);
and U1613 (N_1613,N_1477,N_1501);
or U1614 (N_1614,N_1584,N_1481);
xor U1615 (N_1615,N_1588,N_1436);
and U1616 (N_1616,N_1442,N_1418);
xor U1617 (N_1617,N_1556,N_1518);
nor U1618 (N_1618,N_1515,N_1502);
nor U1619 (N_1619,N_1546,N_1536);
nor U1620 (N_1620,N_1578,N_1550);
or U1621 (N_1621,N_1459,N_1456);
or U1622 (N_1622,N_1585,N_1579);
nor U1623 (N_1623,N_1464,N_1530);
and U1624 (N_1624,N_1597,N_1492);
nand U1625 (N_1625,N_1419,N_1431);
xor U1626 (N_1626,N_1504,N_1505);
nand U1627 (N_1627,N_1426,N_1594);
nor U1628 (N_1628,N_1521,N_1469);
or U1629 (N_1629,N_1405,N_1460);
and U1630 (N_1630,N_1577,N_1586);
or U1631 (N_1631,N_1434,N_1554);
nor U1632 (N_1632,N_1541,N_1499);
xor U1633 (N_1633,N_1582,N_1472);
nand U1634 (N_1634,N_1497,N_1439);
nor U1635 (N_1635,N_1486,N_1479);
xnor U1636 (N_1636,N_1543,N_1587);
nor U1637 (N_1637,N_1403,N_1427);
xnor U1638 (N_1638,N_1533,N_1534);
or U1639 (N_1639,N_1462,N_1495);
nor U1640 (N_1640,N_1409,N_1450);
nor U1641 (N_1641,N_1498,N_1448);
or U1642 (N_1642,N_1451,N_1467);
nor U1643 (N_1643,N_1511,N_1411);
nor U1644 (N_1644,N_1414,N_1444);
nor U1645 (N_1645,N_1555,N_1508);
nand U1646 (N_1646,N_1466,N_1574);
and U1647 (N_1647,N_1482,N_1532);
and U1648 (N_1648,N_1510,N_1552);
or U1649 (N_1649,N_1413,N_1443);
and U1650 (N_1650,N_1474,N_1512);
or U1651 (N_1651,N_1598,N_1461);
nor U1652 (N_1652,N_1494,N_1542);
xnor U1653 (N_1653,N_1484,N_1402);
or U1654 (N_1654,N_1522,N_1483);
or U1655 (N_1655,N_1539,N_1463);
and U1656 (N_1656,N_1488,N_1468);
nand U1657 (N_1657,N_1458,N_1599);
nand U1658 (N_1658,N_1452,N_1563);
nand U1659 (N_1659,N_1420,N_1412);
nor U1660 (N_1660,N_1506,N_1592);
or U1661 (N_1661,N_1473,N_1516);
and U1662 (N_1662,N_1548,N_1491);
nand U1663 (N_1663,N_1581,N_1519);
or U1664 (N_1664,N_1576,N_1560);
and U1665 (N_1665,N_1417,N_1524);
and U1666 (N_1666,N_1440,N_1537);
nand U1667 (N_1667,N_1400,N_1476);
nand U1668 (N_1668,N_1593,N_1437);
nand U1669 (N_1669,N_1490,N_1429);
or U1670 (N_1670,N_1583,N_1595);
nand U1671 (N_1671,N_1570,N_1507);
and U1672 (N_1672,N_1545,N_1547);
nor U1673 (N_1673,N_1596,N_1553);
nand U1674 (N_1674,N_1404,N_1493);
nor U1675 (N_1675,N_1513,N_1557);
or U1676 (N_1676,N_1528,N_1422);
or U1677 (N_1677,N_1471,N_1503);
nor U1678 (N_1678,N_1509,N_1485);
and U1679 (N_1679,N_1441,N_1580);
xnor U1680 (N_1680,N_1424,N_1478);
nor U1681 (N_1681,N_1438,N_1589);
xnor U1682 (N_1682,N_1549,N_1435);
nor U1683 (N_1683,N_1446,N_1416);
nand U1684 (N_1684,N_1480,N_1487);
and U1685 (N_1685,N_1562,N_1428);
or U1686 (N_1686,N_1454,N_1496);
or U1687 (N_1687,N_1433,N_1590);
and U1688 (N_1688,N_1526,N_1421);
nor U1689 (N_1689,N_1455,N_1544);
and U1690 (N_1690,N_1561,N_1401);
or U1691 (N_1691,N_1430,N_1571);
xnor U1692 (N_1692,N_1514,N_1423);
xor U1693 (N_1693,N_1529,N_1535);
and U1694 (N_1694,N_1573,N_1520);
and U1695 (N_1695,N_1569,N_1559);
or U1696 (N_1696,N_1432,N_1572);
or U1697 (N_1697,N_1575,N_1470);
nor U1698 (N_1698,N_1540,N_1406);
or U1699 (N_1699,N_1525,N_1410);
nor U1700 (N_1700,N_1530,N_1493);
xnor U1701 (N_1701,N_1493,N_1430);
or U1702 (N_1702,N_1572,N_1499);
or U1703 (N_1703,N_1457,N_1522);
or U1704 (N_1704,N_1483,N_1548);
nor U1705 (N_1705,N_1551,N_1403);
and U1706 (N_1706,N_1497,N_1486);
or U1707 (N_1707,N_1499,N_1437);
or U1708 (N_1708,N_1446,N_1568);
nand U1709 (N_1709,N_1463,N_1585);
xnor U1710 (N_1710,N_1500,N_1516);
and U1711 (N_1711,N_1577,N_1582);
or U1712 (N_1712,N_1579,N_1589);
or U1713 (N_1713,N_1454,N_1415);
xor U1714 (N_1714,N_1465,N_1523);
and U1715 (N_1715,N_1541,N_1422);
nor U1716 (N_1716,N_1460,N_1593);
xnor U1717 (N_1717,N_1576,N_1579);
and U1718 (N_1718,N_1567,N_1585);
or U1719 (N_1719,N_1417,N_1571);
or U1720 (N_1720,N_1443,N_1570);
or U1721 (N_1721,N_1559,N_1469);
and U1722 (N_1722,N_1440,N_1510);
or U1723 (N_1723,N_1492,N_1513);
and U1724 (N_1724,N_1528,N_1526);
nand U1725 (N_1725,N_1592,N_1471);
xor U1726 (N_1726,N_1445,N_1524);
or U1727 (N_1727,N_1449,N_1430);
nand U1728 (N_1728,N_1484,N_1411);
or U1729 (N_1729,N_1439,N_1503);
or U1730 (N_1730,N_1542,N_1502);
nand U1731 (N_1731,N_1534,N_1556);
xor U1732 (N_1732,N_1518,N_1515);
and U1733 (N_1733,N_1456,N_1478);
and U1734 (N_1734,N_1579,N_1429);
nor U1735 (N_1735,N_1420,N_1480);
xnor U1736 (N_1736,N_1495,N_1535);
nand U1737 (N_1737,N_1428,N_1585);
and U1738 (N_1738,N_1447,N_1504);
or U1739 (N_1739,N_1406,N_1408);
nand U1740 (N_1740,N_1500,N_1569);
or U1741 (N_1741,N_1503,N_1431);
and U1742 (N_1742,N_1408,N_1479);
xnor U1743 (N_1743,N_1555,N_1557);
xnor U1744 (N_1744,N_1485,N_1545);
nor U1745 (N_1745,N_1474,N_1461);
or U1746 (N_1746,N_1482,N_1413);
xor U1747 (N_1747,N_1599,N_1580);
xor U1748 (N_1748,N_1576,N_1448);
nor U1749 (N_1749,N_1510,N_1557);
and U1750 (N_1750,N_1574,N_1409);
nand U1751 (N_1751,N_1599,N_1481);
or U1752 (N_1752,N_1535,N_1596);
nand U1753 (N_1753,N_1478,N_1564);
nand U1754 (N_1754,N_1430,N_1543);
nor U1755 (N_1755,N_1434,N_1408);
nor U1756 (N_1756,N_1425,N_1555);
or U1757 (N_1757,N_1451,N_1483);
nor U1758 (N_1758,N_1589,N_1533);
nand U1759 (N_1759,N_1470,N_1432);
nand U1760 (N_1760,N_1501,N_1558);
and U1761 (N_1761,N_1420,N_1548);
nand U1762 (N_1762,N_1485,N_1502);
nand U1763 (N_1763,N_1450,N_1539);
nor U1764 (N_1764,N_1567,N_1575);
and U1765 (N_1765,N_1406,N_1426);
and U1766 (N_1766,N_1584,N_1441);
xor U1767 (N_1767,N_1432,N_1508);
nor U1768 (N_1768,N_1484,N_1584);
nand U1769 (N_1769,N_1500,N_1534);
nor U1770 (N_1770,N_1541,N_1502);
or U1771 (N_1771,N_1520,N_1508);
nand U1772 (N_1772,N_1487,N_1579);
nor U1773 (N_1773,N_1565,N_1508);
nand U1774 (N_1774,N_1431,N_1576);
or U1775 (N_1775,N_1596,N_1444);
nand U1776 (N_1776,N_1437,N_1405);
nand U1777 (N_1777,N_1528,N_1581);
nand U1778 (N_1778,N_1505,N_1539);
and U1779 (N_1779,N_1459,N_1558);
nand U1780 (N_1780,N_1579,N_1438);
xnor U1781 (N_1781,N_1507,N_1458);
or U1782 (N_1782,N_1488,N_1452);
xnor U1783 (N_1783,N_1429,N_1530);
nor U1784 (N_1784,N_1474,N_1523);
or U1785 (N_1785,N_1595,N_1569);
nand U1786 (N_1786,N_1535,N_1579);
and U1787 (N_1787,N_1588,N_1402);
or U1788 (N_1788,N_1586,N_1475);
and U1789 (N_1789,N_1528,N_1513);
and U1790 (N_1790,N_1519,N_1545);
and U1791 (N_1791,N_1480,N_1499);
xnor U1792 (N_1792,N_1598,N_1477);
nand U1793 (N_1793,N_1418,N_1470);
nand U1794 (N_1794,N_1553,N_1514);
xnor U1795 (N_1795,N_1576,N_1532);
and U1796 (N_1796,N_1588,N_1568);
nand U1797 (N_1797,N_1526,N_1565);
xnor U1798 (N_1798,N_1471,N_1452);
nor U1799 (N_1799,N_1575,N_1451);
nor U1800 (N_1800,N_1677,N_1793);
and U1801 (N_1801,N_1712,N_1620);
nor U1802 (N_1802,N_1726,N_1735);
xnor U1803 (N_1803,N_1766,N_1701);
nand U1804 (N_1804,N_1621,N_1676);
or U1805 (N_1805,N_1619,N_1708);
or U1806 (N_1806,N_1670,N_1633);
nand U1807 (N_1807,N_1664,N_1787);
or U1808 (N_1808,N_1660,N_1648);
nor U1809 (N_1809,N_1673,N_1613);
nand U1810 (N_1810,N_1601,N_1703);
nand U1811 (N_1811,N_1602,N_1728);
xnor U1812 (N_1812,N_1763,N_1653);
nor U1813 (N_1813,N_1666,N_1767);
nand U1814 (N_1814,N_1682,N_1744);
nor U1815 (N_1815,N_1651,N_1760);
nor U1816 (N_1816,N_1680,N_1674);
or U1817 (N_1817,N_1699,N_1709);
and U1818 (N_1818,N_1610,N_1698);
xnor U1819 (N_1819,N_1759,N_1671);
or U1820 (N_1820,N_1717,N_1625);
nand U1821 (N_1821,N_1650,N_1719);
or U1822 (N_1822,N_1738,N_1631);
nor U1823 (N_1823,N_1654,N_1771);
xnor U1824 (N_1824,N_1694,N_1706);
and U1825 (N_1825,N_1705,N_1618);
nor U1826 (N_1826,N_1605,N_1757);
and U1827 (N_1827,N_1755,N_1643);
and U1828 (N_1828,N_1634,N_1713);
and U1829 (N_1829,N_1715,N_1740);
nand U1830 (N_1830,N_1749,N_1663);
or U1831 (N_1831,N_1630,N_1737);
nand U1832 (N_1832,N_1781,N_1641);
or U1833 (N_1833,N_1731,N_1796);
nor U1834 (N_1834,N_1734,N_1690);
nand U1835 (N_1835,N_1762,N_1697);
nor U1836 (N_1836,N_1727,N_1606);
nand U1837 (N_1837,N_1730,N_1733);
or U1838 (N_1838,N_1704,N_1675);
nor U1839 (N_1839,N_1732,N_1642);
and U1840 (N_1840,N_1638,N_1722);
nor U1841 (N_1841,N_1747,N_1729);
nand U1842 (N_1842,N_1702,N_1721);
nand U1843 (N_1843,N_1761,N_1799);
nor U1844 (N_1844,N_1668,N_1776);
and U1845 (N_1845,N_1659,N_1775);
or U1846 (N_1846,N_1724,N_1758);
and U1847 (N_1847,N_1783,N_1743);
or U1848 (N_1848,N_1672,N_1644);
nand U1849 (N_1849,N_1750,N_1782);
nor U1850 (N_1850,N_1636,N_1778);
nand U1851 (N_1851,N_1752,N_1617);
nand U1852 (N_1852,N_1628,N_1753);
nor U1853 (N_1853,N_1632,N_1692);
and U1854 (N_1854,N_1718,N_1741);
and U1855 (N_1855,N_1607,N_1689);
nor U1856 (N_1856,N_1754,N_1637);
and U1857 (N_1857,N_1612,N_1695);
nand U1858 (N_1858,N_1794,N_1661);
or U1859 (N_1859,N_1797,N_1795);
and U1860 (N_1860,N_1647,N_1720);
nor U1861 (N_1861,N_1627,N_1700);
or U1862 (N_1862,N_1774,N_1611);
nor U1863 (N_1863,N_1746,N_1624);
nand U1864 (N_1864,N_1745,N_1646);
xor U1865 (N_1865,N_1614,N_1769);
nand U1866 (N_1866,N_1764,N_1678);
xor U1867 (N_1867,N_1652,N_1786);
nand U1868 (N_1868,N_1667,N_1603);
or U1869 (N_1869,N_1645,N_1788);
xnor U1870 (N_1870,N_1725,N_1789);
nand U1871 (N_1871,N_1691,N_1657);
or U1872 (N_1872,N_1655,N_1748);
nor U1873 (N_1873,N_1777,N_1785);
and U1874 (N_1874,N_1669,N_1609);
or U1875 (N_1875,N_1791,N_1790);
nand U1876 (N_1876,N_1792,N_1736);
nand U1877 (N_1877,N_1658,N_1656);
or U1878 (N_1878,N_1649,N_1626);
nor U1879 (N_1879,N_1772,N_1688);
nor U1880 (N_1880,N_1768,N_1770);
and U1881 (N_1881,N_1640,N_1623);
or U1882 (N_1882,N_1716,N_1798);
nand U1883 (N_1883,N_1756,N_1684);
nor U1884 (N_1884,N_1615,N_1665);
xnor U1885 (N_1885,N_1784,N_1685);
nand U1886 (N_1886,N_1707,N_1773);
and U1887 (N_1887,N_1779,N_1608);
and U1888 (N_1888,N_1751,N_1765);
and U1889 (N_1889,N_1686,N_1687);
xnor U1890 (N_1890,N_1681,N_1604);
or U1891 (N_1891,N_1780,N_1693);
and U1892 (N_1892,N_1679,N_1639);
and U1893 (N_1893,N_1662,N_1600);
nand U1894 (N_1894,N_1742,N_1683);
nand U1895 (N_1895,N_1714,N_1696);
or U1896 (N_1896,N_1635,N_1622);
nand U1897 (N_1897,N_1739,N_1629);
and U1898 (N_1898,N_1723,N_1711);
nand U1899 (N_1899,N_1616,N_1710);
nand U1900 (N_1900,N_1680,N_1661);
or U1901 (N_1901,N_1762,N_1736);
or U1902 (N_1902,N_1726,N_1731);
and U1903 (N_1903,N_1791,N_1708);
nor U1904 (N_1904,N_1661,N_1715);
nand U1905 (N_1905,N_1700,N_1755);
and U1906 (N_1906,N_1755,N_1792);
nand U1907 (N_1907,N_1750,N_1699);
or U1908 (N_1908,N_1674,N_1664);
or U1909 (N_1909,N_1639,N_1615);
and U1910 (N_1910,N_1720,N_1768);
nand U1911 (N_1911,N_1639,N_1738);
nand U1912 (N_1912,N_1648,N_1774);
or U1913 (N_1913,N_1723,N_1669);
and U1914 (N_1914,N_1710,N_1728);
nor U1915 (N_1915,N_1701,N_1628);
nor U1916 (N_1916,N_1646,N_1730);
and U1917 (N_1917,N_1705,N_1602);
nand U1918 (N_1918,N_1690,N_1785);
xnor U1919 (N_1919,N_1727,N_1674);
or U1920 (N_1920,N_1601,N_1799);
xnor U1921 (N_1921,N_1657,N_1787);
and U1922 (N_1922,N_1724,N_1775);
nor U1923 (N_1923,N_1668,N_1774);
nor U1924 (N_1924,N_1682,N_1648);
and U1925 (N_1925,N_1701,N_1745);
nor U1926 (N_1926,N_1654,N_1727);
or U1927 (N_1927,N_1668,N_1693);
or U1928 (N_1928,N_1700,N_1732);
and U1929 (N_1929,N_1761,N_1677);
nor U1930 (N_1930,N_1602,N_1781);
or U1931 (N_1931,N_1663,N_1675);
nor U1932 (N_1932,N_1624,N_1649);
and U1933 (N_1933,N_1629,N_1602);
or U1934 (N_1934,N_1639,N_1799);
nand U1935 (N_1935,N_1747,N_1601);
nor U1936 (N_1936,N_1639,N_1749);
xor U1937 (N_1937,N_1638,N_1702);
nand U1938 (N_1938,N_1720,N_1615);
and U1939 (N_1939,N_1748,N_1690);
xnor U1940 (N_1940,N_1789,N_1609);
xor U1941 (N_1941,N_1793,N_1690);
and U1942 (N_1942,N_1752,N_1633);
nand U1943 (N_1943,N_1705,N_1652);
nand U1944 (N_1944,N_1736,N_1636);
nand U1945 (N_1945,N_1743,N_1630);
nand U1946 (N_1946,N_1753,N_1602);
and U1947 (N_1947,N_1658,N_1643);
or U1948 (N_1948,N_1657,N_1668);
nor U1949 (N_1949,N_1723,N_1777);
nand U1950 (N_1950,N_1604,N_1758);
nor U1951 (N_1951,N_1794,N_1636);
or U1952 (N_1952,N_1746,N_1759);
xor U1953 (N_1953,N_1732,N_1622);
nor U1954 (N_1954,N_1776,N_1677);
xor U1955 (N_1955,N_1643,N_1649);
xnor U1956 (N_1956,N_1758,N_1730);
nor U1957 (N_1957,N_1698,N_1622);
or U1958 (N_1958,N_1621,N_1650);
nor U1959 (N_1959,N_1736,N_1626);
nor U1960 (N_1960,N_1613,N_1705);
and U1961 (N_1961,N_1638,N_1723);
nor U1962 (N_1962,N_1670,N_1635);
and U1963 (N_1963,N_1662,N_1681);
or U1964 (N_1964,N_1756,N_1733);
nand U1965 (N_1965,N_1695,N_1681);
and U1966 (N_1966,N_1728,N_1729);
and U1967 (N_1967,N_1725,N_1695);
or U1968 (N_1968,N_1772,N_1753);
and U1969 (N_1969,N_1698,N_1634);
nand U1970 (N_1970,N_1699,N_1719);
nor U1971 (N_1971,N_1638,N_1674);
nand U1972 (N_1972,N_1725,N_1686);
nand U1973 (N_1973,N_1644,N_1799);
or U1974 (N_1974,N_1669,N_1656);
and U1975 (N_1975,N_1648,N_1641);
nand U1976 (N_1976,N_1726,N_1700);
or U1977 (N_1977,N_1616,N_1622);
or U1978 (N_1978,N_1605,N_1781);
nor U1979 (N_1979,N_1617,N_1673);
or U1980 (N_1980,N_1679,N_1604);
or U1981 (N_1981,N_1799,N_1716);
xor U1982 (N_1982,N_1748,N_1722);
nand U1983 (N_1983,N_1787,N_1610);
nor U1984 (N_1984,N_1745,N_1601);
xor U1985 (N_1985,N_1634,N_1613);
nand U1986 (N_1986,N_1625,N_1603);
nand U1987 (N_1987,N_1770,N_1694);
or U1988 (N_1988,N_1728,N_1650);
xnor U1989 (N_1989,N_1752,N_1737);
nor U1990 (N_1990,N_1756,N_1649);
xnor U1991 (N_1991,N_1666,N_1717);
and U1992 (N_1992,N_1770,N_1744);
nor U1993 (N_1993,N_1608,N_1750);
and U1994 (N_1994,N_1655,N_1754);
nand U1995 (N_1995,N_1685,N_1729);
and U1996 (N_1996,N_1771,N_1659);
or U1997 (N_1997,N_1655,N_1665);
nor U1998 (N_1998,N_1646,N_1760);
nand U1999 (N_1999,N_1674,N_1791);
nand U2000 (N_2000,N_1816,N_1916);
xnor U2001 (N_2001,N_1886,N_1964);
nor U2002 (N_2002,N_1919,N_1823);
or U2003 (N_2003,N_1857,N_1882);
or U2004 (N_2004,N_1880,N_1972);
or U2005 (N_2005,N_1856,N_1812);
and U2006 (N_2006,N_1832,N_1965);
nor U2007 (N_2007,N_1883,N_1879);
nor U2008 (N_2008,N_1997,N_1830);
and U2009 (N_2009,N_1860,N_1910);
xnor U2010 (N_2010,N_1822,N_1989);
or U2011 (N_2011,N_1953,N_1956);
nand U2012 (N_2012,N_1825,N_1975);
nor U2013 (N_2013,N_1990,N_1954);
and U2014 (N_2014,N_1834,N_1870);
and U2015 (N_2015,N_1839,N_1831);
or U2016 (N_2016,N_1889,N_1957);
nor U2017 (N_2017,N_1829,N_1846);
and U2018 (N_2018,N_1898,N_1927);
nor U2019 (N_2019,N_1915,N_1895);
nand U2020 (N_2020,N_1819,N_1904);
nand U2021 (N_2021,N_1917,N_1960);
nand U2022 (N_2022,N_1841,N_1948);
xor U2023 (N_2023,N_1867,N_1902);
nand U2024 (N_2024,N_1912,N_1827);
and U2025 (N_2025,N_1852,N_1801);
or U2026 (N_2026,N_1980,N_1963);
nor U2027 (N_2027,N_1973,N_1878);
and U2028 (N_2028,N_1942,N_1875);
nor U2029 (N_2029,N_1851,N_1946);
nand U2030 (N_2030,N_1890,N_1808);
nand U2031 (N_2031,N_1842,N_1970);
xor U2032 (N_2032,N_1961,N_1920);
or U2033 (N_2033,N_1874,N_1992);
nand U2034 (N_2034,N_1840,N_1907);
and U2035 (N_2035,N_1873,N_1941);
nor U2036 (N_2036,N_1893,N_1810);
and U2037 (N_2037,N_1943,N_1858);
and U2038 (N_2038,N_1971,N_1921);
nand U2039 (N_2039,N_1894,N_1807);
or U2040 (N_2040,N_1968,N_1996);
nand U2041 (N_2041,N_1981,N_1962);
nand U2042 (N_2042,N_1911,N_1803);
and U2043 (N_2043,N_1924,N_1897);
nand U2044 (N_2044,N_1855,N_1872);
nor U2045 (N_2045,N_1844,N_1861);
xnor U2046 (N_2046,N_1887,N_1929);
and U2047 (N_2047,N_1982,N_1836);
or U2048 (N_2048,N_1955,N_1853);
or U2049 (N_2049,N_1939,N_1802);
or U2050 (N_2050,N_1966,N_1938);
and U2051 (N_2051,N_1935,N_1926);
nor U2052 (N_2052,N_1848,N_1871);
nor U2053 (N_2053,N_1993,N_1945);
nor U2054 (N_2054,N_1985,N_1837);
nor U2055 (N_2055,N_1923,N_1815);
or U2056 (N_2056,N_1959,N_1913);
or U2057 (N_2057,N_1940,N_1811);
xnor U2058 (N_2058,N_1978,N_1928);
nor U2059 (N_2059,N_1958,N_1925);
xnor U2060 (N_2060,N_1849,N_1826);
or U2061 (N_2061,N_1877,N_1865);
nor U2062 (N_2062,N_1933,N_1833);
nor U2063 (N_2063,N_1999,N_1864);
nand U2064 (N_2064,N_1896,N_1901);
nor U2065 (N_2065,N_1906,N_1850);
nor U2066 (N_2066,N_1914,N_1814);
and U2067 (N_2067,N_1828,N_1838);
or U2068 (N_2068,N_1888,N_1909);
nor U2069 (N_2069,N_1800,N_1951);
or U2070 (N_2070,N_1949,N_1932);
nor U2071 (N_2071,N_1847,N_1986);
nand U2072 (N_2072,N_1854,N_1995);
and U2073 (N_2073,N_1922,N_1862);
nand U2074 (N_2074,N_1843,N_1863);
nor U2075 (N_2075,N_1821,N_1845);
nand U2076 (N_2076,N_1930,N_1891);
nand U2077 (N_2077,N_1869,N_1952);
nand U2078 (N_2078,N_1818,N_1892);
or U2079 (N_2079,N_1820,N_1977);
nor U2080 (N_2080,N_1866,N_1969);
or U2081 (N_2081,N_1813,N_1900);
nor U2082 (N_2082,N_1947,N_1974);
or U2083 (N_2083,N_1988,N_1806);
or U2084 (N_2084,N_1998,N_1984);
and U2085 (N_2085,N_1983,N_1835);
nor U2086 (N_2086,N_1868,N_1885);
nand U2087 (N_2087,N_1908,N_1824);
or U2088 (N_2088,N_1987,N_1967);
or U2089 (N_2089,N_1976,N_1979);
and U2090 (N_2090,N_1817,N_1918);
or U2091 (N_2091,N_1881,N_1884);
nand U2092 (N_2092,N_1876,N_1804);
or U2093 (N_2093,N_1905,N_1937);
nand U2094 (N_2094,N_1991,N_1931);
or U2095 (N_2095,N_1805,N_1899);
nand U2096 (N_2096,N_1950,N_1994);
xor U2097 (N_2097,N_1934,N_1809);
nor U2098 (N_2098,N_1859,N_1936);
nor U2099 (N_2099,N_1944,N_1903);
and U2100 (N_2100,N_1854,N_1916);
or U2101 (N_2101,N_1891,N_1971);
and U2102 (N_2102,N_1974,N_1805);
nand U2103 (N_2103,N_1896,N_1847);
nand U2104 (N_2104,N_1939,N_1846);
xor U2105 (N_2105,N_1881,N_1838);
or U2106 (N_2106,N_1953,N_1959);
nor U2107 (N_2107,N_1994,N_1914);
or U2108 (N_2108,N_1830,N_1802);
or U2109 (N_2109,N_1983,N_1988);
nor U2110 (N_2110,N_1862,N_1806);
xor U2111 (N_2111,N_1954,N_1835);
and U2112 (N_2112,N_1902,N_1947);
and U2113 (N_2113,N_1925,N_1913);
or U2114 (N_2114,N_1955,N_1923);
nor U2115 (N_2115,N_1895,N_1809);
nand U2116 (N_2116,N_1815,N_1901);
nand U2117 (N_2117,N_1955,N_1846);
nand U2118 (N_2118,N_1998,N_1836);
or U2119 (N_2119,N_1829,N_1876);
and U2120 (N_2120,N_1913,N_1985);
and U2121 (N_2121,N_1990,N_1968);
or U2122 (N_2122,N_1898,N_1957);
and U2123 (N_2123,N_1922,N_1828);
nand U2124 (N_2124,N_1930,N_1850);
nand U2125 (N_2125,N_1816,N_1875);
and U2126 (N_2126,N_1882,N_1803);
or U2127 (N_2127,N_1922,N_1952);
and U2128 (N_2128,N_1971,N_1937);
and U2129 (N_2129,N_1904,N_1860);
nor U2130 (N_2130,N_1856,N_1875);
or U2131 (N_2131,N_1923,N_1855);
or U2132 (N_2132,N_1998,N_1833);
nor U2133 (N_2133,N_1853,N_1856);
and U2134 (N_2134,N_1811,N_1957);
nor U2135 (N_2135,N_1999,N_1949);
nand U2136 (N_2136,N_1927,N_1971);
xnor U2137 (N_2137,N_1887,N_1955);
or U2138 (N_2138,N_1835,N_1865);
nor U2139 (N_2139,N_1952,N_1955);
and U2140 (N_2140,N_1952,N_1991);
nand U2141 (N_2141,N_1870,N_1925);
xnor U2142 (N_2142,N_1837,N_1905);
or U2143 (N_2143,N_1994,N_1835);
and U2144 (N_2144,N_1806,N_1986);
xor U2145 (N_2145,N_1950,N_1915);
nor U2146 (N_2146,N_1950,N_1948);
or U2147 (N_2147,N_1985,N_1815);
or U2148 (N_2148,N_1916,N_1800);
or U2149 (N_2149,N_1812,N_1908);
nand U2150 (N_2150,N_1890,N_1868);
nand U2151 (N_2151,N_1875,N_1973);
or U2152 (N_2152,N_1931,N_1805);
and U2153 (N_2153,N_1829,N_1857);
or U2154 (N_2154,N_1860,N_1923);
or U2155 (N_2155,N_1869,N_1803);
nand U2156 (N_2156,N_1881,N_1849);
nor U2157 (N_2157,N_1840,N_1896);
and U2158 (N_2158,N_1970,N_1908);
xnor U2159 (N_2159,N_1838,N_1965);
nand U2160 (N_2160,N_1878,N_1866);
nand U2161 (N_2161,N_1882,N_1868);
and U2162 (N_2162,N_1938,N_1988);
and U2163 (N_2163,N_1918,N_1973);
or U2164 (N_2164,N_1955,N_1905);
nand U2165 (N_2165,N_1864,N_1889);
and U2166 (N_2166,N_1875,N_1981);
and U2167 (N_2167,N_1971,N_1874);
nand U2168 (N_2168,N_1803,N_1969);
xor U2169 (N_2169,N_1817,N_1901);
nor U2170 (N_2170,N_1804,N_1844);
xnor U2171 (N_2171,N_1940,N_1874);
xnor U2172 (N_2172,N_1979,N_1929);
nand U2173 (N_2173,N_1883,N_1984);
and U2174 (N_2174,N_1807,N_1844);
nand U2175 (N_2175,N_1894,N_1972);
nor U2176 (N_2176,N_1980,N_1984);
xor U2177 (N_2177,N_1841,N_1960);
or U2178 (N_2178,N_1849,N_1965);
nor U2179 (N_2179,N_1856,N_1840);
and U2180 (N_2180,N_1984,N_1938);
nand U2181 (N_2181,N_1845,N_1960);
nand U2182 (N_2182,N_1896,N_1971);
nor U2183 (N_2183,N_1871,N_1842);
nor U2184 (N_2184,N_1973,N_1936);
or U2185 (N_2185,N_1892,N_1820);
xor U2186 (N_2186,N_1854,N_1861);
and U2187 (N_2187,N_1802,N_1999);
nand U2188 (N_2188,N_1999,N_1848);
xor U2189 (N_2189,N_1982,N_1988);
and U2190 (N_2190,N_1998,N_1814);
nand U2191 (N_2191,N_1849,N_1948);
nor U2192 (N_2192,N_1870,N_1942);
nand U2193 (N_2193,N_1803,N_1991);
nor U2194 (N_2194,N_1888,N_1916);
nor U2195 (N_2195,N_1900,N_1950);
or U2196 (N_2196,N_1843,N_1865);
or U2197 (N_2197,N_1921,N_1840);
and U2198 (N_2198,N_1882,N_1861);
or U2199 (N_2199,N_1865,N_1887);
and U2200 (N_2200,N_2174,N_2101);
nor U2201 (N_2201,N_2183,N_2052);
xor U2202 (N_2202,N_2188,N_2000);
nor U2203 (N_2203,N_2193,N_2049);
nand U2204 (N_2204,N_2152,N_2067);
nand U2205 (N_2205,N_2068,N_2001);
nand U2206 (N_2206,N_2189,N_2180);
nor U2207 (N_2207,N_2177,N_2140);
or U2208 (N_2208,N_2121,N_2036);
nor U2209 (N_2209,N_2047,N_2161);
nand U2210 (N_2210,N_2061,N_2113);
nor U2211 (N_2211,N_2195,N_2029);
xor U2212 (N_2212,N_2099,N_2066);
and U2213 (N_2213,N_2042,N_2055);
or U2214 (N_2214,N_2133,N_2185);
nor U2215 (N_2215,N_2178,N_2154);
and U2216 (N_2216,N_2004,N_2169);
nand U2217 (N_2217,N_2132,N_2163);
nor U2218 (N_2218,N_2083,N_2059);
nor U2219 (N_2219,N_2127,N_2142);
xor U2220 (N_2220,N_2153,N_2119);
or U2221 (N_2221,N_2072,N_2198);
and U2222 (N_2222,N_2139,N_2071);
and U2223 (N_2223,N_2184,N_2038);
nand U2224 (N_2224,N_2176,N_2135);
or U2225 (N_2225,N_2013,N_2051);
nor U2226 (N_2226,N_2079,N_2024);
and U2227 (N_2227,N_2171,N_2023);
xnor U2228 (N_2228,N_2063,N_2073);
nor U2229 (N_2229,N_2090,N_2111);
nor U2230 (N_2230,N_2157,N_2081);
or U2231 (N_2231,N_2043,N_2026);
nor U2232 (N_2232,N_2158,N_2129);
xnor U2233 (N_2233,N_2074,N_2010);
nand U2234 (N_2234,N_2164,N_2143);
nand U2235 (N_2235,N_2002,N_2065);
and U2236 (N_2236,N_2162,N_2062);
nor U2237 (N_2237,N_2109,N_2092);
nor U2238 (N_2238,N_2018,N_2098);
xnor U2239 (N_2239,N_2091,N_2034);
and U2240 (N_2240,N_2033,N_2182);
or U2241 (N_2241,N_2147,N_2089);
or U2242 (N_2242,N_2041,N_2100);
or U2243 (N_2243,N_2136,N_2032);
or U2244 (N_2244,N_2012,N_2076);
nand U2245 (N_2245,N_2186,N_2145);
xor U2246 (N_2246,N_2197,N_2087);
nor U2247 (N_2247,N_2137,N_2181);
xor U2248 (N_2248,N_2194,N_2120);
nand U2249 (N_2249,N_2116,N_2156);
nand U2250 (N_2250,N_2011,N_2144);
nand U2251 (N_2251,N_2126,N_2115);
and U2252 (N_2252,N_2085,N_2103);
nor U2253 (N_2253,N_2117,N_2007);
nor U2254 (N_2254,N_2016,N_2020);
and U2255 (N_2255,N_2187,N_2168);
nand U2256 (N_2256,N_2138,N_2053);
nand U2257 (N_2257,N_2070,N_2075);
xnor U2258 (N_2258,N_2050,N_2096);
xor U2259 (N_2259,N_2167,N_2095);
nand U2260 (N_2260,N_2112,N_2106);
nand U2261 (N_2261,N_2009,N_2166);
xnor U2262 (N_2262,N_2003,N_2035);
nand U2263 (N_2263,N_2077,N_2086);
xor U2264 (N_2264,N_2199,N_2039);
and U2265 (N_2265,N_2110,N_2040);
xor U2266 (N_2266,N_2118,N_2125);
nand U2267 (N_2267,N_2141,N_2123);
or U2268 (N_2268,N_2082,N_2015);
nand U2269 (N_2269,N_2021,N_2030);
nand U2270 (N_2270,N_2192,N_2064);
and U2271 (N_2271,N_2150,N_2102);
nand U2272 (N_2272,N_2108,N_2148);
nor U2273 (N_2273,N_2160,N_2037);
nand U2274 (N_2274,N_2069,N_2093);
nand U2275 (N_2275,N_2155,N_2149);
nor U2276 (N_2276,N_2172,N_2190);
nand U2277 (N_2277,N_2122,N_2008);
nand U2278 (N_2278,N_2107,N_2173);
nor U2279 (N_2279,N_2165,N_2019);
or U2280 (N_2280,N_2058,N_2151);
xor U2281 (N_2281,N_2078,N_2159);
and U2282 (N_2282,N_2027,N_2105);
nand U2283 (N_2283,N_2080,N_2031);
nor U2284 (N_2284,N_2088,N_2006);
nand U2285 (N_2285,N_2046,N_2170);
or U2286 (N_2286,N_2114,N_2104);
or U2287 (N_2287,N_2060,N_2025);
nand U2288 (N_2288,N_2054,N_2094);
and U2289 (N_2289,N_2134,N_2175);
nand U2290 (N_2290,N_2196,N_2044);
and U2291 (N_2291,N_2179,N_2057);
or U2292 (N_2292,N_2048,N_2014);
and U2293 (N_2293,N_2084,N_2146);
or U2294 (N_2294,N_2191,N_2028);
or U2295 (N_2295,N_2017,N_2045);
xor U2296 (N_2296,N_2130,N_2097);
nand U2297 (N_2297,N_2131,N_2124);
and U2298 (N_2298,N_2128,N_2005);
nor U2299 (N_2299,N_2022,N_2056);
and U2300 (N_2300,N_2187,N_2072);
and U2301 (N_2301,N_2155,N_2164);
and U2302 (N_2302,N_2046,N_2045);
nand U2303 (N_2303,N_2113,N_2041);
or U2304 (N_2304,N_2147,N_2084);
nor U2305 (N_2305,N_2081,N_2089);
nor U2306 (N_2306,N_2003,N_2049);
nor U2307 (N_2307,N_2132,N_2031);
and U2308 (N_2308,N_2023,N_2043);
nor U2309 (N_2309,N_2140,N_2183);
or U2310 (N_2310,N_2199,N_2063);
xor U2311 (N_2311,N_2106,N_2160);
and U2312 (N_2312,N_2142,N_2086);
nor U2313 (N_2313,N_2030,N_2194);
nand U2314 (N_2314,N_2000,N_2091);
and U2315 (N_2315,N_2150,N_2196);
or U2316 (N_2316,N_2163,N_2012);
or U2317 (N_2317,N_2177,N_2016);
and U2318 (N_2318,N_2157,N_2079);
nand U2319 (N_2319,N_2056,N_2072);
and U2320 (N_2320,N_2028,N_2110);
and U2321 (N_2321,N_2105,N_2021);
nand U2322 (N_2322,N_2025,N_2115);
xnor U2323 (N_2323,N_2152,N_2142);
nor U2324 (N_2324,N_2040,N_2070);
nor U2325 (N_2325,N_2042,N_2093);
xnor U2326 (N_2326,N_2055,N_2064);
and U2327 (N_2327,N_2004,N_2052);
nand U2328 (N_2328,N_2172,N_2132);
or U2329 (N_2329,N_2181,N_2174);
nor U2330 (N_2330,N_2145,N_2069);
or U2331 (N_2331,N_2049,N_2116);
and U2332 (N_2332,N_2175,N_2136);
nor U2333 (N_2333,N_2142,N_2023);
or U2334 (N_2334,N_2128,N_2114);
nand U2335 (N_2335,N_2119,N_2095);
nand U2336 (N_2336,N_2055,N_2184);
or U2337 (N_2337,N_2095,N_2172);
or U2338 (N_2338,N_2087,N_2167);
or U2339 (N_2339,N_2065,N_2023);
nor U2340 (N_2340,N_2125,N_2003);
xnor U2341 (N_2341,N_2122,N_2191);
nand U2342 (N_2342,N_2147,N_2144);
or U2343 (N_2343,N_2041,N_2045);
or U2344 (N_2344,N_2059,N_2119);
or U2345 (N_2345,N_2190,N_2126);
nor U2346 (N_2346,N_2087,N_2000);
and U2347 (N_2347,N_2108,N_2004);
nor U2348 (N_2348,N_2064,N_2103);
or U2349 (N_2349,N_2065,N_2108);
and U2350 (N_2350,N_2176,N_2076);
or U2351 (N_2351,N_2032,N_2040);
or U2352 (N_2352,N_2035,N_2056);
nand U2353 (N_2353,N_2147,N_2116);
nor U2354 (N_2354,N_2189,N_2125);
nor U2355 (N_2355,N_2008,N_2129);
nor U2356 (N_2356,N_2114,N_2068);
nor U2357 (N_2357,N_2099,N_2166);
or U2358 (N_2358,N_2136,N_2171);
or U2359 (N_2359,N_2102,N_2067);
or U2360 (N_2360,N_2049,N_2013);
nand U2361 (N_2361,N_2004,N_2149);
nor U2362 (N_2362,N_2112,N_2187);
nor U2363 (N_2363,N_2115,N_2039);
nor U2364 (N_2364,N_2047,N_2068);
and U2365 (N_2365,N_2196,N_2190);
nor U2366 (N_2366,N_2005,N_2072);
nand U2367 (N_2367,N_2113,N_2131);
nor U2368 (N_2368,N_2004,N_2000);
and U2369 (N_2369,N_2120,N_2028);
nor U2370 (N_2370,N_2058,N_2188);
and U2371 (N_2371,N_2059,N_2193);
or U2372 (N_2372,N_2176,N_2098);
or U2373 (N_2373,N_2020,N_2194);
or U2374 (N_2374,N_2197,N_2190);
nand U2375 (N_2375,N_2158,N_2194);
and U2376 (N_2376,N_2193,N_2024);
or U2377 (N_2377,N_2175,N_2053);
xor U2378 (N_2378,N_2107,N_2017);
nand U2379 (N_2379,N_2028,N_2157);
nand U2380 (N_2380,N_2033,N_2065);
and U2381 (N_2381,N_2165,N_2057);
nand U2382 (N_2382,N_2149,N_2064);
and U2383 (N_2383,N_2153,N_2148);
and U2384 (N_2384,N_2184,N_2185);
and U2385 (N_2385,N_2067,N_2107);
nand U2386 (N_2386,N_2054,N_2097);
nand U2387 (N_2387,N_2090,N_2097);
or U2388 (N_2388,N_2009,N_2125);
nand U2389 (N_2389,N_2097,N_2030);
nor U2390 (N_2390,N_2083,N_2099);
xor U2391 (N_2391,N_2003,N_2101);
nor U2392 (N_2392,N_2088,N_2055);
xor U2393 (N_2393,N_2174,N_2104);
nand U2394 (N_2394,N_2089,N_2159);
and U2395 (N_2395,N_2026,N_2170);
and U2396 (N_2396,N_2078,N_2135);
and U2397 (N_2397,N_2017,N_2042);
and U2398 (N_2398,N_2128,N_2198);
nand U2399 (N_2399,N_2024,N_2078);
nor U2400 (N_2400,N_2386,N_2262);
nor U2401 (N_2401,N_2297,N_2361);
xor U2402 (N_2402,N_2318,N_2391);
or U2403 (N_2403,N_2239,N_2285);
or U2404 (N_2404,N_2338,N_2368);
nor U2405 (N_2405,N_2237,N_2217);
nand U2406 (N_2406,N_2218,N_2380);
xnor U2407 (N_2407,N_2290,N_2332);
nor U2408 (N_2408,N_2291,N_2273);
nor U2409 (N_2409,N_2261,N_2233);
and U2410 (N_2410,N_2203,N_2214);
nor U2411 (N_2411,N_2309,N_2231);
or U2412 (N_2412,N_2207,N_2326);
nand U2413 (N_2413,N_2349,N_2255);
nand U2414 (N_2414,N_2346,N_2335);
and U2415 (N_2415,N_2360,N_2362);
nand U2416 (N_2416,N_2256,N_2305);
nor U2417 (N_2417,N_2209,N_2234);
or U2418 (N_2418,N_2287,N_2222);
or U2419 (N_2419,N_2320,N_2369);
or U2420 (N_2420,N_2229,N_2279);
nor U2421 (N_2421,N_2334,N_2339);
or U2422 (N_2422,N_2296,N_2243);
and U2423 (N_2423,N_2212,N_2206);
xor U2424 (N_2424,N_2205,N_2388);
nor U2425 (N_2425,N_2284,N_2280);
or U2426 (N_2426,N_2215,N_2242);
and U2427 (N_2427,N_2396,N_2352);
and U2428 (N_2428,N_2308,N_2228);
nor U2429 (N_2429,N_2383,N_2213);
and U2430 (N_2430,N_2378,N_2289);
nor U2431 (N_2431,N_2248,N_2359);
or U2432 (N_2432,N_2202,N_2258);
nor U2433 (N_2433,N_2348,N_2253);
and U2434 (N_2434,N_2288,N_2221);
nor U2435 (N_2435,N_2204,N_2224);
and U2436 (N_2436,N_2393,N_2268);
nand U2437 (N_2437,N_2330,N_2249);
or U2438 (N_2438,N_2398,N_2272);
nor U2439 (N_2439,N_2385,N_2327);
nand U2440 (N_2440,N_2357,N_2364);
nor U2441 (N_2441,N_2246,N_2342);
and U2442 (N_2442,N_2282,N_2216);
and U2443 (N_2443,N_2363,N_2238);
nand U2444 (N_2444,N_2276,N_2211);
or U2445 (N_2445,N_2267,N_2337);
nand U2446 (N_2446,N_2354,N_2208);
and U2447 (N_2447,N_2251,N_2254);
and U2448 (N_2448,N_2333,N_2370);
nor U2449 (N_2449,N_2384,N_2374);
or U2450 (N_2450,N_2247,N_2340);
nand U2451 (N_2451,N_2270,N_2390);
nor U2452 (N_2452,N_2293,N_2394);
and U2453 (N_2453,N_2307,N_2371);
or U2454 (N_2454,N_2274,N_2319);
nand U2455 (N_2455,N_2292,N_2266);
nor U2456 (N_2456,N_2225,N_2250);
xor U2457 (N_2457,N_2325,N_2372);
nor U2458 (N_2458,N_2200,N_2397);
nand U2459 (N_2459,N_2316,N_2263);
nor U2460 (N_2460,N_2245,N_2355);
nand U2461 (N_2461,N_2336,N_2295);
nand U2462 (N_2462,N_2381,N_2235);
nand U2463 (N_2463,N_2244,N_2392);
nor U2464 (N_2464,N_2311,N_2313);
and U2465 (N_2465,N_2257,N_2230);
nand U2466 (N_2466,N_2303,N_2240);
nor U2467 (N_2467,N_2219,N_2350);
nor U2468 (N_2468,N_2345,N_2281);
nand U2469 (N_2469,N_2310,N_2278);
or U2470 (N_2470,N_2399,N_2223);
or U2471 (N_2471,N_2347,N_2252);
nand U2472 (N_2472,N_2353,N_2201);
nand U2473 (N_2473,N_2283,N_2220);
and U2474 (N_2474,N_2294,N_2324);
or U2475 (N_2475,N_2375,N_2317);
xnor U2476 (N_2476,N_2264,N_2300);
or U2477 (N_2477,N_2376,N_2298);
and U2478 (N_2478,N_2379,N_2299);
nor U2479 (N_2479,N_2344,N_2389);
nand U2480 (N_2480,N_2227,N_2387);
nor U2481 (N_2481,N_2366,N_2271);
xnor U2482 (N_2482,N_2210,N_2323);
or U2483 (N_2483,N_2226,N_2259);
or U2484 (N_2484,N_2286,N_2306);
nand U2485 (N_2485,N_2358,N_2269);
nand U2486 (N_2486,N_2341,N_2356);
and U2487 (N_2487,N_2277,N_2265);
nor U2488 (N_2488,N_2329,N_2312);
xor U2489 (N_2489,N_2351,N_2304);
and U2490 (N_2490,N_2241,N_2367);
or U2491 (N_2491,N_2232,N_2328);
and U2492 (N_2492,N_2314,N_2301);
nand U2493 (N_2493,N_2302,N_2373);
nor U2494 (N_2494,N_2365,N_2343);
or U2495 (N_2495,N_2275,N_2331);
and U2496 (N_2496,N_2322,N_2236);
and U2497 (N_2497,N_2395,N_2315);
or U2498 (N_2498,N_2260,N_2377);
or U2499 (N_2499,N_2321,N_2382);
and U2500 (N_2500,N_2350,N_2382);
and U2501 (N_2501,N_2394,N_2257);
nor U2502 (N_2502,N_2353,N_2316);
nor U2503 (N_2503,N_2349,N_2391);
nand U2504 (N_2504,N_2276,N_2385);
nand U2505 (N_2505,N_2238,N_2223);
nand U2506 (N_2506,N_2391,N_2327);
nand U2507 (N_2507,N_2399,N_2379);
and U2508 (N_2508,N_2332,N_2347);
or U2509 (N_2509,N_2229,N_2369);
and U2510 (N_2510,N_2243,N_2226);
nor U2511 (N_2511,N_2372,N_2285);
or U2512 (N_2512,N_2302,N_2275);
or U2513 (N_2513,N_2398,N_2305);
or U2514 (N_2514,N_2259,N_2286);
or U2515 (N_2515,N_2327,N_2386);
nand U2516 (N_2516,N_2244,N_2373);
nor U2517 (N_2517,N_2320,N_2212);
nor U2518 (N_2518,N_2249,N_2345);
or U2519 (N_2519,N_2351,N_2210);
and U2520 (N_2520,N_2277,N_2305);
or U2521 (N_2521,N_2201,N_2261);
nor U2522 (N_2522,N_2330,N_2378);
nand U2523 (N_2523,N_2380,N_2227);
or U2524 (N_2524,N_2342,N_2272);
nand U2525 (N_2525,N_2269,N_2334);
or U2526 (N_2526,N_2289,N_2395);
nand U2527 (N_2527,N_2317,N_2285);
or U2528 (N_2528,N_2345,N_2254);
nand U2529 (N_2529,N_2221,N_2224);
xnor U2530 (N_2530,N_2365,N_2274);
and U2531 (N_2531,N_2318,N_2295);
nand U2532 (N_2532,N_2254,N_2315);
and U2533 (N_2533,N_2314,N_2208);
and U2534 (N_2534,N_2375,N_2217);
nor U2535 (N_2535,N_2369,N_2336);
and U2536 (N_2536,N_2389,N_2399);
nor U2537 (N_2537,N_2313,N_2218);
and U2538 (N_2538,N_2249,N_2271);
xor U2539 (N_2539,N_2387,N_2251);
nand U2540 (N_2540,N_2353,N_2314);
nor U2541 (N_2541,N_2303,N_2208);
and U2542 (N_2542,N_2231,N_2354);
or U2543 (N_2543,N_2201,N_2323);
nor U2544 (N_2544,N_2373,N_2303);
nand U2545 (N_2545,N_2311,N_2254);
and U2546 (N_2546,N_2224,N_2349);
nor U2547 (N_2547,N_2399,N_2364);
and U2548 (N_2548,N_2368,N_2263);
or U2549 (N_2549,N_2229,N_2264);
and U2550 (N_2550,N_2351,N_2305);
nor U2551 (N_2551,N_2372,N_2283);
or U2552 (N_2552,N_2229,N_2294);
nor U2553 (N_2553,N_2395,N_2215);
xor U2554 (N_2554,N_2239,N_2380);
nor U2555 (N_2555,N_2309,N_2203);
or U2556 (N_2556,N_2208,N_2345);
and U2557 (N_2557,N_2227,N_2241);
nand U2558 (N_2558,N_2383,N_2247);
nand U2559 (N_2559,N_2238,N_2385);
or U2560 (N_2560,N_2245,N_2396);
and U2561 (N_2561,N_2246,N_2360);
and U2562 (N_2562,N_2317,N_2201);
nor U2563 (N_2563,N_2256,N_2369);
nand U2564 (N_2564,N_2395,N_2290);
or U2565 (N_2565,N_2373,N_2220);
nand U2566 (N_2566,N_2218,N_2209);
nor U2567 (N_2567,N_2368,N_2253);
or U2568 (N_2568,N_2265,N_2248);
nor U2569 (N_2569,N_2205,N_2299);
or U2570 (N_2570,N_2253,N_2306);
nor U2571 (N_2571,N_2202,N_2341);
xor U2572 (N_2572,N_2246,N_2249);
nand U2573 (N_2573,N_2203,N_2208);
nand U2574 (N_2574,N_2379,N_2266);
or U2575 (N_2575,N_2393,N_2301);
nor U2576 (N_2576,N_2338,N_2308);
and U2577 (N_2577,N_2202,N_2392);
nor U2578 (N_2578,N_2227,N_2330);
nor U2579 (N_2579,N_2318,N_2202);
and U2580 (N_2580,N_2223,N_2228);
or U2581 (N_2581,N_2327,N_2395);
nor U2582 (N_2582,N_2254,N_2238);
nand U2583 (N_2583,N_2203,N_2397);
nand U2584 (N_2584,N_2256,N_2347);
or U2585 (N_2585,N_2279,N_2296);
nand U2586 (N_2586,N_2375,N_2313);
nand U2587 (N_2587,N_2213,N_2341);
nor U2588 (N_2588,N_2209,N_2318);
nor U2589 (N_2589,N_2326,N_2259);
nand U2590 (N_2590,N_2236,N_2343);
or U2591 (N_2591,N_2251,N_2318);
or U2592 (N_2592,N_2240,N_2319);
nor U2593 (N_2593,N_2262,N_2366);
or U2594 (N_2594,N_2399,N_2338);
nand U2595 (N_2595,N_2375,N_2291);
or U2596 (N_2596,N_2306,N_2343);
xnor U2597 (N_2597,N_2298,N_2346);
or U2598 (N_2598,N_2235,N_2283);
nand U2599 (N_2599,N_2397,N_2280);
nor U2600 (N_2600,N_2595,N_2597);
and U2601 (N_2601,N_2468,N_2483);
nand U2602 (N_2602,N_2439,N_2482);
nand U2603 (N_2603,N_2427,N_2415);
nor U2604 (N_2604,N_2453,N_2425);
or U2605 (N_2605,N_2551,N_2591);
or U2606 (N_2606,N_2519,N_2447);
nand U2607 (N_2607,N_2501,N_2525);
nand U2608 (N_2608,N_2517,N_2410);
xor U2609 (N_2609,N_2492,N_2516);
or U2610 (N_2610,N_2476,N_2592);
or U2611 (N_2611,N_2546,N_2424);
and U2612 (N_2612,N_2426,N_2544);
or U2613 (N_2613,N_2481,N_2520);
and U2614 (N_2614,N_2474,N_2448);
or U2615 (N_2615,N_2547,N_2454);
and U2616 (N_2616,N_2580,N_2464);
and U2617 (N_2617,N_2495,N_2573);
nor U2618 (N_2618,N_2477,N_2534);
xor U2619 (N_2619,N_2512,N_2434);
or U2620 (N_2620,N_2506,N_2437);
nand U2621 (N_2621,N_2560,N_2462);
and U2622 (N_2622,N_2507,N_2574);
xor U2623 (N_2623,N_2478,N_2496);
nand U2624 (N_2624,N_2504,N_2555);
nand U2625 (N_2625,N_2406,N_2451);
xor U2626 (N_2626,N_2589,N_2473);
nand U2627 (N_2627,N_2443,N_2433);
xor U2628 (N_2628,N_2577,N_2570);
or U2629 (N_2629,N_2400,N_2444);
xor U2630 (N_2630,N_2442,N_2561);
or U2631 (N_2631,N_2508,N_2461);
or U2632 (N_2632,N_2562,N_2419);
or U2633 (N_2633,N_2423,N_2408);
and U2634 (N_2634,N_2584,N_2490);
xor U2635 (N_2635,N_2449,N_2550);
or U2636 (N_2636,N_2450,N_2485);
nand U2637 (N_2637,N_2553,N_2554);
or U2638 (N_2638,N_2446,N_2533);
or U2639 (N_2639,N_2532,N_2575);
and U2640 (N_2640,N_2421,N_2515);
xnor U2641 (N_2641,N_2431,N_2536);
nand U2642 (N_2642,N_2404,N_2432);
and U2643 (N_2643,N_2489,N_2548);
and U2644 (N_2644,N_2526,N_2572);
xnor U2645 (N_2645,N_2499,N_2552);
nor U2646 (N_2646,N_2440,N_2565);
nand U2647 (N_2647,N_2529,N_2488);
nor U2648 (N_2648,N_2503,N_2409);
or U2649 (N_2649,N_2586,N_2564);
nor U2650 (N_2650,N_2556,N_2445);
and U2651 (N_2651,N_2510,N_2559);
nor U2652 (N_2652,N_2417,N_2469);
nor U2653 (N_2653,N_2568,N_2537);
nor U2654 (N_2654,N_2545,N_2502);
or U2655 (N_2655,N_2518,N_2522);
xnor U2656 (N_2656,N_2405,N_2514);
nor U2657 (N_2657,N_2416,N_2500);
or U2658 (N_2658,N_2505,N_2466);
nor U2659 (N_2659,N_2498,N_2598);
nor U2660 (N_2660,N_2470,N_2588);
nor U2661 (N_2661,N_2558,N_2458);
nor U2662 (N_2662,N_2467,N_2491);
and U2663 (N_2663,N_2402,N_2528);
and U2664 (N_2664,N_2494,N_2413);
nand U2665 (N_2665,N_2549,N_2484);
and U2666 (N_2666,N_2583,N_2414);
and U2667 (N_2667,N_2541,N_2422);
nand U2668 (N_2668,N_2487,N_2531);
or U2669 (N_2669,N_2566,N_2540);
and U2670 (N_2670,N_2582,N_2441);
nand U2671 (N_2671,N_2457,N_2428);
or U2672 (N_2672,N_2438,N_2535);
nand U2673 (N_2673,N_2456,N_2571);
and U2674 (N_2674,N_2480,N_2542);
xor U2675 (N_2675,N_2569,N_2578);
or U2676 (N_2676,N_2435,N_2593);
or U2677 (N_2677,N_2418,N_2472);
nand U2678 (N_2678,N_2594,N_2563);
or U2679 (N_2679,N_2509,N_2539);
or U2680 (N_2680,N_2581,N_2479);
nor U2681 (N_2681,N_2513,N_2521);
nand U2682 (N_2682,N_2411,N_2497);
nand U2683 (N_2683,N_2587,N_2596);
and U2684 (N_2684,N_2530,N_2599);
nand U2685 (N_2685,N_2459,N_2576);
or U2686 (N_2686,N_2557,N_2524);
nand U2687 (N_2687,N_2452,N_2493);
or U2688 (N_2688,N_2475,N_2401);
xnor U2689 (N_2689,N_2430,N_2527);
or U2690 (N_2690,N_2465,N_2403);
or U2691 (N_2691,N_2579,N_2471);
and U2692 (N_2692,N_2567,N_2463);
and U2693 (N_2693,N_2429,N_2585);
nor U2694 (N_2694,N_2523,N_2538);
nor U2695 (N_2695,N_2436,N_2412);
or U2696 (N_2696,N_2420,N_2407);
and U2697 (N_2697,N_2486,N_2543);
and U2698 (N_2698,N_2460,N_2511);
or U2699 (N_2699,N_2455,N_2590);
xor U2700 (N_2700,N_2493,N_2508);
and U2701 (N_2701,N_2431,N_2538);
and U2702 (N_2702,N_2456,N_2573);
nor U2703 (N_2703,N_2419,N_2512);
or U2704 (N_2704,N_2572,N_2503);
and U2705 (N_2705,N_2415,N_2569);
and U2706 (N_2706,N_2547,N_2569);
or U2707 (N_2707,N_2422,N_2496);
or U2708 (N_2708,N_2565,N_2515);
or U2709 (N_2709,N_2426,N_2463);
nor U2710 (N_2710,N_2440,N_2587);
nor U2711 (N_2711,N_2424,N_2429);
nand U2712 (N_2712,N_2447,N_2587);
xnor U2713 (N_2713,N_2450,N_2410);
nor U2714 (N_2714,N_2485,N_2424);
xnor U2715 (N_2715,N_2567,N_2445);
or U2716 (N_2716,N_2438,N_2521);
and U2717 (N_2717,N_2541,N_2491);
nand U2718 (N_2718,N_2588,N_2438);
nor U2719 (N_2719,N_2542,N_2414);
xnor U2720 (N_2720,N_2597,N_2582);
nand U2721 (N_2721,N_2474,N_2500);
nor U2722 (N_2722,N_2423,N_2522);
nor U2723 (N_2723,N_2486,N_2553);
xor U2724 (N_2724,N_2563,N_2567);
xnor U2725 (N_2725,N_2401,N_2553);
nand U2726 (N_2726,N_2542,N_2594);
nand U2727 (N_2727,N_2421,N_2464);
nand U2728 (N_2728,N_2416,N_2453);
nand U2729 (N_2729,N_2508,N_2589);
or U2730 (N_2730,N_2501,N_2458);
nand U2731 (N_2731,N_2505,N_2508);
nor U2732 (N_2732,N_2535,N_2427);
or U2733 (N_2733,N_2486,N_2568);
and U2734 (N_2734,N_2513,N_2449);
or U2735 (N_2735,N_2472,N_2428);
and U2736 (N_2736,N_2422,N_2512);
or U2737 (N_2737,N_2489,N_2459);
and U2738 (N_2738,N_2529,N_2493);
xnor U2739 (N_2739,N_2595,N_2482);
and U2740 (N_2740,N_2432,N_2464);
nand U2741 (N_2741,N_2478,N_2406);
and U2742 (N_2742,N_2569,N_2556);
and U2743 (N_2743,N_2410,N_2408);
nor U2744 (N_2744,N_2478,N_2583);
nor U2745 (N_2745,N_2460,N_2519);
nand U2746 (N_2746,N_2544,N_2421);
or U2747 (N_2747,N_2437,N_2550);
and U2748 (N_2748,N_2402,N_2598);
xnor U2749 (N_2749,N_2451,N_2530);
and U2750 (N_2750,N_2460,N_2561);
nor U2751 (N_2751,N_2414,N_2523);
and U2752 (N_2752,N_2588,N_2499);
nor U2753 (N_2753,N_2439,N_2523);
nand U2754 (N_2754,N_2497,N_2545);
and U2755 (N_2755,N_2410,N_2422);
and U2756 (N_2756,N_2547,N_2542);
or U2757 (N_2757,N_2489,N_2586);
nor U2758 (N_2758,N_2512,N_2467);
xnor U2759 (N_2759,N_2480,N_2484);
nor U2760 (N_2760,N_2571,N_2596);
nand U2761 (N_2761,N_2522,N_2417);
or U2762 (N_2762,N_2513,N_2493);
nor U2763 (N_2763,N_2537,N_2599);
and U2764 (N_2764,N_2505,N_2472);
or U2765 (N_2765,N_2534,N_2469);
and U2766 (N_2766,N_2428,N_2512);
nand U2767 (N_2767,N_2526,N_2483);
or U2768 (N_2768,N_2431,N_2569);
nor U2769 (N_2769,N_2461,N_2450);
nor U2770 (N_2770,N_2400,N_2549);
or U2771 (N_2771,N_2528,N_2540);
xor U2772 (N_2772,N_2476,N_2497);
xnor U2773 (N_2773,N_2567,N_2500);
and U2774 (N_2774,N_2571,N_2483);
nor U2775 (N_2775,N_2531,N_2422);
or U2776 (N_2776,N_2434,N_2532);
nand U2777 (N_2777,N_2588,N_2423);
nor U2778 (N_2778,N_2509,N_2409);
nor U2779 (N_2779,N_2566,N_2407);
or U2780 (N_2780,N_2401,N_2574);
nor U2781 (N_2781,N_2447,N_2524);
xnor U2782 (N_2782,N_2439,N_2574);
nand U2783 (N_2783,N_2549,N_2562);
nand U2784 (N_2784,N_2426,N_2576);
or U2785 (N_2785,N_2552,N_2563);
nand U2786 (N_2786,N_2534,N_2459);
or U2787 (N_2787,N_2409,N_2530);
and U2788 (N_2788,N_2517,N_2451);
nor U2789 (N_2789,N_2559,N_2546);
xnor U2790 (N_2790,N_2554,N_2445);
nand U2791 (N_2791,N_2465,N_2458);
nand U2792 (N_2792,N_2475,N_2471);
and U2793 (N_2793,N_2532,N_2441);
nand U2794 (N_2794,N_2591,N_2553);
and U2795 (N_2795,N_2563,N_2542);
nand U2796 (N_2796,N_2439,N_2507);
xnor U2797 (N_2797,N_2598,N_2403);
or U2798 (N_2798,N_2434,N_2437);
or U2799 (N_2799,N_2420,N_2529);
nand U2800 (N_2800,N_2672,N_2616);
nor U2801 (N_2801,N_2699,N_2769);
and U2802 (N_2802,N_2650,N_2741);
nor U2803 (N_2803,N_2747,N_2702);
and U2804 (N_2804,N_2754,N_2762);
nor U2805 (N_2805,N_2749,N_2736);
xnor U2806 (N_2806,N_2631,N_2728);
nor U2807 (N_2807,N_2618,N_2644);
nand U2808 (N_2808,N_2692,N_2784);
xnor U2809 (N_2809,N_2770,N_2629);
or U2810 (N_2810,N_2658,N_2601);
and U2811 (N_2811,N_2767,N_2655);
xnor U2812 (N_2812,N_2796,N_2607);
nand U2813 (N_2813,N_2630,N_2662);
nor U2814 (N_2814,N_2606,N_2712);
nand U2815 (N_2815,N_2775,N_2757);
nor U2816 (N_2816,N_2697,N_2759);
and U2817 (N_2817,N_2676,N_2647);
nand U2818 (N_2818,N_2758,N_2623);
xnor U2819 (N_2819,N_2788,N_2792);
xor U2820 (N_2820,N_2635,N_2772);
nor U2821 (N_2821,N_2642,N_2654);
nand U2822 (N_2822,N_2782,N_2790);
nand U2823 (N_2823,N_2619,N_2681);
or U2824 (N_2824,N_2717,N_2738);
or U2825 (N_2825,N_2696,N_2704);
xnor U2826 (N_2826,N_2660,N_2646);
and U2827 (N_2827,N_2708,N_2764);
xnor U2828 (N_2828,N_2724,N_2611);
or U2829 (N_2829,N_2703,N_2726);
nand U2830 (N_2830,N_2636,N_2670);
nor U2831 (N_2831,N_2604,N_2760);
nor U2832 (N_2832,N_2682,N_2729);
or U2833 (N_2833,N_2771,N_2612);
or U2834 (N_2834,N_2637,N_2665);
and U2835 (N_2835,N_2657,N_2698);
nor U2836 (N_2836,N_2765,N_2716);
and U2837 (N_2837,N_2661,N_2689);
and U2838 (N_2838,N_2732,N_2600);
nor U2839 (N_2839,N_2648,N_2735);
xor U2840 (N_2840,N_2615,N_2641);
and U2841 (N_2841,N_2779,N_2627);
and U2842 (N_2842,N_2668,N_2628);
and U2843 (N_2843,N_2742,N_2687);
nand U2844 (N_2844,N_2713,N_2781);
nor U2845 (N_2845,N_2626,N_2667);
nand U2846 (N_2846,N_2603,N_2797);
and U2847 (N_2847,N_2707,N_2643);
nor U2848 (N_2848,N_2622,N_2746);
nand U2849 (N_2849,N_2679,N_2617);
or U2850 (N_2850,N_2649,N_2602);
nor U2851 (N_2851,N_2798,N_2783);
nor U2852 (N_2852,N_2691,N_2730);
nand U2853 (N_2853,N_2686,N_2663);
nand U2854 (N_2854,N_2799,N_2723);
or U2855 (N_2855,N_2632,N_2659);
nor U2856 (N_2856,N_2669,N_2763);
and U2857 (N_2857,N_2620,N_2621);
and U2858 (N_2858,N_2674,N_2768);
or U2859 (N_2859,N_2785,N_2720);
or U2860 (N_2860,N_2651,N_2778);
xnor U2861 (N_2861,N_2718,N_2680);
nand U2862 (N_2862,N_2605,N_2734);
nand U2863 (N_2863,N_2761,N_2656);
and U2864 (N_2864,N_2795,N_2613);
or U2865 (N_2865,N_2777,N_2733);
nor U2866 (N_2866,N_2693,N_2752);
nor U2867 (N_2867,N_2700,N_2743);
nand U2868 (N_2868,N_2710,N_2721);
and U2869 (N_2869,N_2695,N_2624);
or U2870 (N_2870,N_2694,N_2675);
xor U2871 (N_2871,N_2673,N_2714);
and U2872 (N_2872,N_2705,N_2671);
nand U2873 (N_2873,N_2652,N_2653);
and U2874 (N_2874,N_2634,N_2731);
or U2875 (N_2875,N_2678,N_2639);
and U2876 (N_2876,N_2719,N_2740);
nor U2877 (N_2877,N_2727,N_2633);
and U2878 (N_2878,N_2638,N_2614);
nand U2879 (N_2879,N_2793,N_2755);
and U2880 (N_2880,N_2608,N_2745);
nand U2881 (N_2881,N_2690,N_2794);
nand U2882 (N_2882,N_2756,N_2610);
or U2883 (N_2883,N_2753,N_2645);
or U2884 (N_2884,N_2773,N_2789);
and U2885 (N_2885,N_2737,N_2776);
nand U2886 (N_2886,N_2744,N_2748);
and U2887 (N_2887,N_2786,N_2688);
xor U2888 (N_2888,N_2791,N_2640);
nor U2889 (N_2889,N_2711,N_2715);
and U2890 (N_2890,N_2722,N_2701);
nor U2891 (N_2891,N_2709,N_2664);
or U2892 (N_2892,N_2787,N_2677);
or U2893 (N_2893,N_2683,N_2685);
nor U2894 (N_2894,N_2666,N_2625);
and U2895 (N_2895,N_2706,N_2751);
and U2896 (N_2896,N_2766,N_2774);
nor U2897 (N_2897,N_2750,N_2725);
nand U2898 (N_2898,N_2739,N_2609);
or U2899 (N_2899,N_2780,N_2684);
nand U2900 (N_2900,N_2698,N_2638);
and U2901 (N_2901,N_2697,N_2676);
and U2902 (N_2902,N_2685,N_2704);
or U2903 (N_2903,N_2730,N_2703);
xor U2904 (N_2904,N_2794,N_2632);
nand U2905 (N_2905,N_2730,N_2634);
or U2906 (N_2906,N_2776,N_2660);
xor U2907 (N_2907,N_2731,N_2736);
or U2908 (N_2908,N_2738,N_2774);
nand U2909 (N_2909,N_2770,N_2663);
and U2910 (N_2910,N_2617,N_2701);
xnor U2911 (N_2911,N_2629,N_2711);
nor U2912 (N_2912,N_2791,N_2607);
nor U2913 (N_2913,N_2762,N_2633);
nor U2914 (N_2914,N_2630,N_2769);
nor U2915 (N_2915,N_2705,N_2626);
nand U2916 (N_2916,N_2614,N_2765);
and U2917 (N_2917,N_2624,N_2638);
or U2918 (N_2918,N_2734,N_2626);
nand U2919 (N_2919,N_2605,N_2634);
and U2920 (N_2920,N_2694,N_2721);
or U2921 (N_2921,N_2794,N_2682);
or U2922 (N_2922,N_2777,N_2767);
nand U2923 (N_2923,N_2624,N_2753);
nand U2924 (N_2924,N_2766,N_2613);
nand U2925 (N_2925,N_2666,N_2752);
and U2926 (N_2926,N_2717,N_2713);
xnor U2927 (N_2927,N_2713,N_2732);
and U2928 (N_2928,N_2765,N_2680);
nor U2929 (N_2929,N_2617,N_2647);
nor U2930 (N_2930,N_2653,N_2673);
xor U2931 (N_2931,N_2779,N_2766);
or U2932 (N_2932,N_2749,N_2706);
nand U2933 (N_2933,N_2643,N_2646);
and U2934 (N_2934,N_2637,N_2781);
and U2935 (N_2935,N_2724,N_2750);
and U2936 (N_2936,N_2678,N_2656);
nand U2937 (N_2937,N_2772,N_2619);
and U2938 (N_2938,N_2618,N_2725);
or U2939 (N_2939,N_2783,N_2657);
or U2940 (N_2940,N_2698,N_2764);
nand U2941 (N_2941,N_2793,N_2704);
nor U2942 (N_2942,N_2673,N_2670);
and U2943 (N_2943,N_2773,N_2704);
nor U2944 (N_2944,N_2721,N_2757);
and U2945 (N_2945,N_2632,N_2604);
and U2946 (N_2946,N_2775,N_2611);
and U2947 (N_2947,N_2684,N_2682);
or U2948 (N_2948,N_2660,N_2661);
or U2949 (N_2949,N_2753,N_2631);
nor U2950 (N_2950,N_2708,N_2640);
xnor U2951 (N_2951,N_2738,N_2711);
and U2952 (N_2952,N_2715,N_2624);
xor U2953 (N_2953,N_2651,N_2604);
or U2954 (N_2954,N_2620,N_2676);
nor U2955 (N_2955,N_2687,N_2673);
and U2956 (N_2956,N_2768,N_2770);
or U2957 (N_2957,N_2674,N_2725);
nand U2958 (N_2958,N_2667,N_2650);
nand U2959 (N_2959,N_2740,N_2645);
and U2960 (N_2960,N_2637,N_2644);
and U2961 (N_2961,N_2601,N_2760);
nand U2962 (N_2962,N_2608,N_2758);
nor U2963 (N_2963,N_2660,N_2761);
xnor U2964 (N_2964,N_2698,N_2752);
and U2965 (N_2965,N_2797,N_2600);
and U2966 (N_2966,N_2631,N_2628);
nand U2967 (N_2967,N_2628,N_2706);
or U2968 (N_2968,N_2760,N_2794);
xor U2969 (N_2969,N_2693,N_2713);
or U2970 (N_2970,N_2636,N_2738);
and U2971 (N_2971,N_2681,N_2655);
and U2972 (N_2972,N_2625,N_2758);
nand U2973 (N_2973,N_2662,N_2605);
or U2974 (N_2974,N_2778,N_2703);
nor U2975 (N_2975,N_2683,N_2743);
nor U2976 (N_2976,N_2757,N_2607);
xor U2977 (N_2977,N_2722,N_2695);
or U2978 (N_2978,N_2731,N_2773);
and U2979 (N_2979,N_2753,N_2684);
xnor U2980 (N_2980,N_2615,N_2670);
nand U2981 (N_2981,N_2764,N_2704);
or U2982 (N_2982,N_2645,N_2661);
or U2983 (N_2983,N_2606,N_2708);
nand U2984 (N_2984,N_2636,N_2677);
nor U2985 (N_2985,N_2619,N_2724);
or U2986 (N_2986,N_2618,N_2707);
nand U2987 (N_2987,N_2625,N_2621);
and U2988 (N_2988,N_2777,N_2734);
nand U2989 (N_2989,N_2723,N_2618);
or U2990 (N_2990,N_2704,N_2621);
nor U2991 (N_2991,N_2728,N_2785);
or U2992 (N_2992,N_2667,N_2701);
nor U2993 (N_2993,N_2719,N_2630);
nand U2994 (N_2994,N_2738,N_2633);
or U2995 (N_2995,N_2635,N_2690);
or U2996 (N_2996,N_2673,N_2753);
or U2997 (N_2997,N_2790,N_2707);
nor U2998 (N_2998,N_2632,N_2766);
and U2999 (N_2999,N_2624,N_2689);
or UO_0 (O_0,N_2802,N_2805);
and UO_1 (O_1,N_2894,N_2973);
nand UO_2 (O_2,N_2829,N_2853);
nand UO_3 (O_3,N_2851,N_2856);
and UO_4 (O_4,N_2911,N_2825);
and UO_5 (O_5,N_2890,N_2954);
nor UO_6 (O_6,N_2884,N_2883);
and UO_7 (O_7,N_2907,N_2918);
nand UO_8 (O_8,N_2960,N_2925);
nor UO_9 (O_9,N_2833,N_2878);
and UO_10 (O_10,N_2940,N_2821);
or UO_11 (O_11,N_2835,N_2882);
nor UO_12 (O_12,N_2866,N_2898);
nor UO_13 (O_13,N_2921,N_2932);
or UO_14 (O_14,N_2948,N_2803);
xor UO_15 (O_15,N_2994,N_2974);
nor UO_16 (O_16,N_2844,N_2951);
and UO_17 (O_17,N_2813,N_2831);
nand UO_18 (O_18,N_2822,N_2809);
nor UO_19 (O_19,N_2826,N_2859);
nor UO_20 (O_20,N_2817,N_2855);
and UO_21 (O_21,N_2942,N_2820);
xnor UO_22 (O_22,N_2819,N_2810);
and UO_23 (O_23,N_2931,N_2958);
nand UO_24 (O_24,N_2947,N_2916);
or UO_25 (O_25,N_2956,N_2967);
or UO_26 (O_26,N_2879,N_2804);
and UO_27 (O_27,N_2935,N_2945);
or UO_28 (O_28,N_2961,N_2834);
and UO_29 (O_29,N_2902,N_2816);
nor UO_30 (O_30,N_2842,N_2910);
nor UO_31 (O_31,N_2887,N_2992);
or UO_32 (O_32,N_2926,N_2801);
and UO_33 (O_33,N_2872,N_2892);
or UO_34 (O_34,N_2936,N_2905);
nand UO_35 (O_35,N_2899,N_2857);
or UO_36 (O_36,N_2852,N_2854);
nand UO_37 (O_37,N_2895,N_2888);
nand UO_38 (O_38,N_2846,N_2847);
and UO_39 (O_39,N_2998,N_2873);
and UO_40 (O_40,N_2996,N_2862);
or UO_41 (O_41,N_2995,N_2848);
nand UO_42 (O_42,N_2949,N_2966);
or UO_43 (O_43,N_2811,N_2987);
and UO_44 (O_44,N_2923,N_2999);
nor UO_45 (O_45,N_2818,N_2955);
nor UO_46 (O_46,N_2850,N_2893);
nor UO_47 (O_47,N_2843,N_2800);
or UO_48 (O_48,N_2927,N_2946);
nor UO_49 (O_49,N_2912,N_2944);
nor UO_50 (O_50,N_2929,N_2827);
and UO_51 (O_51,N_2900,N_2934);
nand UO_52 (O_52,N_2979,N_2824);
nand UO_53 (O_53,N_2908,N_2832);
nor UO_54 (O_54,N_2904,N_2922);
or UO_55 (O_55,N_2864,N_2814);
nand UO_56 (O_56,N_2930,N_2889);
xnor UO_57 (O_57,N_2913,N_2867);
nand UO_58 (O_58,N_2975,N_2875);
or UO_59 (O_59,N_2978,N_2840);
nand UO_60 (O_60,N_2919,N_2953);
or UO_61 (O_61,N_2982,N_2830);
nor UO_62 (O_62,N_2896,N_2986);
nor UO_63 (O_63,N_2976,N_2984);
nand UO_64 (O_64,N_2876,N_2849);
and UO_65 (O_65,N_2965,N_2968);
or UO_66 (O_66,N_2962,N_2828);
xor UO_67 (O_67,N_2980,N_2808);
nand UO_68 (O_68,N_2957,N_2812);
or UO_69 (O_69,N_2988,N_2891);
nand UO_70 (O_70,N_2920,N_2970);
nor UO_71 (O_71,N_2815,N_2997);
xor UO_72 (O_72,N_2880,N_2928);
and UO_73 (O_73,N_2985,N_2877);
nand UO_74 (O_74,N_2903,N_2981);
xor UO_75 (O_75,N_2963,N_2993);
and UO_76 (O_76,N_2917,N_2991);
xor UO_77 (O_77,N_2901,N_2906);
xor UO_78 (O_78,N_2941,N_2909);
nand UO_79 (O_79,N_2937,N_2989);
xnor UO_80 (O_80,N_2869,N_2914);
nand UO_81 (O_81,N_2885,N_2806);
or UO_82 (O_82,N_2838,N_2924);
and UO_83 (O_83,N_2977,N_2841);
or UO_84 (O_84,N_2990,N_2839);
and UO_85 (O_85,N_2939,N_2881);
nor UO_86 (O_86,N_2969,N_2952);
or UO_87 (O_87,N_2972,N_2861);
nand UO_88 (O_88,N_2933,N_2863);
or UO_89 (O_89,N_2964,N_2897);
nor UO_90 (O_90,N_2938,N_2971);
or UO_91 (O_91,N_2837,N_2868);
and UO_92 (O_92,N_2845,N_2959);
nand UO_93 (O_93,N_2983,N_2871);
nand UO_94 (O_94,N_2823,N_2870);
and UO_95 (O_95,N_2836,N_2943);
xnor UO_96 (O_96,N_2865,N_2874);
or UO_97 (O_97,N_2950,N_2886);
nor UO_98 (O_98,N_2858,N_2915);
nor UO_99 (O_99,N_2860,N_2807);
nand UO_100 (O_100,N_2948,N_2890);
nor UO_101 (O_101,N_2893,N_2922);
or UO_102 (O_102,N_2994,N_2818);
nor UO_103 (O_103,N_2899,N_2882);
nor UO_104 (O_104,N_2896,N_2803);
xor UO_105 (O_105,N_2920,N_2830);
and UO_106 (O_106,N_2914,N_2865);
nor UO_107 (O_107,N_2967,N_2919);
and UO_108 (O_108,N_2953,N_2893);
or UO_109 (O_109,N_2821,N_2893);
and UO_110 (O_110,N_2969,N_2961);
nand UO_111 (O_111,N_2825,N_2897);
nor UO_112 (O_112,N_2836,N_2872);
or UO_113 (O_113,N_2977,N_2910);
or UO_114 (O_114,N_2992,N_2969);
or UO_115 (O_115,N_2851,N_2941);
or UO_116 (O_116,N_2942,N_2964);
nor UO_117 (O_117,N_2848,N_2816);
or UO_118 (O_118,N_2971,N_2835);
or UO_119 (O_119,N_2815,N_2853);
nand UO_120 (O_120,N_2827,N_2801);
nor UO_121 (O_121,N_2943,N_2870);
and UO_122 (O_122,N_2804,N_2812);
nand UO_123 (O_123,N_2846,N_2804);
nor UO_124 (O_124,N_2858,N_2902);
nand UO_125 (O_125,N_2989,N_2957);
and UO_126 (O_126,N_2853,N_2950);
nand UO_127 (O_127,N_2898,N_2959);
or UO_128 (O_128,N_2899,N_2965);
or UO_129 (O_129,N_2964,N_2967);
xnor UO_130 (O_130,N_2930,N_2979);
nor UO_131 (O_131,N_2970,N_2812);
nor UO_132 (O_132,N_2801,N_2871);
or UO_133 (O_133,N_2916,N_2862);
and UO_134 (O_134,N_2950,N_2801);
and UO_135 (O_135,N_2859,N_2811);
nor UO_136 (O_136,N_2811,N_2881);
nor UO_137 (O_137,N_2927,N_2997);
and UO_138 (O_138,N_2824,N_2990);
nor UO_139 (O_139,N_2974,N_2992);
and UO_140 (O_140,N_2940,N_2921);
nor UO_141 (O_141,N_2848,N_2844);
nor UO_142 (O_142,N_2940,N_2874);
nand UO_143 (O_143,N_2820,N_2830);
nor UO_144 (O_144,N_2870,N_2830);
nand UO_145 (O_145,N_2906,N_2885);
and UO_146 (O_146,N_2992,N_2902);
nand UO_147 (O_147,N_2950,N_2990);
and UO_148 (O_148,N_2929,N_2800);
or UO_149 (O_149,N_2940,N_2984);
nor UO_150 (O_150,N_2876,N_2954);
nor UO_151 (O_151,N_2971,N_2994);
nand UO_152 (O_152,N_2897,N_2967);
nor UO_153 (O_153,N_2827,N_2919);
and UO_154 (O_154,N_2996,N_2911);
or UO_155 (O_155,N_2901,N_2899);
or UO_156 (O_156,N_2845,N_2905);
xor UO_157 (O_157,N_2978,N_2952);
nand UO_158 (O_158,N_2921,N_2836);
and UO_159 (O_159,N_2999,N_2890);
nor UO_160 (O_160,N_2883,N_2811);
and UO_161 (O_161,N_2929,N_2984);
or UO_162 (O_162,N_2982,N_2961);
nor UO_163 (O_163,N_2828,N_2996);
or UO_164 (O_164,N_2925,N_2817);
and UO_165 (O_165,N_2862,N_2965);
or UO_166 (O_166,N_2971,N_2847);
or UO_167 (O_167,N_2977,N_2806);
xnor UO_168 (O_168,N_2939,N_2821);
xor UO_169 (O_169,N_2988,N_2886);
nand UO_170 (O_170,N_2970,N_2952);
and UO_171 (O_171,N_2910,N_2815);
or UO_172 (O_172,N_2800,N_2839);
and UO_173 (O_173,N_2898,N_2862);
or UO_174 (O_174,N_2835,N_2936);
nand UO_175 (O_175,N_2909,N_2847);
nand UO_176 (O_176,N_2889,N_2877);
and UO_177 (O_177,N_2931,N_2993);
nand UO_178 (O_178,N_2851,N_2964);
and UO_179 (O_179,N_2978,N_2943);
nor UO_180 (O_180,N_2891,N_2984);
or UO_181 (O_181,N_2802,N_2971);
or UO_182 (O_182,N_2963,N_2910);
and UO_183 (O_183,N_2881,N_2993);
or UO_184 (O_184,N_2960,N_2912);
nand UO_185 (O_185,N_2935,N_2949);
nor UO_186 (O_186,N_2922,N_2824);
nor UO_187 (O_187,N_2975,N_2958);
nor UO_188 (O_188,N_2896,N_2853);
or UO_189 (O_189,N_2958,N_2938);
and UO_190 (O_190,N_2903,N_2921);
xnor UO_191 (O_191,N_2804,N_2970);
or UO_192 (O_192,N_2844,N_2825);
and UO_193 (O_193,N_2825,N_2840);
nor UO_194 (O_194,N_2865,N_2994);
nand UO_195 (O_195,N_2986,N_2985);
nand UO_196 (O_196,N_2806,N_2941);
and UO_197 (O_197,N_2810,N_2927);
nand UO_198 (O_198,N_2944,N_2907);
nand UO_199 (O_199,N_2828,N_2852);
nand UO_200 (O_200,N_2939,N_2801);
nor UO_201 (O_201,N_2918,N_2915);
and UO_202 (O_202,N_2804,N_2865);
and UO_203 (O_203,N_2853,N_2920);
and UO_204 (O_204,N_2877,N_2899);
nor UO_205 (O_205,N_2954,N_2934);
xor UO_206 (O_206,N_2816,N_2885);
nor UO_207 (O_207,N_2866,N_2810);
or UO_208 (O_208,N_2868,N_2918);
or UO_209 (O_209,N_2910,N_2911);
nand UO_210 (O_210,N_2950,N_2861);
and UO_211 (O_211,N_2885,N_2810);
and UO_212 (O_212,N_2968,N_2934);
nor UO_213 (O_213,N_2862,N_2910);
nand UO_214 (O_214,N_2975,N_2865);
nand UO_215 (O_215,N_2954,N_2834);
nand UO_216 (O_216,N_2999,N_2814);
or UO_217 (O_217,N_2830,N_2921);
or UO_218 (O_218,N_2916,N_2857);
nand UO_219 (O_219,N_2824,N_2911);
nand UO_220 (O_220,N_2994,N_2804);
nor UO_221 (O_221,N_2879,N_2958);
and UO_222 (O_222,N_2823,N_2932);
xnor UO_223 (O_223,N_2955,N_2885);
or UO_224 (O_224,N_2926,N_2939);
xor UO_225 (O_225,N_2915,N_2988);
and UO_226 (O_226,N_2852,N_2841);
or UO_227 (O_227,N_2845,N_2882);
or UO_228 (O_228,N_2825,N_2829);
nor UO_229 (O_229,N_2889,N_2800);
or UO_230 (O_230,N_2845,N_2824);
nor UO_231 (O_231,N_2824,N_2825);
nand UO_232 (O_232,N_2836,N_2927);
nor UO_233 (O_233,N_2927,N_2895);
nor UO_234 (O_234,N_2842,N_2847);
and UO_235 (O_235,N_2833,N_2896);
nor UO_236 (O_236,N_2880,N_2943);
or UO_237 (O_237,N_2800,N_2887);
nand UO_238 (O_238,N_2844,N_2935);
xnor UO_239 (O_239,N_2981,N_2892);
nor UO_240 (O_240,N_2854,N_2987);
nand UO_241 (O_241,N_2825,N_2827);
or UO_242 (O_242,N_2859,N_2911);
nor UO_243 (O_243,N_2877,N_2831);
or UO_244 (O_244,N_2848,N_2979);
nand UO_245 (O_245,N_2883,N_2851);
and UO_246 (O_246,N_2993,N_2982);
and UO_247 (O_247,N_2813,N_2916);
xnor UO_248 (O_248,N_2990,N_2806);
nand UO_249 (O_249,N_2904,N_2900);
and UO_250 (O_250,N_2812,N_2897);
xor UO_251 (O_251,N_2935,N_2992);
nor UO_252 (O_252,N_2896,N_2842);
nor UO_253 (O_253,N_2858,N_2864);
and UO_254 (O_254,N_2952,N_2862);
and UO_255 (O_255,N_2832,N_2989);
nor UO_256 (O_256,N_2996,N_2868);
nand UO_257 (O_257,N_2931,N_2888);
nor UO_258 (O_258,N_2820,N_2907);
and UO_259 (O_259,N_2993,N_2890);
nor UO_260 (O_260,N_2898,N_2851);
or UO_261 (O_261,N_2959,N_2953);
nand UO_262 (O_262,N_2961,N_2822);
nor UO_263 (O_263,N_2887,N_2946);
nand UO_264 (O_264,N_2899,N_2830);
xor UO_265 (O_265,N_2835,N_2995);
and UO_266 (O_266,N_2853,N_2890);
nor UO_267 (O_267,N_2990,N_2852);
nand UO_268 (O_268,N_2947,N_2955);
nand UO_269 (O_269,N_2893,N_2980);
and UO_270 (O_270,N_2801,N_2892);
nand UO_271 (O_271,N_2824,N_2901);
nand UO_272 (O_272,N_2988,N_2866);
nor UO_273 (O_273,N_2862,N_2925);
xor UO_274 (O_274,N_2846,N_2968);
nor UO_275 (O_275,N_2976,N_2880);
nor UO_276 (O_276,N_2999,N_2869);
xnor UO_277 (O_277,N_2946,N_2842);
nor UO_278 (O_278,N_2918,N_2954);
and UO_279 (O_279,N_2913,N_2988);
or UO_280 (O_280,N_2994,N_2822);
or UO_281 (O_281,N_2916,N_2849);
nor UO_282 (O_282,N_2951,N_2831);
xor UO_283 (O_283,N_2844,N_2886);
or UO_284 (O_284,N_2852,N_2825);
xnor UO_285 (O_285,N_2825,N_2832);
and UO_286 (O_286,N_2906,N_2866);
and UO_287 (O_287,N_2992,N_2892);
or UO_288 (O_288,N_2990,N_2977);
and UO_289 (O_289,N_2994,N_2900);
or UO_290 (O_290,N_2926,N_2866);
nor UO_291 (O_291,N_2875,N_2927);
and UO_292 (O_292,N_2916,N_2951);
nor UO_293 (O_293,N_2915,N_2917);
or UO_294 (O_294,N_2901,N_2828);
and UO_295 (O_295,N_2807,N_2995);
or UO_296 (O_296,N_2809,N_2826);
or UO_297 (O_297,N_2920,N_2828);
nand UO_298 (O_298,N_2823,N_2895);
or UO_299 (O_299,N_2812,N_2814);
nor UO_300 (O_300,N_2867,N_2808);
and UO_301 (O_301,N_2815,N_2917);
xor UO_302 (O_302,N_2923,N_2844);
nor UO_303 (O_303,N_2853,N_2979);
or UO_304 (O_304,N_2902,N_2825);
nor UO_305 (O_305,N_2826,N_2904);
and UO_306 (O_306,N_2823,N_2986);
nor UO_307 (O_307,N_2870,N_2923);
or UO_308 (O_308,N_2964,N_2856);
xnor UO_309 (O_309,N_2839,N_2826);
nor UO_310 (O_310,N_2841,N_2886);
nand UO_311 (O_311,N_2915,N_2877);
and UO_312 (O_312,N_2971,N_2868);
and UO_313 (O_313,N_2876,N_2948);
nand UO_314 (O_314,N_2839,N_2866);
and UO_315 (O_315,N_2897,N_2861);
and UO_316 (O_316,N_2850,N_2961);
nor UO_317 (O_317,N_2877,N_2843);
nor UO_318 (O_318,N_2924,N_2871);
or UO_319 (O_319,N_2933,N_2878);
nand UO_320 (O_320,N_2846,N_2907);
nor UO_321 (O_321,N_2875,N_2895);
nand UO_322 (O_322,N_2974,N_2902);
or UO_323 (O_323,N_2858,N_2949);
nand UO_324 (O_324,N_2969,N_2809);
nor UO_325 (O_325,N_2946,N_2938);
nand UO_326 (O_326,N_2839,N_2994);
xnor UO_327 (O_327,N_2944,N_2826);
nand UO_328 (O_328,N_2908,N_2848);
and UO_329 (O_329,N_2849,N_2872);
nor UO_330 (O_330,N_2873,N_2893);
nand UO_331 (O_331,N_2865,N_2818);
or UO_332 (O_332,N_2894,N_2968);
nor UO_333 (O_333,N_2935,N_2976);
and UO_334 (O_334,N_2934,N_2810);
nand UO_335 (O_335,N_2926,N_2963);
and UO_336 (O_336,N_2873,N_2905);
nand UO_337 (O_337,N_2979,N_2952);
or UO_338 (O_338,N_2984,N_2901);
nor UO_339 (O_339,N_2833,N_2916);
xnor UO_340 (O_340,N_2813,N_2800);
and UO_341 (O_341,N_2805,N_2827);
and UO_342 (O_342,N_2821,N_2846);
xnor UO_343 (O_343,N_2811,N_2850);
and UO_344 (O_344,N_2834,N_2987);
and UO_345 (O_345,N_2893,N_2983);
and UO_346 (O_346,N_2800,N_2866);
xnor UO_347 (O_347,N_2823,N_2816);
xor UO_348 (O_348,N_2865,N_2894);
and UO_349 (O_349,N_2880,N_2844);
nor UO_350 (O_350,N_2973,N_2877);
nand UO_351 (O_351,N_2800,N_2987);
or UO_352 (O_352,N_2805,N_2869);
or UO_353 (O_353,N_2800,N_2961);
or UO_354 (O_354,N_2914,N_2937);
nand UO_355 (O_355,N_2967,N_2859);
xor UO_356 (O_356,N_2877,N_2808);
and UO_357 (O_357,N_2949,N_2865);
nor UO_358 (O_358,N_2907,N_2956);
nand UO_359 (O_359,N_2993,N_2896);
nor UO_360 (O_360,N_2905,N_2931);
and UO_361 (O_361,N_2809,N_2942);
nor UO_362 (O_362,N_2954,N_2952);
and UO_363 (O_363,N_2929,N_2932);
and UO_364 (O_364,N_2871,N_2934);
xor UO_365 (O_365,N_2932,N_2834);
and UO_366 (O_366,N_2996,N_2938);
and UO_367 (O_367,N_2974,N_2806);
nor UO_368 (O_368,N_2950,N_2812);
nand UO_369 (O_369,N_2882,N_2929);
nor UO_370 (O_370,N_2957,N_2925);
or UO_371 (O_371,N_2854,N_2942);
xor UO_372 (O_372,N_2880,N_2974);
nor UO_373 (O_373,N_2808,N_2886);
nor UO_374 (O_374,N_2843,N_2874);
and UO_375 (O_375,N_2960,N_2969);
nor UO_376 (O_376,N_2846,N_2905);
nor UO_377 (O_377,N_2806,N_2849);
nor UO_378 (O_378,N_2806,N_2952);
or UO_379 (O_379,N_2840,N_2842);
xor UO_380 (O_380,N_2968,N_2971);
or UO_381 (O_381,N_2824,N_2809);
or UO_382 (O_382,N_2984,N_2989);
nand UO_383 (O_383,N_2882,N_2802);
or UO_384 (O_384,N_2897,N_2893);
and UO_385 (O_385,N_2867,N_2869);
nand UO_386 (O_386,N_2820,N_2878);
and UO_387 (O_387,N_2816,N_2915);
and UO_388 (O_388,N_2983,N_2994);
nor UO_389 (O_389,N_2937,N_2845);
nand UO_390 (O_390,N_2923,N_2860);
or UO_391 (O_391,N_2820,N_2842);
nand UO_392 (O_392,N_2891,N_2961);
xnor UO_393 (O_393,N_2999,N_2973);
xnor UO_394 (O_394,N_2817,N_2982);
and UO_395 (O_395,N_2831,N_2936);
nor UO_396 (O_396,N_2905,N_2887);
nor UO_397 (O_397,N_2873,N_2851);
nor UO_398 (O_398,N_2859,N_2819);
or UO_399 (O_399,N_2921,N_2823);
nand UO_400 (O_400,N_2863,N_2842);
nand UO_401 (O_401,N_2920,N_2934);
and UO_402 (O_402,N_2941,N_2826);
or UO_403 (O_403,N_2804,N_2888);
xnor UO_404 (O_404,N_2913,N_2883);
and UO_405 (O_405,N_2851,N_2836);
xnor UO_406 (O_406,N_2922,N_2819);
nand UO_407 (O_407,N_2907,N_2903);
nor UO_408 (O_408,N_2877,N_2815);
nor UO_409 (O_409,N_2939,N_2971);
or UO_410 (O_410,N_2996,N_2949);
nor UO_411 (O_411,N_2830,N_2866);
nand UO_412 (O_412,N_2837,N_2832);
nand UO_413 (O_413,N_2895,N_2985);
nand UO_414 (O_414,N_2962,N_2866);
and UO_415 (O_415,N_2868,N_2829);
nor UO_416 (O_416,N_2940,N_2819);
and UO_417 (O_417,N_2987,N_2966);
and UO_418 (O_418,N_2826,N_2875);
or UO_419 (O_419,N_2915,N_2828);
or UO_420 (O_420,N_2816,N_2812);
or UO_421 (O_421,N_2941,N_2812);
nor UO_422 (O_422,N_2969,N_2901);
nand UO_423 (O_423,N_2869,N_2874);
and UO_424 (O_424,N_2871,N_2961);
nand UO_425 (O_425,N_2996,N_2802);
nand UO_426 (O_426,N_2856,N_2807);
nor UO_427 (O_427,N_2832,N_2901);
or UO_428 (O_428,N_2802,N_2888);
nand UO_429 (O_429,N_2943,N_2885);
or UO_430 (O_430,N_2986,N_2812);
and UO_431 (O_431,N_2996,N_2821);
nand UO_432 (O_432,N_2980,N_2812);
or UO_433 (O_433,N_2820,N_2857);
and UO_434 (O_434,N_2832,N_2919);
nor UO_435 (O_435,N_2991,N_2834);
and UO_436 (O_436,N_2864,N_2826);
nand UO_437 (O_437,N_2887,N_2975);
nand UO_438 (O_438,N_2929,N_2818);
or UO_439 (O_439,N_2800,N_2893);
or UO_440 (O_440,N_2802,N_2800);
or UO_441 (O_441,N_2860,N_2831);
and UO_442 (O_442,N_2965,N_2837);
or UO_443 (O_443,N_2999,N_2987);
or UO_444 (O_444,N_2833,N_2855);
nand UO_445 (O_445,N_2974,N_2963);
or UO_446 (O_446,N_2908,N_2917);
nor UO_447 (O_447,N_2939,N_2839);
nor UO_448 (O_448,N_2843,N_2908);
nor UO_449 (O_449,N_2876,N_2932);
and UO_450 (O_450,N_2939,N_2995);
or UO_451 (O_451,N_2952,N_2915);
and UO_452 (O_452,N_2904,N_2824);
and UO_453 (O_453,N_2825,N_2956);
nor UO_454 (O_454,N_2967,N_2829);
xnor UO_455 (O_455,N_2944,N_2882);
nor UO_456 (O_456,N_2888,N_2815);
nor UO_457 (O_457,N_2854,N_2871);
or UO_458 (O_458,N_2858,N_2920);
and UO_459 (O_459,N_2975,N_2879);
or UO_460 (O_460,N_2962,N_2871);
and UO_461 (O_461,N_2865,N_2833);
nor UO_462 (O_462,N_2828,N_2883);
nor UO_463 (O_463,N_2929,N_2848);
nor UO_464 (O_464,N_2820,N_2898);
xnor UO_465 (O_465,N_2922,N_2866);
nor UO_466 (O_466,N_2901,N_2929);
nor UO_467 (O_467,N_2944,N_2998);
nor UO_468 (O_468,N_2981,N_2930);
nor UO_469 (O_469,N_2969,N_2810);
or UO_470 (O_470,N_2945,N_2918);
or UO_471 (O_471,N_2960,N_2818);
and UO_472 (O_472,N_2832,N_2899);
or UO_473 (O_473,N_2967,N_2836);
or UO_474 (O_474,N_2981,N_2893);
xnor UO_475 (O_475,N_2960,N_2913);
xor UO_476 (O_476,N_2963,N_2920);
xnor UO_477 (O_477,N_2801,N_2975);
xnor UO_478 (O_478,N_2801,N_2822);
and UO_479 (O_479,N_2946,N_2919);
nand UO_480 (O_480,N_2955,N_2873);
xor UO_481 (O_481,N_2866,N_2909);
nor UO_482 (O_482,N_2943,N_2909);
nand UO_483 (O_483,N_2814,N_2943);
or UO_484 (O_484,N_2828,N_2941);
or UO_485 (O_485,N_2965,N_2891);
and UO_486 (O_486,N_2910,N_2844);
and UO_487 (O_487,N_2906,N_2849);
or UO_488 (O_488,N_2828,N_2894);
or UO_489 (O_489,N_2870,N_2825);
or UO_490 (O_490,N_2985,N_2873);
or UO_491 (O_491,N_2957,N_2973);
xor UO_492 (O_492,N_2938,N_2965);
nand UO_493 (O_493,N_2895,N_2972);
nand UO_494 (O_494,N_2961,N_2957);
nand UO_495 (O_495,N_2925,N_2894);
nor UO_496 (O_496,N_2979,N_2929);
or UO_497 (O_497,N_2808,N_2874);
and UO_498 (O_498,N_2981,N_2816);
or UO_499 (O_499,N_2951,N_2965);
endmodule