module basic_1500_15000_2000_120_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1153,In_514);
xor U1 (N_1,In_1298,In_491);
or U2 (N_2,In_250,In_469);
xor U3 (N_3,In_1099,In_822);
xor U4 (N_4,In_972,In_1082);
xnor U5 (N_5,In_654,In_1268);
or U6 (N_6,In_1151,In_1025);
nor U7 (N_7,In_466,In_122);
xor U8 (N_8,In_370,In_1178);
nor U9 (N_9,In_618,In_869);
nor U10 (N_10,In_587,In_719);
or U11 (N_11,In_20,In_754);
xnor U12 (N_12,In_652,In_728);
nor U13 (N_13,In_148,In_190);
or U14 (N_14,In_264,In_211);
or U15 (N_15,In_1001,In_1220);
and U16 (N_16,In_1224,In_1282);
nand U17 (N_17,In_1048,In_276);
or U18 (N_18,In_546,In_1445);
and U19 (N_19,In_731,In_93);
nand U20 (N_20,In_156,In_794);
xor U21 (N_21,In_1402,In_207);
and U22 (N_22,In_146,In_1032);
nor U23 (N_23,In_477,In_675);
nand U24 (N_24,In_55,In_1364);
or U25 (N_25,In_1020,In_479);
nand U26 (N_26,In_116,In_159);
or U27 (N_27,In_134,In_259);
or U28 (N_28,In_1333,In_68);
and U29 (N_29,In_1129,In_298);
and U30 (N_30,In_953,In_164);
xor U31 (N_31,In_225,In_1334);
or U32 (N_32,In_1095,In_402);
nand U33 (N_33,In_829,In_13);
nor U34 (N_34,In_413,In_1269);
nor U35 (N_35,In_346,In_1258);
nor U36 (N_36,In_204,In_397);
xor U37 (N_37,In_228,In_559);
or U38 (N_38,In_896,In_305);
xor U39 (N_39,In_65,In_1492);
or U40 (N_40,In_1144,In_455);
xnor U41 (N_41,In_1302,In_100);
nand U42 (N_42,In_147,In_1218);
and U43 (N_43,In_169,In_806);
xor U44 (N_44,In_1011,In_783);
and U45 (N_45,In_565,In_846);
nor U46 (N_46,In_7,In_1311);
or U47 (N_47,In_932,In_10);
nand U48 (N_48,In_1076,In_1022);
nand U49 (N_49,In_336,In_1264);
xor U50 (N_50,In_18,In_762);
nor U51 (N_51,In_1132,In_103);
or U52 (N_52,In_1243,In_309);
nor U53 (N_53,In_805,In_838);
or U54 (N_54,In_649,In_1131);
xor U55 (N_55,In_179,In_1139);
nand U56 (N_56,In_620,In_784);
and U57 (N_57,In_1475,In_1351);
or U58 (N_58,In_934,In_258);
nor U59 (N_59,In_1013,In_1309);
or U60 (N_60,In_185,In_123);
xnor U61 (N_61,In_1394,In_1157);
or U62 (N_62,In_590,In_683);
nand U63 (N_63,In_102,In_1284);
and U64 (N_64,In_378,In_234);
or U65 (N_65,In_767,In_905);
nor U66 (N_66,In_448,In_1400);
xor U67 (N_67,In_700,In_1100);
xor U68 (N_68,In_308,In_903);
nand U69 (N_69,In_173,In_673);
nor U70 (N_70,In_129,In_271);
or U71 (N_71,In_394,In_873);
xnor U72 (N_72,In_1440,In_458);
or U73 (N_73,In_484,In_1241);
nand U74 (N_74,In_876,In_1225);
xnor U75 (N_75,In_1083,In_686);
or U76 (N_76,In_361,In_854);
xnor U77 (N_77,In_819,In_354);
and U78 (N_78,In_142,In_1398);
or U79 (N_79,In_1140,In_1372);
nor U80 (N_80,In_687,In_1156);
or U81 (N_81,In_1188,In_1433);
or U82 (N_82,In_1193,In_922);
and U83 (N_83,In_193,In_297);
xor U84 (N_84,In_752,In_1229);
nand U85 (N_85,In_760,In_1391);
or U86 (N_86,In_1421,In_320);
and U87 (N_87,In_301,In_918);
nand U88 (N_88,In_718,In_1273);
xnor U89 (N_89,In_1341,In_128);
nor U90 (N_90,In_1181,In_456);
or U91 (N_91,In_613,In_488);
nand U92 (N_92,In_1145,In_31);
or U93 (N_93,In_1033,In_81);
and U94 (N_94,In_1069,In_534);
and U95 (N_95,In_383,In_1327);
nor U96 (N_96,In_615,In_818);
nor U97 (N_97,In_280,In_1496);
and U98 (N_98,In_189,In_1194);
and U99 (N_99,In_1430,In_1190);
and U100 (N_100,In_715,In_1164);
or U101 (N_101,In_176,In_645);
and U102 (N_102,In_1245,In_847);
and U103 (N_103,In_586,In_1409);
nor U104 (N_104,In_1427,In_22);
nor U105 (N_105,In_1003,In_1036);
nor U106 (N_106,In_1169,In_461);
or U107 (N_107,In_1230,In_1465);
or U108 (N_108,In_303,In_1071);
and U109 (N_109,In_571,In_1425);
and U110 (N_110,In_1493,In_981);
or U111 (N_111,In_1010,In_746);
nand U112 (N_112,In_210,In_1210);
or U113 (N_113,In_524,In_1007);
nor U114 (N_114,In_338,In_509);
nand U115 (N_115,In_1175,In_622);
nor U116 (N_116,In_1466,In_262);
or U117 (N_117,In_37,In_294);
nand U118 (N_118,In_1166,In_1287);
xnor U119 (N_119,In_240,In_591);
xor U120 (N_120,In_892,In_403);
nand U121 (N_121,In_1081,In_826);
nand U122 (N_122,In_1205,In_243);
nor U123 (N_123,In_835,In_725);
or U124 (N_124,In_812,In_828);
nand U125 (N_125,In_1142,In_504);
xnor U126 (N_126,In_1317,In_412);
xor U127 (N_127,In_322,In_833);
and U128 (N_128,In_580,In_200);
nor U129 (N_129,In_520,In_328);
nor U130 (N_130,In_143,In_1461);
or U131 (N_131,In_499,In_1079);
and U132 (N_132,In_438,In_1395);
or U133 (N_133,In_732,In_741);
nand U134 (N_134,In_1328,N_62);
nor U135 (N_135,In_886,In_795);
and U136 (N_136,In_555,In_518);
xnor U137 (N_137,In_220,In_655);
xor U138 (N_138,In_542,N_85);
nor U139 (N_139,In_95,In_44);
xnor U140 (N_140,N_49,N_50);
xnor U141 (N_141,In_78,In_1426);
or U142 (N_142,In_744,In_417);
and U143 (N_143,In_1014,N_113);
xnor U144 (N_144,In_676,In_939);
nor U145 (N_145,In_1252,In_365);
and U146 (N_146,In_959,In_664);
nand U147 (N_147,In_115,N_116);
nand U148 (N_148,In_713,In_63);
and U149 (N_149,In_1000,In_1050);
nand U150 (N_150,In_1450,In_1452);
nand U151 (N_151,In_787,In_1247);
and U152 (N_152,In_6,In_1367);
xnor U153 (N_153,N_64,In_1113);
and U154 (N_154,In_678,N_81);
nand U155 (N_155,In_1111,In_607);
nand U156 (N_156,In_925,In_1172);
xnor U157 (N_157,In_647,In_895);
or U158 (N_158,In_1259,In_74);
and U159 (N_159,In_1349,In_1017);
and U160 (N_160,In_743,In_487);
and U161 (N_161,In_1057,In_1209);
or U162 (N_162,In_398,In_948);
nor U163 (N_163,In_1326,In_372);
xor U164 (N_164,In_1110,In_757);
and U165 (N_165,In_792,In_1217);
nand U166 (N_166,In_168,In_530);
nand U167 (N_167,In_29,N_0);
xnor U168 (N_168,In_1257,In_371);
nor U169 (N_169,N_69,In_1361);
nor U170 (N_170,In_334,In_685);
or U171 (N_171,In_203,In_19);
or U172 (N_172,In_340,In_138);
or U173 (N_173,In_317,N_7);
nand U174 (N_174,In_1385,In_381);
nor U175 (N_175,In_353,In_3);
and U176 (N_176,In_593,In_496);
and U177 (N_177,In_990,In_949);
or U178 (N_178,In_539,In_1215);
xor U179 (N_179,In_682,In_121);
and U180 (N_180,In_1293,In_1377);
nor U181 (N_181,N_22,In_126);
nor U182 (N_182,In_1,N_107);
and U183 (N_183,In_307,In_437);
nand U184 (N_184,In_804,In_526);
or U185 (N_185,In_118,In_9);
and U186 (N_186,In_1077,In_815);
nand U187 (N_187,In_473,In_1278);
nor U188 (N_188,In_942,In_1275);
nor U189 (N_189,In_908,In_135);
nor U190 (N_190,In_809,In_375);
nor U191 (N_191,N_4,In_1294);
and U192 (N_192,In_366,In_286);
nand U193 (N_193,In_766,In_1337);
nand U194 (N_194,In_1167,In_951);
or U195 (N_195,In_493,In_80);
or U196 (N_196,In_1468,In_1219);
and U197 (N_197,N_94,In_201);
nand U198 (N_198,In_849,In_527);
or U199 (N_199,In_306,In_82);
xnor U200 (N_200,In_1114,In_161);
nor U201 (N_201,In_941,In_299);
nor U202 (N_202,In_551,In_864);
xor U203 (N_203,N_84,In_246);
xor U204 (N_204,In_114,In_429);
nand U205 (N_205,In_1052,N_91);
and U206 (N_206,In_653,In_1488);
and U207 (N_207,In_763,In_119);
and U208 (N_208,In_523,In_58);
nand U209 (N_209,In_572,In_1420);
or U210 (N_210,In_411,In_1438);
or U211 (N_211,In_889,In_721);
nand U212 (N_212,In_1090,In_577);
nor U213 (N_213,In_1499,In_41);
nor U214 (N_214,In_1080,In_60);
nand U215 (N_215,In_1448,In_1141);
nand U216 (N_216,In_221,In_807);
nor U217 (N_217,In_658,In_104);
nor U218 (N_218,In_1116,In_266);
nor U219 (N_219,In_1335,In_127);
and U220 (N_220,In_634,In_1092);
nand U221 (N_221,In_1378,In_573);
or U222 (N_222,N_31,In_667);
nand U223 (N_223,In_450,In_1031);
and U224 (N_224,In_661,In_515);
xnor U225 (N_225,In_1306,In_242);
and U226 (N_226,In_1308,In_946);
nand U227 (N_227,In_474,In_1104);
nor U228 (N_228,In_773,In_933);
xor U229 (N_229,N_71,In_1256);
nand U230 (N_230,In_1254,In_871);
nor U231 (N_231,In_196,In_730);
nor U232 (N_232,In_960,In_130);
or U233 (N_233,In_1159,In_1271);
and U234 (N_234,In_916,In_772);
nand U235 (N_235,In_926,In_1304);
xor U236 (N_236,In_1118,In_629);
nor U237 (N_237,In_1418,In_395);
xor U238 (N_238,In_418,In_1449);
or U239 (N_239,In_1432,In_1383);
xor U240 (N_240,In_775,In_722);
nand U241 (N_241,In_1356,N_106);
or U242 (N_242,In_1348,In_409);
or U243 (N_243,In_106,In_950);
nand U244 (N_244,In_735,In_929);
nor U245 (N_245,In_1174,In_384);
or U246 (N_246,In_1086,In_602);
and U247 (N_247,In_1009,In_440);
or U248 (N_248,In_628,In_512);
and U249 (N_249,In_915,In_1212);
xnor U250 (N_250,In_1015,In_252);
and U251 (N_251,In_1312,In_594);
or U252 (N_252,N_156,In_811);
or U253 (N_253,In_475,In_1158);
nand U254 (N_254,In_316,In_98);
nor U255 (N_255,In_983,In_907);
or U256 (N_256,In_810,In_633);
nand U257 (N_257,In_902,In_837);
or U258 (N_258,N_112,In_556);
or U259 (N_259,In_677,In_1314);
nand U260 (N_260,In_1147,In_1442);
nand U261 (N_261,In_1018,In_938);
nand U262 (N_262,In_83,In_274);
and U263 (N_263,N_211,In_261);
xnor U264 (N_264,In_1486,In_1272);
nand U265 (N_265,In_231,In_786);
or U266 (N_266,In_842,In_25);
nand U267 (N_267,N_77,In_1125);
or U268 (N_268,In_637,In_1371);
or U269 (N_269,In_845,In_858);
and U270 (N_270,In_890,In_570);
or U271 (N_271,In_552,N_243);
nor U272 (N_272,In_690,In_603);
or U273 (N_273,In_356,In_1093);
nand U274 (N_274,In_1244,N_171);
nor U275 (N_275,In_643,N_42);
or U276 (N_276,In_608,In_780);
and U277 (N_277,N_56,In_610);
and U278 (N_278,In_1406,In_363);
nand U279 (N_279,In_1123,N_215);
and U280 (N_280,In_117,In_1060);
and U281 (N_281,In_1399,In_1105);
xnor U282 (N_282,In_335,In_1459);
xor U283 (N_283,In_1265,In_1183);
and U284 (N_284,In_583,In_49);
and U285 (N_285,In_1321,In_698);
or U286 (N_286,N_144,In_92);
nor U287 (N_287,N_123,In_1035);
and U288 (N_288,In_944,In_35);
nor U289 (N_289,In_714,In_597);
and U290 (N_290,N_138,In_21);
nand U291 (N_291,N_90,In_140);
or U292 (N_292,In_898,In_963);
and U293 (N_293,In_152,N_2);
nand U294 (N_294,In_879,In_1270);
and U295 (N_295,In_133,In_1061);
nand U296 (N_296,In_257,N_108);
xor U297 (N_297,In_368,N_75);
nor U298 (N_298,N_231,In_505);
or U299 (N_299,In_489,In_814);
and U300 (N_300,In_1323,In_436);
or U301 (N_301,In_575,N_222);
nor U302 (N_302,N_38,In_836);
xor U303 (N_303,N_76,In_1299);
nor U304 (N_304,N_210,N_100);
or U305 (N_305,In_498,In_1006);
xnor U306 (N_306,In_965,In_521);
nor U307 (N_307,In_566,N_79);
nand U308 (N_308,In_1390,In_471);
and U309 (N_309,In_592,In_43);
and U310 (N_310,N_213,N_217);
xnor U311 (N_311,In_840,In_1059);
nand U312 (N_312,In_1024,N_147);
and U313 (N_313,In_832,In_1133);
or U314 (N_314,In_33,In_1097);
xor U315 (N_315,N_89,In_1366);
nand U316 (N_316,In_1115,In_312);
or U317 (N_317,In_851,In_734);
nand U318 (N_318,In_45,In_171);
and U319 (N_319,In_163,N_247);
nand U320 (N_320,In_205,In_779);
nand U321 (N_321,In_1039,N_120);
nand U322 (N_322,N_186,In_973);
and U323 (N_323,In_359,In_1277);
or U324 (N_324,In_971,In_468);
or U325 (N_325,In_808,In_1091);
xor U326 (N_326,In_1297,In_285);
or U327 (N_327,N_128,In_52);
xnor U328 (N_328,In_222,In_663);
xnor U329 (N_329,In_1474,In_14);
and U330 (N_330,In_263,N_32);
or U331 (N_331,In_90,In_1191);
xor U332 (N_332,N_151,In_759);
and U333 (N_333,In_1227,N_18);
nand U334 (N_334,In_680,In_1384);
xor U335 (N_335,In_111,In_51);
and U336 (N_336,In_1417,In_860);
xnor U337 (N_337,In_444,In_727);
nand U338 (N_338,In_253,In_238);
nand U339 (N_339,N_1,N_207);
nor U340 (N_340,In_1480,In_1303);
and U341 (N_341,In_920,In_1292);
and U342 (N_342,N_61,N_114);
and U343 (N_343,In_549,In_332);
and U344 (N_344,In_416,In_789);
or U345 (N_345,In_1439,In_1016);
nand U346 (N_346,In_209,In_961);
or U347 (N_347,N_11,In_289);
xor U348 (N_348,N_238,In_689);
nor U349 (N_349,In_958,In_674);
nand U350 (N_350,In_1063,In_1495);
xor U351 (N_351,In_1376,In_318);
nand U352 (N_352,In_668,In_1414);
and U353 (N_353,In_1246,In_12);
and U354 (N_354,In_962,In_994);
nor U355 (N_355,N_40,In_564);
and U356 (N_356,N_46,In_563);
xnor U357 (N_357,In_707,In_226);
nand U358 (N_358,In_349,N_239);
nand U359 (N_359,In_186,In_265);
xor U360 (N_360,N_216,In_1030);
or U361 (N_361,In_998,In_66);
xnor U362 (N_362,In_1038,In_576);
nand U363 (N_363,In_1049,N_166);
and U364 (N_364,N_19,N_233);
or U365 (N_365,N_70,In_358);
xnor U366 (N_366,In_940,In_476);
nor U367 (N_367,In_1332,N_33);
or U368 (N_368,In_883,N_45);
nand U369 (N_369,In_342,In_1162);
and U370 (N_370,In_921,N_199);
or U371 (N_371,In_296,In_778);
nor U372 (N_372,In_904,In_155);
nand U373 (N_373,N_93,In_600);
nand U374 (N_374,In_1261,N_21);
nand U375 (N_375,In_192,N_260);
and U376 (N_376,N_347,N_55);
nand U377 (N_377,In_1434,In_1074);
xnor U378 (N_378,In_1248,In_1481);
nand U379 (N_379,In_414,In_268);
or U380 (N_380,N_92,In_53);
or U381 (N_381,In_1324,In_1460);
nor U382 (N_382,N_34,N_311);
nor U383 (N_383,In_39,In_1435);
and U384 (N_384,In_292,N_230);
and U385 (N_385,In_646,N_264);
and U386 (N_386,In_914,In_327);
or U387 (N_387,In_0,In_84);
and U388 (N_388,N_68,In_701);
and U389 (N_389,N_328,In_287);
nor U390 (N_390,In_89,In_431);
nand U391 (N_391,In_1149,In_34);
xnor U392 (N_392,In_233,In_439);
or U393 (N_393,N_259,In_671);
or U394 (N_394,In_445,In_1109);
and U395 (N_395,In_1165,In_1029);
nor U396 (N_396,In_1410,N_117);
or U397 (N_397,N_150,In_183);
nor U398 (N_398,In_1026,In_433);
and U399 (N_399,N_188,In_1331);
and U400 (N_400,In_868,In_877);
and U401 (N_401,In_1128,N_195);
xor U402 (N_402,In_753,In_30);
and U403 (N_403,In_379,N_327);
nor U404 (N_404,In_230,In_401);
xnor U405 (N_405,In_1476,In_1008);
nor U406 (N_406,In_880,In_955);
xnor U407 (N_407,In_1479,In_1424);
or U408 (N_408,In_1301,N_221);
nand U409 (N_409,N_160,In_295);
or U410 (N_410,In_279,In_40);
nand U411 (N_411,In_350,In_373);
and U412 (N_412,In_1281,N_372);
nor U413 (N_413,In_691,In_470);
xor U414 (N_414,In_139,In_1455);
xnor U415 (N_415,In_936,N_290);
and U416 (N_416,In_393,In_1161);
or U417 (N_417,In_1373,In_856);
or U418 (N_418,In_170,In_1358);
xor U419 (N_419,In_1042,N_110);
and U420 (N_420,In_314,In_151);
nand U421 (N_421,In_87,In_641);
and U422 (N_422,In_777,N_127);
nand U423 (N_423,N_262,In_1407);
nand U424 (N_424,N_284,In_382);
nor U425 (N_425,In_823,N_170);
nor U426 (N_426,N_252,In_723);
or U427 (N_427,In_717,In_1005);
nand U428 (N_428,N_28,In_1375);
xor U429 (N_429,N_88,In_1267);
or U430 (N_430,In_1340,N_334);
nand U431 (N_431,In_75,N_78);
and U432 (N_432,N_339,In_1472);
nand U433 (N_433,N_303,In_545);
nor U434 (N_434,N_344,In_11);
nand U435 (N_435,In_463,N_336);
xnor U436 (N_436,In_913,N_245);
nand U437 (N_437,In_584,N_299);
nand U438 (N_438,In_931,In_852);
nand U439 (N_439,In_162,In_1211);
nand U440 (N_440,In_333,N_118);
xor U441 (N_441,In_1451,N_39);
nand U442 (N_442,N_96,In_799);
nand U443 (N_443,In_1473,In_300);
or U444 (N_444,In_884,In_141);
nor U445 (N_445,In_976,In_219);
nand U446 (N_446,In_213,In_748);
nor U447 (N_447,In_1397,N_300);
or U448 (N_448,In_987,N_346);
or U449 (N_449,In_270,In_107);
xnor U450 (N_450,In_331,In_1365);
xor U451 (N_451,In_227,N_25);
nand U452 (N_452,In_400,In_1396);
and U453 (N_453,N_340,In_540);
nor U454 (N_454,N_155,N_149);
or U455 (N_455,N_99,In_323);
nand U456 (N_456,In_1054,In_785);
xnor U457 (N_457,In_132,N_366);
xor U458 (N_458,In_181,In_178);
or U459 (N_459,In_765,In_648);
nand U460 (N_460,In_313,N_20);
and U461 (N_461,In_831,N_318);
xnor U462 (N_462,In_267,In_761);
nand U463 (N_463,In_1386,In_1198);
xnor U464 (N_464,N_219,In_467);
and U465 (N_465,In_642,N_240);
xor U466 (N_466,In_348,In_1249);
and U467 (N_467,N_298,In_59);
nand U468 (N_468,In_459,In_670);
nand U469 (N_469,N_183,N_270);
xnor U470 (N_470,In_195,In_1200);
nand U471 (N_471,In_578,N_133);
nor U472 (N_472,In_404,In_1088);
nand U473 (N_473,In_462,N_57);
xor U474 (N_474,In_1345,In_442);
nor U475 (N_475,N_129,In_351);
nor U476 (N_476,In_1250,In_216);
nand U477 (N_477,In_969,In_405);
or U478 (N_478,In_153,In_867);
nand U479 (N_479,In_1041,In_255);
or U480 (N_480,In_1416,In_109);
nand U481 (N_481,N_200,In_1235);
or U482 (N_482,In_339,In_755);
or U483 (N_483,N_321,In_64);
nand U484 (N_484,In_954,In_517);
or U485 (N_485,In_165,In_17);
xor U486 (N_486,In_232,In_1168);
or U487 (N_487,N_162,N_98);
nand U488 (N_488,In_432,In_560);
nand U489 (N_489,N_235,In_702);
nand U490 (N_490,In_1431,In_711);
or U491 (N_491,In_167,In_202);
or U492 (N_492,In_1320,In_704);
nand U493 (N_493,In_1160,In_321);
and U494 (N_494,In_325,In_672);
nor U495 (N_495,In_105,In_749);
and U496 (N_496,In_1401,In_605);
nor U497 (N_497,N_175,In_218);
xor U498 (N_498,In_745,In_1313);
and U499 (N_499,In_1405,In_197);
nor U500 (N_500,N_192,In_574);
nor U501 (N_501,In_606,N_329);
nor U502 (N_502,In_235,In_1369);
nand U503 (N_503,N_146,N_208);
nor U504 (N_504,N_24,In_1073);
xor U505 (N_505,N_60,In_770);
and U506 (N_506,In_736,In_1187);
or U507 (N_507,In_1392,In_588);
or U508 (N_508,In_61,N_442);
xnor U509 (N_509,In_579,In_1223);
xnor U510 (N_510,In_1286,In_595);
and U511 (N_511,In_891,N_445);
nor U512 (N_512,In_1477,In_71);
nor U513 (N_513,In_324,N_422);
xor U514 (N_514,In_507,In_516);
nand U515 (N_515,N_206,N_27);
nor U516 (N_516,In_930,N_393);
nand U517 (N_517,In_791,N_286);
xnor U518 (N_518,In_1360,In_175);
nor U519 (N_519,In_1240,In_739);
or U520 (N_520,In_73,In_1199);
nor U521 (N_521,In_999,In_1154);
nor U522 (N_522,In_326,In_1089);
xor U523 (N_523,In_793,N_410);
or U524 (N_524,In_94,N_495);
and U525 (N_525,In_329,In_32);
nand U526 (N_526,In_1350,N_212);
nor U527 (N_527,N_296,N_457);
and U528 (N_528,In_1279,In_697);
or U529 (N_529,N_381,In_154);
and U530 (N_530,In_885,N_378);
xnor U531 (N_531,N_464,In_1290);
and U532 (N_532,In_979,In_1437);
nor U533 (N_533,N_325,N_470);
nor U534 (N_534,N_281,N_400);
xor U535 (N_535,In_589,In_1467);
and U536 (N_536,N_320,In_1180);
nand U537 (N_537,N_452,N_261);
and U538 (N_538,In_239,N_363);
xor U539 (N_539,In_750,N_242);
nand U540 (N_540,In_251,In_501);
and U541 (N_541,N_278,In_710);
nor U542 (N_542,In_1056,In_859);
or U543 (N_543,N_354,In_212);
and U544 (N_544,N_295,N_225);
or U545 (N_545,N_185,N_310);
xor U546 (N_546,N_271,In_928);
xnor U547 (N_547,In_269,N_388);
and U548 (N_548,In_621,N_44);
xnor U549 (N_549,In_131,In_1478);
or U550 (N_550,N_267,N_164);
xor U551 (N_551,In_991,In_457);
or U552 (N_552,In_345,In_424);
nand U553 (N_553,In_1415,N_283);
xnor U554 (N_554,N_244,In_1216);
xor U555 (N_555,In_149,In_1260);
or U556 (N_556,N_480,In_1491);
nor U557 (N_557,In_443,In_968);
or U558 (N_558,In_453,In_1138);
nor U559 (N_559,In_1428,In_69);
nand U560 (N_560,In_1120,In_1464);
or U561 (N_561,In_273,N_35);
nand U562 (N_562,In_1127,In_893);
nand U563 (N_563,N_36,In_1315);
nor U564 (N_564,N_135,In_1487);
nor U565 (N_565,In_1055,In_347);
nand U566 (N_566,N_418,In_482);
xor U567 (N_567,In_839,In_86);
or U568 (N_568,In_709,In_460);
and U569 (N_569,N_424,In_428);
nand U570 (N_570,In_427,N_269);
or U571 (N_571,In_781,In_611);
xnor U572 (N_572,In_535,In_364);
or U573 (N_573,N_438,In_391);
xnor U574 (N_574,N_172,In_900);
or U575 (N_575,In_1288,In_1186);
nand U576 (N_576,N_288,In_76);
xnor U577 (N_577,N_343,In_1023);
and U578 (N_578,N_37,In_901);
nor U579 (N_579,In_330,N_83);
or U580 (N_580,In_820,N_437);
and U581 (N_581,In_769,N_483);
and U582 (N_582,N_158,In_626);
nor U583 (N_583,In_585,In_1047);
xnor U584 (N_584,In_729,In_472);
xor U585 (N_585,In_882,N_458);
or U586 (N_586,In_581,N_414);
xnor U587 (N_587,N_292,In_875);
nor U588 (N_588,In_237,N_429);
nor U589 (N_589,N_430,In_124);
nor U590 (N_590,In_706,In_1253);
and U591 (N_591,In_1204,N_74);
nor U592 (N_592,In_277,In_343);
xnor U593 (N_593,In_97,In_157);
nor U594 (N_594,In_452,N_126);
or U595 (N_595,N_391,N_349);
nand U596 (N_596,N_370,N_130);
xor U597 (N_597,N_481,In_802);
xor U598 (N_598,N_258,In_341);
nand U599 (N_599,In_862,In_260);
nand U600 (N_600,In_88,N_23);
or U601 (N_601,In_927,In_1339);
nor U602 (N_602,In_311,N_73);
xnor U603 (N_603,N_308,In_848);
or U604 (N_604,In_844,In_878);
nor U605 (N_605,In_604,In_26);
nand U606 (N_606,N_229,In_492);
nand U607 (N_607,N_291,N_53);
nand U608 (N_608,N_364,In_249);
nand U609 (N_609,In_813,In_695);
and U610 (N_610,N_80,N_473);
nand U611 (N_611,In_62,N_468);
and U612 (N_612,In_8,N_397);
or U613 (N_613,In_906,N_279);
and U614 (N_614,N_479,N_141);
xnor U615 (N_615,N_122,In_304);
nor U616 (N_616,In_1040,N_392);
nand U617 (N_617,N_312,In_1213);
xor U618 (N_618,N_494,In_1300);
xnor U619 (N_619,N_365,In_1148);
nor U620 (N_620,N_371,In_1353);
xnor U621 (N_621,In_110,In_217);
nand U622 (N_622,N_373,N_478);
and U623 (N_623,In_275,N_41);
and U624 (N_624,In_974,N_189);
or U625 (N_625,In_380,N_237);
nor U626 (N_626,In_1354,In_389);
nand U627 (N_627,In_989,N_273);
and U628 (N_628,In_1182,N_256);
nand U629 (N_629,In_419,In_1126);
and U630 (N_630,In_150,In_1316);
xor U631 (N_631,In_1085,N_482);
xor U632 (N_632,N_459,N_181);
nand U633 (N_633,N_178,N_228);
nand U634 (N_634,In_1346,In_1359);
or U635 (N_635,In_1196,N_305);
nor U636 (N_636,In_1490,In_47);
and U637 (N_637,N_167,N_377);
or U638 (N_638,N_331,N_168);
or U639 (N_639,In_1471,N_622);
and U640 (N_640,In_1102,N_275);
nand U641 (N_641,In_911,In_1363);
xor U642 (N_642,In_790,N_157);
nor U643 (N_643,N_599,N_220);
or U644 (N_644,In_978,N_454);
or U645 (N_645,N_236,In_1108);
nor U646 (N_646,In_1489,In_223);
nor U647 (N_647,N_379,N_426);
and U648 (N_648,In_272,In_1135);
or U649 (N_649,In_1236,In_1497);
nand U650 (N_650,N_348,In_774);
nand U651 (N_651,N_597,In_747);
nand U652 (N_652,In_1336,N_567);
and U653 (N_653,In_396,N_335);
and U654 (N_654,In_1285,N_169);
xor U655 (N_655,In_627,N_30);
or U656 (N_656,In_1441,In_733);
nand U657 (N_657,N_619,In_282);
nand U658 (N_658,N_460,In_1347);
xnor U659 (N_659,In_481,N_399);
and U660 (N_660,In_1028,N_10);
and U661 (N_661,In_1098,In_614);
and U662 (N_662,In_1289,N_578);
nand U663 (N_663,In_843,In_48);
nand U664 (N_664,N_405,N_203);
or U665 (N_665,N_505,N_601);
or U666 (N_666,In_797,In_742);
or U667 (N_667,N_582,In_631);
nand U668 (N_668,N_154,In_137);
and U669 (N_669,In_1357,In_206);
and U670 (N_670,In_554,In_1381);
nor U671 (N_671,In_187,In_693);
and U672 (N_672,In_1185,In_705);
and U673 (N_673,In_870,In_977);
nand U674 (N_674,N_255,N_466);
nand U675 (N_675,N_427,In_1155);
nor U676 (N_676,N_12,In_410);
nor U677 (N_677,In_422,In_1206);
or U678 (N_678,In_1101,N_115);
nand U679 (N_679,In_23,In_1498);
nor U680 (N_680,In_101,N_179);
or U681 (N_681,N_226,N_274);
and U682 (N_682,N_585,N_304);
and U683 (N_683,In_247,N_605);
and U684 (N_684,In_174,N_608);
and U685 (N_685,N_249,N_15);
and U686 (N_686,In_758,N_173);
and U687 (N_687,In_659,In_367);
or U688 (N_688,N_485,In_1403);
nand U689 (N_689,N_374,N_276);
or U690 (N_690,In_42,In_120);
xor U691 (N_691,N_584,In_992);
xnor U692 (N_692,In_598,In_975);
or U693 (N_693,In_855,In_553);
xnor U694 (N_694,In_360,In_194);
xor U695 (N_695,N_234,In_408);
or U696 (N_696,N_176,N_534);
xnor U697 (N_697,N_367,In_1058);
nand U698 (N_698,N_294,N_326);
or U699 (N_699,N_491,In_522);
nor U700 (N_700,In_688,In_1344);
or U701 (N_701,N_125,N_148);
nand U702 (N_702,In_543,In_290);
nand U703 (N_703,N_48,In_525);
xnor U704 (N_704,N_502,In_782);
xnor U705 (N_705,N_5,In_756);
nand U706 (N_706,N_82,In_957);
or U707 (N_707,N_152,N_520);
nand U708 (N_708,N_499,N_59);
and U709 (N_709,In_986,In_937);
xor U710 (N_710,N_496,N_561);
nor U711 (N_711,N_9,In_866);
and U712 (N_712,In_1422,N_14);
and U713 (N_713,N_433,In_740);
nor U714 (N_714,In_1043,N_518);
or U715 (N_715,In_1233,In_800);
nand U716 (N_716,In_1117,N_47);
nor U717 (N_717,N_194,N_517);
nand U718 (N_718,In_635,N_431);
or U719 (N_719,In_1456,In_224);
or U720 (N_720,In_465,In_256);
xor U721 (N_721,N_620,In_319);
nand U722 (N_722,N_511,N_111);
nand U723 (N_723,N_493,N_359);
xnor U724 (N_724,In_984,In_863);
or U725 (N_725,N_432,N_415);
nor U726 (N_726,N_87,N_306);
nor U727 (N_727,N_409,N_263);
and U728 (N_728,N_202,In_1202);
and U729 (N_729,In_1112,N_436);
nor U730 (N_730,N_3,In_2);
nor U731 (N_731,N_184,N_515);
nand U732 (N_732,In_1189,In_712);
nand U733 (N_733,In_1062,N_412);
and U734 (N_734,N_557,In_861);
nand U735 (N_735,N_214,N_248);
nor U736 (N_736,In_660,In_214);
nor U737 (N_737,In_38,In_1355);
xor U738 (N_738,N_280,N_309);
or U739 (N_739,In_980,N_564);
xor U740 (N_740,N_560,N_142);
or U741 (N_741,N_467,N_501);
and U742 (N_742,N_223,In_344);
nand U743 (N_743,N_97,In_538);
nor U744 (N_744,N_317,In_352);
xor U745 (N_745,N_587,In_1280);
xnor U746 (N_746,In_1274,N_182);
nand U747 (N_747,In_1121,N_516);
nor U748 (N_748,In_1067,In_708);
nor U749 (N_749,In_1170,N_227);
or U750 (N_750,N_610,N_440);
xnor U751 (N_751,In_1343,In_966);
and U752 (N_752,N_562,In_125);
or U753 (N_753,In_1084,In_426);
xnor U754 (N_754,N_209,N_16);
nor U755 (N_755,N_497,In_912);
nor U756 (N_756,In_281,N_568);
nand U757 (N_757,In_1064,N_655);
and U758 (N_758,N_742,In_816);
or U759 (N_759,N_549,N_319);
and U760 (N_760,In_454,In_1429);
or U761 (N_761,N_537,N_419);
nor U762 (N_762,In_215,In_1307);
or U763 (N_763,In_1380,N_352);
and U764 (N_764,In_982,N_682);
nor U765 (N_765,N_333,N_692);
xnor U766 (N_766,In_993,In_1352);
xor U767 (N_767,In_1469,In_1137);
nor U768 (N_768,In_1179,N_523);
and U769 (N_769,N_205,N_598);
and U770 (N_770,N_361,In_446);
and U771 (N_771,N_193,N_103);
xnor U772 (N_772,N_729,N_621);
and U773 (N_773,In_768,In_1119);
or U774 (N_774,N_639,N_246);
and U775 (N_775,N_736,N_699);
xor U776 (N_776,In_434,In_636);
or U777 (N_777,In_1107,In_1176);
and U778 (N_778,N_661,N_553);
and U779 (N_779,In_624,N_132);
and U780 (N_780,In_684,N_580);
nor U781 (N_781,N_615,N_664);
nor U782 (N_782,N_66,N_648);
nand U783 (N_783,In_337,In_1004);
nand U784 (N_784,N_686,N_119);
xnor U785 (N_785,In_1412,In_657);
or U786 (N_786,N_554,N_688);
nor U787 (N_787,In_387,N_250);
nor U788 (N_788,N_428,In_1457);
xor U789 (N_789,N_201,N_576);
or U790 (N_790,N_708,N_488);
or U791 (N_791,N_384,In_441);
or U792 (N_792,N_555,N_532);
nor U793 (N_793,N_724,In_166);
and U794 (N_794,N_421,N_625);
and U795 (N_795,In_737,In_1065);
or U796 (N_796,N_735,N_659);
nand U797 (N_797,N_538,N_423);
nand U798 (N_798,In_399,In_1239);
xnor U799 (N_799,In_1046,In_716);
xnor U800 (N_800,N_647,In_548);
nor U801 (N_801,In_430,In_1173);
or U802 (N_802,N_471,In_632);
nor U803 (N_803,In_1305,In_1214);
or U804 (N_804,N_86,In_390);
xnor U805 (N_805,N_282,N_741);
and U806 (N_806,In_1171,In_536);
xnor U807 (N_807,In_865,N_498);
and U808 (N_808,N_611,In_485);
nand U809 (N_809,In_544,N_330);
or U810 (N_810,N_606,In_1291);
or U811 (N_811,In_464,In_1484);
or U812 (N_812,N_671,In_245);
nand U813 (N_813,In_1404,In_964);
xnor U814 (N_814,In_798,N_590);
xor U815 (N_815,In_1152,N_508);
or U816 (N_816,In_550,N_600);
or U817 (N_817,N_633,N_663);
and U818 (N_818,In_1045,In_1318);
xnor U819 (N_819,In_1226,N_696);
nor U820 (N_820,N_342,N_43);
nor U821 (N_821,N_588,In_478);
xor U822 (N_822,In_1379,N_657);
and U823 (N_823,N_642,In_995);
nand U824 (N_824,In_897,In_1087);
xnor U825 (N_825,In_532,In_494);
and U826 (N_826,In_1338,N_707);
and U827 (N_827,In_490,N_652);
nor U828 (N_828,N_500,N_572);
nor U829 (N_829,N_302,In_952);
nand U830 (N_830,N_701,In_28);
or U831 (N_831,In_547,In_640);
and U832 (N_832,N_187,In_887);
nor U833 (N_833,N_137,N_17);
and U834 (N_834,N_738,N_6);
and U835 (N_835,N_583,In_623);
nand U836 (N_836,N_434,In_850);
and U837 (N_837,N_717,N_574);
nand U838 (N_838,N_533,N_743);
nand U839 (N_839,N_65,In_392);
and U840 (N_840,N_265,In_894);
nand U841 (N_841,N_643,In_208);
xnor U842 (N_842,In_27,In_1096);
and U843 (N_843,N_713,N_632);
and U844 (N_844,In_46,N_631);
nor U845 (N_845,In_541,N_541);
nor U846 (N_846,In_449,In_248);
or U847 (N_847,In_619,In_970);
or U848 (N_848,N_301,N_586);
and U849 (N_849,N_623,In_15);
or U850 (N_850,N_559,N_51);
nand U851 (N_851,N_104,In_1150);
nor U852 (N_852,In_751,N_272);
nand U853 (N_853,N_737,In_284);
nor U854 (N_854,In_67,N_477);
nand U855 (N_855,N_649,N_672);
xor U856 (N_856,N_139,N_629);
xor U857 (N_857,In_1197,N_566);
nand U858 (N_858,N_548,N_638);
xor U859 (N_859,In_945,N_700);
nor U860 (N_860,N_604,N_29);
nor U861 (N_861,N_232,In_1221);
nand U862 (N_862,In_596,In_997);
xor U863 (N_863,In_1124,In_1094);
nor U864 (N_864,In_24,In_771);
xor U865 (N_865,N_720,In_528);
or U866 (N_866,N_131,N_640);
or U867 (N_867,N_287,N_727);
and U868 (N_868,In_537,N_704);
xnor U869 (N_869,N_540,In_283);
nor U870 (N_870,N_730,N_413);
nand U871 (N_871,In_1368,N_161);
nand U872 (N_872,N_662,In_377);
xor U873 (N_873,N_218,N_636);
nand U874 (N_874,N_524,N_407);
and U875 (N_875,In_956,In_188);
xnor U876 (N_876,In_1012,In_108);
xnor U877 (N_877,In_1362,In_803);
or U878 (N_878,In_692,N_703);
or U879 (N_879,N_866,N_709);
nor U880 (N_880,N_812,N_474);
nor U881 (N_881,In_1184,N_776);
nor U882 (N_882,N_544,N_492);
nand U883 (N_883,N_577,N_358);
and U884 (N_884,N_277,In_899);
nor U885 (N_885,N_140,In_1002);
and U886 (N_886,N_761,N_396);
and U887 (N_887,N_627,In_1207);
nand U888 (N_888,In_177,In_315);
nor U889 (N_889,In_1462,In_724);
and U890 (N_890,N_832,N_674);
or U891 (N_891,In_1136,N_26);
xnor U892 (N_892,N_803,N_487);
xnor U893 (N_893,In_1389,In_738);
nand U894 (N_894,In_1342,In_796);
and U895 (N_895,In_244,N_375);
or U896 (N_896,In_531,N_385);
nand U897 (N_897,In_502,N_792);
or U898 (N_898,N_801,N_596);
xnor U899 (N_899,In_1027,N_617);
or U900 (N_900,In_1228,In_609);
and U901 (N_901,In_1419,N_775);
and U902 (N_902,In_1262,N_472);
and U903 (N_903,N_289,N_448);
or U904 (N_904,In_357,In_435);
and U905 (N_905,N_689,N_241);
nand U906 (N_906,In_198,In_644);
xor U907 (N_907,N_522,N_777);
or U908 (N_908,In_1446,N_360);
and U909 (N_909,N_833,N_716);
and U910 (N_910,N_749,In_1237);
nand U911 (N_911,N_824,In_776);
or U912 (N_912,N_844,N_747);
nand U913 (N_913,N_771,N_780);
nor U914 (N_914,N_594,In_1325);
nand U915 (N_915,N_507,N_563);
or U916 (N_916,N_644,In_113);
nand U917 (N_917,In_310,In_1037);
and U918 (N_918,In_451,In_420);
nor U919 (N_919,N_102,In_1393);
and U920 (N_920,N_796,N_441);
nand U921 (N_921,N_859,In_669);
nor U922 (N_922,N_355,In_415);
and U923 (N_923,N_63,N_867);
and U924 (N_924,In_666,In_1122);
nand U925 (N_925,N_368,N_536);
nor U926 (N_926,In_1106,In_1388);
nand U927 (N_927,N_718,N_871);
nor U928 (N_928,N_543,In_888);
nor U929 (N_929,N_855,In_726);
or U930 (N_930,In_924,N_769);
nor U931 (N_931,N_791,N_854);
nand U932 (N_932,N_745,N_751);
and U933 (N_933,N_710,N_726);
xnor U934 (N_934,N_545,In_423);
nand U935 (N_935,In_788,N_817);
nand U936 (N_936,N_788,In_54);
or U937 (N_937,N_687,N_253);
nand U938 (N_938,N_313,N_733);
and U939 (N_939,N_752,N_630);
nand U940 (N_940,N_679,N_180);
nor U941 (N_941,N_853,N_637);
and U942 (N_942,In_355,In_72);
xor U943 (N_943,N_174,N_351);
nand U944 (N_944,In_720,N_772);
and U945 (N_945,N_846,N_697);
or U946 (N_946,In_158,In_236);
nand U947 (N_947,N_322,In_1413);
and U948 (N_948,N_257,N_658);
nand U949 (N_949,In_625,In_529);
and U950 (N_950,In_681,N_475);
and U951 (N_951,N_865,In_70);
xor U952 (N_952,In_1453,N_569);
and U953 (N_953,In_1066,N_756);
xor U954 (N_954,N_109,N_754);
nand U955 (N_955,N_874,N_589);
and U956 (N_956,N_764,In_558);
nor U957 (N_957,N_197,In_1044);
nor U958 (N_958,In_824,N_465);
nand U959 (N_959,N_635,N_618);
xnor U960 (N_960,N_163,In_1411);
or U961 (N_961,N_849,In_639);
nor U962 (N_962,In_1436,In_699);
or U963 (N_963,In_425,In_386);
or U964 (N_964,N_711,In_696);
nor U965 (N_965,In_182,In_1053);
nor U966 (N_966,N_13,N_607);
xor U967 (N_967,N_525,In_1078);
xnor U968 (N_968,N_748,N_739);
xnor U969 (N_969,In_985,N_356);
xor U970 (N_970,N_750,N_417);
or U971 (N_971,N_852,N_105);
nand U972 (N_972,N_857,In_909);
xor U973 (N_973,N_834,In_1485);
xnor U974 (N_974,In_1322,N_469);
or U975 (N_975,In_519,In_144);
nor U976 (N_976,In_1458,N_556);
and U977 (N_977,N_695,N_683);
xnor U978 (N_978,N_451,N_760);
and U979 (N_979,N_869,N_705);
and U980 (N_980,In_881,N_136);
nand U981 (N_981,N_667,In_57);
nor U982 (N_982,In_1329,N_612);
and U983 (N_983,N_251,In_1021);
and U984 (N_984,N_830,N_847);
xor U985 (N_985,In_1374,N_676);
xor U986 (N_986,N_721,N_822);
nand U987 (N_987,N_159,N_616);
and U988 (N_988,In_191,In_172);
or U989 (N_989,N_864,In_1447);
xor U990 (N_990,In_1283,N_529);
nand U991 (N_991,N_565,N_840);
xor U992 (N_992,In_947,N_678);
nor U993 (N_993,N_490,N_425);
xnor U994 (N_994,N_758,N_539);
nor U995 (N_995,In_96,In_1034);
or U996 (N_996,In_4,In_362);
or U997 (N_997,N_702,N_394);
nor U998 (N_998,N_268,N_8);
or U999 (N_999,In_503,N_453);
nor U1000 (N_1000,N_933,N_337);
nor U1001 (N_1001,N_972,N_862);
or U1002 (N_1002,N_506,N_573);
xor U1003 (N_1003,In_510,N_919);
and U1004 (N_1004,N_911,In_77);
or U1005 (N_1005,N_967,N_794);
and U1006 (N_1006,N_602,N_836);
xnor U1007 (N_1007,N_907,N_285);
xnor U1008 (N_1008,N_974,N_930);
nand U1009 (N_1009,N_786,N_654);
or U1010 (N_1010,N_550,N_153);
xor U1011 (N_1011,N_858,N_793);
xnor U1012 (N_1012,N_134,N_798);
xnor U1013 (N_1013,N_592,N_953);
and U1014 (N_1014,N_935,N_839);
or U1015 (N_1015,In_85,N_902);
and U1016 (N_1016,N_819,N_814);
nor U1017 (N_1017,N_677,N_759);
nand U1018 (N_1018,N_825,N_634);
and U1019 (N_1019,In_612,N_324);
xnor U1020 (N_1020,N_946,N_691);
nand U1021 (N_1021,N_401,In_1068);
nor U1022 (N_1022,N_797,In_630);
nor U1023 (N_1023,N_893,N_811);
nand U1024 (N_1024,N_673,In_1494);
or U1025 (N_1025,In_872,In_1310);
and U1026 (N_1026,In_1051,In_910);
or U1027 (N_1027,N_781,N_443);
nor U1028 (N_1028,N_552,N_787);
xor U1029 (N_1029,In_1192,N_821);
or U1030 (N_1030,N_316,In_1130);
xnor U1031 (N_1031,N_904,N_975);
nor U1032 (N_1032,In_293,N_341);
and U1033 (N_1033,N_357,In_923);
nor U1034 (N_1034,N_446,In_486);
nor U1035 (N_1035,N_693,N_961);
and U1036 (N_1036,In_1370,N_991);
nand U1037 (N_1037,N_850,N_762);
nand U1038 (N_1038,In_406,N_338);
or U1039 (N_1039,N_571,N_404);
xnor U1040 (N_1040,N_928,N_723);
and U1041 (N_1041,N_143,N_684);
nor U1042 (N_1042,In_1222,In_241);
xor U1043 (N_1043,N_996,In_679);
nand U1044 (N_1044,N_712,N_783);
and U1045 (N_1045,N_909,N_362);
nand U1046 (N_1046,N_997,In_199);
nand U1047 (N_1047,N_595,N_765);
or U1048 (N_1048,N_121,N_389);
and U1049 (N_1049,N_614,N_963);
nor U1050 (N_1050,N_945,N_818);
or U1051 (N_1051,In_369,N_528);
xor U1052 (N_1052,N_350,N_675);
nor U1053 (N_1053,In_1203,In_254);
xor U1054 (N_1054,N_806,N_929);
and U1055 (N_1055,N_680,N_753);
and U1056 (N_1056,N_802,N_646);
xnor U1057 (N_1057,N_992,N_734);
and U1058 (N_1058,In_1208,N_345);
nand U1059 (N_1059,N_987,N_435);
nor U1060 (N_1060,N_921,N_486);
xnor U1061 (N_1061,In_919,N_641);
or U1062 (N_1062,N_983,N_837);
xnor U1063 (N_1063,N_462,N_732);
xnor U1064 (N_1064,N_936,N_519);
nand U1065 (N_1065,In_184,N_913);
or U1066 (N_1066,N_145,N_484);
or U1067 (N_1067,N_804,In_302);
or U1068 (N_1068,N_690,N_978);
nor U1069 (N_1069,N_884,N_789);
nor U1070 (N_1070,N_899,N_959);
xnor U1071 (N_1071,N_944,N_456);
nor U1072 (N_1072,N_509,N_224);
xnor U1073 (N_1073,N_873,N_503);
and U1074 (N_1074,N_934,In_561);
nor U1075 (N_1075,N_740,N_694);
or U1076 (N_1076,N_960,N_897);
and U1077 (N_1077,In_1444,N_903);
and U1078 (N_1078,N_353,N_942);
or U1079 (N_1079,In_569,N_845);
nor U1080 (N_1080,N_810,N_581);
xnor U1081 (N_1081,N_514,N_757);
and U1082 (N_1082,N_912,N_950);
and U1083 (N_1083,In_1482,In_1330);
and U1084 (N_1084,In_1295,N_593);
xnor U1085 (N_1085,N_746,In_662);
and U1086 (N_1086,N_398,N_842);
and U1087 (N_1087,N_755,N_900);
or U1088 (N_1088,N_315,In_99);
nor U1089 (N_1089,N_332,N_624);
or U1090 (N_1090,N_547,In_1382);
and U1091 (N_1091,N_922,N_917);
nor U1092 (N_1092,N_861,N_785);
nor U1093 (N_1093,In_1072,N_665);
or U1094 (N_1094,N_823,N_535);
or U1095 (N_1095,N_603,N_863);
xnor U1096 (N_1096,N_957,In_650);
nand U1097 (N_1097,In_506,N_820);
xnor U1098 (N_1098,N_925,In_582);
nand U1099 (N_1099,N_725,N_376);
nand U1100 (N_1100,N_773,N_976);
nor U1101 (N_1101,N_895,In_967);
nor U1102 (N_1102,In_374,N_489);
nor U1103 (N_1103,N_843,In_801);
nor U1104 (N_1104,N_931,In_1143);
or U1105 (N_1105,N_886,In_1195);
nor U1106 (N_1106,In_1255,In_601);
xor U1107 (N_1107,N_254,N_406);
nand U1108 (N_1108,In_1146,In_483);
nand U1109 (N_1109,In_56,N_681);
nor U1110 (N_1110,In_694,N_570);
or U1111 (N_1111,In_1238,N_990);
and U1112 (N_1112,N_513,In_1163);
xnor U1113 (N_1113,N_790,N_651);
nor U1114 (N_1114,In_853,N_941);
or U1115 (N_1115,N_728,N_954);
and U1116 (N_1116,In_160,N_970);
or U1117 (N_1117,N_191,N_980);
nor U1118 (N_1118,N_715,N_952);
nand U1119 (N_1119,In_508,N_878);
and U1120 (N_1120,N_977,N_198);
nand U1121 (N_1121,N_964,N_981);
xnor U1122 (N_1122,In_145,In_665);
nor U1123 (N_1123,In_16,N_851);
xnor U1124 (N_1124,N_766,N_190);
or U1125 (N_1125,N_1007,N_1105);
nor U1126 (N_1126,N_1001,N_905);
nor U1127 (N_1127,N_910,In_557);
and U1128 (N_1128,N_1016,N_95);
xor U1129 (N_1129,N_124,In_500);
nand U1130 (N_1130,N_875,N_1117);
or U1131 (N_1131,N_1011,N_993);
or U1132 (N_1132,N_390,N_880);
xnor U1133 (N_1133,In_1408,N_656);
nand U1134 (N_1134,N_955,In_825);
and U1135 (N_1135,N_591,N_626);
nand U1136 (N_1136,N_891,N_965);
nand U1137 (N_1137,N_660,N_888);
or U1138 (N_1138,N_1102,In_385);
and U1139 (N_1139,N_1110,N_889);
or U1140 (N_1140,N_476,N_1108);
nand U1141 (N_1141,N_1065,N_731);
nor U1142 (N_1142,N_1088,N_1003);
nand U1143 (N_1143,N_940,N_1036);
nor U1144 (N_1144,N_204,N_827);
nand U1145 (N_1145,N_1020,N_763);
and U1146 (N_1146,N_1033,N_1069);
xnor U1147 (N_1147,N_971,N_885);
and U1148 (N_1148,In_638,N_314);
xor U1149 (N_1149,N_896,N_1055);
xor U1150 (N_1150,N_416,N_1101);
nand U1151 (N_1151,In_407,In_841);
or U1152 (N_1152,N_1090,N_504);
and U1153 (N_1153,N_1100,N_1045);
or U1154 (N_1154,In_599,N_1025);
nand U1155 (N_1155,N_1053,N_1059);
nor U1156 (N_1156,In_1177,N_72);
and U1157 (N_1157,N_898,N_795);
nor U1158 (N_1158,N_1037,In_917);
nand U1159 (N_1159,N_883,N_444);
xnor U1160 (N_1160,N_461,N_609);
and U1161 (N_1161,N_1062,N_1091);
or U1162 (N_1162,N_1082,In_1443);
or U1163 (N_1163,N_799,N_685);
and U1164 (N_1164,N_1005,N_915);
nand U1165 (N_1165,N_1081,N_807);
nor U1166 (N_1166,In_112,N_542);
or U1167 (N_1167,In_616,N_949);
xnor U1168 (N_1168,N_669,N_58);
xnor U1169 (N_1169,N_877,N_1122);
and U1170 (N_1170,N_449,N_531);
nand U1171 (N_1171,In_229,N_1123);
xor U1172 (N_1172,N_1073,N_323);
nand U1173 (N_1173,N_1095,N_808);
nand U1174 (N_1174,N_382,N_628);
or U1175 (N_1175,In_1423,N_653);
and U1176 (N_1176,In_857,N_876);
nand U1177 (N_1177,N_1019,In_562);
and U1178 (N_1178,In_1075,N_1089);
nor U1179 (N_1179,N_968,N_927);
or U1180 (N_1180,N_768,N_714);
or U1181 (N_1181,In_1251,N_882);
xor U1182 (N_1182,N_988,N_266);
and U1183 (N_1183,N_1018,N_1056);
and U1184 (N_1184,In_1276,N_1014);
xor U1185 (N_1185,In_497,N_439);
and U1186 (N_1186,N_1121,N_1047);
xnor U1187 (N_1187,N_879,In_50);
and U1188 (N_1188,In_278,N_307);
xnor U1189 (N_1189,N_1046,N_948);
or U1190 (N_1190,N_1060,N_1028);
and U1191 (N_1191,N_923,N_1077);
nand U1192 (N_1192,In_180,In_447);
or U1193 (N_1193,N_813,N_1035);
nor U1194 (N_1194,N_1039,N_926);
nor U1195 (N_1195,N_1083,N_1087);
or U1196 (N_1196,In_513,N_575);
nand U1197 (N_1197,In_1463,N_579);
xor U1198 (N_1198,N_829,N_939);
and U1199 (N_1199,N_848,In_1232);
nand U1200 (N_1200,N_924,N_838);
xnor U1201 (N_1201,N_958,N_860);
nand U1202 (N_1202,N_1048,N_670);
nand U1203 (N_1203,N_1058,N_984);
or U1204 (N_1204,In_1070,N_1093);
nor U1205 (N_1205,N_1104,N_1043);
xor U1206 (N_1206,N_870,N_982);
nor U1207 (N_1207,N_744,N_979);
and U1208 (N_1208,N_1099,N_784);
or U1209 (N_1209,N_1012,In_703);
xor U1210 (N_1210,N_908,N_521);
xnor U1211 (N_1211,N_196,N_998);
nor U1212 (N_1212,In_1134,N_779);
and U1213 (N_1213,N_1071,N_1098);
xnor U1214 (N_1214,N_856,N_1031);
xor U1215 (N_1215,N_1006,In_830);
and U1216 (N_1216,N_774,N_386);
xnor U1217 (N_1217,N_1076,In_1103);
and U1218 (N_1218,In_1019,N_293);
or U1219 (N_1219,In_817,N_1116);
nor U1220 (N_1220,In_1231,In_79);
xor U1221 (N_1221,N_1040,N_1109);
or U1222 (N_1222,N_369,N_986);
nand U1223 (N_1223,In_996,In_1470);
nand U1224 (N_1224,In_376,N_512);
nand U1225 (N_1225,N_1017,N_916);
or U1226 (N_1226,N_297,N_1074);
xnor U1227 (N_1227,N_890,N_1124);
or U1228 (N_1228,N_951,N_1067);
or U1229 (N_1229,N_1111,N_892);
and U1230 (N_1230,N_408,In_1201);
xnor U1231 (N_1231,N_1118,In_567);
and U1232 (N_1232,In_988,N_1008);
or U1233 (N_1233,N_613,N_938);
nand U1234 (N_1234,N_932,N_767);
nor U1235 (N_1235,In_651,In_495);
nand U1236 (N_1236,N_666,N_706);
and U1237 (N_1237,N_558,In_1454);
and U1238 (N_1238,N_650,N_901);
nand U1239 (N_1239,N_1106,N_177);
xnor U1240 (N_1240,N_947,N_1119);
nor U1241 (N_1241,In_568,N_937);
and U1242 (N_1242,N_956,N_815);
nor U1243 (N_1243,In_421,N_1084);
nand U1244 (N_1244,N_411,In_1263);
or U1245 (N_1245,N_1038,N_828);
or U1246 (N_1246,N_1096,N_989);
nor U1247 (N_1247,N_1044,In_656);
nand U1248 (N_1248,N_395,N_1054);
nand U1249 (N_1249,In_834,In_821);
or U1250 (N_1250,N_809,N_1128);
and U1251 (N_1251,In_874,N_1237);
nand U1252 (N_1252,N_1161,N_1185);
nor U1253 (N_1253,In_1242,N_914);
and U1254 (N_1254,N_1156,N_1176);
nand U1255 (N_1255,N_52,N_1114);
xor U1256 (N_1256,N_920,N_1203);
xor U1257 (N_1257,N_1245,N_1080);
xnor U1258 (N_1258,N_1009,N_1248);
and U1259 (N_1259,N_1216,N_1032);
nand U1260 (N_1260,N_1224,N_1192);
xnor U1261 (N_1261,N_1079,N_1097);
xnor U1262 (N_1262,In_1483,In_288);
or U1263 (N_1263,N_510,N_1230);
and U1264 (N_1264,N_999,N_1193);
and U1265 (N_1265,N_1160,N_1198);
and U1266 (N_1266,N_826,N_546);
xor U1267 (N_1267,N_1175,N_383);
or U1268 (N_1268,In_91,N_1139);
nand U1269 (N_1269,N_966,N_1143);
nand U1270 (N_1270,N_1194,N_1120);
nand U1271 (N_1271,N_1042,N_1092);
or U1272 (N_1272,N_1182,N_1165);
and U1273 (N_1273,N_1241,N_770);
or U1274 (N_1274,In_1234,N_1004);
and U1275 (N_1275,N_1236,N_1146);
and U1276 (N_1276,N_1243,N_1141);
or U1277 (N_1277,N_1112,In_1266);
nor U1278 (N_1278,N_1240,N_1162);
nand U1279 (N_1279,N_719,In_388);
nor U1280 (N_1280,N_1187,In_1296);
xor U1281 (N_1281,N_1221,N_1177);
or U1282 (N_1282,N_1228,N_841);
or U1283 (N_1283,N_1196,N_450);
nor U1284 (N_1284,N_1179,N_668);
nand U1285 (N_1285,N_1075,N_1225);
nor U1286 (N_1286,N_887,N_1041);
and U1287 (N_1287,N_1142,N_403);
and U1288 (N_1288,N_1068,N_1158);
xor U1289 (N_1289,N_1219,N_1132);
nand U1290 (N_1290,N_872,N_969);
nand U1291 (N_1291,N_1234,N_1178);
xnor U1292 (N_1292,N_835,N_1205);
xnor U1293 (N_1293,N_1051,N_1029);
or U1294 (N_1294,N_1078,N_1061);
nand U1295 (N_1295,N_1227,N_1222);
xor U1296 (N_1296,N_1147,N_1170);
xnor U1297 (N_1297,N_1206,N_1244);
or U1298 (N_1298,N_994,N_1167);
xor U1299 (N_1299,In_533,In_5);
and U1300 (N_1300,N_1201,N_1214);
or U1301 (N_1301,N_1024,N_1235);
nand U1302 (N_1302,N_1163,N_1034);
xnor U1303 (N_1303,N_1013,N_1223);
xnor U1304 (N_1304,N_420,In_136);
xor U1305 (N_1305,N_1151,N_868);
xor U1306 (N_1306,N_1173,N_380);
and U1307 (N_1307,N_1188,N_1207);
xnor U1308 (N_1308,N_1233,N_1231);
or U1309 (N_1309,N_985,N_1202);
and U1310 (N_1310,N_1213,N_1021);
xor U1311 (N_1311,N_1057,N_962);
xnor U1312 (N_1312,N_1180,N_67);
xnor U1313 (N_1313,N_1218,N_1166);
nor U1314 (N_1314,N_1115,N_805);
or U1315 (N_1315,N_1149,N_1140);
nand U1316 (N_1316,N_831,N_1215);
or U1317 (N_1317,N_455,N_1131);
or U1318 (N_1318,N_1152,N_1086);
nand U1319 (N_1319,N_1211,In_617);
and U1320 (N_1320,In_1319,N_1107);
and U1321 (N_1321,N_943,N_463);
nor U1322 (N_1322,N_1150,N_1154);
and U1323 (N_1323,N_527,N_1052);
or U1324 (N_1324,N_1125,N_645);
or U1325 (N_1325,N_800,N_1226);
and U1326 (N_1326,N_1200,In_935);
or U1327 (N_1327,N_1050,N_1094);
or U1328 (N_1328,N_1072,N_1186);
and U1329 (N_1329,N_1148,N_1030);
and U1330 (N_1330,N_526,N_1195);
or U1331 (N_1331,N_1103,N_1210);
nand U1332 (N_1332,N_1066,N_1168);
nand U1333 (N_1333,N_816,N_1212);
and U1334 (N_1334,N_1208,N_1063);
xor U1335 (N_1335,N_881,N_551);
nand U1336 (N_1336,N_165,N_1064);
nand U1337 (N_1337,N_1183,N_1153);
nor U1338 (N_1338,N_101,N_918);
xor U1339 (N_1339,N_1027,N_1209);
xnor U1340 (N_1340,N_1133,N_1164);
nand U1341 (N_1341,N_1189,N_1190);
nor U1342 (N_1342,N_1238,N_1002);
nor U1343 (N_1343,N_1113,N_1136);
and U1344 (N_1344,N_1000,N_1204);
or U1345 (N_1345,N_1184,N_1134);
nor U1346 (N_1346,N_1239,N_1242);
xor U1347 (N_1347,N_1217,N_1169);
xnor U1348 (N_1348,N_1127,N_1247);
nand U1349 (N_1349,N_1191,N_1085);
and U1350 (N_1350,N_1144,N_1137);
or U1351 (N_1351,In_36,N_1172);
nor U1352 (N_1352,N_1126,N_1220);
or U1353 (N_1353,N_1129,N_1010);
or U1354 (N_1354,N_54,N_530);
nor U1355 (N_1355,N_1159,N_1171);
or U1356 (N_1356,N_402,In_1387);
xnor U1357 (N_1357,N_1181,N_1049);
nand U1358 (N_1358,In_480,N_1174);
nor U1359 (N_1359,N_1249,N_722);
nand U1360 (N_1360,In_764,N_894);
nand U1361 (N_1361,N_447,N_1246);
or U1362 (N_1362,In_943,N_1015);
nor U1363 (N_1363,N_1138,N_1229);
and U1364 (N_1364,N_995,N_1023);
nor U1365 (N_1365,N_1197,N_778);
xor U1366 (N_1366,N_387,In_291);
xor U1367 (N_1367,N_973,N_1135);
and U1368 (N_1368,N_1130,N_1155);
and U1369 (N_1369,In_511,N_698);
xnor U1370 (N_1370,N_1026,N_1232);
xnor U1371 (N_1371,N_1157,N_1199);
nand U1372 (N_1372,N_782,N_1070);
or U1373 (N_1373,N_1145,N_906);
or U1374 (N_1374,In_827,N_1022);
nor U1375 (N_1375,N_1345,N_1310);
xor U1376 (N_1376,N_1305,N_1291);
or U1377 (N_1377,N_1263,N_1318);
nor U1378 (N_1378,N_1299,N_1368);
nor U1379 (N_1379,N_1272,N_1326);
or U1380 (N_1380,N_1269,N_1265);
nor U1381 (N_1381,N_1302,N_1324);
or U1382 (N_1382,N_1282,N_1301);
nor U1383 (N_1383,N_1293,N_1297);
and U1384 (N_1384,N_1338,N_1335);
nand U1385 (N_1385,N_1333,N_1268);
and U1386 (N_1386,N_1309,N_1270);
nand U1387 (N_1387,N_1294,N_1349);
nor U1388 (N_1388,N_1279,N_1350);
nor U1389 (N_1389,N_1277,N_1300);
nand U1390 (N_1390,N_1348,N_1353);
or U1391 (N_1391,N_1339,N_1303);
nand U1392 (N_1392,N_1330,N_1374);
nand U1393 (N_1393,N_1355,N_1253);
or U1394 (N_1394,N_1284,N_1273);
and U1395 (N_1395,N_1357,N_1316);
and U1396 (N_1396,N_1288,N_1295);
nor U1397 (N_1397,N_1271,N_1281);
nand U1398 (N_1398,N_1364,N_1278);
nor U1399 (N_1399,N_1343,N_1358);
and U1400 (N_1400,N_1274,N_1256);
and U1401 (N_1401,N_1369,N_1275);
and U1402 (N_1402,N_1262,N_1306);
nand U1403 (N_1403,N_1367,N_1311);
and U1404 (N_1404,N_1313,N_1250);
nor U1405 (N_1405,N_1362,N_1354);
and U1406 (N_1406,N_1312,N_1258);
nor U1407 (N_1407,N_1259,N_1261);
xor U1408 (N_1408,N_1337,N_1283);
or U1409 (N_1409,N_1257,N_1356);
nand U1410 (N_1410,N_1327,N_1361);
xnor U1411 (N_1411,N_1292,N_1359);
or U1412 (N_1412,N_1370,N_1317);
or U1413 (N_1413,N_1314,N_1342);
xnor U1414 (N_1414,N_1307,N_1267);
xor U1415 (N_1415,N_1373,N_1344);
and U1416 (N_1416,N_1308,N_1336);
nand U1417 (N_1417,N_1266,N_1315);
and U1418 (N_1418,N_1365,N_1319);
nand U1419 (N_1419,N_1351,N_1304);
nand U1420 (N_1420,N_1280,N_1322);
xnor U1421 (N_1421,N_1352,N_1346);
or U1422 (N_1422,N_1334,N_1341);
nand U1423 (N_1423,N_1252,N_1290);
or U1424 (N_1424,N_1251,N_1372);
nor U1425 (N_1425,N_1260,N_1320);
and U1426 (N_1426,N_1289,N_1298);
and U1427 (N_1427,N_1285,N_1254);
or U1428 (N_1428,N_1332,N_1255);
xnor U1429 (N_1429,N_1360,N_1371);
nand U1430 (N_1430,N_1321,N_1323);
xnor U1431 (N_1431,N_1329,N_1296);
or U1432 (N_1432,N_1276,N_1331);
nor U1433 (N_1433,N_1287,N_1340);
nor U1434 (N_1434,N_1325,N_1328);
and U1435 (N_1435,N_1366,N_1264);
nand U1436 (N_1436,N_1347,N_1363);
nand U1437 (N_1437,N_1286,N_1332);
xnor U1438 (N_1438,N_1274,N_1312);
nand U1439 (N_1439,N_1360,N_1292);
nor U1440 (N_1440,N_1261,N_1341);
nand U1441 (N_1441,N_1279,N_1364);
and U1442 (N_1442,N_1310,N_1281);
and U1443 (N_1443,N_1279,N_1323);
nand U1444 (N_1444,N_1309,N_1264);
nor U1445 (N_1445,N_1334,N_1357);
nor U1446 (N_1446,N_1281,N_1276);
and U1447 (N_1447,N_1373,N_1358);
and U1448 (N_1448,N_1331,N_1299);
xnor U1449 (N_1449,N_1326,N_1369);
or U1450 (N_1450,N_1282,N_1332);
nand U1451 (N_1451,N_1336,N_1307);
or U1452 (N_1452,N_1268,N_1355);
or U1453 (N_1453,N_1282,N_1295);
nor U1454 (N_1454,N_1360,N_1354);
or U1455 (N_1455,N_1284,N_1372);
xnor U1456 (N_1456,N_1360,N_1257);
nand U1457 (N_1457,N_1311,N_1278);
xor U1458 (N_1458,N_1370,N_1250);
or U1459 (N_1459,N_1269,N_1281);
and U1460 (N_1460,N_1296,N_1259);
nand U1461 (N_1461,N_1359,N_1309);
xor U1462 (N_1462,N_1295,N_1305);
xor U1463 (N_1463,N_1263,N_1250);
and U1464 (N_1464,N_1326,N_1261);
or U1465 (N_1465,N_1271,N_1371);
and U1466 (N_1466,N_1316,N_1299);
or U1467 (N_1467,N_1306,N_1348);
nor U1468 (N_1468,N_1361,N_1254);
nand U1469 (N_1469,N_1282,N_1327);
nand U1470 (N_1470,N_1360,N_1337);
or U1471 (N_1471,N_1355,N_1363);
or U1472 (N_1472,N_1276,N_1349);
and U1473 (N_1473,N_1334,N_1355);
and U1474 (N_1474,N_1284,N_1289);
and U1475 (N_1475,N_1359,N_1302);
and U1476 (N_1476,N_1282,N_1255);
and U1477 (N_1477,N_1301,N_1281);
and U1478 (N_1478,N_1372,N_1265);
nand U1479 (N_1479,N_1334,N_1343);
and U1480 (N_1480,N_1260,N_1322);
and U1481 (N_1481,N_1262,N_1298);
nor U1482 (N_1482,N_1339,N_1257);
nand U1483 (N_1483,N_1265,N_1336);
nand U1484 (N_1484,N_1339,N_1373);
nand U1485 (N_1485,N_1308,N_1337);
or U1486 (N_1486,N_1301,N_1368);
xnor U1487 (N_1487,N_1262,N_1320);
xnor U1488 (N_1488,N_1367,N_1261);
xnor U1489 (N_1489,N_1339,N_1259);
xnor U1490 (N_1490,N_1335,N_1269);
or U1491 (N_1491,N_1368,N_1359);
nand U1492 (N_1492,N_1278,N_1332);
and U1493 (N_1493,N_1374,N_1250);
and U1494 (N_1494,N_1355,N_1316);
nand U1495 (N_1495,N_1252,N_1256);
nand U1496 (N_1496,N_1371,N_1311);
and U1497 (N_1497,N_1308,N_1317);
nand U1498 (N_1498,N_1254,N_1266);
and U1499 (N_1499,N_1338,N_1255);
nor U1500 (N_1500,N_1487,N_1466);
xnor U1501 (N_1501,N_1428,N_1398);
and U1502 (N_1502,N_1380,N_1495);
or U1503 (N_1503,N_1378,N_1381);
or U1504 (N_1504,N_1409,N_1471);
nor U1505 (N_1505,N_1403,N_1469);
or U1506 (N_1506,N_1486,N_1436);
and U1507 (N_1507,N_1411,N_1439);
nor U1508 (N_1508,N_1431,N_1413);
and U1509 (N_1509,N_1451,N_1489);
xor U1510 (N_1510,N_1477,N_1414);
or U1511 (N_1511,N_1400,N_1499);
or U1512 (N_1512,N_1449,N_1440);
nor U1513 (N_1513,N_1425,N_1459);
nand U1514 (N_1514,N_1438,N_1401);
nand U1515 (N_1515,N_1422,N_1404);
and U1516 (N_1516,N_1375,N_1435);
or U1517 (N_1517,N_1393,N_1391);
nor U1518 (N_1518,N_1498,N_1458);
nand U1519 (N_1519,N_1397,N_1441);
nand U1520 (N_1520,N_1427,N_1483);
xnor U1521 (N_1521,N_1389,N_1454);
nor U1522 (N_1522,N_1446,N_1452);
nand U1523 (N_1523,N_1415,N_1388);
or U1524 (N_1524,N_1384,N_1470);
xnor U1525 (N_1525,N_1417,N_1426);
and U1526 (N_1526,N_1416,N_1410);
nand U1527 (N_1527,N_1450,N_1464);
xnor U1528 (N_1528,N_1432,N_1394);
and U1529 (N_1529,N_1424,N_1396);
and U1530 (N_1530,N_1395,N_1379);
xnor U1531 (N_1531,N_1376,N_1443);
xnor U1532 (N_1532,N_1484,N_1488);
nor U1533 (N_1533,N_1387,N_1497);
nand U1534 (N_1534,N_1453,N_1455);
and U1535 (N_1535,N_1399,N_1406);
nor U1536 (N_1536,N_1481,N_1480);
xor U1537 (N_1537,N_1468,N_1460);
or U1538 (N_1538,N_1493,N_1437);
and U1539 (N_1539,N_1474,N_1448);
nand U1540 (N_1540,N_1476,N_1402);
nand U1541 (N_1541,N_1478,N_1482);
nor U1542 (N_1542,N_1479,N_1492);
nand U1543 (N_1543,N_1423,N_1473);
nand U1544 (N_1544,N_1385,N_1465);
nand U1545 (N_1545,N_1485,N_1472);
and U1546 (N_1546,N_1457,N_1491);
and U1547 (N_1547,N_1445,N_1419);
or U1548 (N_1548,N_1390,N_1463);
xor U1549 (N_1549,N_1418,N_1377);
or U1550 (N_1550,N_1447,N_1494);
nand U1551 (N_1551,N_1434,N_1405);
or U1552 (N_1552,N_1475,N_1496);
xor U1553 (N_1553,N_1382,N_1412);
xor U1554 (N_1554,N_1407,N_1490);
and U1555 (N_1555,N_1442,N_1456);
or U1556 (N_1556,N_1461,N_1467);
and U1557 (N_1557,N_1420,N_1430);
or U1558 (N_1558,N_1421,N_1386);
xnor U1559 (N_1559,N_1462,N_1433);
nor U1560 (N_1560,N_1408,N_1429);
and U1561 (N_1561,N_1392,N_1383);
and U1562 (N_1562,N_1444,N_1406);
nor U1563 (N_1563,N_1459,N_1493);
xnor U1564 (N_1564,N_1458,N_1454);
nand U1565 (N_1565,N_1499,N_1450);
or U1566 (N_1566,N_1468,N_1379);
or U1567 (N_1567,N_1452,N_1380);
nor U1568 (N_1568,N_1401,N_1376);
or U1569 (N_1569,N_1487,N_1380);
xnor U1570 (N_1570,N_1497,N_1419);
xnor U1571 (N_1571,N_1447,N_1406);
nand U1572 (N_1572,N_1454,N_1481);
xnor U1573 (N_1573,N_1409,N_1497);
or U1574 (N_1574,N_1418,N_1441);
and U1575 (N_1575,N_1424,N_1497);
or U1576 (N_1576,N_1387,N_1421);
nor U1577 (N_1577,N_1427,N_1448);
and U1578 (N_1578,N_1381,N_1469);
or U1579 (N_1579,N_1413,N_1424);
nor U1580 (N_1580,N_1429,N_1468);
nand U1581 (N_1581,N_1483,N_1408);
nand U1582 (N_1582,N_1422,N_1424);
nor U1583 (N_1583,N_1425,N_1452);
xor U1584 (N_1584,N_1439,N_1486);
xor U1585 (N_1585,N_1450,N_1385);
or U1586 (N_1586,N_1423,N_1483);
nor U1587 (N_1587,N_1491,N_1447);
xor U1588 (N_1588,N_1449,N_1469);
nor U1589 (N_1589,N_1399,N_1430);
nand U1590 (N_1590,N_1414,N_1438);
xor U1591 (N_1591,N_1461,N_1407);
nor U1592 (N_1592,N_1451,N_1383);
nand U1593 (N_1593,N_1439,N_1399);
xnor U1594 (N_1594,N_1495,N_1479);
xor U1595 (N_1595,N_1426,N_1467);
nand U1596 (N_1596,N_1379,N_1418);
and U1597 (N_1597,N_1457,N_1432);
nor U1598 (N_1598,N_1410,N_1419);
and U1599 (N_1599,N_1478,N_1457);
and U1600 (N_1600,N_1377,N_1498);
or U1601 (N_1601,N_1474,N_1449);
nor U1602 (N_1602,N_1448,N_1431);
or U1603 (N_1603,N_1491,N_1464);
or U1604 (N_1604,N_1382,N_1421);
or U1605 (N_1605,N_1423,N_1389);
xnor U1606 (N_1606,N_1493,N_1441);
xnor U1607 (N_1607,N_1483,N_1410);
nand U1608 (N_1608,N_1456,N_1459);
nor U1609 (N_1609,N_1489,N_1446);
or U1610 (N_1610,N_1396,N_1459);
or U1611 (N_1611,N_1463,N_1399);
nor U1612 (N_1612,N_1458,N_1406);
and U1613 (N_1613,N_1385,N_1443);
xor U1614 (N_1614,N_1478,N_1460);
or U1615 (N_1615,N_1435,N_1482);
or U1616 (N_1616,N_1486,N_1480);
nand U1617 (N_1617,N_1479,N_1387);
or U1618 (N_1618,N_1397,N_1477);
nor U1619 (N_1619,N_1435,N_1405);
nand U1620 (N_1620,N_1377,N_1463);
nand U1621 (N_1621,N_1394,N_1429);
nor U1622 (N_1622,N_1382,N_1426);
nor U1623 (N_1623,N_1389,N_1434);
xnor U1624 (N_1624,N_1381,N_1432);
xnor U1625 (N_1625,N_1513,N_1571);
or U1626 (N_1626,N_1525,N_1558);
nor U1627 (N_1627,N_1579,N_1545);
xor U1628 (N_1628,N_1538,N_1501);
or U1629 (N_1629,N_1605,N_1606);
xor U1630 (N_1630,N_1512,N_1618);
or U1631 (N_1631,N_1603,N_1516);
and U1632 (N_1632,N_1622,N_1546);
nor U1633 (N_1633,N_1540,N_1612);
and U1634 (N_1634,N_1541,N_1511);
xor U1635 (N_1635,N_1562,N_1569);
xnor U1636 (N_1636,N_1535,N_1598);
and U1637 (N_1637,N_1514,N_1506);
xor U1638 (N_1638,N_1608,N_1578);
nor U1639 (N_1639,N_1509,N_1537);
nand U1640 (N_1640,N_1566,N_1533);
xnor U1641 (N_1641,N_1576,N_1522);
and U1642 (N_1642,N_1609,N_1549);
nor U1643 (N_1643,N_1568,N_1543);
nand U1644 (N_1644,N_1610,N_1584);
nand U1645 (N_1645,N_1583,N_1559);
nand U1646 (N_1646,N_1515,N_1620);
nand U1647 (N_1647,N_1539,N_1553);
nand U1648 (N_1648,N_1532,N_1586);
nand U1649 (N_1649,N_1526,N_1611);
nand U1650 (N_1650,N_1548,N_1534);
nor U1651 (N_1651,N_1556,N_1616);
nor U1652 (N_1652,N_1504,N_1527);
nand U1653 (N_1653,N_1563,N_1574);
nor U1654 (N_1654,N_1589,N_1524);
and U1655 (N_1655,N_1623,N_1575);
and U1656 (N_1656,N_1502,N_1555);
or U1657 (N_1657,N_1594,N_1518);
xnor U1658 (N_1658,N_1596,N_1550);
nor U1659 (N_1659,N_1593,N_1508);
and U1660 (N_1660,N_1591,N_1551);
nand U1661 (N_1661,N_1536,N_1587);
nor U1662 (N_1662,N_1500,N_1600);
and U1663 (N_1663,N_1531,N_1581);
or U1664 (N_1664,N_1590,N_1602);
nand U1665 (N_1665,N_1604,N_1592);
xnor U1666 (N_1666,N_1544,N_1624);
and U1667 (N_1667,N_1554,N_1520);
xor U1668 (N_1668,N_1547,N_1607);
or U1669 (N_1669,N_1530,N_1621);
and U1670 (N_1670,N_1588,N_1517);
nor U1671 (N_1671,N_1580,N_1528);
nand U1672 (N_1672,N_1585,N_1505);
nor U1673 (N_1673,N_1595,N_1507);
xor U1674 (N_1674,N_1519,N_1619);
nand U1675 (N_1675,N_1552,N_1557);
nor U1676 (N_1676,N_1573,N_1613);
and U1677 (N_1677,N_1564,N_1523);
or U1678 (N_1678,N_1582,N_1561);
nand U1679 (N_1679,N_1617,N_1503);
xnor U1680 (N_1680,N_1597,N_1567);
and U1681 (N_1681,N_1570,N_1572);
nor U1682 (N_1682,N_1565,N_1614);
nand U1683 (N_1683,N_1577,N_1510);
xor U1684 (N_1684,N_1615,N_1599);
nor U1685 (N_1685,N_1601,N_1521);
xor U1686 (N_1686,N_1560,N_1542);
nor U1687 (N_1687,N_1529,N_1530);
and U1688 (N_1688,N_1609,N_1569);
nor U1689 (N_1689,N_1530,N_1533);
and U1690 (N_1690,N_1512,N_1534);
and U1691 (N_1691,N_1597,N_1601);
nor U1692 (N_1692,N_1606,N_1534);
or U1693 (N_1693,N_1558,N_1531);
nand U1694 (N_1694,N_1553,N_1500);
xnor U1695 (N_1695,N_1551,N_1555);
nand U1696 (N_1696,N_1602,N_1585);
or U1697 (N_1697,N_1541,N_1564);
and U1698 (N_1698,N_1541,N_1587);
or U1699 (N_1699,N_1571,N_1520);
and U1700 (N_1700,N_1576,N_1588);
nor U1701 (N_1701,N_1512,N_1518);
nor U1702 (N_1702,N_1554,N_1516);
nor U1703 (N_1703,N_1594,N_1621);
nand U1704 (N_1704,N_1528,N_1536);
xnor U1705 (N_1705,N_1519,N_1578);
nor U1706 (N_1706,N_1568,N_1601);
or U1707 (N_1707,N_1527,N_1563);
or U1708 (N_1708,N_1567,N_1585);
or U1709 (N_1709,N_1552,N_1579);
and U1710 (N_1710,N_1504,N_1606);
nand U1711 (N_1711,N_1534,N_1538);
nand U1712 (N_1712,N_1566,N_1583);
nand U1713 (N_1713,N_1611,N_1509);
and U1714 (N_1714,N_1527,N_1614);
nor U1715 (N_1715,N_1594,N_1540);
and U1716 (N_1716,N_1590,N_1587);
xor U1717 (N_1717,N_1586,N_1577);
or U1718 (N_1718,N_1506,N_1588);
or U1719 (N_1719,N_1612,N_1600);
nand U1720 (N_1720,N_1586,N_1555);
xnor U1721 (N_1721,N_1612,N_1522);
xnor U1722 (N_1722,N_1621,N_1604);
nand U1723 (N_1723,N_1524,N_1533);
and U1724 (N_1724,N_1598,N_1613);
nand U1725 (N_1725,N_1501,N_1552);
nor U1726 (N_1726,N_1582,N_1517);
or U1727 (N_1727,N_1568,N_1510);
xor U1728 (N_1728,N_1545,N_1524);
xor U1729 (N_1729,N_1583,N_1510);
nor U1730 (N_1730,N_1513,N_1517);
nand U1731 (N_1731,N_1510,N_1596);
nor U1732 (N_1732,N_1503,N_1608);
and U1733 (N_1733,N_1524,N_1505);
or U1734 (N_1734,N_1521,N_1537);
or U1735 (N_1735,N_1524,N_1622);
xnor U1736 (N_1736,N_1518,N_1581);
xnor U1737 (N_1737,N_1581,N_1542);
nor U1738 (N_1738,N_1624,N_1512);
xnor U1739 (N_1739,N_1556,N_1520);
or U1740 (N_1740,N_1610,N_1604);
nand U1741 (N_1741,N_1524,N_1580);
and U1742 (N_1742,N_1528,N_1604);
xor U1743 (N_1743,N_1541,N_1508);
and U1744 (N_1744,N_1537,N_1575);
nor U1745 (N_1745,N_1524,N_1612);
and U1746 (N_1746,N_1584,N_1563);
or U1747 (N_1747,N_1578,N_1620);
and U1748 (N_1748,N_1599,N_1606);
nor U1749 (N_1749,N_1550,N_1541);
or U1750 (N_1750,N_1625,N_1727);
and U1751 (N_1751,N_1649,N_1643);
nor U1752 (N_1752,N_1629,N_1737);
nor U1753 (N_1753,N_1646,N_1680);
xnor U1754 (N_1754,N_1627,N_1660);
nand U1755 (N_1755,N_1715,N_1731);
or U1756 (N_1756,N_1691,N_1749);
and U1757 (N_1757,N_1708,N_1694);
nor U1758 (N_1758,N_1639,N_1710);
or U1759 (N_1759,N_1650,N_1725);
and U1760 (N_1760,N_1656,N_1735);
nand U1761 (N_1761,N_1695,N_1661);
or U1762 (N_1762,N_1642,N_1729);
nand U1763 (N_1763,N_1640,N_1700);
nor U1764 (N_1764,N_1652,N_1736);
or U1765 (N_1765,N_1733,N_1673);
or U1766 (N_1766,N_1684,N_1686);
nor U1767 (N_1767,N_1742,N_1716);
xor U1768 (N_1768,N_1666,N_1672);
nor U1769 (N_1769,N_1712,N_1698);
and U1770 (N_1770,N_1676,N_1654);
nor U1771 (N_1771,N_1638,N_1683);
xor U1772 (N_1772,N_1718,N_1740);
nor U1773 (N_1773,N_1667,N_1688);
nor U1774 (N_1774,N_1677,N_1635);
or U1775 (N_1775,N_1664,N_1647);
or U1776 (N_1776,N_1662,N_1719);
nor U1777 (N_1777,N_1732,N_1633);
xnor U1778 (N_1778,N_1746,N_1747);
or U1779 (N_1779,N_1702,N_1692);
nand U1780 (N_1780,N_1657,N_1713);
nor U1781 (N_1781,N_1645,N_1711);
xor U1782 (N_1782,N_1701,N_1641);
xor U1783 (N_1783,N_1714,N_1628);
xnor U1784 (N_1784,N_1696,N_1659);
xor U1785 (N_1785,N_1723,N_1699);
nand U1786 (N_1786,N_1674,N_1730);
and U1787 (N_1787,N_1720,N_1685);
or U1788 (N_1788,N_1644,N_1734);
nand U1789 (N_1789,N_1626,N_1728);
nand U1790 (N_1790,N_1726,N_1675);
nand U1791 (N_1791,N_1738,N_1653);
xnor U1792 (N_1792,N_1631,N_1678);
nor U1793 (N_1793,N_1705,N_1704);
xor U1794 (N_1794,N_1709,N_1744);
nor U1795 (N_1795,N_1697,N_1668);
xnor U1796 (N_1796,N_1670,N_1651);
nand U1797 (N_1797,N_1706,N_1630);
xnor U1798 (N_1798,N_1748,N_1743);
nor U1799 (N_1799,N_1717,N_1679);
and U1800 (N_1800,N_1739,N_1669);
nand U1801 (N_1801,N_1632,N_1636);
xor U1802 (N_1802,N_1648,N_1665);
or U1803 (N_1803,N_1687,N_1724);
nor U1804 (N_1804,N_1655,N_1693);
nor U1805 (N_1805,N_1671,N_1681);
and U1806 (N_1806,N_1663,N_1690);
xor U1807 (N_1807,N_1722,N_1721);
xnor U1808 (N_1808,N_1682,N_1634);
nand U1809 (N_1809,N_1703,N_1745);
or U1810 (N_1810,N_1689,N_1707);
nor U1811 (N_1811,N_1741,N_1637);
or U1812 (N_1812,N_1658,N_1625);
or U1813 (N_1813,N_1749,N_1649);
nor U1814 (N_1814,N_1669,N_1661);
nor U1815 (N_1815,N_1653,N_1700);
and U1816 (N_1816,N_1713,N_1629);
nand U1817 (N_1817,N_1630,N_1671);
nor U1818 (N_1818,N_1642,N_1687);
or U1819 (N_1819,N_1715,N_1655);
nor U1820 (N_1820,N_1640,N_1736);
nand U1821 (N_1821,N_1679,N_1731);
and U1822 (N_1822,N_1658,N_1629);
or U1823 (N_1823,N_1662,N_1729);
nor U1824 (N_1824,N_1739,N_1713);
or U1825 (N_1825,N_1692,N_1730);
xor U1826 (N_1826,N_1633,N_1678);
or U1827 (N_1827,N_1638,N_1705);
and U1828 (N_1828,N_1709,N_1726);
nand U1829 (N_1829,N_1657,N_1668);
and U1830 (N_1830,N_1715,N_1683);
nor U1831 (N_1831,N_1668,N_1727);
nor U1832 (N_1832,N_1700,N_1692);
nand U1833 (N_1833,N_1636,N_1678);
nand U1834 (N_1834,N_1708,N_1717);
nor U1835 (N_1835,N_1650,N_1718);
or U1836 (N_1836,N_1721,N_1747);
or U1837 (N_1837,N_1707,N_1724);
nor U1838 (N_1838,N_1749,N_1724);
xnor U1839 (N_1839,N_1626,N_1642);
nand U1840 (N_1840,N_1685,N_1698);
xor U1841 (N_1841,N_1646,N_1718);
and U1842 (N_1842,N_1701,N_1730);
and U1843 (N_1843,N_1717,N_1680);
or U1844 (N_1844,N_1675,N_1719);
or U1845 (N_1845,N_1655,N_1658);
xnor U1846 (N_1846,N_1674,N_1707);
nand U1847 (N_1847,N_1627,N_1708);
or U1848 (N_1848,N_1725,N_1712);
and U1849 (N_1849,N_1630,N_1639);
xor U1850 (N_1850,N_1734,N_1699);
or U1851 (N_1851,N_1635,N_1712);
and U1852 (N_1852,N_1628,N_1724);
xor U1853 (N_1853,N_1674,N_1684);
nor U1854 (N_1854,N_1742,N_1656);
xnor U1855 (N_1855,N_1697,N_1679);
nor U1856 (N_1856,N_1705,N_1670);
and U1857 (N_1857,N_1691,N_1684);
nand U1858 (N_1858,N_1714,N_1727);
and U1859 (N_1859,N_1725,N_1641);
nor U1860 (N_1860,N_1636,N_1656);
and U1861 (N_1861,N_1701,N_1705);
nand U1862 (N_1862,N_1705,N_1685);
nand U1863 (N_1863,N_1659,N_1733);
nor U1864 (N_1864,N_1749,N_1712);
xnor U1865 (N_1865,N_1631,N_1659);
or U1866 (N_1866,N_1657,N_1638);
xnor U1867 (N_1867,N_1718,N_1721);
or U1868 (N_1868,N_1661,N_1682);
nand U1869 (N_1869,N_1662,N_1647);
or U1870 (N_1870,N_1633,N_1630);
or U1871 (N_1871,N_1672,N_1708);
nand U1872 (N_1872,N_1648,N_1646);
nand U1873 (N_1873,N_1749,N_1733);
nor U1874 (N_1874,N_1713,N_1715);
nor U1875 (N_1875,N_1801,N_1811);
nand U1876 (N_1876,N_1864,N_1794);
xor U1877 (N_1877,N_1853,N_1762);
or U1878 (N_1878,N_1838,N_1804);
xor U1879 (N_1879,N_1815,N_1823);
nor U1880 (N_1880,N_1757,N_1750);
nand U1881 (N_1881,N_1786,N_1816);
or U1882 (N_1882,N_1751,N_1819);
nor U1883 (N_1883,N_1840,N_1774);
nor U1884 (N_1884,N_1769,N_1812);
and U1885 (N_1885,N_1813,N_1835);
nor U1886 (N_1886,N_1800,N_1780);
or U1887 (N_1887,N_1841,N_1767);
and U1888 (N_1888,N_1770,N_1870);
nand U1889 (N_1889,N_1868,N_1779);
nor U1890 (N_1890,N_1825,N_1756);
nor U1891 (N_1891,N_1759,N_1781);
nor U1892 (N_1892,N_1810,N_1836);
or U1893 (N_1893,N_1854,N_1760);
nand U1894 (N_1894,N_1833,N_1778);
nor U1895 (N_1895,N_1847,N_1837);
xor U1896 (N_1896,N_1845,N_1849);
nand U1897 (N_1897,N_1758,N_1826);
nand U1898 (N_1898,N_1796,N_1807);
xnor U1899 (N_1899,N_1871,N_1867);
and U1900 (N_1900,N_1761,N_1782);
or U1901 (N_1901,N_1828,N_1798);
nand U1902 (N_1902,N_1834,N_1844);
nor U1903 (N_1903,N_1785,N_1772);
and U1904 (N_1904,N_1866,N_1817);
nor U1905 (N_1905,N_1842,N_1831);
and U1906 (N_1906,N_1763,N_1806);
or U1907 (N_1907,N_1843,N_1795);
or U1908 (N_1908,N_1765,N_1852);
nand U1909 (N_1909,N_1754,N_1846);
xnor U1910 (N_1910,N_1802,N_1752);
nand U1911 (N_1911,N_1792,N_1872);
nand U1912 (N_1912,N_1859,N_1776);
xor U1913 (N_1913,N_1829,N_1803);
or U1914 (N_1914,N_1809,N_1793);
xor U1915 (N_1915,N_1827,N_1865);
and U1916 (N_1916,N_1773,N_1851);
nor U1917 (N_1917,N_1771,N_1874);
nand U1918 (N_1918,N_1862,N_1830);
nand U1919 (N_1919,N_1850,N_1775);
nand U1920 (N_1920,N_1755,N_1784);
and U1921 (N_1921,N_1789,N_1839);
nor U1922 (N_1922,N_1860,N_1873);
nor U1923 (N_1923,N_1855,N_1799);
nor U1924 (N_1924,N_1805,N_1777);
xor U1925 (N_1925,N_1821,N_1820);
or U1926 (N_1926,N_1766,N_1824);
nand U1927 (N_1927,N_1863,N_1818);
xnor U1928 (N_1928,N_1790,N_1869);
xnor U1929 (N_1929,N_1787,N_1791);
and U1930 (N_1930,N_1783,N_1768);
xnor U1931 (N_1931,N_1861,N_1822);
or U1932 (N_1932,N_1764,N_1858);
nand U1933 (N_1933,N_1856,N_1797);
xor U1934 (N_1934,N_1832,N_1808);
or U1935 (N_1935,N_1857,N_1788);
nand U1936 (N_1936,N_1814,N_1848);
nor U1937 (N_1937,N_1753,N_1821);
and U1938 (N_1938,N_1757,N_1809);
xnor U1939 (N_1939,N_1798,N_1854);
or U1940 (N_1940,N_1846,N_1778);
nand U1941 (N_1941,N_1750,N_1850);
xnor U1942 (N_1942,N_1755,N_1840);
nand U1943 (N_1943,N_1764,N_1806);
or U1944 (N_1944,N_1829,N_1770);
nor U1945 (N_1945,N_1831,N_1871);
nor U1946 (N_1946,N_1842,N_1777);
nor U1947 (N_1947,N_1859,N_1863);
nand U1948 (N_1948,N_1785,N_1789);
and U1949 (N_1949,N_1850,N_1791);
nand U1950 (N_1950,N_1770,N_1761);
and U1951 (N_1951,N_1782,N_1825);
nand U1952 (N_1952,N_1807,N_1856);
xnor U1953 (N_1953,N_1827,N_1837);
nand U1954 (N_1954,N_1846,N_1845);
nor U1955 (N_1955,N_1874,N_1867);
nor U1956 (N_1956,N_1842,N_1868);
nand U1957 (N_1957,N_1763,N_1848);
and U1958 (N_1958,N_1804,N_1813);
xnor U1959 (N_1959,N_1790,N_1788);
nor U1960 (N_1960,N_1813,N_1855);
nor U1961 (N_1961,N_1792,N_1801);
xnor U1962 (N_1962,N_1760,N_1856);
xor U1963 (N_1963,N_1790,N_1872);
nand U1964 (N_1964,N_1778,N_1752);
or U1965 (N_1965,N_1826,N_1808);
nor U1966 (N_1966,N_1865,N_1839);
nand U1967 (N_1967,N_1830,N_1750);
xnor U1968 (N_1968,N_1816,N_1873);
and U1969 (N_1969,N_1816,N_1867);
and U1970 (N_1970,N_1858,N_1779);
xnor U1971 (N_1971,N_1780,N_1804);
or U1972 (N_1972,N_1815,N_1774);
nor U1973 (N_1973,N_1854,N_1861);
xnor U1974 (N_1974,N_1751,N_1792);
or U1975 (N_1975,N_1821,N_1816);
nand U1976 (N_1976,N_1795,N_1788);
xnor U1977 (N_1977,N_1848,N_1856);
nor U1978 (N_1978,N_1837,N_1803);
or U1979 (N_1979,N_1834,N_1874);
or U1980 (N_1980,N_1820,N_1830);
and U1981 (N_1981,N_1758,N_1764);
or U1982 (N_1982,N_1873,N_1865);
nor U1983 (N_1983,N_1764,N_1842);
nand U1984 (N_1984,N_1808,N_1831);
nor U1985 (N_1985,N_1835,N_1791);
nand U1986 (N_1986,N_1795,N_1846);
or U1987 (N_1987,N_1805,N_1834);
and U1988 (N_1988,N_1757,N_1836);
xor U1989 (N_1989,N_1788,N_1854);
nor U1990 (N_1990,N_1831,N_1844);
xor U1991 (N_1991,N_1796,N_1782);
xor U1992 (N_1992,N_1753,N_1874);
and U1993 (N_1993,N_1817,N_1752);
nand U1994 (N_1994,N_1845,N_1835);
or U1995 (N_1995,N_1869,N_1793);
xnor U1996 (N_1996,N_1784,N_1872);
xnor U1997 (N_1997,N_1867,N_1836);
nand U1998 (N_1998,N_1766,N_1841);
xnor U1999 (N_1999,N_1826,N_1857);
xnor U2000 (N_2000,N_1999,N_1912);
nand U2001 (N_2001,N_1916,N_1929);
xor U2002 (N_2002,N_1906,N_1924);
xor U2003 (N_2003,N_1974,N_1927);
or U2004 (N_2004,N_1996,N_1940);
xnor U2005 (N_2005,N_1959,N_1898);
or U2006 (N_2006,N_1909,N_1914);
nor U2007 (N_2007,N_1879,N_1971);
xnor U2008 (N_2008,N_1951,N_1993);
and U2009 (N_2009,N_1917,N_1964);
nand U2010 (N_2010,N_1876,N_1968);
nor U2011 (N_2011,N_1979,N_1960);
xor U2012 (N_2012,N_1995,N_1885);
xor U2013 (N_2013,N_1893,N_1926);
or U2014 (N_2014,N_1928,N_1990);
and U2015 (N_2015,N_1899,N_1976);
nor U2016 (N_2016,N_1961,N_1887);
and U2017 (N_2017,N_1967,N_1910);
or U2018 (N_2018,N_1883,N_1985);
nand U2019 (N_2019,N_1884,N_1925);
nand U2020 (N_2020,N_1994,N_1945);
xnor U2021 (N_2021,N_1892,N_1918);
xor U2022 (N_2022,N_1958,N_1950);
and U2023 (N_2023,N_1880,N_1989);
and U2024 (N_2024,N_1983,N_1966);
or U2025 (N_2025,N_1939,N_1923);
and U2026 (N_2026,N_1878,N_1987);
nand U2027 (N_2027,N_1963,N_1882);
and U2028 (N_2028,N_1890,N_1970);
and U2029 (N_2029,N_1919,N_1997);
nor U2030 (N_2030,N_1953,N_1956);
xnor U2031 (N_2031,N_1930,N_1935);
or U2032 (N_2032,N_1915,N_1904);
xor U2033 (N_2033,N_1900,N_1891);
or U2034 (N_2034,N_1881,N_1911);
nand U2035 (N_2035,N_1902,N_1957);
or U2036 (N_2036,N_1920,N_1877);
nor U2037 (N_2037,N_1955,N_1942);
nor U2038 (N_2038,N_1936,N_1980);
xor U2039 (N_2039,N_1888,N_1886);
or U2040 (N_2040,N_1889,N_1897);
or U2041 (N_2041,N_1938,N_1949);
or U2042 (N_2042,N_1895,N_1975);
xnor U2043 (N_2043,N_1943,N_1903);
nand U2044 (N_2044,N_1875,N_1972);
nor U2045 (N_2045,N_1947,N_1896);
or U2046 (N_2046,N_1933,N_1937);
and U2047 (N_2047,N_1977,N_1991);
nand U2048 (N_2048,N_1934,N_1986);
xor U2049 (N_2049,N_1922,N_1907);
and U2050 (N_2050,N_1931,N_1982);
nand U2051 (N_2051,N_1894,N_1984);
and U2052 (N_2052,N_1978,N_1981);
or U2053 (N_2053,N_1969,N_1948);
and U2054 (N_2054,N_1901,N_1905);
nand U2055 (N_2055,N_1921,N_1954);
xor U2056 (N_2056,N_1962,N_1952);
xor U2057 (N_2057,N_1932,N_1973);
and U2058 (N_2058,N_1988,N_1908);
nor U2059 (N_2059,N_1946,N_1998);
nor U2060 (N_2060,N_1965,N_1992);
and U2061 (N_2061,N_1941,N_1944);
or U2062 (N_2062,N_1913,N_1931);
nor U2063 (N_2063,N_1889,N_1974);
nor U2064 (N_2064,N_1926,N_1999);
and U2065 (N_2065,N_1984,N_1939);
or U2066 (N_2066,N_1951,N_1961);
or U2067 (N_2067,N_1896,N_1968);
nand U2068 (N_2068,N_1948,N_1936);
and U2069 (N_2069,N_1950,N_1946);
and U2070 (N_2070,N_1969,N_1986);
nor U2071 (N_2071,N_1987,N_1950);
and U2072 (N_2072,N_1989,N_1893);
xor U2073 (N_2073,N_1911,N_1905);
nor U2074 (N_2074,N_1950,N_1964);
nor U2075 (N_2075,N_1903,N_1959);
xor U2076 (N_2076,N_1917,N_1916);
xor U2077 (N_2077,N_1921,N_1999);
xor U2078 (N_2078,N_1974,N_1991);
nor U2079 (N_2079,N_1915,N_1926);
nand U2080 (N_2080,N_1983,N_1929);
nor U2081 (N_2081,N_1877,N_1997);
or U2082 (N_2082,N_1913,N_1939);
and U2083 (N_2083,N_1995,N_1880);
or U2084 (N_2084,N_1914,N_1968);
nor U2085 (N_2085,N_1963,N_1931);
and U2086 (N_2086,N_1997,N_1979);
nand U2087 (N_2087,N_1932,N_1951);
nor U2088 (N_2088,N_1922,N_1971);
or U2089 (N_2089,N_1972,N_1905);
nor U2090 (N_2090,N_1952,N_1966);
nor U2091 (N_2091,N_1913,N_1969);
xnor U2092 (N_2092,N_1926,N_1981);
or U2093 (N_2093,N_1917,N_1950);
and U2094 (N_2094,N_1972,N_1944);
xnor U2095 (N_2095,N_1904,N_1958);
xnor U2096 (N_2096,N_1912,N_1950);
nand U2097 (N_2097,N_1923,N_1908);
nor U2098 (N_2098,N_1900,N_1911);
nor U2099 (N_2099,N_1930,N_1990);
and U2100 (N_2100,N_1918,N_1894);
and U2101 (N_2101,N_1921,N_1937);
nor U2102 (N_2102,N_1941,N_1905);
nor U2103 (N_2103,N_1955,N_1976);
nand U2104 (N_2104,N_1915,N_1963);
nor U2105 (N_2105,N_1996,N_1878);
nor U2106 (N_2106,N_1892,N_1995);
and U2107 (N_2107,N_1895,N_1921);
or U2108 (N_2108,N_1939,N_1956);
and U2109 (N_2109,N_1989,N_1921);
or U2110 (N_2110,N_1905,N_1876);
nand U2111 (N_2111,N_1929,N_1888);
or U2112 (N_2112,N_1908,N_1899);
nor U2113 (N_2113,N_1914,N_1883);
xnor U2114 (N_2114,N_1926,N_1918);
xnor U2115 (N_2115,N_1887,N_1893);
nand U2116 (N_2116,N_1895,N_1965);
and U2117 (N_2117,N_1910,N_1941);
or U2118 (N_2118,N_1918,N_1997);
nand U2119 (N_2119,N_1927,N_1981);
or U2120 (N_2120,N_1949,N_1902);
xnor U2121 (N_2121,N_1908,N_1960);
and U2122 (N_2122,N_1972,N_1984);
or U2123 (N_2123,N_1950,N_1886);
nand U2124 (N_2124,N_1992,N_1882);
xnor U2125 (N_2125,N_2076,N_2118);
nor U2126 (N_2126,N_2005,N_2047);
nand U2127 (N_2127,N_2002,N_2006);
nand U2128 (N_2128,N_2083,N_2065);
nand U2129 (N_2129,N_2011,N_2110);
and U2130 (N_2130,N_2067,N_2014);
nand U2131 (N_2131,N_2060,N_2030);
nor U2132 (N_2132,N_2013,N_2081);
nand U2133 (N_2133,N_2048,N_2029);
and U2134 (N_2134,N_2106,N_2102);
nand U2135 (N_2135,N_2026,N_2079);
or U2136 (N_2136,N_2043,N_2050);
xnor U2137 (N_2137,N_2115,N_2095);
and U2138 (N_2138,N_2044,N_2027);
or U2139 (N_2139,N_2109,N_2046);
nor U2140 (N_2140,N_2022,N_2008);
xnor U2141 (N_2141,N_2096,N_2069);
and U2142 (N_2142,N_2054,N_2035);
or U2143 (N_2143,N_2052,N_2103);
nor U2144 (N_2144,N_2017,N_2012);
and U2145 (N_2145,N_2073,N_2078);
nor U2146 (N_2146,N_2116,N_2028);
xnor U2147 (N_2147,N_2124,N_2113);
or U2148 (N_2148,N_2021,N_2009);
and U2149 (N_2149,N_2056,N_2020);
and U2150 (N_2150,N_2120,N_2034);
or U2151 (N_2151,N_2107,N_2084);
and U2152 (N_2152,N_2100,N_2068);
nor U2153 (N_2153,N_2112,N_2074);
and U2154 (N_2154,N_2049,N_2121);
and U2155 (N_2155,N_2114,N_2055);
or U2156 (N_2156,N_2061,N_2038);
nand U2157 (N_2157,N_2098,N_2123);
and U2158 (N_2158,N_2031,N_2033);
xnor U2159 (N_2159,N_2037,N_2091);
xnor U2160 (N_2160,N_2023,N_2045);
xnor U2161 (N_2161,N_2062,N_2080);
nand U2162 (N_2162,N_2122,N_2041);
or U2163 (N_2163,N_2066,N_2000);
xor U2164 (N_2164,N_2001,N_2004);
nand U2165 (N_2165,N_2039,N_2119);
xor U2166 (N_2166,N_2003,N_2092);
or U2167 (N_2167,N_2019,N_2111);
or U2168 (N_2168,N_2086,N_2070);
xor U2169 (N_2169,N_2082,N_2087);
nand U2170 (N_2170,N_2072,N_2090);
xor U2171 (N_2171,N_2099,N_2007);
xnor U2172 (N_2172,N_2117,N_2089);
nor U2173 (N_2173,N_2032,N_2053);
nand U2174 (N_2174,N_2077,N_2024);
or U2175 (N_2175,N_2097,N_2104);
xnor U2176 (N_2176,N_2064,N_2057);
and U2177 (N_2177,N_2088,N_2085);
and U2178 (N_2178,N_2025,N_2071);
nand U2179 (N_2179,N_2094,N_2093);
nor U2180 (N_2180,N_2063,N_2016);
or U2181 (N_2181,N_2040,N_2018);
nand U2182 (N_2182,N_2010,N_2059);
and U2183 (N_2183,N_2101,N_2015);
or U2184 (N_2184,N_2075,N_2036);
and U2185 (N_2185,N_2058,N_2042);
and U2186 (N_2186,N_2051,N_2105);
and U2187 (N_2187,N_2108,N_2031);
or U2188 (N_2188,N_2056,N_2081);
nor U2189 (N_2189,N_2037,N_2006);
xnor U2190 (N_2190,N_2073,N_2093);
and U2191 (N_2191,N_2018,N_2028);
nor U2192 (N_2192,N_2103,N_2000);
or U2193 (N_2193,N_2007,N_2115);
nand U2194 (N_2194,N_2094,N_2046);
nand U2195 (N_2195,N_2088,N_2004);
and U2196 (N_2196,N_2043,N_2119);
nand U2197 (N_2197,N_2092,N_2039);
or U2198 (N_2198,N_2077,N_2034);
xor U2199 (N_2199,N_2011,N_2116);
or U2200 (N_2200,N_2119,N_2094);
and U2201 (N_2201,N_2068,N_2014);
nor U2202 (N_2202,N_2047,N_2115);
nor U2203 (N_2203,N_2080,N_2044);
or U2204 (N_2204,N_2097,N_2055);
nand U2205 (N_2205,N_2048,N_2060);
or U2206 (N_2206,N_2042,N_2053);
and U2207 (N_2207,N_2009,N_2002);
xor U2208 (N_2208,N_2099,N_2052);
and U2209 (N_2209,N_2007,N_2005);
nand U2210 (N_2210,N_2034,N_2056);
nand U2211 (N_2211,N_2097,N_2101);
or U2212 (N_2212,N_2018,N_2036);
nand U2213 (N_2213,N_2003,N_2095);
and U2214 (N_2214,N_2034,N_2019);
nand U2215 (N_2215,N_2067,N_2040);
xor U2216 (N_2216,N_2084,N_2014);
or U2217 (N_2217,N_2074,N_2064);
nand U2218 (N_2218,N_2072,N_2087);
nor U2219 (N_2219,N_2041,N_2087);
xor U2220 (N_2220,N_2100,N_2034);
xor U2221 (N_2221,N_2062,N_2107);
and U2222 (N_2222,N_2067,N_2003);
nand U2223 (N_2223,N_2047,N_2048);
nor U2224 (N_2224,N_2028,N_2069);
nand U2225 (N_2225,N_2011,N_2090);
or U2226 (N_2226,N_2101,N_2041);
xor U2227 (N_2227,N_2015,N_2039);
nand U2228 (N_2228,N_2071,N_2004);
nand U2229 (N_2229,N_2019,N_2080);
or U2230 (N_2230,N_2084,N_2091);
xnor U2231 (N_2231,N_2064,N_2037);
xnor U2232 (N_2232,N_2025,N_2016);
or U2233 (N_2233,N_2056,N_2109);
nand U2234 (N_2234,N_2079,N_2007);
xor U2235 (N_2235,N_2080,N_2040);
or U2236 (N_2236,N_2019,N_2016);
and U2237 (N_2237,N_2031,N_2111);
or U2238 (N_2238,N_2030,N_2104);
or U2239 (N_2239,N_2109,N_2001);
or U2240 (N_2240,N_2050,N_2062);
and U2241 (N_2241,N_2122,N_2092);
nor U2242 (N_2242,N_2051,N_2032);
nor U2243 (N_2243,N_2050,N_2067);
nand U2244 (N_2244,N_2101,N_2001);
and U2245 (N_2245,N_2068,N_2006);
nand U2246 (N_2246,N_2053,N_2033);
nand U2247 (N_2247,N_2090,N_2001);
and U2248 (N_2248,N_2034,N_2066);
nand U2249 (N_2249,N_2038,N_2055);
nor U2250 (N_2250,N_2205,N_2217);
nor U2251 (N_2251,N_2231,N_2180);
nand U2252 (N_2252,N_2243,N_2151);
and U2253 (N_2253,N_2200,N_2213);
and U2254 (N_2254,N_2245,N_2157);
nand U2255 (N_2255,N_2128,N_2125);
or U2256 (N_2256,N_2147,N_2235);
or U2257 (N_2257,N_2139,N_2177);
nor U2258 (N_2258,N_2249,N_2211);
xor U2259 (N_2259,N_2229,N_2215);
nand U2260 (N_2260,N_2218,N_2175);
nor U2261 (N_2261,N_2248,N_2222);
and U2262 (N_2262,N_2210,N_2165);
nor U2263 (N_2263,N_2127,N_2206);
nor U2264 (N_2264,N_2159,N_2209);
nand U2265 (N_2265,N_2226,N_2244);
nor U2266 (N_2266,N_2191,N_2169);
nor U2267 (N_2267,N_2144,N_2152);
and U2268 (N_2268,N_2131,N_2190);
nor U2269 (N_2269,N_2193,N_2212);
nand U2270 (N_2270,N_2216,N_2197);
xor U2271 (N_2271,N_2220,N_2207);
xnor U2272 (N_2272,N_2136,N_2202);
nand U2273 (N_2273,N_2163,N_2146);
xnor U2274 (N_2274,N_2201,N_2134);
xnor U2275 (N_2275,N_2203,N_2236);
nor U2276 (N_2276,N_2178,N_2137);
or U2277 (N_2277,N_2237,N_2182);
and U2278 (N_2278,N_2142,N_2247);
nand U2279 (N_2279,N_2219,N_2214);
nand U2280 (N_2280,N_2238,N_2183);
xnor U2281 (N_2281,N_2126,N_2170);
and U2282 (N_2282,N_2154,N_2241);
or U2283 (N_2283,N_2171,N_2228);
nor U2284 (N_2284,N_2138,N_2192);
nor U2285 (N_2285,N_2162,N_2240);
and U2286 (N_2286,N_2155,N_2179);
nor U2287 (N_2287,N_2189,N_2242);
and U2288 (N_2288,N_2196,N_2184);
or U2289 (N_2289,N_2188,N_2135);
nand U2290 (N_2290,N_2230,N_2232);
nor U2291 (N_2291,N_2141,N_2181);
nand U2292 (N_2292,N_2156,N_2132);
or U2293 (N_2293,N_2161,N_2221);
nor U2294 (N_2294,N_2172,N_2129);
or U2295 (N_2295,N_2140,N_2174);
nor U2296 (N_2296,N_2186,N_2160);
nand U2297 (N_2297,N_2167,N_2158);
nand U2298 (N_2298,N_2224,N_2176);
nor U2299 (N_2299,N_2168,N_2164);
or U2300 (N_2300,N_2233,N_2149);
xnor U2301 (N_2301,N_2227,N_2145);
or U2302 (N_2302,N_2173,N_2223);
and U2303 (N_2303,N_2194,N_2246);
and U2304 (N_2304,N_2239,N_2166);
and U2305 (N_2305,N_2143,N_2199);
nand U2306 (N_2306,N_2133,N_2195);
or U2307 (N_2307,N_2148,N_2150);
xor U2308 (N_2308,N_2225,N_2153);
nand U2309 (N_2309,N_2187,N_2208);
and U2310 (N_2310,N_2130,N_2204);
nor U2311 (N_2311,N_2198,N_2185);
nor U2312 (N_2312,N_2234,N_2200);
and U2313 (N_2313,N_2232,N_2175);
or U2314 (N_2314,N_2162,N_2203);
nor U2315 (N_2315,N_2176,N_2210);
nor U2316 (N_2316,N_2146,N_2224);
or U2317 (N_2317,N_2193,N_2181);
xor U2318 (N_2318,N_2231,N_2240);
xor U2319 (N_2319,N_2148,N_2152);
nand U2320 (N_2320,N_2155,N_2184);
nor U2321 (N_2321,N_2127,N_2159);
or U2322 (N_2322,N_2194,N_2229);
xor U2323 (N_2323,N_2173,N_2159);
and U2324 (N_2324,N_2137,N_2130);
nand U2325 (N_2325,N_2143,N_2139);
nand U2326 (N_2326,N_2213,N_2144);
xor U2327 (N_2327,N_2230,N_2245);
nor U2328 (N_2328,N_2239,N_2237);
and U2329 (N_2329,N_2196,N_2126);
xnor U2330 (N_2330,N_2185,N_2173);
and U2331 (N_2331,N_2203,N_2224);
and U2332 (N_2332,N_2172,N_2128);
xnor U2333 (N_2333,N_2186,N_2221);
or U2334 (N_2334,N_2210,N_2248);
nor U2335 (N_2335,N_2249,N_2136);
or U2336 (N_2336,N_2240,N_2227);
or U2337 (N_2337,N_2145,N_2243);
or U2338 (N_2338,N_2133,N_2216);
nor U2339 (N_2339,N_2156,N_2229);
nand U2340 (N_2340,N_2222,N_2187);
or U2341 (N_2341,N_2205,N_2189);
nand U2342 (N_2342,N_2176,N_2168);
xor U2343 (N_2343,N_2228,N_2248);
or U2344 (N_2344,N_2193,N_2154);
xnor U2345 (N_2345,N_2241,N_2190);
xnor U2346 (N_2346,N_2128,N_2132);
xor U2347 (N_2347,N_2143,N_2147);
and U2348 (N_2348,N_2129,N_2243);
nor U2349 (N_2349,N_2145,N_2213);
nor U2350 (N_2350,N_2160,N_2211);
nor U2351 (N_2351,N_2222,N_2204);
and U2352 (N_2352,N_2142,N_2174);
nand U2353 (N_2353,N_2146,N_2180);
or U2354 (N_2354,N_2241,N_2187);
nand U2355 (N_2355,N_2223,N_2236);
xnor U2356 (N_2356,N_2150,N_2157);
xnor U2357 (N_2357,N_2125,N_2160);
or U2358 (N_2358,N_2186,N_2140);
nand U2359 (N_2359,N_2170,N_2188);
or U2360 (N_2360,N_2223,N_2148);
and U2361 (N_2361,N_2155,N_2206);
and U2362 (N_2362,N_2211,N_2151);
or U2363 (N_2363,N_2176,N_2243);
and U2364 (N_2364,N_2199,N_2132);
and U2365 (N_2365,N_2221,N_2182);
nand U2366 (N_2366,N_2155,N_2180);
xor U2367 (N_2367,N_2181,N_2234);
nor U2368 (N_2368,N_2193,N_2146);
or U2369 (N_2369,N_2187,N_2173);
nand U2370 (N_2370,N_2246,N_2169);
nor U2371 (N_2371,N_2239,N_2156);
nor U2372 (N_2372,N_2159,N_2206);
xnor U2373 (N_2373,N_2165,N_2245);
or U2374 (N_2374,N_2142,N_2181);
nand U2375 (N_2375,N_2266,N_2353);
and U2376 (N_2376,N_2338,N_2263);
xor U2377 (N_2377,N_2306,N_2260);
or U2378 (N_2378,N_2331,N_2283);
xor U2379 (N_2379,N_2366,N_2288);
nand U2380 (N_2380,N_2372,N_2364);
nor U2381 (N_2381,N_2250,N_2294);
nand U2382 (N_2382,N_2360,N_2320);
or U2383 (N_2383,N_2254,N_2335);
nand U2384 (N_2384,N_2268,N_2359);
xnor U2385 (N_2385,N_2362,N_2354);
nor U2386 (N_2386,N_2351,N_2319);
and U2387 (N_2387,N_2334,N_2316);
and U2388 (N_2388,N_2305,N_2270);
and U2389 (N_2389,N_2285,N_2258);
xor U2390 (N_2390,N_2337,N_2284);
nand U2391 (N_2391,N_2256,N_2328);
or U2392 (N_2392,N_2251,N_2315);
and U2393 (N_2393,N_2259,N_2336);
and U2394 (N_2394,N_2355,N_2255);
and U2395 (N_2395,N_2343,N_2369);
nor U2396 (N_2396,N_2357,N_2253);
or U2397 (N_2397,N_2296,N_2265);
nand U2398 (N_2398,N_2257,N_2282);
nor U2399 (N_2399,N_2365,N_2304);
or U2400 (N_2400,N_2347,N_2278);
and U2401 (N_2401,N_2277,N_2329);
or U2402 (N_2402,N_2301,N_2314);
and U2403 (N_2403,N_2363,N_2302);
and U2404 (N_2404,N_2345,N_2293);
and U2405 (N_2405,N_2318,N_2325);
xnor U2406 (N_2406,N_2321,N_2344);
or U2407 (N_2407,N_2332,N_2341);
xor U2408 (N_2408,N_2307,N_2326);
nand U2409 (N_2409,N_2356,N_2300);
or U2410 (N_2410,N_2348,N_2297);
nand U2411 (N_2411,N_2350,N_2371);
and U2412 (N_2412,N_2261,N_2311);
nor U2413 (N_2413,N_2339,N_2290);
and U2414 (N_2414,N_2313,N_2291);
nand U2415 (N_2415,N_2346,N_2308);
nor U2416 (N_2416,N_2323,N_2340);
nand U2417 (N_2417,N_2272,N_2262);
or U2418 (N_2418,N_2269,N_2333);
xnor U2419 (N_2419,N_2295,N_2374);
xnor U2420 (N_2420,N_2281,N_2317);
nor U2421 (N_2421,N_2324,N_2370);
nand U2422 (N_2422,N_2299,N_2330);
nor U2423 (N_2423,N_2273,N_2310);
or U2424 (N_2424,N_2312,N_2264);
nor U2425 (N_2425,N_2303,N_2275);
nor U2426 (N_2426,N_2276,N_2274);
xor U2427 (N_2427,N_2342,N_2287);
nor U2428 (N_2428,N_2367,N_2368);
nor U2429 (N_2429,N_2373,N_2292);
xor U2430 (N_2430,N_2298,N_2271);
and U2431 (N_2431,N_2327,N_2309);
nand U2432 (N_2432,N_2358,N_2286);
xnor U2433 (N_2433,N_2289,N_2252);
xor U2434 (N_2434,N_2279,N_2361);
and U2435 (N_2435,N_2322,N_2280);
xnor U2436 (N_2436,N_2352,N_2349);
nand U2437 (N_2437,N_2267,N_2295);
nor U2438 (N_2438,N_2267,N_2280);
xnor U2439 (N_2439,N_2362,N_2322);
nor U2440 (N_2440,N_2330,N_2341);
or U2441 (N_2441,N_2277,N_2310);
nor U2442 (N_2442,N_2315,N_2338);
nor U2443 (N_2443,N_2275,N_2341);
xnor U2444 (N_2444,N_2278,N_2355);
xnor U2445 (N_2445,N_2292,N_2288);
or U2446 (N_2446,N_2252,N_2284);
nor U2447 (N_2447,N_2295,N_2310);
xor U2448 (N_2448,N_2316,N_2336);
or U2449 (N_2449,N_2356,N_2302);
nor U2450 (N_2450,N_2252,N_2314);
xnor U2451 (N_2451,N_2322,N_2351);
or U2452 (N_2452,N_2287,N_2288);
or U2453 (N_2453,N_2353,N_2350);
nor U2454 (N_2454,N_2300,N_2363);
nor U2455 (N_2455,N_2349,N_2303);
or U2456 (N_2456,N_2348,N_2282);
nand U2457 (N_2457,N_2299,N_2253);
xor U2458 (N_2458,N_2260,N_2287);
xor U2459 (N_2459,N_2365,N_2322);
nor U2460 (N_2460,N_2329,N_2273);
and U2461 (N_2461,N_2252,N_2307);
nor U2462 (N_2462,N_2307,N_2303);
xor U2463 (N_2463,N_2272,N_2306);
xnor U2464 (N_2464,N_2327,N_2323);
nand U2465 (N_2465,N_2319,N_2265);
and U2466 (N_2466,N_2308,N_2259);
xnor U2467 (N_2467,N_2323,N_2369);
xor U2468 (N_2468,N_2312,N_2365);
xor U2469 (N_2469,N_2288,N_2320);
nand U2470 (N_2470,N_2365,N_2284);
or U2471 (N_2471,N_2295,N_2273);
nor U2472 (N_2472,N_2345,N_2343);
and U2473 (N_2473,N_2288,N_2270);
or U2474 (N_2474,N_2260,N_2367);
nand U2475 (N_2475,N_2259,N_2297);
nand U2476 (N_2476,N_2281,N_2294);
and U2477 (N_2477,N_2334,N_2312);
nand U2478 (N_2478,N_2362,N_2346);
or U2479 (N_2479,N_2250,N_2357);
or U2480 (N_2480,N_2347,N_2355);
or U2481 (N_2481,N_2262,N_2351);
and U2482 (N_2482,N_2343,N_2258);
nand U2483 (N_2483,N_2256,N_2372);
and U2484 (N_2484,N_2364,N_2336);
or U2485 (N_2485,N_2270,N_2341);
nor U2486 (N_2486,N_2286,N_2327);
nor U2487 (N_2487,N_2296,N_2369);
nor U2488 (N_2488,N_2344,N_2357);
or U2489 (N_2489,N_2307,N_2263);
xor U2490 (N_2490,N_2251,N_2371);
and U2491 (N_2491,N_2368,N_2357);
or U2492 (N_2492,N_2278,N_2292);
or U2493 (N_2493,N_2293,N_2359);
or U2494 (N_2494,N_2258,N_2280);
nand U2495 (N_2495,N_2308,N_2358);
nand U2496 (N_2496,N_2298,N_2301);
nand U2497 (N_2497,N_2350,N_2296);
nand U2498 (N_2498,N_2361,N_2269);
xor U2499 (N_2499,N_2315,N_2320);
xnor U2500 (N_2500,N_2405,N_2388);
or U2501 (N_2501,N_2493,N_2454);
and U2502 (N_2502,N_2437,N_2458);
and U2503 (N_2503,N_2400,N_2434);
nand U2504 (N_2504,N_2429,N_2385);
and U2505 (N_2505,N_2441,N_2477);
xnor U2506 (N_2506,N_2491,N_2425);
nand U2507 (N_2507,N_2481,N_2455);
nand U2508 (N_2508,N_2460,N_2499);
nand U2509 (N_2509,N_2389,N_2485);
or U2510 (N_2510,N_2421,N_2480);
nor U2511 (N_2511,N_2418,N_2475);
nor U2512 (N_2512,N_2449,N_2376);
and U2513 (N_2513,N_2392,N_2431);
nand U2514 (N_2514,N_2423,N_2432);
and U2515 (N_2515,N_2445,N_2462);
or U2516 (N_2516,N_2446,N_2414);
nor U2517 (N_2517,N_2417,N_2468);
or U2518 (N_2518,N_2474,N_2488);
nand U2519 (N_2519,N_2416,N_2494);
or U2520 (N_2520,N_2433,N_2479);
xnor U2521 (N_2521,N_2470,N_2476);
nand U2522 (N_2522,N_2490,N_2391);
xnor U2523 (N_2523,N_2419,N_2492);
or U2524 (N_2524,N_2386,N_2447);
xnor U2525 (N_2525,N_2375,N_2390);
and U2526 (N_2526,N_2412,N_2487);
and U2527 (N_2527,N_2444,N_2422);
and U2528 (N_2528,N_2408,N_2436);
or U2529 (N_2529,N_2430,N_2463);
nand U2530 (N_2530,N_2413,N_2497);
xor U2531 (N_2531,N_2409,N_2489);
xor U2532 (N_2532,N_2381,N_2404);
nand U2533 (N_2533,N_2452,N_2456);
and U2534 (N_2534,N_2435,N_2402);
or U2535 (N_2535,N_2387,N_2399);
nor U2536 (N_2536,N_2415,N_2420);
xor U2537 (N_2537,N_2380,N_2465);
xnor U2538 (N_2538,N_2466,N_2383);
nor U2539 (N_2539,N_2484,N_2378);
and U2540 (N_2540,N_2496,N_2442);
and U2541 (N_2541,N_2478,N_2467);
or U2542 (N_2542,N_2398,N_2457);
nor U2543 (N_2543,N_2411,N_2450);
nand U2544 (N_2544,N_2410,N_2473);
and U2545 (N_2545,N_2471,N_2451);
xor U2546 (N_2546,N_2483,N_2384);
nand U2547 (N_2547,N_2424,N_2407);
nand U2548 (N_2548,N_2438,N_2377);
nor U2549 (N_2549,N_2498,N_2439);
or U2550 (N_2550,N_2464,N_2428);
or U2551 (N_2551,N_2443,N_2395);
nand U2552 (N_2552,N_2448,N_2382);
and U2553 (N_2553,N_2403,N_2397);
nand U2554 (N_2554,N_2440,N_2472);
nand U2555 (N_2555,N_2459,N_2396);
nand U2556 (N_2556,N_2401,N_2427);
xor U2557 (N_2557,N_2469,N_2495);
or U2558 (N_2558,N_2486,N_2394);
nand U2559 (N_2559,N_2406,N_2482);
nor U2560 (N_2560,N_2461,N_2453);
xnor U2561 (N_2561,N_2379,N_2393);
nor U2562 (N_2562,N_2426,N_2410);
xor U2563 (N_2563,N_2383,N_2440);
nor U2564 (N_2564,N_2488,N_2409);
nand U2565 (N_2565,N_2396,N_2482);
or U2566 (N_2566,N_2433,N_2442);
nor U2567 (N_2567,N_2404,N_2498);
and U2568 (N_2568,N_2468,N_2487);
or U2569 (N_2569,N_2401,N_2416);
xnor U2570 (N_2570,N_2490,N_2376);
nand U2571 (N_2571,N_2379,N_2376);
and U2572 (N_2572,N_2432,N_2444);
nor U2573 (N_2573,N_2498,N_2447);
and U2574 (N_2574,N_2491,N_2430);
nor U2575 (N_2575,N_2409,N_2411);
or U2576 (N_2576,N_2477,N_2475);
or U2577 (N_2577,N_2406,N_2455);
nand U2578 (N_2578,N_2483,N_2468);
xnor U2579 (N_2579,N_2440,N_2467);
and U2580 (N_2580,N_2441,N_2378);
nor U2581 (N_2581,N_2416,N_2409);
nor U2582 (N_2582,N_2417,N_2425);
and U2583 (N_2583,N_2465,N_2409);
xor U2584 (N_2584,N_2485,N_2413);
nand U2585 (N_2585,N_2417,N_2396);
xor U2586 (N_2586,N_2420,N_2467);
and U2587 (N_2587,N_2486,N_2493);
or U2588 (N_2588,N_2495,N_2485);
or U2589 (N_2589,N_2459,N_2457);
and U2590 (N_2590,N_2389,N_2401);
and U2591 (N_2591,N_2396,N_2468);
nor U2592 (N_2592,N_2421,N_2424);
nand U2593 (N_2593,N_2458,N_2447);
or U2594 (N_2594,N_2482,N_2438);
nor U2595 (N_2595,N_2499,N_2428);
and U2596 (N_2596,N_2394,N_2382);
nand U2597 (N_2597,N_2408,N_2412);
or U2598 (N_2598,N_2404,N_2376);
nor U2599 (N_2599,N_2470,N_2471);
xor U2600 (N_2600,N_2422,N_2450);
xnor U2601 (N_2601,N_2397,N_2378);
nor U2602 (N_2602,N_2433,N_2467);
or U2603 (N_2603,N_2490,N_2484);
nor U2604 (N_2604,N_2397,N_2431);
nand U2605 (N_2605,N_2406,N_2459);
and U2606 (N_2606,N_2486,N_2487);
xnor U2607 (N_2607,N_2465,N_2375);
xnor U2608 (N_2608,N_2476,N_2397);
nor U2609 (N_2609,N_2420,N_2379);
nand U2610 (N_2610,N_2436,N_2462);
xnor U2611 (N_2611,N_2402,N_2493);
and U2612 (N_2612,N_2375,N_2447);
or U2613 (N_2613,N_2443,N_2464);
nor U2614 (N_2614,N_2404,N_2418);
nand U2615 (N_2615,N_2489,N_2453);
and U2616 (N_2616,N_2470,N_2481);
nand U2617 (N_2617,N_2422,N_2376);
or U2618 (N_2618,N_2398,N_2469);
nor U2619 (N_2619,N_2439,N_2477);
or U2620 (N_2620,N_2439,N_2496);
and U2621 (N_2621,N_2440,N_2462);
xor U2622 (N_2622,N_2428,N_2463);
xor U2623 (N_2623,N_2473,N_2467);
nand U2624 (N_2624,N_2464,N_2494);
and U2625 (N_2625,N_2616,N_2504);
nand U2626 (N_2626,N_2586,N_2529);
or U2627 (N_2627,N_2533,N_2609);
or U2628 (N_2628,N_2590,N_2549);
or U2629 (N_2629,N_2508,N_2623);
nand U2630 (N_2630,N_2536,N_2524);
or U2631 (N_2631,N_2597,N_2520);
and U2632 (N_2632,N_2617,N_2543);
nand U2633 (N_2633,N_2606,N_2601);
nand U2634 (N_2634,N_2621,N_2512);
nor U2635 (N_2635,N_2534,N_2619);
and U2636 (N_2636,N_2569,N_2605);
nand U2637 (N_2637,N_2525,N_2603);
nor U2638 (N_2638,N_2584,N_2620);
or U2639 (N_2639,N_2596,N_2588);
xor U2640 (N_2640,N_2546,N_2509);
nor U2641 (N_2641,N_2541,N_2622);
nor U2642 (N_2642,N_2612,N_2511);
nand U2643 (N_2643,N_2510,N_2558);
and U2644 (N_2644,N_2537,N_2552);
nand U2645 (N_2645,N_2604,N_2581);
and U2646 (N_2646,N_2513,N_2530);
nand U2647 (N_2647,N_2560,N_2618);
and U2648 (N_2648,N_2565,N_2578);
or U2649 (N_2649,N_2564,N_2580);
or U2650 (N_2650,N_2514,N_2582);
nand U2651 (N_2651,N_2556,N_2506);
or U2652 (N_2652,N_2554,N_2548);
and U2653 (N_2653,N_2515,N_2579);
and U2654 (N_2654,N_2518,N_2539);
nand U2655 (N_2655,N_2531,N_2503);
xor U2656 (N_2656,N_2550,N_2502);
nand U2657 (N_2657,N_2575,N_2519);
nand U2658 (N_2658,N_2551,N_2613);
or U2659 (N_2659,N_2540,N_2545);
xor U2660 (N_2660,N_2572,N_2532);
and U2661 (N_2661,N_2583,N_2611);
xnor U2662 (N_2662,N_2555,N_2610);
nand U2663 (N_2663,N_2595,N_2528);
xnor U2664 (N_2664,N_2563,N_2598);
nand U2665 (N_2665,N_2585,N_2559);
nand U2666 (N_2666,N_2547,N_2592);
or U2667 (N_2667,N_2501,N_2523);
or U2668 (N_2668,N_2602,N_2587);
nor U2669 (N_2669,N_2561,N_2567);
or U2670 (N_2670,N_2591,N_2544);
xor U2671 (N_2671,N_2600,N_2599);
and U2672 (N_2672,N_2589,N_2574);
xor U2673 (N_2673,N_2542,N_2527);
nand U2674 (N_2674,N_2571,N_2607);
nand U2675 (N_2675,N_2538,N_2500);
nor U2676 (N_2676,N_2516,N_2614);
nor U2677 (N_2677,N_2557,N_2517);
xor U2678 (N_2678,N_2521,N_2526);
nand U2679 (N_2679,N_2566,N_2570);
nand U2680 (N_2680,N_2507,N_2573);
nor U2681 (N_2681,N_2535,N_2576);
nand U2682 (N_2682,N_2505,N_2615);
xnor U2683 (N_2683,N_2553,N_2594);
nand U2684 (N_2684,N_2562,N_2577);
nand U2685 (N_2685,N_2608,N_2568);
and U2686 (N_2686,N_2593,N_2624);
xnor U2687 (N_2687,N_2522,N_2508);
nor U2688 (N_2688,N_2556,N_2606);
xor U2689 (N_2689,N_2504,N_2599);
xor U2690 (N_2690,N_2606,N_2566);
or U2691 (N_2691,N_2526,N_2578);
and U2692 (N_2692,N_2567,N_2534);
nand U2693 (N_2693,N_2597,N_2524);
nand U2694 (N_2694,N_2512,N_2600);
or U2695 (N_2695,N_2531,N_2609);
or U2696 (N_2696,N_2585,N_2519);
or U2697 (N_2697,N_2550,N_2533);
or U2698 (N_2698,N_2510,N_2536);
nor U2699 (N_2699,N_2503,N_2521);
nand U2700 (N_2700,N_2513,N_2533);
nand U2701 (N_2701,N_2587,N_2543);
nor U2702 (N_2702,N_2521,N_2530);
xor U2703 (N_2703,N_2579,N_2600);
or U2704 (N_2704,N_2613,N_2517);
xor U2705 (N_2705,N_2611,N_2529);
or U2706 (N_2706,N_2506,N_2621);
xor U2707 (N_2707,N_2592,N_2617);
or U2708 (N_2708,N_2542,N_2540);
or U2709 (N_2709,N_2501,N_2590);
and U2710 (N_2710,N_2540,N_2512);
xnor U2711 (N_2711,N_2581,N_2561);
nor U2712 (N_2712,N_2512,N_2572);
xnor U2713 (N_2713,N_2505,N_2530);
nand U2714 (N_2714,N_2591,N_2572);
and U2715 (N_2715,N_2502,N_2606);
nor U2716 (N_2716,N_2506,N_2596);
or U2717 (N_2717,N_2524,N_2622);
and U2718 (N_2718,N_2510,N_2550);
or U2719 (N_2719,N_2608,N_2570);
or U2720 (N_2720,N_2522,N_2584);
and U2721 (N_2721,N_2512,N_2525);
or U2722 (N_2722,N_2521,N_2571);
xor U2723 (N_2723,N_2560,N_2605);
or U2724 (N_2724,N_2502,N_2526);
nor U2725 (N_2725,N_2602,N_2564);
and U2726 (N_2726,N_2564,N_2598);
nand U2727 (N_2727,N_2545,N_2510);
xnor U2728 (N_2728,N_2533,N_2597);
or U2729 (N_2729,N_2619,N_2530);
and U2730 (N_2730,N_2584,N_2559);
and U2731 (N_2731,N_2534,N_2615);
nand U2732 (N_2732,N_2506,N_2570);
nor U2733 (N_2733,N_2560,N_2606);
nand U2734 (N_2734,N_2506,N_2575);
and U2735 (N_2735,N_2546,N_2607);
and U2736 (N_2736,N_2544,N_2582);
and U2737 (N_2737,N_2508,N_2576);
nor U2738 (N_2738,N_2547,N_2588);
xnor U2739 (N_2739,N_2593,N_2602);
xor U2740 (N_2740,N_2574,N_2596);
or U2741 (N_2741,N_2614,N_2604);
or U2742 (N_2742,N_2505,N_2534);
xnor U2743 (N_2743,N_2598,N_2614);
xnor U2744 (N_2744,N_2591,N_2588);
nor U2745 (N_2745,N_2550,N_2529);
or U2746 (N_2746,N_2562,N_2558);
and U2747 (N_2747,N_2582,N_2580);
nand U2748 (N_2748,N_2586,N_2556);
or U2749 (N_2749,N_2513,N_2550);
xnor U2750 (N_2750,N_2714,N_2682);
or U2751 (N_2751,N_2625,N_2695);
or U2752 (N_2752,N_2707,N_2648);
and U2753 (N_2753,N_2705,N_2700);
and U2754 (N_2754,N_2637,N_2634);
or U2755 (N_2755,N_2679,N_2687);
nor U2756 (N_2756,N_2745,N_2702);
xor U2757 (N_2757,N_2749,N_2657);
xnor U2758 (N_2758,N_2631,N_2704);
and U2759 (N_2759,N_2706,N_2680);
or U2760 (N_2760,N_2727,N_2711);
or U2761 (N_2761,N_2661,N_2746);
nand U2762 (N_2762,N_2676,N_2710);
or U2763 (N_2763,N_2653,N_2670);
or U2764 (N_2764,N_2739,N_2668);
nand U2765 (N_2765,N_2662,N_2681);
xor U2766 (N_2766,N_2658,N_2688);
nand U2767 (N_2767,N_2719,N_2630);
nand U2768 (N_2768,N_2717,N_2722);
nor U2769 (N_2769,N_2674,N_2667);
and U2770 (N_2770,N_2747,N_2652);
nand U2771 (N_2771,N_2659,N_2744);
nand U2772 (N_2772,N_2693,N_2684);
or U2773 (N_2773,N_2708,N_2715);
and U2774 (N_2774,N_2642,N_2728);
xnor U2775 (N_2775,N_2703,N_2692);
or U2776 (N_2776,N_2701,N_2633);
nand U2777 (N_2777,N_2683,N_2641);
and U2778 (N_2778,N_2685,N_2632);
and U2779 (N_2779,N_2736,N_2650);
nor U2780 (N_2780,N_2643,N_2742);
xnor U2781 (N_2781,N_2656,N_2644);
nor U2782 (N_2782,N_2748,N_2636);
and U2783 (N_2783,N_2729,N_2665);
xor U2784 (N_2784,N_2645,N_2698);
or U2785 (N_2785,N_2664,N_2699);
nor U2786 (N_2786,N_2639,N_2732);
and U2787 (N_2787,N_2626,N_2627);
nand U2788 (N_2788,N_2669,N_2694);
nor U2789 (N_2789,N_2638,N_2716);
and U2790 (N_2790,N_2696,N_2628);
or U2791 (N_2791,N_2690,N_2723);
and U2792 (N_2792,N_2646,N_2629);
nand U2793 (N_2793,N_2671,N_2660);
or U2794 (N_2794,N_2725,N_2709);
xnor U2795 (N_2795,N_2743,N_2635);
and U2796 (N_2796,N_2673,N_2666);
or U2797 (N_2797,N_2649,N_2735);
nor U2798 (N_2798,N_2724,N_2686);
nand U2799 (N_2799,N_2689,N_2730);
xnor U2800 (N_2800,N_2733,N_2731);
and U2801 (N_2801,N_2655,N_2720);
nand U2802 (N_2802,N_2713,N_2738);
nand U2803 (N_2803,N_2737,N_2640);
or U2804 (N_2804,N_2678,N_2718);
or U2805 (N_2805,N_2651,N_2726);
or U2806 (N_2806,N_2721,N_2712);
nor U2807 (N_2807,N_2734,N_2741);
xor U2808 (N_2808,N_2697,N_2675);
nor U2809 (N_2809,N_2647,N_2740);
nor U2810 (N_2810,N_2691,N_2677);
nand U2811 (N_2811,N_2654,N_2672);
and U2812 (N_2812,N_2663,N_2674);
and U2813 (N_2813,N_2714,N_2676);
or U2814 (N_2814,N_2703,N_2644);
and U2815 (N_2815,N_2731,N_2684);
nor U2816 (N_2816,N_2736,N_2677);
or U2817 (N_2817,N_2702,N_2676);
nand U2818 (N_2818,N_2727,N_2738);
xnor U2819 (N_2819,N_2697,N_2736);
or U2820 (N_2820,N_2734,N_2729);
or U2821 (N_2821,N_2678,N_2724);
or U2822 (N_2822,N_2733,N_2670);
or U2823 (N_2823,N_2742,N_2626);
or U2824 (N_2824,N_2726,N_2739);
nor U2825 (N_2825,N_2748,N_2663);
nand U2826 (N_2826,N_2634,N_2749);
and U2827 (N_2827,N_2704,N_2685);
nand U2828 (N_2828,N_2717,N_2649);
xnor U2829 (N_2829,N_2714,N_2636);
and U2830 (N_2830,N_2634,N_2734);
or U2831 (N_2831,N_2628,N_2728);
and U2832 (N_2832,N_2651,N_2642);
nand U2833 (N_2833,N_2732,N_2745);
and U2834 (N_2834,N_2638,N_2720);
nor U2835 (N_2835,N_2645,N_2734);
and U2836 (N_2836,N_2683,N_2701);
and U2837 (N_2837,N_2704,N_2682);
or U2838 (N_2838,N_2742,N_2699);
nand U2839 (N_2839,N_2721,N_2743);
or U2840 (N_2840,N_2733,N_2745);
nand U2841 (N_2841,N_2710,N_2654);
nand U2842 (N_2842,N_2739,N_2727);
and U2843 (N_2843,N_2725,N_2666);
or U2844 (N_2844,N_2652,N_2703);
xor U2845 (N_2845,N_2633,N_2651);
and U2846 (N_2846,N_2678,N_2730);
or U2847 (N_2847,N_2676,N_2729);
nor U2848 (N_2848,N_2666,N_2710);
and U2849 (N_2849,N_2690,N_2743);
xor U2850 (N_2850,N_2684,N_2643);
nor U2851 (N_2851,N_2653,N_2654);
and U2852 (N_2852,N_2703,N_2645);
nor U2853 (N_2853,N_2656,N_2628);
or U2854 (N_2854,N_2699,N_2641);
and U2855 (N_2855,N_2734,N_2632);
nand U2856 (N_2856,N_2701,N_2737);
nor U2857 (N_2857,N_2655,N_2740);
xor U2858 (N_2858,N_2735,N_2730);
nor U2859 (N_2859,N_2684,N_2666);
and U2860 (N_2860,N_2642,N_2702);
xnor U2861 (N_2861,N_2679,N_2720);
xor U2862 (N_2862,N_2634,N_2666);
xnor U2863 (N_2863,N_2726,N_2717);
or U2864 (N_2864,N_2673,N_2650);
nand U2865 (N_2865,N_2647,N_2706);
xor U2866 (N_2866,N_2745,N_2647);
nor U2867 (N_2867,N_2637,N_2697);
or U2868 (N_2868,N_2640,N_2746);
and U2869 (N_2869,N_2628,N_2726);
nor U2870 (N_2870,N_2698,N_2633);
nor U2871 (N_2871,N_2635,N_2724);
nand U2872 (N_2872,N_2639,N_2716);
and U2873 (N_2873,N_2679,N_2650);
nand U2874 (N_2874,N_2715,N_2701);
xnor U2875 (N_2875,N_2822,N_2821);
or U2876 (N_2876,N_2862,N_2802);
and U2877 (N_2877,N_2838,N_2750);
nand U2878 (N_2878,N_2858,N_2786);
or U2879 (N_2879,N_2801,N_2847);
nor U2880 (N_2880,N_2871,N_2792);
xor U2881 (N_2881,N_2850,N_2845);
and U2882 (N_2882,N_2760,N_2874);
nand U2883 (N_2883,N_2853,N_2754);
nor U2884 (N_2884,N_2791,N_2798);
nor U2885 (N_2885,N_2873,N_2859);
and U2886 (N_2886,N_2826,N_2811);
or U2887 (N_2887,N_2755,N_2774);
or U2888 (N_2888,N_2825,N_2766);
and U2889 (N_2889,N_2863,N_2815);
or U2890 (N_2890,N_2833,N_2848);
xnor U2891 (N_2891,N_2816,N_2856);
nor U2892 (N_2892,N_2780,N_2790);
nor U2893 (N_2893,N_2849,N_2767);
nand U2894 (N_2894,N_2860,N_2776);
and U2895 (N_2895,N_2857,N_2819);
or U2896 (N_2896,N_2793,N_2828);
and U2897 (N_2897,N_2830,N_2762);
nor U2898 (N_2898,N_2832,N_2800);
nor U2899 (N_2899,N_2779,N_2770);
nand U2900 (N_2900,N_2768,N_2757);
or U2901 (N_2901,N_2788,N_2806);
nand U2902 (N_2902,N_2820,N_2783);
and U2903 (N_2903,N_2843,N_2759);
nor U2904 (N_2904,N_2872,N_2855);
nand U2905 (N_2905,N_2807,N_2772);
nor U2906 (N_2906,N_2851,N_2799);
nor U2907 (N_2907,N_2829,N_2869);
nor U2908 (N_2908,N_2787,N_2784);
or U2909 (N_2909,N_2814,N_2778);
nand U2910 (N_2910,N_2756,N_2823);
nor U2911 (N_2911,N_2868,N_2804);
or U2912 (N_2912,N_2824,N_2752);
and U2913 (N_2913,N_2846,N_2865);
or U2914 (N_2914,N_2782,N_2769);
or U2915 (N_2915,N_2864,N_2773);
nor U2916 (N_2916,N_2866,N_2867);
or U2917 (N_2917,N_2809,N_2831);
xnor U2918 (N_2918,N_2777,N_2781);
xor U2919 (N_2919,N_2844,N_2861);
or U2920 (N_2920,N_2870,N_2771);
nand U2921 (N_2921,N_2797,N_2834);
nor U2922 (N_2922,N_2805,N_2854);
or U2923 (N_2923,N_2764,N_2841);
xnor U2924 (N_2924,N_2842,N_2758);
and U2925 (N_2925,N_2818,N_2836);
nand U2926 (N_2926,N_2813,N_2751);
nand U2927 (N_2927,N_2763,N_2785);
xor U2928 (N_2928,N_2840,N_2837);
or U2929 (N_2929,N_2803,N_2852);
or U2930 (N_2930,N_2794,N_2835);
nor U2931 (N_2931,N_2795,N_2761);
nor U2932 (N_2932,N_2789,N_2839);
and U2933 (N_2933,N_2808,N_2796);
nor U2934 (N_2934,N_2765,N_2812);
and U2935 (N_2935,N_2753,N_2810);
nor U2936 (N_2936,N_2827,N_2775);
xor U2937 (N_2937,N_2817,N_2801);
and U2938 (N_2938,N_2791,N_2863);
xor U2939 (N_2939,N_2833,N_2807);
and U2940 (N_2940,N_2795,N_2809);
xnor U2941 (N_2941,N_2758,N_2786);
xor U2942 (N_2942,N_2763,N_2861);
xor U2943 (N_2943,N_2777,N_2799);
or U2944 (N_2944,N_2776,N_2834);
nand U2945 (N_2945,N_2812,N_2783);
or U2946 (N_2946,N_2772,N_2860);
nand U2947 (N_2947,N_2760,N_2841);
nor U2948 (N_2948,N_2865,N_2794);
nor U2949 (N_2949,N_2774,N_2845);
or U2950 (N_2950,N_2782,N_2872);
nand U2951 (N_2951,N_2819,N_2864);
xor U2952 (N_2952,N_2853,N_2838);
nand U2953 (N_2953,N_2752,N_2871);
or U2954 (N_2954,N_2863,N_2818);
nor U2955 (N_2955,N_2768,N_2857);
nand U2956 (N_2956,N_2783,N_2801);
or U2957 (N_2957,N_2785,N_2816);
nor U2958 (N_2958,N_2776,N_2813);
and U2959 (N_2959,N_2804,N_2829);
nor U2960 (N_2960,N_2799,N_2776);
nand U2961 (N_2961,N_2874,N_2863);
or U2962 (N_2962,N_2855,N_2853);
nand U2963 (N_2963,N_2754,N_2845);
nand U2964 (N_2964,N_2839,N_2790);
nor U2965 (N_2965,N_2812,N_2817);
or U2966 (N_2966,N_2798,N_2841);
and U2967 (N_2967,N_2836,N_2860);
or U2968 (N_2968,N_2857,N_2792);
nand U2969 (N_2969,N_2807,N_2842);
nand U2970 (N_2970,N_2860,N_2750);
or U2971 (N_2971,N_2854,N_2796);
or U2972 (N_2972,N_2868,N_2818);
and U2973 (N_2973,N_2763,N_2782);
xnor U2974 (N_2974,N_2869,N_2872);
nand U2975 (N_2975,N_2787,N_2789);
and U2976 (N_2976,N_2823,N_2804);
xnor U2977 (N_2977,N_2872,N_2779);
nand U2978 (N_2978,N_2852,N_2771);
and U2979 (N_2979,N_2765,N_2786);
xnor U2980 (N_2980,N_2866,N_2790);
nand U2981 (N_2981,N_2813,N_2864);
or U2982 (N_2982,N_2843,N_2820);
and U2983 (N_2983,N_2846,N_2754);
and U2984 (N_2984,N_2868,N_2807);
nand U2985 (N_2985,N_2868,N_2851);
and U2986 (N_2986,N_2812,N_2835);
and U2987 (N_2987,N_2761,N_2790);
or U2988 (N_2988,N_2775,N_2812);
and U2989 (N_2989,N_2814,N_2822);
and U2990 (N_2990,N_2759,N_2841);
and U2991 (N_2991,N_2764,N_2856);
nand U2992 (N_2992,N_2774,N_2828);
nand U2993 (N_2993,N_2750,N_2780);
or U2994 (N_2994,N_2829,N_2853);
xor U2995 (N_2995,N_2787,N_2774);
nor U2996 (N_2996,N_2839,N_2871);
or U2997 (N_2997,N_2754,N_2833);
xor U2998 (N_2998,N_2809,N_2760);
nor U2999 (N_2999,N_2868,N_2863);
nand U3000 (N_3000,N_2916,N_2915);
or U3001 (N_3001,N_2983,N_2879);
and U3002 (N_3002,N_2901,N_2882);
and U3003 (N_3003,N_2949,N_2965);
nor U3004 (N_3004,N_2903,N_2975);
nor U3005 (N_3005,N_2981,N_2957);
xnor U3006 (N_3006,N_2988,N_2911);
and U3007 (N_3007,N_2907,N_2942);
nor U3008 (N_3008,N_2927,N_2997);
and U3009 (N_3009,N_2960,N_2996);
and U3010 (N_3010,N_2945,N_2888);
and U3011 (N_3011,N_2920,N_2939);
nor U3012 (N_3012,N_2971,N_2946);
xnor U3013 (N_3013,N_2897,N_2961);
and U3014 (N_3014,N_2919,N_2885);
nor U3015 (N_3015,N_2998,N_2964);
nand U3016 (N_3016,N_2953,N_2900);
or U3017 (N_3017,N_2967,N_2954);
nor U3018 (N_3018,N_2928,N_2896);
and U3019 (N_3019,N_2973,N_2962);
xnor U3020 (N_3020,N_2922,N_2979);
xor U3021 (N_3021,N_2895,N_2958);
xor U3022 (N_3022,N_2972,N_2930);
nand U3023 (N_3023,N_2969,N_2952);
nand U3024 (N_3024,N_2877,N_2898);
nor U3025 (N_3025,N_2985,N_2974);
nor U3026 (N_3026,N_2935,N_2899);
or U3027 (N_3027,N_2984,N_2918);
or U3028 (N_3028,N_2932,N_2948);
nor U3029 (N_3029,N_2941,N_2880);
nor U3030 (N_3030,N_2884,N_2940);
nand U3031 (N_3031,N_2914,N_2990);
or U3032 (N_3032,N_2943,N_2937);
or U3033 (N_3033,N_2950,N_2933);
xnor U3034 (N_3034,N_2970,N_2992);
nor U3035 (N_3035,N_2994,N_2980);
xor U3036 (N_3036,N_2966,N_2878);
or U3037 (N_3037,N_2959,N_2881);
xnor U3038 (N_3038,N_2923,N_2883);
nor U3039 (N_3039,N_2987,N_2904);
nor U3040 (N_3040,N_2989,N_2912);
and U3041 (N_3041,N_2906,N_2889);
and U3042 (N_3042,N_2931,N_2934);
and U3043 (N_3043,N_2956,N_2910);
xor U3044 (N_3044,N_2993,N_2894);
nor U3045 (N_3045,N_2929,N_2947);
and U3046 (N_3046,N_2908,N_2925);
xnor U3047 (N_3047,N_2955,N_2976);
nand U3048 (N_3048,N_2909,N_2876);
or U3049 (N_3049,N_2887,N_2951);
and U3050 (N_3050,N_2986,N_2982);
and U3051 (N_3051,N_2886,N_2890);
or U3052 (N_3052,N_2905,N_2944);
and U3053 (N_3053,N_2913,N_2963);
and U3054 (N_3054,N_2924,N_2893);
or U3055 (N_3055,N_2921,N_2938);
xnor U3056 (N_3056,N_2926,N_2991);
or U3057 (N_3057,N_2936,N_2968);
and U3058 (N_3058,N_2977,N_2978);
nor U3059 (N_3059,N_2995,N_2999);
nor U3060 (N_3060,N_2875,N_2891);
xor U3061 (N_3061,N_2917,N_2902);
xnor U3062 (N_3062,N_2892,N_2957);
nand U3063 (N_3063,N_2879,N_2966);
nand U3064 (N_3064,N_2934,N_2963);
and U3065 (N_3065,N_2953,N_2948);
nand U3066 (N_3066,N_2893,N_2996);
xor U3067 (N_3067,N_2929,N_2942);
nor U3068 (N_3068,N_2951,N_2921);
xor U3069 (N_3069,N_2983,N_2958);
xor U3070 (N_3070,N_2996,N_2969);
nor U3071 (N_3071,N_2988,N_2970);
xor U3072 (N_3072,N_2878,N_2877);
xor U3073 (N_3073,N_2992,N_2916);
and U3074 (N_3074,N_2903,N_2885);
and U3075 (N_3075,N_2928,N_2878);
and U3076 (N_3076,N_2905,N_2940);
xor U3077 (N_3077,N_2881,N_2965);
nand U3078 (N_3078,N_2949,N_2936);
or U3079 (N_3079,N_2883,N_2895);
and U3080 (N_3080,N_2897,N_2986);
xnor U3081 (N_3081,N_2924,N_2950);
or U3082 (N_3082,N_2911,N_2949);
nor U3083 (N_3083,N_2882,N_2903);
xor U3084 (N_3084,N_2949,N_2993);
nor U3085 (N_3085,N_2934,N_2906);
xor U3086 (N_3086,N_2944,N_2875);
or U3087 (N_3087,N_2937,N_2905);
nor U3088 (N_3088,N_2990,N_2971);
and U3089 (N_3089,N_2954,N_2957);
xnor U3090 (N_3090,N_2967,N_2992);
nor U3091 (N_3091,N_2945,N_2943);
nor U3092 (N_3092,N_2908,N_2918);
and U3093 (N_3093,N_2894,N_2981);
nand U3094 (N_3094,N_2961,N_2917);
nor U3095 (N_3095,N_2956,N_2963);
and U3096 (N_3096,N_2880,N_2886);
nand U3097 (N_3097,N_2917,N_2896);
and U3098 (N_3098,N_2927,N_2977);
or U3099 (N_3099,N_2926,N_2892);
xnor U3100 (N_3100,N_2962,N_2916);
xor U3101 (N_3101,N_2901,N_2941);
and U3102 (N_3102,N_2961,N_2959);
nor U3103 (N_3103,N_2963,N_2939);
or U3104 (N_3104,N_2947,N_2959);
nor U3105 (N_3105,N_2939,N_2908);
nand U3106 (N_3106,N_2877,N_2984);
xnor U3107 (N_3107,N_2956,N_2946);
or U3108 (N_3108,N_2922,N_2895);
and U3109 (N_3109,N_2899,N_2967);
or U3110 (N_3110,N_2897,N_2908);
or U3111 (N_3111,N_2888,N_2900);
nand U3112 (N_3112,N_2915,N_2925);
nand U3113 (N_3113,N_2989,N_2891);
or U3114 (N_3114,N_2906,N_2951);
nor U3115 (N_3115,N_2913,N_2936);
xor U3116 (N_3116,N_2941,N_2995);
nand U3117 (N_3117,N_2899,N_2903);
or U3118 (N_3118,N_2945,N_2886);
or U3119 (N_3119,N_2983,N_2992);
or U3120 (N_3120,N_2979,N_2914);
nand U3121 (N_3121,N_2918,N_2969);
and U3122 (N_3122,N_2905,N_2966);
and U3123 (N_3123,N_2972,N_2928);
nor U3124 (N_3124,N_2918,N_2914);
xor U3125 (N_3125,N_3040,N_3048);
and U3126 (N_3126,N_3075,N_3026);
nand U3127 (N_3127,N_3007,N_3120);
and U3128 (N_3128,N_3116,N_3091);
nand U3129 (N_3129,N_3098,N_3093);
nor U3130 (N_3130,N_3101,N_3035);
xor U3131 (N_3131,N_3059,N_3025);
and U3132 (N_3132,N_3060,N_3013);
and U3133 (N_3133,N_3081,N_3003);
and U3134 (N_3134,N_3084,N_3062);
or U3135 (N_3135,N_3045,N_3119);
xor U3136 (N_3136,N_3011,N_3115);
xor U3137 (N_3137,N_3089,N_3055);
nand U3138 (N_3138,N_3010,N_3124);
nor U3139 (N_3139,N_3073,N_3009);
and U3140 (N_3140,N_3018,N_3014);
or U3141 (N_3141,N_3042,N_3051);
nand U3142 (N_3142,N_3108,N_3032);
or U3143 (N_3143,N_3123,N_3106);
nand U3144 (N_3144,N_3076,N_3004);
nor U3145 (N_3145,N_3069,N_3020);
and U3146 (N_3146,N_3029,N_3005);
and U3147 (N_3147,N_3087,N_3114);
nor U3148 (N_3148,N_3057,N_3046);
nand U3149 (N_3149,N_3015,N_3067);
and U3150 (N_3150,N_3061,N_3041);
and U3151 (N_3151,N_3028,N_3037);
and U3152 (N_3152,N_3117,N_3111);
or U3153 (N_3153,N_3053,N_3094);
or U3154 (N_3154,N_3002,N_3070);
nor U3155 (N_3155,N_3085,N_3049);
or U3156 (N_3156,N_3109,N_3024);
and U3157 (N_3157,N_3065,N_3110);
or U3158 (N_3158,N_3099,N_3064);
xor U3159 (N_3159,N_3052,N_3031);
or U3160 (N_3160,N_3021,N_3056);
and U3161 (N_3161,N_3122,N_3030);
xor U3162 (N_3162,N_3012,N_3092);
or U3163 (N_3163,N_3066,N_3090);
xnor U3164 (N_3164,N_3027,N_3113);
xor U3165 (N_3165,N_3078,N_3107);
xor U3166 (N_3166,N_3100,N_3086);
xor U3167 (N_3167,N_3121,N_3112);
and U3168 (N_3168,N_3033,N_3036);
nor U3169 (N_3169,N_3097,N_3017);
and U3170 (N_3170,N_3006,N_3063);
or U3171 (N_3171,N_3054,N_3039);
or U3172 (N_3172,N_3043,N_3104);
and U3173 (N_3173,N_3102,N_3071);
and U3174 (N_3174,N_3008,N_3105);
and U3175 (N_3175,N_3016,N_3074);
nor U3176 (N_3176,N_3072,N_3023);
or U3177 (N_3177,N_3038,N_3080);
and U3178 (N_3178,N_3068,N_3047);
and U3179 (N_3179,N_3096,N_3058);
nand U3180 (N_3180,N_3019,N_3000);
nor U3181 (N_3181,N_3050,N_3082);
nor U3182 (N_3182,N_3118,N_3095);
xor U3183 (N_3183,N_3088,N_3079);
or U3184 (N_3184,N_3077,N_3103);
or U3185 (N_3185,N_3001,N_3044);
nor U3186 (N_3186,N_3022,N_3083);
xnor U3187 (N_3187,N_3034,N_3019);
or U3188 (N_3188,N_3002,N_3113);
nor U3189 (N_3189,N_3066,N_3116);
or U3190 (N_3190,N_3007,N_3023);
nor U3191 (N_3191,N_3077,N_3099);
xnor U3192 (N_3192,N_3103,N_3076);
xnor U3193 (N_3193,N_3002,N_3015);
nand U3194 (N_3194,N_3096,N_3063);
xor U3195 (N_3195,N_3086,N_3087);
nand U3196 (N_3196,N_3086,N_3080);
xnor U3197 (N_3197,N_3112,N_3073);
nand U3198 (N_3198,N_3114,N_3044);
or U3199 (N_3199,N_3027,N_3105);
nor U3200 (N_3200,N_3049,N_3006);
nand U3201 (N_3201,N_3087,N_3074);
and U3202 (N_3202,N_3034,N_3064);
nand U3203 (N_3203,N_3061,N_3019);
xnor U3204 (N_3204,N_3068,N_3106);
nand U3205 (N_3205,N_3055,N_3079);
or U3206 (N_3206,N_3088,N_3064);
nor U3207 (N_3207,N_3043,N_3070);
nand U3208 (N_3208,N_3113,N_3074);
xnor U3209 (N_3209,N_3007,N_3067);
or U3210 (N_3210,N_3116,N_3030);
nand U3211 (N_3211,N_3046,N_3088);
nor U3212 (N_3212,N_3041,N_3105);
xor U3213 (N_3213,N_3093,N_3051);
xor U3214 (N_3214,N_3109,N_3075);
nor U3215 (N_3215,N_3031,N_3065);
nand U3216 (N_3216,N_3058,N_3027);
and U3217 (N_3217,N_3053,N_3116);
and U3218 (N_3218,N_3009,N_3092);
xor U3219 (N_3219,N_3090,N_3003);
nor U3220 (N_3220,N_3077,N_3031);
and U3221 (N_3221,N_3086,N_3084);
nor U3222 (N_3222,N_3017,N_3014);
and U3223 (N_3223,N_3104,N_3107);
nand U3224 (N_3224,N_3119,N_3070);
nor U3225 (N_3225,N_3091,N_3081);
or U3226 (N_3226,N_3032,N_3073);
nand U3227 (N_3227,N_3083,N_3046);
and U3228 (N_3228,N_3076,N_3045);
and U3229 (N_3229,N_3074,N_3066);
or U3230 (N_3230,N_3088,N_3119);
and U3231 (N_3231,N_3004,N_3106);
or U3232 (N_3232,N_3034,N_3001);
nor U3233 (N_3233,N_3119,N_3008);
nand U3234 (N_3234,N_3117,N_3021);
nor U3235 (N_3235,N_3053,N_3016);
nor U3236 (N_3236,N_3102,N_3031);
and U3237 (N_3237,N_3118,N_3036);
xor U3238 (N_3238,N_3013,N_3084);
and U3239 (N_3239,N_3055,N_3025);
or U3240 (N_3240,N_3067,N_3081);
nand U3241 (N_3241,N_3022,N_3107);
nor U3242 (N_3242,N_3033,N_3006);
and U3243 (N_3243,N_3026,N_3106);
and U3244 (N_3244,N_3012,N_3032);
xnor U3245 (N_3245,N_3103,N_3017);
nand U3246 (N_3246,N_3076,N_3097);
nor U3247 (N_3247,N_3117,N_3032);
nand U3248 (N_3248,N_3048,N_3015);
or U3249 (N_3249,N_3012,N_3050);
xnor U3250 (N_3250,N_3140,N_3158);
nand U3251 (N_3251,N_3244,N_3131);
or U3252 (N_3252,N_3172,N_3247);
or U3253 (N_3253,N_3141,N_3211);
and U3254 (N_3254,N_3183,N_3249);
xnor U3255 (N_3255,N_3219,N_3170);
and U3256 (N_3256,N_3215,N_3130);
or U3257 (N_3257,N_3159,N_3194);
xnor U3258 (N_3258,N_3163,N_3237);
and U3259 (N_3259,N_3205,N_3182);
or U3260 (N_3260,N_3236,N_3226);
nand U3261 (N_3261,N_3225,N_3148);
or U3262 (N_3262,N_3238,N_3241);
or U3263 (N_3263,N_3229,N_3231);
nand U3264 (N_3264,N_3185,N_3196);
and U3265 (N_3265,N_3144,N_3217);
and U3266 (N_3266,N_3227,N_3228);
and U3267 (N_3267,N_3221,N_3125);
xnor U3268 (N_3268,N_3129,N_3186);
nor U3269 (N_3269,N_3188,N_3150);
and U3270 (N_3270,N_3192,N_3223);
nand U3271 (N_3271,N_3179,N_3127);
xnor U3272 (N_3272,N_3166,N_3209);
xor U3273 (N_3273,N_3137,N_3126);
or U3274 (N_3274,N_3146,N_3195);
or U3275 (N_3275,N_3178,N_3191);
or U3276 (N_3276,N_3245,N_3175);
or U3277 (N_3277,N_3128,N_3153);
and U3278 (N_3278,N_3152,N_3207);
nor U3279 (N_3279,N_3160,N_3136);
nand U3280 (N_3280,N_3190,N_3233);
or U3281 (N_3281,N_3212,N_3216);
and U3282 (N_3282,N_3210,N_3214);
nand U3283 (N_3283,N_3218,N_3248);
and U3284 (N_3284,N_3142,N_3246);
or U3285 (N_3285,N_3174,N_3168);
xor U3286 (N_3286,N_3134,N_3222);
or U3287 (N_3287,N_3187,N_3177);
or U3288 (N_3288,N_3198,N_3138);
or U3289 (N_3289,N_3235,N_3173);
and U3290 (N_3290,N_3180,N_3242);
or U3291 (N_3291,N_3243,N_3147);
xor U3292 (N_3292,N_3201,N_3240);
and U3293 (N_3293,N_3230,N_3213);
xor U3294 (N_3294,N_3232,N_3189);
and U3295 (N_3295,N_3200,N_3206);
or U3296 (N_3296,N_3165,N_3167);
and U3297 (N_3297,N_3176,N_3169);
and U3298 (N_3298,N_3143,N_3184);
nand U3299 (N_3299,N_3204,N_3224);
nand U3300 (N_3300,N_3162,N_3203);
and U3301 (N_3301,N_3149,N_3155);
and U3302 (N_3302,N_3145,N_3157);
xor U3303 (N_3303,N_3208,N_3156);
and U3304 (N_3304,N_3202,N_3133);
nor U3305 (N_3305,N_3239,N_3139);
and U3306 (N_3306,N_3151,N_3164);
nand U3307 (N_3307,N_3154,N_3197);
or U3308 (N_3308,N_3199,N_3193);
or U3309 (N_3309,N_3181,N_3220);
xor U3310 (N_3310,N_3161,N_3234);
xor U3311 (N_3311,N_3132,N_3171);
nand U3312 (N_3312,N_3135,N_3242);
nand U3313 (N_3313,N_3175,N_3210);
nand U3314 (N_3314,N_3128,N_3143);
nor U3315 (N_3315,N_3190,N_3197);
xnor U3316 (N_3316,N_3174,N_3132);
or U3317 (N_3317,N_3128,N_3139);
and U3318 (N_3318,N_3174,N_3157);
xor U3319 (N_3319,N_3223,N_3199);
xnor U3320 (N_3320,N_3246,N_3140);
nor U3321 (N_3321,N_3188,N_3130);
and U3322 (N_3322,N_3140,N_3145);
nor U3323 (N_3323,N_3194,N_3215);
or U3324 (N_3324,N_3201,N_3163);
or U3325 (N_3325,N_3167,N_3151);
or U3326 (N_3326,N_3204,N_3138);
xor U3327 (N_3327,N_3209,N_3133);
nand U3328 (N_3328,N_3242,N_3248);
nor U3329 (N_3329,N_3133,N_3242);
xnor U3330 (N_3330,N_3135,N_3198);
or U3331 (N_3331,N_3133,N_3162);
and U3332 (N_3332,N_3220,N_3134);
and U3333 (N_3333,N_3168,N_3238);
and U3334 (N_3334,N_3164,N_3245);
nand U3335 (N_3335,N_3221,N_3181);
nand U3336 (N_3336,N_3205,N_3160);
xnor U3337 (N_3337,N_3165,N_3173);
xnor U3338 (N_3338,N_3167,N_3126);
nor U3339 (N_3339,N_3203,N_3156);
and U3340 (N_3340,N_3193,N_3243);
xor U3341 (N_3341,N_3143,N_3172);
xor U3342 (N_3342,N_3141,N_3164);
nand U3343 (N_3343,N_3188,N_3204);
nand U3344 (N_3344,N_3130,N_3183);
nand U3345 (N_3345,N_3167,N_3164);
nand U3346 (N_3346,N_3137,N_3155);
and U3347 (N_3347,N_3223,N_3146);
and U3348 (N_3348,N_3153,N_3139);
or U3349 (N_3349,N_3205,N_3129);
nand U3350 (N_3350,N_3243,N_3218);
nand U3351 (N_3351,N_3211,N_3221);
and U3352 (N_3352,N_3133,N_3174);
and U3353 (N_3353,N_3192,N_3240);
xor U3354 (N_3354,N_3235,N_3143);
and U3355 (N_3355,N_3225,N_3170);
and U3356 (N_3356,N_3145,N_3141);
and U3357 (N_3357,N_3202,N_3148);
nor U3358 (N_3358,N_3244,N_3158);
or U3359 (N_3359,N_3219,N_3131);
nor U3360 (N_3360,N_3176,N_3167);
or U3361 (N_3361,N_3237,N_3139);
or U3362 (N_3362,N_3179,N_3244);
nand U3363 (N_3363,N_3218,N_3234);
and U3364 (N_3364,N_3187,N_3167);
nor U3365 (N_3365,N_3125,N_3164);
xnor U3366 (N_3366,N_3249,N_3178);
xnor U3367 (N_3367,N_3149,N_3229);
or U3368 (N_3368,N_3140,N_3176);
nor U3369 (N_3369,N_3146,N_3188);
and U3370 (N_3370,N_3200,N_3161);
and U3371 (N_3371,N_3207,N_3170);
and U3372 (N_3372,N_3244,N_3202);
and U3373 (N_3373,N_3219,N_3220);
nor U3374 (N_3374,N_3225,N_3149);
and U3375 (N_3375,N_3304,N_3301);
and U3376 (N_3376,N_3312,N_3255);
xor U3377 (N_3377,N_3278,N_3279);
nor U3378 (N_3378,N_3261,N_3257);
nor U3379 (N_3379,N_3330,N_3299);
or U3380 (N_3380,N_3265,N_3311);
or U3381 (N_3381,N_3339,N_3315);
and U3382 (N_3382,N_3251,N_3262);
nor U3383 (N_3383,N_3294,N_3324);
or U3384 (N_3384,N_3317,N_3291);
xor U3385 (N_3385,N_3270,N_3296);
or U3386 (N_3386,N_3292,N_3367);
or U3387 (N_3387,N_3309,N_3276);
or U3388 (N_3388,N_3325,N_3268);
nand U3389 (N_3389,N_3346,N_3253);
nor U3390 (N_3390,N_3345,N_3374);
and U3391 (N_3391,N_3342,N_3281);
or U3392 (N_3392,N_3308,N_3333);
nand U3393 (N_3393,N_3359,N_3297);
and U3394 (N_3394,N_3365,N_3335);
nand U3395 (N_3395,N_3254,N_3344);
or U3396 (N_3396,N_3316,N_3290);
nor U3397 (N_3397,N_3372,N_3258);
nand U3398 (N_3398,N_3352,N_3250);
nand U3399 (N_3399,N_3334,N_3322);
nand U3400 (N_3400,N_3373,N_3332);
xor U3401 (N_3401,N_3306,N_3313);
and U3402 (N_3402,N_3277,N_3267);
xor U3403 (N_3403,N_3310,N_3326);
nand U3404 (N_3404,N_3269,N_3369);
nor U3405 (N_3405,N_3314,N_3273);
xor U3406 (N_3406,N_3289,N_3356);
and U3407 (N_3407,N_3363,N_3275);
and U3408 (N_3408,N_3327,N_3295);
xor U3409 (N_3409,N_3364,N_3368);
nor U3410 (N_3410,N_3321,N_3272);
nand U3411 (N_3411,N_3357,N_3338);
and U3412 (N_3412,N_3348,N_3293);
nor U3413 (N_3413,N_3302,N_3288);
xnor U3414 (N_3414,N_3271,N_3260);
xnor U3415 (N_3415,N_3264,N_3266);
nor U3416 (N_3416,N_3328,N_3337);
nor U3417 (N_3417,N_3303,N_3358);
or U3418 (N_3418,N_3280,N_3274);
xor U3419 (N_3419,N_3361,N_3347);
or U3420 (N_3420,N_3319,N_3331);
and U3421 (N_3421,N_3362,N_3343);
and U3422 (N_3422,N_3351,N_3341);
nor U3423 (N_3423,N_3298,N_3336);
nor U3424 (N_3424,N_3371,N_3286);
nor U3425 (N_3425,N_3329,N_3283);
and U3426 (N_3426,N_3300,N_3360);
nand U3427 (N_3427,N_3366,N_3259);
nand U3428 (N_3428,N_3340,N_3285);
or U3429 (N_3429,N_3263,N_3284);
xor U3430 (N_3430,N_3307,N_3252);
nor U3431 (N_3431,N_3305,N_3287);
xor U3432 (N_3432,N_3282,N_3353);
and U3433 (N_3433,N_3355,N_3323);
and U3434 (N_3434,N_3318,N_3349);
nor U3435 (N_3435,N_3320,N_3354);
nand U3436 (N_3436,N_3370,N_3350);
nand U3437 (N_3437,N_3256,N_3250);
or U3438 (N_3438,N_3286,N_3336);
or U3439 (N_3439,N_3264,N_3300);
or U3440 (N_3440,N_3256,N_3323);
nor U3441 (N_3441,N_3297,N_3318);
xnor U3442 (N_3442,N_3346,N_3295);
and U3443 (N_3443,N_3344,N_3310);
nand U3444 (N_3444,N_3355,N_3270);
nor U3445 (N_3445,N_3305,N_3336);
xor U3446 (N_3446,N_3362,N_3287);
xnor U3447 (N_3447,N_3329,N_3274);
and U3448 (N_3448,N_3321,N_3288);
nor U3449 (N_3449,N_3307,N_3320);
xnor U3450 (N_3450,N_3292,N_3333);
nand U3451 (N_3451,N_3372,N_3370);
nand U3452 (N_3452,N_3323,N_3320);
nand U3453 (N_3453,N_3350,N_3277);
nand U3454 (N_3454,N_3344,N_3306);
nor U3455 (N_3455,N_3315,N_3290);
or U3456 (N_3456,N_3374,N_3311);
xnor U3457 (N_3457,N_3293,N_3354);
nand U3458 (N_3458,N_3268,N_3280);
nor U3459 (N_3459,N_3254,N_3331);
or U3460 (N_3460,N_3305,N_3343);
or U3461 (N_3461,N_3274,N_3316);
or U3462 (N_3462,N_3307,N_3319);
or U3463 (N_3463,N_3316,N_3358);
nand U3464 (N_3464,N_3270,N_3267);
nand U3465 (N_3465,N_3307,N_3369);
nand U3466 (N_3466,N_3316,N_3327);
nand U3467 (N_3467,N_3269,N_3250);
nand U3468 (N_3468,N_3337,N_3264);
xor U3469 (N_3469,N_3255,N_3267);
or U3470 (N_3470,N_3275,N_3265);
xnor U3471 (N_3471,N_3344,N_3267);
nand U3472 (N_3472,N_3272,N_3341);
xnor U3473 (N_3473,N_3373,N_3308);
nor U3474 (N_3474,N_3263,N_3309);
or U3475 (N_3475,N_3260,N_3327);
or U3476 (N_3476,N_3343,N_3326);
nor U3477 (N_3477,N_3319,N_3338);
nor U3478 (N_3478,N_3317,N_3367);
xor U3479 (N_3479,N_3334,N_3256);
or U3480 (N_3480,N_3294,N_3295);
xnor U3481 (N_3481,N_3344,N_3342);
nor U3482 (N_3482,N_3364,N_3336);
or U3483 (N_3483,N_3275,N_3278);
or U3484 (N_3484,N_3357,N_3347);
and U3485 (N_3485,N_3359,N_3312);
nor U3486 (N_3486,N_3329,N_3282);
nand U3487 (N_3487,N_3293,N_3320);
or U3488 (N_3488,N_3270,N_3256);
nand U3489 (N_3489,N_3259,N_3355);
nand U3490 (N_3490,N_3268,N_3299);
xnor U3491 (N_3491,N_3282,N_3307);
xnor U3492 (N_3492,N_3367,N_3285);
nor U3493 (N_3493,N_3341,N_3286);
nor U3494 (N_3494,N_3312,N_3321);
and U3495 (N_3495,N_3288,N_3374);
nor U3496 (N_3496,N_3362,N_3272);
nor U3497 (N_3497,N_3257,N_3256);
xnor U3498 (N_3498,N_3292,N_3254);
nor U3499 (N_3499,N_3340,N_3297);
and U3500 (N_3500,N_3440,N_3452);
and U3501 (N_3501,N_3448,N_3376);
or U3502 (N_3502,N_3477,N_3499);
nor U3503 (N_3503,N_3444,N_3435);
and U3504 (N_3504,N_3425,N_3472);
nor U3505 (N_3505,N_3410,N_3466);
nand U3506 (N_3506,N_3380,N_3432);
or U3507 (N_3507,N_3388,N_3485);
nor U3508 (N_3508,N_3465,N_3497);
or U3509 (N_3509,N_3384,N_3389);
or U3510 (N_3510,N_3430,N_3375);
or U3511 (N_3511,N_3421,N_3399);
or U3512 (N_3512,N_3428,N_3447);
nor U3513 (N_3513,N_3438,N_3488);
nor U3514 (N_3514,N_3392,N_3473);
or U3515 (N_3515,N_3489,N_3431);
or U3516 (N_3516,N_3442,N_3419);
or U3517 (N_3517,N_3398,N_3397);
nand U3518 (N_3518,N_3385,N_3457);
and U3519 (N_3519,N_3411,N_3403);
xor U3520 (N_3520,N_3391,N_3394);
nor U3521 (N_3521,N_3422,N_3451);
or U3522 (N_3522,N_3417,N_3481);
or U3523 (N_3523,N_3426,N_3407);
or U3524 (N_3524,N_3436,N_3483);
xnor U3525 (N_3525,N_3406,N_3445);
xnor U3526 (N_3526,N_3454,N_3402);
or U3527 (N_3527,N_3458,N_3460);
or U3528 (N_3528,N_3416,N_3487);
nor U3529 (N_3529,N_3490,N_3495);
or U3530 (N_3530,N_3378,N_3462);
nand U3531 (N_3531,N_3491,N_3474);
xor U3532 (N_3532,N_3382,N_3449);
nand U3533 (N_3533,N_3441,N_3455);
nand U3534 (N_3534,N_3401,N_3479);
xor U3535 (N_3535,N_3467,N_3492);
xor U3536 (N_3536,N_3482,N_3446);
or U3537 (N_3537,N_3461,N_3476);
nor U3538 (N_3538,N_3470,N_3450);
and U3539 (N_3539,N_3456,N_3478);
or U3540 (N_3540,N_3409,N_3433);
nor U3541 (N_3541,N_3439,N_3393);
nand U3542 (N_3542,N_3443,N_3434);
and U3543 (N_3543,N_3464,N_3396);
and U3544 (N_3544,N_3423,N_3437);
nand U3545 (N_3545,N_3414,N_3420);
nor U3546 (N_3546,N_3379,N_3424);
nand U3547 (N_3547,N_3453,N_3475);
nor U3548 (N_3548,N_3383,N_3387);
and U3549 (N_3549,N_3390,N_3377);
or U3550 (N_3550,N_3484,N_3486);
nand U3551 (N_3551,N_3408,N_3386);
xnor U3552 (N_3552,N_3405,N_3395);
and U3553 (N_3553,N_3494,N_3429);
and U3554 (N_3554,N_3415,N_3413);
nor U3555 (N_3555,N_3498,N_3381);
xnor U3556 (N_3556,N_3493,N_3468);
xnor U3557 (N_3557,N_3418,N_3469);
or U3558 (N_3558,N_3496,N_3459);
nand U3559 (N_3559,N_3471,N_3400);
or U3560 (N_3560,N_3412,N_3427);
and U3561 (N_3561,N_3463,N_3480);
xor U3562 (N_3562,N_3404,N_3394);
nand U3563 (N_3563,N_3469,N_3492);
xnor U3564 (N_3564,N_3499,N_3433);
xor U3565 (N_3565,N_3440,N_3425);
and U3566 (N_3566,N_3452,N_3406);
nor U3567 (N_3567,N_3377,N_3430);
nor U3568 (N_3568,N_3441,N_3409);
or U3569 (N_3569,N_3433,N_3403);
xor U3570 (N_3570,N_3448,N_3457);
or U3571 (N_3571,N_3390,N_3421);
and U3572 (N_3572,N_3477,N_3402);
nand U3573 (N_3573,N_3443,N_3467);
and U3574 (N_3574,N_3411,N_3468);
xnor U3575 (N_3575,N_3434,N_3465);
and U3576 (N_3576,N_3425,N_3383);
and U3577 (N_3577,N_3416,N_3462);
and U3578 (N_3578,N_3466,N_3435);
nand U3579 (N_3579,N_3378,N_3487);
nor U3580 (N_3580,N_3483,N_3495);
xnor U3581 (N_3581,N_3479,N_3496);
nor U3582 (N_3582,N_3425,N_3393);
and U3583 (N_3583,N_3487,N_3462);
or U3584 (N_3584,N_3386,N_3394);
xor U3585 (N_3585,N_3416,N_3414);
and U3586 (N_3586,N_3436,N_3404);
nor U3587 (N_3587,N_3471,N_3458);
xnor U3588 (N_3588,N_3483,N_3474);
nand U3589 (N_3589,N_3488,N_3380);
or U3590 (N_3590,N_3475,N_3469);
nand U3591 (N_3591,N_3455,N_3377);
nor U3592 (N_3592,N_3426,N_3488);
xnor U3593 (N_3593,N_3463,N_3483);
nor U3594 (N_3594,N_3387,N_3424);
xor U3595 (N_3595,N_3406,N_3398);
or U3596 (N_3596,N_3485,N_3428);
xnor U3597 (N_3597,N_3427,N_3431);
xnor U3598 (N_3598,N_3466,N_3473);
or U3599 (N_3599,N_3445,N_3474);
nor U3600 (N_3600,N_3464,N_3459);
nor U3601 (N_3601,N_3483,N_3439);
nand U3602 (N_3602,N_3446,N_3479);
nor U3603 (N_3603,N_3405,N_3436);
nand U3604 (N_3604,N_3398,N_3499);
and U3605 (N_3605,N_3389,N_3404);
and U3606 (N_3606,N_3494,N_3407);
nor U3607 (N_3607,N_3473,N_3460);
xnor U3608 (N_3608,N_3462,N_3485);
and U3609 (N_3609,N_3452,N_3482);
or U3610 (N_3610,N_3386,N_3477);
nand U3611 (N_3611,N_3473,N_3464);
nand U3612 (N_3612,N_3451,N_3458);
and U3613 (N_3613,N_3406,N_3391);
nand U3614 (N_3614,N_3379,N_3417);
xnor U3615 (N_3615,N_3498,N_3473);
xor U3616 (N_3616,N_3403,N_3445);
and U3617 (N_3617,N_3414,N_3442);
nand U3618 (N_3618,N_3432,N_3478);
and U3619 (N_3619,N_3420,N_3405);
or U3620 (N_3620,N_3475,N_3478);
nand U3621 (N_3621,N_3462,N_3389);
nor U3622 (N_3622,N_3489,N_3386);
nor U3623 (N_3623,N_3402,N_3483);
nor U3624 (N_3624,N_3426,N_3466);
nand U3625 (N_3625,N_3611,N_3614);
nand U3626 (N_3626,N_3590,N_3610);
and U3627 (N_3627,N_3523,N_3600);
or U3628 (N_3628,N_3511,N_3571);
nor U3629 (N_3629,N_3572,N_3503);
and U3630 (N_3630,N_3609,N_3547);
nand U3631 (N_3631,N_3607,N_3588);
or U3632 (N_3632,N_3550,N_3556);
nor U3633 (N_3633,N_3591,N_3531);
and U3634 (N_3634,N_3502,N_3530);
xor U3635 (N_3635,N_3592,N_3535);
nand U3636 (N_3636,N_3622,N_3606);
or U3637 (N_3637,N_3562,N_3568);
nand U3638 (N_3638,N_3524,N_3534);
or U3639 (N_3639,N_3520,N_3576);
nand U3640 (N_3640,N_3578,N_3595);
xnor U3641 (N_3641,N_3537,N_3546);
nor U3642 (N_3642,N_3623,N_3549);
or U3643 (N_3643,N_3616,N_3510);
nor U3644 (N_3644,N_3528,N_3594);
nand U3645 (N_3645,N_3565,N_3620);
and U3646 (N_3646,N_3533,N_3564);
nand U3647 (N_3647,N_3601,N_3604);
nand U3648 (N_3648,N_3559,N_3573);
nor U3649 (N_3649,N_3599,N_3612);
xor U3650 (N_3650,N_3508,N_3555);
or U3651 (N_3651,N_3536,N_3558);
or U3652 (N_3652,N_3596,N_3589);
xnor U3653 (N_3653,N_3522,N_3529);
or U3654 (N_3654,N_3618,N_3552);
xnor U3655 (N_3655,N_3527,N_3624);
nand U3656 (N_3656,N_3526,N_3563);
nor U3657 (N_3657,N_3541,N_3539);
and U3658 (N_3658,N_3551,N_3515);
nand U3659 (N_3659,N_3575,N_3542);
or U3660 (N_3660,N_3506,N_3574);
nand U3661 (N_3661,N_3521,N_3593);
xnor U3662 (N_3662,N_3605,N_3514);
and U3663 (N_3663,N_3580,N_3587);
nor U3664 (N_3664,N_3519,N_3567);
and U3665 (N_3665,N_3516,N_3615);
and U3666 (N_3666,N_3570,N_3543);
and U3667 (N_3667,N_3548,N_3617);
nor U3668 (N_3668,N_3585,N_3557);
and U3669 (N_3669,N_3544,N_3561);
nand U3670 (N_3670,N_3598,N_3619);
xor U3671 (N_3671,N_3608,N_3540);
nand U3672 (N_3672,N_3554,N_3613);
xnor U3673 (N_3673,N_3500,N_3525);
and U3674 (N_3674,N_3577,N_3603);
and U3675 (N_3675,N_3602,N_3581);
or U3676 (N_3676,N_3507,N_3501);
and U3677 (N_3677,N_3579,N_3597);
and U3678 (N_3678,N_3584,N_3566);
and U3679 (N_3679,N_3621,N_3545);
or U3680 (N_3680,N_3504,N_3569);
xor U3681 (N_3681,N_3517,N_3505);
nor U3682 (N_3682,N_3538,N_3582);
and U3683 (N_3683,N_3583,N_3560);
or U3684 (N_3684,N_3512,N_3553);
nor U3685 (N_3685,N_3513,N_3586);
or U3686 (N_3686,N_3509,N_3518);
xor U3687 (N_3687,N_3532,N_3502);
nand U3688 (N_3688,N_3623,N_3509);
or U3689 (N_3689,N_3595,N_3609);
nand U3690 (N_3690,N_3622,N_3546);
nor U3691 (N_3691,N_3558,N_3616);
nor U3692 (N_3692,N_3567,N_3607);
or U3693 (N_3693,N_3578,N_3573);
xor U3694 (N_3694,N_3516,N_3601);
xnor U3695 (N_3695,N_3616,N_3597);
or U3696 (N_3696,N_3513,N_3506);
nor U3697 (N_3697,N_3586,N_3512);
or U3698 (N_3698,N_3608,N_3593);
or U3699 (N_3699,N_3614,N_3548);
or U3700 (N_3700,N_3514,N_3567);
nor U3701 (N_3701,N_3516,N_3540);
xnor U3702 (N_3702,N_3589,N_3562);
nor U3703 (N_3703,N_3606,N_3602);
xor U3704 (N_3704,N_3580,N_3545);
and U3705 (N_3705,N_3506,N_3575);
nor U3706 (N_3706,N_3527,N_3571);
xor U3707 (N_3707,N_3587,N_3577);
or U3708 (N_3708,N_3617,N_3615);
xor U3709 (N_3709,N_3619,N_3553);
or U3710 (N_3710,N_3582,N_3618);
nor U3711 (N_3711,N_3542,N_3613);
nor U3712 (N_3712,N_3595,N_3612);
or U3713 (N_3713,N_3624,N_3617);
xnor U3714 (N_3714,N_3618,N_3535);
nor U3715 (N_3715,N_3549,N_3535);
and U3716 (N_3716,N_3601,N_3608);
nor U3717 (N_3717,N_3534,N_3596);
nor U3718 (N_3718,N_3578,N_3553);
and U3719 (N_3719,N_3614,N_3580);
and U3720 (N_3720,N_3532,N_3533);
nor U3721 (N_3721,N_3516,N_3506);
or U3722 (N_3722,N_3525,N_3604);
and U3723 (N_3723,N_3518,N_3536);
nor U3724 (N_3724,N_3549,N_3601);
xor U3725 (N_3725,N_3563,N_3539);
xnor U3726 (N_3726,N_3527,N_3504);
nor U3727 (N_3727,N_3549,N_3572);
nand U3728 (N_3728,N_3556,N_3621);
nor U3729 (N_3729,N_3540,N_3620);
nor U3730 (N_3730,N_3602,N_3571);
nor U3731 (N_3731,N_3576,N_3514);
nor U3732 (N_3732,N_3516,N_3588);
nand U3733 (N_3733,N_3601,N_3546);
xnor U3734 (N_3734,N_3589,N_3518);
nor U3735 (N_3735,N_3618,N_3539);
and U3736 (N_3736,N_3505,N_3605);
xor U3737 (N_3737,N_3503,N_3606);
nor U3738 (N_3738,N_3502,N_3554);
and U3739 (N_3739,N_3611,N_3551);
and U3740 (N_3740,N_3542,N_3547);
xor U3741 (N_3741,N_3553,N_3533);
or U3742 (N_3742,N_3503,N_3506);
or U3743 (N_3743,N_3537,N_3563);
nor U3744 (N_3744,N_3610,N_3573);
or U3745 (N_3745,N_3611,N_3607);
or U3746 (N_3746,N_3530,N_3515);
nor U3747 (N_3747,N_3618,N_3508);
nor U3748 (N_3748,N_3503,N_3513);
and U3749 (N_3749,N_3568,N_3503);
nor U3750 (N_3750,N_3669,N_3743);
nor U3751 (N_3751,N_3665,N_3663);
or U3752 (N_3752,N_3685,N_3659);
or U3753 (N_3753,N_3668,N_3634);
and U3754 (N_3754,N_3637,N_3684);
nor U3755 (N_3755,N_3735,N_3734);
and U3756 (N_3756,N_3626,N_3651);
xor U3757 (N_3757,N_3691,N_3713);
nand U3758 (N_3758,N_3690,N_3656);
or U3759 (N_3759,N_3701,N_3687);
or U3760 (N_3760,N_3672,N_3712);
nand U3761 (N_3761,N_3740,N_3636);
nand U3762 (N_3762,N_3653,N_3658);
or U3763 (N_3763,N_3662,N_3689);
nor U3764 (N_3764,N_3698,N_3670);
and U3765 (N_3765,N_3650,N_3729);
nor U3766 (N_3766,N_3652,N_3639);
and U3767 (N_3767,N_3741,N_3705);
nor U3768 (N_3768,N_3686,N_3746);
nand U3769 (N_3769,N_3649,N_3676);
and U3770 (N_3770,N_3654,N_3661);
and U3771 (N_3771,N_3696,N_3707);
and U3772 (N_3772,N_3648,N_3719);
and U3773 (N_3773,N_3709,N_3688);
nand U3774 (N_3774,N_3633,N_3694);
and U3775 (N_3775,N_3703,N_3657);
nor U3776 (N_3776,N_3716,N_3682);
xor U3777 (N_3777,N_3715,N_3644);
nor U3778 (N_3778,N_3680,N_3660);
xor U3779 (N_3779,N_3631,N_3630);
xor U3780 (N_3780,N_3679,N_3722);
nor U3781 (N_3781,N_3711,N_3635);
nor U3782 (N_3782,N_3738,N_3732);
xor U3783 (N_3783,N_3748,N_3728);
nor U3784 (N_3784,N_3717,N_3692);
nand U3785 (N_3785,N_3744,N_3641);
nand U3786 (N_3786,N_3693,N_3667);
and U3787 (N_3787,N_3706,N_3697);
nand U3788 (N_3788,N_3643,N_3745);
and U3789 (N_3789,N_3723,N_3724);
xor U3790 (N_3790,N_3671,N_3645);
or U3791 (N_3791,N_3721,N_3675);
and U3792 (N_3792,N_3625,N_3733);
and U3793 (N_3793,N_3677,N_3683);
and U3794 (N_3794,N_3695,N_3655);
and U3795 (N_3795,N_3726,N_3749);
nand U3796 (N_3796,N_3731,N_3730);
nor U3797 (N_3797,N_3628,N_3666);
nor U3798 (N_3798,N_3646,N_3642);
nor U3799 (N_3799,N_3629,N_3673);
nor U3800 (N_3800,N_3627,N_3708);
nor U3801 (N_3801,N_3702,N_3718);
nor U3802 (N_3802,N_3725,N_3647);
nand U3803 (N_3803,N_3742,N_3640);
nor U3804 (N_3804,N_3674,N_3737);
nand U3805 (N_3805,N_3704,N_3678);
nand U3806 (N_3806,N_3714,N_3736);
or U3807 (N_3807,N_3727,N_3664);
xnor U3808 (N_3808,N_3700,N_3699);
nor U3809 (N_3809,N_3747,N_3638);
and U3810 (N_3810,N_3632,N_3710);
nand U3811 (N_3811,N_3739,N_3720);
nor U3812 (N_3812,N_3681,N_3692);
or U3813 (N_3813,N_3717,N_3638);
xnor U3814 (N_3814,N_3695,N_3694);
nor U3815 (N_3815,N_3720,N_3731);
xnor U3816 (N_3816,N_3699,N_3651);
nor U3817 (N_3817,N_3647,N_3631);
nor U3818 (N_3818,N_3648,N_3632);
nor U3819 (N_3819,N_3668,N_3701);
nand U3820 (N_3820,N_3659,N_3697);
xor U3821 (N_3821,N_3645,N_3670);
or U3822 (N_3822,N_3747,N_3669);
nand U3823 (N_3823,N_3744,N_3630);
nand U3824 (N_3824,N_3628,N_3656);
and U3825 (N_3825,N_3687,N_3735);
nor U3826 (N_3826,N_3645,N_3675);
nand U3827 (N_3827,N_3664,N_3707);
xnor U3828 (N_3828,N_3730,N_3627);
nor U3829 (N_3829,N_3648,N_3635);
or U3830 (N_3830,N_3641,N_3691);
or U3831 (N_3831,N_3626,N_3631);
xor U3832 (N_3832,N_3734,N_3684);
and U3833 (N_3833,N_3704,N_3655);
xnor U3834 (N_3834,N_3681,N_3660);
nand U3835 (N_3835,N_3642,N_3710);
xor U3836 (N_3836,N_3718,N_3721);
or U3837 (N_3837,N_3645,N_3700);
or U3838 (N_3838,N_3744,N_3644);
nand U3839 (N_3839,N_3742,N_3660);
or U3840 (N_3840,N_3740,N_3663);
xnor U3841 (N_3841,N_3686,N_3650);
or U3842 (N_3842,N_3626,N_3700);
nor U3843 (N_3843,N_3717,N_3712);
and U3844 (N_3844,N_3738,N_3676);
xnor U3845 (N_3845,N_3725,N_3669);
nor U3846 (N_3846,N_3670,N_3709);
nand U3847 (N_3847,N_3682,N_3701);
nand U3848 (N_3848,N_3703,N_3742);
nor U3849 (N_3849,N_3724,N_3657);
and U3850 (N_3850,N_3683,N_3666);
or U3851 (N_3851,N_3681,N_3629);
nand U3852 (N_3852,N_3673,N_3724);
nand U3853 (N_3853,N_3709,N_3695);
nand U3854 (N_3854,N_3677,N_3705);
nor U3855 (N_3855,N_3662,N_3656);
nand U3856 (N_3856,N_3717,N_3629);
nor U3857 (N_3857,N_3660,N_3687);
xnor U3858 (N_3858,N_3726,N_3660);
or U3859 (N_3859,N_3704,N_3657);
or U3860 (N_3860,N_3636,N_3717);
xor U3861 (N_3861,N_3698,N_3747);
xor U3862 (N_3862,N_3712,N_3749);
and U3863 (N_3863,N_3666,N_3679);
nand U3864 (N_3864,N_3627,N_3630);
nand U3865 (N_3865,N_3680,N_3748);
nor U3866 (N_3866,N_3645,N_3697);
nor U3867 (N_3867,N_3734,N_3741);
xnor U3868 (N_3868,N_3669,N_3667);
nor U3869 (N_3869,N_3722,N_3632);
xor U3870 (N_3870,N_3626,N_3721);
or U3871 (N_3871,N_3720,N_3660);
or U3872 (N_3872,N_3643,N_3698);
nand U3873 (N_3873,N_3628,N_3704);
and U3874 (N_3874,N_3685,N_3698);
and U3875 (N_3875,N_3817,N_3777);
xnor U3876 (N_3876,N_3872,N_3838);
and U3877 (N_3877,N_3860,N_3802);
and U3878 (N_3878,N_3796,N_3867);
or U3879 (N_3879,N_3836,N_3840);
and U3880 (N_3880,N_3770,N_3847);
nand U3881 (N_3881,N_3816,N_3789);
nand U3882 (N_3882,N_3807,N_3805);
or U3883 (N_3883,N_3823,N_3843);
and U3884 (N_3884,N_3791,N_3773);
nor U3885 (N_3885,N_3835,N_3839);
and U3886 (N_3886,N_3788,N_3768);
xor U3887 (N_3887,N_3818,N_3819);
or U3888 (N_3888,N_3866,N_3795);
nand U3889 (N_3889,N_3824,N_3855);
xor U3890 (N_3890,N_3756,N_3798);
nand U3891 (N_3891,N_3842,N_3794);
nor U3892 (N_3892,N_3810,N_3772);
and U3893 (N_3893,N_3859,N_3830);
nor U3894 (N_3894,N_3752,N_3760);
xnor U3895 (N_3895,N_3787,N_3856);
or U3896 (N_3896,N_3779,N_3755);
and U3897 (N_3897,N_3766,N_3797);
nand U3898 (N_3898,N_3869,N_3828);
or U3899 (N_3899,N_3769,N_3775);
nand U3900 (N_3900,N_3845,N_3833);
and U3901 (N_3901,N_3870,N_3774);
xnor U3902 (N_3902,N_3849,N_3783);
nor U3903 (N_3903,N_3785,N_3829);
or U3904 (N_3904,N_3864,N_3868);
nand U3905 (N_3905,N_3753,N_3861);
or U3906 (N_3906,N_3808,N_3832);
nand U3907 (N_3907,N_3801,N_3762);
and U3908 (N_3908,N_3800,N_3792);
nand U3909 (N_3909,N_3822,N_3811);
and U3910 (N_3910,N_3793,N_3821);
nand U3911 (N_3911,N_3825,N_3831);
xor U3912 (N_3912,N_3764,N_3809);
nor U3913 (N_3913,N_3862,N_3765);
nor U3914 (N_3914,N_3781,N_3812);
nor U3915 (N_3915,N_3790,N_3786);
nor U3916 (N_3916,N_3767,N_3776);
nand U3917 (N_3917,N_3863,N_3757);
xnor U3918 (N_3918,N_3761,N_3803);
nor U3919 (N_3919,N_3754,N_3782);
nor U3920 (N_3920,N_3763,N_3851);
or U3921 (N_3921,N_3844,N_3778);
nor U3922 (N_3922,N_3814,N_3871);
or U3923 (N_3923,N_3837,N_3751);
nor U3924 (N_3924,N_3799,N_3780);
xor U3925 (N_3925,N_3841,N_3750);
xnor U3926 (N_3926,N_3852,N_3865);
xnor U3927 (N_3927,N_3813,N_3826);
or U3928 (N_3928,N_3804,N_3758);
or U3929 (N_3929,N_3846,N_3857);
nand U3930 (N_3930,N_3771,N_3854);
or U3931 (N_3931,N_3759,N_3873);
and U3932 (N_3932,N_3834,N_3874);
or U3933 (N_3933,N_3848,N_3858);
nand U3934 (N_3934,N_3820,N_3806);
nand U3935 (N_3935,N_3827,N_3784);
xnor U3936 (N_3936,N_3815,N_3853);
and U3937 (N_3937,N_3850,N_3798);
xor U3938 (N_3938,N_3874,N_3869);
and U3939 (N_3939,N_3807,N_3832);
nand U3940 (N_3940,N_3842,N_3757);
and U3941 (N_3941,N_3776,N_3836);
and U3942 (N_3942,N_3835,N_3836);
xnor U3943 (N_3943,N_3813,N_3807);
nand U3944 (N_3944,N_3868,N_3858);
xnor U3945 (N_3945,N_3800,N_3771);
xor U3946 (N_3946,N_3849,N_3751);
or U3947 (N_3947,N_3798,N_3844);
and U3948 (N_3948,N_3863,N_3758);
and U3949 (N_3949,N_3790,N_3777);
nor U3950 (N_3950,N_3823,N_3846);
or U3951 (N_3951,N_3763,N_3750);
nor U3952 (N_3952,N_3778,N_3766);
xnor U3953 (N_3953,N_3820,N_3755);
nand U3954 (N_3954,N_3788,N_3824);
and U3955 (N_3955,N_3830,N_3823);
nor U3956 (N_3956,N_3757,N_3824);
xor U3957 (N_3957,N_3775,N_3869);
nor U3958 (N_3958,N_3863,N_3778);
nand U3959 (N_3959,N_3809,N_3862);
xor U3960 (N_3960,N_3867,N_3795);
and U3961 (N_3961,N_3851,N_3812);
xnor U3962 (N_3962,N_3751,N_3772);
and U3963 (N_3963,N_3857,N_3799);
xor U3964 (N_3964,N_3775,N_3761);
and U3965 (N_3965,N_3847,N_3816);
nand U3966 (N_3966,N_3793,N_3811);
xnor U3967 (N_3967,N_3867,N_3846);
xnor U3968 (N_3968,N_3786,N_3785);
xor U3969 (N_3969,N_3776,N_3853);
or U3970 (N_3970,N_3857,N_3786);
or U3971 (N_3971,N_3770,N_3759);
xor U3972 (N_3972,N_3850,N_3808);
nand U3973 (N_3973,N_3837,N_3766);
and U3974 (N_3974,N_3864,N_3863);
and U3975 (N_3975,N_3803,N_3769);
xnor U3976 (N_3976,N_3784,N_3755);
xnor U3977 (N_3977,N_3819,N_3784);
nor U3978 (N_3978,N_3774,N_3787);
nor U3979 (N_3979,N_3750,N_3826);
nand U3980 (N_3980,N_3843,N_3836);
and U3981 (N_3981,N_3772,N_3829);
and U3982 (N_3982,N_3863,N_3809);
nor U3983 (N_3983,N_3803,N_3782);
and U3984 (N_3984,N_3833,N_3785);
nand U3985 (N_3985,N_3865,N_3807);
nor U3986 (N_3986,N_3809,N_3777);
or U3987 (N_3987,N_3864,N_3770);
nand U3988 (N_3988,N_3854,N_3751);
or U3989 (N_3989,N_3801,N_3807);
and U3990 (N_3990,N_3766,N_3827);
xor U3991 (N_3991,N_3800,N_3812);
nor U3992 (N_3992,N_3821,N_3830);
and U3993 (N_3993,N_3811,N_3852);
nor U3994 (N_3994,N_3777,N_3827);
nor U3995 (N_3995,N_3828,N_3752);
nor U3996 (N_3996,N_3788,N_3765);
nor U3997 (N_3997,N_3762,N_3832);
and U3998 (N_3998,N_3839,N_3775);
nor U3999 (N_3999,N_3823,N_3860);
nand U4000 (N_4000,N_3988,N_3941);
and U4001 (N_4001,N_3924,N_3934);
or U4002 (N_4002,N_3887,N_3970);
xnor U4003 (N_4003,N_3906,N_3915);
and U4004 (N_4004,N_3935,N_3946);
or U4005 (N_4005,N_3967,N_3968);
nor U4006 (N_4006,N_3947,N_3897);
xnor U4007 (N_4007,N_3954,N_3990);
nand U4008 (N_4008,N_3945,N_3917);
nor U4009 (N_4009,N_3931,N_3922);
xnor U4010 (N_4010,N_3936,N_3949);
nand U4011 (N_4011,N_3888,N_3977);
nor U4012 (N_4012,N_3933,N_3926);
xor U4013 (N_4013,N_3901,N_3910);
xor U4014 (N_4014,N_3973,N_3983);
or U4015 (N_4015,N_3965,N_3994);
and U4016 (N_4016,N_3878,N_3944);
and U4017 (N_4017,N_3892,N_3991);
xnor U4018 (N_4018,N_3995,N_3918);
xor U4019 (N_4019,N_3951,N_3952);
nand U4020 (N_4020,N_3900,N_3928);
xnor U4021 (N_4021,N_3987,N_3920);
xor U4022 (N_4022,N_3879,N_3907);
xnor U4023 (N_4023,N_3989,N_3911);
nor U4024 (N_4024,N_3891,N_3895);
nor U4025 (N_4025,N_3963,N_3883);
nand U4026 (N_4026,N_3956,N_3916);
xnor U4027 (N_4027,N_3961,N_3993);
nor U4028 (N_4028,N_3962,N_3996);
or U4029 (N_4029,N_3974,N_3955);
nand U4030 (N_4030,N_3925,N_3903);
or U4031 (N_4031,N_3904,N_3981);
xnor U4032 (N_4032,N_3948,N_3882);
xor U4033 (N_4033,N_3953,N_3930);
nor U4034 (N_4034,N_3889,N_3921);
and U4035 (N_4035,N_3905,N_3942);
and U4036 (N_4036,N_3959,N_3884);
nor U4037 (N_4037,N_3880,N_3923);
xnor U4038 (N_4038,N_3937,N_3877);
and U4039 (N_4039,N_3982,N_3976);
or U4040 (N_4040,N_3908,N_3972);
and U4041 (N_4041,N_3978,N_3984);
and U4042 (N_4042,N_3890,N_3875);
and U4043 (N_4043,N_3985,N_3881);
xor U4044 (N_4044,N_3927,N_3999);
or U4045 (N_4045,N_3943,N_3898);
nand U4046 (N_4046,N_3966,N_3902);
nand U4047 (N_4047,N_3919,N_3894);
and U4048 (N_4048,N_3940,N_3997);
xnor U4049 (N_4049,N_3939,N_3957);
nor U4050 (N_4050,N_3876,N_3893);
or U4051 (N_4051,N_3885,N_3969);
nor U4052 (N_4052,N_3986,N_3979);
nor U4053 (N_4053,N_3899,N_3992);
xor U4054 (N_4054,N_3998,N_3932);
and U4055 (N_4055,N_3909,N_3971);
nor U4056 (N_4056,N_3964,N_3938);
nand U4057 (N_4057,N_3975,N_3913);
or U4058 (N_4058,N_3912,N_3950);
xnor U4059 (N_4059,N_3896,N_3960);
nor U4060 (N_4060,N_3958,N_3929);
and U4061 (N_4061,N_3980,N_3914);
and U4062 (N_4062,N_3886,N_3893);
or U4063 (N_4063,N_3922,N_3887);
or U4064 (N_4064,N_3883,N_3938);
nand U4065 (N_4065,N_3932,N_3908);
nand U4066 (N_4066,N_3989,N_3877);
and U4067 (N_4067,N_3928,N_3993);
or U4068 (N_4068,N_3938,N_3877);
nor U4069 (N_4069,N_3923,N_3878);
or U4070 (N_4070,N_3950,N_3965);
or U4071 (N_4071,N_3995,N_3881);
nor U4072 (N_4072,N_3936,N_3897);
or U4073 (N_4073,N_3905,N_3988);
or U4074 (N_4074,N_3947,N_3926);
nand U4075 (N_4075,N_3929,N_3919);
xor U4076 (N_4076,N_3941,N_3880);
nor U4077 (N_4077,N_3914,N_3999);
and U4078 (N_4078,N_3961,N_3976);
or U4079 (N_4079,N_3922,N_3947);
xnor U4080 (N_4080,N_3969,N_3991);
or U4081 (N_4081,N_3996,N_3882);
nor U4082 (N_4082,N_3875,N_3984);
and U4083 (N_4083,N_3896,N_3939);
nor U4084 (N_4084,N_3877,N_3984);
and U4085 (N_4085,N_3921,N_3993);
xor U4086 (N_4086,N_3972,N_3971);
xor U4087 (N_4087,N_3997,N_3932);
xor U4088 (N_4088,N_3995,N_3903);
nand U4089 (N_4089,N_3965,N_3897);
or U4090 (N_4090,N_3993,N_3883);
or U4091 (N_4091,N_3913,N_3936);
nand U4092 (N_4092,N_3916,N_3927);
and U4093 (N_4093,N_3961,N_3998);
xor U4094 (N_4094,N_3931,N_3978);
nand U4095 (N_4095,N_3885,N_3921);
and U4096 (N_4096,N_3994,N_3943);
xor U4097 (N_4097,N_3974,N_3969);
nor U4098 (N_4098,N_3980,N_3915);
nor U4099 (N_4099,N_3882,N_3898);
or U4100 (N_4100,N_3985,N_3970);
and U4101 (N_4101,N_3961,N_3949);
or U4102 (N_4102,N_3972,N_3952);
xor U4103 (N_4103,N_3964,N_3888);
xnor U4104 (N_4104,N_3914,N_3885);
and U4105 (N_4105,N_3890,N_3956);
and U4106 (N_4106,N_3947,N_3973);
xnor U4107 (N_4107,N_3977,N_3907);
nand U4108 (N_4108,N_3972,N_3960);
or U4109 (N_4109,N_3892,N_3943);
nor U4110 (N_4110,N_3930,N_3951);
and U4111 (N_4111,N_3934,N_3908);
or U4112 (N_4112,N_3964,N_3943);
nor U4113 (N_4113,N_3905,N_3920);
nand U4114 (N_4114,N_3915,N_3946);
and U4115 (N_4115,N_3992,N_3907);
nor U4116 (N_4116,N_3972,N_3955);
or U4117 (N_4117,N_3888,N_3966);
or U4118 (N_4118,N_3993,N_3965);
xnor U4119 (N_4119,N_3880,N_3896);
nand U4120 (N_4120,N_3949,N_3994);
nor U4121 (N_4121,N_3970,N_3980);
xor U4122 (N_4122,N_3914,N_3894);
xor U4123 (N_4123,N_3996,N_3955);
or U4124 (N_4124,N_3951,N_3955);
and U4125 (N_4125,N_4121,N_4090);
nand U4126 (N_4126,N_4094,N_4018);
and U4127 (N_4127,N_4076,N_4029);
and U4128 (N_4128,N_4039,N_4108);
xor U4129 (N_4129,N_4034,N_4114);
or U4130 (N_4130,N_4031,N_4104);
and U4131 (N_4131,N_4122,N_4019);
xor U4132 (N_4132,N_4096,N_4040);
nor U4133 (N_4133,N_4092,N_4097);
or U4134 (N_4134,N_4016,N_4058);
nand U4135 (N_4135,N_4075,N_4084);
xnor U4136 (N_4136,N_4071,N_4102);
nor U4137 (N_4137,N_4007,N_4059);
and U4138 (N_4138,N_4005,N_4107);
nand U4139 (N_4139,N_4116,N_4006);
or U4140 (N_4140,N_4026,N_4074);
nor U4141 (N_4141,N_4036,N_4078);
and U4142 (N_4142,N_4115,N_4060);
xor U4143 (N_4143,N_4064,N_4087);
nor U4144 (N_4144,N_4048,N_4027);
nand U4145 (N_4145,N_4095,N_4055);
xor U4146 (N_4146,N_4099,N_4035);
xnor U4147 (N_4147,N_4088,N_4014);
nand U4148 (N_4148,N_4054,N_4082);
nor U4149 (N_4149,N_4089,N_4083);
nor U4150 (N_4150,N_4008,N_4056);
or U4151 (N_4151,N_4119,N_4070);
nand U4152 (N_4152,N_4047,N_4004);
nand U4153 (N_4153,N_4021,N_4112);
nor U4154 (N_4154,N_4098,N_4003);
nor U4155 (N_4155,N_4022,N_4028);
nand U4156 (N_4156,N_4023,N_4010);
nand U4157 (N_4157,N_4067,N_4113);
nand U4158 (N_4158,N_4065,N_4117);
and U4159 (N_4159,N_4009,N_4015);
or U4160 (N_4160,N_4025,N_4063);
or U4161 (N_4161,N_4110,N_4000);
xor U4162 (N_4162,N_4043,N_4077);
nor U4163 (N_4163,N_4017,N_4086);
xnor U4164 (N_4164,N_4069,N_4002);
xnor U4165 (N_4165,N_4081,N_4066);
nor U4166 (N_4166,N_4053,N_4041);
or U4167 (N_4167,N_4050,N_4120);
or U4168 (N_4168,N_4032,N_4044);
or U4169 (N_4169,N_4052,N_4020);
nand U4170 (N_4170,N_4024,N_4072);
nor U4171 (N_4171,N_4037,N_4106);
or U4172 (N_4172,N_4051,N_4049);
xnor U4173 (N_4173,N_4013,N_4045);
and U4174 (N_4174,N_4079,N_4062);
and U4175 (N_4175,N_4001,N_4011);
nor U4176 (N_4176,N_4033,N_4080);
xor U4177 (N_4177,N_4101,N_4046);
or U4178 (N_4178,N_4038,N_4068);
or U4179 (N_4179,N_4118,N_4057);
and U4180 (N_4180,N_4085,N_4105);
xor U4181 (N_4181,N_4093,N_4091);
nor U4182 (N_4182,N_4109,N_4030);
xor U4183 (N_4183,N_4100,N_4012);
nor U4184 (N_4184,N_4042,N_4073);
and U4185 (N_4185,N_4123,N_4103);
nor U4186 (N_4186,N_4124,N_4111);
nand U4187 (N_4187,N_4061,N_4115);
xor U4188 (N_4188,N_4028,N_4056);
or U4189 (N_4189,N_4018,N_4067);
xnor U4190 (N_4190,N_4041,N_4090);
and U4191 (N_4191,N_4087,N_4027);
nand U4192 (N_4192,N_4111,N_4028);
and U4193 (N_4193,N_4110,N_4097);
nand U4194 (N_4194,N_4072,N_4112);
xnor U4195 (N_4195,N_4111,N_4066);
nor U4196 (N_4196,N_4023,N_4108);
nor U4197 (N_4197,N_4070,N_4036);
nand U4198 (N_4198,N_4015,N_4027);
or U4199 (N_4199,N_4051,N_4087);
and U4200 (N_4200,N_4109,N_4013);
nor U4201 (N_4201,N_4063,N_4086);
xor U4202 (N_4202,N_4101,N_4027);
nand U4203 (N_4203,N_4030,N_4098);
and U4204 (N_4204,N_4030,N_4115);
or U4205 (N_4205,N_4008,N_4068);
xor U4206 (N_4206,N_4020,N_4102);
nand U4207 (N_4207,N_4033,N_4029);
xor U4208 (N_4208,N_4038,N_4070);
nor U4209 (N_4209,N_4056,N_4030);
xor U4210 (N_4210,N_4007,N_4124);
nor U4211 (N_4211,N_4012,N_4089);
or U4212 (N_4212,N_4033,N_4085);
nand U4213 (N_4213,N_4011,N_4095);
nor U4214 (N_4214,N_4013,N_4084);
xnor U4215 (N_4215,N_4105,N_4084);
or U4216 (N_4216,N_4040,N_4054);
nand U4217 (N_4217,N_4115,N_4089);
nor U4218 (N_4218,N_4078,N_4023);
and U4219 (N_4219,N_4038,N_4035);
and U4220 (N_4220,N_4061,N_4040);
or U4221 (N_4221,N_4093,N_4025);
and U4222 (N_4222,N_4008,N_4074);
xnor U4223 (N_4223,N_4040,N_4105);
or U4224 (N_4224,N_4116,N_4107);
xnor U4225 (N_4225,N_4030,N_4081);
or U4226 (N_4226,N_4023,N_4022);
xor U4227 (N_4227,N_4081,N_4104);
nand U4228 (N_4228,N_4032,N_4066);
and U4229 (N_4229,N_4111,N_4039);
nor U4230 (N_4230,N_4079,N_4081);
or U4231 (N_4231,N_4105,N_4093);
xor U4232 (N_4232,N_4107,N_4077);
or U4233 (N_4233,N_4001,N_4086);
xnor U4234 (N_4234,N_4019,N_4082);
nand U4235 (N_4235,N_4049,N_4085);
or U4236 (N_4236,N_4049,N_4075);
nor U4237 (N_4237,N_4054,N_4045);
and U4238 (N_4238,N_4092,N_4070);
nand U4239 (N_4239,N_4079,N_4122);
nor U4240 (N_4240,N_4113,N_4045);
or U4241 (N_4241,N_4082,N_4009);
and U4242 (N_4242,N_4044,N_4014);
nor U4243 (N_4243,N_4001,N_4090);
and U4244 (N_4244,N_4096,N_4031);
and U4245 (N_4245,N_4107,N_4003);
and U4246 (N_4246,N_4045,N_4072);
xnor U4247 (N_4247,N_4120,N_4091);
and U4248 (N_4248,N_4091,N_4031);
xor U4249 (N_4249,N_4121,N_4030);
nand U4250 (N_4250,N_4148,N_4141);
and U4251 (N_4251,N_4202,N_4208);
xnor U4252 (N_4252,N_4126,N_4157);
or U4253 (N_4253,N_4171,N_4220);
or U4254 (N_4254,N_4209,N_4230);
and U4255 (N_4255,N_4164,N_4145);
nor U4256 (N_4256,N_4216,N_4215);
xor U4257 (N_4257,N_4237,N_4182);
nor U4258 (N_4258,N_4243,N_4205);
or U4259 (N_4259,N_4178,N_4140);
or U4260 (N_4260,N_4206,N_4218);
xor U4261 (N_4261,N_4161,N_4191);
or U4262 (N_4262,N_4244,N_4210);
nor U4263 (N_4263,N_4195,N_4173);
xnor U4264 (N_4264,N_4163,N_4127);
or U4265 (N_4265,N_4132,N_4165);
nor U4266 (N_4266,N_4174,N_4176);
nand U4267 (N_4267,N_4144,N_4128);
nor U4268 (N_4268,N_4185,N_4125);
xor U4269 (N_4269,N_4135,N_4188);
xor U4270 (N_4270,N_4151,N_4219);
and U4271 (N_4271,N_4226,N_4129);
nor U4272 (N_4272,N_4175,N_4196);
nor U4273 (N_4273,N_4180,N_4203);
xnor U4274 (N_4274,N_4130,N_4168);
and U4275 (N_4275,N_4194,N_4235);
or U4276 (N_4276,N_4149,N_4166);
or U4277 (N_4277,N_4142,N_4183);
nor U4278 (N_4278,N_4238,N_4192);
nor U4279 (N_4279,N_4233,N_4225);
nor U4280 (N_4280,N_4207,N_4227);
or U4281 (N_4281,N_4158,N_4241);
nor U4282 (N_4282,N_4187,N_4172);
and U4283 (N_4283,N_4181,N_4186);
or U4284 (N_4284,N_4143,N_4248);
and U4285 (N_4285,N_4224,N_4246);
nor U4286 (N_4286,N_4217,N_4245);
nand U4287 (N_4287,N_4242,N_4147);
xor U4288 (N_4288,N_4213,N_4247);
xnor U4289 (N_4289,N_4170,N_4228);
nor U4290 (N_4290,N_4160,N_4136);
nand U4291 (N_4291,N_4197,N_4159);
nand U4292 (N_4292,N_4189,N_4138);
or U4293 (N_4293,N_4146,N_4199);
and U4294 (N_4294,N_4198,N_4154);
nand U4295 (N_4295,N_4156,N_4167);
and U4296 (N_4296,N_4211,N_4162);
xor U4297 (N_4297,N_4133,N_4239);
and U4298 (N_4298,N_4177,N_4184);
nor U4299 (N_4299,N_4231,N_4212);
nor U4300 (N_4300,N_4236,N_4201);
nor U4301 (N_4301,N_4214,N_4222);
nor U4302 (N_4302,N_4169,N_4240);
or U4303 (N_4303,N_4179,N_4137);
xnor U4304 (N_4304,N_4204,N_4249);
or U4305 (N_4305,N_4131,N_4152);
xor U4306 (N_4306,N_4190,N_4232);
or U4307 (N_4307,N_4193,N_4139);
and U4308 (N_4308,N_4155,N_4221);
or U4309 (N_4309,N_4234,N_4200);
nor U4310 (N_4310,N_4150,N_4229);
nand U4311 (N_4311,N_4223,N_4134);
nor U4312 (N_4312,N_4153,N_4221);
and U4313 (N_4313,N_4130,N_4195);
xnor U4314 (N_4314,N_4242,N_4161);
and U4315 (N_4315,N_4193,N_4155);
or U4316 (N_4316,N_4172,N_4247);
or U4317 (N_4317,N_4238,N_4146);
or U4318 (N_4318,N_4171,N_4149);
xnor U4319 (N_4319,N_4167,N_4132);
nor U4320 (N_4320,N_4234,N_4137);
nor U4321 (N_4321,N_4138,N_4140);
nand U4322 (N_4322,N_4206,N_4209);
or U4323 (N_4323,N_4138,N_4148);
and U4324 (N_4324,N_4184,N_4148);
nor U4325 (N_4325,N_4211,N_4234);
nand U4326 (N_4326,N_4153,N_4207);
or U4327 (N_4327,N_4204,N_4230);
or U4328 (N_4328,N_4184,N_4225);
or U4329 (N_4329,N_4225,N_4218);
or U4330 (N_4330,N_4181,N_4225);
nor U4331 (N_4331,N_4197,N_4238);
nor U4332 (N_4332,N_4137,N_4187);
nand U4333 (N_4333,N_4234,N_4218);
and U4334 (N_4334,N_4209,N_4179);
or U4335 (N_4335,N_4177,N_4219);
xnor U4336 (N_4336,N_4191,N_4153);
and U4337 (N_4337,N_4186,N_4223);
or U4338 (N_4338,N_4140,N_4196);
xnor U4339 (N_4339,N_4148,N_4226);
xor U4340 (N_4340,N_4191,N_4151);
nor U4341 (N_4341,N_4135,N_4221);
and U4342 (N_4342,N_4181,N_4142);
nand U4343 (N_4343,N_4129,N_4220);
nor U4344 (N_4344,N_4132,N_4218);
or U4345 (N_4345,N_4214,N_4154);
nor U4346 (N_4346,N_4189,N_4246);
and U4347 (N_4347,N_4174,N_4155);
nand U4348 (N_4348,N_4237,N_4207);
and U4349 (N_4349,N_4130,N_4220);
and U4350 (N_4350,N_4240,N_4167);
nand U4351 (N_4351,N_4236,N_4248);
nor U4352 (N_4352,N_4224,N_4210);
nor U4353 (N_4353,N_4241,N_4151);
and U4354 (N_4354,N_4147,N_4165);
or U4355 (N_4355,N_4134,N_4184);
and U4356 (N_4356,N_4125,N_4238);
nor U4357 (N_4357,N_4127,N_4210);
nor U4358 (N_4358,N_4205,N_4159);
nand U4359 (N_4359,N_4221,N_4165);
or U4360 (N_4360,N_4179,N_4139);
nor U4361 (N_4361,N_4132,N_4235);
xor U4362 (N_4362,N_4201,N_4241);
xor U4363 (N_4363,N_4233,N_4215);
or U4364 (N_4364,N_4223,N_4245);
nor U4365 (N_4365,N_4156,N_4141);
or U4366 (N_4366,N_4129,N_4235);
or U4367 (N_4367,N_4147,N_4181);
and U4368 (N_4368,N_4178,N_4220);
xnor U4369 (N_4369,N_4182,N_4135);
xor U4370 (N_4370,N_4234,N_4191);
and U4371 (N_4371,N_4138,N_4248);
nand U4372 (N_4372,N_4152,N_4186);
xnor U4373 (N_4373,N_4245,N_4249);
and U4374 (N_4374,N_4142,N_4163);
nand U4375 (N_4375,N_4283,N_4346);
or U4376 (N_4376,N_4332,N_4269);
xor U4377 (N_4377,N_4339,N_4287);
nand U4378 (N_4378,N_4360,N_4281);
nand U4379 (N_4379,N_4306,N_4337);
and U4380 (N_4380,N_4359,N_4267);
nand U4381 (N_4381,N_4295,N_4369);
or U4382 (N_4382,N_4373,N_4338);
xor U4383 (N_4383,N_4284,N_4351);
nand U4384 (N_4384,N_4307,N_4303);
nand U4385 (N_4385,N_4263,N_4370);
nand U4386 (N_4386,N_4341,N_4314);
nor U4387 (N_4387,N_4288,N_4368);
xor U4388 (N_4388,N_4273,N_4353);
nand U4389 (N_4389,N_4251,N_4312);
or U4390 (N_4390,N_4255,N_4323);
or U4391 (N_4391,N_4271,N_4278);
nand U4392 (N_4392,N_4342,N_4347);
xnor U4393 (N_4393,N_4321,N_4334);
nand U4394 (N_4394,N_4358,N_4279);
and U4395 (N_4395,N_4266,N_4354);
nor U4396 (N_4396,N_4309,N_4292);
xor U4397 (N_4397,N_4363,N_4280);
nand U4398 (N_4398,N_4374,N_4301);
or U4399 (N_4399,N_4275,N_4258);
xnor U4400 (N_4400,N_4305,N_4331);
or U4401 (N_4401,N_4298,N_4274);
and U4402 (N_4402,N_4286,N_4344);
nand U4403 (N_4403,N_4343,N_4311);
and U4404 (N_4404,N_4316,N_4264);
nand U4405 (N_4405,N_4329,N_4367);
and U4406 (N_4406,N_4362,N_4262);
or U4407 (N_4407,N_4261,N_4348);
and U4408 (N_4408,N_4313,N_4304);
xnor U4409 (N_4409,N_4361,N_4350);
or U4410 (N_4410,N_4296,N_4308);
or U4411 (N_4411,N_4325,N_4330);
nor U4412 (N_4412,N_4340,N_4366);
or U4413 (N_4413,N_4320,N_4282);
nand U4414 (N_4414,N_4268,N_4357);
and U4415 (N_4415,N_4291,N_4328);
or U4416 (N_4416,N_4276,N_4277);
xnor U4417 (N_4417,N_4345,N_4315);
and U4418 (N_4418,N_4364,N_4336);
nand U4419 (N_4419,N_4293,N_4257);
and U4420 (N_4420,N_4352,N_4371);
nor U4421 (N_4421,N_4327,N_4302);
and U4422 (N_4422,N_4285,N_4270);
nor U4423 (N_4423,N_4365,N_4318);
nor U4424 (N_4424,N_4319,N_4256);
and U4425 (N_4425,N_4290,N_4254);
xnor U4426 (N_4426,N_4356,N_4259);
or U4427 (N_4427,N_4349,N_4310);
xor U4428 (N_4428,N_4294,N_4297);
and U4429 (N_4429,N_4289,N_4300);
xor U4430 (N_4430,N_4250,N_4299);
nor U4431 (N_4431,N_4252,N_4326);
xnor U4432 (N_4432,N_4322,N_4253);
nand U4433 (N_4433,N_4260,N_4335);
xor U4434 (N_4434,N_4265,N_4372);
nor U4435 (N_4435,N_4355,N_4272);
or U4436 (N_4436,N_4333,N_4317);
and U4437 (N_4437,N_4324,N_4297);
nor U4438 (N_4438,N_4294,N_4371);
xnor U4439 (N_4439,N_4362,N_4279);
nand U4440 (N_4440,N_4299,N_4313);
xor U4441 (N_4441,N_4296,N_4365);
nand U4442 (N_4442,N_4332,N_4280);
nand U4443 (N_4443,N_4268,N_4279);
nor U4444 (N_4444,N_4360,N_4267);
nor U4445 (N_4445,N_4304,N_4262);
and U4446 (N_4446,N_4343,N_4278);
xor U4447 (N_4447,N_4292,N_4341);
nor U4448 (N_4448,N_4287,N_4337);
nor U4449 (N_4449,N_4308,N_4320);
xor U4450 (N_4450,N_4259,N_4371);
xnor U4451 (N_4451,N_4265,N_4254);
and U4452 (N_4452,N_4334,N_4276);
or U4453 (N_4453,N_4362,N_4319);
or U4454 (N_4454,N_4337,N_4281);
nor U4455 (N_4455,N_4287,N_4350);
or U4456 (N_4456,N_4321,N_4269);
nor U4457 (N_4457,N_4353,N_4352);
xor U4458 (N_4458,N_4307,N_4254);
or U4459 (N_4459,N_4263,N_4303);
nor U4460 (N_4460,N_4268,N_4371);
nor U4461 (N_4461,N_4309,N_4287);
nor U4462 (N_4462,N_4292,N_4358);
xnor U4463 (N_4463,N_4284,N_4340);
nor U4464 (N_4464,N_4360,N_4279);
nor U4465 (N_4465,N_4305,N_4366);
xnor U4466 (N_4466,N_4278,N_4311);
nand U4467 (N_4467,N_4373,N_4323);
nand U4468 (N_4468,N_4291,N_4360);
or U4469 (N_4469,N_4285,N_4364);
xor U4470 (N_4470,N_4363,N_4344);
or U4471 (N_4471,N_4270,N_4373);
xnor U4472 (N_4472,N_4342,N_4369);
or U4473 (N_4473,N_4342,N_4253);
nand U4474 (N_4474,N_4276,N_4331);
nor U4475 (N_4475,N_4255,N_4254);
nor U4476 (N_4476,N_4308,N_4356);
and U4477 (N_4477,N_4253,N_4339);
nor U4478 (N_4478,N_4366,N_4373);
nor U4479 (N_4479,N_4350,N_4306);
or U4480 (N_4480,N_4340,N_4297);
xor U4481 (N_4481,N_4282,N_4333);
nand U4482 (N_4482,N_4354,N_4299);
xnor U4483 (N_4483,N_4341,N_4361);
or U4484 (N_4484,N_4270,N_4268);
and U4485 (N_4485,N_4250,N_4300);
nand U4486 (N_4486,N_4350,N_4290);
or U4487 (N_4487,N_4350,N_4332);
xnor U4488 (N_4488,N_4345,N_4310);
or U4489 (N_4489,N_4304,N_4357);
xnor U4490 (N_4490,N_4355,N_4297);
or U4491 (N_4491,N_4288,N_4296);
xor U4492 (N_4492,N_4299,N_4367);
xnor U4493 (N_4493,N_4273,N_4292);
or U4494 (N_4494,N_4332,N_4301);
nand U4495 (N_4495,N_4260,N_4290);
or U4496 (N_4496,N_4270,N_4348);
nor U4497 (N_4497,N_4328,N_4333);
nor U4498 (N_4498,N_4334,N_4280);
xor U4499 (N_4499,N_4345,N_4333);
nand U4500 (N_4500,N_4499,N_4421);
or U4501 (N_4501,N_4418,N_4412);
nor U4502 (N_4502,N_4419,N_4416);
and U4503 (N_4503,N_4485,N_4380);
xor U4504 (N_4504,N_4422,N_4417);
and U4505 (N_4505,N_4453,N_4435);
nor U4506 (N_4506,N_4486,N_4441);
or U4507 (N_4507,N_4444,N_4414);
xor U4508 (N_4508,N_4405,N_4382);
nand U4509 (N_4509,N_4388,N_4452);
nor U4510 (N_4510,N_4477,N_4396);
xor U4511 (N_4511,N_4428,N_4451);
and U4512 (N_4512,N_4464,N_4469);
nand U4513 (N_4513,N_4415,N_4454);
or U4514 (N_4514,N_4439,N_4401);
nand U4515 (N_4515,N_4407,N_4455);
nor U4516 (N_4516,N_4438,N_4430);
xor U4517 (N_4517,N_4381,N_4434);
or U4518 (N_4518,N_4449,N_4402);
or U4519 (N_4519,N_4375,N_4465);
nor U4520 (N_4520,N_4457,N_4466);
nor U4521 (N_4521,N_4397,N_4400);
xor U4522 (N_4522,N_4424,N_4493);
or U4523 (N_4523,N_4394,N_4403);
and U4524 (N_4524,N_4391,N_4461);
xor U4525 (N_4525,N_4495,N_4488);
or U4526 (N_4526,N_4420,N_4497);
nor U4527 (N_4527,N_4459,N_4487);
or U4528 (N_4528,N_4409,N_4474);
and U4529 (N_4529,N_4462,N_4491);
and U4530 (N_4530,N_4468,N_4489);
nor U4531 (N_4531,N_4390,N_4478);
and U4532 (N_4532,N_4450,N_4445);
nor U4533 (N_4533,N_4483,N_4399);
nor U4534 (N_4534,N_4404,N_4426);
xnor U4535 (N_4535,N_4432,N_4446);
nand U4536 (N_4536,N_4392,N_4482);
and U4537 (N_4537,N_4378,N_4431);
nand U4538 (N_4538,N_4494,N_4429);
or U4539 (N_4539,N_4475,N_4467);
nor U4540 (N_4540,N_4470,N_4498);
or U4541 (N_4541,N_4410,N_4490);
xor U4542 (N_4542,N_4377,N_4387);
nor U4543 (N_4543,N_4379,N_4386);
nor U4544 (N_4544,N_4437,N_4398);
and U4545 (N_4545,N_4383,N_4458);
or U4546 (N_4546,N_4460,N_4476);
or U4547 (N_4547,N_4479,N_4376);
nand U4548 (N_4548,N_4440,N_4472);
or U4549 (N_4549,N_4408,N_4427);
and U4550 (N_4550,N_4456,N_4473);
or U4551 (N_4551,N_4496,N_4425);
nand U4552 (N_4552,N_4492,N_4463);
xnor U4553 (N_4553,N_4448,N_4423);
and U4554 (N_4554,N_4411,N_4436);
nor U4555 (N_4555,N_4406,N_4389);
nand U4556 (N_4556,N_4447,N_4443);
nand U4557 (N_4557,N_4433,N_4413);
xor U4558 (N_4558,N_4442,N_4385);
nor U4559 (N_4559,N_4384,N_4393);
nor U4560 (N_4560,N_4471,N_4484);
or U4561 (N_4561,N_4480,N_4395);
xnor U4562 (N_4562,N_4481,N_4485);
nand U4563 (N_4563,N_4459,N_4379);
or U4564 (N_4564,N_4405,N_4497);
xnor U4565 (N_4565,N_4481,N_4429);
and U4566 (N_4566,N_4430,N_4449);
nor U4567 (N_4567,N_4480,N_4460);
xnor U4568 (N_4568,N_4492,N_4404);
nand U4569 (N_4569,N_4421,N_4375);
nand U4570 (N_4570,N_4392,N_4441);
and U4571 (N_4571,N_4499,N_4397);
xnor U4572 (N_4572,N_4375,N_4473);
nand U4573 (N_4573,N_4402,N_4383);
nand U4574 (N_4574,N_4496,N_4422);
nor U4575 (N_4575,N_4472,N_4416);
and U4576 (N_4576,N_4487,N_4384);
nand U4577 (N_4577,N_4426,N_4470);
xor U4578 (N_4578,N_4396,N_4487);
and U4579 (N_4579,N_4430,N_4421);
nand U4580 (N_4580,N_4479,N_4486);
nor U4581 (N_4581,N_4469,N_4492);
nor U4582 (N_4582,N_4391,N_4453);
nand U4583 (N_4583,N_4448,N_4380);
nand U4584 (N_4584,N_4431,N_4466);
and U4585 (N_4585,N_4481,N_4375);
or U4586 (N_4586,N_4379,N_4475);
or U4587 (N_4587,N_4459,N_4396);
nand U4588 (N_4588,N_4382,N_4468);
nand U4589 (N_4589,N_4453,N_4387);
and U4590 (N_4590,N_4435,N_4467);
or U4591 (N_4591,N_4383,N_4389);
nand U4592 (N_4592,N_4409,N_4378);
nand U4593 (N_4593,N_4384,N_4396);
nor U4594 (N_4594,N_4422,N_4457);
nor U4595 (N_4595,N_4470,N_4480);
nor U4596 (N_4596,N_4382,N_4426);
or U4597 (N_4597,N_4395,N_4396);
xnor U4598 (N_4598,N_4420,N_4454);
nand U4599 (N_4599,N_4421,N_4476);
xnor U4600 (N_4600,N_4426,N_4400);
nand U4601 (N_4601,N_4422,N_4493);
or U4602 (N_4602,N_4453,N_4446);
nor U4603 (N_4603,N_4485,N_4401);
xnor U4604 (N_4604,N_4448,N_4387);
xnor U4605 (N_4605,N_4446,N_4381);
and U4606 (N_4606,N_4479,N_4493);
or U4607 (N_4607,N_4395,N_4415);
nor U4608 (N_4608,N_4471,N_4384);
or U4609 (N_4609,N_4446,N_4413);
or U4610 (N_4610,N_4377,N_4376);
xnor U4611 (N_4611,N_4420,N_4482);
xnor U4612 (N_4612,N_4424,N_4405);
or U4613 (N_4613,N_4477,N_4408);
nand U4614 (N_4614,N_4403,N_4409);
nor U4615 (N_4615,N_4485,N_4479);
nor U4616 (N_4616,N_4407,N_4477);
and U4617 (N_4617,N_4473,N_4381);
nand U4618 (N_4618,N_4453,N_4431);
nand U4619 (N_4619,N_4391,N_4450);
xnor U4620 (N_4620,N_4469,N_4410);
nand U4621 (N_4621,N_4422,N_4395);
nor U4622 (N_4622,N_4387,N_4437);
nor U4623 (N_4623,N_4396,N_4423);
nor U4624 (N_4624,N_4432,N_4495);
xnor U4625 (N_4625,N_4551,N_4587);
xnor U4626 (N_4626,N_4594,N_4604);
nand U4627 (N_4627,N_4568,N_4612);
nand U4628 (N_4628,N_4523,N_4585);
nor U4629 (N_4629,N_4580,N_4577);
xor U4630 (N_4630,N_4552,N_4592);
and U4631 (N_4631,N_4615,N_4623);
nor U4632 (N_4632,N_4617,N_4547);
nand U4633 (N_4633,N_4569,N_4528);
or U4634 (N_4634,N_4504,N_4567);
or U4635 (N_4635,N_4514,N_4555);
or U4636 (N_4636,N_4583,N_4517);
nand U4637 (N_4637,N_4564,N_4513);
xnor U4638 (N_4638,N_4500,N_4520);
nor U4639 (N_4639,N_4549,N_4571);
xnor U4640 (N_4640,N_4598,N_4545);
xnor U4641 (N_4641,N_4595,N_4565);
and U4642 (N_4642,N_4588,N_4526);
xor U4643 (N_4643,N_4573,N_4611);
or U4644 (N_4644,N_4518,N_4525);
nor U4645 (N_4645,N_4559,N_4579);
or U4646 (N_4646,N_4596,N_4516);
nand U4647 (N_4647,N_4554,N_4581);
xnor U4648 (N_4648,N_4521,N_4561);
and U4649 (N_4649,N_4553,N_4622);
and U4650 (N_4650,N_4540,N_4616);
xnor U4651 (N_4651,N_4619,N_4572);
nor U4652 (N_4652,N_4614,N_4519);
nand U4653 (N_4653,N_4597,N_4546);
or U4654 (N_4654,N_4515,N_4531);
or U4655 (N_4655,N_4624,N_4591);
nand U4656 (N_4656,N_4590,N_4505);
and U4657 (N_4657,N_4532,N_4541);
and U4658 (N_4658,N_4562,N_4503);
and U4659 (N_4659,N_4509,N_4511);
xor U4660 (N_4660,N_4602,N_4610);
and U4661 (N_4661,N_4584,N_4535);
nor U4662 (N_4662,N_4548,N_4536);
nor U4663 (N_4663,N_4578,N_4539);
or U4664 (N_4664,N_4601,N_4543);
nor U4665 (N_4665,N_4538,N_4533);
and U4666 (N_4666,N_4558,N_4556);
xnor U4667 (N_4667,N_4608,N_4512);
or U4668 (N_4668,N_4586,N_4560);
nor U4669 (N_4669,N_4607,N_4605);
xnor U4670 (N_4670,N_4507,N_4534);
nand U4671 (N_4671,N_4527,N_4576);
or U4672 (N_4672,N_4599,N_4501);
nor U4673 (N_4673,N_4537,N_4570);
or U4674 (N_4674,N_4524,N_4557);
xnor U4675 (N_4675,N_4574,N_4510);
and U4676 (N_4676,N_4621,N_4508);
or U4677 (N_4677,N_4575,N_4542);
xor U4678 (N_4678,N_4613,N_4618);
nor U4679 (N_4679,N_4593,N_4502);
xnor U4680 (N_4680,N_4589,N_4529);
or U4681 (N_4681,N_4606,N_4522);
nand U4682 (N_4682,N_4600,N_4566);
xor U4683 (N_4683,N_4563,N_4603);
and U4684 (N_4684,N_4506,N_4582);
nand U4685 (N_4685,N_4544,N_4609);
xor U4686 (N_4686,N_4620,N_4550);
xnor U4687 (N_4687,N_4530,N_4513);
and U4688 (N_4688,N_4547,N_4507);
xnor U4689 (N_4689,N_4573,N_4600);
nand U4690 (N_4690,N_4602,N_4612);
nor U4691 (N_4691,N_4600,N_4570);
and U4692 (N_4692,N_4529,N_4520);
or U4693 (N_4693,N_4534,N_4529);
nor U4694 (N_4694,N_4612,N_4621);
nand U4695 (N_4695,N_4594,N_4555);
and U4696 (N_4696,N_4618,N_4578);
or U4697 (N_4697,N_4568,N_4563);
or U4698 (N_4698,N_4502,N_4563);
nand U4699 (N_4699,N_4519,N_4605);
nand U4700 (N_4700,N_4514,N_4550);
and U4701 (N_4701,N_4513,N_4572);
nor U4702 (N_4702,N_4563,N_4600);
nor U4703 (N_4703,N_4575,N_4576);
and U4704 (N_4704,N_4545,N_4608);
nand U4705 (N_4705,N_4507,N_4623);
or U4706 (N_4706,N_4500,N_4613);
nand U4707 (N_4707,N_4500,N_4596);
nor U4708 (N_4708,N_4586,N_4543);
nor U4709 (N_4709,N_4555,N_4550);
nor U4710 (N_4710,N_4606,N_4502);
nand U4711 (N_4711,N_4543,N_4518);
nand U4712 (N_4712,N_4533,N_4501);
and U4713 (N_4713,N_4599,N_4542);
or U4714 (N_4714,N_4613,N_4507);
xor U4715 (N_4715,N_4557,N_4535);
xor U4716 (N_4716,N_4532,N_4611);
and U4717 (N_4717,N_4550,N_4529);
xnor U4718 (N_4718,N_4504,N_4547);
nor U4719 (N_4719,N_4572,N_4511);
and U4720 (N_4720,N_4548,N_4554);
xnor U4721 (N_4721,N_4593,N_4567);
xnor U4722 (N_4722,N_4581,N_4524);
xnor U4723 (N_4723,N_4601,N_4555);
xnor U4724 (N_4724,N_4569,N_4570);
xnor U4725 (N_4725,N_4622,N_4527);
nor U4726 (N_4726,N_4511,N_4584);
nand U4727 (N_4727,N_4588,N_4617);
and U4728 (N_4728,N_4573,N_4538);
and U4729 (N_4729,N_4576,N_4548);
or U4730 (N_4730,N_4591,N_4533);
and U4731 (N_4731,N_4564,N_4574);
nor U4732 (N_4732,N_4541,N_4548);
nor U4733 (N_4733,N_4595,N_4594);
and U4734 (N_4734,N_4567,N_4502);
or U4735 (N_4735,N_4548,N_4561);
xnor U4736 (N_4736,N_4623,N_4558);
nor U4737 (N_4737,N_4500,N_4580);
xnor U4738 (N_4738,N_4611,N_4555);
xor U4739 (N_4739,N_4556,N_4537);
or U4740 (N_4740,N_4502,N_4508);
nand U4741 (N_4741,N_4593,N_4574);
nor U4742 (N_4742,N_4569,N_4609);
nor U4743 (N_4743,N_4606,N_4542);
nand U4744 (N_4744,N_4605,N_4586);
and U4745 (N_4745,N_4582,N_4510);
and U4746 (N_4746,N_4577,N_4523);
nand U4747 (N_4747,N_4610,N_4622);
and U4748 (N_4748,N_4531,N_4557);
or U4749 (N_4749,N_4544,N_4566);
nand U4750 (N_4750,N_4691,N_4634);
and U4751 (N_4751,N_4745,N_4671);
xor U4752 (N_4752,N_4736,N_4660);
or U4753 (N_4753,N_4677,N_4697);
nand U4754 (N_4754,N_4642,N_4692);
nand U4755 (N_4755,N_4662,N_4629);
or U4756 (N_4756,N_4733,N_4718);
xor U4757 (N_4757,N_4647,N_4650);
nor U4758 (N_4758,N_4705,N_4641);
and U4759 (N_4759,N_4659,N_4701);
or U4760 (N_4760,N_4675,N_4749);
nand U4761 (N_4761,N_4698,N_4648);
and U4762 (N_4762,N_4730,N_4737);
xnor U4763 (N_4763,N_4638,N_4681);
and U4764 (N_4764,N_4672,N_4635);
nand U4765 (N_4765,N_4680,N_4683);
and U4766 (N_4766,N_4741,N_4711);
or U4767 (N_4767,N_4673,N_4731);
or U4768 (N_4768,N_4664,N_4747);
nand U4769 (N_4769,N_4655,N_4684);
xor U4770 (N_4770,N_4654,N_4667);
nor U4771 (N_4771,N_4669,N_4685);
nor U4772 (N_4772,N_4627,N_4740);
nor U4773 (N_4773,N_4657,N_4636);
and U4774 (N_4774,N_4693,N_4632);
nand U4775 (N_4775,N_4744,N_4716);
and U4776 (N_4776,N_4727,N_4656);
nand U4777 (N_4777,N_4703,N_4728);
and U4778 (N_4778,N_4742,N_4732);
xor U4779 (N_4779,N_4652,N_4707);
nor U4780 (N_4780,N_4689,N_4708);
nand U4781 (N_4781,N_4658,N_4688);
nor U4782 (N_4782,N_4670,N_4640);
or U4783 (N_4783,N_4713,N_4700);
nand U4784 (N_4784,N_4738,N_4726);
nand U4785 (N_4785,N_4729,N_4663);
or U4786 (N_4786,N_4706,N_4714);
nand U4787 (N_4787,N_4702,N_4651);
and U4788 (N_4788,N_4628,N_4739);
and U4789 (N_4789,N_4710,N_4719);
xnor U4790 (N_4790,N_4717,N_4653);
nand U4791 (N_4791,N_4746,N_4676);
xor U4792 (N_4792,N_4645,N_4625);
or U4793 (N_4793,N_4626,N_4687);
nor U4794 (N_4794,N_4722,N_4643);
and U4795 (N_4795,N_4720,N_4725);
nand U4796 (N_4796,N_4712,N_4735);
nor U4797 (N_4797,N_4724,N_4633);
nor U4798 (N_4798,N_4630,N_4679);
nand U4799 (N_4799,N_4649,N_4678);
and U4800 (N_4800,N_4690,N_4695);
and U4801 (N_4801,N_4668,N_4743);
nand U4802 (N_4802,N_4637,N_4661);
nor U4803 (N_4803,N_4631,N_4694);
xor U4804 (N_4804,N_4715,N_4686);
or U4805 (N_4805,N_4644,N_4665);
xor U4806 (N_4806,N_4723,N_4666);
nor U4807 (N_4807,N_4709,N_4704);
and U4808 (N_4808,N_4699,N_4674);
and U4809 (N_4809,N_4721,N_4682);
and U4810 (N_4810,N_4696,N_4734);
xor U4811 (N_4811,N_4646,N_4639);
nor U4812 (N_4812,N_4748,N_4717);
nand U4813 (N_4813,N_4747,N_4668);
or U4814 (N_4814,N_4638,N_4736);
and U4815 (N_4815,N_4700,N_4652);
and U4816 (N_4816,N_4733,N_4749);
nand U4817 (N_4817,N_4653,N_4729);
nand U4818 (N_4818,N_4683,N_4713);
or U4819 (N_4819,N_4740,N_4730);
or U4820 (N_4820,N_4670,N_4709);
and U4821 (N_4821,N_4704,N_4725);
or U4822 (N_4822,N_4677,N_4684);
and U4823 (N_4823,N_4690,N_4646);
nand U4824 (N_4824,N_4721,N_4663);
nor U4825 (N_4825,N_4673,N_4700);
or U4826 (N_4826,N_4714,N_4721);
or U4827 (N_4827,N_4680,N_4638);
nand U4828 (N_4828,N_4712,N_4723);
or U4829 (N_4829,N_4734,N_4738);
or U4830 (N_4830,N_4693,N_4686);
nand U4831 (N_4831,N_4717,N_4652);
nor U4832 (N_4832,N_4749,N_4732);
and U4833 (N_4833,N_4725,N_4688);
and U4834 (N_4834,N_4641,N_4733);
or U4835 (N_4835,N_4742,N_4667);
and U4836 (N_4836,N_4635,N_4696);
xnor U4837 (N_4837,N_4634,N_4682);
and U4838 (N_4838,N_4682,N_4700);
or U4839 (N_4839,N_4668,N_4695);
nor U4840 (N_4840,N_4632,N_4725);
xnor U4841 (N_4841,N_4639,N_4737);
or U4842 (N_4842,N_4708,N_4634);
nand U4843 (N_4843,N_4712,N_4698);
nand U4844 (N_4844,N_4708,N_4676);
nand U4845 (N_4845,N_4660,N_4681);
xnor U4846 (N_4846,N_4694,N_4740);
nor U4847 (N_4847,N_4726,N_4668);
and U4848 (N_4848,N_4729,N_4655);
and U4849 (N_4849,N_4714,N_4697);
xor U4850 (N_4850,N_4704,N_4717);
nand U4851 (N_4851,N_4631,N_4716);
and U4852 (N_4852,N_4690,N_4729);
xor U4853 (N_4853,N_4720,N_4689);
nor U4854 (N_4854,N_4713,N_4720);
or U4855 (N_4855,N_4701,N_4710);
and U4856 (N_4856,N_4665,N_4735);
nand U4857 (N_4857,N_4709,N_4705);
nand U4858 (N_4858,N_4736,N_4637);
xnor U4859 (N_4859,N_4687,N_4644);
and U4860 (N_4860,N_4708,N_4652);
and U4861 (N_4861,N_4642,N_4733);
xor U4862 (N_4862,N_4738,N_4664);
or U4863 (N_4863,N_4663,N_4648);
xnor U4864 (N_4864,N_4645,N_4673);
nor U4865 (N_4865,N_4702,N_4682);
nor U4866 (N_4866,N_4735,N_4722);
nor U4867 (N_4867,N_4650,N_4644);
or U4868 (N_4868,N_4628,N_4705);
or U4869 (N_4869,N_4710,N_4627);
or U4870 (N_4870,N_4675,N_4659);
or U4871 (N_4871,N_4699,N_4722);
or U4872 (N_4872,N_4682,N_4638);
nor U4873 (N_4873,N_4731,N_4629);
nor U4874 (N_4874,N_4709,N_4679);
nor U4875 (N_4875,N_4774,N_4851);
xor U4876 (N_4876,N_4825,N_4872);
nor U4877 (N_4877,N_4780,N_4782);
and U4878 (N_4878,N_4795,N_4755);
nand U4879 (N_4879,N_4813,N_4778);
or U4880 (N_4880,N_4751,N_4758);
nand U4881 (N_4881,N_4840,N_4800);
and U4882 (N_4882,N_4806,N_4862);
xnor U4883 (N_4883,N_4819,N_4803);
nor U4884 (N_4884,N_4759,N_4841);
or U4885 (N_4885,N_4839,N_4761);
xor U4886 (N_4886,N_4866,N_4850);
or U4887 (N_4887,N_4865,N_4811);
and U4888 (N_4888,N_4873,N_4855);
xnor U4889 (N_4889,N_4821,N_4805);
nand U4890 (N_4890,N_4833,N_4820);
xor U4891 (N_4891,N_4854,N_4786);
nand U4892 (N_4892,N_4763,N_4760);
or U4893 (N_4893,N_4775,N_4858);
nand U4894 (N_4894,N_4766,N_4861);
and U4895 (N_4895,N_4767,N_4859);
xnor U4896 (N_4896,N_4797,N_4871);
nand U4897 (N_4897,N_4785,N_4874);
nor U4898 (N_4898,N_4799,N_4753);
nand U4899 (N_4899,N_4818,N_4779);
xnor U4900 (N_4900,N_4777,N_4822);
nor U4901 (N_4901,N_4792,N_4781);
and U4902 (N_4902,N_4809,N_4828);
xnor U4903 (N_4903,N_4768,N_4824);
and U4904 (N_4904,N_4867,N_4817);
or U4905 (N_4905,N_4816,N_4765);
nand U4906 (N_4906,N_4752,N_4804);
and U4907 (N_4907,N_4791,N_4847);
nand U4908 (N_4908,N_4807,N_4832);
nor U4909 (N_4909,N_4798,N_4794);
nand U4910 (N_4910,N_4756,N_4848);
nor U4911 (N_4911,N_4864,N_4790);
nor U4912 (N_4912,N_4796,N_4757);
nand U4913 (N_4913,N_4764,N_4773);
and U4914 (N_4914,N_4829,N_4801);
xnor U4915 (N_4915,N_4869,N_4769);
nor U4916 (N_4916,N_4835,N_4783);
or U4917 (N_4917,N_4750,N_4772);
or U4918 (N_4918,N_4868,N_4771);
xnor U4919 (N_4919,N_4836,N_4843);
xor U4920 (N_4920,N_4837,N_4793);
and U4921 (N_4921,N_4838,N_4844);
or U4922 (N_4922,N_4754,N_4815);
nor U4923 (N_4923,N_4857,N_4852);
nand U4924 (N_4924,N_4812,N_4856);
xor U4925 (N_4925,N_4789,N_4810);
and U4926 (N_4926,N_4784,N_4842);
or U4927 (N_4927,N_4762,N_4860);
xnor U4928 (N_4928,N_4770,N_4802);
xor U4929 (N_4929,N_4831,N_4788);
nand U4930 (N_4930,N_4826,N_4814);
nor U4931 (N_4931,N_4827,N_4853);
nor U4932 (N_4932,N_4823,N_4776);
nand U4933 (N_4933,N_4870,N_4787);
nand U4934 (N_4934,N_4808,N_4834);
nand U4935 (N_4935,N_4830,N_4849);
xnor U4936 (N_4936,N_4863,N_4846);
or U4937 (N_4937,N_4845,N_4843);
nand U4938 (N_4938,N_4768,N_4834);
or U4939 (N_4939,N_4824,N_4763);
nor U4940 (N_4940,N_4867,N_4856);
nor U4941 (N_4941,N_4766,N_4865);
and U4942 (N_4942,N_4805,N_4766);
nand U4943 (N_4943,N_4835,N_4764);
or U4944 (N_4944,N_4854,N_4859);
xor U4945 (N_4945,N_4826,N_4760);
nand U4946 (N_4946,N_4866,N_4806);
nand U4947 (N_4947,N_4866,N_4858);
nor U4948 (N_4948,N_4789,N_4868);
xnor U4949 (N_4949,N_4756,N_4780);
and U4950 (N_4950,N_4801,N_4788);
xor U4951 (N_4951,N_4811,N_4786);
xor U4952 (N_4952,N_4770,N_4771);
nand U4953 (N_4953,N_4813,N_4851);
nor U4954 (N_4954,N_4776,N_4872);
or U4955 (N_4955,N_4802,N_4762);
nor U4956 (N_4956,N_4853,N_4773);
nand U4957 (N_4957,N_4810,N_4768);
nand U4958 (N_4958,N_4859,N_4803);
or U4959 (N_4959,N_4853,N_4839);
nand U4960 (N_4960,N_4793,N_4809);
or U4961 (N_4961,N_4837,N_4857);
nand U4962 (N_4962,N_4845,N_4818);
nand U4963 (N_4963,N_4874,N_4764);
nand U4964 (N_4964,N_4861,N_4776);
or U4965 (N_4965,N_4766,N_4760);
xor U4966 (N_4966,N_4783,N_4786);
xor U4967 (N_4967,N_4829,N_4820);
or U4968 (N_4968,N_4843,N_4754);
or U4969 (N_4969,N_4856,N_4849);
xor U4970 (N_4970,N_4786,N_4818);
xnor U4971 (N_4971,N_4774,N_4800);
and U4972 (N_4972,N_4867,N_4789);
or U4973 (N_4973,N_4830,N_4833);
xnor U4974 (N_4974,N_4817,N_4828);
or U4975 (N_4975,N_4819,N_4774);
and U4976 (N_4976,N_4796,N_4799);
nand U4977 (N_4977,N_4816,N_4761);
nand U4978 (N_4978,N_4859,N_4773);
xnor U4979 (N_4979,N_4850,N_4817);
xnor U4980 (N_4980,N_4780,N_4830);
nor U4981 (N_4981,N_4818,N_4855);
nor U4982 (N_4982,N_4822,N_4865);
nand U4983 (N_4983,N_4859,N_4796);
and U4984 (N_4984,N_4768,N_4798);
nand U4985 (N_4985,N_4759,N_4760);
xor U4986 (N_4986,N_4858,N_4759);
and U4987 (N_4987,N_4810,N_4840);
xor U4988 (N_4988,N_4851,N_4778);
xor U4989 (N_4989,N_4825,N_4765);
and U4990 (N_4990,N_4852,N_4850);
nand U4991 (N_4991,N_4795,N_4803);
and U4992 (N_4992,N_4775,N_4794);
xor U4993 (N_4993,N_4779,N_4802);
and U4994 (N_4994,N_4873,N_4810);
nor U4995 (N_4995,N_4813,N_4772);
xor U4996 (N_4996,N_4852,N_4846);
xor U4997 (N_4997,N_4797,N_4862);
nand U4998 (N_4998,N_4837,N_4780);
xnor U4999 (N_4999,N_4835,N_4817);
and U5000 (N_5000,N_4988,N_4877);
and U5001 (N_5001,N_4943,N_4974);
nand U5002 (N_5002,N_4977,N_4963);
nand U5003 (N_5003,N_4980,N_4927);
nand U5004 (N_5004,N_4999,N_4917);
xnor U5005 (N_5005,N_4968,N_4948);
and U5006 (N_5006,N_4887,N_4907);
and U5007 (N_5007,N_4909,N_4918);
or U5008 (N_5008,N_4978,N_4990);
and U5009 (N_5009,N_4912,N_4895);
or U5010 (N_5010,N_4890,N_4994);
nand U5011 (N_5011,N_4901,N_4889);
or U5012 (N_5012,N_4965,N_4992);
or U5013 (N_5013,N_4923,N_4906);
nor U5014 (N_5014,N_4921,N_4949);
xnor U5015 (N_5015,N_4944,N_4882);
nand U5016 (N_5016,N_4914,N_4883);
xor U5017 (N_5017,N_4931,N_4956);
or U5018 (N_5018,N_4955,N_4985);
or U5019 (N_5019,N_4934,N_4935);
and U5020 (N_5020,N_4982,N_4892);
nand U5021 (N_5021,N_4998,N_4938);
xnor U5022 (N_5022,N_4881,N_4996);
or U5023 (N_5023,N_4919,N_4973);
nand U5024 (N_5024,N_4908,N_4904);
and U5025 (N_5025,N_4975,N_4941);
nand U5026 (N_5026,N_4928,N_4954);
nand U5027 (N_5027,N_4983,N_4897);
nand U5028 (N_5028,N_4997,N_4959);
or U5029 (N_5029,N_4960,N_4879);
xor U5030 (N_5030,N_4969,N_4979);
xnor U5031 (N_5031,N_4878,N_4971);
and U5032 (N_5032,N_4900,N_4920);
nor U5033 (N_5033,N_4984,N_4940);
or U5034 (N_5034,N_4942,N_4896);
and U5035 (N_5035,N_4905,N_4953);
nand U5036 (N_5036,N_4946,N_4936);
nor U5037 (N_5037,N_4903,N_4924);
nand U5038 (N_5038,N_4958,N_4893);
xnor U5039 (N_5039,N_4894,N_4930);
nand U5040 (N_5040,N_4876,N_4947);
nor U5041 (N_5041,N_4880,N_4964);
xor U5042 (N_5042,N_4966,N_4925);
and U5043 (N_5043,N_4967,N_4898);
nand U5044 (N_5044,N_4995,N_4976);
or U5045 (N_5045,N_4884,N_4939);
nor U5046 (N_5046,N_4957,N_4989);
and U5047 (N_5047,N_4886,N_4970);
nor U5048 (N_5048,N_4932,N_4987);
nor U5049 (N_5049,N_4981,N_4937);
or U5050 (N_5050,N_4916,N_4922);
xnor U5051 (N_5051,N_4888,N_4915);
or U5052 (N_5052,N_4951,N_4945);
and U5053 (N_5053,N_4961,N_4993);
xnor U5054 (N_5054,N_4891,N_4929);
nand U5055 (N_5055,N_4902,N_4885);
and U5056 (N_5056,N_4972,N_4952);
nor U5057 (N_5057,N_4910,N_4899);
and U5058 (N_5058,N_4875,N_4991);
nand U5059 (N_5059,N_4950,N_4926);
nor U5060 (N_5060,N_4933,N_4911);
and U5061 (N_5061,N_4986,N_4962);
nand U5062 (N_5062,N_4913,N_4980);
or U5063 (N_5063,N_4919,N_4910);
nand U5064 (N_5064,N_4973,N_4996);
xnor U5065 (N_5065,N_4878,N_4919);
nor U5066 (N_5066,N_4995,N_4938);
xnor U5067 (N_5067,N_4933,N_4879);
nand U5068 (N_5068,N_4894,N_4987);
nand U5069 (N_5069,N_4919,N_4954);
nor U5070 (N_5070,N_4989,N_4998);
and U5071 (N_5071,N_4892,N_4958);
and U5072 (N_5072,N_4932,N_4942);
and U5073 (N_5073,N_4959,N_4969);
or U5074 (N_5074,N_4961,N_4882);
and U5075 (N_5075,N_4968,N_4979);
nand U5076 (N_5076,N_4967,N_4943);
and U5077 (N_5077,N_4921,N_4945);
or U5078 (N_5078,N_4955,N_4963);
xnor U5079 (N_5079,N_4910,N_4917);
nand U5080 (N_5080,N_4890,N_4900);
or U5081 (N_5081,N_4923,N_4966);
and U5082 (N_5082,N_4977,N_4950);
or U5083 (N_5083,N_4938,N_4985);
nor U5084 (N_5084,N_4962,N_4897);
nor U5085 (N_5085,N_4932,N_4978);
or U5086 (N_5086,N_4958,N_4956);
and U5087 (N_5087,N_4903,N_4894);
and U5088 (N_5088,N_4896,N_4910);
or U5089 (N_5089,N_4927,N_4911);
and U5090 (N_5090,N_4879,N_4942);
or U5091 (N_5091,N_4971,N_4958);
nand U5092 (N_5092,N_4880,N_4919);
nand U5093 (N_5093,N_4976,N_4985);
or U5094 (N_5094,N_4957,N_4906);
nor U5095 (N_5095,N_4942,N_4889);
nand U5096 (N_5096,N_4954,N_4882);
nand U5097 (N_5097,N_4935,N_4888);
or U5098 (N_5098,N_4883,N_4987);
or U5099 (N_5099,N_4890,N_4899);
nand U5100 (N_5100,N_4969,N_4932);
or U5101 (N_5101,N_4922,N_4978);
nand U5102 (N_5102,N_4977,N_4886);
xor U5103 (N_5103,N_4909,N_4912);
xnor U5104 (N_5104,N_4987,N_4881);
xnor U5105 (N_5105,N_4978,N_4942);
nor U5106 (N_5106,N_4895,N_4979);
xor U5107 (N_5107,N_4977,N_4879);
or U5108 (N_5108,N_4997,N_4958);
nor U5109 (N_5109,N_4883,N_4989);
xnor U5110 (N_5110,N_4880,N_4923);
xor U5111 (N_5111,N_4956,N_4892);
or U5112 (N_5112,N_4973,N_4913);
or U5113 (N_5113,N_4911,N_4979);
nor U5114 (N_5114,N_4927,N_4897);
nor U5115 (N_5115,N_4983,N_4966);
or U5116 (N_5116,N_4878,N_4992);
or U5117 (N_5117,N_4967,N_4996);
xnor U5118 (N_5118,N_4931,N_4982);
and U5119 (N_5119,N_4938,N_4933);
xnor U5120 (N_5120,N_4973,N_4957);
nor U5121 (N_5121,N_4940,N_4944);
xnor U5122 (N_5122,N_4942,N_4928);
xor U5123 (N_5123,N_4889,N_4978);
nor U5124 (N_5124,N_4945,N_4905);
and U5125 (N_5125,N_5023,N_5067);
and U5126 (N_5126,N_5088,N_5013);
and U5127 (N_5127,N_5097,N_5071);
and U5128 (N_5128,N_5074,N_5114);
nand U5129 (N_5129,N_5115,N_5066);
nand U5130 (N_5130,N_5031,N_5007);
and U5131 (N_5131,N_5014,N_5054);
and U5132 (N_5132,N_5117,N_5116);
nor U5133 (N_5133,N_5111,N_5049);
xnor U5134 (N_5134,N_5019,N_5038);
xor U5135 (N_5135,N_5072,N_5087);
and U5136 (N_5136,N_5077,N_5080);
xor U5137 (N_5137,N_5010,N_5005);
xor U5138 (N_5138,N_5075,N_5092);
nand U5139 (N_5139,N_5078,N_5002);
nor U5140 (N_5140,N_5095,N_5001);
xor U5141 (N_5141,N_5045,N_5032);
nor U5142 (N_5142,N_5044,N_5119);
or U5143 (N_5143,N_5083,N_5026);
nor U5144 (N_5144,N_5096,N_5086);
xnor U5145 (N_5145,N_5076,N_5039);
xnor U5146 (N_5146,N_5004,N_5106);
or U5147 (N_5147,N_5108,N_5028);
and U5148 (N_5148,N_5048,N_5041);
or U5149 (N_5149,N_5120,N_5124);
or U5150 (N_5150,N_5061,N_5123);
or U5151 (N_5151,N_5091,N_5015);
nor U5152 (N_5152,N_5112,N_5018);
xor U5153 (N_5153,N_5052,N_5105);
nand U5154 (N_5154,N_5000,N_5094);
nand U5155 (N_5155,N_5047,N_5058);
xnor U5156 (N_5156,N_5104,N_5056);
xor U5157 (N_5157,N_5089,N_5034);
and U5158 (N_5158,N_5102,N_5110);
xnor U5159 (N_5159,N_5008,N_5122);
xnor U5160 (N_5160,N_5079,N_5098);
or U5161 (N_5161,N_5073,N_5059);
xor U5162 (N_5162,N_5020,N_5011);
and U5163 (N_5163,N_5006,N_5036);
nand U5164 (N_5164,N_5069,N_5063);
nand U5165 (N_5165,N_5084,N_5021);
xnor U5166 (N_5166,N_5033,N_5012);
or U5167 (N_5167,N_5082,N_5107);
and U5168 (N_5168,N_5027,N_5070);
nand U5169 (N_5169,N_5113,N_5053);
nand U5170 (N_5170,N_5060,N_5093);
and U5171 (N_5171,N_5037,N_5103);
or U5172 (N_5172,N_5009,N_5057);
nand U5173 (N_5173,N_5118,N_5090);
nand U5174 (N_5174,N_5030,N_5046);
and U5175 (N_5175,N_5024,N_5035);
nand U5176 (N_5176,N_5064,N_5042);
and U5177 (N_5177,N_5050,N_5062);
xnor U5178 (N_5178,N_5017,N_5022);
and U5179 (N_5179,N_5043,N_5055);
xnor U5180 (N_5180,N_5081,N_5065);
xnor U5181 (N_5181,N_5016,N_5025);
or U5182 (N_5182,N_5029,N_5003);
nor U5183 (N_5183,N_5068,N_5100);
nor U5184 (N_5184,N_5101,N_5085);
or U5185 (N_5185,N_5051,N_5099);
nand U5186 (N_5186,N_5040,N_5109);
or U5187 (N_5187,N_5121,N_5124);
or U5188 (N_5188,N_5055,N_5024);
or U5189 (N_5189,N_5021,N_5076);
or U5190 (N_5190,N_5120,N_5013);
or U5191 (N_5191,N_5029,N_5067);
and U5192 (N_5192,N_5079,N_5062);
and U5193 (N_5193,N_5037,N_5031);
nand U5194 (N_5194,N_5062,N_5073);
xor U5195 (N_5195,N_5006,N_5035);
or U5196 (N_5196,N_5110,N_5044);
or U5197 (N_5197,N_5068,N_5019);
nor U5198 (N_5198,N_5086,N_5100);
nand U5199 (N_5199,N_5121,N_5067);
nand U5200 (N_5200,N_5058,N_5022);
nand U5201 (N_5201,N_5009,N_5017);
nor U5202 (N_5202,N_5122,N_5067);
nor U5203 (N_5203,N_5010,N_5105);
xor U5204 (N_5204,N_5095,N_5115);
nand U5205 (N_5205,N_5110,N_5121);
nand U5206 (N_5206,N_5068,N_5087);
xor U5207 (N_5207,N_5073,N_5000);
and U5208 (N_5208,N_5117,N_5029);
nor U5209 (N_5209,N_5055,N_5094);
nand U5210 (N_5210,N_5043,N_5019);
and U5211 (N_5211,N_5035,N_5098);
xnor U5212 (N_5212,N_5038,N_5042);
or U5213 (N_5213,N_5017,N_5067);
nand U5214 (N_5214,N_5040,N_5016);
or U5215 (N_5215,N_5037,N_5044);
and U5216 (N_5216,N_5100,N_5124);
and U5217 (N_5217,N_5114,N_5079);
and U5218 (N_5218,N_5092,N_5085);
and U5219 (N_5219,N_5034,N_5063);
or U5220 (N_5220,N_5019,N_5046);
nor U5221 (N_5221,N_5042,N_5035);
or U5222 (N_5222,N_5008,N_5005);
or U5223 (N_5223,N_5008,N_5072);
or U5224 (N_5224,N_5112,N_5119);
nand U5225 (N_5225,N_5056,N_5028);
or U5226 (N_5226,N_5083,N_5013);
nand U5227 (N_5227,N_5083,N_5037);
or U5228 (N_5228,N_5043,N_5057);
and U5229 (N_5229,N_5043,N_5036);
nand U5230 (N_5230,N_5041,N_5082);
nor U5231 (N_5231,N_5087,N_5094);
nor U5232 (N_5232,N_5020,N_5094);
xnor U5233 (N_5233,N_5001,N_5023);
and U5234 (N_5234,N_5115,N_5048);
and U5235 (N_5235,N_5055,N_5015);
nor U5236 (N_5236,N_5071,N_5076);
nand U5237 (N_5237,N_5114,N_5112);
nor U5238 (N_5238,N_5026,N_5052);
xnor U5239 (N_5239,N_5114,N_5118);
xor U5240 (N_5240,N_5002,N_5060);
nand U5241 (N_5241,N_5109,N_5060);
nand U5242 (N_5242,N_5048,N_5067);
xnor U5243 (N_5243,N_5007,N_5038);
nor U5244 (N_5244,N_5044,N_5072);
xor U5245 (N_5245,N_5036,N_5012);
and U5246 (N_5246,N_5074,N_5039);
nor U5247 (N_5247,N_5097,N_5103);
nor U5248 (N_5248,N_5059,N_5046);
nor U5249 (N_5249,N_5111,N_5032);
nand U5250 (N_5250,N_5246,N_5164);
xor U5251 (N_5251,N_5151,N_5226);
and U5252 (N_5252,N_5178,N_5241);
or U5253 (N_5253,N_5239,N_5180);
nand U5254 (N_5254,N_5244,N_5165);
nand U5255 (N_5255,N_5135,N_5140);
xor U5256 (N_5256,N_5249,N_5125);
xnor U5257 (N_5257,N_5170,N_5136);
xor U5258 (N_5258,N_5203,N_5128);
and U5259 (N_5259,N_5227,N_5219);
nor U5260 (N_5260,N_5235,N_5197);
and U5261 (N_5261,N_5234,N_5162);
nand U5262 (N_5262,N_5130,N_5231);
and U5263 (N_5263,N_5242,N_5179);
nor U5264 (N_5264,N_5199,N_5171);
and U5265 (N_5265,N_5218,N_5212);
nor U5266 (N_5266,N_5163,N_5202);
nand U5267 (N_5267,N_5193,N_5190);
nand U5268 (N_5268,N_5154,N_5138);
nand U5269 (N_5269,N_5172,N_5209);
nand U5270 (N_5270,N_5191,N_5177);
and U5271 (N_5271,N_5215,N_5147);
xor U5272 (N_5272,N_5213,N_5194);
and U5273 (N_5273,N_5168,N_5236);
and U5274 (N_5274,N_5158,N_5208);
nor U5275 (N_5275,N_5232,N_5224);
nand U5276 (N_5276,N_5206,N_5181);
nand U5277 (N_5277,N_5211,N_5229);
or U5278 (N_5278,N_5173,N_5167);
xor U5279 (N_5279,N_5148,N_5186);
or U5280 (N_5280,N_5214,N_5131);
nor U5281 (N_5281,N_5225,N_5153);
xnor U5282 (N_5282,N_5223,N_5156);
or U5283 (N_5283,N_5245,N_5169);
or U5284 (N_5284,N_5185,N_5204);
or U5285 (N_5285,N_5238,N_5230);
nand U5286 (N_5286,N_5237,N_5139);
or U5287 (N_5287,N_5221,N_5207);
nand U5288 (N_5288,N_5195,N_5188);
nor U5289 (N_5289,N_5192,N_5141);
and U5290 (N_5290,N_5137,N_5233);
xor U5291 (N_5291,N_5248,N_5142);
and U5292 (N_5292,N_5149,N_5127);
and U5293 (N_5293,N_5200,N_5144);
nand U5294 (N_5294,N_5134,N_5146);
and U5295 (N_5295,N_5176,N_5157);
nor U5296 (N_5296,N_5166,N_5205);
and U5297 (N_5297,N_5220,N_5183);
and U5298 (N_5298,N_5155,N_5198);
or U5299 (N_5299,N_5161,N_5129);
or U5300 (N_5300,N_5243,N_5182);
xnor U5301 (N_5301,N_5160,N_5196);
or U5302 (N_5302,N_5145,N_5132);
and U5303 (N_5303,N_5152,N_5143);
and U5304 (N_5304,N_5216,N_5175);
and U5305 (N_5305,N_5174,N_5133);
or U5306 (N_5306,N_5126,N_5189);
and U5307 (N_5307,N_5184,N_5150);
nor U5308 (N_5308,N_5187,N_5217);
nor U5309 (N_5309,N_5201,N_5247);
or U5310 (N_5310,N_5222,N_5210);
nor U5311 (N_5311,N_5228,N_5240);
nand U5312 (N_5312,N_5159,N_5204);
xor U5313 (N_5313,N_5132,N_5244);
and U5314 (N_5314,N_5190,N_5196);
and U5315 (N_5315,N_5134,N_5197);
and U5316 (N_5316,N_5186,N_5195);
nand U5317 (N_5317,N_5180,N_5189);
nand U5318 (N_5318,N_5180,N_5231);
xor U5319 (N_5319,N_5155,N_5150);
or U5320 (N_5320,N_5138,N_5221);
nand U5321 (N_5321,N_5215,N_5187);
and U5322 (N_5322,N_5219,N_5231);
xnor U5323 (N_5323,N_5173,N_5241);
and U5324 (N_5324,N_5151,N_5197);
nor U5325 (N_5325,N_5230,N_5173);
or U5326 (N_5326,N_5203,N_5153);
xor U5327 (N_5327,N_5236,N_5179);
nor U5328 (N_5328,N_5206,N_5221);
xor U5329 (N_5329,N_5146,N_5159);
nor U5330 (N_5330,N_5249,N_5225);
nor U5331 (N_5331,N_5249,N_5208);
or U5332 (N_5332,N_5212,N_5240);
or U5333 (N_5333,N_5211,N_5129);
xor U5334 (N_5334,N_5190,N_5166);
nand U5335 (N_5335,N_5244,N_5159);
nor U5336 (N_5336,N_5165,N_5166);
or U5337 (N_5337,N_5135,N_5130);
or U5338 (N_5338,N_5233,N_5249);
xor U5339 (N_5339,N_5145,N_5185);
nand U5340 (N_5340,N_5212,N_5135);
or U5341 (N_5341,N_5128,N_5168);
nor U5342 (N_5342,N_5135,N_5174);
nand U5343 (N_5343,N_5242,N_5181);
nor U5344 (N_5344,N_5190,N_5199);
xor U5345 (N_5345,N_5132,N_5233);
or U5346 (N_5346,N_5214,N_5193);
nor U5347 (N_5347,N_5228,N_5157);
and U5348 (N_5348,N_5185,N_5182);
or U5349 (N_5349,N_5190,N_5216);
or U5350 (N_5350,N_5168,N_5249);
nand U5351 (N_5351,N_5203,N_5222);
or U5352 (N_5352,N_5225,N_5184);
or U5353 (N_5353,N_5157,N_5221);
nor U5354 (N_5354,N_5165,N_5140);
or U5355 (N_5355,N_5227,N_5206);
nand U5356 (N_5356,N_5222,N_5221);
xor U5357 (N_5357,N_5247,N_5143);
xor U5358 (N_5358,N_5216,N_5228);
or U5359 (N_5359,N_5138,N_5223);
or U5360 (N_5360,N_5166,N_5242);
or U5361 (N_5361,N_5205,N_5247);
xor U5362 (N_5362,N_5178,N_5195);
nand U5363 (N_5363,N_5230,N_5234);
or U5364 (N_5364,N_5130,N_5189);
nand U5365 (N_5365,N_5185,N_5239);
xor U5366 (N_5366,N_5213,N_5159);
nor U5367 (N_5367,N_5146,N_5238);
nor U5368 (N_5368,N_5133,N_5128);
nor U5369 (N_5369,N_5248,N_5178);
and U5370 (N_5370,N_5248,N_5207);
nor U5371 (N_5371,N_5134,N_5177);
or U5372 (N_5372,N_5239,N_5201);
xnor U5373 (N_5373,N_5248,N_5181);
nor U5374 (N_5374,N_5149,N_5161);
or U5375 (N_5375,N_5302,N_5278);
and U5376 (N_5376,N_5283,N_5298);
xnor U5377 (N_5377,N_5254,N_5364);
and U5378 (N_5378,N_5332,N_5284);
xnor U5379 (N_5379,N_5367,N_5337);
xnor U5380 (N_5380,N_5296,N_5366);
nand U5381 (N_5381,N_5311,N_5357);
nand U5382 (N_5382,N_5279,N_5318);
or U5383 (N_5383,N_5313,N_5307);
and U5384 (N_5384,N_5358,N_5286);
nor U5385 (N_5385,N_5312,N_5350);
nor U5386 (N_5386,N_5320,N_5263);
nor U5387 (N_5387,N_5285,N_5370);
and U5388 (N_5388,N_5309,N_5356);
and U5389 (N_5389,N_5329,N_5333);
nor U5390 (N_5390,N_5251,N_5342);
nor U5391 (N_5391,N_5314,N_5335);
or U5392 (N_5392,N_5346,N_5322);
nor U5393 (N_5393,N_5294,N_5310);
and U5394 (N_5394,N_5303,N_5272);
and U5395 (N_5395,N_5345,N_5280);
xor U5396 (N_5396,N_5273,N_5261);
xor U5397 (N_5397,N_5324,N_5252);
and U5398 (N_5398,N_5316,N_5300);
nand U5399 (N_5399,N_5372,N_5266);
and U5400 (N_5400,N_5321,N_5349);
or U5401 (N_5401,N_5374,N_5269);
and U5402 (N_5402,N_5361,N_5327);
or U5403 (N_5403,N_5275,N_5338);
xor U5404 (N_5404,N_5362,N_5336);
or U5405 (N_5405,N_5258,N_5369);
nand U5406 (N_5406,N_5267,N_5293);
nand U5407 (N_5407,N_5257,N_5353);
and U5408 (N_5408,N_5325,N_5290);
and U5409 (N_5409,N_5326,N_5264);
or U5410 (N_5410,N_5347,N_5323);
or U5411 (N_5411,N_5304,N_5271);
and U5412 (N_5412,N_5355,N_5295);
nor U5413 (N_5413,N_5330,N_5343);
xnor U5414 (N_5414,N_5354,N_5351);
or U5415 (N_5415,N_5253,N_5334);
and U5416 (N_5416,N_5339,N_5373);
or U5417 (N_5417,N_5262,N_5291);
and U5418 (N_5418,N_5292,N_5319);
nor U5419 (N_5419,N_5315,N_5365);
nand U5420 (N_5420,N_5297,N_5268);
nand U5421 (N_5421,N_5259,N_5348);
and U5422 (N_5422,N_5317,N_5363);
and U5423 (N_5423,N_5305,N_5352);
nor U5424 (N_5424,N_5299,N_5341);
nor U5425 (N_5425,N_5331,N_5368);
and U5426 (N_5426,N_5360,N_5301);
xor U5427 (N_5427,N_5277,N_5288);
nor U5428 (N_5428,N_5328,N_5265);
and U5429 (N_5429,N_5359,N_5306);
nor U5430 (N_5430,N_5371,N_5282);
and U5431 (N_5431,N_5276,N_5274);
or U5432 (N_5432,N_5281,N_5255);
nor U5433 (N_5433,N_5344,N_5289);
xor U5434 (N_5434,N_5340,N_5260);
nor U5435 (N_5435,N_5287,N_5250);
or U5436 (N_5436,N_5308,N_5270);
and U5437 (N_5437,N_5256,N_5291);
nor U5438 (N_5438,N_5322,N_5323);
and U5439 (N_5439,N_5251,N_5333);
and U5440 (N_5440,N_5371,N_5285);
or U5441 (N_5441,N_5332,N_5363);
xor U5442 (N_5442,N_5320,N_5363);
nor U5443 (N_5443,N_5352,N_5291);
and U5444 (N_5444,N_5292,N_5334);
nor U5445 (N_5445,N_5263,N_5272);
xor U5446 (N_5446,N_5302,N_5270);
nand U5447 (N_5447,N_5359,N_5298);
and U5448 (N_5448,N_5336,N_5287);
or U5449 (N_5449,N_5364,N_5288);
and U5450 (N_5450,N_5363,N_5299);
and U5451 (N_5451,N_5307,N_5359);
nor U5452 (N_5452,N_5356,N_5265);
and U5453 (N_5453,N_5281,N_5336);
nand U5454 (N_5454,N_5266,N_5343);
and U5455 (N_5455,N_5316,N_5304);
and U5456 (N_5456,N_5317,N_5327);
and U5457 (N_5457,N_5337,N_5250);
or U5458 (N_5458,N_5348,N_5351);
and U5459 (N_5459,N_5351,N_5276);
nor U5460 (N_5460,N_5284,N_5350);
and U5461 (N_5461,N_5263,N_5361);
or U5462 (N_5462,N_5332,N_5301);
or U5463 (N_5463,N_5254,N_5256);
nor U5464 (N_5464,N_5268,N_5299);
nor U5465 (N_5465,N_5260,N_5310);
and U5466 (N_5466,N_5302,N_5269);
and U5467 (N_5467,N_5306,N_5304);
nand U5468 (N_5468,N_5359,N_5285);
nand U5469 (N_5469,N_5373,N_5298);
xor U5470 (N_5470,N_5281,N_5333);
xnor U5471 (N_5471,N_5285,N_5352);
or U5472 (N_5472,N_5343,N_5260);
xor U5473 (N_5473,N_5279,N_5296);
and U5474 (N_5474,N_5260,N_5313);
and U5475 (N_5475,N_5354,N_5250);
and U5476 (N_5476,N_5255,N_5292);
or U5477 (N_5477,N_5280,N_5305);
xor U5478 (N_5478,N_5313,N_5332);
or U5479 (N_5479,N_5353,N_5320);
xnor U5480 (N_5480,N_5364,N_5308);
nand U5481 (N_5481,N_5272,N_5348);
xor U5482 (N_5482,N_5271,N_5308);
xnor U5483 (N_5483,N_5260,N_5354);
and U5484 (N_5484,N_5321,N_5254);
xor U5485 (N_5485,N_5252,N_5351);
nor U5486 (N_5486,N_5258,N_5343);
xnor U5487 (N_5487,N_5334,N_5274);
nor U5488 (N_5488,N_5322,N_5305);
nor U5489 (N_5489,N_5286,N_5265);
nor U5490 (N_5490,N_5352,N_5299);
nor U5491 (N_5491,N_5346,N_5266);
xnor U5492 (N_5492,N_5270,N_5329);
xnor U5493 (N_5493,N_5352,N_5250);
or U5494 (N_5494,N_5275,N_5334);
nand U5495 (N_5495,N_5333,N_5266);
xnor U5496 (N_5496,N_5272,N_5365);
or U5497 (N_5497,N_5308,N_5255);
nor U5498 (N_5498,N_5270,N_5256);
and U5499 (N_5499,N_5365,N_5308);
or U5500 (N_5500,N_5458,N_5393);
or U5501 (N_5501,N_5481,N_5433);
xor U5502 (N_5502,N_5435,N_5400);
nand U5503 (N_5503,N_5434,N_5467);
xor U5504 (N_5504,N_5406,N_5407);
or U5505 (N_5505,N_5475,N_5487);
nor U5506 (N_5506,N_5402,N_5454);
or U5507 (N_5507,N_5381,N_5494);
xor U5508 (N_5508,N_5392,N_5482);
xor U5509 (N_5509,N_5491,N_5399);
xor U5510 (N_5510,N_5438,N_5391);
nor U5511 (N_5511,N_5470,N_5476);
and U5512 (N_5512,N_5429,N_5414);
and U5513 (N_5513,N_5445,N_5442);
xor U5514 (N_5514,N_5449,N_5468);
and U5515 (N_5515,N_5410,N_5462);
and U5516 (N_5516,N_5428,N_5375);
nand U5517 (N_5517,N_5387,N_5473);
or U5518 (N_5518,N_5466,N_5437);
nor U5519 (N_5519,N_5484,N_5424);
xor U5520 (N_5520,N_5453,N_5384);
xor U5521 (N_5521,N_5403,N_5499);
and U5522 (N_5522,N_5451,N_5418);
nand U5523 (N_5523,N_5404,N_5452);
nor U5524 (N_5524,N_5379,N_5408);
nand U5525 (N_5525,N_5465,N_5448);
nor U5526 (N_5526,N_5380,N_5432);
and U5527 (N_5527,N_5478,N_5385);
nand U5528 (N_5528,N_5405,N_5456);
nand U5529 (N_5529,N_5457,N_5441);
and U5530 (N_5530,N_5490,N_5469);
or U5531 (N_5531,N_5413,N_5386);
and U5532 (N_5532,N_5383,N_5394);
nand U5533 (N_5533,N_5425,N_5398);
xnor U5534 (N_5534,N_5420,N_5388);
and U5535 (N_5535,N_5471,N_5417);
xnor U5536 (N_5536,N_5443,N_5464);
and U5537 (N_5537,N_5497,N_5423);
or U5538 (N_5538,N_5498,N_5382);
nand U5539 (N_5539,N_5463,N_5492);
xnor U5540 (N_5540,N_5415,N_5430);
nor U5541 (N_5541,N_5422,N_5376);
and U5542 (N_5542,N_5489,N_5421);
xor U5543 (N_5543,N_5397,N_5419);
or U5544 (N_5544,N_5488,N_5444);
or U5545 (N_5545,N_5495,N_5460);
nand U5546 (N_5546,N_5396,N_5411);
and U5547 (N_5547,N_5401,N_5440);
and U5548 (N_5548,N_5483,N_5446);
nand U5549 (N_5549,N_5395,N_5459);
or U5550 (N_5550,N_5455,N_5431);
nand U5551 (N_5551,N_5496,N_5377);
nand U5552 (N_5552,N_5416,N_5409);
nand U5553 (N_5553,N_5486,N_5479);
nand U5554 (N_5554,N_5378,N_5472);
nor U5555 (N_5555,N_5493,N_5474);
nand U5556 (N_5556,N_5390,N_5439);
nor U5557 (N_5557,N_5447,N_5480);
nor U5558 (N_5558,N_5427,N_5477);
or U5559 (N_5559,N_5461,N_5426);
nor U5560 (N_5560,N_5389,N_5436);
nor U5561 (N_5561,N_5485,N_5412);
and U5562 (N_5562,N_5450,N_5463);
or U5563 (N_5563,N_5442,N_5463);
nor U5564 (N_5564,N_5496,N_5489);
nand U5565 (N_5565,N_5454,N_5495);
nor U5566 (N_5566,N_5492,N_5443);
xnor U5567 (N_5567,N_5427,N_5431);
nor U5568 (N_5568,N_5466,N_5377);
and U5569 (N_5569,N_5456,N_5440);
and U5570 (N_5570,N_5392,N_5436);
xor U5571 (N_5571,N_5497,N_5470);
and U5572 (N_5572,N_5490,N_5387);
and U5573 (N_5573,N_5424,N_5492);
and U5574 (N_5574,N_5485,N_5378);
nor U5575 (N_5575,N_5439,N_5492);
nor U5576 (N_5576,N_5416,N_5419);
nor U5577 (N_5577,N_5400,N_5481);
xnor U5578 (N_5578,N_5441,N_5421);
or U5579 (N_5579,N_5447,N_5427);
nand U5580 (N_5580,N_5440,N_5408);
nand U5581 (N_5581,N_5460,N_5411);
nor U5582 (N_5582,N_5425,N_5390);
xor U5583 (N_5583,N_5377,N_5388);
and U5584 (N_5584,N_5421,N_5438);
nor U5585 (N_5585,N_5415,N_5480);
or U5586 (N_5586,N_5460,N_5497);
xnor U5587 (N_5587,N_5493,N_5445);
xnor U5588 (N_5588,N_5437,N_5407);
xnor U5589 (N_5589,N_5424,N_5382);
and U5590 (N_5590,N_5411,N_5406);
and U5591 (N_5591,N_5408,N_5455);
and U5592 (N_5592,N_5440,N_5446);
and U5593 (N_5593,N_5428,N_5401);
nand U5594 (N_5594,N_5491,N_5444);
nor U5595 (N_5595,N_5390,N_5441);
nor U5596 (N_5596,N_5471,N_5439);
and U5597 (N_5597,N_5425,N_5427);
nand U5598 (N_5598,N_5435,N_5394);
nor U5599 (N_5599,N_5385,N_5459);
and U5600 (N_5600,N_5451,N_5445);
nand U5601 (N_5601,N_5499,N_5482);
or U5602 (N_5602,N_5450,N_5408);
nand U5603 (N_5603,N_5439,N_5381);
xor U5604 (N_5604,N_5425,N_5448);
nand U5605 (N_5605,N_5421,N_5445);
and U5606 (N_5606,N_5476,N_5393);
xnor U5607 (N_5607,N_5452,N_5386);
nor U5608 (N_5608,N_5399,N_5444);
xnor U5609 (N_5609,N_5468,N_5386);
or U5610 (N_5610,N_5401,N_5412);
or U5611 (N_5611,N_5427,N_5388);
or U5612 (N_5612,N_5492,N_5461);
or U5613 (N_5613,N_5452,N_5494);
or U5614 (N_5614,N_5446,N_5493);
nor U5615 (N_5615,N_5498,N_5401);
nor U5616 (N_5616,N_5476,N_5404);
nor U5617 (N_5617,N_5392,N_5393);
and U5618 (N_5618,N_5409,N_5450);
and U5619 (N_5619,N_5430,N_5426);
or U5620 (N_5620,N_5406,N_5472);
xor U5621 (N_5621,N_5398,N_5457);
nand U5622 (N_5622,N_5451,N_5385);
nor U5623 (N_5623,N_5397,N_5426);
and U5624 (N_5624,N_5462,N_5393);
and U5625 (N_5625,N_5521,N_5567);
xnor U5626 (N_5626,N_5538,N_5615);
and U5627 (N_5627,N_5548,N_5512);
or U5628 (N_5628,N_5598,N_5610);
nand U5629 (N_5629,N_5570,N_5504);
and U5630 (N_5630,N_5537,N_5568);
xor U5631 (N_5631,N_5583,N_5579);
nand U5632 (N_5632,N_5531,N_5585);
xnor U5633 (N_5633,N_5618,N_5557);
nor U5634 (N_5634,N_5516,N_5520);
and U5635 (N_5635,N_5576,N_5543);
xor U5636 (N_5636,N_5549,N_5526);
xnor U5637 (N_5637,N_5573,N_5574);
and U5638 (N_5638,N_5571,N_5612);
and U5639 (N_5639,N_5536,N_5519);
nand U5640 (N_5640,N_5578,N_5503);
nand U5641 (N_5641,N_5550,N_5547);
nor U5642 (N_5642,N_5500,N_5590);
nand U5643 (N_5643,N_5624,N_5593);
nand U5644 (N_5644,N_5605,N_5559);
and U5645 (N_5645,N_5600,N_5502);
or U5646 (N_5646,N_5565,N_5603);
or U5647 (N_5647,N_5551,N_5561);
xor U5648 (N_5648,N_5611,N_5554);
nor U5649 (N_5649,N_5616,N_5544);
or U5650 (N_5650,N_5556,N_5621);
or U5651 (N_5651,N_5541,N_5528);
or U5652 (N_5652,N_5606,N_5511);
and U5653 (N_5653,N_5555,N_5507);
and U5654 (N_5654,N_5532,N_5607);
nor U5655 (N_5655,N_5501,N_5510);
and U5656 (N_5656,N_5533,N_5540);
nor U5657 (N_5657,N_5518,N_5523);
and U5658 (N_5658,N_5546,N_5595);
and U5659 (N_5659,N_5539,N_5614);
nand U5660 (N_5660,N_5506,N_5535);
nand U5661 (N_5661,N_5589,N_5545);
and U5662 (N_5662,N_5596,N_5552);
and U5663 (N_5663,N_5558,N_5602);
nand U5664 (N_5664,N_5563,N_5594);
nor U5665 (N_5665,N_5517,N_5623);
xnor U5666 (N_5666,N_5613,N_5586);
xor U5667 (N_5667,N_5542,N_5597);
nand U5668 (N_5668,N_5620,N_5527);
and U5669 (N_5669,N_5530,N_5508);
xor U5670 (N_5670,N_5505,N_5588);
xor U5671 (N_5671,N_5591,N_5587);
nand U5672 (N_5672,N_5529,N_5580);
and U5673 (N_5673,N_5599,N_5617);
xor U5674 (N_5674,N_5525,N_5619);
and U5675 (N_5675,N_5560,N_5509);
nor U5676 (N_5676,N_5608,N_5622);
or U5677 (N_5677,N_5534,N_5572);
xnor U5678 (N_5678,N_5575,N_5562);
xor U5679 (N_5679,N_5601,N_5569);
xnor U5680 (N_5680,N_5604,N_5514);
xnor U5681 (N_5681,N_5609,N_5515);
nor U5682 (N_5682,N_5513,N_5524);
xor U5683 (N_5683,N_5582,N_5581);
nand U5684 (N_5684,N_5577,N_5584);
xor U5685 (N_5685,N_5566,N_5592);
or U5686 (N_5686,N_5564,N_5522);
nand U5687 (N_5687,N_5553,N_5534);
nand U5688 (N_5688,N_5564,N_5587);
nor U5689 (N_5689,N_5544,N_5513);
xor U5690 (N_5690,N_5568,N_5617);
nand U5691 (N_5691,N_5561,N_5513);
or U5692 (N_5692,N_5512,N_5609);
or U5693 (N_5693,N_5590,N_5595);
nor U5694 (N_5694,N_5528,N_5593);
nand U5695 (N_5695,N_5554,N_5624);
and U5696 (N_5696,N_5518,N_5554);
or U5697 (N_5697,N_5589,N_5505);
nor U5698 (N_5698,N_5503,N_5537);
nand U5699 (N_5699,N_5554,N_5590);
or U5700 (N_5700,N_5561,N_5614);
or U5701 (N_5701,N_5554,N_5571);
or U5702 (N_5702,N_5557,N_5527);
or U5703 (N_5703,N_5517,N_5516);
and U5704 (N_5704,N_5528,N_5549);
or U5705 (N_5705,N_5592,N_5540);
nor U5706 (N_5706,N_5587,N_5520);
or U5707 (N_5707,N_5620,N_5617);
nor U5708 (N_5708,N_5503,N_5567);
xor U5709 (N_5709,N_5602,N_5567);
nand U5710 (N_5710,N_5570,N_5583);
xnor U5711 (N_5711,N_5504,N_5597);
and U5712 (N_5712,N_5558,N_5510);
nor U5713 (N_5713,N_5509,N_5590);
nand U5714 (N_5714,N_5536,N_5590);
xor U5715 (N_5715,N_5518,N_5575);
and U5716 (N_5716,N_5571,N_5585);
nand U5717 (N_5717,N_5571,N_5509);
xor U5718 (N_5718,N_5511,N_5504);
nor U5719 (N_5719,N_5552,N_5553);
nor U5720 (N_5720,N_5509,N_5615);
nand U5721 (N_5721,N_5555,N_5512);
and U5722 (N_5722,N_5613,N_5533);
nand U5723 (N_5723,N_5519,N_5513);
or U5724 (N_5724,N_5526,N_5590);
or U5725 (N_5725,N_5601,N_5542);
nand U5726 (N_5726,N_5570,N_5547);
nor U5727 (N_5727,N_5612,N_5606);
or U5728 (N_5728,N_5522,N_5505);
xnor U5729 (N_5729,N_5597,N_5614);
or U5730 (N_5730,N_5560,N_5609);
or U5731 (N_5731,N_5513,N_5610);
or U5732 (N_5732,N_5600,N_5505);
and U5733 (N_5733,N_5526,N_5571);
nor U5734 (N_5734,N_5564,N_5520);
or U5735 (N_5735,N_5564,N_5535);
and U5736 (N_5736,N_5603,N_5529);
or U5737 (N_5737,N_5513,N_5502);
nand U5738 (N_5738,N_5580,N_5528);
and U5739 (N_5739,N_5624,N_5515);
nor U5740 (N_5740,N_5529,N_5517);
nor U5741 (N_5741,N_5503,N_5538);
xor U5742 (N_5742,N_5550,N_5573);
nand U5743 (N_5743,N_5504,N_5517);
or U5744 (N_5744,N_5564,N_5548);
nand U5745 (N_5745,N_5566,N_5507);
or U5746 (N_5746,N_5616,N_5522);
nand U5747 (N_5747,N_5517,N_5552);
nor U5748 (N_5748,N_5565,N_5521);
nor U5749 (N_5749,N_5599,N_5502);
xor U5750 (N_5750,N_5712,N_5625);
nand U5751 (N_5751,N_5638,N_5708);
xor U5752 (N_5752,N_5646,N_5657);
xor U5753 (N_5753,N_5734,N_5694);
nand U5754 (N_5754,N_5651,N_5682);
nand U5755 (N_5755,N_5659,N_5701);
or U5756 (N_5756,N_5660,N_5663);
and U5757 (N_5757,N_5650,N_5669);
or U5758 (N_5758,N_5671,N_5749);
nor U5759 (N_5759,N_5632,N_5661);
or U5760 (N_5760,N_5656,N_5692);
nor U5761 (N_5761,N_5736,N_5639);
nand U5762 (N_5762,N_5667,N_5677);
nand U5763 (N_5763,N_5709,N_5680);
nand U5764 (N_5764,N_5704,N_5630);
nor U5765 (N_5765,N_5652,N_5728);
and U5766 (N_5766,N_5637,N_5733);
nor U5767 (N_5767,N_5732,N_5634);
nor U5768 (N_5768,N_5741,N_5668);
or U5769 (N_5769,N_5626,N_5722);
nor U5770 (N_5770,N_5628,N_5745);
and U5771 (N_5771,N_5719,N_5711);
nor U5772 (N_5772,N_5642,N_5687);
nor U5773 (N_5773,N_5735,N_5631);
and U5774 (N_5774,N_5698,N_5730);
or U5775 (N_5775,N_5744,N_5739);
or U5776 (N_5776,N_5643,N_5679);
or U5777 (N_5777,N_5673,N_5716);
nand U5778 (N_5778,N_5695,N_5681);
nor U5779 (N_5779,N_5636,N_5747);
or U5780 (N_5780,N_5635,N_5738);
and U5781 (N_5781,N_5721,N_5743);
xor U5782 (N_5782,N_5714,N_5737);
or U5783 (N_5783,N_5720,N_5648);
or U5784 (N_5784,N_5700,N_5693);
or U5785 (N_5785,N_5665,N_5678);
nand U5786 (N_5786,N_5666,N_5746);
or U5787 (N_5787,N_5702,N_5629);
or U5788 (N_5788,N_5710,N_5726);
nor U5789 (N_5789,N_5647,N_5748);
and U5790 (N_5790,N_5633,N_5627);
nand U5791 (N_5791,N_5691,N_5703);
xnor U5792 (N_5792,N_5705,N_5723);
or U5793 (N_5793,N_5729,N_5644);
nand U5794 (N_5794,N_5645,N_5683);
nor U5795 (N_5795,N_5672,N_5641);
nor U5796 (N_5796,N_5649,N_5707);
nand U5797 (N_5797,N_5706,N_5688);
nor U5798 (N_5798,N_5699,N_5697);
nand U5799 (N_5799,N_5674,N_5654);
nand U5800 (N_5800,N_5696,N_5715);
xnor U5801 (N_5801,N_5742,N_5725);
nor U5802 (N_5802,N_5718,N_5724);
xor U5803 (N_5803,N_5686,N_5655);
nor U5804 (N_5804,N_5731,N_5670);
xor U5805 (N_5805,N_5727,N_5658);
xor U5806 (N_5806,N_5675,N_5685);
or U5807 (N_5807,N_5713,N_5653);
or U5808 (N_5808,N_5684,N_5662);
xor U5809 (N_5809,N_5690,N_5717);
or U5810 (N_5810,N_5740,N_5689);
xor U5811 (N_5811,N_5664,N_5640);
or U5812 (N_5812,N_5676,N_5644);
and U5813 (N_5813,N_5647,N_5637);
xnor U5814 (N_5814,N_5722,N_5633);
xor U5815 (N_5815,N_5671,N_5668);
nor U5816 (N_5816,N_5717,N_5699);
nand U5817 (N_5817,N_5688,N_5642);
xor U5818 (N_5818,N_5739,N_5703);
or U5819 (N_5819,N_5685,N_5634);
nor U5820 (N_5820,N_5664,N_5670);
or U5821 (N_5821,N_5719,N_5700);
nand U5822 (N_5822,N_5703,N_5651);
nand U5823 (N_5823,N_5627,N_5708);
xnor U5824 (N_5824,N_5711,N_5733);
xor U5825 (N_5825,N_5717,N_5727);
xnor U5826 (N_5826,N_5661,N_5689);
xor U5827 (N_5827,N_5666,N_5683);
nand U5828 (N_5828,N_5685,N_5672);
xor U5829 (N_5829,N_5703,N_5676);
xor U5830 (N_5830,N_5749,N_5665);
nand U5831 (N_5831,N_5698,N_5655);
xor U5832 (N_5832,N_5648,N_5710);
nand U5833 (N_5833,N_5740,N_5682);
xnor U5834 (N_5834,N_5735,N_5730);
xor U5835 (N_5835,N_5694,N_5715);
and U5836 (N_5836,N_5737,N_5749);
and U5837 (N_5837,N_5706,N_5703);
nor U5838 (N_5838,N_5689,N_5649);
or U5839 (N_5839,N_5740,N_5650);
nand U5840 (N_5840,N_5700,N_5694);
and U5841 (N_5841,N_5713,N_5712);
and U5842 (N_5842,N_5749,N_5733);
and U5843 (N_5843,N_5632,N_5700);
nand U5844 (N_5844,N_5631,N_5709);
nor U5845 (N_5845,N_5732,N_5674);
or U5846 (N_5846,N_5745,N_5672);
nand U5847 (N_5847,N_5671,N_5723);
nor U5848 (N_5848,N_5689,N_5673);
nor U5849 (N_5849,N_5704,N_5726);
and U5850 (N_5850,N_5644,N_5722);
and U5851 (N_5851,N_5689,N_5716);
nor U5852 (N_5852,N_5649,N_5650);
nor U5853 (N_5853,N_5739,N_5652);
nand U5854 (N_5854,N_5692,N_5671);
or U5855 (N_5855,N_5748,N_5667);
or U5856 (N_5856,N_5713,N_5656);
nor U5857 (N_5857,N_5684,N_5687);
xor U5858 (N_5858,N_5721,N_5678);
xnor U5859 (N_5859,N_5692,N_5711);
or U5860 (N_5860,N_5724,N_5685);
and U5861 (N_5861,N_5734,N_5692);
xnor U5862 (N_5862,N_5743,N_5690);
nand U5863 (N_5863,N_5632,N_5635);
xnor U5864 (N_5864,N_5699,N_5743);
nand U5865 (N_5865,N_5646,N_5738);
or U5866 (N_5866,N_5632,N_5704);
nand U5867 (N_5867,N_5711,N_5723);
and U5868 (N_5868,N_5690,N_5661);
xor U5869 (N_5869,N_5681,N_5650);
nand U5870 (N_5870,N_5639,N_5652);
nor U5871 (N_5871,N_5738,N_5690);
nor U5872 (N_5872,N_5664,N_5644);
and U5873 (N_5873,N_5662,N_5633);
nor U5874 (N_5874,N_5719,N_5722);
nand U5875 (N_5875,N_5752,N_5842);
nand U5876 (N_5876,N_5764,N_5852);
nand U5877 (N_5877,N_5869,N_5756);
nor U5878 (N_5878,N_5784,N_5793);
xor U5879 (N_5879,N_5754,N_5782);
or U5880 (N_5880,N_5772,N_5812);
nor U5881 (N_5881,N_5801,N_5779);
xor U5882 (N_5882,N_5773,N_5849);
nor U5883 (N_5883,N_5800,N_5861);
or U5884 (N_5884,N_5817,N_5848);
xnor U5885 (N_5885,N_5765,N_5873);
nor U5886 (N_5886,N_5831,N_5826);
nor U5887 (N_5887,N_5838,N_5818);
nand U5888 (N_5888,N_5802,N_5868);
and U5889 (N_5889,N_5872,N_5792);
and U5890 (N_5890,N_5769,N_5836);
nand U5891 (N_5891,N_5790,N_5846);
xor U5892 (N_5892,N_5770,N_5858);
or U5893 (N_5893,N_5821,N_5803);
or U5894 (N_5894,N_5761,N_5820);
nor U5895 (N_5895,N_5796,N_5808);
or U5896 (N_5896,N_5867,N_5751);
xnor U5897 (N_5897,N_5777,N_5798);
nand U5898 (N_5898,N_5788,N_5766);
and U5899 (N_5899,N_5755,N_5822);
or U5900 (N_5900,N_5813,N_5843);
xnor U5901 (N_5901,N_5827,N_5864);
nand U5902 (N_5902,N_5799,N_5816);
or U5903 (N_5903,N_5865,N_5795);
and U5904 (N_5904,N_5760,N_5762);
xnor U5905 (N_5905,N_5841,N_5758);
and U5906 (N_5906,N_5797,N_5791);
or U5907 (N_5907,N_5856,N_5809);
nand U5908 (N_5908,N_5763,N_5805);
or U5909 (N_5909,N_5767,N_5845);
nor U5910 (N_5910,N_5815,N_5750);
nand U5911 (N_5911,N_5854,N_5871);
and U5912 (N_5912,N_5794,N_5810);
xor U5913 (N_5913,N_5804,N_5862);
nand U5914 (N_5914,N_5857,N_5850);
nor U5915 (N_5915,N_5823,N_5870);
xor U5916 (N_5916,N_5829,N_5771);
or U5917 (N_5917,N_5847,N_5819);
xnor U5918 (N_5918,N_5859,N_5806);
or U5919 (N_5919,N_5783,N_5757);
xor U5920 (N_5920,N_5759,N_5853);
xnor U5921 (N_5921,N_5775,N_5866);
xnor U5922 (N_5922,N_5830,N_5814);
nand U5923 (N_5923,N_5837,N_5753);
nand U5924 (N_5924,N_5781,N_5824);
or U5925 (N_5925,N_5786,N_5785);
xor U5926 (N_5926,N_5833,N_5778);
nand U5927 (N_5927,N_5811,N_5851);
nand U5928 (N_5928,N_5825,N_5863);
nor U5929 (N_5929,N_5776,N_5834);
nand U5930 (N_5930,N_5768,N_5828);
or U5931 (N_5931,N_5860,N_5835);
xor U5932 (N_5932,N_5780,N_5789);
nand U5933 (N_5933,N_5874,N_5787);
or U5934 (N_5934,N_5855,N_5844);
nand U5935 (N_5935,N_5832,N_5839);
xor U5936 (N_5936,N_5774,N_5807);
nand U5937 (N_5937,N_5840,N_5814);
and U5938 (N_5938,N_5872,N_5870);
or U5939 (N_5939,N_5780,N_5867);
and U5940 (N_5940,N_5795,N_5809);
nand U5941 (N_5941,N_5817,N_5783);
xor U5942 (N_5942,N_5796,N_5751);
or U5943 (N_5943,N_5803,N_5867);
and U5944 (N_5944,N_5769,N_5794);
nand U5945 (N_5945,N_5853,N_5811);
and U5946 (N_5946,N_5797,N_5801);
xnor U5947 (N_5947,N_5801,N_5770);
and U5948 (N_5948,N_5765,N_5858);
xnor U5949 (N_5949,N_5762,N_5761);
and U5950 (N_5950,N_5820,N_5772);
xnor U5951 (N_5951,N_5775,N_5767);
nand U5952 (N_5952,N_5751,N_5813);
nor U5953 (N_5953,N_5829,N_5784);
xnor U5954 (N_5954,N_5823,N_5753);
or U5955 (N_5955,N_5783,N_5756);
nor U5956 (N_5956,N_5870,N_5838);
or U5957 (N_5957,N_5752,N_5775);
or U5958 (N_5958,N_5814,N_5779);
and U5959 (N_5959,N_5780,N_5776);
nor U5960 (N_5960,N_5831,N_5780);
and U5961 (N_5961,N_5852,N_5763);
xor U5962 (N_5962,N_5799,N_5752);
xor U5963 (N_5963,N_5774,N_5845);
xnor U5964 (N_5964,N_5757,N_5825);
nand U5965 (N_5965,N_5814,N_5870);
or U5966 (N_5966,N_5847,N_5811);
or U5967 (N_5967,N_5865,N_5841);
xor U5968 (N_5968,N_5848,N_5853);
nand U5969 (N_5969,N_5756,N_5815);
nor U5970 (N_5970,N_5860,N_5817);
nand U5971 (N_5971,N_5869,N_5760);
xor U5972 (N_5972,N_5765,N_5774);
xnor U5973 (N_5973,N_5818,N_5788);
and U5974 (N_5974,N_5831,N_5821);
and U5975 (N_5975,N_5860,N_5792);
or U5976 (N_5976,N_5793,N_5844);
nand U5977 (N_5977,N_5830,N_5844);
or U5978 (N_5978,N_5873,N_5803);
nand U5979 (N_5979,N_5845,N_5835);
and U5980 (N_5980,N_5869,N_5847);
or U5981 (N_5981,N_5797,N_5796);
and U5982 (N_5982,N_5845,N_5806);
nor U5983 (N_5983,N_5850,N_5828);
nand U5984 (N_5984,N_5809,N_5764);
xnor U5985 (N_5985,N_5859,N_5863);
or U5986 (N_5986,N_5753,N_5768);
or U5987 (N_5987,N_5854,N_5789);
or U5988 (N_5988,N_5830,N_5756);
nor U5989 (N_5989,N_5859,N_5846);
or U5990 (N_5990,N_5810,N_5753);
nor U5991 (N_5991,N_5835,N_5855);
and U5992 (N_5992,N_5794,N_5840);
or U5993 (N_5993,N_5845,N_5841);
nand U5994 (N_5994,N_5761,N_5812);
or U5995 (N_5995,N_5870,N_5772);
or U5996 (N_5996,N_5837,N_5756);
and U5997 (N_5997,N_5843,N_5821);
nor U5998 (N_5998,N_5785,N_5820);
or U5999 (N_5999,N_5867,N_5762);
nor U6000 (N_6000,N_5934,N_5921);
and U6001 (N_6001,N_5927,N_5995);
and U6002 (N_6002,N_5942,N_5945);
nor U6003 (N_6003,N_5981,N_5959);
xnor U6004 (N_6004,N_5930,N_5939);
nand U6005 (N_6005,N_5929,N_5974);
nand U6006 (N_6006,N_5931,N_5887);
or U6007 (N_6007,N_5966,N_5989);
nor U6008 (N_6008,N_5976,N_5902);
and U6009 (N_6009,N_5968,N_5965);
nor U6010 (N_6010,N_5890,N_5960);
nor U6011 (N_6011,N_5940,N_5971);
or U6012 (N_6012,N_5954,N_5952);
nor U6013 (N_6013,N_5967,N_5932);
nor U6014 (N_6014,N_5910,N_5913);
and U6015 (N_6015,N_5912,N_5889);
or U6016 (N_6016,N_5922,N_5969);
xnor U6017 (N_6017,N_5920,N_5951);
nand U6018 (N_6018,N_5992,N_5899);
xor U6019 (N_6019,N_5955,N_5944);
nor U6020 (N_6020,N_5987,N_5916);
or U6021 (N_6021,N_5915,N_5982);
xor U6022 (N_6022,N_5886,N_5879);
nand U6023 (N_6023,N_5880,N_5990);
nor U6024 (N_6024,N_5958,N_5897);
nor U6025 (N_6025,N_5948,N_5893);
xnor U6026 (N_6026,N_5972,N_5875);
nor U6027 (N_6027,N_5923,N_5894);
nand U6028 (N_6028,N_5993,N_5947);
or U6029 (N_6029,N_5996,N_5973);
and U6030 (N_6030,N_5888,N_5956);
nand U6031 (N_6031,N_5891,N_5878);
nor U6032 (N_6032,N_5949,N_5918);
and U6033 (N_6033,N_5986,N_5914);
nor U6034 (N_6034,N_5896,N_5957);
nand U6035 (N_6035,N_5928,N_5963);
or U6036 (N_6036,N_5881,N_5883);
xor U6037 (N_6037,N_5905,N_5877);
nand U6038 (N_6038,N_5911,N_5898);
or U6039 (N_6039,N_5926,N_5984);
xnor U6040 (N_6040,N_5950,N_5937);
and U6041 (N_6041,N_5909,N_5980);
nand U6042 (N_6042,N_5991,N_5941);
nor U6043 (N_6043,N_5903,N_5964);
xnor U6044 (N_6044,N_5876,N_5975);
or U6045 (N_6045,N_5983,N_5994);
and U6046 (N_6046,N_5884,N_5978);
nor U6047 (N_6047,N_5999,N_5953);
and U6048 (N_6048,N_5900,N_5882);
nor U6049 (N_6049,N_5892,N_5936);
nor U6050 (N_6050,N_5998,N_5907);
and U6051 (N_6051,N_5988,N_5935);
and U6052 (N_6052,N_5997,N_5895);
and U6053 (N_6053,N_5908,N_5985);
nand U6054 (N_6054,N_5906,N_5962);
and U6055 (N_6055,N_5917,N_5943);
xor U6056 (N_6056,N_5885,N_5970);
nand U6057 (N_6057,N_5977,N_5961);
or U6058 (N_6058,N_5946,N_5904);
and U6059 (N_6059,N_5925,N_5901);
xor U6060 (N_6060,N_5938,N_5933);
and U6061 (N_6061,N_5979,N_5919);
nand U6062 (N_6062,N_5924,N_5884);
and U6063 (N_6063,N_5954,N_5948);
nor U6064 (N_6064,N_5897,N_5947);
nor U6065 (N_6065,N_5972,N_5966);
nor U6066 (N_6066,N_5878,N_5915);
nand U6067 (N_6067,N_5883,N_5970);
or U6068 (N_6068,N_5889,N_5981);
and U6069 (N_6069,N_5930,N_5898);
xor U6070 (N_6070,N_5893,N_5909);
xor U6071 (N_6071,N_5994,N_5954);
xnor U6072 (N_6072,N_5968,N_5966);
and U6073 (N_6073,N_5963,N_5941);
nor U6074 (N_6074,N_5894,N_5896);
nand U6075 (N_6075,N_5910,N_5997);
and U6076 (N_6076,N_5887,N_5986);
or U6077 (N_6077,N_5986,N_5915);
nand U6078 (N_6078,N_5909,N_5902);
xor U6079 (N_6079,N_5957,N_5991);
and U6080 (N_6080,N_5960,N_5963);
and U6081 (N_6081,N_5932,N_5984);
xor U6082 (N_6082,N_5950,N_5992);
or U6083 (N_6083,N_5904,N_5886);
or U6084 (N_6084,N_5892,N_5989);
nor U6085 (N_6085,N_5887,N_5926);
or U6086 (N_6086,N_5909,N_5963);
and U6087 (N_6087,N_5963,N_5913);
or U6088 (N_6088,N_5905,N_5944);
nand U6089 (N_6089,N_5986,N_5932);
nand U6090 (N_6090,N_5883,N_5927);
nor U6091 (N_6091,N_5920,N_5996);
or U6092 (N_6092,N_5979,N_5929);
xor U6093 (N_6093,N_5893,N_5902);
or U6094 (N_6094,N_5970,N_5915);
nand U6095 (N_6095,N_5882,N_5988);
xnor U6096 (N_6096,N_5977,N_5922);
nand U6097 (N_6097,N_5896,N_5989);
xor U6098 (N_6098,N_5986,N_5960);
or U6099 (N_6099,N_5888,N_5925);
nor U6100 (N_6100,N_5951,N_5955);
and U6101 (N_6101,N_5909,N_5988);
nand U6102 (N_6102,N_5918,N_5899);
nand U6103 (N_6103,N_5997,N_5916);
xor U6104 (N_6104,N_5970,N_5960);
and U6105 (N_6105,N_5891,N_5932);
nor U6106 (N_6106,N_5946,N_5910);
nor U6107 (N_6107,N_5956,N_5984);
and U6108 (N_6108,N_5970,N_5878);
and U6109 (N_6109,N_5958,N_5934);
or U6110 (N_6110,N_5891,N_5992);
or U6111 (N_6111,N_5920,N_5878);
or U6112 (N_6112,N_5948,N_5897);
or U6113 (N_6113,N_5893,N_5886);
xnor U6114 (N_6114,N_5937,N_5911);
nand U6115 (N_6115,N_5977,N_5897);
xnor U6116 (N_6116,N_5910,N_5885);
and U6117 (N_6117,N_5954,N_5880);
xnor U6118 (N_6118,N_5957,N_5875);
and U6119 (N_6119,N_5888,N_5884);
nor U6120 (N_6120,N_5906,N_5913);
nand U6121 (N_6121,N_5979,N_5959);
nand U6122 (N_6122,N_5942,N_5895);
xnor U6123 (N_6123,N_5920,N_5875);
nand U6124 (N_6124,N_5960,N_5924);
and U6125 (N_6125,N_6118,N_6022);
nand U6126 (N_6126,N_6034,N_6048);
xnor U6127 (N_6127,N_6049,N_6013);
nor U6128 (N_6128,N_6018,N_6116);
xnor U6129 (N_6129,N_6062,N_6037);
or U6130 (N_6130,N_6088,N_6072);
or U6131 (N_6131,N_6066,N_6039);
xor U6132 (N_6132,N_6094,N_6036);
nor U6133 (N_6133,N_6108,N_6053);
nand U6134 (N_6134,N_6083,N_6006);
xnor U6135 (N_6135,N_6026,N_6014);
or U6136 (N_6136,N_6112,N_6106);
or U6137 (N_6137,N_6033,N_6040);
xor U6138 (N_6138,N_6016,N_6110);
and U6139 (N_6139,N_6114,N_6024);
nand U6140 (N_6140,N_6002,N_6020);
and U6141 (N_6141,N_6044,N_6052);
xnor U6142 (N_6142,N_6085,N_6084);
nand U6143 (N_6143,N_6068,N_6025);
or U6144 (N_6144,N_6071,N_6031);
and U6145 (N_6145,N_6001,N_6007);
nor U6146 (N_6146,N_6050,N_6059);
and U6147 (N_6147,N_6117,N_6086);
or U6148 (N_6148,N_6087,N_6065);
nand U6149 (N_6149,N_6092,N_6069);
xor U6150 (N_6150,N_6122,N_6028);
and U6151 (N_6151,N_6082,N_6099);
nor U6152 (N_6152,N_6113,N_6100);
or U6153 (N_6153,N_6077,N_6124);
xor U6154 (N_6154,N_6058,N_6035);
or U6155 (N_6155,N_6095,N_6096);
and U6156 (N_6156,N_6063,N_6019);
nor U6157 (N_6157,N_6093,N_6073);
nor U6158 (N_6158,N_6107,N_6023);
nor U6159 (N_6159,N_6115,N_6098);
xor U6160 (N_6160,N_6027,N_6080);
nand U6161 (N_6161,N_6089,N_6057);
or U6162 (N_6162,N_6032,N_6038);
or U6163 (N_6163,N_6119,N_6079);
nor U6164 (N_6164,N_6012,N_6067);
xnor U6165 (N_6165,N_6015,N_6060);
xor U6166 (N_6166,N_6104,N_6074);
xnor U6167 (N_6167,N_6091,N_6005);
and U6168 (N_6168,N_6055,N_6064);
and U6169 (N_6169,N_6041,N_6105);
xnor U6170 (N_6170,N_6003,N_6004);
xnor U6171 (N_6171,N_6030,N_6021);
or U6172 (N_6172,N_6090,N_6123);
and U6173 (N_6173,N_6010,N_6097);
xor U6174 (N_6174,N_6054,N_6046);
or U6175 (N_6175,N_6120,N_6009);
nor U6176 (N_6176,N_6102,N_6045);
or U6177 (N_6177,N_6078,N_6029);
or U6178 (N_6178,N_6061,N_6075);
nand U6179 (N_6179,N_6056,N_6109);
nor U6180 (N_6180,N_6008,N_6101);
nor U6181 (N_6181,N_6047,N_6076);
xor U6182 (N_6182,N_6111,N_6051);
xnor U6183 (N_6183,N_6017,N_6081);
or U6184 (N_6184,N_6043,N_6121);
nor U6185 (N_6185,N_6070,N_6103);
or U6186 (N_6186,N_6000,N_6011);
xor U6187 (N_6187,N_6042,N_6122);
and U6188 (N_6188,N_6090,N_6088);
nor U6189 (N_6189,N_6014,N_6109);
nor U6190 (N_6190,N_6077,N_6098);
or U6191 (N_6191,N_6040,N_6092);
nor U6192 (N_6192,N_6052,N_6072);
nor U6193 (N_6193,N_6000,N_6013);
nand U6194 (N_6194,N_6035,N_6085);
nand U6195 (N_6195,N_6121,N_6074);
and U6196 (N_6196,N_6099,N_6085);
nand U6197 (N_6197,N_6118,N_6120);
and U6198 (N_6198,N_6044,N_6106);
nand U6199 (N_6199,N_6078,N_6102);
and U6200 (N_6200,N_6075,N_6016);
nand U6201 (N_6201,N_6101,N_6089);
or U6202 (N_6202,N_6086,N_6033);
xnor U6203 (N_6203,N_6022,N_6024);
or U6204 (N_6204,N_6089,N_6012);
nor U6205 (N_6205,N_6030,N_6065);
xor U6206 (N_6206,N_6036,N_6013);
and U6207 (N_6207,N_6035,N_6095);
nor U6208 (N_6208,N_6009,N_6004);
nor U6209 (N_6209,N_6017,N_6087);
and U6210 (N_6210,N_6120,N_6079);
and U6211 (N_6211,N_6115,N_6123);
or U6212 (N_6212,N_6047,N_6057);
nand U6213 (N_6213,N_6113,N_6124);
and U6214 (N_6214,N_6025,N_6070);
and U6215 (N_6215,N_6072,N_6112);
and U6216 (N_6216,N_6085,N_6055);
and U6217 (N_6217,N_6018,N_6017);
or U6218 (N_6218,N_6124,N_6050);
or U6219 (N_6219,N_6048,N_6071);
and U6220 (N_6220,N_6097,N_6080);
or U6221 (N_6221,N_6058,N_6008);
nand U6222 (N_6222,N_6039,N_6058);
nand U6223 (N_6223,N_6097,N_6115);
xnor U6224 (N_6224,N_6043,N_6059);
xnor U6225 (N_6225,N_6119,N_6102);
nand U6226 (N_6226,N_6093,N_6058);
and U6227 (N_6227,N_6069,N_6085);
nand U6228 (N_6228,N_6098,N_6073);
nor U6229 (N_6229,N_6020,N_6029);
xor U6230 (N_6230,N_6013,N_6020);
xnor U6231 (N_6231,N_6122,N_6084);
or U6232 (N_6232,N_6061,N_6066);
xor U6233 (N_6233,N_6069,N_6041);
nand U6234 (N_6234,N_6038,N_6045);
or U6235 (N_6235,N_6111,N_6045);
nand U6236 (N_6236,N_6109,N_6087);
or U6237 (N_6237,N_6084,N_6003);
and U6238 (N_6238,N_6034,N_6040);
nor U6239 (N_6239,N_6101,N_6058);
and U6240 (N_6240,N_6111,N_6046);
or U6241 (N_6241,N_6021,N_6089);
nor U6242 (N_6242,N_6107,N_6108);
or U6243 (N_6243,N_6074,N_6120);
xnor U6244 (N_6244,N_6094,N_6043);
and U6245 (N_6245,N_6002,N_6058);
xor U6246 (N_6246,N_6057,N_6026);
nor U6247 (N_6247,N_6044,N_6100);
nor U6248 (N_6248,N_6057,N_6032);
nor U6249 (N_6249,N_6087,N_6046);
xor U6250 (N_6250,N_6131,N_6230);
nor U6251 (N_6251,N_6151,N_6129);
nor U6252 (N_6252,N_6150,N_6158);
and U6253 (N_6253,N_6127,N_6139);
or U6254 (N_6254,N_6181,N_6223);
and U6255 (N_6255,N_6191,N_6170);
and U6256 (N_6256,N_6206,N_6198);
nand U6257 (N_6257,N_6217,N_6134);
and U6258 (N_6258,N_6167,N_6161);
nand U6259 (N_6259,N_6226,N_6200);
nor U6260 (N_6260,N_6140,N_6211);
or U6261 (N_6261,N_6188,N_6147);
nor U6262 (N_6262,N_6239,N_6241);
xor U6263 (N_6263,N_6232,N_6195);
nor U6264 (N_6264,N_6172,N_6235);
nor U6265 (N_6265,N_6125,N_6160);
and U6266 (N_6266,N_6197,N_6224);
xor U6267 (N_6267,N_6152,N_6185);
xnor U6268 (N_6268,N_6182,N_6174);
and U6269 (N_6269,N_6209,N_6229);
and U6270 (N_6270,N_6225,N_6218);
xnor U6271 (N_6271,N_6221,N_6242);
or U6272 (N_6272,N_6141,N_6190);
xnor U6273 (N_6273,N_6228,N_6154);
or U6274 (N_6274,N_6138,N_6192);
xor U6275 (N_6275,N_6149,N_6248);
nand U6276 (N_6276,N_6219,N_6184);
and U6277 (N_6277,N_6240,N_6136);
nand U6278 (N_6278,N_6178,N_6207);
or U6279 (N_6279,N_6231,N_6186);
or U6280 (N_6280,N_6133,N_6233);
nand U6281 (N_6281,N_6130,N_6204);
and U6282 (N_6282,N_6215,N_6165);
nand U6283 (N_6283,N_6214,N_6246);
nand U6284 (N_6284,N_6213,N_6205);
xor U6285 (N_6285,N_6238,N_6244);
or U6286 (N_6286,N_6171,N_6202);
or U6287 (N_6287,N_6146,N_6163);
xor U6288 (N_6288,N_6196,N_6143);
nand U6289 (N_6289,N_6245,N_6208);
nor U6290 (N_6290,N_6237,N_6159);
xor U6291 (N_6291,N_6135,N_6201);
nor U6292 (N_6292,N_6155,N_6128);
or U6293 (N_6293,N_6243,N_6212);
nor U6294 (N_6294,N_6168,N_6234);
xnor U6295 (N_6295,N_6210,N_6145);
xnor U6296 (N_6296,N_6144,N_6169);
nor U6297 (N_6297,N_6187,N_6203);
or U6298 (N_6298,N_6222,N_6164);
xor U6299 (N_6299,N_6249,N_6193);
nand U6300 (N_6300,N_6247,N_6194);
nor U6301 (N_6301,N_6148,N_6236);
and U6302 (N_6302,N_6179,N_6153);
nand U6303 (N_6303,N_6137,N_6199);
and U6304 (N_6304,N_6175,N_6177);
nand U6305 (N_6305,N_6189,N_6166);
nand U6306 (N_6306,N_6173,N_6176);
and U6307 (N_6307,N_6162,N_6220);
nand U6308 (N_6308,N_6227,N_6157);
nor U6309 (N_6309,N_6180,N_6156);
nand U6310 (N_6310,N_6126,N_6142);
or U6311 (N_6311,N_6183,N_6216);
nand U6312 (N_6312,N_6132,N_6174);
xor U6313 (N_6313,N_6173,N_6197);
or U6314 (N_6314,N_6198,N_6176);
nand U6315 (N_6315,N_6248,N_6147);
nor U6316 (N_6316,N_6134,N_6152);
and U6317 (N_6317,N_6173,N_6160);
xnor U6318 (N_6318,N_6138,N_6195);
xor U6319 (N_6319,N_6230,N_6193);
or U6320 (N_6320,N_6174,N_6227);
xnor U6321 (N_6321,N_6165,N_6141);
nor U6322 (N_6322,N_6186,N_6169);
nand U6323 (N_6323,N_6243,N_6127);
and U6324 (N_6324,N_6137,N_6128);
nor U6325 (N_6325,N_6146,N_6169);
nor U6326 (N_6326,N_6239,N_6186);
xor U6327 (N_6327,N_6249,N_6176);
nor U6328 (N_6328,N_6249,N_6241);
nor U6329 (N_6329,N_6186,N_6174);
nor U6330 (N_6330,N_6128,N_6201);
xor U6331 (N_6331,N_6130,N_6182);
or U6332 (N_6332,N_6216,N_6213);
nor U6333 (N_6333,N_6200,N_6234);
and U6334 (N_6334,N_6135,N_6244);
or U6335 (N_6335,N_6126,N_6169);
xnor U6336 (N_6336,N_6144,N_6126);
and U6337 (N_6337,N_6168,N_6231);
nand U6338 (N_6338,N_6172,N_6142);
xor U6339 (N_6339,N_6132,N_6126);
nor U6340 (N_6340,N_6147,N_6201);
nor U6341 (N_6341,N_6243,N_6219);
nand U6342 (N_6342,N_6201,N_6208);
xor U6343 (N_6343,N_6130,N_6151);
nand U6344 (N_6344,N_6228,N_6158);
or U6345 (N_6345,N_6148,N_6129);
and U6346 (N_6346,N_6150,N_6133);
and U6347 (N_6347,N_6160,N_6211);
or U6348 (N_6348,N_6132,N_6162);
and U6349 (N_6349,N_6198,N_6210);
nor U6350 (N_6350,N_6211,N_6221);
nor U6351 (N_6351,N_6158,N_6213);
xor U6352 (N_6352,N_6185,N_6132);
nand U6353 (N_6353,N_6186,N_6241);
nand U6354 (N_6354,N_6249,N_6127);
or U6355 (N_6355,N_6176,N_6192);
nand U6356 (N_6356,N_6237,N_6149);
nand U6357 (N_6357,N_6193,N_6217);
or U6358 (N_6358,N_6177,N_6134);
xnor U6359 (N_6359,N_6184,N_6210);
nand U6360 (N_6360,N_6237,N_6170);
or U6361 (N_6361,N_6201,N_6243);
or U6362 (N_6362,N_6133,N_6209);
nand U6363 (N_6363,N_6208,N_6168);
xor U6364 (N_6364,N_6163,N_6229);
or U6365 (N_6365,N_6219,N_6200);
or U6366 (N_6366,N_6183,N_6149);
or U6367 (N_6367,N_6239,N_6134);
or U6368 (N_6368,N_6229,N_6157);
or U6369 (N_6369,N_6214,N_6158);
nand U6370 (N_6370,N_6219,N_6171);
nand U6371 (N_6371,N_6241,N_6171);
nor U6372 (N_6372,N_6228,N_6156);
nor U6373 (N_6373,N_6218,N_6152);
or U6374 (N_6374,N_6238,N_6225);
and U6375 (N_6375,N_6318,N_6340);
and U6376 (N_6376,N_6310,N_6267);
or U6377 (N_6377,N_6280,N_6304);
and U6378 (N_6378,N_6329,N_6328);
and U6379 (N_6379,N_6322,N_6303);
and U6380 (N_6380,N_6314,N_6299);
nand U6381 (N_6381,N_6251,N_6356);
nor U6382 (N_6382,N_6273,N_6301);
or U6383 (N_6383,N_6282,N_6334);
xnor U6384 (N_6384,N_6275,N_6362);
xnor U6385 (N_6385,N_6263,N_6349);
nand U6386 (N_6386,N_6372,N_6353);
nand U6387 (N_6387,N_6320,N_6288);
nand U6388 (N_6388,N_6339,N_6250);
xor U6389 (N_6389,N_6291,N_6338);
nand U6390 (N_6390,N_6271,N_6326);
nor U6391 (N_6391,N_6346,N_6341);
xor U6392 (N_6392,N_6278,N_6295);
nor U6393 (N_6393,N_6313,N_6360);
nor U6394 (N_6394,N_6311,N_6281);
and U6395 (N_6395,N_6364,N_6266);
nor U6396 (N_6396,N_6309,N_6367);
nand U6397 (N_6397,N_6294,N_6293);
or U6398 (N_6398,N_6358,N_6373);
nand U6399 (N_6399,N_6359,N_6256);
xnor U6400 (N_6400,N_6371,N_6283);
xor U6401 (N_6401,N_6289,N_6255);
nand U6402 (N_6402,N_6369,N_6350);
or U6403 (N_6403,N_6302,N_6316);
and U6404 (N_6404,N_6305,N_6296);
or U6405 (N_6405,N_6317,N_6374);
nand U6406 (N_6406,N_6297,N_6269);
or U6407 (N_6407,N_6306,N_6337);
or U6408 (N_6408,N_6276,N_6270);
or U6409 (N_6409,N_6253,N_6254);
and U6410 (N_6410,N_6319,N_6327);
and U6411 (N_6411,N_6286,N_6352);
nand U6412 (N_6412,N_6307,N_6298);
xor U6413 (N_6413,N_6284,N_6261);
xor U6414 (N_6414,N_6324,N_6325);
or U6415 (N_6415,N_6312,N_6321);
and U6416 (N_6416,N_6257,N_6354);
or U6417 (N_6417,N_6330,N_6323);
xnor U6418 (N_6418,N_6260,N_6259);
nor U6419 (N_6419,N_6366,N_6351);
and U6420 (N_6420,N_6335,N_6331);
nor U6421 (N_6421,N_6264,N_6308);
xnor U6422 (N_6422,N_6347,N_6274);
xor U6423 (N_6423,N_6361,N_6343);
xnor U6424 (N_6424,N_6355,N_6290);
nand U6425 (N_6425,N_6262,N_6370);
nand U6426 (N_6426,N_6292,N_6348);
xnor U6427 (N_6427,N_6336,N_6363);
nor U6428 (N_6428,N_6277,N_6258);
xor U6429 (N_6429,N_6333,N_6252);
xor U6430 (N_6430,N_6365,N_6315);
nand U6431 (N_6431,N_6342,N_6268);
and U6432 (N_6432,N_6300,N_6332);
xnor U6433 (N_6433,N_6368,N_6285);
or U6434 (N_6434,N_6345,N_6357);
xor U6435 (N_6435,N_6279,N_6344);
nor U6436 (N_6436,N_6265,N_6272);
xnor U6437 (N_6437,N_6287,N_6303);
or U6438 (N_6438,N_6292,N_6311);
and U6439 (N_6439,N_6357,N_6365);
nand U6440 (N_6440,N_6316,N_6295);
and U6441 (N_6441,N_6312,N_6270);
nor U6442 (N_6442,N_6336,N_6345);
nand U6443 (N_6443,N_6365,N_6368);
xnor U6444 (N_6444,N_6349,N_6279);
nand U6445 (N_6445,N_6372,N_6361);
xor U6446 (N_6446,N_6307,N_6310);
nand U6447 (N_6447,N_6364,N_6298);
nor U6448 (N_6448,N_6273,N_6346);
and U6449 (N_6449,N_6312,N_6295);
or U6450 (N_6450,N_6282,N_6368);
or U6451 (N_6451,N_6341,N_6361);
or U6452 (N_6452,N_6307,N_6287);
xor U6453 (N_6453,N_6369,N_6295);
nand U6454 (N_6454,N_6335,N_6354);
nand U6455 (N_6455,N_6344,N_6299);
and U6456 (N_6456,N_6373,N_6338);
or U6457 (N_6457,N_6309,N_6353);
nor U6458 (N_6458,N_6274,N_6350);
and U6459 (N_6459,N_6353,N_6314);
xor U6460 (N_6460,N_6272,N_6345);
nor U6461 (N_6461,N_6304,N_6347);
nor U6462 (N_6462,N_6337,N_6328);
nor U6463 (N_6463,N_6275,N_6305);
xnor U6464 (N_6464,N_6369,N_6273);
nor U6465 (N_6465,N_6291,N_6275);
nor U6466 (N_6466,N_6254,N_6361);
xnor U6467 (N_6467,N_6328,N_6344);
or U6468 (N_6468,N_6296,N_6339);
xor U6469 (N_6469,N_6266,N_6278);
nand U6470 (N_6470,N_6262,N_6275);
nor U6471 (N_6471,N_6298,N_6311);
and U6472 (N_6472,N_6329,N_6326);
and U6473 (N_6473,N_6289,N_6327);
and U6474 (N_6474,N_6269,N_6306);
or U6475 (N_6475,N_6328,N_6293);
and U6476 (N_6476,N_6256,N_6270);
or U6477 (N_6477,N_6266,N_6362);
xor U6478 (N_6478,N_6363,N_6342);
xor U6479 (N_6479,N_6319,N_6270);
or U6480 (N_6480,N_6283,N_6364);
and U6481 (N_6481,N_6309,N_6251);
nand U6482 (N_6482,N_6370,N_6286);
xnor U6483 (N_6483,N_6372,N_6294);
or U6484 (N_6484,N_6359,N_6327);
nor U6485 (N_6485,N_6310,N_6331);
nor U6486 (N_6486,N_6297,N_6356);
nand U6487 (N_6487,N_6368,N_6331);
and U6488 (N_6488,N_6373,N_6276);
and U6489 (N_6489,N_6294,N_6350);
nand U6490 (N_6490,N_6282,N_6305);
nor U6491 (N_6491,N_6276,N_6318);
nor U6492 (N_6492,N_6298,N_6324);
nor U6493 (N_6493,N_6269,N_6343);
and U6494 (N_6494,N_6339,N_6268);
or U6495 (N_6495,N_6355,N_6261);
and U6496 (N_6496,N_6250,N_6357);
and U6497 (N_6497,N_6362,N_6308);
or U6498 (N_6498,N_6323,N_6334);
nor U6499 (N_6499,N_6265,N_6268);
or U6500 (N_6500,N_6450,N_6478);
and U6501 (N_6501,N_6439,N_6459);
xnor U6502 (N_6502,N_6412,N_6461);
xnor U6503 (N_6503,N_6383,N_6400);
xor U6504 (N_6504,N_6436,N_6470);
nor U6505 (N_6505,N_6446,N_6378);
xor U6506 (N_6506,N_6421,N_6396);
nand U6507 (N_6507,N_6460,N_6486);
xnor U6508 (N_6508,N_6402,N_6494);
or U6509 (N_6509,N_6492,N_6465);
or U6510 (N_6510,N_6405,N_6448);
and U6511 (N_6511,N_6379,N_6420);
nor U6512 (N_6512,N_6417,N_6476);
nor U6513 (N_6513,N_6406,N_6415);
or U6514 (N_6514,N_6388,N_6475);
nand U6515 (N_6515,N_6426,N_6471);
nand U6516 (N_6516,N_6449,N_6385);
and U6517 (N_6517,N_6483,N_6482);
or U6518 (N_6518,N_6466,N_6389);
and U6519 (N_6519,N_6463,N_6481);
nor U6520 (N_6520,N_6452,N_6462);
nand U6521 (N_6521,N_6432,N_6485);
nor U6522 (N_6522,N_6380,N_6435);
nand U6523 (N_6523,N_6422,N_6382);
nor U6524 (N_6524,N_6403,N_6376);
xnor U6525 (N_6525,N_6407,N_6458);
or U6526 (N_6526,N_6454,N_6427);
nor U6527 (N_6527,N_6445,N_6440);
nor U6528 (N_6528,N_6423,N_6387);
xnor U6529 (N_6529,N_6437,N_6392);
or U6530 (N_6530,N_6438,N_6425);
xor U6531 (N_6531,N_6457,N_6408);
xor U6532 (N_6532,N_6384,N_6409);
or U6533 (N_6533,N_6499,N_6473);
nand U6534 (N_6534,N_6493,N_6398);
nor U6535 (N_6535,N_6416,N_6419);
nor U6536 (N_6536,N_6429,N_6431);
and U6537 (N_6537,N_6455,N_6443);
nor U6538 (N_6538,N_6434,N_6498);
nand U6539 (N_6539,N_6451,N_6430);
nand U6540 (N_6540,N_6444,N_6488);
and U6541 (N_6541,N_6395,N_6472);
nor U6542 (N_6542,N_6484,N_6386);
xor U6543 (N_6543,N_6391,N_6424);
nand U6544 (N_6544,N_6487,N_6410);
nor U6545 (N_6545,N_6394,N_6397);
xnor U6546 (N_6546,N_6393,N_6399);
xnor U6547 (N_6547,N_6411,N_6418);
or U6548 (N_6548,N_6404,N_6442);
nor U6549 (N_6549,N_6467,N_6497);
nor U6550 (N_6550,N_6490,N_6468);
or U6551 (N_6551,N_6456,N_6413);
nor U6552 (N_6552,N_6377,N_6469);
nand U6553 (N_6553,N_6390,N_6401);
nand U6554 (N_6554,N_6441,N_6495);
or U6555 (N_6555,N_6453,N_6479);
and U6556 (N_6556,N_6464,N_6414);
nor U6557 (N_6557,N_6375,N_6381);
xnor U6558 (N_6558,N_6496,N_6480);
nor U6559 (N_6559,N_6491,N_6489);
xnor U6560 (N_6560,N_6477,N_6447);
nor U6561 (N_6561,N_6433,N_6474);
or U6562 (N_6562,N_6428,N_6396);
or U6563 (N_6563,N_6405,N_6467);
and U6564 (N_6564,N_6408,N_6472);
and U6565 (N_6565,N_6384,N_6492);
xnor U6566 (N_6566,N_6479,N_6420);
or U6567 (N_6567,N_6410,N_6406);
nor U6568 (N_6568,N_6440,N_6399);
nor U6569 (N_6569,N_6478,N_6462);
or U6570 (N_6570,N_6442,N_6449);
or U6571 (N_6571,N_6442,N_6429);
and U6572 (N_6572,N_6485,N_6421);
nand U6573 (N_6573,N_6457,N_6388);
and U6574 (N_6574,N_6472,N_6452);
nor U6575 (N_6575,N_6487,N_6460);
xor U6576 (N_6576,N_6439,N_6476);
xor U6577 (N_6577,N_6495,N_6415);
nor U6578 (N_6578,N_6489,N_6434);
nor U6579 (N_6579,N_6486,N_6427);
or U6580 (N_6580,N_6452,N_6438);
and U6581 (N_6581,N_6429,N_6444);
nand U6582 (N_6582,N_6477,N_6487);
nor U6583 (N_6583,N_6446,N_6392);
xnor U6584 (N_6584,N_6420,N_6435);
xnor U6585 (N_6585,N_6381,N_6477);
nand U6586 (N_6586,N_6414,N_6413);
xnor U6587 (N_6587,N_6409,N_6404);
and U6588 (N_6588,N_6440,N_6379);
xor U6589 (N_6589,N_6497,N_6446);
and U6590 (N_6590,N_6407,N_6468);
nand U6591 (N_6591,N_6474,N_6484);
or U6592 (N_6592,N_6385,N_6383);
xor U6593 (N_6593,N_6421,N_6379);
nand U6594 (N_6594,N_6376,N_6382);
xnor U6595 (N_6595,N_6474,N_6405);
and U6596 (N_6596,N_6426,N_6389);
or U6597 (N_6597,N_6418,N_6447);
and U6598 (N_6598,N_6482,N_6448);
or U6599 (N_6599,N_6462,N_6480);
or U6600 (N_6600,N_6454,N_6494);
xnor U6601 (N_6601,N_6401,N_6422);
xnor U6602 (N_6602,N_6392,N_6431);
nand U6603 (N_6603,N_6381,N_6463);
or U6604 (N_6604,N_6381,N_6487);
nor U6605 (N_6605,N_6467,N_6451);
nor U6606 (N_6606,N_6399,N_6443);
xor U6607 (N_6607,N_6381,N_6469);
nand U6608 (N_6608,N_6408,N_6474);
nand U6609 (N_6609,N_6434,N_6404);
or U6610 (N_6610,N_6428,N_6421);
nand U6611 (N_6611,N_6429,N_6446);
nand U6612 (N_6612,N_6448,N_6443);
nand U6613 (N_6613,N_6466,N_6419);
nand U6614 (N_6614,N_6465,N_6484);
and U6615 (N_6615,N_6478,N_6493);
nor U6616 (N_6616,N_6442,N_6498);
nand U6617 (N_6617,N_6388,N_6436);
and U6618 (N_6618,N_6403,N_6496);
xnor U6619 (N_6619,N_6471,N_6475);
xnor U6620 (N_6620,N_6489,N_6398);
nand U6621 (N_6621,N_6456,N_6473);
or U6622 (N_6622,N_6383,N_6411);
or U6623 (N_6623,N_6389,N_6429);
nand U6624 (N_6624,N_6381,N_6397);
xnor U6625 (N_6625,N_6529,N_6589);
or U6626 (N_6626,N_6548,N_6603);
nand U6627 (N_6627,N_6518,N_6597);
or U6628 (N_6628,N_6581,N_6604);
and U6629 (N_6629,N_6623,N_6577);
nand U6630 (N_6630,N_6504,N_6594);
or U6631 (N_6631,N_6533,N_6563);
nand U6632 (N_6632,N_6515,N_6556);
xnor U6633 (N_6633,N_6500,N_6510);
nand U6634 (N_6634,N_6585,N_6574);
nor U6635 (N_6635,N_6570,N_6580);
nor U6636 (N_6636,N_6517,N_6615);
and U6637 (N_6637,N_6506,N_6572);
nand U6638 (N_6638,N_6546,N_6535);
or U6639 (N_6639,N_6525,N_6593);
xor U6640 (N_6640,N_6607,N_6592);
xnor U6641 (N_6641,N_6598,N_6549);
xor U6642 (N_6642,N_6537,N_6606);
xor U6643 (N_6643,N_6599,N_6539);
or U6644 (N_6644,N_6505,N_6612);
nor U6645 (N_6645,N_6501,N_6600);
nand U6646 (N_6646,N_6555,N_6605);
nor U6647 (N_6647,N_6530,N_6565);
xnor U6648 (N_6648,N_6602,N_6516);
and U6649 (N_6649,N_6571,N_6553);
xnor U6650 (N_6650,N_6620,N_6512);
and U6651 (N_6651,N_6601,N_6568);
and U6652 (N_6652,N_6519,N_6559);
nor U6653 (N_6653,N_6511,N_6547);
xor U6654 (N_6654,N_6520,N_6619);
nand U6655 (N_6655,N_6590,N_6595);
nor U6656 (N_6656,N_6528,N_6586);
nand U6657 (N_6657,N_6610,N_6621);
xor U6658 (N_6658,N_6618,N_6608);
nand U6659 (N_6659,N_6526,N_6507);
and U6660 (N_6660,N_6567,N_6617);
or U6661 (N_6661,N_6521,N_6522);
and U6662 (N_6662,N_6575,N_6564);
or U6663 (N_6663,N_6588,N_6622);
or U6664 (N_6664,N_6558,N_6616);
or U6665 (N_6665,N_6536,N_6583);
and U6666 (N_6666,N_6545,N_6532);
or U6667 (N_6667,N_6569,N_6527);
and U6668 (N_6668,N_6609,N_6523);
and U6669 (N_6669,N_6503,N_6543);
xor U6670 (N_6670,N_6587,N_6578);
nor U6671 (N_6671,N_6566,N_6502);
nand U6672 (N_6672,N_6531,N_6613);
or U6673 (N_6673,N_6560,N_6557);
nand U6674 (N_6674,N_6544,N_6551);
and U6675 (N_6675,N_6534,N_6538);
nor U6676 (N_6676,N_6591,N_6552);
and U6677 (N_6677,N_6573,N_6562);
and U6678 (N_6678,N_6541,N_6596);
nand U6679 (N_6679,N_6508,N_6576);
and U6680 (N_6680,N_6542,N_6624);
xor U6681 (N_6681,N_6561,N_6513);
nand U6682 (N_6682,N_6554,N_6550);
or U6683 (N_6683,N_6509,N_6524);
nor U6684 (N_6684,N_6614,N_6579);
nor U6685 (N_6685,N_6611,N_6582);
or U6686 (N_6686,N_6540,N_6514);
xnor U6687 (N_6687,N_6584,N_6545);
nor U6688 (N_6688,N_6611,N_6560);
xnor U6689 (N_6689,N_6579,N_6568);
nor U6690 (N_6690,N_6515,N_6527);
and U6691 (N_6691,N_6553,N_6606);
nand U6692 (N_6692,N_6504,N_6596);
and U6693 (N_6693,N_6592,N_6530);
nand U6694 (N_6694,N_6503,N_6587);
or U6695 (N_6695,N_6624,N_6555);
or U6696 (N_6696,N_6586,N_6613);
and U6697 (N_6697,N_6560,N_6607);
and U6698 (N_6698,N_6517,N_6505);
nor U6699 (N_6699,N_6618,N_6534);
xor U6700 (N_6700,N_6520,N_6581);
nor U6701 (N_6701,N_6598,N_6532);
xnor U6702 (N_6702,N_6518,N_6553);
or U6703 (N_6703,N_6518,N_6555);
nor U6704 (N_6704,N_6501,N_6610);
nand U6705 (N_6705,N_6565,N_6578);
nand U6706 (N_6706,N_6587,N_6520);
nor U6707 (N_6707,N_6531,N_6512);
nor U6708 (N_6708,N_6563,N_6550);
nand U6709 (N_6709,N_6612,N_6618);
nand U6710 (N_6710,N_6502,N_6624);
or U6711 (N_6711,N_6519,N_6514);
or U6712 (N_6712,N_6581,N_6618);
nand U6713 (N_6713,N_6547,N_6512);
and U6714 (N_6714,N_6577,N_6585);
or U6715 (N_6715,N_6567,N_6523);
and U6716 (N_6716,N_6513,N_6618);
and U6717 (N_6717,N_6606,N_6597);
xor U6718 (N_6718,N_6503,N_6574);
or U6719 (N_6719,N_6539,N_6547);
or U6720 (N_6720,N_6600,N_6575);
or U6721 (N_6721,N_6573,N_6624);
nand U6722 (N_6722,N_6575,N_6551);
nor U6723 (N_6723,N_6603,N_6509);
xor U6724 (N_6724,N_6506,N_6534);
or U6725 (N_6725,N_6603,N_6516);
nor U6726 (N_6726,N_6558,N_6518);
nor U6727 (N_6727,N_6539,N_6505);
and U6728 (N_6728,N_6611,N_6586);
and U6729 (N_6729,N_6558,N_6606);
nand U6730 (N_6730,N_6559,N_6546);
or U6731 (N_6731,N_6620,N_6555);
or U6732 (N_6732,N_6588,N_6531);
and U6733 (N_6733,N_6566,N_6623);
or U6734 (N_6734,N_6578,N_6582);
xnor U6735 (N_6735,N_6609,N_6621);
and U6736 (N_6736,N_6512,N_6606);
or U6737 (N_6737,N_6507,N_6613);
nor U6738 (N_6738,N_6605,N_6548);
nand U6739 (N_6739,N_6595,N_6600);
or U6740 (N_6740,N_6577,N_6557);
xor U6741 (N_6741,N_6538,N_6585);
xor U6742 (N_6742,N_6587,N_6600);
and U6743 (N_6743,N_6585,N_6558);
nor U6744 (N_6744,N_6616,N_6517);
or U6745 (N_6745,N_6606,N_6508);
nor U6746 (N_6746,N_6517,N_6531);
xnor U6747 (N_6747,N_6528,N_6573);
nor U6748 (N_6748,N_6568,N_6586);
xnor U6749 (N_6749,N_6594,N_6571);
nand U6750 (N_6750,N_6641,N_6630);
and U6751 (N_6751,N_6686,N_6740);
or U6752 (N_6752,N_6644,N_6657);
and U6753 (N_6753,N_6748,N_6733);
and U6754 (N_6754,N_6711,N_6675);
and U6755 (N_6755,N_6636,N_6690);
or U6756 (N_6756,N_6685,N_6701);
or U6757 (N_6757,N_6672,N_6739);
nor U6758 (N_6758,N_6716,N_6745);
xnor U6759 (N_6759,N_6667,N_6735);
or U6760 (N_6760,N_6679,N_6628);
xor U6761 (N_6761,N_6741,N_6749);
and U6762 (N_6762,N_6687,N_6652);
and U6763 (N_6763,N_6696,N_6684);
nand U6764 (N_6764,N_6699,N_6646);
nand U6765 (N_6765,N_6702,N_6625);
and U6766 (N_6766,N_6736,N_6634);
or U6767 (N_6767,N_6724,N_6746);
or U6768 (N_6768,N_6719,N_6703);
nor U6769 (N_6769,N_6718,N_6656);
nor U6770 (N_6770,N_6632,N_6695);
nor U6771 (N_6771,N_6654,N_6665);
nand U6772 (N_6772,N_6638,N_6707);
and U6773 (N_6773,N_6659,N_6706);
or U6774 (N_6774,N_6631,N_6726);
xor U6775 (N_6775,N_6626,N_6712);
or U6776 (N_6776,N_6693,N_6629);
xor U6777 (N_6777,N_6710,N_6663);
and U6778 (N_6778,N_6671,N_6744);
xor U6779 (N_6779,N_6689,N_6678);
or U6780 (N_6780,N_6691,N_6677);
nand U6781 (N_6781,N_6698,N_6694);
nand U6782 (N_6782,N_6662,N_6727);
nor U6783 (N_6783,N_6633,N_6688);
or U6784 (N_6784,N_6715,N_6720);
or U6785 (N_6785,N_6729,N_6664);
xnor U6786 (N_6786,N_6673,N_6668);
nand U6787 (N_6787,N_6674,N_6647);
nand U6788 (N_6788,N_6692,N_6700);
nand U6789 (N_6789,N_6653,N_6639);
or U6790 (N_6790,N_6645,N_6637);
nand U6791 (N_6791,N_6730,N_6697);
nor U6792 (N_6792,N_6705,N_6721);
and U6793 (N_6793,N_6627,N_6722);
nor U6794 (N_6794,N_6643,N_6670);
nand U6795 (N_6795,N_6642,N_6723);
nand U6796 (N_6796,N_6635,N_6649);
or U6797 (N_6797,N_6640,N_6655);
nor U6798 (N_6798,N_6728,N_6704);
and U6799 (N_6799,N_6660,N_6683);
and U6800 (N_6800,N_6734,N_6658);
xnor U6801 (N_6801,N_6666,N_6725);
and U6802 (N_6802,N_6742,N_6713);
nor U6803 (N_6803,N_6717,N_6680);
nor U6804 (N_6804,N_6732,N_6650);
nor U6805 (N_6805,N_6648,N_6669);
or U6806 (N_6806,N_6651,N_6743);
and U6807 (N_6807,N_6676,N_6714);
xor U6808 (N_6808,N_6661,N_6747);
nor U6809 (N_6809,N_6709,N_6737);
xor U6810 (N_6810,N_6731,N_6681);
nor U6811 (N_6811,N_6682,N_6708);
nor U6812 (N_6812,N_6738,N_6720);
xnor U6813 (N_6813,N_6720,N_6702);
and U6814 (N_6814,N_6696,N_6703);
and U6815 (N_6815,N_6714,N_6626);
nor U6816 (N_6816,N_6686,N_6721);
nor U6817 (N_6817,N_6667,N_6645);
and U6818 (N_6818,N_6691,N_6649);
xnor U6819 (N_6819,N_6729,N_6698);
nor U6820 (N_6820,N_6691,N_6646);
nand U6821 (N_6821,N_6731,N_6640);
or U6822 (N_6822,N_6721,N_6729);
nor U6823 (N_6823,N_6734,N_6700);
xnor U6824 (N_6824,N_6692,N_6720);
nand U6825 (N_6825,N_6650,N_6635);
xor U6826 (N_6826,N_6728,N_6636);
nor U6827 (N_6827,N_6730,N_6628);
and U6828 (N_6828,N_6731,N_6661);
nor U6829 (N_6829,N_6744,N_6734);
or U6830 (N_6830,N_6660,N_6640);
nand U6831 (N_6831,N_6668,N_6730);
or U6832 (N_6832,N_6738,N_6734);
nor U6833 (N_6833,N_6727,N_6651);
xnor U6834 (N_6834,N_6652,N_6738);
nor U6835 (N_6835,N_6631,N_6693);
and U6836 (N_6836,N_6627,N_6665);
or U6837 (N_6837,N_6670,N_6709);
and U6838 (N_6838,N_6745,N_6673);
xor U6839 (N_6839,N_6728,N_6727);
or U6840 (N_6840,N_6659,N_6748);
or U6841 (N_6841,N_6641,N_6628);
and U6842 (N_6842,N_6642,N_6658);
nor U6843 (N_6843,N_6725,N_6652);
nand U6844 (N_6844,N_6705,N_6673);
nand U6845 (N_6845,N_6710,N_6707);
nor U6846 (N_6846,N_6684,N_6735);
xor U6847 (N_6847,N_6655,N_6712);
and U6848 (N_6848,N_6721,N_6719);
or U6849 (N_6849,N_6702,N_6684);
or U6850 (N_6850,N_6676,N_6638);
nor U6851 (N_6851,N_6655,N_6727);
or U6852 (N_6852,N_6700,N_6741);
xor U6853 (N_6853,N_6646,N_6643);
nor U6854 (N_6854,N_6721,N_6737);
and U6855 (N_6855,N_6706,N_6631);
and U6856 (N_6856,N_6687,N_6688);
and U6857 (N_6857,N_6653,N_6681);
nand U6858 (N_6858,N_6651,N_6627);
nor U6859 (N_6859,N_6658,N_6686);
xor U6860 (N_6860,N_6637,N_6725);
or U6861 (N_6861,N_6712,N_6651);
or U6862 (N_6862,N_6639,N_6729);
and U6863 (N_6863,N_6729,N_6736);
or U6864 (N_6864,N_6678,N_6679);
nor U6865 (N_6865,N_6726,N_6730);
or U6866 (N_6866,N_6697,N_6679);
nand U6867 (N_6867,N_6718,N_6706);
nand U6868 (N_6868,N_6747,N_6683);
nand U6869 (N_6869,N_6714,N_6685);
nand U6870 (N_6870,N_6694,N_6648);
or U6871 (N_6871,N_6678,N_6723);
nor U6872 (N_6872,N_6717,N_6666);
xor U6873 (N_6873,N_6632,N_6746);
nand U6874 (N_6874,N_6710,N_6638);
nor U6875 (N_6875,N_6854,N_6765);
and U6876 (N_6876,N_6817,N_6828);
or U6877 (N_6877,N_6849,N_6803);
xor U6878 (N_6878,N_6779,N_6750);
or U6879 (N_6879,N_6818,N_6841);
and U6880 (N_6880,N_6773,N_6850);
and U6881 (N_6881,N_6756,N_6822);
nor U6882 (N_6882,N_6859,N_6766);
xor U6883 (N_6883,N_6860,N_6867);
and U6884 (N_6884,N_6753,N_6870);
nor U6885 (N_6885,N_6783,N_6833);
or U6886 (N_6886,N_6769,N_6866);
nand U6887 (N_6887,N_6839,N_6838);
nor U6888 (N_6888,N_6791,N_6847);
and U6889 (N_6889,N_6865,N_6869);
and U6890 (N_6890,N_6805,N_6855);
or U6891 (N_6891,N_6794,N_6844);
and U6892 (N_6892,N_6806,N_6864);
nor U6893 (N_6893,N_6792,N_6785);
xor U6894 (N_6894,N_6758,N_6771);
and U6895 (N_6895,N_6772,N_6786);
nor U6896 (N_6896,N_6809,N_6760);
xnor U6897 (N_6897,N_6853,N_6781);
nand U6898 (N_6898,N_6762,N_6840);
nor U6899 (N_6899,N_6813,N_6775);
nor U6900 (N_6900,N_6825,N_6845);
xnor U6901 (N_6901,N_6842,N_6757);
or U6902 (N_6902,N_6861,N_6768);
nand U6903 (N_6903,N_6862,N_6836);
nor U6904 (N_6904,N_6800,N_6852);
nand U6905 (N_6905,N_6846,N_6872);
nor U6906 (N_6906,N_6777,N_6798);
and U6907 (N_6907,N_6812,N_6807);
nor U6908 (N_6908,N_6826,N_6797);
or U6909 (N_6909,N_6752,N_6767);
or U6910 (N_6910,N_6830,N_6814);
and U6911 (N_6911,N_6790,N_6751);
xor U6912 (N_6912,N_6823,N_6759);
nand U6913 (N_6913,N_6801,N_6843);
and U6914 (N_6914,N_6778,N_6804);
nand U6915 (N_6915,N_6782,N_6821);
nand U6916 (N_6916,N_6856,N_6784);
or U6917 (N_6917,N_6874,N_6787);
nor U6918 (N_6918,N_6763,N_6873);
nand U6919 (N_6919,N_6835,N_6811);
and U6920 (N_6920,N_6810,N_6776);
xnor U6921 (N_6921,N_6802,N_6851);
nand U6922 (N_6922,N_6868,N_6820);
or U6923 (N_6923,N_6755,N_6774);
nand U6924 (N_6924,N_6754,N_6834);
nand U6925 (N_6925,N_6789,N_6796);
xnor U6926 (N_6926,N_6764,N_6871);
and U6927 (N_6927,N_6831,N_6780);
nand U6928 (N_6928,N_6858,N_6815);
and U6929 (N_6929,N_6863,N_6827);
xor U6930 (N_6930,N_6795,N_6824);
xnor U6931 (N_6931,N_6837,N_6819);
xnor U6932 (N_6932,N_6770,N_6808);
and U6933 (N_6933,N_6788,N_6857);
or U6934 (N_6934,N_6793,N_6761);
nand U6935 (N_6935,N_6799,N_6816);
and U6936 (N_6936,N_6832,N_6848);
xnor U6937 (N_6937,N_6829,N_6858);
nor U6938 (N_6938,N_6833,N_6867);
xnor U6939 (N_6939,N_6758,N_6750);
or U6940 (N_6940,N_6853,N_6807);
and U6941 (N_6941,N_6868,N_6782);
nor U6942 (N_6942,N_6861,N_6752);
nor U6943 (N_6943,N_6862,N_6774);
xnor U6944 (N_6944,N_6839,N_6843);
nand U6945 (N_6945,N_6811,N_6858);
or U6946 (N_6946,N_6821,N_6842);
and U6947 (N_6947,N_6805,N_6799);
nor U6948 (N_6948,N_6755,N_6804);
nor U6949 (N_6949,N_6807,N_6796);
xor U6950 (N_6950,N_6791,N_6813);
or U6951 (N_6951,N_6853,N_6788);
xor U6952 (N_6952,N_6860,N_6812);
or U6953 (N_6953,N_6798,N_6787);
nand U6954 (N_6954,N_6797,N_6861);
nor U6955 (N_6955,N_6794,N_6850);
xor U6956 (N_6956,N_6761,N_6873);
xnor U6957 (N_6957,N_6766,N_6765);
or U6958 (N_6958,N_6818,N_6777);
nand U6959 (N_6959,N_6763,N_6791);
xnor U6960 (N_6960,N_6846,N_6843);
nand U6961 (N_6961,N_6763,N_6853);
nor U6962 (N_6962,N_6811,N_6859);
xnor U6963 (N_6963,N_6827,N_6781);
xnor U6964 (N_6964,N_6826,N_6763);
nor U6965 (N_6965,N_6795,N_6761);
xnor U6966 (N_6966,N_6803,N_6858);
nand U6967 (N_6967,N_6830,N_6823);
xnor U6968 (N_6968,N_6763,N_6799);
nand U6969 (N_6969,N_6857,N_6859);
or U6970 (N_6970,N_6801,N_6769);
nand U6971 (N_6971,N_6823,N_6772);
xnor U6972 (N_6972,N_6841,N_6763);
and U6973 (N_6973,N_6767,N_6758);
nor U6974 (N_6974,N_6838,N_6797);
nor U6975 (N_6975,N_6761,N_6778);
nor U6976 (N_6976,N_6802,N_6817);
nand U6977 (N_6977,N_6776,N_6766);
nor U6978 (N_6978,N_6862,N_6849);
or U6979 (N_6979,N_6860,N_6792);
xnor U6980 (N_6980,N_6757,N_6775);
or U6981 (N_6981,N_6752,N_6788);
and U6982 (N_6982,N_6789,N_6780);
xor U6983 (N_6983,N_6826,N_6872);
nor U6984 (N_6984,N_6847,N_6788);
xor U6985 (N_6985,N_6803,N_6847);
or U6986 (N_6986,N_6828,N_6776);
nand U6987 (N_6987,N_6823,N_6828);
nand U6988 (N_6988,N_6853,N_6769);
nor U6989 (N_6989,N_6848,N_6755);
and U6990 (N_6990,N_6865,N_6868);
xor U6991 (N_6991,N_6818,N_6851);
nor U6992 (N_6992,N_6870,N_6848);
nor U6993 (N_6993,N_6795,N_6857);
nor U6994 (N_6994,N_6787,N_6781);
nor U6995 (N_6995,N_6847,N_6850);
nand U6996 (N_6996,N_6780,N_6870);
or U6997 (N_6997,N_6764,N_6807);
nor U6998 (N_6998,N_6871,N_6858);
and U6999 (N_6999,N_6850,N_6862);
or U7000 (N_7000,N_6887,N_6970);
nand U7001 (N_7001,N_6955,N_6953);
nand U7002 (N_7002,N_6975,N_6910);
nand U7003 (N_7003,N_6878,N_6945);
or U7004 (N_7004,N_6974,N_6891);
and U7005 (N_7005,N_6981,N_6909);
and U7006 (N_7006,N_6886,N_6983);
nand U7007 (N_7007,N_6932,N_6935);
or U7008 (N_7008,N_6913,N_6994);
or U7009 (N_7009,N_6950,N_6982);
nand U7010 (N_7010,N_6942,N_6962);
nand U7011 (N_7011,N_6918,N_6896);
xor U7012 (N_7012,N_6991,N_6968);
nor U7013 (N_7013,N_6965,N_6890);
nand U7014 (N_7014,N_6972,N_6897);
nor U7015 (N_7015,N_6901,N_6904);
nor U7016 (N_7016,N_6907,N_6908);
and U7017 (N_7017,N_6951,N_6927);
xnor U7018 (N_7018,N_6941,N_6880);
nor U7019 (N_7019,N_6936,N_6917);
and U7020 (N_7020,N_6928,N_6961);
nor U7021 (N_7021,N_6999,N_6979);
xor U7022 (N_7022,N_6929,N_6906);
xor U7023 (N_7023,N_6894,N_6933);
or U7024 (N_7024,N_6985,N_6895);
nand U7025 (N_7025,N_6958,N_6947);
xor U7026 (N_7026,N_6960,N_6969);
nand U7027 (N_7027,N_6898,N_6875);
xor U7028 (N_7028,N_6892,N_6877);
nor U7029 (N_7029,N_6912,N_6915);
or U7030 (N_7030,N_6964,N_6989);
nor U7031 (N_7031,N_6940,N_6923);
or U7032 (N_7032,N_6924,N_6967);
xnor U7033 (N_7033,N_6971,N_6879);
and U7034 (N_7034,N_6963,N_6977);
nand U7035 (N_7035,N_6956,N_6899);
or U7036 (N_7036,N_6926,N_6902);
xor U7037 (N_7037,N_6993,N_6934);
nand U7038 (N_7038,N_6937,N_6905);
and U7039 (N_7039,N_6944,N_6914);
xnor U7040 (N_7040,N_6996,N_6986);
nor U7041 (N_7041,N_6952,N_6921);
nand U7042 (N_7042,N_6916,N_6882);
nand U7043 (N_7043,N_6925,N_6980);
xor U7044 (N_7044,N_6998,N_6903);
or U7045 (N_7045,N_6943,N_6946);
nand U7046 (N_7046,N_6954,N_6922);
or U7047 (N_7047,N_6997,N_6995);
and U7048 (N_7048,N_6939,N_6919);
nand U7049 (N_7049,N_6888,N_6990);
nand U7050 (N_7050,N_6893,N_6966);
nand U7051 (N_7051,N_6930,N_6876);
and U7052 (N_7052,N_6911,N_6959);
or U7053 (N_7053,N_6992,N_6984);
xnor U7054 (N_7054,N_6885,N_6987);
xnor U7055 (N_7055,N_6988,N_6948);
and U7056 (N_7056,N_6938,N_6881);
or U7057 (N_7057,N_6978,N_6931);
nand U7058 (N_7058,N_6973,N_6883);
xnor U7059 (N_7059,N_6889,N_6920);
and U7060 (N_7060,N_6884,N_6957);
xnor U7061 (N_7061,N_6976,N_6900);
or U7062 (N_7062,N_6949,N_6965);
nor U7063 (N_7063,N_6926,N_6877);
and U7064 (N_7064,N_6931,N_6901);
nand U7065 (N_7065,N_6970,N_6990);
and U7066 (N_7066,N_6963,N_6879);
or U7067 (N_7067,N_6895,N_6992);
and U7068 (N_7068,N_6939,N_6937);
nand U7069 (N_7069,N_6953,N_6967);
xnor U7070 (N_7070,N_6929,N_6931);
xor U7071 (N_7071,N_6904,N_6916);
and U7072 (N_7072,N_6897,N_6978);
xor U7073 (N_7073,N_6996,N_6928);
xnor U7074 (N_7074,N_6973,N_6914);
or U7075 (N_7075,N_6997,N_6981);
xnor U7076 (N_7076,N_6919,N_6915);
nand U7077 (N_7077,N_6937,N_6914);
xnor U7078 (N_7078,N_6923,N_6898);
nor U7079 (N_7079,N_6995,N_6945);
and U7080 (N_7080,N_6922,N_6944);
or U7081 (N_7081,N_6985,N_6947);
xnor U7082 (N_7082,N_6919,N_6966);
xor U7083 (N_7083,N_6961,N_6885);
nor U7084 (N_7084,N_6886,N_6925);
or U7085 (N_7085,N_6977,N_6970);
nand U7086 (N_7086,N_6892,N_6930);
or U7087 (N_7087,N_6896,N_6887);
xnor U7088 (N_7088,N_6920,N_6971);
nand U7089 (N_7089,N_6916,N_6883);
nand U7090 (N_7090,N_6896,N_6987);
nor U7091 (N_7091,N_6890,N_6982);
nor U7092 (N_7092,N_6909,N_6892);
nand U7093 (N_7093,N_6892,N_6961);
or U7094 (N_7094,N_6912,N_6955);
and U7095 (N_7095,N_6920,N_6978);
or U7096 (N_7096,N_6915,N_6991);
xor U7097 (N_7097,N_6943,N_6931);
or U7098 (N_7098,N_6933,N_6937);
nor U7099 (N_7099,N_6949,N_6881);
or U7100 (N_7100,N_6932,N_6902);
or U7101 (N_7101,N_6890,N_6975);
xor U7102 (N_7102,N_6915,N_6954);
and U7103 (N_7103,N_6902,N_6918);
nor U7104 (N_7104,N_6979,N_6940);
xnor U7105 (N_7105,N_6884,N_6910);
or U7106 (N_7106,N_6902,N_6933);
or U7107 (N_7107,N_6956,N_6993);
xnor U7108 (N_7108,N_6892,N_6941);
and U7109 (N_7109,N_6896,N_6968);
xor U7110 (N_7110,N_6961,N_6972);
xor U7111 (N_7111,N_6980,N_6972);
and U7112 (N_7112,N_6883,N_6988);
or U7113 (N_7113,N_6886,N_6898);
and U7114 (N_7114,N_6907,N_6897);
nand U7115 (N_7115,N_6980,N_6912);
or U7116 (N_7116,N_6906,N_6898);
and U7117 (N_7117,N_6977,N_6964);
and U7118 (N_7118,N_6890,N_6952);
and U7119 (N_7119,N_6984,N_6916);
nand U7120 (N_7120,N_6892,N_6975);
nand U7121 (N_7121,N_6927,N_6908);
and U7122 (N_7122,N_6894,N_6982);
nand U7123 (N_7123,N_6971,N_6905);
nand U7124 (N_7124,N_6953,N_6927);
nand U7125 (N_7125,N_7056,N_7059);
and U7126 (N_7126,N_7016,N_7009);
or U7127 (N_7127,N_7001,N_7003);
nand U7128 (N_7128,N_7031,N_7034);
xor U7129 (N_7129,N_7044,N_7049);
or U7130 (N_7130,N_7086,N_7105);
nor U7131 (N_7131,N_7068,N_7089);
or U7132 (N_7132,N_7000,N_7083);
and U7133 (N_7133,N_7052,N_7117);
and U7134 (N_7134,N_7028,N_7048);
nand U7135 (N_7135,N_7027,N_7074);
or U7136 (N_7136,N_7093,N_7085);
nand U7137 (N_7137,N_7110,N_7022);
nor U7138 (N_7138,N_7007,N_7036);
and U7139 (N_7139,N_7047,N_7039);
xor U7140 (N_7140,N_7062,N_7106);
or U7141 (N_7141,N_7051,N_7077);
nand U7142 (N_7142,N_7090,N_7116);
nor U7143 (N_7143,N_7020,N_7054);
and U7144 (N_7144,N_7094,N_7072);
nand U7145 (N_7145,N_7014,N_7121);
and U7146 (N_7146,N_7026,N_7021);
xnor U7147 (N_7147,N_7099,N_7008);
xnor U7148 (N_7148,N_7108,N_7046);
nor U7149 (N_7149,N_7064,N_7053);
or U7150 (N_7150,N_7019,N_7012);
or U7151 (N_7151,N_7010,N_7073);
nor U7152 (N_7152,N_7042,N_7100);
and U7153 (N_7153,N_7033,N_7002);
xnor U7154 (N_7154,N_7004,N_7115);
xnor U7155 (N_7155,N_7124,N_7055);
or U7156 (N_7156,N_7113,N_7104);
nand U7157 (N_7157,N_7017,N_7030);
xor U7158 (N_7158,N_7025,N_7095);
nand U7159 (N_7159,N_7066,N_7102);
nand U7160 (N_7160,N_7013,N_7081);
and U7161 (N_7161,N_7037,N_7069);
xor U7162 (N_7162,N_7123,N_7006);
or U7163 (N_7163,N_7065,N_7096);
xor U7164 (N_7164,N_7067,N_7101);
nand U7165 (N_7165,N_7088,N_7005);
or U7166 (N_7166,N_7071,N_7114);
nand U7167 (N_7167,N_7103,N_7078);
and U7168 (N_7168,N_7058,N_7061);
nor U7169 (N_7169,N_7018,N_7091);
nand U7170 (N_7170,N_7079,N_7038);
nor U7171 (N_7171,N_7119,N_7092);
or U7172 (N_7172,N_7111,N_7075);
and U7173 (N_7173,N_7024,N_7087);
or U7174 (N_7174,N_7063,N_7070);
and U7175 (N_7175,N_7023,N_7029);
or U7176 (N_7176,N_7050,N_7109);
or U7177 (N_7177,N_7057,N_7107);
nand U7178 (N_7178,N_7041,N_7035);
nand U7179 (N_7179,N_7060,N_7118);
and U7180 (N_7180,N_7120,N_7082);
xnor U7181 (N_7181,N_7080,N_7097);
or U7182 (N_7182,N_7011,N_7122);
nand U7183 (N_7183,N_7043,N_7112);
and U7184 (N_7184,N_7045,N_7084);
or U7185 (N_7185,N_7015,N_7040);
or U7186 (N_7186,N_7076,N_7098);
and U7187 (N_7187,N_7032,N_7107);
and U7188 (N_7188,N_7024,N_7007);
nor U7189 (N_7189,N_7104,N_7059);
and U7190 (N_7190,N_7007,N_7078);
nand U7191 (N_7191,N_7034,N_7106);
or U7192 (N_7192,N_7082,N_7061);
nor U7193 (N_7193,N_7089,N_7077);
nor U7194 (N_7194,N_7010,N_7112);
xor U7195 (N_7195,N_7061,N_7014);
or U7196 (N_7196,N_7035,N_7055);
nand U7197 (N_7197,N_7076,N_7099);
nor U7198 (N_7198,N_7034,N_7062);
or U7199 (N_7199,N_7038,N_7040);
nor U7200 (N_7200,N_7033,N_7022);
or U7201 (N_7201,N_7115,N_7062);
xor U7202 (N_7202,N_7017,N_7011);
xor U7203 (N_7203,N_7007,N_7115);
xnor U7204 (N_7204,N_7039,N_7101);
and U7205 (N_7205,N_7046,N_7115);
xnor U7206 (N_7206,N_7000,N_7035);
and U7207 (N_7207,N_7080,N_7102);
and U7208 (N_7208,N_7054,N_7012);
xnor U7209 (N_7209,N_7117,N_7005);
nor U7210 (N_7210,N_7028,N_7036);
and U7211 (N_7211,N_7019,N_7091);
and U7212 (N_7212,N_7004,N_7050);
and U7213 (N_7213,N_7008,N_7096);
or U7214 (N_7214,N_7019,N_7041);
nor U7215 (N_7215,N_7096,N_7041);
nand U7216 (N_7216,N_7004,N_7121);
nor U7217 (N_7217,N_7047,N_7063);
nand U7218 (N_7218,N_7063,N_7064);
xor U7219 (N_7219,N_7045,N_7076);
or U7220 (N_7220,N_7012,N_7101);
nand U7221 (N_7221,N_7039,N_7061);
nand U7222 (N_7222,N_7016,N_7093);
or U7223 (N_7223,N_7021,N_7096);
or U7224 (N_7224,N_7006,N_7057);
nor U7225 (N_7225,N_7049,N_7081);
xor U7226 (N_7226,N_7020,N_7122);
and U7227 (N_7227,N_7106,N_7001);
nand U7228 (N_7228,N_7039,N_7037);
or U7229 (N_7229,N_7094,N_7040);
nor U7230 (N_7230,N_7080,N_7071);
nor U7231 (N_7231,N_7117,N_7023);
and U7232 (N_7232,N_7022,N_7122);
and U7233 (N_7233,N_7046,N_7040);
and U7234 (N_7234,N_7006,N_7068);
or U7235 (N_7235,N_7122,N_7065);
nand U7236 (N_7236,N_7048,N_7026);
and U7237 (N_7237,N_7063,N_7059);
or U7238 (N_7238,N_7074,N_7099);
and U7239 (N_7239,N_7119,N_7021);
xor U7240 (N_7240,N_7117,N_7066);
nor U7241 (N_7241,N_7088,N_7045);
xnor U7242 (N_7242,N_7044,N_7112);
xnor U7243 (N_7243,N_7030,N_7008);
or U7244 (N_7244,N_7066,N_7032);
nor U7245 (N_7245,N_7017,N_7054);
or U7246 (N_7246,N_7035,N_7117);
and U7247 (N_7247,N_7005,N_7012);
xnor U7248 (N_7248,N_7079,N_7107);
nor U7249 (N_7249,N_7071,N_7112);
xor U7250 (N_7250,N_7248,N_7222);
xor U7251 (N_7251,N_7164,N_7189);
or U7252 (N_7252,N_7132,N_7231);
xnor U7253 (N_7253,N_7171,N_7249);
or U7254 (N_7254,N_7142,N_7191);
xnor U7255 (N_7255,N_7243,N_7161);
nand U7256 (N_7256,N_7160,N_7175);
nand U7257 (N_7257,N_7199,N_7190);
nor U7258 (N_7258,N_7170,N_7185);
or U7259 (N_7259,N_7215,N_7207);
xnor U7260 (N_7260,N_7219,N_7147);
xnor U7261 (N_7261,N_7157,N_7182);
or U7262 (N_7262,N_7172,N_7127);
nand U7263 (N_7263,N_7224,N_7174);
and U7264 (N_7264,N_7134,N_7146);
nand U7265 (N_7265,N_7208,N_7247);
xor U7266 (N_7266,N_7201,N_7144);
nor U7267 (N_7267,N_7131,N_7230);
xnor U7268 (N_7268,N_7218,N_7209);
nor U7269 (N_7269,N_7244,N_7139);
or U7270 (N_7270,N_7153,N_7188);
xnor U7271 (N_7271,N_7204,N_7177);
nand U7272 (N_7272,N_7141,N_7135);
nor U7273 (N_7273,N_7228,N_7136);
and U7274 (N_7274,N_7206,N_7179);
xnor U7275 (N_7275,N_7221,N_7167);
nand U7276 (N_7276,N_7126,N_7125);
or U7277 (N_7277,N_7168,N_7194);
or U7278 (N_7278,N_7183,N_7233);
nor U7279 (N_7279,N_7166,N_7220);
and U7280 (N_7280,N_7216,N_7187);
or U7281 (N_7281,N_7178,N_7212);
nand U7282 (N_7282,N_7181,N_7197);
or U7283 (N_7283,N_7137,N_7225);
nor U7284 (N_7284,N_7217,N_7202);
nor U7285 (N_7285,N_7128,N_7173);
xor U7286 (N_7286,N_7234,N_7223);
and U7287 (N_7287,N_7198,N_7129);
nand U7288 (N_7288,N_7195,N_7239);
xor U7289 (N_7289,N_7158,N_7232);
nand U7290 (N_7290,N_7162,N_7138);
nor U7291 (N_7291,N_7133,N_7169);
or U7292 (N_7292,N_7163,N_7238);
or U7293 (N_7293,N_7246,N_7203);
nor U7294 (N_7294,N_7165,N_7242);
or U7295 (N_7295,N_7130,N_7155);
and U7296 (N_7296,N_7150,N_7152);
nand U7297 (N_7297,N_7235,N_7236);
xnor U7298 (N_7298,N_7240,N_7193);
nand U7299 (N_7299,N_7205,N_7211);
or U7300 (N_7300,N_7159,N_7180);
and U7301 (N_7301,N_7241,N_7176);
xnor U7302 (N_7302,N_7186,N_7210);
xnor U7303 (N_7303,N_7226,N_7184);
and U7304 (N_7304,N_7140,N_7229);
nand U7305 (N_7305,N_7151,N_7237);
xor U7306 (N_7306,N_7192,N_7227);
or U7307 (N_7307,N_7149,N_7200);
or U7308 (N_7308,N_7214,N_7145);
or U7309 (N_7309,N_7196,N_7156);
and U7310 (N_7310,N_7213,N_7148);
nand U7311 (N_7311,N_7245,N_7154);
nand U7312 (N_7312,N_7143,N_7172);
xnor U7313 (N_7313,N_7197,N_7248);
xnor U7314 (N_7314,N_7202,N_7144);
xnor U7315 (N_7315,N_7199,N_7189);
nor U7316 (N_7316,N_7126,N_7130);
nor U7317 (N_7317,N_7179,N_7172);
xor U7318 (N_7318,N_7247,N_7190);
xor U7319 (N_7319,N_7205,N_7206);
nor U7320 (N_7320,N_7229,N_7197);
and U7321 (N_7321,N_7245,N_7230);
or U7322 (N_7322,N_7242,N_7243);
xnor U7323 (N_7323,N_7198,N_7242);
or U7324 (N_7324,N_7184,N_7225);
or U7325 (N_7325,N_7188,N_7136);
nor U7326 (N_7326,N_7181,N_7143);
and U7327 (N_7327,N_7172,N_7169);
nand U7328 (N_7328,N_7242,N_7152);
nand U7329 (N_7329,N_7226,N_7175);
xor U7330 (N_7330,N_7178,N_7214);
and U7331 (N_7331,N_7246,N_7159);
and U7332 (N_7332,N_7138,N_7148);
or U7333 (N_7333,N_7128,N_7183);
xnor U7334 (N_7334,N_7211,N_7152);
nand U7335 (N_7335,N_7228,N_7249);
or U7336 (N_7336,N_7234,N_7184);
and U7337 (N_7337,N_7212,N_7161);
and U7338 (N_7338,N_7134,N_7213);
or U7339 (N_7339,N_7204,N_7229);
or U7340 (N_7340,N_7153,N_7198);
and U7341 (N_7341,N_7228,N_7181);
or U7342 (N_7342,N_7226,N_7247);
xnor U7343 (N_7343,N_7233,N_7175);
and U7344 (N_7344,N_7139,N_7192);
nor U7345 (N_7345,N_7167,N_7186);
nor U7346 (N_7346,N_7140,N_7162);
nand U7347 (N_7347,N_7238,N_7223);
nor U7348 (N_7348,N_7131,N_7185);
or U7349 (N_7349,N_7129,N_7244);
or U7350 (N_7350,N_7241,N_7133);
nand U7351 (N_7351,N_7159,N_7234);
or U7352 (N_7352,N_7167,N_7197);
nor U7353 (N_7353,N_7171,N_7240);
nor U7354 (N_7354,N_7241,N_7243);
nand U7355 (N_7355,N_7194,N_7172);
nor U7356 (N_7356,N_7168,N_7203);
nor U7357 (N_7357,N_7185,N_7220);
nand U7358 (N_7358,N_7222,N_7139);
xor U7359 (N_7359,N_7138,N_7146);
nor U7360 (N_7360,N_7129,N_7205);
xor U7361 (N_7361,N_7145,N_7131);
or U7362 (N_7362,N_7190,N_7159);
nor U7363 (N_7363,N_7222,N_7242);
or U7364 (N_7364,N_7205,N_7125);
and U7365 (N_7365,N_7173,N_7160);
nor U7366 (N_7366,N_7125,N_7136);
nor U7367 (N_7367,N_7155,N_7162);
xnor U7368 (N_7368,N_7154,N_7181);
or U7369 (N_7369,N_7138,N_7125);
and U7370 (N_7370,N_7184,N_7201);
xnor U7371 (N_7371,N_7180,N_7129);
or U7372 (N_7372,N_7167,N_7157);
nor U7373 (N_7373,N_7200,N_7188);
nor U7374 (N_7374,N_7218,N_7133);
and U7375 (N_7375,N_7280,N_7343);
nand U7376 (N_7376,N_7359,N_7301);
nand U7377 (N_7377,N_7335,N_7320);
and U7378 (N_7378,N_7300,N_7288);
or U7379 (N_7379,N_7332,N_7291);
and U7380 (N_7380,N_7303,N_7258);
nand U7381 (N_7381,N_7261,N_7340);
xnor U7382 (N_7382,N_7355,N_7294);
nor U7383 (N_7383,N_7313,N_7341);
and U7384 (N_7384,N_7366,N_7297);
nand U7385 (N_7385,N_7350,N_7357);
and U7386 (N_7386,N_7283,N_7268);
nor U7387 (N_7387,N_7356,N_7310);
and U7388 (N_7388,N_7339,N_7323);
or U7389 (N_7389,N_7374,N_7277);
nor U7390 (N_7390,N_7269,N_7278);
and U7391 (N_7391,N_7284,N_7317);
or U7392 (N_7392,N_7290,N_7270);
and U7393 (N_7393,N_7309,N_7315);
nand U7394 (N_7394,N_7327,N_7305);
nor U7395 (N_7395,N_7252,N_7279);
nor U7396 (N_7396,N_7285,N_7308);
or U7397 (N_7397,N_7292,N_7336);
and U7398 (N_7398,N_7250,N_7259);
nor U7399 (N_7399,N_7299,N_7345);
xnor U7400 (N_7400,N_7267,N_7364);
nand U7401 (N_7401,N_7334,N_7253);
and U7402 (N_7402,N_7266,N_7352);
and U7403 (N_7403,N_7321,N_7371);
nand U7404 (N_7404,N_7351,N_7368);
and U7405 (N_7405,N_7281,N_7337);
and U7406 (N_7406,N_7295,N_7342);
nor U7407 (N_7407,N_7331,N_7326);
xor U7408 (N_7408,N_7346,N_7263);
xnor U7409 (N_7409,N_7318,N_7264);
nor U7410 (N_7410,N_7276,N_7272);
and U7411 (N_7411,N_7286,N_7256);
xnor U7412 (N_7412,N_7365,N_7372);
xor U7413 (N_7413,N_7348,N_7370);
and U7414 (N_7414,N_7293,N_7373);
nand U7415 (N_7415,N_7306,N_7273);
nand U7416 (N_7416,N_7353,N_7265);
nor U7417 (N_7417,N_7330,N_7262);
and U7418 (N_7418,N_7324,N_7328);
xnor U7419 (N_7419,N_7255,N_7333);
nand U7420 (N_7420,N_7338,N_7287);
nand U7421 (N_7421,N_7251,N_7329);
nand U7422 (N_7422,N_7296,N_7361);
nand U7423 (N_7423,N_7260,N_7275);
nand U7424 (N_7424,N_7358,N_7316);
nand U7425 (N_7425,N_7271,N_7347);
nand U7426 (N_7426,N_7312,N_7367);
and U7427 (N_7427,N_7349,N_7298);
xnor U7428 (N_7428,N_7362,N_7257);
nand U7429 (N_7429,N_7319,N_7369);
and U7430 (N_7430,N_7304,N_7360);
xor U7431 (N_7431,N_7302,N_7325);
nand U7432 (N_7432,N_7363,N_7274);
and U7433 (N_7433,N_7322,N_7282);
or U7434 (N_7434,N_7254,N_7314);
or U7435 (N_7435,N_7344,N_7307);
nand U7436 (N_7436,N_7311,N_7354);
nor U7437 (N_7437,N_7289,N_7346);
or U7438 (N_7438,N_7301,N_7313);
nand U7439 (N_7439,N_7307,N_7353);
and U7440 (N_7440,N_7317,N_7323);
nor U7441 (N_7441,N_7310,N_7323);
nand U7442 (N_7442,N_7286,N_7327);
xnor U7443 (N_7443,N_7354,N_7358);
or U7444 (N_7444,N_7309,N_7290);
xnor U7445 (N_7445,N_7366,N_7360);
and U7446 (N_7446,N_7281,N_7269);
xnor U7447 (N_7447,N_7277,N_7267);
and U7448 (N_7448,N_7292,N_7256);
xor U7449 (N_7449,N_7306,N_7253);
xor U7450 (N_7450,N_7343,N_7349);
nand U7451 (N_7451,N_7335,N_7299);
nor U7452 (N_7452,N_7310,N_7301);
nand U7453 (N_7453,N_7261,N_7312);
nor U7454 (N_7454,N_7338,N_7268);
or U7455 (N_7455,N_7307,N_7366);
and U7456 (N_7456,N_7267,N_7320);
or U7457 (N_7457,N_7297,N_7264);
nor U7458 (N_7458,N_7351,N_7270);
nor U7459 (N_7459,N_7310,N_7348);
nor U7460 (N_7460,N_7333,N_7360);
nor U7461 (N_7461,N_7346,N_7276);
or U7462 (N_7462,N_7300,N_7276);
and U7463 (N_7463,N_7273,N_7330);
xor U7464 (N_7464,N_7338,N_7288);
or U7465 (N_7465,N_7312,N_7307);
and U7466 (N_7466,N_7268,N_7292);
xnor U7467 (N_7467,N_7286,N_7325);
nand U7468 (N_7468,N_7371,N_7303);
nor U7469 (N_7469,N_7274,N_7272);
and U7470 (N_7470,N_7370,N_7359);
nand U7471 (N_7471,N_7291,N_7260);
nand U7472 (N_7472,N_7268,N_7330);
nor U7473 (N_7473,N_7370,N_7360);
xnor U7474 (N_7474,N_7263,N_7286);
and U7475 (N_7475,N_7279,N_7349);
nor U7476 (N_7476,N_7310,N_7364);
or U7477 (N_7477,N_7309,N_7359);
or U7478 (N_7478,N_7260,N_7366);
nor U7479 (N_7479,N_7299,N_7358);
xnor U7480 (N_7480,N_7352,N_7326);
nor U7481 (N_7481,N_7347,N_7316);
xnor U7482 (N_7482,N_7324,N_7305);
or U7483 (N_7483,N_7271,N_7313);
nor U7484 (N_7484,N_7348,N_7293);
nor U7485 (N_7485,N_7347,N_7315);
or U7486 (N_7486,N_7266,N_7254);
and U7487 (N_7487,N_7320,N_7354);
nand U7488 (N_7488,N_7259,N_7334);
nor U7489 (N_7489,N_7268,N_7253);
nor U7490 (N_7490,N_7355,N_7318);
and U7491 (N_7491,N_7335,N_7357);
nand U7492 (N_7492,N_7359,N_7305);
nand U7493 (N_7493,N_7335,N_7374);
nand U7494 (N_7494,N_7277,N_7335);
and U7495 (N_7495,N_7343,N_7309);
nand U7496 (N_7496,N_7369,N_7361);
nand U7497 (N_7497,N_7342,N_7354);
xnor U7498 (N_7498,N_7270,N_7341);
and U7499 (N_7499,N_7320,N_7319);
or U7500 (N_7500,N_7422,N_7390);
and U7501 (N_7501,N_7380,N_7404);
and U7502 (N_7502,N_7385,N_7439);
nand U7503 (N_7503,N_7387,N_7396);
and U7504 (N_7504,N_7400,N_7491);
xor U7505 (N_7505,N_7457,N_7458);
nor U7506 (N_7506,N_7436,N_7379);
and U7507 (N_7507,N_7426,N_7493);
nor U7508 (N_7508,N_7450,N_7402);
and U7509 (N_7509,N_7453,N_7437);
or U7510 (N_7510,N_7466,N_7412);
xor U7511 (N_7511,N_7376,N_7494);
or U7512 (N_7512,N_7451,N_7469);
nor U7513 (N_7513,N_7428,N_7397);
nand U7514 (N_7514,N_7405,N_7415);
and U7515 (N_7515,N_7394,N_7395);
nor U7516 (N_7516,N_7375,N_7401);
nand U7517 (N_7517,N_7483,N_7485);
and U7518 (N_7518,N_7406,N_7459);
nor U7519 (N_7519,N_7496,N_7393);
xor U7520 (N_7520,N_7490,N_7416);
xor U7521 (N_7521,N_7381,N_7431);
or U7522 (N_7522,N_7468,N_7389);
and U7523 (N_7523,N_7482,N_7448);
nand U7524 (N_7524,N_7471,N_7445);
xor U7525 (N_7525,N_7425,N_7498);
and U7526 (N_7526,N_7441,N_7408);
nor U7527 (N_7527,N_7444,N_7424);
nor U7528 (N_7528,N_7454,N_7432);
and U7529 (N_7529,N_7442,N_7449);
nand U7530 (N_7530,N_7465,N_7446);
nor U7531 (N_7531,N_7492,N_7481);
nand U7532 (N_7532,N_7480,N_7399);
or U7533 (N_7533,N_7430,N_7418);
nand U7534 (N_7534,N_7391,N_7377);
nor U7535 (N_7535,N_7479,N_7433);
nand U7536 (N_7536,N_7427,N_7487);
nor U7537 (N_7537,N_7420,N_7435);
or U7538 (N_7538,N_7411,N_7499);
nand U7539 (N_7539,N_7434,N_7409);
or U7540 (N_7540,N_7407,N_7478);
nand U7541 (N_7541,N_7475,N_7382);
nor U7542 (N_7542,N_7440,N_7474);
xor U7543 (N_7543,N_7472,N_7477);
and U7544 (N_7544,N_7388,N_7410);
nor U7545 (N_7545,N_7460,N_7455);
and U7546 (N_7546,N_7429,N_7476);
nor U7547 (N_7547,N_7419,N_7421);
nand U7548 (N_7548,N_7414,N_7417);
nor U7549 (N_7549,N_7452,N_7464);
nor U7550 (N_7550,N_7470,N_7462);
nand U7551 (N_7551,N_7378,N_7392);
xnor U7552 (N_7552,N_7456,N_7484);
and U7553 (N_7553,N_7489,N_7403);
or U7554 (N_7554,N_7486,N_7447);
xnor U7555 (N_7555,N_7473,N_7461);
nor U7556 (N_7556,N_7495,N_7384);
and U7557 (N_7557,N_7497,N_7413);
and U7558 (N_7558,N_7443,N_7467);
xor U7559 (N_7559,N_7438,N_7488);
nand U7560 (N_7560,N_7398,N_7383);
nor U7561 (N_7561,N_7386,N_7463);
xnor U7562 (N_7562,N_7423,N_7380);
xnor U7563 (N_7563,N_7442,N_7421);
xnor U7564 (N_7564,N_7451,N_7418);
xor U7565 (N_7565,N_7421,N_7445);
and U7566 (N_7566,N_7495,N_7447);
xor U7567 (N_7567,N_7414,N_7399);
or U7568 (N_7568,N_7472,N_7437);
and U7569 (N_7569,N_7404,N_7445);
and U7570 (N_7570,N_7499,N_7410);
nor U7571 (N_7571,N_7386,N_7497);
or U7572 (N_7572,N_7382,N_7469);
nand U7573 (N_7573,N_7379,N_7499);
or U7574 (N_7574,N_7438,N_7422);
and U7575 (N_7575,N_7403,N_7402);
nor U7576 (N_7576,N_7463,N_7437);
or U7577 (N_7577,N_7390,N_7488);
xnor U7578 (N_7578,N_7378,N_7388);
and U7579 (N_7579,N_7460,N_7397);
and U7580 (N_7580,N_7439,N_7456);
xor U7581 (N_7581,N_7383,N_7425);
or U7582 (N_7582,N_7446,N_7426);
nand U7583 (N_7583,N_7403,N_7378);
xnor U7584 (N_7584,N_7467,N_7418);
or U7585 (N_7585,N_7430,N_7471);
or U7586 (N_7586,N_7422,N_7489);
or U7587 (N_7587,N_7453,N_7444);
xor U7588 (N_7588,N_7478,N_7387);
and U7589 (N_7589,N_7488,N_7375);
nor U7590 (N_7590,N_7457,N_7455);
xor U7591 (N_7591,N_7380,N_7494);
xor U7592 (N_7592,N_7432,N_7382);
xnor U7593 (N_7593,N_7474,N_7424);
nor U7594 (N_7594,N_7459,N_7471);
or U7595 (N_7595,N_7497,N_7489);
and U7596 (N_7596,N_7441,N_7448);
nor U7597 (N_7597,N_7461,N_7393);
nor U7598 (N_7598,N_7455,N_7414);
xor U7599 (N_7599,N_7441,N_7478);
or U7600 (N_7600,N_7495,N_7424);
and U7601 (N_7601,N_7427,N_7470);
nand U7602 (N_7602,N_7420,N_7408);
and U7603 (N_7603,N_7409,N_7470);
nor U7604 (N_7604,N_7398,N_7447);
xor U7605 (N_7605,N_7378,N_7461);
nand U7606 (N_7606,N_7416,N_7442);
and U7607 (N_7607,N_7402,N_7470);
and U7608 (N_7608,N_7429,N_7391);
xor U7609 (N_7609,N_7499,N_7387);
nand U7610 (N_7610,N_7473,N_7410);
nand U7611 (N_7611,N_7471,N_7446);
or U7612 (N_7612,N_7396,N_7463);
nor U7613 (N_7613,N_7418,N_7464);
xnor U7614 (N_7614,N_7451,N_7466);
and U7615 (N_7615,N_7478,N_7460);
xor U7616 (N_7616,N_7398,N_7405);
nor U7617 (N_7617,N_7412,N_7480);
xor U7618 (N_7618,N_7469,N_7390);
xnor U7619 (N_7619,N_7492,N_7436);
and U7620 (N_7620,N_7445,N_7478);
xnor U7621 (N_7621,N_7494,N_7472);
and U7622 (N_7622,N_7402,N_7421);
and U7623 (N_7623,N_7442,N_7450);
xor U7624 (N_7624,N_7376,N_7478);
and U7625 (N_7625,N_7522,N_7607);
nand U7626 (N_7626,N_7581,N_7507);
nor U7627 (N_7627,N_7527,N_7531);
and U7628 (N_7628,N_7547,N_7594);
nor U7629 (N_7629,N_7583,N_7603);
or U7630 (N_7630,N_7598,N_7509);
or U7631 (N_7631,N_7536,N_7579);
xor U7632 (N_7632,N_7503,N_7608);
or U7633 (N_7633,N_7596,N_7618);
nor U7634 (N_7634,N_7568,N_7512);
nand U7635 (N_7635,N_7595,N_7622);
nand U7636 (N_7636,N_7524,N_7575);
nor U7637 (N_7637,N_7535,N_7610);
xor U7638 (N_7638,N_7556,N_7580);
or U7639 (N_7639,N_7571,N_7553);
and U7640 (N_7640,N_7533,N_7506);
nor U7641 (N_7641,N_7572,N_7514);
nor U7642 (N_7642,N_7541,N_7578);
xnor U7643 (N_7643,N_7567,N_7609);
nand U7644 (N_7644,N_7582,N_7534);
and U7645 (N_7645,N_7601,N_7517);
and U7646 (N_7646,N_7584,N_7604);
nor U7647 (N_7647,N_7550,N_7552);
or U7648 (N_7648,N_7569,N_7516);
xor U7649 (N_7649,N_7544,N_7562);
nand U7650 (N_7650,N_7508,N_7558);
nor U7651 (N_7651,N_7505,N_7559);
xnor U7652 (N_7652,N_7530,N_7617);
nor U7653 (N_7653,N_7591,N_7525);
and U7654 (N_7654,N_7624,N_7611);
or U7655 (N_7655,N_7540,N_7551);
or U7656 (N_7656,N_7621,N_7585);
or U7657 (N_7657,N_7549,N_7519);
and U7658 (N_7658,N_7560,N_7502);
and U7659 (N_7659,N_7538,N_7542);
and U7660 (N_7660,N_7504,N_7532);
nand U7661 (N_7661,N_7526,N_7586);
and U7662 (N_7662,N_7501,N_7619);
and U7663 (N_7663,N_7613,N_7513);
and U7664 (N_7664,N_7587,N_7529);
and U7665 (N_7665,N_7557,N_7570);
or U7666 (N_7666,N_7592,N_7563);
or U7667 (N_7667,N_7593,N_7599);
nor U7668 (N_7668,N_7510,N_7623);
or U7669 (N_7669,N_7515,N_7588);
and U7670 (N_7670,N_7528,N_7555);
xnor U7671 (N_7671,N_7566,N_7564);
nor U7672 (N_7672,N_7602,N_7521);
and U7673 (N_7673,N_7577,N_7573);
nor U7674 (N_7674,N_7612,N_7589);
nor U7675 (N_7675,N_7554,N_7600);
xor U7676 (N_7676,N_7520,N_7616);
or U7677 (N_7677,N_7605,N_7574);
and U7678 (N_7678,N_7548,N_7614);
nor U7679 (N_7679,N_7537,N_7561);
xnor U7680 (N_7680,N_7597,N_7539);
nor U7681 (N_7681,N_7511,N_7590);
and U7682 (N_7682,N_7546,N_7576);
nor U7683 (N_7683,N_7620,N_7523);
and U7684 (N_7684,N_7606,N_7545);
xnor U7685 (N_7685,N_7543,N_7500);
or U7686 (N_7686,N_7615,N_7518);
nor U7687 (N_7687,N_7565,N_7582);
and U7688 (N_7688,N_7556,N_7605);
or U7689 (N_7689,N_7553,N_7558);
nand U7690 (N_7690,N_7563,N_7529);
and U7691 (N_7691,N_7501,N_7500);
or U7692 (N_7692,N_7550,N_7571);
nor U7693 (N_7693,N_7574,N_7526);
xor U7694 (N_7694,N_7509,N_7599);
and U7695 (N_7695,N_7550,N_7608);
nand U7696 (N_7696,N_7603,N_7607);
and U7697 (N_7697,N_7604,N_7531);
nand U7698 (N_7698,N_7571,N_7578);
or U7699 (N_7699,N_7587,N_7509);
and U7700 (N_7700,N_7595,N_7521);
and U7701 (N_7701,N_7577,N_7501);
or U7702 (N_7702,N_7532,N_7582);
and U7703 (N_7703,N_7513,N_7560);
or U7704 (N_7704,N_7514,N_7620);
nor U7705 (N_7705,N_7574,N_7510);
nand U7706 (N_7706,N_7610,N_7548);
nand U7707 (N_7707,N_7552,N_7502);
or U7708 (N_7708,N_7545,N_7603);
nor U7709 (N_7709,N_7581,N_7577);
or U7710 (N_7710,N_7568,N_7521);
nand U7711 (N_7711,N_7516,N_7611);
nor U7712 (N_7712,N_7514,N_7541);
xor U7713 (N_7713,N_7556,N_7529);
nand U7714 (N_7714,N_7571,N_7511);
nand U7715 (N_7715,N_7572,N_7555);
or U7716 (N_7716,N_7572,N_7578);
nand U7717 (N_7717,N_7593,N_7506);
xnor U7718 (N_7718,N_7586,N_7565);
nand U7719 (N_7719,N_7534,N_7539);
or U7720 (N_7720,N_7591,N_7541);
xor U7721 (N_7721,N_7602,N_7592);
nor U7722 (N_7722,N_7524,N_7588);
nor U7723 (N_7723,N_7593,N_7597);
nand U7724 (N_7724,N_7595,N_7564);
and U7725 (N_7725,N_7522,N_7576);
nand U7726 (N_7726,N_7504,N_7599);
xnor U7727 (N_7727,N_7592,N_7505);
xnor U7728 (N_7728,N_7546,N_7613);
and U7729 (N_7729,N_7597,N_7510);
and U7730 (N_7730,N_7531,N_7586);
nand U7731 (N_7731,N_7609,N_7501);
xor U7732 (N_7732,N_7584,N_7538);
xor U7733 (N_7733,N_7585,N_7549);
or U7734 (N_7734,N_7607,N_7567);
nor U7735 (N_7735,N_7521,N_7567);
xor U7736 (N_7736,N_7552,N_7574);
xor U7737 (N_7737,N_7517,N_7547);
xor U7738 (N_7738,N_7573,N_7579);
nand U7739 (N_7739,N_7602,N_7604);
nand U7740 (N_7740,N_7510,N_7584);
nor U7741 (N_7741,N_7557,N_7578);
xor U7742 (N_7742,N_7622,N_7590);
nand U7743 (N_7743,N_7542,N_7585);
and U7744 (N_7744,N_7618,N_7538);
xnor U7745 (N_7745,N_7575,N_7609);
nor U7746 (N_7746,N_7560,N_7589);
and U7747 (N_7747,N_7535,N_7520);
nor U7748 (N_7748,N_7577,N_7615);
or U7749 (N_7749,N_7503,N_7610);
xor U7750 (N_7750,N_7668,N_7722);
nand U7751 (N_7751,N_7742,N_7633);
or U7752 (N_7752,N_7697,N_7738);
xnor U7753 (N_7753,N_7708,N_7703);
nor U7754 (N_7754,N_7684,N_7639);
or U7755 (N_7755,N_7718,N_7655);
nand U7756 (N_7756,N_7665,N_7712);
and U7757 (N_7757,N_7680,N_7667);
nor U7758 (N_7758,N_7659,N_7692);
or U7759 (N_7759,N_7647,N_7646);
nor U7760 (N_7760,N_7634,N_7716);
and U7761 (N_7761,N_7746,N_7686);
or U7762 (N_7762,N_7625,N_7706);
and U7763 (N_7763,N_7663,N_7656);
or U7764 (N_7764,N_7630,N_7707);
and U7765 (N_7765,N_7711,N_7715);
nor U7766 (N_7766,N_7724,N_7710);
or U7767 (N_7767,N_7632,N_7700);
nand U7768 (N_7768,N_7652,N_7627);
xnor U7769 (N_7769,N_7705,N_7720);
nor U7770 (N_7770,N_7645,N_7679);
nand U7771 (N_7771,N_7674,N_7628);
or U7772 (N_7772,N_7733,N_7666);
xnor U7773 (N_7773,N_7719,N_7696);
or U7774 (N_7774,N_7734,N_7648);
or U7775 (N_7775,N_7640,N_7717);
or U7776 (N_7776,N_7727,N_7664);
and U7777 (N_7777,N_7730,N_7635);
or U7778 (N_7778,N_7739,N_7695);
and U7779 (N_7779,N_7747,N_7642);
xnor U7780 (N_7780,N_7660,N_7682);
or U7781 (N_7781,N_7694,N_7744);
xnor U7782 (N_7782,N_7657,N_7670);
or U7783 (N_7783,N_7702,N_7721);
and U7784 (N_7784,N_7681,N_7678);
xor U7785 (N_7785,N_7672,N_7709);
and U7786 (N_7786,N_7626,N_7661);
xor U7787 (N_7787,N_7745,N_7748);
xnor U7788 (N_7788,N_7690,N_7729);
and U7789 (N_7789,N_7735,N_7728);
nor U7790 (N_7790,N_7654,N_7637);
nand U7791 (N_7791,N_7731,N_7673);
nand U7792 (N_7792,N_7685,N_7701);
nor U7793 (N_7793,N_7693,N_7723);
and U7794 (N_7794,N_7740,N_7725);
and U7795 (N_7795,N_7698,N_7741);
xnor U7796 (N_7796,N_7638,N_7650);
nor U7797 (N_7797,N_7676,N_7649);
xor U7798 (N_7798,N_7704,N_7688);
and U7799 (N_7799,N_7658,N_7653);
xor U7800 (N_7800,N_7671,N_7687);
or U7801 (N_7801,N_7736,N_7726);
nor U7802 (N_7802,N_7749,N_7644);
and U7803 (N_7803,N_7629,N_7643);
xor U7804 (N_7804,N_7641,N_7713);
or U7805 (N_7805,N_7631,N_7732);
xnor U7806 (N_7806,N_7737,N_7651);
nor U7807 (N_7807,N_7714,N_7675);
and U7808 (N_7808,N_7691,N_7689);
or U7809 (N_7809,N_7699,N_7636);
nor U7810 (N_7810,N_7677,N_7662);
xnor U7811 (N_7811,N_7669,N_7743);
nand U7812 (N_7812,N_7683,N_7711);
nor U7813 (N_7813,N_7687,N_7652);
xnor U7814 (N_7814,N_7665,N_7735);
or U7815 (N_7815,N_7664,N_7741);
nor U7816 (N_7816,N_7719,N_7640);
or U7817 (N_7817,N_7739,N_7676);
and U7818 (N_7818,N_7718,N_7711);
nand U7819 (N_7819,N_7675,N_7718);
or U7820 (N_7820,N_7630,N_7629);
xnor U7821 (N_7821,N_7747,N_7660);
and U7822 (N_7822,N_7714,N_7718);
and U7823 (N_7823,N_7686,N_7736);
and U7824 (N_7824,N_7660,N_7673);
xnor U7825 (N_7825,N_7701,N_7639);
and U7826 (N_7826,N_7666,N_7700);
nand U7827 (N_7827,N_7636,N_7646);
and U7828 (N_7828,N_7746,N_7736);
xor U7829 (N_7829,N_7671,N_7741);
or U7830 (N_7830,N_7718,N_7650);
or U7831 (N_7831,N_7627,N_7746);
and U7832 (N_7832,N_7706,N_7682);
nand U7833 (N_7833,N_7711,N_7680);
nor U7834 (N_7834,N_7701,N_7636);
or U7835 (N_7835,N_7716,N_7678);
nand U7836 (N_7836,N_7739,N_7698);
xnor U7837 (N_7837,N_7671,N_7689);
or U7838 (N_7838,N_7728,N_7662);
or U7839 (N_7839,N_7668,N_7635);
and U7840 (N_7840,N_7675,N_7676);
nand U7841 (N_7841,N_7667,N_7673);
and U7842 (N_7842,N_7625,N_7724);
nor U7843 (N_7843,N_7675,N_7681);
or U7844 (N_7844,N_7642,N_7721);
nand U7845 (N_7845,N_7719,N_7635);
nand U7846 (N_7846,N_7655,N_7700);
and U7847 (N_7847,N_7703,N_7629);
nand U7848 (N_7848,N_7729,N_7635);
and U7849 (N_7849,N_7690,N_7648);
xor U7850 (N_7850,N_7649,N_7700);
xor U7851 (N_7851,N_7715,N_7666);
and U7852 (N_7852,N_7732,N_7701);
nor U7853 (N_7853,N_7748,N_7687);
and U7854 (N_7854,N_7643,N_7627);
xor U7855 (N_7855,N_7709,N_7708);
and U7856 (N_7856,N_7710,N_7687);
nor U7857 (N_7857,N_7689,N_7687);
and U7858 (N_7858,N_7721,N_7626);
or U7859 (N_7859,N_7647,N_7632);
xnor U7860 (N_7860,N_7666,N_7656);
and U7861 (N_7861,N_7673,N_7729);
xnor U7862 (N_7862,N_7677,N_7698);
and U7863 (N_7863,N_7641,N_7654);
and U7864 (N_7864,N_7727,N_7739);
or U7865 (N_7865,N_7661,N_7640);
nand U7866 (N_7866,N_7707,N_7736);
or U7867 (N_7867,N_7699,N_7685);
nand U7868 (N_7868,N_7697,N_7685);
nand U7869 (N_7869,N_7630,N_7674);
nand U7870 (N_7870,N_7652,N_7674);
or U7871 (N_7871,N_7733,N_7704);
and U7872 (N_7872,N_7642,N_7697);
xor U7873 (N_7873,N_7675,N_7644);
or U7874 (N_7874,N_7716,N_7736);
nand U7875 (N_7875,N_7842,N_7770);
xnor U7876 (N_7876,N_7817,N_7820);
nor U7877 (N_7877,N_7858,N_7867);
nor U7878 (N_7878,N_7807,N_7821);
nor U7879 (N_7879,N_7855,N_7778);
nand U7880 (N_7880,N_7774,N_7750);
nand U7881 (N_7881,N_7791,N_7805);
xor U7882 (N_7882,N_7872,N_7763);
and U7883 (N_7883,N_7822,N_7852);
nand U7884 (N_7884,N_7755,N_7794);
nor U7885 (N_7885,N_7874,N_7818);
xor U7886 (N_7886,N_7766,N_7839);
nor U7887 (N_7887,N_7809,N_7857);
and U7888 (N_7888,N_7767,N_7771);
nor U7889 (N_7889,N_7776,N_7832);
or U7890 (N_7890,N_7803,N_7854);
nand U7891 (N_7891,N_7873,N_7861);
nor U7892 (N_7892,N_7765,N_7793);
nand U7893 (N_7893,N_7851,N_7865);
or U7894 (N_7894,N_7823,N_7845);
nor U7895 (N_7895,N_7816,N_7824);
nand U7896 (N_7896,N_7813,N_7780);
and U7897 (N_7897,N_7826,N_7764);
and U7898 (N_7898,N_7801,N_7753);
nor U7899 (N_7899,N_7869,N_7843);
or U7900 (N_7900,N_7830,N_7758);
nor U7901 (N_7901,N_7859,N_7761);
xor U7902 (N_7902,N_7775,N_7837);
and U7903 (N_7903,N_7819,N_7762);
nor U7904 (N_7904,N_7777,N_7783);
and U7905 (N_7905,N_7847,N_7784);
nand U7906 (N_7906,N_7797,N_7863);
nand U7907 (N_7907,N_7785,N_7773);
xor U7908 (N_7908,N_7808,N_7871);
xnor U7909 (N_7909,N_7757,N_7759);
xor U7910 (N_7910,N_7835,N_7789);
xor U7911 (N_7911,N_7782,N_7825);
xor U7912 (N_7912,N_7868,N_7840);
nor U7913 (N_7913,N_7829,N_7870);
xor U7914 (N_7914,N_7834,N_7800);
xor U7915 (N_7915,N_7751,N_7804);
xnor U7916 (N_7916,N_7798,N_7853);
nand U7917 (N_7917,N_7752,N_7796);
xor U7918 (N_7918,N_7787,N_7848);
or U7919 (N_7919,N_7781,N_7844);
nor U7920 (N_7920,N_7792,N_7849);
and U7921 (N_7921,N_7772,N_7856);
nand U7922 (N_7922,N_7828,N_7769);
xor U7923 (N_7923,N_7866,N_7790);
nor U7924 (N_7924,N_7810,N_7846);
nor U7925 (N_7925,N_7799,N_7841);
or U7926 (N_7926,N_7812,N_7788);
nand U7927 (N_7927,N_7760,N_7779);
nand U7928 (N_7928,N_7838,N_7850);
or U7929 (N_7929,N_7831,N_7836);
nor U7930 (N_7930,N_7802,N_7754);
nor U7931 (N_7931,N_7795,N_7806);
or U7932 (N_7932,N_7814,N_7756);
and U7933 (N_7933,N_7811,N_7860);
or U7934 (N_7934,N_7815,N_7862);
and U7935 (N_7935,N_7864,N_7827);
or U7936 (N_7936,N_7786,N_7833);
or U7937 (N_7937,N_7768,N_7835);
xnor U7938 (N_7938,N_7807,N_7785);
and U7939 (N_7939,N_7852,N_7821);
or U7940 (N_7940,N_7761,N_7873);
or U7941 (N_7941,N_7858,N_7849);
nor U7942 (N_7942,N_7817,N_7765);
xnor U7943 (N_7943,N_7848,N_7754);
or U7944 (N_7944,N_7756,N_7757);
nand U7945 (N_7945,N_7862,N_7791);
and U7946 (N_7946,N_7805,N_7750);
or U7947 (N_7947,N_7800,N_7797);
nand U7948 (N_7948,N_7772,N_7859);
and U7949 (N_7949,N_7848,N_7814);
and U7950 (N_7950,N_7770,N_7848);
and U7951 (N_7951,N_7871,N_7864);
xnor U7952 (N_7952,N_7874,N_7777);
or U7953 (N_7953,N_7868,N_7870);
and U7954 (N_7954,N_7870,N_7776);
xor U7955 (N_7955,N_7787,N_7816);
nand U7956 (N_7956,N_7793,N_7815);
and U7957 (N_7957,N_7787,N_7827);
xnor U7958 (N_7958,N_7766,N_7770);
nand U7959 (N_7959,N_7820,N_7863);
nand U7960 (N_7960,N_7794,N_7837);
nand U7961 (N_7961,N_7874,N_7871);
xor U7962 (N_7962,N_7792,N_7779);
xor U7963 (N_7963,N_7833,N_7842);
or U7964 (N_7964,N_7772,N_7822);
xnor U7965 (N_7965,N_7771,N_7793);
and U7966 (N_7966,N_7843,N_7776);
and U7967 (N_7967,N_7771,N_7754);
nand U7968 (N_7968,N_7794,N_7831);
or U7969 (N_7969,N_7785,N_7839);
and U7970 (N_7970,N_7755,N_7799);
and U7971 (N_7971,N_7785,N_7750);
xnor U7972 (N_7972,N_7753,N_7758);
nor U7973 (N_7973,N_7750,N_7786);
nand U7974 (N_7974,N_7763,N_7757);
nand U7975 (N_7975,N_7804,N_7789);
or U7976 (N_7976,N_7863,N_7776);
and U7977 (N_7977,N_7859,N_7837);
or U7978 (N_7978,N_7770,N_7772);
xor U7979 (N_7979,N_7874,N_7793);
and U7980 (N_7980,N_7775,N_7776);
or U7981 (N_7981,N_7859,N_7846);
and U7982 (N_7982,N_7831,N_7759);
xnor U7983 (N_7983,N_7805,N_7795);
and U7984 (N_7984,N_7757,N_7795);
and U7985 (N_7985,N_7799,N_7855);
nor U7986 (N_7986,N_7813,N_7765);
or U7987 (N_7987,N_7814,N_7811);
nand U7988 (N_7988,N_7758,N_7782);
nand U7989 (N_7989,N_7815,N_7858);
nor U7990 (N_7990,N_7867,N_7837);
xnor U7991 (N_7991,N_7771,N_7821);
and U7992 (N_7992,N_7870,N_7867);
nor U7993 (N_7993,N_7830,N_7819);
xnor U7994 (N_7994,N_7772,N_7805);
and U7995 (N_7995,N_7836,N_7810);
xor U7996 (N_7996,N_7805,N_7810);
nand U7997 (N_7997,N_7776,N_7758);
or U7998 (N_7998,N_7774,N_7843);
or U7999 (N_7999,N_7792,N_7851);
nand U8000 (N_8000,N_7997,N_7887);
or U8001 (N_8001,N_7880,N_7953);
nor U8002 (N_8002,N_7954,N_7921);
xnor U8003 (N_8003,N_7964,N_7984);
and U8004 (N_8004,N_7989,N_7971);
nor U8005 (N_8005,N_7993,N_7894);
nor U8006 (N_8006,N_7878,N_7898);
nor U8007 (N_8007,N_7966,N_7947);
and U8008 (N_8008,N_7919,N_7977);
and U8009 (N_8009,N_7937,N_7890);
xnor U8010 (N_8010,N_7913,N_7920);
nand U8011 (N_8011,N_7892,N_7899);
or U8012 (N_8012,N_7960,N_7918);
xnor U8013 (N_8013,N_7967,N_7876);
or U8014 (N_8014,N_7986,N_7902);
and U8015 (N_8015,N_7914,N_7886);
or U8016 (N_8016,N_7957,N_7978);
nand U8017 (N_8017,N_7992,N_7934);
nor U8018 (N_8018,N_7924,N_7955);
and U8019 (N_8019,N_7976,N_7936);
xor U8020 (N_8020,N_7942,N_7969);
or U8021 (N_8021,N_7926,N_7963);
or U8022 (N_8022,N_7940,N_7904);
xnor U8023 (N_8023,N_7888,N_7943);
nor U8024 (N_8024,N_7990,N_7962);
nand U8025 (N_8025,N_7911,N_7879);
nand U8026 (N_8026,N_7952,N_7991);
nand U8027 (N_8027,N_7973,N_7999);
and U8028 (N_8028,N_7938,N_7896);
or U8029 (N_8029,N_7889,N_7956);
nand U8030 (N_8030,N_7891,N_7965);
and U8031 (N_8031,N_7959,N_7996);
nand U8032 (N_8032,N_7928,N_7895);
and U8033 (N_8033,N_7941,N_7910);
nand U8034 (N_8034,N_7980,N_7922);
nand U8035 (N_8035,N_7987,N_7968);
xnor U8036 (N_8036,N_7961,N_7877);
or U8037 (N_8037,N_7900,N_7906);
xor U8038 (N_8038,N_7939,N_7985);
nor U8039 (N_8039,N_7923,N_7884);
nand U8040 (N_8040,N_7945,N_7998);
nor U8041 (N_8041,N_7930,N_7903);
nor U8042 (N_8042,N_7883,N_7907);
and U8043 (N_8043,N_7982,N_7983);
nand U8044 (N_8044,N_7915,N_7901);
nor U8045 (N_8045,N_7909,N_7935);
nand U8046 (N_8046,N_7979,N_7975);
xor U8047 (N_8047,N_7927,N_7948);
nor U8048 (N_8048,N_7882,N_7974);
xnor U8049 (N_8049,N_7981,N_7925);
nor U8050 (N_8050,N_7995,N_7929);
xnor U8051 (N_8051,N_7885,N_7908);
xnor U8052 (N_8052,N_7972,N_7893);
and U8053 (N_8053,N_7912,N_7946);
and U8054 (N_8054,N_7917,N_7970);
nor U8055 (N_8055,N_7988,N_7944);
and U8056 (N_8056,N_7958,N_7881);
or U8057 (N_8057,N_7905,N_7875);
nand U8058 (N_8058,N_7951,N_7932);
or U8059 (N_8059,N_7931,N_7897);
and U8060 (N_8060,N_7994,N_7949);
xnor U8061 (N_8061,N_7933,N_7950);
xnor U8062 (N_8062,N_7916,N_7959);
nand U8063 (N_8063,N_7926,N_7974);
xnor U8064 (N_8064,N_7964,N_7931);
nand U8065 (N_8065,N_7959,N_7915);
or U8066 (N_8066,N_7915,N_7981);
or U8067 (N_8067,N_7992,N_7981);
nand U8068 (N_8068,N_7884,N_7922);
or U8069 (N_8069,N_7943,N_7920);
and U8070 (N_8070,N_7890,N_7932);
xor U8071 (N_8071,N_7877,N_7925);
nor U8072 (N_8072,N_7985,N_7888);
nand U8073 (N_8073,N_7914,N_7905);
xnor U8074 (N_8074,N_7977,N_7964);
xor U8075 (N_8075,N_7953,N_7904);
or U8076 (N_8076,N_7881,N_7891);
xnor U8077 (N_8077,N_7875,N_7903);
nand U8078 (N_8078,N_7968,N_7969);
xor U8079 (N_8079,N_7878,N_7917);
nand U8080 (N_8080,N_7914,N_7987);
nor U8081 (N_8081,N_7894,N_7954);
xnor U8082 (N_8082,N_7999,N_7941);
or U8083 (N_8083,N_7996,N_7921);
nand U8084 (N_8084,N_7901,N_7973);
or U8085 (N_8085,N_7933,N_7962);
xnor U8086 (N_8086,N_7876,N_7907);
xor U8087 (N_8087,N_7887,N_7937);
nand U8088 (N_8088,N_7971,N_7993);
and U8089 (N_8089,N_7996,N_7999);
nor U8090 (N_8090,N_7979,N_7973);
xnor U8091 (N_8091,N_7902,N_7957);
xor U8092 (N_8092,N_7914,N_7994);
nand U8093 (N_8093,N_7978,N_7992);
nand U8094 (N_8094,N_7890,N_7944);
nor U8095 (N_8095,N_7952,N_7921);
nand U8096 (N_8096,N_7942,N_7914);
nand U8097 (N_8097,N_7960,N_7888);
nand U8098 (N_8098,N_7980,N_7900);
nor U8099 (N_8099,N_7971,N_7910);
nor U8100 (N_8100,N_7948,N_7998);
nor U8101 (N_8101,N_7941,N_7956);
or U8102 (N_8102,N_7912,N_7879);
nand U8103 (N_8103,N_7954,N_7990);
or U8104 (N_8104,N_7898,N_7915);
xnor U8105 (N_8105,N_7941,N_7933);
nand U8106 (N_8106,N_7986,N_7983);
or U8107 (N_8107,N_7967,N_7997);
nand U8108 (N_8108,N_7924,N_7957);
nor U8109 (N_8109,N_7917,N_7909);
xnor U8110 (N_8110,N_7902,N_7900);
and U8111 (N_8111,N_7902,N_7956);
nand U8112 (N_8112,N_7891,N_7875);
xnor U8113 (N_8113,N_7921,N_7956);
or U8114 (N_8114,N_7910,N_7899);
xnor U8115 (N_8115,N_7895,N_7956);
xor U8116 (N_8116,N_7965,N_7897);
nand U8117 (N_8117,N_7985,N_7923);
nor U8118 (N_8118,N_7974,N_7976);
nor U8119 (N_8119,N_7979,N_7936);
or U8120 (N_8120,N_7963,N_7996);
nor U8121 (N_8121,N_7955,N_7949);
nor U8122 (N_8122,N_7953,N_7999);
nor U8123 (N_8123,N_7978,N_7949);
nor U8124 (N_8124,N_7886,N_7878);
or U8125 (N_8125,N_8004,N_8069);
nand U8126 (N_8126,N_8087,N_8106);
xnor U8127 (N_8127,N_8060,N_8113);
or U8128 (N_8128,N_8033,N_8108);
nor U8129 (N_8129,N_8048,N_8056);
nor U8130 (N_8130,N_8027,N_8121);
xor U8131 (N_8131,N_8035,N_8052);
or U8132 (N_8132,N_8111,N_8079);
nand U8133 (N_8133,N_8014,N_8039);
nand U8134 (N_8134,N_8116,N_8074);
and U8135 (N_8135,N_8012,N_8112);
and U8136 (N_8136,N_8088,N_8100);
nand U8137 (N_8137,N_8076,N_8024);
and U8138 (N_8138,N_8009,N_8018);
xor U8139 (N_8139,N_8065,N_8097);
and U8140 (N_8140,N_8021,N_8075);
or U8141 (N_8141,N_8054,N_8062);
nand U8142 (N_8142,N_8019,N_8059);
nor U8143 (N_8143,N_8083,N_8026);
or U8144 (N_8144,N_8045,N_8109);
nor U8145 (N_8145,N_8023,N_8030);
nor U8146 (N_8146,N_8119,N_8118);
and U8147 (N_8147,N_8006,N_8049);
or U8148 (N_8148,N_8029,N_8115);
nand U8149 (N_8149,N_8080,N_8025);
xor U8150 (N_8150,N_8068,N_8007);
nand U8151 (N_8151,N_8082,N_8042);
and U8152 (N_8152,N_8064,N_8067);
xnor U8153 (N_8153,N_8038,N_8050);
and U8154 (N_8154,N_8124,N_8031);
or U8155 (N_8155,N_8095,N_8053);
nand U8156 (N_8156,N_8013,N_8010);
xnor U8157 (N_8157,N_8047,N_8017);
or U8158 (N_8158,N_8005,N_8036);
and U8159 (N_8159,N_8022,N_8084);
and U8160 (N_8160,N_8044,N_8107);
and U8161 (N_8161,N_8070,N_8020);
and U8162 (N_8162,N_8094,N_8120);
nand U8163 (N_8163,N_8090,N_8066);
xor U8164 (N_8164,N_8046,N_8071);
nand U8165 (N_8165,N_8101,N_8081);
or U8166 (N_8166,N_8098,N_8077);
xnor U8167 (N_8167,N_8015,N_8117);
nand U8168 (N_8168,N_8089,N_8099);
nor U8169 (N_8169,N_8057,N_8016);
xnor U8170 (N_8170,N_8061,N_8086);
and U8171 (N_8171,N_8093,N_8008);
or U8172 (N_8172,N_8073,N_8028);
and U8173 (N_8173,N_8102,N_8096);
and U8174 (N_8174,N_8037,N_8040);
xnor U8175 (N_8175,N_8041,N_8055);
xor U8176 (N_8176,N_8032,N_8003);
nand U8177 (N_8177,N_8104,N_8103);
xnor U8178 (N_8178,N_8091,N_8051);
nand U8179 (N_8179,N_8110,N_8085);
and U8180 (N_8180,N_8011,N_8063);
xor U8181 (N_8181,N_8123,N_8034);
and U8182 (N_8182,N_8043,N_8000);
and U8183 (N_8183,N_8105,N_8001);
xor U8184 (N_8184,N_8078,N_8058);
or U8185 (N_8185,N_8114,N_8002);
and U8186 (N_8186,N_8122,N_8092);
nor U8187 (N_8187,N_8072,N_8031);
or U8188 (N_8188,N_8013,N_8114);
nand U8189 (N_8189,N_8050,N_8000);
nand U8190 (N_8190,N_8101,N_8084);
or U8191 (N_8191,N_8109,N_8074);
nor U8192 (N_8192,N_8083,N_8005);
nor U8193 (N_8193,N_8030,N_8066);
xnor U8194 (N_8194,N_8029,N_8042);
nor U8195 (N_8195,N_8039,N_8012);
and U8196 (N_8196,N_8019,N_8124);
xnor U8197 (N_8197,N_8039,N_8113);
and U8198 (N_8198,N_8121,N_8075);
nand U8199 (N_8199,N_8085,N_8002);
and U8200 (N_8200,N_8094,N_8118);
nand U8201 (N_8201,N_8032,N_8092);
nor U8202 (N_8202,N_8003,N_8079);
and U8203 (N_8203,N_8095,N_8025);
and U8204 (N_8204,N_8085,N_8051);
nand U8205 (N_8205,N_8056,N_8036);
xnor U8206 (N_8206,N_8072,N_8017);
nand U8207 (N_8207,N_8093,N_8106);
nand U8208 (N_8208,N_8015,N_8080);
nand U8209 (N_8209,N_8017,N_8102);
xor U8210 (N_8210,N_8026,N_8106);
and U8211 (N_8211,N_8081,N_8003);
and U8212 (N_8212,N_8123,N_8066);
nand U8213 (N_8213,N_8064,N_8050);
or U8214 (N_8214,N_8108,N_8010);
and U8215 (N_8215,N_8078,N_8085);
nor U8216 (N_8216,N_8026,N_8076);
and U8217 (N_8217,N_8088,N_8118);
and U8218 (N_8218,N_8032,N_8101);
or U8219 (N_8219,N_8012,N_8106);
or U8220 (N_8220,N_8104,N_8096);
or U8221 (N_8221,N_8072,N_8111);
nand U8222 (N_8222,N_8003,N_8056);
nand U8223 (N_8223,N_8091,N_8105);
and U8224 (N_8224,N_8110,N_8074);
nor U8225 (N_8225,N_8067,N_8001);
and U8226 (N_8226,N_8115,N_8088);
nand U8227 (N_8227,N_8037,N_8003);
nand U8228 (N_8228,N_8106,N_8098);
xnor U8229 (N_8229,N_8067,N_8120);
nor U8230 (N_8230,N_8058,N_8015);
xor U8231 (N_8231,N_8111,N_8061);
nand U8232 (N_8232,N_8104,N_8098);
xor U8233 (N_8233,N_8049,N_8099);
or U8234 (N_8234,N_8068,N_8003);
nand U8235 (N_8235,N_8009,N_8011);
and U8236 (N_8236,N_8102,N_8118);
and U8237 (N_8237,N_8008,N_8064);
or U8238 (N_8238,N_8040,N_8075);
nand U8239 (N_8239,N_8107,N_8051);
nand U8240 (N_8240,N_8094,N_8100);
xnor U8241 (N_8241,N_8052,N_8050);
xor U8242 (N_8242,N_8029,N_8074);
xnor U8243 (N_8243,N_8082,N_8116);
or U8244 (N_8244,N_8062,N_8036);
nor U8245 (N_8245,N_8053,N_8055);
nor U8246 (N_8246,N_8066,N_8082);
or U8247 (N_8247,N_8069,N_8076);
or U8248 (N_8248,N_8124,N_8095);
nor U8249 (N_8249,N_8050,N_8069);
nand U8250 (N_8250,N_8135,N_8229);
xor U8251 (N_8251,N_8149,N_8155);
nor U8252 (N_8252,N_8125,N_8202);
nand U8253 (N_8253,N_8129,N_8194);
or U8254 (N_8254,N_8249,N_8225);
and U8255 (N_8255,N_8219,N_8172);
nor U8256 (N_8256,N_8232,N_8164);
and U8257 (N_8257,N_8142,N_8151);
and U8258 (N_8258,N_8235,N_8183);
or U8259 (N_8259,N_8127,N_8133);
or U8260 (N_8260,N_8178,N_8213);
xnor U8261 (N_8261,N_8247,N_8246);
or U8262 (N_8262,N_8205,N_8243);
nor U8263 (N_8263,N_8131,N_8198);
or U8264 (N_8264,N_8216,N_8166);
nand U8265 (N_8265,N_8210,N_8214);
nand U8266 (N_8266,N_8208,N_8146);
nand U8267 (N_8267,N_8211,N_8148);
or U8268 (N_8268,N_8222,N_8185);
xor U8269 (N_8269,N_8157,N_8224);
nor U8270 (N_8270,N_8245,N_8215);
nor U8271 (N_8271,N_8203,N_8218);
nand U8272 (N_8272,N_8207,N_8152);
nand U8273 (N_8273,N_8163,N_8159);
nand U8274 (N_8274,N_8136,N_8165);
nand U8275 (N_8275,N_8236,N_8223);
and U8276 (N_8276,N_8195,N_8189);
xnor U8277 (N_8277,N_8170,N_8181);
nand U8278 (N_8278,N_8242,N_8184);
or U8279 (N_8279,N_8179,N_8197);
nand U8280 (N_8280,N_8143,N_8226);
nor U8281 (N_8281,N_8201,N_8233);
nor U8282 (N_8282,N_8134,N_8173);
nor U8283 (N_8283,N_8180,N_8227);
nand U8284 (N_8284,N_8239,N_8231);
or U8285 (N_8285,N_8191,N_8153);
xor U8286 (N_8286,N_8209,N_8190);
xor U8287 (N_8287,N_8187,N_8182);
xor U8288 (N_8288,N_8169,N_8137);
and U8289 (N_8289,N_8175,N_8196);
and U8290 (N_8290,N_8150,N_8217);
nand U8291 (N_8291,N_8171,N_8186);
and U8292 (N_8292,N_8220,N_8139);
xor U8293 (N_8293,N_8193,N_8176);
xnor U8294 (N_8294,N_8132,N_8240);
nand U8295 (N_8295,N_8162,N_8168);
nor U8296 (N_8296,N_8230,N_8130);
and U8297 (N_8297,N_8212,N_8237);
nand U8298 (N_8298,N_8177,N_8126);
and U8299 (N_8299,N_8141,N_8167);
and U8300 (N_8300,N_8174,N_8248);
xnor U8301 (N_8301,N_8128,N_8147);
nor U8302 (N_8302,N_8144,N_8206);
nand U8303 (N_8303,N_8138,N_8140);
and U8304 (N_8304,N_8158,N_8160);
and U8305 (N_8305,N_8234,N_8238);
nand U8306 (N_8306,N_8244,N_8204);
and U8307 (N_8307,N_8200,N_8199);
or U8308 (N_8308,N_8154,N_8228);
xnor U8309 (N_8309,N_8241,N_8156);
nand U8310 (N_8310,N_8145,N_8188);
xor U8311 (N_8311,N_8221,N_8161);
nor U8312 (N_8312,N_8192,N_8168);
xor U8313 (N_8313,N_8129,N_8184);
nor U8314 (N_8314,N_8204,N_8145);
nand U8315 (N_8315,N_8155,N_8200);
xor U8316 (N_8316,N_8221,N_8194);
and U8317 (N_8317,N_8148,N_8192);
and U8318 (N_8318,N_8213,N_8185);
or U8319 (N_8319,N_8129,N_8193);
nor U8320 (N_8320,N_8223,N_8197);
or U8321 (N_8321,N_8174,N_8175);
xor U8322 (N_8322,N_8182,N_8228);
xnor U8323 (N_8323,N_8168,N_8157);
nand U8324 (N_8324,N_8205,N_8247);
nand U8325 (N_8325,N_8179,N_8128);
and U8326 (N_8326,N_8159,N_8204);
nand U8327 (N_8327,N_8135,N_8181);
and U8328 (N_8328,N_8189,N_8204);
nor U8329 (N_8329,N_8173,N_8167);
xnor U8330 (N_8330,N_8159,N_8245);
nor U8331 (N_8331,N_8203,N_8229);
xnor U8332 (N_8332,N_8154,N_8214);
or U8333 (N_8333,N_8192,N_8208);
nor U8334 (N_8334,N_8208,N_8230);
or U8335 (N_8335,N_8160,N_8240);
nand U8336 (N_8336,N_8197,N_8137);
or U8337 (N_8337,N_8208,N_8242);
nand U8338 (N_8338,N_8171,N_8204);
nand U8339 (N_8339,N_8190,N_8235);
or U8340 (N_8340,N_8188,N_8129);
nor U8341 (N_8341,N_8239,N_8216);
xor U8342 (N_8342,N_8144,N_8189);
or U8343 (N_8343,N_8141,N_8234);
nor U8344 (N_8344,N_8210,N_8219);
nand U8345 (N_8345,N_8166,N_8134);
nand U8346 (N_8346,N_8249,N_8142);
nand U8347 (N_8347,N_8235,N_8138);
xnor U8348 (N_8348,N_8183,N_8169);
nor U8349 (N_8349,N_8175,N_8245);
nand U8350 (N_8350,N_8179,N_8181);
or U8351 (N_8351,N_8180,N_8215);
xor U8352 (N_8352,N_8222,N_8241);
xor U8353 (N_8353,N_8164,N_8231);
or U8354 (N_8354,N_8241,N_8159);
nand U8355 (N_8355,N_8181,N_8203);
nand U8356 (N_8356,N_8224,N_8136);
xor U8357 (N_8357,N_8142,N_8159);
nor U8358 (N_8358,N_8231,N_8210);
or U8359 (N_8359,N_8189,N_8133);
nand U8360 (N_8360,N_8223,N_8193);
or U8361 (N_8361,N_8164,N_8241);
and U8362 (N_8362,N_8198,N_8221);
and U8363 (N_8363,N_8180,N_8245);
and U8364 (N_8364,N_8147,N_8140);
or U8365 (N_8365,N_8185,N_8178);
and U8366 (N_8366,N_8164,N_8221);
and U8367 (N_8367,N_8205,N_8200);
nand U8368 (N_8368,N_8146,N_8199);
nand U8369 (N_8369,N_8147,N_8174);
or U8370 (N_8370,N_8144,N_8177);
or U8371 (N_8371,N_8170,N_8153);
nor U8372 (N_8372,N_8200,N_8159);
nor U8373 (N_8373,N_8131,N_8168);
and U8374 (N_8374,N_8227,N_8159);
nor U8375 (N_8375,N_8368,N_8260);
nor U8376 (N_8376,N_8363,N_8259);
or U8377 (N_8377,N_8352,N_8314);
xor U8378 (N_8378,N_8350,N_8264);
and U8379 (N_8379,N_8373,N_8346);
xor U8380 (N_8380,N_8374,N_8337);
and U8381 (N_8381,N_8256,N_8334);
nor U8382 (N_8382,N_8299,N_8253);
and U8383 (N_8383,N_8269,N_8330);
nand U8384 (N_8384,N_8336,N_8284);
and U8385 (N_8385,N_8370,N_8295);
nor U8386 (N_8386,N_8328,N_8265);
or U8387 (N_8387,N_8323,N_8358);
and U8388 (N_8388,N_8304,N_8278);
xor U8389 (N_8389,N_8303,N_8339);
or U8390 (N_8390,N_8254,N_8322);
xor U8391 (N_8391,N_8309,N_8296);
and U8392 (N_8392,N_8372,N_8273);
or U8393 (N_8393,N_8355,N_8349);
xnor U8394 (N_8394,N_8366,N_8294);
nor U8395 (N_8395,N_8266,N_8283);
and U8396 (N_8396,N_8255,N_8258);
nor U8397 (N_8397,N_8300,N_8301);
xor U8398 (N_8398,N_8289,N_8308);
and U8399 (N_8399,N_8292,N_8325);
or U8400 (N_8400,N_8343,N_8362);
or U8401 (N_8401,N_8310,N_8293);
nand U8402 (N_8402,N_8371,N_8275);
or U8403 (N_8403,N_8298,N_8319);
nor U8404 (N_8404,N_8267,N_8340);
nor U8405 (N_8405,N_8307,N_8338);
nor U8406 (N_8406,N_8287,N_8361);
or U8407 (N_8407,N_8280,N_8274);
or U8408 (N_8408,N_8270,N_8252);
xor U8409 (N_8409,N_8364,N_8351);
and U8410 (N_8410,N_8291,N_8342);
or U8411 (N_8411,N_8261,N_8297);
nand U8412 (N_8412,N_8354,N_8302);
nor U8413 (N_8413,N_8332,N_8320);
xnor U8414 (N_8414,N_8272,N_8359);
or U8415 (N_8415,N_8286,N_8324);
or U8416 (N_8416,N_8277,N_8285);
and U8417 (N_8417,N_8347,N_8251);
nor U8418 (N_8418,N_8268,N_8276);
nand U8419 (N_8419,N_8345,N_8353);
and U8420 (N_8420,N_8341,N_8279);
or U8421 (N_8421,N_8311,N_8288);
nor U8422 (N_8422,N_8306,N_8263);
nor U8423 (N_8423,N_8331,N_8257);
or U8424 (N_8424,N_8318,N_8369);
and U8425 (N_8425,N_8282,N_8326);
and U8426 (N_8426,N_8365,N_8271);
nor U8427 (N_8427,N_8348,N_8344);
nor U8428 (N_8428,N_8262,N_8335);
or U8429 (N_8429,N_8333,N_8316);
xnor U8430 (N_8430,N_8312,N_8357);
nand U8431 (N_8431,N_8305,N_8327);
nor U8432 (N_8432,N_8315,N_8290);
nand U8433 (N_8433,N_8367,N_8250);
nor U8434 (N_8434,N_8313,N_8317);
or U8435 (N_8435,N_8360,N_8281);
nand U8436 (N_8436,N_8329,N_8356);
nand U8437 (N_8437,N_8321,N_8333);
xor U8438 (N_8438,N_8315,N_8373);
and U8439 (N_8439,N_8278,N_8296);
and U8440 (N_8440,N_8333,N_8372);
or U8441 (N_8441,N_8270,N_8295);
nand U8442 (N_8442,N_8305,N_8274);
xor U8443 (N_8443,N_8254,N_8306);
nor U8444 (N_8444,N_8258,N_8365);
xor U8445 (N_8445,N_8356,N_8359);
and U8446 (N_8446,N_8336,N_8250);
or U8447 (N_8447,N_8266,N_8280);
nor U8448 (N_8448,N_8342,N_8298);
nor U8449 (N_8449,N_8301,N_8308);
nand U8450 (N_8450,N_8285,N_8325);
nand U8451 (N_8451,N_8289,N_8362);
nor U8452 (N_8452,N_8302,N_8310);
xnor U8453 (N_8453,N_8334,N_8327);
nor U8454 (N_8454,N_8351,N_8349);
or U8455 (N_8455,N_8271,N_8285);
or U8456 (N_8456,N_8364,N_8255);
or U8457 (N_8457,N_8261,N_8324);
nor U8458 (N_8458,N_8273,N_8340);
or U8459 (N_8459,N_8256,N_8265);
xor U8460 (N_8460,N_8352,N_8325);
and U8461 (N_8461,N_8362,N_8286);
and U8462 (N_8462,N_8302,N_8371);
and U8463 (N_8463,N_8291,N_8338);
or U8464 (N_8464,N_8360,N_8276);
xnor U8465 (N_8465,N_8267,N_8348);
nand U8466 (N_8466,N_8295,N_8327);
nor U8467 (N_8467,N_8313,N_8285);
and U8468 (N_8468,N_8348,N_8264);
xor U8469 (N_8469,N_8358,N_8308);
or U8470 (N_8470,N_8318,N_8336);
or U8471 (N_8471,N_8373,N_8339);
and U8472 (N_8472,N_8347,N_8331);
nor U8473 (N_8473,N_8338,N_8288);
or U8474 (N_8474,N_8285,N_8318);
xnor U8475 (N_8475,N_8250,N_8261);
or U8476 (N_8476,N_8305,N_8270);
xor U8477 (N_8477,N_8276,N_8374);
or U8478 (N_8478,N_8260,N_8367);
nor U8479 (N_8479,N_8337,N_8367);
or U8480 (N_8480,N_8343,N_8292);
or U8481 (N_8481,N_8251,N_8349);
or U8482 (N_8482,N_8311,N_8330);
and U8483 (N_8483,N_8267,N_8329);
nor U8484 (N_8484,N_8373,N_8280);
or U8485 (N_8485,N_8353,N_8374);
nand U8486 (N_8486,N_8262,N_8259);
and U8487 (N_8487,N_8352,N_8272);
nor U8488 (N_8488,N_8260,N_8302);
or U8489 (N_8489,N_8255,N_8295);
xor U8490 (N_8490,N_8326,N_8337);
nand U8491 (N_8491,N_8350,N_8316);
xnor U8492 (N_8492,N_8297,N_8363);
or U8493 (N_8493,N_8309,N_8262);
nand U8494 (N_8494,N_8267,N_8332);
and U8495 (N_8495,N_8256,N_8255);
nor U8496 (N_8496,N_8354,N_8363);
xor U8497 (N_8497,N_8362,N_8294);
or U8498 (N_8498,N_8309,N_8306);
and U8499 (N_8499,N_8266,N_8259);
nor U8500 (N_8500,N_8388,N_8490);
and U8501 (N_8501,N_8412,N_8403);
and U8502 (N_8502,N_8437,N_8424);
xor U8503 (N_8503,N_8466,N_8494);
and U8504 (N_8504,N_8486,N_8391);
xnor U8505 (N_8505,N_8382,N_8418);
or U8506 (N_8506,N_8489,N_8478);
and U8507 (N_8507,N_8465,N_8433);
xor U8508 (N_8508,N_8386,N_8428);
xor U8509 (N_8509,N_8458,N_8463);
or U8510 (N_8510,N_8392,N_8434);
and U8511 (N_8511,N_8449,N_8447);
xnor U8512 (N_8512,N_8396,N_8380);
and U8513 (N_8513,N_8499,N_8409);
xnor U8514 (N_8514,N_8444,N_8479);
xnor U8515 (N_8515,N_8404,N_8453);
xnor U8516 (N_8516,N_8473,N_8413);
nand U8517 (N_8517,N_8474,N_8410);
or U8518 (N_8518,N_8414,N_8416);
and U8519 (N_8519,N_8468,N_8495);
and U8520 (N_8520,N_8487,N_8464);
xnor U8521 (N_8521,N_8484,N_8422);
and U8522 (N_8522,N_8405,N_8398);
nor U8523 (N_8523,N_8470,N_8407);
or U8524 (N_8524,N_8402,N_8378);
nand U8525 (N_8525,N_8445,N_8452);
or U8526 (N_8526,N_8488,N_8485);
or U8527 (N_8527,N_8435,N_8469);
or U8528 (N_8528,N_8451,N_8411);
nand U8529 (N_8529,N_8441,N_8450);
or U8530 (N_8530,N_8429,N_8419);
and U8531 (N_8531,N_8446,N_8493);
and U8532 (N_8532,N_8483,N_8415);
nand U8533 (N_8533,N_8482,N_8421);
and U8534 (N_8534,N_8472,N_8467);
and U8535 (N_8535,N_8420,N_8389);
xor U8536 (N_8536,N_8423,N_8491);
nor U8537 (N_8537,N_8408,N_8436);
or U8538 (N_8538,N_8397,N_8461);
or U8539 (N_8539,N_8400,N_8431);
or U8540 (N_8540,N_8496,N_8454);
nor U8541 (N_8541,N_8492,N_8475);
or U8542 (N_8542,N_8377,N_8476);
nand U8543 (N_8543,N_8390,N_8383);
and U8544 (N_8544,N_8406,N_8471);
nand U8545 (N_8545,N_8498,N_8425);
nor U8546 (N_8546,N_8440,N_8426);
nor U8547 (N_8547,N_8394,N_8480);
or U8548 (N_8548,N_8399,N_8427);
xor U8549 (N_8549,N_8457,N_8442);
and U8550 (N_8550,N_8455,N_8439);
or U8551 (N_8551,N_8381,N_8448);
xnor U8552 (N_8552,N_8393,N_8430);
nor U8553 (N_8553,N_8376,N_8375);
nand U8554 (N_8554,N_8385,N_8438);
nand U8555 (N_8555,N_8460,N_8477);
xor U8556 (N_8556,N_8417,N_8432);
nor U8557 (N_8557,N_8456,N_8379);
nor U8558 (N_8558,N_8497,N_8462);
nand U8559 (N_8559,N_8443,N_8387);
nand U8560 (N_8560,N_8401,N_8459);
xor U8561 (N_8561,N_8481,N_8384);
or U8562 (N_8562,N_8395,N_8428);
or U8563 (N_8563,N_8429,N_8389);
or U8564 (N_8564,N_8420,N_8415);
and U8565 (N_8565,N_8387,N_8401);
or U8566 (N_8566,N_8466,N_8421);
nor U8567 (N_8567,N_8403,N_8391);
nand U8568 (N_8568,N_8443,N_8406);
nor U8569 (N_8569,N_8494,N_8388);
or U8570 (N_8570,N_8462,N_8378);
or U8571 (N_8571,N_8376,N_8493);
xor U8572 (N_8572,N_8477,N_8495);
nor U8573 (N_8573,N_8454,N_8413);
nor U8574 (N_8574,N_8457,N_8429);
and U8575 (N_8575,N_8476,N_8493);
nor U8576 (N_8576,N_8475,N_8403);
nor U8577 (N_8577,N_8399,N_8481);
nand U8578 (N_8578,N_8437,N_8400);
xnor U8579 (N_8579,N_8438,N_8470);
xnor U8580 (N_8580,N_8453,N_8393);
xnor U8581 (N_8581,N_8460,N_8388);
nand U8582 (N_8582,N_8478,N_8467);
and U8583 (N_8583,N_8456,N_8400);
and U8584 (N_8584,N_8418,N_8389);
or U8585 (N_8585,N_8484,N_8380);
nor U8586 (N_8586,N_8411,N_8473);
or U8587 (N_8587,N_8465,N_8489);
and U8588 (N_8588,N_8493,N_8494);
or U8589 (N_8589,N_8392,N_8413);
nor U8590 (N_8590,N_8417,N_8444);
nor U8591 (N_8591,N_8411,N_8488);
nor U8592 (N_8592,N_8442,N_8489);
nand U8593 (N_8593,N_8455,N_8413);
and U8594 (N_8594,N_8380,N_8415);
xor U8595 (N_8595,N_8476,N_8491);
xor U8596 (N_8596,N_8429,N_8439);
and U8597 (N_8597,N_8390,N_8391);
or U8598 (N_8598,N_8419,N_8465);
nand U8599 (N_8599,N_8478,N_8388);
xor U8600 (N_8600,N_8455,N_8419);
nand U8601 (N_8601,N_8471,N_8455);
nor U8602 (N_8602,N_8423,N_8428);
nor U8603 (N_8603,N_8447,N_8395);
nor U8604 (N_8604,N_8457,N_8384);
nor U8605 (N_8605,N_8417,N_8385);
and U8606 (N_8606,N_8390,N_8386);
or U8607 (N_8607,N_8452,N_8498);
and U8608 (N_8608,N_8419,N_8382);
xnor U8609 (N_8609,N_8482,N_8383);
nand U8610 (N_8610,N_8406,N_8395);
or U8611 (N_8611,N_8455,N_8479);
nand U8612 (N_8612,N_8382,N_8463);
or U8613 (N_8613,N_8478,N_8412);
and U8614 (N_8614,N_8389,N_8403);
nand U8615 (N_8615,N_8451,N_8436);
nor U8616 (N_8616,N_8498,N_8497);
nand U8617 (N_8617,N_8387,N_8464);
nand U8618 (N_8618,N_8382,N_8431);
nor U8619 (N_8619,N_8381,N_8391);
and U8620 (N_8620,N_8487,N_8400);
and U8621 (N_8621,N_8449,N_8481);
and U8622 (N_8622,N_8451,N_8475);
nor U8623 (N_8623,N_8492,N_8381);
and U8624 (N_8624,N_8393,N_8495);
xor U8625 (N_8625,N_8523,N_8512);
nand U8626 (N_8626,N_8582,N_8563);
xnor U8627 (N_8627,N_8560,N_8578);
xor U8628 (N_8628,N_8588,N_8538);
nand U8629 (N_8629,N_8610,N_8573);
nand U8630 (N_8630,N_8541,N_8525);
nor U8631 (N_8631,N_8594,N_8619);
or U8632 (N_8632,N_8535,N_8599);
or U8633 (N_8633,N_8587,N_8576);
nor U8634 (N_8634,N_8571,N_8540);
xor U8635 (N_8635,N_8604,N_8609);
nand U8636 (N_8636,N_8569,N_8621);
nor U8637 (N_8637,N_8583,N_8592);
and U8638 (N_8638,N_8553,N_8600);
xor U8639 (N_8639,N_8518,N_8590);
nand U8640 (N_8640,N_8534,N_8612);
xor U8641 (N_8641,N_8572,N_8566);
xnor U8642 (N_8642,N_8562,N_8550);
or U8643 (N_8643,N_8543,N_8602);
nor U8644 (N_8644,N_8589,N_8605);
nand U8645 (N_8645,N_8527,N_8515);
xor U8646 (N_8646,N_8558,N_8584);
or U8647 (N_8647,N_8507,N_8537);
xor U8648 (N_8648,N_8520,N_8547);
xor U8649 (N_8649,N_8519,N_8581);
xnor U8650 (N_8650,N_8500,N_8528);
xor U8651 (N_8651,N_8598,N_8579);
or U8652 (N_8652,N_8622,N_8516);
nor U8653 (N_8653,N_8561,N_8595);
xor U8654 (N_8654,N_8568,N_8586);
nor U8655 (N_8655,N_8601,N_8533);
nand U8656 (N_8656,N_8510,N_8508);
and U8657 (N_8657,N_8521,N_8616);
nand U8658 (N_8658,N_8552,N_8574);
and U8659 (N_8659,N_8608,N_8603);
xnor U8660 (N_8660,N_8539,N_8585);
or U8661 (N_8661,N_8506,N_8530);
nand U8662 (N_8662,N_8613,N_8524);
or U8663 (N_8663,N_8570,N_8511);
or U8664 (N_8664,N_8514,N_8551);
nand U8665 (N_8665,N_8591,N_8546);
xnor U8666 (N_8666,N_8624,N_8596);
nor U8667 (N_8667,N_8614,N_8556);
nor U8668 (N_8668,N_8501,N_8504);
nand U8669 (N_8669,N_8567,N_8536);
nor U8670 (N_8670,N_8620,N_8503);
or U8671 (N_8671,N_8580,N_8522);
nand U8672 (N_8672,N_8542,N_8526);
or U8673 (N_8673,N_8611,N_8513);
or U8674 (N_8674,N_8607,N_8517);
nand U8675 (N_8675,N_8615,N_8531);
or U8676 (N_8676,N_8593,N_8509);
or U8677 (N_8677,N_8565,N_8554);
and U8678 (N_8678,N_8505,N_8548);
nand U8679 (N_8679,N_8564,N_8557);
or U8680 (N_8680,N_8618,N_8559);
xnor U8681 (N_8681,N_8577,N_8606);
xor U8682 (N_8682,N_8617,N_8555);
xor U8683 (N_8683,N_8623,N_8597);
and U8684 (N_8684,N_8502,N_8545);
or U8685 (N_8685,N_8549,N_8575);
nor U8686 (N_8686,N_8544,N_8532);
nand U8687 (N_8687,N_8529,N_8571);
xnor U8688 (N_8688,N_8515,N_8556);
and U8689 (N_8689,N_8537,N_8536);
xnor U8690 (N_8690,N_8503,N_8532);
and U8691 (N_8691,N_8606,N_8551);
or U8692 (N_8692,N_8536,N_8606);
nand U8693 (N_8693,N_8610,N_8615);
and U8694 (N_8694,N_8513,N_8535);
nand U8695 (N_8695,N_8616,N_8580);
nand U8696 (N_8696,N_8589,N_8576);
nor U8697 (N_8697,N_8543,N_8606);
and U8698 (N_8698,N_8586,N_8529);
nand U8699 (N_8699,N_8523,N_8527);
and U8700 (N_8700,N_8522,N_8578);
or U8701 (N_8701,N_8546,N_8509);
and U8702 (N_8702,N_8529,N_8525);
nand U8703 (N_8703,N_8579,N_8548);
and U8704 (N_8704,N_8563,N_8550);
or U8705 (N_8705,N_8537,N_8510);
nand U8706 (N_8706,N_8588,N_8563);
xor U8707 (N_8707,N_8601,N_8554);
nor U8708 (N_8708,N_8591,N_8611);
and U8709 (N_8709,N_8539,N_8579);
or U8710 (N_8710,N_8609,N_8532);
or U8711 (N_8711,N_8613,N_8581);
xnor U8712 (N_8712,N_8619,N_8620);
nand U8713 (N_8713,N_8526,N_8534);
nor U8714 (N_8714,N_8524,N_8583);
nor U8715 (N_8715,N_8614,N_8568);
nor U8716 (N_8716,N_8603,N_8589);
nor U8717 (N_8717,N_8515,N_8618);
nand U8718 (N_8718,N_8574,N_8531);
xor U8719 (N_8719,N_8544,N_8565);
xnor U8720 (N_8720,N_8531,N_8510);
nor U8721 (N_8721,N_8597,N_8540);
nor U8722 (N_8722,N_8569,N_8623);
and U8723 (N_8723,N_8522,N_8593);
or U8724 (N_8724,N_8591,N_8619);
nor U8725 (N_8725,N_8542,N_8581);
nor U8726 (N_8726,N_8581,N_8553);
xor U8727 (N_8727,N_8525,N_8549);
or U8728 (N_8728,N_8600,N_8587);
xor U8729 (N_8729,N_8617,N_8557);
nand U8730 (N_8730,N_8530,N_8615);
nor U8731 (N_8731,N_8609,N_8614);
nor U8732 (N_8732,N_8521,N_8531);
and U8733 (N_8733,N_8564,N_8521);
xnor U8734 (N_8734,N_8580,N_8575);
nor U8735 (N_8735,N_8594,N_8592);
nand U8736 (N_8736,N_8504,N_8580);
nand U8737 (N_8737,N_8604,N_8501);
nand U8738 (N_8738,N_8556,N_8542);
and U8739 (N_8739,N_8539,N_8517);
or U8740 (N_8740,N_8621,N_8520);
nand U8741 (N_8741,N_8550,N_8614);
nor U8742 (N_8742,N_8594,N_8529);
nand U8743 (N_8743,N_8512,N_8508);
and U8744 (N_8744,N_8578,N_8623);
and U8745 (N_8745,N_8533,N_8545);
and U8746 (N_8746,N_8618,N_8533);
and U8747 (N_8747,N_8557,N_8587);
nand U8748 (N_8748,N_8535,N_8515);
xor U8749 (N_8749,N_8582,N_8544);
nor U8750 (N_8750,N_8676,N_8677);
or U8751 (N_8751,N_8700,N_8675);
nor U8752 (N_8752,N_8661,N_8667);
nand U8753 (N_8753,N_8704,N_8663);
and U8754 (N_8754,N_8708,N_8695);
nand U8755 (N_8755,N_8674,N_8659);
and U8756 (N_8756,N_8688,N_8653);
and U8757 (N_8757,N_8724,N_8636);
or U8758 (N_8758,N_8687,N_8734);
xor U8759 (N_8759,N_8739,N_8694);
nor U8760 (N_8760,N_8629,N_8671);
xnor U8761 (N_8761,N_8628,N_8635);
or U8762 (N_8762,N_8703,N_8637);
and U8763 (N_8763,N_8710,N_8746);
and U8764 (N_8764,N_8642,N_8714);
or U8765 (N_8765,N_8657,N_8699);
or U8766 (N_8766,N_8728,N_8691);
nand U8767 (N_8767,N_8723,N_8626);
xor U8768 (N_8768,N_8705,N_8670);
or U8769 (N_8769,N_8721,N_8655);
and U8770 (N_8770,N_8693,N_8646);
or U8771 (N_8771,N_8662,N_8685);
nor U8772 (N_8772,N_8702,N_8740);
and U8773 (N_8773,N_8648,N_8698);
xnor U8774 (N_8774,N_8684,N_8744);
or U8775 (N_8775,N_8664,N_8747);
nor U8776 (N_8776,N_8741,N_8689);
or U8777 (N_8777,N_8641,N_8697);
or U8778 (N_8778,N_8665,N_8715);
xnor U8779 (N_8779,N_8720,N_8745);
or U8780 (N_8780,N_8660,N_8634);
and U8781 (N_8781,N_8706,N_8749);
or U8782 (N_8782,N_8748,N_8658);
and U8783 (N_8783,N_8649,N_8709);
xnor U8784 (N_8784,N_8718,N_8743);
or U8785 (N_8785,N_8729,N_8656);
nand U8786 (N_8786,N_8669,N_8683);
xor U8787 (N_8787,N_8726,N_8736);
and U8788 (N_8788,N_8645,N_8668);
xnor U8789 (N_8789,N_8742,N_8666);
xor U8790 (N_8790,N_8650,N_8672);
xor U8791 (N_8791,N_8643,N_8630);
or U8792 (N_8792,N_8678,N_8632);
or U8793 (N_8793,N_8696,N_8713);
and U8794 (N_8794,N_8639,N_8631);
and U8795 (N_8795,N_8652,N_8707);
xor U8796 (N_8796,N_8673,N_8682);
nand U8797 (N_8797,N_8686,N_8681);
nand U8798 (N_8798,N_8633,N_8732);
nand U8799 (N_8799,N_8680,N_8719);
nand U8800 (N_8800,N_8711,N_8651);
or U8801 (N_8801,N_8737,N_8647);
nor U8802 (N_8802,N_8712,N_8644);
and U8803 (N_8803,N_8716,N_8679);
and U8804 (N_8804,N_8731,N_8640);
xnor U8805 (N_8805,N_8654,N_8625);
nand U8806 (N_8806,N_8627,N_8638);
and U8807 (N_8807,N_8725,N_8738);
nor U8808 (N_8808,N_8692,N_8701);
nor U8809 (N_8809,N_8733,N_8717);
and U8810 (N_8810,N_8722,N_8735);
xnor U8811 (N_8811,N_8730,N_8690);
or U8812 (N_8812,N_8727,N_8632);
nor U8813 (N_8813,N_8721,N_8695);
or U8814 (N_8814,N_8679,N_8725);
xor U8815 (N_8815,N_8711,N_8663);
or U8816 (N_8816,N_8654,N_8745);
nand U8817 (N_8817,N_8707,N_8635);
or U8818 (N_8818,N_8691,N_8635);
xnor U8819 (N_8819,N_8700,N_8679);
xnor U8820 (N_8820,N_8708,N_8747);
and U8821 (N_8821,N_8691,N_8697);
or U8822 (N_8822,N_8670,N_8716);
and U8823 (N_8823,N_8749,N_8663);
nor U8824 (N_8824,N_8682,N_8730);
and U8825 (N_8825,N_8720,N_8685);
or U8826 (N_8826,N_8740,N_8671);
xor U8827 (N_8827,N_8729,N_8631);
xor U8828 (N_8828,N_8743,N_8638);
nor U8829 (N_8829,N_8634,N_8642);
nor U8830 (N_8830,N_8674,N_8653);
xnor U8831 (N_8831,N_8744,N_8686);
nand U8832 (N_8832,N_8695,N_8675);
nand U8833 (N_8833,N_8742,N_8702);
nand U8834 (N_8834,N_8655,N_8649);
nand U8835 (N_8835,N_8691,N_8678);
and U8836 (N_8836,N_8740,N_8644);
nor U8837 (N_8837,N_8707,N_8639);
nand U8838 (N_8838,N_8693,N_8692);
nor U8839 (N_8839,N_8639,N_8679);
and U8840 (N_8840,N_8710,N_8666);
or U8841 (N_8841,N_8683,N_8651);
nand U8842 (N_8842,N_8700,N_8710);
nor U8843 (N_8843,N_8678,N_8715);
xnor U8844 (N_8844,N_8731,N_8672);
nor U8845 (N_8845,N_8691,N_8695);
nand U8846 (N_8846,N_8663,N_8641);
xnor U8847 (N_8847,N_8642,N_8653);
nor U8848 (N_8848,N_8639,N_8644);
or U8849 (N_8849,N_8733,N_8639);
xnor U8850 (N_8850,N_8685,N_8731);
nand U8851 (N_8851,N_8695,N_8657);
or U8852 (N_8852,N_8659,N_8688);
nor U8853 (N_8853,N_8700,N_8636);
xor U8854 (N_8854,N_8649,N_8628);
nand U8855 (N_8855,N_8638,N_8727);
nor U8856 (N_8856,N_8652,N_8637);
xor U8857 (N_8857,N_8697,N_8711);
xor U8858 (N_8858,N_8626,N_8738);
or U8859 (N_8859,N_8698,N_8669);
nand U8860 (N_8860,N_8746,N_8658);
or U8861 (N_8861,N_8686,N_8696);
xor U8862 (N_8862,N_8649,N_8699);
nand U8863 (N_8863,N_8675,N_8736);
nor U8864 (N_8864,N_8682,N_8639);
xor U8865 (N_8865,N_8675,N_8674);
or U8866 (N_8866,N_8629,N_8663);
and U8867 (N_8867,N_8630,N_8667);
xnor U8868 (N_8868,N_8697,N_8688);
and U8869 (N_8869,N_8653,N_8741);
or U8870 (N_8870,N_8649,N_8719);
and U8871 (N_8871,N_8740,N_8748);
nor U8872 (N_8872,N_8683,N_8625);
xor U8873 (N_8873,N_8657,N_8745);
and U8874 (N_8874,N_8635,N_8732);
xor U8875 (N_8875,N_8773,N_8835);
nor U8876 (N_8876,N_8849,N_8831);
xor U8877 (N_8877,N_8858,N_8846);
nor U8878 (N_8878,N_8832,N_8850);
nand U8879 (N_8879,N_8872,N_8784);
nand U8880 (N_8880,N_8761,N_8775);
nor U8881 (N_8881,N_8801,N_8787);
or U8882 (N_8882,N_8815,N_8799);
and U8883 (N_8883,N_8867,N_8809);
nand U8884 (N_8884,N_8844,N_8873);
nand U8885 (N_8885,N_8774,N_8821);
nand U8886 (N_8886,N_8834,N_8756);
and U8887 (N_8887,N_8788,N_8836);
xor U8888 (N_8888,N_8824,N_8818);
xor U8889 (N_8889,N_8804,N_8786);
and U8890 (N_8890,N_8793,N_8826);
or U8891 (N_8891,N_8862,N_8857);
xor U8892 (N_8892,N_8768,N_8816);
or U8893 (N_8893,N_8822,N_8842);
nand U8894 (N_8894,N_8767,N_8754);
and U8895 (N_8895,N_8874,N_8798);
nand U8896 (N_8896,N_8779,N_8763);
xnor U8897 (N_8897,N_8751,N_8833);
and U8898 (N_8898,N_8861,N_8807);
xnor U8899 (N_8899,N_8752,N_8845);
xnor U8900 (N_8900,N_8771,N_8762);
nand U8901 (N_8901,N_8853,N_8764);
and U8902 (N_8902,N_8854,N_8847);
or U8903 (N_8903,N_8819,N_8828);
nand U8904 (N_8904,N_8813,N_8753);
and U8905 (N_8905,N_8795,N_8770);
xor U8906 (N_8906,N_8797,N_8755);
nor U8907 (N_8907,N_8800,N_8765);
nand U8908 (N_8908,N_8851,N_8805);
and U8909 (N_8909,N_8827,N_8808);
xor U8910 (N_8910,N_8812,N_8869);
nor U8911 (N_8911,N_8790,N_8780);
and U8912 (N_8912,N_8806,N_8823);
nand U8913 (N_8913,N_8766,N_8863);
xor U8914 (N_8914,N_8814,N_8759);
xnor U8915 (N_8915,N_8777,N_8803);
or U8916 (N_8916,N_8852,N_8829);
or U8917 (N_8917,N_8838,N_8782);
and U8918 (N_8918,N_8791,N_8825);
nor U8919 (N_8919,N_8839,N_8785);
xor U8920 (N_8920,N_8859,N_8792);
xor U8921 (N_8921,N_8865,N_8830);
or U8922 (N_8922,N_8781,N_8840);
nor U8923 (N_8923,N_8864,N_8796);
nand U8924 (N_8924,N_8841,N_8760);
xnor U8925 (N_8925,N_8750,N_8776);
or U8926 (N_8926,N_8843,N_8860);
nor U8927 (N_8927,N_8837,N_8802);
and U8928 (N_8928,N_8817,N_8866);
xnor U8929 (N_8929,N_8811,N_8810);
nor U8930 (N_8930,N_8769,N_8868);
and U8931 (N_8931,N_8783,N_8757);
nand U8932 (N_8932,N_8772,N_8758);
nor U8933 (N_8933,N_8855,N_8789);
and U8934 (N_8934,N_8871,N_8848);
xor U8935 (N_8935,N_8794,N_8870);
nand U8936 (N_8936,N_8856,N_8778);
xnor U8937 (N_8937,N_8820,N_8781);
or U8938 (N_8938,N_8813,N_8804);
and U8939 (N_8939,N_8772,N_8849);
nand U8940 (N_8940,N_8775,N_8871);
and U8941 (N_8941,N_8869,N_8759);
nand U8942 (N_8942,N_8821,N_8804);
nand U8943 (N_8943,N_8759,N_8832);
nand U8944 (N_8944,N_8758,N_8865);
nand U8945 (N_8945,N_8759,N_8754);
nor U8946 (N_8946,N_8858,N_8867);
xnor U8947 (N_8947,N_8839,N_8840);
nor U8948 (N_8948,N_8831,N_8860);
and U8949 (N_8949,N_8833,N_8770);
and U8950 (N_8950,N_8750,N_8835);
and U8951 (N_8951,N_8758,N_8762);
nor U8952 (N_8952,N_8836,N_8821);
or U8953 (N_8953,N_8803,N_8779);
nor U8954 (N_8954,N_8808,N_8764);
or U8955 (N_8955,N_8796,N_8782);
or U8956 (N_8956,N_8818,N_8768);
nand U8957 (N_8957,N_8860,N_8871);
nor U8958 (N_8958,N_8814,N_8811);
xnor U8959 (N_8959,N_8848,N_8810);
nand U8960 (N_8960,N_8777,N_8762);
or U8961 (N_8961,N_8797,N_8761);
xor U8962 (N_8962,N_8824,N_8794);
and U8963 (N_8963,N_8766,N_8762);
nand U8964 (N_8964,N_8791,N_8796);
xnor U8965 (N_8965,N_8754,N_8855);
nand U8966 (N_8966,N_8783,N_8771);
nor U8967 (N_8967,N_8817,N_8800);
or U8968 (N_8968,N_8852,N_8799);
nand U8969 (N_8969,N_8750,N_8768);
nor U8970 (N_8970,N_8841,N_8818);
nand U8971 (N_8971,N_8835,N_8823);
nand U8972 (N_8972,N_8825,N_8829);
or U8973 (N_8973,N_8851,N_8788);
nor U8974 (N_8974,N_8804,N_8765);
xnor U8975 (N_8975,N_8839,N_8850);
nor U8976 (N_8976,N_8764,N_8824);
or U8977 (N_8977,N_8795,N_8850);
and U8978 (N_8978,N_8849,N_8795);
nor U8979 (N_8979,N_8783,N_8766);
or U8980 (N_8980,N_8849,N_8774);
and U8981 (N_8981,N_8806,N_8758);
nor U8982 (N_8982,N_8784,N_8854);
or U8983 (N_8983,N_8808,N_8867);
xor U8984 (N_8984,N_8841,N_8791);
nor U8985 (N_8985,N_8841,N_8769);
nor U8986 (N_8986,N_8812,N_8828);
or U8987 (N_8987,N_8782,N_8764);
or U8988 (N_8988,N_8841,N_8763);
nor U8989 (N_8989,N_8754,N_8751);
nand U8990 (N_8990,N_8754,N_8779);
or U8991 (N_8991,N_8810,N_8849);
xnor U8992 (N_8992,N_8826,N_8841);
nand U8993 (N_8993,N_8826,N_8847);
nor U8994 (N_8994,N_8776,N_8769);
xnor U8995 (N_8995,N_8800,N_8828);
nand U8996 (N_8996,N_8758,N_8814);
xnor U8997 (N_8997,N_8759,N_8862);
nor U8998 (N_8998,N_8791,N_8776);
xnor U8999 (N_8999,N_8753,N_8814);
nand U9000 (N_9000,N_8971,N_8913);
and U9001 (N_9001,N_8999,N_8894);
and U9002 (N_9002,N_8979,N_8990);
and U9003 (N_9003,N_8937,N_8970);
nor U9004 (N_9004,N_8928,N_8958);
or U9005 (N_9005,N_8886,N_8930);
and U9006 (N_9006,N_8939,N_8967);
nand U9007 (N_9007,N_8916,N_8993);
or U9008 (N_9008,N_8922,N_8942);
nand U9009 (N_9009,N_8956,N_8925);
and U9010 (N_9010,N_8936,N_8895);
or U9011 (N_9011,N_8963,N_8888);
xnor U9012 (N_9012,N_8906,N_8978);
nor U9013 (N_9013,N_8950,N_8884);
nor U9014 (N_9014,N_8910,N_8951);
xnor U9015 (N_9015,N_8982,N_8989);
or U9016 (N_9016,N_8965,N_8880);
nor U9017 (N_9017,N_8974,N_8915);
and U9018 (N_9018,N_8875,N_8988);
nor U9019 (N_9019,N_8986,N_8980);
nor U9020 (N_9020,N_8977,N_8998);
or U9021 (N_9021,N_8900,N_8997);
nand U9022 (N_9022,N_8995,N_8973);
nand U9023 (N_9023,N_8972,N_8934);
nand U9024 (N_9024,N_8949,N_8952);
nor U9025 (N_9025,N_8892,N_8896);
xnor U9026 (N_9026,N_8948,N_8898);
xnor U9027 (N_9027,N_8943,N_8897);
nand U9028 (N_9028,N_8953,N_8935);
nor U9029 (N_9029,N_8878,N_8926);
xnor U9030 (N_9030,N_8923,N_8908);
nand U9031 (N_9031,N_8946,N_8904);
xnor U9032 (N_9032,N_8938,N_8921);
nor U9033 (N_9033,N_8924,N_8891);
or U9034 (N_9034,N_8899,N_8905);
and U9035 (N_9035,N_8994,N_8941);
xor U9036 (N_9036,N_8889,N_8885);
nand U9037 (N_9037,N_8945,N_8890);
or U9038 (N_9038,N_8929,N_8976);
nand U9039 (N_9039,N_8918,N_8968);
nor U9040 (N_9040,N_8883,N_8893);
nand U9041 (N_9041,N_8887,N_8933);
and U9042 (N_9042,N_8919,N_8944);
or U9043 (N_9043,N_8907,N_8912);
nand U9044 (N_9044,N_8920,N_8882);
nor U9045 (N_9045,N_8983,N_8959);
xnor U9046 (N_9046,N_8955,N_8992);
nor U9047 (N_9047,N_8984,N_8940);
or U9048 (N_9048,N_8957,N_8996);
nand U9049 (N_9049,N_8947,N_8876);
nand U9050 (N_9050,N_8966,N_8991);
xnor U9051 (N_9051,N_8969,N_8909);
nor U9052 (N_9052,N_8962,N_8954);
or U9053 (N_9053,N_8975,N_8960);
xor U9054 (N_9054,N_8987,N_8917);
and U9055 (N_9055,N_8964,N_8881);
nand U9056 (N_9056,N_8981,N_8877);
or U9057 (N_9057,N_8901,N_8927);
nor U9058 (N_9058,N_8879,N_8903);
xor U9059 (N_9059,N_8961,N_8902);
or U9060 (N_9060,N_8932,N_8931);
or U9061 (N_9061,N_8914,N_8985);
or U9062 (N_9062,N_8911,N_8965);
nor U9063 (N_9063,N_8879,N_8924);
or U9064 (N_9064,N_8903,N_8960);
and U9065 (N_9065,N_8981,N_8925);
and U9066 (N_9066,N_8915,N_8899);
nor U9067 (N_9067,N_8975,N_8993);
nor U9068 (N_9068,N_8900,N_8985);
nand U9069 (N_9069,N_8974,N_8963);
nor U9070 (N_9070,N_8966,N_8970);
nor U9071 (N_9071,N_8917,N_8906);
nand U9072 (N_9072,N_8911,N_8927);
nor U9073 (N_9073,N_8938,N_8882);
xnor U9074 (N_9074,N_8961,N_8955);
nor U9075 (N_9075,N_8990,N_8962);
nor U9076 (N_9076,N_8959,N_8921);
and U9077 (N_9077,N_8896,N_8910);
and U9078 (N_9078,N_8949,N_8946);
or U9079 (N_9079,N_8905,N_8972);
or U9080 (N_9080,N_8988,N_8904);
xor U9081 (N_9081,N_8989,N_8935);
xor U9082 (N_9082,N_8958,N_8917);
nor U9083 (N_9083,N_8939,N_8956);
or U9084 (N_9084,N_8947,N_8954);
or U9085 (N_9085,N_8925,N_8970);
nand U9086 (N_9086,N_8977,N_8908);
and U9087 (N_9087,N_8939,N_8920);
and U9088 (N_9088,N_8998,N_8936);
and U9089 (N_9089,N_8956,N_8884);
and U9090 (N_9090,N_8906,N_8918);
and U9091 (N_9091,N_8980,N_8975);
xnor U9092 (N_9092,N_8884,N_8901);
and U9093 (N_9093,N_8990,N_8952);
nor U9094 (N_9094,N_8984,N_8986);
xor U9095 (N_9095,N_8922,N_8956);
xor U9096 (N_9096,N_8890,N_8952);
and U9097 (N_9097,N_8981,N_8885);
xor U9098 (N_9098,N_8880,N_8910);
nand U9099 (N_9099,N_8880,N_8973);
xor U9100 (N_9100,N_8952,N_8969);
xnor U9101 (N_9101,N_8955,N_8924);
nand U9102 (N_9102,N_8914,N_8889);
or U9103 (N_9103,N_8898,N_8988);
nor U9104 (N_9104,N_8985,N_8899);
nand U9105 (N_9105,N_8926,N_8910);
xnor U9106 (N_9106,N_8997,N_8885);
or U9107 (N_9107,N_8981,N_8916);
or U9108 (N_9108,N_8985,N_8989);
nand U9109 (N_9109,N_8923,N_8899);
nand U9110 (N_9110,N_8913,N_8991);
nand U9111 (N_9111,N_8946,N_8920);
nand U9112 (N_9112,N_8973,N_8937);
or U9113 (N_9113,N_8982,N_8921);
xnor U9114 (N_9114,N_8958,N_8891);
nand U9115 (N_9115,N_8938,N_8991);
xnor U9116 (N_9116,N_8922,N_8937);
nand U9117 (N_9117,N_8925,N_8978);
and U9118 (N_9118,N_8915,N_8892);
nand U9119 (N_9119,N_8918,N_8915);
or U9120 (N_9120,N_8953,N_8926);
nand U9121 (N_9121,N_8943,N_8948);
and U9122 (N_9122,N_8928,N_8964);
or U9123 (N_9123,N_8984,N_8938);
nor U9124 (N_9124,N_8876,N_8917);
nand U9125 (N_9125,N_9069,N_9084);
xnor U9126 (N_9126,N_9067,N_9046);
nor U9127 (N_9127,N_9102,N_9068);
nor U9128 (N_9128,N_9017,N_9080);
xor U9129 (N_9129,N_9100,N_9072);
or U9130 (N_9130,N_9110,N_9105);
nand U9131 (N_9131,N_9076,N_9078);
nor U9132 (N_9132,N_9091,N_9036);
or U9133 (N_9133,N_9090,N_9118);
nor U9134 (N_9134,N_9044,N_9107);
nand U9135 (N_9135,N_9056,N_9075);
nor U9136 (N_9136,N_9094,N_9088);
nand U9137 (N_9137,N_9089,N_9025);
nor U9138 (N_9138,N_9016,N_9121);
or U9139 (N_9139,N_9104,N_9083);
and U9140 (N_9140,N_9002,N_9034);
nand U9141 (N_9141,N_9009,N_9101);
or U9142 (N_9142,N_9086,N_9081);
nor U9143 (N_9143,N_9049,N_9035);
or U9144 (N_9144,N_9023,N_9021);
or U9145 (N_9145,N_9029,N_9063);
and U9146 (N_9146,N_9064,N_9062);
or U9147 (N_9147,N_9116,N_9030);
xnor U9148 (N_9148,N_9115,N_9000);
nor U9149 (N_9149,N_9008,N_9111);
xor U9150 (N_9150,N_9113,N_9099);
or U9151 (N_9151,N_9006,N_9012);
nand U9152 (N_9152,N_9028,N_9092);
nor U9153 (N_9153,N_9114,N_9074);
nand U9154 (N_9154,N_9108,N_9082);
and U9155 (N_9155,N_9058,N_9013);
or U9156 (N_9156,N_9073,N_9117);
or U9157 (N_9157,N_9093,N_9098);
nor U9158 (N_9158,N_9026,N_9004);
and U9159 (N_9159,N_9060,N_9042);
xor U9160 (N_9160,N_9124,N_9031);
and U9161 (N_9161,N_9011,N_9096);
nor U9162 (N_9162,N_9014,N_9003);
nand U9163 (N_9163,N_9033,N_9005);
or U9164 (N_9164,N_9045,N_9055);
nand U9165 (N_9165,N_9057,N_9112);
xnor U9166 (N_9166,N_9070,N_9040);
and U9167 (N_9167,N_9097,N_9120);
or U9168 (N_9168,N_9054,N_9015);
nor U9169 (N_9169,N_9043,N_9103);
or U9170 (N_9170,N_9109,N_9032);
and U9171 (N_9171,N_9047,N_9059);
nor U9172 (N_9172,N_9041,N_9051);
or U9173 (N_9173,N_9053,N_9020);
xnor U9174 (N_9174,N_9039,N_9007);
nor U9175 (N_9175,N_9122,N_9066);
xnor U9176 (N_9176,N_9123,N_9079);
nand U9177 (N_9177,N_9001,N_9037);
nand U9178 (N_9178,N_9119,N_9052);
and U9179 (N_9179,N_9106,N_9050);
nand U9180 (N_9180,N_9077,N_9048);
and U9181 (N_9181,N_9024,N_9022);
or U9182 (N_9182,N_9010,N_9095);
xor U9183 (N_9183,N_9018,N_9087);
nand U9184 (N_9184,N_9019,N_9085);
xnor U9185 (N_9185,N_9027,N_9038);
and U9186 (N_9186,N_9071,N_9061);
xor U9187 (N_9187,N_9065,N_9046);
xor U9188 (N_9188,N_9018,N_9082);
xnor U9189 (N_9189,N_9068,N_9046);
or U9190 (N_9190,N_9078,N_9102);
nor U9191 (N_9191,N_9069,N_9108);
xor U9192 (N_9192,N_9035,N_9118);
nor U9193 (N_9193,N_9076,N_9081);
and U9194 (N_9194,N_9059,N_9088);
nand U9195 (N_9195,N_9116,N_9038);
xor U9196 (N_9196,N_9045,N_9075);
or U9197 (N_9197,N_9059,N_9018);
nand U9198 (N_9198,N_9044,N_9064);
xnor U9199 (N_9199,N_9098,N_9060);
nor U9200 (N_9200,N_9019,N_9060);
xor U9201 (N_9201,N_9098,N_9011);
nand U9202 (N_9202,N_9050,N_9079);
nor U9203 (N_9203,N_9064,N_9116);
xor U9204 (N_9204,N_9029,N_9018);
and U9205 (N_9205,N_9017,N_9067);
xor U9206 (N_9206,N_9015,N_9010);
xnor U9207 (N_9207,N_9124,N_9096);
and U9208 (N_9208,N_9078,N_9042);
or U9209 (N_9209,N_9064,N_9021);
nand U9210 (N_9210,N_9022,N_9014);
xor U9211 (N_9211,N_9120,N_9098);
nor U9212 (N_9212,N_9003,N_9031);
xor U9213 (N_9213,N_9122,N_9016);
or U9214 (N_9214,N_9005,N_9113);
or U9215 (N_9215,N_9032,N_9114);
nor U9216 (N_9216,N_9072,N_9075);
xnor U9217 (N_9217,N_9013,N_9088);
and U9218 (N_9218,N_9057,N_9007);
nor U9219 (N_9219,N_9088,N_9057);
and U9220 (N_9220,N_9020,N_9069);
nand U9221 (N_9221,N_9015,N_9116);
nand U9222 (N_9222,N_9017,N_9098);
nand U9223 (N_9223,N_9099,N_9098);
and U9224 (N_9224,N_9106,N_9051);
xnor U9225 (N_9225,N_9040,N_9098);
nor U9226 (N_9226,N_9027,N_9046);
nand U9227 (N_9227,N_9012,N_9099);
and U9228 (N_9228,N_9059,N_9120);
and U9229 (N_9229,N_9124,N_9043);
nor U9230 (N_9230,N_9114,N_9041);
and U9231 (N_9231,N_9004,N_9095);
nor U9232 (N_9232,N_9058,N_9043);
xor U9233 (N_9233,N_9008,N_9002);
and U9234 (N_9234,N_9055,N_9081);
nand U9235 (N_9235,N_9054,N_9014);
nor U9236 (N_9236,N_9024,N_9063);
and U9237 (N_9237,N_9075,N_9010);
and U9238 (N_9238,N_9106,N_9006);
and U9239 (N_9239,N_9041,N_9091);
nor U9240 (N_9240,N_9012,N_9078);
nor U9241 (N_9241,N_9028,N_9026);
xor U9242 (N_9242,N_9015,N_9094);
xor U9243 (N_9243,N_9045,N_9065);
nand U9244 (N_9244,N_9120,N_9039);
nand U9245 (N_9245,N_9033,N_9118);
nand U9246 (N_9246,N_9010,N_9028);
xor U9247 (N_9247,N_9016,N_9064);
and U9248 (N_9248,N_9110,N_9011);
xnor U9249 (N_9249,N_9063,N_9089);
xnor U9250 (N_9250,N_9244,N_9170);
or U9251 (N_9251,N_9168,N_9203);
nand U9252 (N_9252,N_9177,N_9211);
or U9253 (N_9253,N_9241,N_9149);
nand U9254 (N_9254,N_9141,N_9146);
and U9255 (N_9255,N_9201,N_9166);
xnor U9256 (N_9256,N_9179,N_9212);
nand U9257 (N_9257,N_9202,N_9216);
and U9258 (N_9258,N_9152,N_9140);
nand U9259 (N_9259,N_9249,N_9199);
and U9260 (N_9260,N_9136,N_9198);
nor U9261 (N_9261,N_9157,N_9171);
and U9262 (N_9262,N_9222,N_9173);
nor U9263 (N_9263,N_9151,N_9220);
and U9264 (N_9264,N_9169,N_9224);
xor U9265 (N_9265,N_9207,N_9176);
or U9266 (N_9266,N_9126,N_9232);
and U9267 (N_9267,N_9234,N_9188);
nor U9268 (N_9268,N_9229,N_9191);
nor U9269 (N_9269,N_9133,N_9180);
and U9270 (N_9270,N_9150,N_9143);
or U9271 (N_9271,N_9162,N_9164);
xnor U9272 (N_9272,N_9245,N_9239);
and U9273 (N_9273,N_9206,N_9225);
nand U9274 (N_9274,N_9125,N_9129);
or U9275 (N_9275,N_9155,N_9238);
nor U9276 (N_9276,N_9167,N_9236);
or U9277 (N_9277,N_9217,N_9196);
xor U9278 (N_9278,N_9138,N_9134);
and U9279 (N_9279,N_9161,N_9130);
or U9280 (N_9280,N_9205,N_9128);
nand U9281 (N_9281,N_9156,N_9227);
nor U9282 (N_9282,N_9213,N_9139);
and U9283 (N_9283,N_9178,N_9131);
xor U9284 (N_9284,N_9237,N_9208);
and U9285 (N_9285,N_9153,N_9228);
xor U9286 (N_9286,N_9223,N_9159);
or U9287 (N_9287,N_9235,N_9174);
nand U9288 (N_9288,N_9219,N_9186);
or U9289 (N_9289,N_9172,N_9137);
or U9290 (N_9290,N_9243,N_9194);
and U9291 (N_9291,N_9189,N_9147);
or U9292 (N_9292,N_9165,N_9175);
or U9293 (N_9293,N_9145,N_9190);
or U9294 (N_9294,N_9158,N_9248);
xor U9295 (N_9295,N_9160,N_9184);
xor U9296 (N_9296,N_9233,N_9221);
xor U9297 (N_9297,N_9154,N_9163);
nor U9298 (N_9298,N_9148,N_9209);
xor U9299 (N_9299,N_9187,N_9181);
and U9300 (N_9300,N_9142,N_9192);
nand U9301 (N_9301,N_9204,N_9183);
xnor U9302 (N_9302,N_9200,N_9215);
and U9303 (N_9303,N_9214,N_9135);
or U9304 (N_9304,N_9182,N_9193);
xor U9305 (N_9305,N_9230,N_9247);
nor U9306 (N_9306,N_9231,N_9218);
xor U9307 (N_9307,N_9185,N_9240);
or U9308 (N_9308,N_9246,N_9195);
nand U9309 (N_9309,N_9127,N_9132);
nor U9310 (N_9310,N_9144,N_9210);
or U9311 (N_9311,N_9197,N_9226);
xor U9312 (N_9312,N_9242,N_9182);
or U9313 (N_9313,N_9186,N_9208);
nand U9314 (N_9314,N_9178,N_9175);
and U9315 (N_9315,N_9247,N_9185);
and U9316 (N_9316,N_9235,N_9200);
and U9317 (N_9317,N_9237,N_9210);
and U9318 (N_9318,N_9198,N_9162);
or U9319 (N_9319,N_9224,N_9232);
nor U9320 (N_9320,N_9189,N_9206);
xnor U9321 (N_9321,N_9142,N_9187);
and U9322 (N_9322,N_9183,N_9135);
nand U9323 (N_9323,N_9197,N_9246);
and U9324 (N_9324,N_9173,N_9165);
nand U9325 (N_9325,N_9172,N_9219);
nor U9326 (N_9326,N_9178,N_9236);
nand U9327 (N_9327,N_9179,N_9203);
or U9328 (N_9328,N_9175,N_9243);
nand U9329 (N_9329,N_9156,N_9183);
or U9330 (N_9330,N_9215,N_9146);
nand U9331 (N_9331,N_9189,N_9134);
and U9332 (N_9332,N_9190,N_9131);
nand U9333 (N_9333,N_9131,N_9242);
nor U9334 (N_9334,N_9149,N_9217);
xor U9335 (N_9335,N_9168,N_9207);
nand U9336 (N_9336,N_9140,N_9182);
xnor U9337 (N_9337,N_9167,N_9210);
nand U9338 (N_9338,N_9147,N_9174);
nor U9339 (N_9339,N_9159,N_9152);
and U9340 (N_9340,N_9205,N_9129);
nor U9341 (N_9341,N_9215,N_9140);
and U9342 (N_9342,N_9126,N_9206);
nand U9343 (N_9343,N_9147,N_9178);
nand U9344 (N_9344,N_9206,N_9125);
nand U9345 (N_9345,N_9150,N_9184);
xnor U9346 (N_9346,N_9129,N_9226);
nor U9347 (N_9347,N_9204,N_9158);
nor U9348 (N_9348,N_9167,N_9221);
and U9349 (N_9349,N_9214,N_9228);
nor U9350 (N_9350,N_9185,N_9136);
or U9351 (N_9351,N_9219,N_9152);
and U9352 (N_9352,N_9225,N_9148);
and U9353 (N_9353,N_9205,N_9198);
nor U9354 (N_9354,N_9191,N_9213);
and U9355 (N_9355,N_9202,N_9172);
nand U9356 (N_9356,N_9211,N_9144);
or U9357 (N_9357,N_9233,N_9158);
and U9358 (N_9358,N_9195,N_9174);
nor U9359 (N_9359,N_9211,N_9174);
nor U9360 (N_9360,N_9224,N_9190);
or U9361 (N_9361,N_9135,N_9189);
nor U9362 (N_9362,N_9171,N_9146);
and U9363 (N_9363,N_9247,N_9162);
nand U9364 (N_9364,N_9217,N_9243);
and U9365 (N_9365,N_9207,N_9183);
nor U9366 (N_9366,N_9197,N_9146);
and U9367 (N_9367,N_9141,N_9144);
nor U9368 (N_9368,N_9182,N_9198);
xnor U9369 (N_9369,N_9161,N_9201);
and U9370 (N_9370,N_9176,N_9245);
nand U9371 (N_9371,N_9201,N_9184);
nand U9372 (N_9372,N_9137,N_9245);
xor U9373 (N_9373,N_9180,N_9204);
or U9374 (N_9374,N_9187,N_9135);
nand U9375 (N_9375,N_9313,N_9251);
or U9376 (N_9376,N_9373,N_9324);
and U9377 (N_9377,N_9300,N_9332);
xor U9378 (N_9378,N_9342,N_9357);
nor U9379 (N_9379,N_9295,N_9368);
nand U9380 (N_9380,N_9296,N_9364);
xnor U9381 (N_9381,N_9270,N_9283);
and U9382 (N_9382,N_9292,N_9358);
nor U9383 (N_9383,N_9258,N_9322);
nand U9384 (N_9384,N_9359,N_9309);
and U9385 (N_9385,N_9325,N_9282);
and U9386 (N_9386,N_9260,N_9250);
xnor U9387 (N_9387,N_9262,N_9297);
xor U9388 (N_9388,N_9356,N_9290);
nor U9389 (N_9389,N_9326,N_9320);
xnor U9390 (N_9390,N_9321,N_9365);
nor U9391 (N_9391,N_9318,N_9288);
or U9392 (N_9392,N_9298,N_9311);
nor U9393 (N_9393,N_9354,N_9317);
nor U9394 (N_9394,N_9286,N_9316);
xor U9395 (N_9395,N_9348,N_9355);
nor U9396 (N_9396,N_9363,N_9315);
xor U9397 (N_9397,N_9362,N_9374);
and U9398 (N_9398,N_9310,N_9268);
and U9399 (N_9399,N_9337,N_9269);
nand U9400 (N_9400,N_9289,N_9312);
xnor U9401 (N_9401,N_9346,N_9265);
nor U9402 (N_9402,N_9344,N_9271);
and U9403 (N_9403,N_9284,N_9345);
nor U9404 (N_9404,N_9367,N_9254);
or U9405 (N_9405,N_9275,N_9366);
nor U9406 (N_9406,N_9261,N_9277);
xnor U9407 (N_9407,N_9305,N_9331);
and U9408 (N_9408,N_9336,N_9294);
nor U9409 (N_9409,N_9276,N_9329);
or U9410 (N_9410,N_9338,N_9293);
xnor U9411 (N_9411,N_9303,N_9343);
xor U9412 (N_9412,N_9350,N_9273);
and U9413 (N_9413,N_9352,N_9340);
xnor U9414 (N_9414,N_9301,N_9328);
nand U9415 (N_9415,N_9369,N_9274);
xor U9416 (N_9416,N_9266,N_9361);
nand U9417 (N_9417,N_9333,N_9285);
or U9418 (N_9418,N_9279,N_9308);
or U9419 (N_9419,N_9272,N_9255);
xor U9420 (N_9420,N_9370,N_9259);
xnor U9421 (N_9421,N_9319,N_9252);
xnor U9422 (N_9422,N_9327,N_9304);
xnor U9423 (N_9423,N_9371,N_9341);
or U9424 (N_9424,N_9263,N_9339);
nand U9425 (N_9425,N_9347,N_9349);
nand U9426 (N_9426,N_9302,N_9264);
nor U9427 (N_9427,N_9306,N_9257);
nor U9428 (N_9428,N_9287,N_9281);
nor U9429 (N_9429,N_9267,N_9372);
xor U9430 (N_9430,N_9256,N_9299);
or U9431 (N_9431,N_9360,N_9330);
nand U9432 (N_9432,N_9334,N_9353);
nand U9433 (N_9433,N_9323,N_9291);
xnor U9434 (N_9434,N_9335,N_9278);
and U9435 (N_9435,N_9307,N_9314);
and U9436 (N_9436,N_9280,N_9351);
nand U9437 (N_9437,N_9253,N_9347);
xnor U9438 (N_9438,N_9279,N_9261);
and U9439 (N_9439,N_9271,N_9257);
nor U9440 (N_9440,N_9287,N_9267);
xnor U9441 (N_9441,N_9327,N_9367);
or U9442 (N_9442,N_9330,N_9349);
and U9443 (N_9443,N_9286,N_9257);
and U9444 (N_9444,N_9322,N_9320);
and U9445 (N_9445,N_9293,N_9365);
nor U9446 (N_9446,N_9265,N_9355);
and U9447 (N_9447,N_9326,N_9344);
nand U9448 (N_9448,N_9286,N_9305);
nand U9449 (N_9449,N_9364,N_9336);
nand U9450 (N_9450,N_9299,N_9315);
or U9451 (N_9451,N_9288,N_9281);
xnor U9452 (N_9452,N_9271,N_9280);
or U9453 (N_9453,N_9325,N_9342);
nand U9454 (N_9454,N_9276,N_9308);
nor U9455 (N_9455,N_9370,N_9294);
xor U9456 (N_9456,N_9374,N_9360);
and U9457 (N_9457,N_9348,N_9275);
and U9458 (N_9458,N_9286,N_9307);
and U9459 (N_9459,N_9254,N_9338);
nand U9460 (N_9460,N_9332,N_9311);
nor U9461 (N_9461,N_9300,N_9366);
and U9462 (N_9462,N_9350,N_9364);
xor U9463 (N_9463,N_9354,N_9329);
or U9464 (N_9464,N_9310,N_9311);
nor U9465 (N_9465,N_9370,N_9341);
nand U9466 (N_9466,N_9311,N_9352);
or U9467 (N_9467,N_9285,N_9284);
or U9468 (N_9468,N_9299,N_9259);
or U9469 (N_9469,N_9270,N_9268);
and U9470 (N_9470,N_9357,N_9292);
or U9471 (N_9471,N_9268,N_9324);
and U9472 (N_9472,N_9270,N_9287);
or U9473 (N_9473,N_9354,N_9331);
and U9474 (N_9474,N_9265,N_9357);
and U9475 (N_9475,N_9338,N_9362);
or U9476 (N_9476,N_9365,N_9333);
and U9477 (N_9477,N_9301,N_9302);
and U9478 (N_9478,N_9283,N_9323);
and U9479 (N_9479,N_9307,N_9265);
nor U9480 (N_9480,N_9282,N_9268);
nand U9481 (N_9481,N_9323,N_9319);
or U9482 (N_9482,N_9276,N_9330);
nor U9483 (N_9483,N_9257,N_9373);
xnor U9484 (N_9484,N_9368,N_9294);
or U9485 (N_9485,N_9370,N_9301);
and U9486 (N_9486,N_9349,N_9288);
nand U9487 (N_9487,N_9312,N_9255);
nand U9488 (N_9488,N_9265,N_9264);
nand U9489 (N_9489,N_9333,N_9252);
and U9490 (N_9490,N_9344,N_9307);
and U9491 (N_9491,N_9313,N_9353);
or U9492 (N_9492,N_9346,N_9352);
and U9493 (N_9493,N_9298,N_9371);
or U9494 (N_9494,N_9292,N_9294);
nand U9495 (N_9495,N_9371,N_9352);
nand U9496 (N_9496,N_9265,N_9335);
xnor U9497 (N_9497,N_9278,N_9363);
or U9498 (N_9498,N_9315,N_9285);
nor U9499 (N_9499,N_9364,N_9361);
xnor U9500 (N_9500,N_9465,N_9479);
or U9501 (N_9501,N_9400,N_9386);
xnor U9502 (N_9502,N_9383,N_9435);
nor U9503 (N_9503,N_9451,N_9422);
or U9504 (N_9504,N_9375,N_9411);
and U9505 (N_9505,N_9438,N_9396);
and U9506 (N_9506,N_9489,N_9409);
and U9507 (N_9507,N_9472,N_9379);
xnor U9508 (N_9508,N_9399,N_9495);
or U9509 (N_9509,N_9463,N_9486);
nand U9510 (N_9510,N_9420,N_9405);
nand U9511 (N_9511,N_9434,N_9401);
xor U9512 (N_9512,N_9397,N_9387);
nand U9513 (N_9513,N_9477,N_9490);
xor U9514 (N_9514,N_9398,N_9492);
xnor U9515 (N_9515,N_9458,N_9416);
or U9516 (N_9516,N_9494,N_9402);
nor U9517 (N_9517,N_9413,N_9454);
nand U9518 (N_9518,N_9480,N_9447);
xor U9519 (N_9519,N_9431,N_9470);
xor U9520 (N_9520,N_9432,N_9433);
nor U9521 (N_9521,N_9497,N_9437);
or U9522 (N_9522,N_9421,N_9448);
xor U9523 (N_9523,N_9436,N_9474);
and U9524 (N_9524,N_9429,N_9406);
or U9525 (N_9525,N_9461,N_9456);
or U9526 (N_9526,N_9446,N_9439);
nor U9527 (N_9527,N_9481,N_9393);
nor U9528 (N_9528,N_9426,N_9493);
nor U9529 (N_9529,N_9441,N_9395);
or U9530 (N_9530,N_9430,N_9417);
xnor U9531 (N_9531,N_9491,N_9485);
xnor U9532 (N_9532,N_9462,N_9408);
xnor U9533 (N_9533,N_9415,N_9496);
nand U9534 (N_9534,N_9444,N_9414);
nor U9535 (N_9535,N_9403,N_9450);
nand U9536 (N_9536,N_9487,N_9455);
xnor U9537 (N_9537,N_9483,N_9424);
or U9538 (N_9538,N_9384,N_9380);
nand U9539 (N_9539,N_9428,N_9499);
and U9540 (N_9540,N_9442,N_9376);
nand U9541 (N_9541,N_9469,N_9466);
nor U9542 (N_9542,N_9418,N_9449);
and U9543 (N_9543,N_9457,N_9407);
nor U9544 (N_9544,N_9473,N_9460);
nand U9545 (N_9545,N_9391,N_9471);
or U9546 (N_9546,N_9475,N_9478);
and U9547 (N_9547,N_9381,N_9388);
or U9548 (N_9548,N_9453,N_9445);
or U9549 (N_9549,N_9378,N_9412);
and U9550 (N_9550,N_9392,N_9476);
nand U9551 (N_9551,N_9484,N_9443);
nor U9552 (N_9552,N_9382,N_9394);
nor U9553 (N_9553,N_9482,N_9452);
nand U9554 (N_9554,N_9488,N_9389);
and U9555 (N_9555,N_9498,N_9390);
and U9556 (N_9556,N_9419,N_9377);
and U9557 (N_9557,N_9459,N_9467);
or U9558 (N_9558,N_9468,N_9427);
nor U9559 (N_9559,N_9464,N_9410);
and U9560 (N_9560,N_9423,N_9385);
xor U9561 (N_9561,N_9440,N_9425);
and U9562 (N_9562,N_9404,N_9405);
and U9563 (N_9563,N_9388,N_9486);
nor U9564 (N_9564,N_9484,N_9418);
xnor U9565 (N_9565,N_9408,N_9478);
and U9566 (N_9566,N_9448,N_9485);
nor U9567 (N_9567,N_9484,N_9375);
and U9568 (N_9568,N_9398,N_9424);
and U9569 (N_9569,N_9479,N_9461);
or U9570 (N_9570,N_9497,N_9440);
xnor U9571 (N_9571,N_9424,N_9383);
nand U9572 (N_9572,N_9451,N_9400);
or U9573 (N_9573,N_9496,N_9498);
or U9574 (N_9574,N_9404,N_9388);
and U9575 (N_9575,N_9428,N_9466);
xnor U9576 (N_9576,N_9461,N_9405);
nor U9577 (N_9577,N_9491,N_9471);
xnor U9578 (N_9578,N_9401,N_9402);
nand U9579 (N_9579,N_9383,N_9392);
or U9580 (N_9580,N_9463,N_9390);
and U9581 (N_9581,N_9413,N_9493);
xnor U9582 (N_9582,N_9394,N_9459);
or U9583 (N_9583,N_9473,N_9377);
xor U9584 (N_9584,N_9462,N_9475);
and U9585 (N_9585,N_9495,N_9464);
xor U9586 (N_9586,N_9465,N_9443);
nand U9587 (N_9587,N_9457,N_9408);
xor U9588 (N_9588,N_9493,N_9432);
nor U9589 (N_9589,N_9467,N_9377);
nand U9590 (N_9590,N_9385,N_9449);
xnor U9591 (N_9591,N_9386,N_9378);
and U9592 (N_9592,N_9485,N_9393);
and U9593 (N_9593,N_9427,N_9422);
xnor U9594 (N_9594,N_9419,N_9401);
xnor U9595 (N_9595,N_9470,N_9490);
and U9596 (N_9596,N_9381,N_9448);
xnor U9597 (N_9597,N_9479,N_9471);
nand U9598 (N_9598,N_9488,N_9415);
nand U9599 (N_9599,N_9478,N_9379);
nor U9600 (N_9600,N_9492,N_9470);
nor U9601 (N_9601,N_9411,N_9427);
nor U9602 (N_9602,N_9475,N_9408);
xnor U9603 (N_9603,N_9424,N_9384);
or U9604 (N_9604,N_9408,N_9481);
and U9605 (N_9605,N_9471,N_9396);
and U9606 (N_9606,N_9451,N_9412);
xor U9607 (N_9607,N_9491,N_9481);
and U9608 (N_9608,N_9452,N_9493);
nand U9609 (N_9609,N_9378,N_9495);
and U9610 (N_9610,N_9448,N_9422);
and U9611 (N_9611,N_9390,N_9408);
nor U9612 (N_9612,N_9492,N_9463);
xor U9613 (N_9613,N_9396,N_9477);
xor U9614 (N_9614,N_9379,N_9398);
nor U9615 (N_9615,N_9437,N_9434);
xnor U9616 (N_9616,N_9447,N_9403);
nand U9617 (N_9617,N_9378,N_9464);
or U9618 (N_9618,N_9407,N_9444);
and U9619 (N_9619,N_9461,N_9409);
and U9620 (N_9620,N_9434,N_9438);
nand U9621 (N_9621,N_9466,N_9419);
or U9622 (N_9622,N_9431,N_9381);
nor U9623 (N_9623,N_9490,N_9411);
and U9624 (N_9624,N_9412,N_9443);
xnor U9625 (N_9625,N_9604,N_9599);
xnor U9626 (N_9626,N_9618,N_9501);
xor U9627 (N_9627,N_9548,N_9577);
and U9628 (N_9628,N_9612,N_9603);
nand U9629 (N_9629,N_9594,N_9587);
nor U9630 (N_9630,N_9579,N_9590);
nor U9631 (N_9631,N_9529,N_9609);
nand U9632 (N_9632,N_9586,N_9616);
nor U9633 (N_9633,N_9562,N_9520);
and U9634 (N_9634,N_9506,N_9543);
xnor U9635 (N_9635,N_9546,N_9555);
and U9636 (N_9636,N_9554,N_9611);
or U9637 (N_9637,N_9619,N_9600);
xor U9638 (N_9638,N_9513,N_9621);
nor U9639 (N_9639,N_9522,N_9544);
nor U9640 (N_9640,N_9623,N_9547);
nand U9641 (N_9641,N_9514,N_9568);
nor U9642 (N_9642,N_9518,N_9549);
xnor U9643 (N_9643,N_9596,N_9531);
xor U9644 (N_9644,N_9584,N_9620);
nor U9645 (N_9645,N_9569,N_9558);
nor U9646 (N_9646,N_9615,N_9589);
nor U9647 (N_9647,N_9508,N_9610);
nand U9648 (N_9648,N_9578,N_9606);
xor U9649 (N_9649,N_9510,N_9504);
xnor U9650 (N_9650,N_9527,N_9500);
or U9651 (N_9651,N_9605,N_9571);
nor U9652 (N_9652,N_9567,N_9515);
or U9653 (N_9653,N_9585,N_9557);
nand U9654 (N_9654,N_9521,N_9614);
nor U9655 (N_9655,N_9519,N_9607);
xnor U9656 (N_9656,N_9535,N_9541);
xor U9657 (N_9657,N_9502,N_9553);
or U9658 (N_9658,N_9503,N_9572);
nor U9659 (N_9659,N_9574,N_9517);
nand U9660 (N_9660,N_9564,N_9566);
or U9661 (N_9661,N_9511,N_9561);
nand U9662 (N_9662,N_9598,N_9552);
or U9663 (N_9663,N_9560,N_9582);
and U9664 (N_9664,N_9538,N_9534);
or U9665 (N_9665,N_9575,N_9581);
or U9666 (N_9666,N_9542,N_9576);
and U9667 (N_9667,N_9595,N_9556);
xor U9668 (N_9668,N_9617,N_9525);
or U9669 (N_9669,N_9540,N_9622);
nand U9670 (N_9670,N_9536,N_9509);
or U9671 (N_9671,N_9597,N_9583);
and U9672 (N_9672,N_9613,N_9533);
nor U9673 (N_9673,N_9516,N_9505);
and U9674 (N_9674,N_9539,N_9523);
xor U9675 (N_9675,N_9602,N_9532);
or U9676 (N_9676,N_9570,N_9545);
nor U9677 (N_9677,N_9563,N_9537);
and U9678 (N_9678,N_9526,N_9524);
xnor U9679 (N_9679,N_9565,N_9573);
xnor U9680 (N_9680,N_9593,N_9530);
or U9681 (N_9681,N_9624,N_9592);
and U9682 (N_9682,N_9580,N_9588);
nor U9683 (N_9683,N_9550,N_9591);
nand U9684 (N_9684,N_9528,N_9507);
and U9685 (N_9685,N_9512,N_9551);
or U9686 (N_9686,N_9608,N_9559);
and U9687 (N_9687,N_9601,N_9592);
xnor U9688 (N_9688,N_9547,N_9510);
nand U9689 (N_9689,N_9504,N_9585);
and U9690 (N_9690,N_9622,N_9527);
or U9691 (N_9691,N_9524,N_9533);
and U9692 (N_9692,N_9619,N_9542);
nand U9693 (N_9693,N_9620,N_9581);
xor U9694 (N_9694,N_9601,N_9507);
nor U9695 (N_9695,N_9573,N_9512);
xor U9696 (N_9696,N_9588,N_9564);
nor U9697 (N_9697,N_9565,N_9587);
and U9698 (N_9698,N_9601,N_9555);
and U9699 (N_9699,N_9558,N_9573);
or U9700 (N_9700,N_9503,N_9597);
nand U9701 (N_9701,N_9597,N_9515);
nor U9702 (N_9702,N_9523,N_9549);
nand U9703 (N_9703,N_9500,N_9555);
nor U9704 (N_9704,N_9571,N_9522);
or U9705 (N_9705,N_9604,N_9574);
nand U9706 (N_9706,N_9573,N_9539);
nand U9707 (N_9707,N_9561,N_9573);
or U9708 (N_9708,N_9508,N_9505);
or U9709 (N_9709,N_9546,N_9620);
or U9710 (N_9710,N_9582,N_9557);
xnor U9711 (N_9711,N_9525,N_9502);
nand U9712 (N_9712,N_9573,N_9621);
xor U9713 (N_9713,N_9504,N_9531);
or U9714 (N_9714,N_9624,N_9548);
xnor U9715 (N_9715,N_9547,N_9505);
and U9716 (N_9716,N_9539,N_9565);
nor U9717 (N_9717,N_9592,N_9530);
xnor U9718 (N_9718,N_9516,N_9535);
and U9719 (N_9719,N_9594,N_9610);
or U9720 (N_9720,N_9509,N_9591);
nor U9721 (N_9721,N_9608,N_9540);
or U9722 (N_9722,N_9503,N_9517);
and U9723 (N_9723,N_9621,N_9619);
nor U9724 (N_9724,N_9571,N_9500);
nor U9725 (N_9725,N_9590,N_9525);
or U9726 (N_9726,N_9539,N_9536);
or U9727 (N_9727,N_9517,N_9580);
or U9728 (N_9728,N_9595,N_9592);
nand U9729 (N_9729,N_9596,N_9564);
or U9730 (N_9730,N_9536,N_9568);
nand U9731 (N_9731,N_9570,N_9515);
nor U9732 (N_9732,N_9606,N_9604);
nand U9733 (N_9733,N_9624,N_9528);
and U9734 (N_9734,N_9541,N_9507);
nor U9735 (N_9735,N_9577,N_9621);
nor U9736 (N_9736,N_9570,N_9605);
xor U9737 (N_9737,N_9618,N_9619);
nor U9738 (N_9738,N_9516,N_9558);
nor U9739 (N_9739,N_9612,N_9523);
xor U9740 (N_9740,N_9616,N_9529);
or U9741 (N_9741,N_9540,N_9500);
and U9742 (N_9742,N_9597,N_9507);
and U9743 (N_9743,N_9519,N_9507);
nor U9744 (N_9744,N_9599,N_9510);
nor U9745 (N_9745,N_9617,N_9586);
nand U9746 (N_9746,N_9530,N_9564);
or U9747 (N_9747,N_9501,N_9521);
nand U9748 (N_9748,N_9558,N_9580);
and U9749 (N_9749,N_9618,N_9595);
and U9750 (N_9750,N_9701,N_9726);
xor U9751 (N_9751,N_9749,N_9699);
nor U9752 (N_9752,N_9746,N_9707);
or U9753 (N_9753,N_9661,N_9677);
or U9754 (N_9754,N_9718,N_9671);
xnor U9755 (N_9755,N_9710,N_9630);
and U9756 (N_9756,N_9724,N_9649);
and U9757 (N_9757,N_9629,N_9712);
nor U9758 (N_9758,N_9682,N_9715);
and U9759 (N_9759,N_9665,N_9725);
xnor U9760 (N_9760,N_9678,N_9738);
and U9761 (N_9761,N_9642,N_9662);
nor U9762 (N_9762,N_9713,N_9697);
nor U9763 (N_9763,N_9723,N_9741);
or U9764 (N_9764,N_9721,N_9733);
or U9765 (N_9765,N_9636,N_9643);
and U9766 (N_9766,N_9679,N_9628);
or U9767 (N_9767,N_9703,N_9654);
and U9768 (N_9768,N_9676,N_9748);
and U9769 (N_9769,N_9708,N_9651);
or U9770 (N_9770,N_9664,N_9637);
nand U9771 (N_9771,N_9706,N_9685);
nand U9772 (N_9772,N_9650,N_9625);
nand U9773 (N_9773,N_9694,N_9693);
or U9774 (N_9774,N_9666,N_9641);
or U9775 (N_9775,N_9732,N_9663);
nand U9776 (N_9776,N_9691,N_9696);
nor U9777 (N_9777,N_9742,N_9692);
xor U9778 (N_9778,N_9745,N_9744);
or U9779 (N_9779,N_9743,N_9669);
xor U9780 (N_9780,N_9705,N_9737);
xnor U9781 (N_9781,N_9645,N_9711);
nor U9782 (N_9782,N_9648,N_9735);
and U9783 (N_9783,N_9729,N_9722);
nor U9784 (N_9784,N_9670,N_9709);
or U9785 (N_9785,N_9673,N_9714);
xnor U9786 (N_9786,N_9631,N_9684);
xnor U9787 (N_9787,N_9655,N_9702);
nor U9788 (N_9788,N_9690,N_9652);
and U9789 (N_9789,N_9736,N_9638);
nand U9790 (N_9790,N_9634,N_9657);
nor U9791 (N_9791,N_9647,N_9626);
nand U9792 (N_9792,N_9720,N_9659);
or U9793 (N_9793,N_9717,N_9653);
xor U9794 (N_9794,N_9668,N_9672);
and U9795 (N_9795,N_9686,N_9727);
and U9796 (N_9796,N_9667,N_9739);
nor U9797 (N_9797,N_9704,N_9633);
nand U9798 (N_9798,N_9716,N_9728);
nand U9799 (N_9799,N_9687,N_9646);
nor U9800 (N_9800,N_9730,N_9639);
xor U9801 (N_9801,N_9740,N_9675);
and U9802 (N_9802,N_9644,N_9656);
nor U9803 (N_9803,N_9674,N_9658);
and U9804 (N_9804,N_9640,N_9695);
and U9805 (N_9805,N_9627,N_9689);
nor U9806 (N_9806,N_9734,N_9660);
and U9807 (N_9807,N_9700,N_9683);
nor U9808 (N_9808,N_9632,N_9719);
xor U9809 (N_9809,N_9635,N_9698);
nor U9810 (N_9810,N_9747,N_9680);
nor U9811 (N_9811,N_9681,N_9688);
and U9812 (N_9812,N_9731,N_9650);
nand U9813 (N_9813,N_9696,N_9730);
and U9814 (N_9814,N_9655,N_9653);
and U9815 (N_9815,N_9731,N_9696);
xor U9816 (N_9816,N_9725,N_9675);
or U9817 (N_9817,N_9683,N_9627);
nor U9818 (N_9818,N_9718,N_9716);
nand U9819 (N_9819,N_9653,N_9739);
and U9820 (N_9820,N_9698,N_9703);
or U9821 (N_9821,N_9734,N_9713);
nor U9822 (N_9822,N_9626,N_9700);
xnor U9823 (N_9823,N_9653,N_9663);
nor U9824 (N_9824,N_9653,N_9746);
or U9825 (N_9825,N_9708,N_9647);
or U9826 (N_9826,N_9645,N_9732);
and U9827 (N_9827,N_9663,N_9649);
nor U9828 (N_9828,N_9726,N_9670);
nor U9829 (N_9829,N_9702,N_9713);
or U9830 (N_9830,N_9713,N_9718);
or U9831 (N_9831,N_9743,N_9712);
xor U9832 (N_9832,N_9709,N_9696);
nand U9833 (N_9833,N_9702,N_9731);
or U9834 (N_9834,N_9643,N_9740);
xnor U9835 (N_9835,N_9630,N_9658);
or U9836 (N_9836,N_9630,N_9639);
nand U9837 (N_9837,N_9659,N_9637);
nor U9838 (N_9838,N_9732,N_9644);
xnor U9839 (N_9839,N_9646,N_9708);
or U9840 (N_9840,N_9733,N_9636);
xnor U9841 (N_9841,N_9693,N_9652);
xor U9842 (N_9842,N_9731,N_9673);
and U9843 (N_9843,N_9635,N_9651);
xor U9844 (N_9844,N_9669,N_9682);
or U9845 (N_9845,N_9653,N_9630);
nor U9846 (N_9846,N_9692,N_9709);
nor U9847 (N_9847,N_9682,N_9729);
xor U9848 (N_9848,N_9665,N_9728);
and U9849 (N_9849,N_9700,N_9702);
nand U9850 (N_9850,N_9629,N_9647);
xnor U9851 (N_9851,N_9675,N_9713);
nand U9852 (N_9852,N_9693,N_9699);
nor U9853 (N_9853,N_9710,N_9680);
and U9854 (N_9854,N_9676,N_9708);
or U9855 (N_9855,N_9723,N_9689);
nand U9856 (N_9856,N_9682,N_9704);
or U9857 (N_9857,N_9635,N_9662);
nand U9858 (N_9858,N_9693,N_9657);
xor U9859 (N_9859,N_9653,N_9641);
and U9860 (N_9860,N_9738,N_9734);
nor U9861 (N_9861,N_9685,N_9729);
xnor U9862 (N_9862,N_9728,N_9732);
nand U9863 (N_9863,N_9725,N_9731);
and U9864 (N_9864,N_9691,N_9667);
nor U9865 (N_9865,N_9645,N_9654);
or U9866 (N_9866,N_9704,N_9731);
nor U9867 (N_9867,N_9721,N_9720);
xor U9868 (N_9868,N_9683,N_9729);
nand U9869 (N_9869,N_9744,N_9700);
and U9870 (N_9870,N_9746,N_9628);
xor U9871 (N_9871,N_9696,N_9650);
nand U9872 (N_9872,N_9696,N_9699);
nor U9873 (N_9873,N_9671,N_9709);
nand U9874 (N_9874,N_9706,N_9719);
and U9875 (N_9875,N_9829,N_9764);
and U9876 (N_9876,N_9785,N_9778);
nor U9877 (N_9877,N_9750,N_9768);
nor U9878 (N_9878,N_9824,N_9855);
and U9879 (N_9879,N_9849,N_9852);
and U9880 (N_9880,N_9847,N_9751);
xor U9881 (N_9881,N_9822,N_9802);
or U9882 (N_9882,N_9873,N_9830);
or U9883 (N_9883,N_9866,N_9780);
nor U9884 (N_9884,N_9783,N_9801);
or U9885 (N_9885,N_9871,N_9781);
and U9886 (N_9886,N_9858,N_9752);
nand U9887 (N_9887,N_9777,N_9809);
nand U9888 (N_9888,N_9821,N_9825);
or U9889 (N_9889,N_9754,N_9812);
and U9890 (N_9890,N_9838,N_9857);
and U9891 (N_9891,N_9850,N_9846);
nor U9892 (N_9892,N_9795,N_9808);
nor U9893 (N_9893,N_9776,N_9782);
xor U9894 (N_9894,N_9842,N_9819);
or U9895 (N_9895,N_9772,N_9791);
nand U9896 (N_9896,N_9757,N_9870);
nand U9897 (N_9897,N_9820,N_9798);
xor U9898 (N_9898,N_9815,N_9839);
nor U9899 (N_9899,N_9771,N_9811);
or U9900 (N_9900,N_9787,N_9863);
and U9901 (N_9901,N_9859,N_9869);
and U9902 (N_9902,N_9853,N_9827);
or U9903 (N_9903,N_9845,N_9769);
nor U9904 (N_9904,N_9759,N_9800);
and U9905 (N_9905,N_9814,N_9861);
and U9906 (N_9906,N_9790,N_9799);
and U9907 (N_9907,N_9793,N_9753);
and U9908 (N_9908,N_9779,N_9837);
nand U9909 (N_9909,N_9774,N_9760);
and U9910 (N_9910,N_9756,N_9834);
and U9911 (N_9911,N_9796,N_9841);
or U9912 (N_9912,N_9810,N_9817);
or U9913 (N_9913,N_9864,N_9797);
or U9914 (N_9914,N_9851,N_9843);
and U9915 (N_9915,N_9868,N_9806);
nor U9916 (N_9916,N_9788,N_9818);
nor U9917 (N_9917,N_9775,N_9804);
xnor U9918 (N_9918,N_9833,N_9807);
xnor U9919 (N_9919,N_9835,N_9758);
nor U9920 (N_9920,N_9786,N_9826);
nand U9921 (N_9921,N_9766,N_9816);
xor U9922 (N_9922,N_9773,N_9836);
nor U9923 (N_9923,N_9867,N_9792);
and U9924 (N_9924,N_9840,N_9803);
nor U9925 (N_9925,N_9770,N_9805);
nand U9926 (N_9926,N_9874,N_9854);
and U9927 (N_9927,N_9862,N_9831);
xor U9928 (N_9928,N_9848,N_9761);
or U9929 (N_9929,N_9784,N_9789);
xnor U9930 (N_9930,N_9828,N_9767);
or U9931 (N_9931,N_9762,N_9813);
or U9932 (N_9932,N_9823,N_9794);
or U9933 (N_9933,N_9755,N_9844);
and U9934 (N_9934,N_9765,N_9856);
or U9935 (N_9935,N_9832,N_9860);
xnor U9936 (N_9936,N_9872,N_9865);
xor U9937 (N_9937,N_9763,N_9833);
and U9938 (N_9938,N_9817,N_9846);
or U9939 (N_9939,N_9801,N_9752);
nor U9940 (N_9940,N_9849,N_9758);
and U9941 (N_9941,N_9786,N_9793);
xnor U9942 (N_9942,N_9754,N_9848);
or U9943 (N_9943,N_9821,N_9843);
nand U9944 (N_9944,N_9823,N_9765);
or U9945 (N_9945,N_9835,N_9802);
nor U9946 (N_9946,N_9804,N_9834);
xnor U9947 (N_9947,N_9756,N_9841);
nand U9948 (N_9948,N_9852,N_9756);
xor U9949 (N_9949,N_9841,N_9795);
nor U9950 (N_9950,N_9773,N_9787);
xor U9951 (N_9951,N_9792,N_9793);
xor U9952 (N_9952,N_9766,N_9822);
nor U9953 (N_9953,N_9758,N_9799);
and U9954 (N_9954,N_9787,N_9755);
or U9955 (N_9955,N_9775,N_9832);
nor U9956 (N_9956,N_9844,N_9766);
nor U9957 (N_9957,N_9759,N_9858);
or U9958 (N_9958,N_9837,N_9826);
nand U9959 (N_9959,N_9862,N_9823);
or U9960 (N_9960,N_9831,N_9764);
nor U9961 (N_9961,N_9750,N_9818);
xnor U9962 (N_9962,N_9854,N_9785);
nand U9963 (N_9963,N_9752,N_9871);
xnor U9964 (N_9964,N_9860,N_9829);
and U9965 (N_9965,N_9836,N_9837);
xnor U9966 (N_9966,N_9785,N_9789);
nor U9967 (N_9967,N_9766,N_9752);
and U9968 (N_9968,N_9758,N_9808);
or U9969 (N_9969,N_9862,N_9767);
or U9970 (N_9970,N_9815,N_9780);
and U9971 (N_9971,N_9783,N_9770);
nand U9972 (N_9972,N_9786,N_9780);
and U9973 (N_9973,N_9824,N_9858);
xor U9974 (N_9974,N_9873,N_9799);
nand U9975 (N_9975,N_9788,N_9827);
and U9976 (N_9976,N_9848,N_9792);
nand U9977 (N_9977,N_9867,N_9755);
nor U9978 (N_9978,N_9776,N_9777);
nand U9979 (N_9979,N_9762,N_9848);
nand U9980 (N_9980,N_9857,N_9823);
nor U9981 (N_9981,N_9860,N_9855);
or U9982 (N_9982,N_9866,N_9840);
xnor U9983 (N_9983,N_9788,N_9808);
and U9984 (N_9984,N_9837,N_9843);
or U9985 (N_9985,N_9807,N_9770);
nor U9986 (N_9986,N_9794,N_9825);
xor U9987 (N_9987,N_9828,N_9849);
nor U9988 (N_9988,N_9782,N_9764);
xnor U9989 (N_9989,N_9850,N_9864);
or U9990 (N_9990,N_9764,N_9816);
nor U9991 (N_9991,N_9774,N_9808);
and U9992 (N_9992,N_9854,N_9863);
xnor U9993 (N_9993,N_9847,N_9778);
and U9994 (N_9994,N_9806,N_9833);
nor U9995 (N_9995,N_9755,N_9855);
nor U9996 (N_9996,N_9870,N_9841);
xnor U9997 (N_9997,N_9765,N_9869);
nor U9998 (N_9998,N_9812,N_9798);
and U9999 (N_9999,N_9760,N_9842);
and U10000 (N_10000,N_9886,N_9883);
nand U10001 (N_10001,N_9888,N_9922);
or U10002 (N_10002,N_9892,N_9992);
nor U10003 (N_10003,N_9944,N_9965);
nor U10004 (N_10004,N_9941,N_9942);
or U10005 (N_10005,N_9929,N_9917);
or U10006 (N_10006,N_9951,N_9936);
and U10007 (N_10007,N_9998,N_9899);
xnor U10008 (N_10008,N_9963,N_9981);
or U10009 (N_10009,N_9945,N_9916);
and U10010 (N_10010,N_9970,N_9926);
nand U10011 (N_10011,N_9960,N_9962);
xor U10012 (N_10012,N_9933,N_9972);
nor U10013 (N_10013,N_9993,N_9911);
nor U10014 (N_10014,N_9976,N_9928);
or U10015 (N_10015,N_9894,N_9907);
xnor U10016 (N_10016,N_9909,N_9905);
xor U10017 (N_10017,N_9947,N_9968);
or U10018 (N_10018,N_9983,N_9977);
and U10019 (N_10019,N_9914,N_9950);
nor U10020 (N_10020,N_9966,N_9915);
and U10021 (N_10021,N_9989,N_9994);
nor U10022 (N_10022,N_9953,N_9991);
xor U10023 (N_10023,N_9887,N_9997);
xor U10024 (N_10024,N_9974,N_9988);
or U10025 (N_10025,N_9878,N_9876);
or U10026 (N_10026,N_9875,N_9990);
and U10027 (N_10027,N_9967,N_9919);
and U10028 (N_10028,N_9898,N_9978);
xnor U10029 (N_10029,N_9987,N_9938);
or U10030 (N_10030,N_9900,N_9985);
and U10031 (N_10031,N_9920,N_9979);
nor U10032 (N_10032,N_9889,N_9903);
or U10033 (N_10033,N_9952,N_9999);
and U10034 (N_10034,N_9904,N_9996);
and U10035 (N_10035,N_9902,N_9946);
nand U10036 (N_10036,N_9956,N_9927);
and U10037 (N_10037,N_9884,N_9969);
nand U10038 (N_10038,N_9885,N_9908);
xnor U10039 (N_10039,N_9921,N_9975);
or U10040 (N_10040,N_9986,N_9877);
and U10041 (N_10041,N_9935,N_9939);
nand U10042 (N_10042,N_9943,N_9954);
nand U10043 (N_10043,N_9995,N_9913);
nor U10044 (N_10044,N_9958,N_9932);
nor U10045 (N_10045,N_9910,N_9973);
xnor U10046 (N_10046,N_9982,N_9971);
nor U10047 (N_10047,N_9964,N_9957);
nor U10048 (N_10048,N_9923,N_9980);
and U10049 (N_10049,N_9906,N_9882);
nand U10050 (N_10050,N_9879,N_9925);
xor U10051 (N_10051,N_9881,N_9891);
and U10052 (N_10052,N_9961,N_9893);
nand U10053 (N_10053,N_9937,N_9918);
and U10054 (N_10054,N_9930,N_9896);
or U10055 (N_10055,N_9880,N_9949);
and U10056 (N_10056,N_9959,N_9897);
nor U10057 (N_10057,N_9895,N_9924);
nor U10058 (N_10058,N_9948,N_9955);
or U10059 (N_10059,N_9890,N_9912);
or U10060 (N_10060,N_9984,N_9934);
and U10061 (N_10061,N_9901,N_9931);
and U10062 (N_10062,N_9940,N_9945);
nand U10063 (N_10063,N_9943,N_9881);
nor U10064 (N_10064,N_9882,N_9881);
nand U10065 (N_10065,N_9989,N_9966);
or U10066 (N_10066,N_9934,N_9992);
xor U10067 (N_10067,N_9977,N_9987);
and U10068 (N_10068,N_9919,N_9886);
and U10069 (N_10069,N_9925,N_9899);
nor U10070 (N_10070,N_9982,N_9993);
or U10071 (N_10071,N_9968,N_9948);
or U10072 (N_10072,N_9891,N_9996);
or U10073 (N_10073,N_9925,N_9891);
nand U10074 (N_10074,N_9892,N_9974);
nand U10075 (N_10075,N_9886,N_9982);
nand U10076 (N_10076,N_9907,N_9987);
nand U10077 (N_10077,N_9988,N_9929);
xnor U10078 (N_10078,N_9936,N_9917);
xor U10079 (N_10079,N_9943,N_9921);
nor U10080 (N_10080,N_9945,N_9909);
or U10081 (N_10081,N_9901,N_9962);
nor U10082 (N_10082,N_9933,N_9948);
or U10083 (N_10083,N_9972,N_9946);
or U10084 (N_10084,N_9892,N_9999);
xor U10085 (N_10085,N_9901,N_9889);
xnor U10086 (N_10086,N_9892,N_9959);
or U10087 (N_10087,N_9928,N_9902);
or U10088 (N_10088,N_9902,N_9951);
xor U10089 (N_10089,N_9894,N_9882);
nor U10090 (N_10090,N_9896,N_9885);
nand U10091 (N_10091,N_9914,N_9973);
xnor U10092 (N_10092,N_9930,N_9891);
nand U10093 (N_10093,N_9944,N_9886);
and U10094 (N_10094,N_9888,N_9967);
and U10095 (N_10095,N_9883,N_9992);
xor U10096 (N_10096,N_9971,N_9943);
and U10097 (N_10097,N_9937,N_9959);
nor U10098 (N_10098,N_9875,N_9976);
xor U10099 (N_10099,N_9905,N_9948);
or U10100 (N_10100,N_9907,N_9957);
nor U10101 (N_10101,N_9994,N_9918);
xor U10102 (N_10102,N_9948,N_9979);
or U10103 (N_10103,N_9915,N_9889);
nor U10104 (N_10104,N_9931,N_9969);
nand U10105 (N_10105,N_9960,N_9924);
nand U10106 (N_10106,N_9924,N_9981);
or U10107 (N_10107,N_9880,N_9980);
xnor U10108 (N_10108,N_9886,N_9900);
nor U10109 (N_10109,N_9956,N_9974);
and U10110 (N_10110,N_9921,N_9958);
nor U10111 (N_10111,N_9911,N_9963);
or U10112 (N_10112,N_9877,N_9935);
and U10113 (N_10113,N_9927,N_9934);
xnor U10114 (N_10114,N_9998,N_9937);
xor U10115 (N_10115,N_9949,N_9884);
or U10116 (N_10116,N_9974,N_9889);
or U10117 (N_10117,N_9939,N_9915);
or U10118 (N_10118,N_9921,N_9933);
or U10119 (N_10119,N_9923,N_9888);
or U10120 (N_10120,N_9965,N_9976);
xor U10121 (N_10121,N_9972,N_9956);
nand U10122 (N_10122,N_9996,N_9959);
nor U10123 (N_10123,N_9926,N_9996);
xnor U10124 (N_10124,N_9900,N_9936);
xor U10125 (N_10125,N_10118,N_10112);
and U10126 (N_10126,N_10016,N_10020);
nor U10127 (N_10127,N_10085,N_10092);
xnor U10128 (N_10128,N_10017,N_10060);
and U10129 (N_10129,N_10030,N_10091);
nor U10130 (N_10130,N_10102,N_10120);
xnor U10131 (N_10131,N_10025,N_10045);
and U10132 (N_10132,N_10070,N_10121);
nand U10133 (N_10133,N_10098,N_10021);
xor U10134 (N_10134,N_10003,N_10095);
nand U10135 (N_10135,N_10004,N_10038);
nand U10136 (N_10136,N_10100,N_10008);
nor U10137 (N_10137,N_10073,N_10062);
nor U10138 (N_10138,N_10012,N_10006);
nor U10139 (N_10139,N_10103,N_10117);
nor U10140 (N_10140,N_10108,N_10011);
nand U10141 (N_10141,N_10055,N_10067);
and U10142 (N_10142,N_10072,N_10093);
xor U10143 (N_10143,N_10054,N_10002);
nand U10144 (N_10144,N_10039,N_10032);
nor U10145 (N_10145,N_10069,N_10050);
or U10146 (N_10146,N_10047,N_10111);
or U10147 (N_10147,N_10087,N_10027);
or U10148 (N_10148,N_10029,N_10049);
or U10149 (N_10149,N_10089,N_10031);
xor U10150 (N_10150,N_10022,N_10059);
xor U10151 (N_10151,N_10097,N_10010);
xnor U10152 (N_10152,N_10099,N_10001);
or U10153 (N_10153,N_10075,N_10051);
and U10154 (N_10154,N_10115,N_10086);
and U10155 (N_10155,N_10122,N_10056);
xnor U10156 (N_10156,N_10015,N_10013);
nand U10157 (N_10157,N_10066,N_10014);
or U10158 (N_10158,N_10081,N_10005);
and U10159 (N_10159,N_10104,N_10018);
nor U10160 (N_10160,N_10034,N_10040);
nand U10161 (N_10161,N_10044,N_10043);
and U10162 (N_10162,N_10065,N_10058);
or U10163 (N_10163,N_10084,N_10079);
nand U10164 (N_10164,N_10033,N_10037);
nor U10165 (N_10165,N_10000,N_10035);
nand U10166 (N_10166,N_10036,N_10094);
and U10167 (N_10167,N_10074,N_10106);
and U10168 (N_10168,N_10064,N_10007);
nand U10169 (N_10169,N_10046,N_10096);
or U10170 (N_10170,N_10090,N_10088);
or U10171 (N_10171,N_10042,N_10071);
or U10172 (N_10172,N_10048,N_10052);
and U10173 (N_10173,N_10124,N_10101);
or U10174 (N_10174,N_10019,N_10063);
and U10175 (N_10175,N_10028,N_10083);
or U10176 (N_10176,N_10109,N_10023);
and U10177 (N_10177,N_10105,N_10068);
or U10178 (N_10178,N_10078,N_10110);
xor U10179 (N_10179,N_10116,N_10009);
and U10180 (N_10180,N_10061,N_10057);
nor U10181 (N_10181,N_10114,N_10026);
or U10182 (N_10182,N_10082,N_10119);
and U10183 (N_10183,N_10113,N_10041);
or U10184 (N_10184,N_10053,N_10107);
and U10185 (N_10185,N_10024,N_10076);
or U10186 (N_10186,N_10077,N_10123);
and U10187 (N_10187,N_10080,N_10121);
and U10188 (N_10188,N_10095,N_10014);
nand U10189 (N_10189,N_10102,N_10013);
or U10190 (N_10190,N_10012,N_10087);
xnor U10191 (N_10191,N_10023,N_10065);
or U10192 (N_10192,N_10019,N_10120);
and U10193 (N_10193,N_10025,N_10094);
nand U10194 (N_10194,N_10051,N_10049);
and U10195 (N_10195,N_10097,N_10085);
or U10196 (N_10196,N_10088,N_10060);
xnor U10197 (N_10197,N_10112,N_10055);
nand U10198 (N_10198,N_10096,N_10013);
xnor U10199 (N_10199,N_10036,N_10024);
or U10200 (N_10200,N_10021,N_10117);
and U10201 (N_10201,N_10034,N_10003);
nand U10202 (N_10202,N_10110,N_10117);
nand U10203 (N_10203,N_10020,N_10085);
and U10204 (N_10204,N_10084,N_10037);
xor U10205 (N_10205,N_10103,N_10056);
and U10206 (N_10206,N_10086,N_10110);
xnor U10207 (N_10207,N_10116,N_10123);
or U10208 (N_10208,N_10105,N_10107);
nor U10209 (N_10209,N_10059,N_10047);
nor U10210 (N_10210,N_10007,N_10038);
xor U10211 (N_10211,N_10113,N_10068);
nor U10212 (N_10212,N_10052,N_10047);
and U10213 (N_10213,N_10067,N_10030);
nor U10214 (N_10214,N_10073,N_10118);
or U10215 (N_10215,N_10091,N_10113);
nand U10216 (N_10216,N_10091,N_10121);
or U10217 (N_10217,N_10069,N_10044);
xnor U10218 (N_10218,N_10026,N_10053);
nand U10219 (N_10219,N_10060,N_10035);
and U10220 (N_10220,N_10107,N_10044);
nor U10221 (N_10221,N_10072,N_10075);
xor U10222 (N_10222,N_10064,N_10099);
or U10223 (N_10223,N_10115,N_10063);
nor U10224 (N_10224,N_10005,N_10007);
and U10225 (N_10225,N_10074,N_10085);
nand U10226 (N_10226,N_10011,N_10041);
or U10227 (N_10227,N_10113,N_10031);
nor U10228 (N_10228,N_10005,N_10111);
or U10229 (N_10229,N_10008,N_10027);
nor U10230 (N_10230,N_10003,N_10065);
nand U10231 (N_10231,N_10038,N_10049);
and U10232 (N_10232,N_10112,N_10063);
or U10233 (N_10233,N_10064,N_10022);
or U10234 (N_10234,N_10056,N_10117);
or U10235 (N_10235,N_10027,N_10082);
and U10236 (N_10236,N_10035,N_10072);
nor U10237 (N_10237,N_10053,N_10040);
xor U10238 (N_10238,N_10094,N_10106);
nand U10239 (N_10239,N_10099,N_10100);
nor U10240 (N_10240,N_10070,N_10051);
nand U10241 (N_10241,N_10123,N_10108);
nor U10242 (N_10242,N_10040,N_10070);
or U10243 (N_10243,N_10008,N_10019);
nand U10244 (N_10244,N_10015,N_10005);
or U10245 (N_10245,N_10013,N_10006);
and U10246 (N_10246,N_10118,N_10123);
or U10247 (N_10247,N_10020,N_10074);
and U10248 (N_10248,N_10079,N_10087);
nor U10249 (N_10249,N_10045,N_10049);
and U10250 (N_10250,N_10143,N_10198);
or U10251 (N_10251,N_10235,N_10209);
or U10252 (N_10252,N_10233,N_10244);
xor U10253 (N_10253,N_10164,N_10222);
or U10254 (N_10254,N_10212,N_10140);
nor U10255 (N_10255,N_10232,N_10202);
nor U10256 (N_10256,N_10204,N_10148);
nor U10257 (N_10257,N_10162,N_10219);
nand U10258 (N_10258,N_10165,N_10210);
or U10259 (N_10259,N_10179,N_10213);
nand U10260 (N_10260,N_10173,N_10223);
xnor U10261 (N_10261,N_10144,N_10182);
and U10262 (N_10262,N_10137,N_10246);
nor U10263 (N_10263,N_10205,N_10201);
xnor U10264 (N_10264,N_10159,N_10203);
nand U10265 (N_10265,N_10239,N_10149);
or U10266 (N_10266,N_10224,N_10183);
nor U10267 (N_10267,N_10237,N_10227);
or U10268 (N_10268,N_10138,N_10166);
and U10269 (N_10269,N_10199,N_10238);
or U10270 (N_10270,N_10163,N_10161);
and U10271 (N_10271,N_10152,N_10142);
nor U10272 (N_10272,N_10128,N_10200);
or U10273 (N_10273,N_10215,N_10195);
nor U10274 (N_10274,N_10171,N_10245);
or U10275 (N_10275,N_10151,N_10176);
and U10276 (N_10276,N_10131,N_10216);
or U10277 (N_10277,N_10247,N_10221);
and U10278 (N_10278,N_10226,N_10242);
and U10279 (N_10279,N_10193,N_10206);
xor U10280 (N_10280,N_10236,N_10129);
or U10281 (N_10281,N_10189,N_10197);
nor U10282 (N_10282,N_10181,N_10207);
xor U10283 (N_10283,N_10187,N_10160);
nand U10284 (N_10284,N_10214,N_10172);
or U10285 (N_10285,N_10241,N_10130);
nor U10286 (N_10286,N_10150,N_10178);
or U10287 (N_10287,N_10184,N_10146);
or U10288 (N_10288,N_10240,N_10220);
nor U10289 (N_10289,N_10135,N_10145);
xor U10290 (N_10290,N_10157,N_10211);
nand U10291 (N_10291,N_10133,N_10234);
or U10292 (N_10292,N_10186,N_10218);
nor U10293 (N_10293,N_10208,N_10249);
xnor U10294 (N_10294,N_10196,N_10231);
or U10295 (N_10295,N_10230,N_10217);
xor U10296 (N_10296,N_10174,N_10229);
nand U10297 (N_10297,N_10136,N_10156);
or U10298 (N_10298,N_10169,N_10177);
xor U10299 (N_10299,N_10168,N_10185);
or U10300 (N_10300,N_10155,N_10134);
or U10301 (N_10301,N_10175,N_10167);
nor U10302 (N_10302,N_10228,N_10125);
nand U10303 (N_10303,N_10243,N_10248);
nand U10304 (N_10304,N_10154,N_10188);
xor U10305 (N_10305,N_10139,N_10132);
nor U10306 (N_10306,N_10141,N_10126);
xor U10307 (N_10307,N_10190,N_10191);
nand U10308 (N_10308,N_10180,N_10225);
or U10309 (N_10309,N_10153,N_10194);
and U10310 (N_10310,N_10158,N_10147);
nand U10311 (N_10311,N_10170,N_10127);
nor U10312 (N_10312,N_10192,N_10225);
xnor U10313 (N_10313,N_10238,N_10156);
and U10314 (N_10314,N_10221,N_10200);
and U10315 (N_10315,N_10173,N_10175);
and U10316 (N_10316,N_10199,N_10146);
nand U10317 (N_10317,N_10245,N_10187);
xor U10318 (N_10318,N_10155,N_10163);
and U10319 (N_10319,N_10136,N_10206);
nand U10320 (N_10320,N_10127,N_10241);
or U10321 (N_10321,N_10138,N_10133);
xnor U10322 (N_10322,N_10150,N_10244);
nand U10323 (N_10323,N_10169,N_10238);
nand U10324 (N_10324,N_10219,N_10246);
and U10325 (N_10325,N_10226,N_10174);
or U10326 (N_10326,N_10194,N_10232);
or U10327 (N_10327,N_10192,N_10143);
nor U10328 (N_10328,N_10132,N_10150);
nand U10329 (N_10329,N_10168,N_10219);
nand U10330 (N_10330,N_10200,N_10237);
or U10331 (N_10331,N_10148,N_10195);
nor U10332 (N_10332,N_10181,N_10246);
or U10333 (N_10333,N_10237,N_10218);
nand U10334 (N_10334,N_10227,N_10133);
nand U10335 (N_10335,N_10212,N_10158);
xor U10336 (N_10336,N_10195,N_10197);
xor U10337 (N_10337,N_10149,N_10171);
xor U10338 (N_10338,N_10142,N_10206);
or U10339 (N_10339,N_10170,N_10166);
nor U10340 (N_10340,N_10231,N_10201);
xor U10341 (N_10341,N_10243,N_10151);
nand U10342 (N_10342,N_10248,N_10187);
or U10343 (N_10343,N_10178,N_10235);
or U10344 (N_10344,N_10188,N_10193);
and U10345 (N_10345,N_10141,N_10180);
and U10346 (N_10346,N_10130,N_10208);
nand U10347 (N_10347,N_10174,N_10240);
or U10348 (N_10348,N_10150,N_10175);
nand U10349 (N_10349,N_10135,N_10231);
xnor U10350 (N_10350,N_10156,N_10186);
nand U10351 (N_10351,N_10244,N_10213);
or U10352 (N_10352,N_10138,N_10141);
xor U10353 (N_10353,N_10231,N_10182);
and U10354 (N_10354,N_10186,N_10205);
nand U10355 (N_10355,N_10172,N_10158);
and U10356 (N_10356,N_10153,N_10169);
nor U10357 (N_10357,N_10239,N_10146);
nor U10358 (N_10358,N_10132,N_10192);
and U10359 (N_10359,N_10135,N_10186);
nor U10360 (N_10360,N_10131,N_10224);
xor U10361 (N_10361,N_10212,N_10242);
nor U10362 (N_10362,N_10216,N_10210);
nand U10363 (N_10363,N_10244,N_10209);
or U10364 (N_10364,N_10193,N_10226);
nand U10365 (N_10365,N_10216,N_10148);
nand U10366 (N_10366,N_10180,N_10145);
nor U10367 (N_10367,N_10141,N_10208);
and U10368 (N_10368,N_10131,N_10234);
and U10369 (N_10369,N_10208,N_10226);
or U10370 (N_10370,N_10203,N_10192);
xnor U10371 (N_10371,N_10224,N_10134);
and U10372 (N_10372,N_10140,N_10216);
or U10373 (N_10373,N_10184,N_10175);
xor U10374 (N_10374,N_10222,N_10204);
or U10375 (N_10375,N_10346,N_10254);
xor U10376 (N_10376,N_10307,N_10342);
nor U10377 (N_10377,N_10351,N_10275);
and U10378 (N_10378,N_10278,N_10335);
and U10379 (N_10379,N_10304,N_10288);
xnor U10380 (N_10380,N_10343,N_10289);
nor U10381 (N_10381,N_10360,N_10314);
nand U10382 (N_10382,N_10340,N_10305);
and U10383 (N_10383,N_10272,N_10258);
nand U10384 (N_10384,N_10253,N_10260);
or U10385 (N_10385,N_10374,N_10287);
or U10386 (N_10386,N_10296,N_10312);
nand U10387 (N_10387,N_10257,N_10334);
or U10388 (N_10388,N_10306,N_10338);
xnor U10389 (N_10389,N_10282,N_10333);
and U10390 (N_10390,N_10316,N_10372);
nor U10391 (N_10391,N_10370,N_10251);
nand U10392 (N_10392,N_10279,N_10269);
xnor U10393 (N_10393,N_10273,N_10271);
or U10394 (N_10394,N_10284,N_10315);
xnor U10395 (N_10395,N_10280,N_10297);
and U10396 (N_10396,N_10294,N_10256);
xor U10397 (N_10397,N_10362,N_10349);
and U10398 (N_10398,N_10301,N_10341);
xnor U10399 (N_10399,N_10292,N_10366);
xor U10400 (N_10400,N_10255,N_10285);
or U10401 (N_10401,N_10295,N_10331);
or U10402 (N_10402,N_10328,N_10265);
nor U10403 (N_10403,N_10252,N_10359);
nand U10404 (N_10404,N_10365,N_10322);
and U10405 (N_10405,N_10319,N_10268);
nand U10406 (N_10406,N_10259,N_10367);
or U10407 (N_10407,N_10302,N_10353);
xnor U10408 (N_10408,N_10320,N_10310);
or U10409 (N_10409,N_10318,N_10337);
nand U10410 (N_10410,N_10313,N_10363);
nor U10411 (N_10411,N_10311,N_10369);
and U10412 (N_10412,N_10281,N_10274);
nor U10413 (N_10413,N_10355,N_10299);
and U10414 (N_10414,N_10347,N_10330);
xnor U10415 (N_10415,N_10354,N_10345);
xnor U10416 (N_10416,N_10358,N_10300);
and U10417 (N_10417,N_10336,N_10332);
nand U10418 (N_10418,N_10368,N_10323);
xor U10419 (N_10419,N_10270,N_10276);
and U10420 (N_10420,N_10293,N_10324);
nand U10421 (N_10421,N_10250,N_10263);
and U10422 (N_10422,N_10290,N_10371);
or U10423 (N_10423,N_10329,N_10344);
nand U10424 (N_10424,N_10267,N_10356);
or U10425 (N_10425,N_10262,N_10350);
nor U10426 (N_10426,N_10361,N_10303);
nand U10427 (N_10427,N_10373,N_10277);
or U10428 (N_10428,N_10321,N_10317);
or U10429 (N_10429,N_10286,N_10266);
nand U10430 (N_10430,N_10357,N_10339);
nor U10431 (N_10431,N_10261,N_10298);
nor U10432 (N_10432,N_10308,N_10291);
xnor U10433 (N_10433,N_10327,N_10364);
nor U10434 (N_10434,N_10352,N_10264);
xnor U10435 (N_10435,N_10348,N_10326);
nor U10436 (N_10436,N_10325,N_10309);
xor U10437 (N_10437,N_10283,N_10308);
nor U10438 (N_10438,N_10293,N_10303);
nand U10439 (N_10439,N_10282,N_10326);
or U10440 (N_10440,N_10294,N_10353);
or U10441 (N_10441,N_10291,N_10343);
and U10442 (N_10442,N_10297,N_10271);
and U10443 (N_10443,N_10365,N_10260);
nor U10444 (N_10444,N_10353,N_10292);
nor U10445 (N_10445,N_10365,N_10253);
xor U10446 (N_10446,N_10360,N_10369);
and U10447 (N_10447,N_10360,N_10302);
xor U10448 (N_10448,N_10274,N_10258);
and U10449 (N_10449,N_10358,N_10371);
nor U10450 (N_10450,N_10288,N_10262);
and U10451 (N_10451,N_10344,N_10326);
xor U10452 (N_10452,N_10348,N_10371);
or U10453 (N_10453,N_10301,N_10297);
or U10454 (N_10454,N_10336,N_10371);
xnor U10455 (N_10455,N_10328,N_10331);
or U10456 (N_10456,N_10312,N_10275);
xnor U10457 (N_10457,N_10277,N_10303);
nor U10458 (N_10458,N_10332,N_10351);
or U10459 (N_10459,N_10308,N_10323);
and U10460 (N_10460,N_10265,N_10348);
nand U10461 (N_10461,N_10334,N_10252);
and U10462 (N_10462,N_10270,N_10306);
xor U10463 (N_10463,N_10295,N_10253);
or U10464 (N_10464,N_10291,N_10351);
nor U10465 (N_10465,N_10256,N_10327);
or U10466 (N_10466,N_10299,N_10348);
and U10467 (N_10467,N_10331,N_10278);
nor U10468 (N_10468,N_10280,N_10253);
nor U10469 (N_10469,N_10343,N_10255);
nor U10470 (N_10470,N_10357,N_10313);
xnor U10471 (N_10471,N_10311,N_10348);
xnor U10472 (N_10472,N_10330,N_10255);
nor U10473 (N_10473,N_10285,N_10329);
xnor U10474 (N_10474,N_10316,N_10257);
or U10475 (N_10475,N_10295,N_10275);
xnor U10476 (N_10476,N_10310,N_10330);
nor U10477 (N_10477,N_10318,N_10320);
or U10478 (N_10478,N_10278,N_10313);
and U10479 (N_10479,N_10347,N_10346);
nand U10480 (N_10480,N_10374,N_10304);
and U10481 (N_10481,N_10352,N_10297);
nor U10482 (N_10482,N_10254,N_10268);
nand U10483 (N_10483,N_10335,N_10316);
or U10484 (N_10484,N_10366,N_10256);
or U10485 (N_10485,N_10278,N_10265);
or U10486 (N_10486,N_10370,N_10297);
nor U10487 (N_10487,N_10321,N_10273);
nand U10488 (N_10488,N_10327,N_10284);
and U10489 (N_10489,N_10298,N_10320);
or U10490 (N_10490,N_10358,N_10273);
nor U10491 (N_10491,N_10260,N_10259);
nor U10492 (N_10492,N_10272,N_10262);
and U10493 (N_10493,N_10368,N_10290);
xnor U10494 (N_10494,N_10281,N_10270);
nand U10495 (N_10495,N_10324,N_10302);
xnor U10496 (N_10496,N_10328,N_10315);
nand U10497 (N_10497,N_10355,N_10301);
nand U10498 (N_10498,N_10321,N_10364);
nor U10499 (N_10499,N_10335,N_10364);
nand U10500 (N_10500,N_10455,N_10463);
and U10501 (N_10501,N_10488,N_10412);
nor U10502 (N_10502,N_10425,N_10396);
and U10503 (N_10503,N_10462,N_10380);
or U10504 (N_10504,N_10395,N_10486);
and U10505 (N_10505,N_10499,N_10427);
xor U10506 (N_10506,N_10430,N_10401);
nor U10507 (N_10507,N_10482,N_10375);
and U10508 (N_10508,N_10406,N_10415);
nor U10509 (N_10509,N_10470,N_10474);
nand U10510 (N_10510,N_10402,N_10400);
xor U10511 (N_10511,N_10460,N_10403);
nand U10512 (N_10512,N_10493,N_10420);
xnor U10513 (N_10513,N_10445,N_10382);
nor U10514 (N_10514,N_10436,N_10461);
and U10515 (N_10515,N_10393,N_10422);
nor U10516 (N_10516,N_10389,N_10405);
and U10517 (N_10517,N_10409,N_10478);
and U10518 (N_10518,N_10448,N_10388);
xnor U10519 (N_10519,N_10469,N_10394);
xor U10520 (N_10520,N_10465,N_10464);
and U10521 (N_10521,N_10379,N_10381);
and U10522 (N_10522,N_10386,N_10492);
or U10523 (N_10523,N_10452,N_10471);
nand U10524 (N_10524,N_10407,N_10477);
nor U10525 (N_10525,N_10467,N_10441);
and U10526 (N_10526,N_10489,N_10392);
or U10527 (N_10527,N_10473,N_10418);
xnor U10528 (N_10528,N_10449,N_10385);
nor U10529 (N_10529,N_10456,N_10475);
nand U10530 (N_10530,N_10431,N_10426);
xnor U10531 (N_10531,N_10495,N_10447);
and U10532 (N_10532,N_10484,N_10480);
or U10533 (N_10533,N_10483,N_10444);
nor U10534 (N_10534,N_10399,N_10421);
xnor U10535 (N_10535,N_10397,N_10432);
xor U10536 (N_10536,N_10408,N_10424);
xor U10537 (N_10537,N_10417,N_10458);
xnor U10538 (N_10538,N_10494,N_10442);
nor U10539 (N_10539,N_10378,N_10479);
xnor U10540 (N_10540,N_10419,N_10451);
or U10541 (N_10541,N_10497,N_10453);
nor U10542 (N_10542,N_10391,N_10446);
nor U10543 (N_10543,N_10496,N_10414);
xnor U10544 (N_10544,N_10466,N_10468);
nor U10545 (N_10545,N_10454,N_10410);
nand U10546 (N_10546,N_10498,N_10491);
or U10547 (N_10547,N_10459,N_10383);
xor U10548 (N_10548,N_10435,N_10428);
and U10549 (N_10549,N_10376,N_10443);
or U10550 (N_10550,N_10411,N_10384);
and U10551 (N_10551,N_10434,N_10485);
nor U10552 (N_10552,N_10390,N_10413);
nor U10553 (N_10553,N_10450,N_10487);
and U10554 (N_10554,N_10377,N_10481);
and U10555 (N_10555,N_10416,N_10457);
or U10556 (N_10556,N_10472,N_10398);
or U10557 (N_10557,N_10476,N_10490);
and U10558 (N_10558,N_10423,N_10429);
or U10559 (N_10559,N_10437,N_10438);
xor U10560 (N_10560,N_10439,N_10404);
and U10561 (N_10561,N_10433,N_10440);
or U10562 (N_10562,N_10387,N_10403);
or U10563 (N_10563,N_10406,N_10466);
and U10564 (N_10564,N_10443,N_10403);
or U10565 (N_10565,N_10388,N_10393);
nor U10566 (N_10566,N_10433,N_10467);
or U10567 (N_10567,N_10492,N_10479);
nand U10568 (N_10568,N_10392,N_10429);
nor U10569 (N_10569,N_10411,N_10399);
or U10570 (N_10570,N_10434,N_10453);
or U10571 (N_10571,N_10484,N_10471);
xnor U10572 (N_10572,N_10397,N_10386);
nand U10573 (N_10573,N_10488,N_10400);
nand U10574 (N_10574,N_10478,N_10475);
nor U10575 (N_10575,N_10490,N_10478);
nor U10576 (N_10576,N_10419,N_10380);
nand U10577 (N_10577,N_10491,N_10427);
nand U10578 (N_10578,N_10433,N_10486);
xor U10579 (N_10579,N_10476,N_10473);
nand U10580 (N_10580,N_10490,N_10391);
or U10581 (N_10581,N_10491,N_10459);
nand U10582 (N_10582,N_10414,N_10457);
and U10583 (N_10583,N_10474,N_10437);
nor U10584 (N_10584,N_10438,N_10458);
nor U10585 (N_10585,N_10461,N_10427);
or U10586 (N_10586,N_10477,N_10389);
nand U10587 (N_10587,N_10417,N_10428);
xor U10588 (N_10588,N_10440,N_10455);
nand U10589 (N_10589,N_10391,N_10420);
xor U10590 (N_10590,N_10419,N_10389);
xnor U10591 (N_10591,N_10427,N_10402);
nand U10592 (N_10592,N_10379,N_10467);
nand U10593 (N_10593,N_10384,N_10487);
or U10594 (N_10594,N_10419,N_10387);
or U10595 (N_10595,N_10487,N_10441);
nand U10596 (N_10596,N_10383,N_10394);
xor U10597 (N_10597,N_10376,N_10467);
and U10598 (N_10598,N_10461,N_10394);
nor U10599 (N_10599,N_10459,N_10464);
nor U10600 (N_10600,N_10487,N_10375);
and U10601 (N_10601,N_10454,N_10464);
xnor U10602 (N_10602,N_10381,N_10455);
xnor U10603 (N_10603,N_10403,N_10379);
xnor U10604 (N_10604,N_10444,N_10473);
nor U10605 (N_10605,N_10408,N_10439);
and U10606 (N_10606,N_10439,N_10390);
and U10607 (N_10607,N_10396,N_10477);
nand U10608 (N_10608,N_10398,N_10494);
nor U10609 (N_10609,N_10384,N_10425);
or U10610 (N_10610,N_10448,N_10487);
nand U10611 (N_10611,N_10461,N_10466);
nor U10612 (N_10612,N_10474,N_10379);
and U10613 (N_10613,N_10379,N_10377);
and U10614 (N_10614,N_10487,N_10404);
nand U10615 (N_10615,N_10492,N_10494);
and U10616 (N_10616,N_10400,N_10468);
nor U10617 (N_10617,N_10398,N_10448);
xor U10618 (N_10618,N_10388,N_10394);
or U10619 (N_10619,N_10495,N_10456);
and U10620 (N_10620,N_10395,N_10425);
nand U10621 (N_10621,N_10442,N_10395);
nand U10622 (N_10622,N_10444,N_10463);
or U10623 (N_10623,N_10378,N_10478);
nand U10624 (N_10624,N_10409,N_10448);
xor U10625 (N_10625,N_10544,N_10529);
xor U10626 (N_10626,N_10598,N_10595);
nand U10627 (N_10627,N_10531,N_10602);
nand U10628 (N_10628,N_10538,N_10579);
and U10629 (N_10629,N_10516,N_10607);
nor U10630 (N_10630,N_10609,N_10572);
and U10631 (N_10631,N_10546,N_10526);
xnor U10632 (N_10632,N_10560,N_10564);
xor U10633 (N_10633,N_10553,N_10588);
nor U10634 (N_10634,N_10583,N_10527);
xnor U10635 (N_10635,N_10556,N_10610);
xnor U10636 (N_10636,N_10541,N_10518);
nor U10637 (N_10637,N_10569,N_10574);
and U10638 (N_10638,N_10501,N_10559);
nand U10639 (N_10639,N_10508,N_10591);
nand U10640 (N_10640,N_10615,N_10562);
and U10641 (N_10641,N_10509,N_10599);
nand U10642 (N_10642,N_10623,N_10597);
and U10643 (N_10643,N_10594,N_10523);
nor U10644 (N_10644,N_10580,N_10507);
nor U10645 (N_10645,N_10521,N_10582);
and U10646 (N_10646,N_10536,N_10601);
nor U10647 (N_10647,N_10571,N_10568);
nor U10648 (N_10648,N_10503,N_10522);
or U10649 (N_10649,N_10510,N_10505);
xor U10650 (N_10650,N_10528,N_10547);
nand U10651 (N_10651,N_10567,N_10617);
nor U10652 (N_10652,N_10624,N_10613);
or U10653 (N_10653,N_10621,N_10515);
nand U10654 (N_10654,N_10577,N_10540);
nor U10655 (N_10655,N_10614,N_10519);
nor U10656 (N_10656,N_10604,N_10539);
or U10657 (N_10657,N_10513,N_10592);
or U10658 (N_10658,N_10514,N_10611);
nor U10659 (N_10659,N_10589,N_10548);
nor U10660 (N_10660,N_10566,N_10576);
nor U10661 (N_10661,N_10587,N_10500);
xor U10662 (N_10662,N_10524,N_10596);
nand U10663 (N_10663,N_10552,N_10561);
xor U10664 (N_10664,N_10586,N_10558);
nor U10665 (N_10665,N_10542,N_10533);
or U10666 (N_10666,N_10545,N_10537);
xor U10667 (N_10667,N_10606,N_10603);
nand U10668 (N_10668,N_10534,N_10578);
nand U10669 (N_10669,N_10570,N_10525);
xnor U10670 (N_10670,N_10549,N_10573);
and U10671 (N_10671,N_10504,N_10590);
and U10672 (N_10672,N_10532,N_10563);
nor U10673 (N_10673,N_10506,N_10618);
nor U10674 (N_10674,N_10554,N_10608);
xor U10675 (N_10675,N_10619,N_10502);
nand U10676 (N_10676,N_10565,N_10535);
nand U10677 (N_10677,N_10512,N_10584);
nand U10678 (N_10678,N_10585,N_10620);
nand U10679 (N_10679,N_10550,N_10555);
nand U10680 (N_10680,N_10517,N_10605);
nand U10681 (N_10681,N_10612,N_10622);
xor U10682 (N_10682,N_10616,N_10511);
xor U10683 (N_10683,N_10557,N_10593);
and U10684 (N_10684,N_10520,N_10581);
nor U10685 (N_10685,N_10575,N_10530);
nor U10686 (N_10686,N_10543,N_10551);
nor U10687 (N_10687,N_10600,N_10554);
nand U10688 (N_10688,N_10544,N_10586);
nand U10689 (N_10689,N_10587,N_10613);
xor U10690 (N_10690,N_10537,N_10514);
nor U10691 (N_10691,N_10581,N_10558);
nand U10692 (N_10692,N_10533,N_10585);
xor U10693 (N_10693,N_10586,N_10582);
or U10694 (N_10694,N_10571,N_10595);
xor U10695 (N_10695,N_10542,N_10524);
nand U10696 (N_10696,N_10530,N_10516);
xnor U10697 (N_10697,N_10563,N_10620);
xor U10698 (N_10698,N_10546,N_10505);
nand U10699 (N_10699,N_10619,N_10573);
nor U10700 (N_10700,N_10578,N_10613);
xor U10701 (N_10701,N_10508,N_10505);
nand U10702 (N_10702,N_10571,N_10522);
or U10703 (N_10703,N_10538,N_10513);
nor U10704 (N_10704,N_10578,N_10581);
nor U10705 (N_10705,N_10621,N_10584);
xor U10706 (N_10706,N_10532,N_10610);
nand U10707 (N_10707,N_10598,N_10501);
nor U10708 (N_10708,N_10553,N_10565);
nor U10709 (N_10709,N_10576,N_10545);
and U10710 (N_10710,N_10525,N_10544);
xor U10711 (N_10711,N_10562,N_10585);
xnor U10712 (N_10712,N_10595,N_10509);
and U10713 (N_10713,N_10500,N_10555);
xnor U10714 (N_10714,N_10566,N_10580);
and U10715 (N_10715,N_10540,N_10590);
xor U10716 (N_10716,N_10602,N_10603);
nor U10717 (N_10717,N_10611,N_10580);
nor U10718 (N_10718,N_10593,N_10521);
nand U10719 (N_10719,N_10601,N_10615);
and U10720 (N_10720,N_10587,N_10570);
or U10721 (N_10721,N_10544,N_10502);
xor U10722 (N_10722,N_10609,N_10521);
and U10723 (N_10723,N_10561,N_10538);
nand U10724 (N_10724,N_10581,N_10535);
and U10725 (N_10725,N_10537,N_10512);
or U10726 (N_10726,N_10591,N_10545);
and U10727 (N_10727,N_10508,N_10506);
xnor U10728 (N_10728,N_10623,N_10533);
nand U10729 (N_10729,N_10528,N_10552);
nor U10730 (N_10730,N_10503,N_10555);
and U10731 (N_10731,N_10604,N_10573);
nor U10732 (N_10732,N_10536,N_10545);
or U10733 (N_10733,N_10544,N_10604);
nand U10734 (N_10734,N_10608,N_10539);
xor U10735 (N_10735,N_10502,N_10533);
nand U10736 (N_10736,N_10541,N_10623);
nand U10737 (N_10737,N_10513,N_10614);
or U10738 (N_10738,N_10587,N_10509);
xor U10739 (N_10739,N_10605,N_10500);
or U10740 (N_10740,N_10569,N_10585);
xor U10741 (N_10741,N_10501,N_10588);
and U10742 (N_10742,N_10584,N_10620);
xnor U10743 (N_10743,N_10603,N_10514);
nor U10744 (N_10744,N_10607,N_10600);
nand U10745 (N_10745,N_10604,N_10505);
nand U10746 (N_10746,N_10563,N_10526);
and U10747 (N_10747,N_10624,N_10618);
nor U10748 (N_10748,N_10587,N_10616);
and U10749 (N_10749,N_10574,N_10599);
or U10750 (N_10750,N_10694,N_10749);
and U10751 (N_10751,N_10738,N_10633);
xnor U10752 (N_10752,N_10682,N_10725);
or U10753 (N_10753,N_10637,N_10693);
or U10754 (N_10754,N_10665,N_10634);
xnor U10755 (N_10755,N_10628,N_10635);
or U10756 (N_10756,N_10746,N_10676);
and U10757 (N_10757,N_10726,N_10681);
or U10758 (N_10758,N_10741,N_10722);
and U10759 (N_10759,N_10699,N_10734);
nand U10760 (N_10760,N_10721,N_10728);
and U10761 (N_10761,N_10745,N_10706);
xnor U10762 (N_10762,N_10642,N_10724);
or U10763 (N_10763,N_10735,N_10648);
nand U10764 (N_10764,N_10672,N_10723);
and U10765 (N_10765,N_10685,N_10684);
nor U10766 (N_10766,N_10652,N_10668);
or U10767 (N_10767,N_10700,N_10687);
nor U10768 (N_10768,N_10670,N_10660);
xnor U10769 (N_10769,N_10698,N_10727);
and U10770 (N_10770,N_10679,N_10743);
nor U10771 (N_10771,N_10653,N_10714);
or U10772 (N_10772,N_10673,N_10658);
and U10773 (N_10773,N_10748,N_10710);
nor U10774 (N_10774,N_10742,N_10733);
xor U10775 (N_10775,N_10664,N_10675);
xor U10776 (N_10776,N_10736,N_10656);
nand U10777 (N_10777,N_10697,N_10715);
or U10778 (N_10778,N_10692,N_10686);
nor U10779 (N_10779,N_10737,N_10646);
xor U10780 (N_10780,N_10667,N_10678);
and U10781 (N_10781,N_10718,N_10732);
nor U10782 (N_10782,N_10747,N_10647);
xnor U10783 (N_10783,N_10671,N_10650);
xnor U10784 (N_10784,N_10707,N_10729);
or U10785 (N_10785,N_10739,N_10627);
xnor U10786 (N_10786,N_10708,N_10689);
and U10787 (N_10787,N_10702,N_10643);
xor U10788 (N_10788,N_10669,N_10740);
or U10789 (N_10789,N_10636,N_10731);
and U10790 (N_10790,N_10630,N_10639);
xor U10791 (N_10791,N_10677,N_10680);
xnor U10792 (N_10792,N_10701,N_10720);
or U10793 (N_10793,N_10631,N_10649);
and U10794 (N_10794,N_10625,N_10629);
and U10795 (N_10795,N_10654,N_10712);
xnor U10796 (N_10796,N_10709,N_10638);
nand U10797 (N_10797,N_10717,N_10662);
or U10798 (N_10798,N_10659,N_10730);
and U10799 (N_10799,N_10645,N_10644);
xnor U10800 (N_10800,N_10655,N_10695);
nor U10801 (N_10801,N_10688,N_10666);
and U10802 (N_10802,N_10626,N_10716);
and U10803 (N_10803,N_10632,N_10674);
xnor U10804 (N_10804,N_10690,N_10691);
or U10805 (N_10805,N_10696,N_10713);
or U10806 (N_10806,N_10661,N_10704);
or U10807 (N_10807,N_10663,N_10703);
xor U10808 (N_10808,N_10651,N_10657);
nor U10809 (N_10809,N_10711,N_10719);
nor U10810 (N_10810,N_10683,N_10744);
or U10811 (N_10811,N_10705,N_10641);
and U10812 (N_10812,N_10640,N_10749);
nand U10813 (N_10813,N_10645,N_10699);
and U10814 (N_10814,N_10748,N_10701);
and U10815 (N_10815,N_10707,N_10692);
nand U10816 (N_10816,N_10643,N_10717);
xor U10817 (N_10817,N_10655,N_10649);
nor U10818 (N_10818,N_10673,N_10702);
xor U10819 (N_10819,N_10720,N_10674);
and U10820 (N_10820,N_10640,N_10698);
and U10821 (N_10821,N_10705,N_10625);
nand U10822 (N_10822,N_10691,N_10735);
and U10823 (N_10823,N_10647,N_10648);
nand U10824 (N_10824,N_10720,N_10630);
nor U10825 (N_10825,N_10676,N_10725);
xnor U10826 (N_10826,N_10674,N_10647);
xor U10827 (N_10827,N_10712,N_10689);
xnor U10828 (N_10828,N_10639,N_10741);
and U10829 (N_10829,N_10665,N_10720);
and U10830 (N_10830,N_10627,N_10695);
nand U10831 (N_10831,N_10651,N_10640);
and U10832 (N_10832,N_10712,N_10630);
xor U10833 (N_10833,N_10748,N_10723);
nor U10834 (N_10834,N_10639,N_10691);
or U10835 (N_10835,N_10713,N_10732);
and U10836 (N_10836,N_10675,N_10655);
or U10837 (N_10837,N_10699,N_10715);
nand U10838 (N_10838,N_10716,N_10728);
or U10839 (N_10839,N_10635,N_10742);
nand U10840 (N_10840,N_10746,N_10710);
and U10841 (N_10841,N_10678,N_10643);
and U10842 (N_10842,N_10661,N_10744);
or U10843 (N_10843,N_10693,N_10739);
nand U10844 (N_10844,N_10685,N_10657);
nor U10845 (N_10845,N_10744,N_10676);
and U10846 (N_10846,N_10653,N_10678);
nand U10847 (N_10847,N_10684,N_10711);
nand U10848 (N_10848,N_10641,N_10697);
nor U10849 (N_10849,N_10671,N_10741);
and U10850 (N_10850,N_10687,N_10740);
or U10851 (N_10851,N_10667,N_10742);
xnor U10852 (N_10852,N_10708,N_10638);
nand U10853 (N_10853,N_10705,N_10643);
nand U10854 (N_10854,N_10727,N_10670);
nor U10855 (N_10855,N_10710,N_10731);
xnor U10856 (N_10856,N_10663,N_10732);
xor U10857 (N_10857,N_10665,N_10723);
xor U10858 (N_10858,N_10704,N_10706);
and U10859 (N_10859,N_10683,N_10730);
nor U10860 (N_10860,N_10670,N_10685);
nand U10861 (N_10861,N_10742,N_10682);
nand U10862 (N_10862,N_10706,N_10738);
nand U10863 (N_10863,N_10728,N_10680);
xnor U10864 (N_10864,N_10674,N_10681);
and U10865 (N_10865,N_10748,N_10735);
xnor U10866 (N_10866,N_10717,N_10696);
nor U10867 (N_10867,N_10731,N_10712);
nor U10868 (N_10868,N_10699,N_10659);
xor U10869 (N_10869,N_10683,N_10636);
or U10870 (N_10870,N_10668,N_10737);
nor U10871 (N_10871,N_10723,N_10693);
nor U10872 (N_10872,N_10651,N_10628);
and U10873 (N_10873,N_10634,N_10719);
or U10874 (N_10874,N_10638,N_10689);
nor U10875 (N_10875,N_10808,N_10781);
nand U10876 (N_10876,N_10853,N_10869);
xnor U10877 (N_10877,N_10795,N_10874);
xnor U10878 (N_10878,N_10842,N_10813);
nand U10879 (N_10879,N_10793,N_10790);
and U10880 (N_10880,N_10837,N_10763);
or U10881 (N_10881,N_10782,N_10772);
xor U10882 (N_10882,N_10819,N_10871);
nor U10883 (N_10883,N_10850,N_10815);
nor U10884 (N_10884,N_10859,N_10811);
and U10885 (N_10885,N_10827,N_10836);
and U10886 (N_10886,N_10833,N_10750);
and U10887 (N_10887,N_10797,N_10840);
and U10888 (N_10888,N_10804,N_10821);
and U10889 (N_10889,N_10768,N_10812);
and U10890 (N_10890,N_10770,N_10826);
and U10891 (N_10891,N_10769,N_10788);
or U10892 (N_10892,N_10818,N_10754);
or U10893 (N_10893,N_10798,N_10847);
xnor U10894 (N_10894,N_10841,N_10868);
or U10895 (N_10895,N_10757,N_10838);
nand U10896 (N_10896,N_10828,N_10823);
xnor U10897 (N_10897,N_10807,N_10830);
and U10898 (N_10898,N_10835,N_10771);
nand U10899 (N_10899,N_10872,N_10831);
nor U10900 (N_10900,N_10861,N_10814);
nor U10901 (N_10901,N_10766,N_10789);
and U10902 (N_10902,N_10761,N_10778);
nand U10903 (N_10903,N_10755,N_10764);
xor U10904 (N_10904,N_10809,N_10864);
nor U10905 (N_10905,N_10780,N_10824);
or U10906 (N_10906,N_10783,N_10794);
nor U10907 (N_10907,N_10796,N_10851);
nand U10908 (N_10908,N_10858,N_10844);
nor U10909 (N_10909,N_10775,N_10839);
or U10910 (N_10910,N_10855,N_10870);
and U10911 (N_10911,N_10786,N_10806);
or U10912 (N_10912,N_10845,N_10856);
nand U10913 (N_10913,N_10832,N_10852);
nor U10914 (N_10914,N_10846,N_10816);
nand U10915 (N_10915,N_10799,N_10863);
xor U10916 (N_10916,N_10817,N_10857);
nand U10917 (N_10917,N_10760,N_10843);
xor U10918 (N_10918,N_10825,N_10829);
nand U10919 (N_10919,N_10751,N_10787);
and U10920 (N_10920,N_10762,N_10805);
nand U10921 (N_10921,N_10784,N_10834);
nand U10922 (N_10922,N_10753,N_10774);
xnor U10923 (N_10923,N_10776,N_10860);
or U10924 (N_10924,N_10822,N_10752);
and U10925 (N_10925,N_10801,N_10866);
xnor U10926 (N_10926,N_10862,N_10800);
nor U10927 (N_10927,N_10849,N_10820);
and U10928 (N_10928,N_10854,N_10758);
nor U10929 (N_10929,N_10773,N_10867);
and U10930 (N_10930,N_10803,N_10865);
or U10931 (N_10931,N_10873,N_10792);
xor U10932 (N_10932,N_10759,N_10785);
or U10933 (N_10933,N_10810,N_10802);
nor U10934 (N_10934,N_10765,N_10848);
xnor U10935 (N_10935,N_10779,N_10777);
nor U10936 (N_10936,N_10767,N_10791);
xor U10937 (N_10937,N_10756,N_10813);
or U10938 (N_10938,N_10844,N_10754);
xnor U10939 (N_10939,N_10806,N_10792);
or U10940 (N_10940,N_10847,N_10824);
nor U10941 (N_10941,N_10765,N_10846);
xor U10942 (N_10942,N_10854,N_10827);
nor U10943 (N_10943,N_10774,N_10815);
or U10944 (N_10944,N_10782,N_10834);
nand U10945 (N_10945,N_10835,N_10811);
nand U10946 (N_10946,N_10815,N_10780);
nor U10947 (N_10947,N_10796,N_10770);
and U10948 (N_10948,N_10785,N_10790);
nand U10949 (N_10949,N_10852,N_10855);
or U10950 (N_10950,N_10849,N_10852);
or U10951 (N_10951,N_10765,N_10835);
nand U10952 (N_10952,N_10787,N_10829);
nor U10953 (N_10953,N_10760,N_10775);
nor U10954 (N_10954,N_10759,N_10773);
xnor U10955 (N_10955,N_10818,N_10760);
nor U10956 (N_10956,N_10756,N_10810);
nand U10957 (N_10957,N_10840,N_10862);
nand U10958 (N_10958,N_10838,N_10750);
xnor U10959 (N_10959,N_10809,N_10854);
nor U10960 (N_10960,N_10769,N_10849);
nor U10961 (N_10961,N_10837,N_10835);
nor U10962 (N_10962,N_10756,N_10774);
or U10963 (N_10963,N_10864,N_10812);
nor U10964 (N_10964,N_10835,N_10830);
xor U10965 (N_10965,N_10825,N_10766);
nor U10966 (N_10966,N_10750,N_10816);
xnor U10967 (N_10967,N_10773,N_10808);
and U10968 (N_10968,N_10849,N_10824);
and U10969 (N_10969,N_10850,N_10779);
nor U10970 (N_10970,N_10840,N_10854);
nand U10971 (N_10971,N_10847,N_10846);
nand U10972 (N_10972,N_10751,N_10848);
and U10973 (N_10973,N_10872,N_10760);
and U10974 (N_10974,N_10832,N_10819);
and U10975 (N_10975,N_10868,N_10872);
nand U10976 (N_10976,N_10848,N_10778);
nor U10977 (N_10977,N_10763,N_10840);
xnor U10978 (N_10978,N_10866,N_10818);
xor U10979 (N_10979,N_10845,N_10857);
and U10980 (N_10980,N_10826,N_10821);
nor U10981 (N_10981,N_10767,N_10838);
and U10982 (N_10982,N_10840,N_10760);
xnor U10983 (N_10983,N_10758,N_10848);
nand U10984 (N_10984,N_10781,N_10851);
nor U10985 (N_10985,N_10835,N_10814);
xnor U10986 (N_10986,N_10818,N_10872);
and U10987 (N_10987,N_10817,N_10847);
or U10988 (N_10988,N_10801,N_10811);
and U10989 (N_10989,N_10764,N_10802);
xor U10990 (N_10990,N_10850,N_10757);
nand U10991 (N_10991,N_10866,N_10777);
and U10992 (N_10992,N_10827,N_10833);
and U10993 (N_10993,N_10762,N_10766);
nor U10994 (N_10994,N_10802,N_10853);
nand U10995 (N_10995,N_10794,N_10836);
nand U10996 (N_10996,N_10799,N_10750);
nor U10997 (N_10997,N_10808,N_10821);
and U10998 (N_10998,N_10873,N_10766);
or U10999 (N_10999,N_10872,N_10809);
xnor U11000 (N_11000,N_10924,N_10901);
nand U11001 (N_11001,N_10923,N_10987);
or U11002 (N_11002,N_10970,N_10892);
nand U11003 (N_11003,N_10975,N_10954);
xor U11004 (N_11004,N_10878,N_10927);
nand U11005 (N_11005,N_10905,N_10896);
and U11006 (N_11006,N_10944,N_10971);
nand U11007 (N_11007,N_10981,N_10952);
nor U11008 (N_11008,N_10904,N_10957);
nor U11009 (N_11009,N_10928,N_10883);
xor U11010 (N_11010,N_10902,N_10933);
and U11011 (N_11011,N_10897,N_10940);
xnor U11012 (N_11012,N_10964,N_10920);
nor U11013 (N_11013,N_10882,N_10982);
and U11014 (N_11014,N_10906,N_10900);
nand U11015 (N_11015,N_10991,N_10946);
xor U11016 (N_11016,N_10989,N_10936);
nand U11017 (N_11017,N_10993,N_10886);
nand U11018 (N_11018,N_10889,N_10921);
xor U11019 (N_11019,N_10979,N_10942);
and U11020 (N_11020,N_10912,N_10876);
nor U11021 (N_11021,N_10884,N_10926);
and U11022 (N_11022,N_10894,N_10974);
and U11023 (N_11023,N_10955,N_10907);
nor U11024 (N_11024,N_10918,N_10973);
and U11025 (N_11025,N_10895,N_10903);
or U11026 (N_11026,N_10958,N_10875);
nor U11027 (N_11027,N_10985,N_10961);
nor U11028 (N_11028,N_10947,N_10916);
xnor U11029 (N_11029,N_10996,N_10948);
or U11030 (N_11030,N_10934,N_10931);
xnor U11031 (N_11031,N_10925,N_10890);
xor U11032 (N_11032,N_10966,N_10891);
or U11033 (N_11033,N_10994,N_10950);
nand U11034 (N_11034,N_10898,N_10909);
xnor U11035 (N_11035,N_10932,N_10963);
or U11036 (N_11036,N_10976,N_10984);
xnor U11037 (N_11037,N_10888,N_10986);
nor U11038 (N_11038,N_10917,N_10911);
or U11039 (N_11039,N_10951,N_10965);
and U11040 (N_11040,N_10879,N_10945);
nand U11041 (N_11041,N_10930,N_10938);
and U11042 (N_11042,N_10943,N_10929);
and U11043 (N_11043,N_10968,N_10969);
nand U11044 (N_11044,N_10983,N_10978);
nor U11045 (N_11045,N_10893,N_10992);
xor U11046 (N_11046,N_10922,N_10962);
or U11047 (N_11047,N_10919,N_10995);
xor U11048 (N_11048,N_10939,N_10960);
nand U11049 (N_11049,N_10877,N_10908);
and U11050 (N_11050,N_10913,N_10959);
or U11051 (N_11051,N_10988,N_10972);
or U11052 (N_11052,N_10880,N_10941);
and U11053 (N_11053,N_10887,N_10881);
xnor U11054 (N_11054,N_10953,N_10999);
or U11055 (N_11055,N_10937,N_10914);
nand U11056 (N_11056,N_10935,N_10980);
or U11057 (N_11057,N_10997,N_10977);
and U11058 (N_11058,N_10899,N_10885);
nor U11059 (N_11059,N_10990,N_10949);
xor U11060 (N_11060,N_10915,N_10967);
and U11061 (N_11061,N_10910,N_10956);
nor U11062 (N_11062,N_10998,N_10989);
and U11063 (N_11063,N_10901,N_10891);
xnor U11064 (N_11064,N_10882,N_10983);
nand U11065 (N_11065,N_10895,N_10905);
xor U11066 (N_11066,N_10933,N_10927);
nor U11067 (N_11067,N_10981,N_10910);
or U11068 (N_11068,N_10889,N_10987);
nand U11069 (N_11069,N_10950,N_10995);
and U11070 (N_11070,N_10890,N_10921);
or U11071 (N_11071,N_10977,N_10911);
nand U11072 (N_11072,N_10966,N_10930);
nor U11073 (N_11073,N_10959,N_10881);
nand U11074 (N_11074,N_10918,N_10916);
and U11075 (N_11075,N_10898,N_10900);
xnor U11076 (N_11076,N_10935,N_10939);
nor U11077 (N_11077,N_10950,N_10989);
nor U11078 (N_11078,N_10898,N_10999);
nand U11079 (N_11079,N_10918,N_10928);
and U11080 (N_11080,N_10908,N_10940);
xor U11081 (N_11081,N_10912,N_10893);
or U11082 (N_11082,N_10972,N_10897);
or U11083 (N_11083,N_10901,N_10978);
and U11084 (N_11084,N_10933,N_10901);
nand U11085 (N_11085,N_10887,N_10979);
or U11086 (N_11086,N_10962,N_10996);
nor U11087 (N_11087,N_10923,N_10875);
and U11088 (N_11088,N_10931,N_10979);
or U11089 (N_11089,N_10877,N_10878);
xor U11090 (N_11090,N_10990,N_10923);
nand U11091 (N_11091,N_10877,N_10987);
nand U11092 (N_11092,N_10953,N_10979);
nor U11093 (N_11093,N_10938,N_10918);
or U11094 (N_11094,N_10957,N_10915);
nor U11095 (N_11095,N_10884,N_10956);
nand U11096 (N_11096,N_10878,N_10920);
nand U11097 (N_11097,N_10938,N_10943);
or U11098 (N_11098,N_10985,N_10942);
and U11099 (N_11099,N_10921,N_10877);
nor U11100 (N_11100,N_10914,N_10902);
or U11101 (N_11101,N_10952,N_10937);
nand U11102 (N_11102,N_10961,N_10965);
nor U11103 (N_11103,N_10914,N_10985);
and U11104 (N_11104,N_10926,N_10961);
xor U11105 (N_11105,N_10954,N_10993);
or U11106 (N_11106,N_10957,N_10879);
nand U11107 (N_11107,N_10979,N_10982);
xor U11108 (N_11108,N_10908,N_10973);
nand U11109 (N_11109,N_10916,N_10997);
or U11110 (N_11110,N_10993,N_10882);
nor U11111 (N_11111,N_10978,N_10997);
or U11112 (N_11112,N_10898,N_10956);
nor U11113 (N_11113,N_10957,N_10987);
nor U11114 (N_11114,N_10909,N_10998);
nor U11115 (N_11115,N_10999,N_10948);
and U11116 (N_11116,N_10990,N_10950);
nand U11117 (N_11117,N_10899,N_10884);
and U11118 (N_11118,N_10932,N_10951);
nor U11119 (N_11119,N_10877,N_10916);
nand U11120 (N_11120,N_10877,N_10883);
nand U11121 (N_11121,N_10977,N_10967);
xor U11122 (N_11122,N_10961,N_10938);
and U11123 (N_11123,N_10932,N_10876);
or U11124 (N_11124,N_10981,N_10990);
or U11125 (N_11125,N_11092,N_11101);
or U11126 (N_11126,N_11048,N_11034);
and U11127 (N_11127,N_11069,N_11041);
nand U11128 (N_11128,N_11060,N_11036);
nand U11129 (N_11129,N_11066,N_11065);
nor U11130 (N_11130,N_11022,N_11073);
xnor U11131 (N_11131,N_11072,N_11021);
and U11132 (N_11132,N_11054,N_11010);
nand U11133 (N_11133,N_11017,N_11042);
nand U11134 (N_11134,N_11002,N_11074);
xor U11135 (N_11135,N_11059,N_11044);
and U11136 (N_11136,N_11116,N_11085);
xnor U11137 (N_11137,N_11061,N_11111);
and U11138 (N_11138,N_11071,N_11007);
nand U11139 (N_11139,N_11086,N_11013);
nand U11140 (N_11140,N_11016,N_11009);
nor U11141 (N_11141,N_11051,N_11115);
nand U11142 (N_11142,N_11000,N_11063);
or U11143 (N_11143,N_11120,N_11037);
xnor U11144 (N_11144,N_11090,N_11075);
or U11145 (N_11145,N_11113,N_11121);
and U11146 (N_11146,N_11100,N_11099);
or U11147 (N_11147,N_11083,N_11039);
and U11148 (N_11148,N_11027,N_11089);
xor U11149 (N_11149,N_11028,N_11064);
nor U11150 (N_11150,N_11106,N_11040);
and U11151 (N_11151,N_11080,N_11087);
nand U11152 (N_11152,N_11038,N_11081);
nand U11153 (N_11153,N_11045,N_11114);
nor U11154 (N_11154,N_11097,N_11110);
nand U11155 (N_11155,N_11014,N_11043);
xor U11156 (N_11156,N_11124,N_11107);
and U11157 (N_11157,N_11095,N_11091);
xor U11158 (N_11158,N_11033,N_11082);
nor U11159 (N_11159,N_11070,N_11122);
or U11160 (N_11160,N_11102,N_11020);
nor U11161 (N_11161,N_11093,N_11052);
and U11162 (N_11162,N_11077,N_11109);
nor U11163 (N_11163,N_11112,N_11050);
nor U11164 (N_11164,N_11118,N_11105);
xnor U11165 (N_11165,N_11053,N_11096);
xnor U11166 (N_11166,N_11015,N_11057);
or U11167 (N_11167,N_11098,N_11049);
xnor U11168 (N_11168,N_11119,N_11046);
or U11169 (N_11169,N_11123,N_11006);
xnor U11170 (N_11170,N_11108,N_11068);
nor U11171 (N_11171,N_11067,N_11078);
and U11172 (N_11172,N_11103,N_11084);
nand U11173 (N_11173,N_11079,N_11062);
nor U11174 (N_11174,N_11024,N_11094);
nand U11175 (N_11175,N_11001,N_11032);
and U11176 (N_11176,N_11008,N_11117);
and U11177 (N_11177,N_11018,N_11029);
and U11178 (N_11178,N_11104,N_11025);
or U11179 (N_11179,N_11031,N_11003);
and U11180 (N_11180,N_11004,N_11058);
nand U11181 (N_11181,N_11030,N_11011);
nor U11182 (N_11182,N_11088,N_11056);
or U11183 (N_11183,N_11012,N_11023);
and U11184 (N_11184,N_11055,N_11026);
and U11185 (N_11185,N_11005,N_11076);
and U11186 (N_11186,N_11035,N_11047);
xnor U11187 (N_11187,N_11019,N_11119);
nand U11188 (N_11188,N_11114,N_11049);
or U11189 (N_11189,N_11004,N_11078);
and U11190 (N_11190,N_11096,N_11010);
or U11191 (N_11191,N_11115,N_11123);
and U11192 (N_11192,N_11101,N_11056);
and U11193 (N_11193,N_11103,N_11034);
nand U11194 (N_11194,N_11004,N_11052);
xor U11195 (N_11195,N_11057,N_11038);
and U11196 (N_11196,N_11121,N_11058);
xnor U11197 (N_11197,N_11028,N_11090);
and U11198 (N_11198,N_11070,N_11102);
nand U11199 (N_11199,N_11031,N_11004);
or U11200 (N_11200,N_11043,N_11108);
xnor U11201 (N_11201,N_11117,N_11021);
xnor U11202 (N_11202,N_11050,N_11015);
and U11203 (N_11203,N_11106,N_11094);
nand U11204 (N_11204,N_11084,N_11058);
and U11205 (N_11205,N_11043,N_11071);
xor U11206 (N_11206,N_11075,N_11062);
nor U11207 (N_11207,N_11121,N_11050);
xor U11208 (N_11208,N_11045,N_11110);
xnor U11209 (N_11209,N_11033,N_11092);
or U11210 (N_11210,N_11058,N_11070);
or U11211 (N_11211,N_11064,N_11037);
and U11212 (N_11212,N_11078,N_11070);
xor U11213 (N_11213,N_11033,N_11049);
nand U11214 (N_11214,N_11054,N_11102);
and U11215 (N_11215,N_11079,N_11111);
and U11216 (N_11216,N_11090,N_11021);
and U11217 (N_11217,N_11045,N_11031);
xor U11218 (N_11218,N_11065,N_11045);
or U11219 (N_11219,N_11008,N_11005);
xnor U11220 (N_11220,N_11123,N_11095);
and U11221 (N_11221,N_11070,N_11040);
or U11222 (N_11222,N_11060,N_11075);
xor U11223 (N_11223,N_11029,N_11073);
nand U11224 (N_11224,N_11008,N_11030);
xnor U11225 (N_11225,N_11036,N_11099);
and U11226 (N_11226,N_11032,N_11062);
xor U11227 (N_11227,N_11114,N_11059);
and U11228 (N_11228,N_11059,N_11071);
nand U11229 (N_11229,N_11065,N_11086);
nand U11230 (N_11230,N_11002,N_11026);
nand U11231 (N_11231,N_11123,N_11032);
and U11232 (N_11232,N_11019,N_11095);
nor U11233 (N_11233,N_11076,N_11068);
or U11234 (N_11234,N_11075,N_11051);
nor U11235 (N_11235,N_11118,N_11116);
nor U11236 (N_11236,N_11106,N_11035);
and U11237 (N_11237,N_11099,N_11004);
nand U11238 (N_11238,N_11001,N_11035);
nand U11239 (N_11239,N_11082,N_11055);
and U11240 (N_11240,N_11123,N_11085);
or U11241 (N_11241,N_11035,N_11118);
nor U11242 (N_11242,N_11108,N_11046);
or U11243 (N_11243,N_11123,N_11057);
xnor U11244 (N_11244,N_11043,N_11052);
nor U11245 (N_11245,N_11042,N_11062);
or U11246 (N_11246,N_11076,N_11066);
nand U11247 (N_11247,N_11004,N_11091);
xor U11248 (N_11248,N_11100,N_11031);
nand U11249 (N_11249,N_11083,N_11084);
nor U11250 (N_11250,N_11234,N_11172);
and U11251 (N_11251,N_11152,N_11212);
nor U11252 (N_11252,N_11247,N_11213);
or U11253 (N_11253,N_11197,N_11216);
nor U11254 (N_11254,N_11170,N_11161);
and U11255 (N_11255,N_11184,N_11174);
nand U11256 (N_11256,N_11147,N_11249);
or U11257 (N_11257,N_11203,N_11201);
nand U11258 (N_11258,N_11204,N_11205);
xor U11259 (N_11259,N_11230,N_11202);
nand U11260 (N_11260,N_11208,N_11138);
xor U11261 (N_11261,N_11215,N_11178);
or U11262 (N_11262,N_11148,N_11164);
xor U11263 (N_11263,N_11224,N_11126);
xor U11264 (N_11264,N_11218,N_11166);
nor U11265 (N_11265,N_11207,N_11221);
nand U11266 (N_11266,N_11136,N_11157);
nor U11267 (N_11267,N_11156,N_11153);
and U11268 (N_11268,N_11169,N_11143);
xnor U11269 (N_11269,N_11195,N_11185);
and U11270 (N_11270,N_11125,N_11181);
xor U11271 (N_11271,N_11248,N_11127);
nor U11272 (N_11272,N_11193,N_11162);
and U11273 (N_11273,N_11151,N_11241);
or U11274 (N_11274,N_11159,N_11155);
nand U11275 (N_11275,N_11149,N_11217);
nor U11276 (N_11276,N_11209,N_11236);
xnor U11277 (N_11277,N_11200,N_11226);
xor U11278 (N_11278,N_11173,N_11239);
xor U11279 (N_11279,N_11129,N_11139);
nor U11280 (N_11280,N_11187,N_11237);
nor U11281 (N_11281,N_11135,N_11219);
or U11282 (N_11282,N_11154,N_11182);
and U11283 (N_11283,N_11214,N_11235);
xnor U11284 (N_11284,N_11171,N_11176);
or U11285 (N_11285,N_11131,N_11243);
xor U11286 (N_11286,N_11229,N_11186);
nand U11287 (N_11287,N_11191,N_11150);
xnor U11288 (N_11288,N_11198,N_11165);
nand U11289 (N_11289,N_11194,N_11188);
and U11290 (N_11290,N_11206,N_11175);
and U11291 (N_11291,N_11223,N_11245);
nand U11292 (N_11292,N_11177,N_11128);
and U11293 (N_11293,N_11225,N_11231);
nand U11294 (N_11294,N_11130,N_11190);
nor U11295 (N_11295,N_11158,N_11242);
and U11296 (N_11296,N_11233,N_11145);
nor U11297 (N_11297,N_11246,N_11220);
and U11298 (N_11298,N_11160,N_11168);
xor U11299 (N_11299,N_11132,N_11142);
nor U11300 (N_11300,N_11167,N_11211);
nand U11301 (N_11301,N_11240,N_11144);
nand U11302 (N_11302,N_11140,N_11232);
or U11303 (N_11303,N_11244,N_11163);
and U11304 (N_11304,N_11222,N_11183);
nor U11305 (N_11305,N_11134,N_11196);
nor U11306 (N_11306,N_11210,N_11228);
nor U11307 (N_11307,N_11192,N_11238);
and U11308 (N_11308,N_11133,N_11137);
or U11309 (N_11309,N_11199,N_11146);
or U11310 (N_11310,N_11179,N_11227);
nor U11311 (N_11311,N_11141,N_11180);
or U11312 (N_11312,N_11189,N_11229);
and U11313 (N_11313,N_11223,N_11240);
or U11314 (N_11314,N_11245,N_11147);
nor U11315 (N_11315,N_11186,N_11207);
nand U11316 (N_11316,N_11182,N_11244);
and U11317 (N_11317,N_11164,N_11163);
nand U11318 (N_11318,N_11208,N_11135);
xor U11319 (N_11319,N_11200,N_11248);
and U11320 (N_11320,N_11227,N_11240);
or U11321 (N_11321,N_11156,N_11125);
xor U11322 (N_11322,N_11207,N_11183);
and U11323 (N_11323,N_11204,N_11237);
nor U11324 (N_11324,N_11160,N_11213);
xor U11325 (N_11325,N_11127,N_11126);
nor U11326 (N_11326,N_11155,N_11182);
xnor U11327 (N_11327,N_11229,N_11147);
and U11328 (N_11328,N_11202,N_11188);
nor U11329 (N_11329,N_11137,N_11209);
nor U11330 (N_11330,N_11215,N_11165);
xnor U11331 (N_11331,N_11234,N_11156);
or U11332 (N_11332,N_11198,N_11247);
nand U11333 (N_11333,N_11137,N_11244);
xor U11334 (N_11334,N_11184,N_11224);
xor U11335 (N_11335,N_11171,N_11133);
nand U11336 (N_11336,N_11226,N_11213);
or U11337 (N_11337,N_11168,N_11150);
xor U11338 (N_11338,N_11156,N_11189);
and U11339 (N_11339,N_11246,N_11200);
or U11340 (N_11340,N_11160,N_11151);
nand U11341 (N_11341,N_11159,N_11209);
nand U11342 (N_11342,N_11235,N_11236);
nor U11343 (N_11343,N_11143,N_11191);
nand U11344 (N_11344,N_11136,N_11194);
or U11345 (N_11345,N_11128,N_11170);
nand U11346 (N_11346,N_11133,N_11233);
and U11347 (N_11347,N_11140,N_11230);
and U11348 (N_11348,N_11183,N_11184);
and U11349 (N_11349,N_11234,N_11219);
nand U11350 (N_11350,N_11184,N_11189);
and U11351 (N_11351,N_11236,N_11190);
nor U11352 (N_11352,N_11209,N_11131);
nand U11353 (N_11353,N_11225,N_11146);
nor U11354 (N_11354,N_11194,N_11231);
or U11355 (N_11355,N_11163,N_11194);
or U11356 (N_11356,N_11198,N_11249);
nor U11357 (N_11357,N_11143,N_11128);
or U11358 (N_11358,N_11176,N_11238);
nand U11359 (N_11359,N_11168,N_11172);
xor U11360 (N_11360,N_11138,N_11184);
and U11361 (N_11361,N_11235,N_11134);
xor U11362 (N_11362,N_11206,N_11160);
nor U11363 (N_11363,N_11247,N_11138);
or U11364 (N_11364,N_11131,N_11128);
nand U11365 (N_11365,N_11143,N_11181);
and U11366 (N_11366,N_11161,N_11234);
and U11367 (N_11367,N_11192,N_11169);
or U11368 (N_11368,N_11181,N_11236);
or U11369 (N_11369,N_11193,N_11216);
nor U11370 (N_11370,N_11156,N_11226);
xor U11371 (N_11371,N_11163,N_11140);
or U11372 (N_11372,N_11171,N_11157);
and U11373 (N_11373,N_11186,N_11212);
or U11374 (N_11374,N_11248,N_11203);
and U11375 (N_11375,N_11369,N_11261);
nor U11376 (N_11376,N_11265,N_11331);
and U11377 (N_11377,N_11338,N_11286);
or U11378 (N_11378,N_11323,N_11270);
nor U11379 (N_11379,N_11357,N_11361);
nand U11380 (N_11380,N_11333,N_11267);
nor U11381 (N_11381,N_11312,N_11302);
nand U11382 (N_11382,N_11356,N_11332);
xnor U11383 (N_11383,N_11273,N_11274);
and U11384 (N_11384,N_11340,N_11282);
nand U11385 (N_11385,N_11255,N_11280);
nor U11386 (N_11386,N_11314,N_11253);
or U11387 (N_11387,N_11349,N_11343);
or U11388 (N_11388,N_11305,N_11359);
nand U11389 (N_11389,N_11345,N_11278);
nand U11390 (N_11390,N_11327,N_11362);
nor U11391 (N_11391,N_11366,N_11372);
nand U11392 (N_11392,N_11289,N_11354);
nor U11393 (N_11393,N_11317,N_11296);
or U11394 (N_11394,N_11271,N_11320);
or U11395 (N_11395,N_11324,N_11308);
xnor U11396 (N_11396,N_11350,N_11304);
or U11397 (N_11397,N_11330,N_11365);
or U11398 (N_11398,N_11313,N_11287);
xnor U11399 (N_11399,N_11281,N_11341);
or U11400 (N_11400,N_11272,N_11326);
nor U11401 (N_11401,N_11254,N_11318);
nor U11402 (N_11402,N_11279,N_11315);
and U11403 (N_11403,N_11351,N_11353);
nand U11404 (N_11404,N_11373,N_11262);
and U11405 (N_11405,N_11346,N_11309);
nor U11406 (N_11406,N_11290,N_11339);
and U11407 (N_11407,N_11257,N_11358);
or U11408 (N_11408,N_11371,N_11367);
nor U11409 (N_11409,N_11301,N_11329);
nor U11410 (N_11410,N_11260,N_11364);
nor U11411 (N_11411,N_11321,N_11292);
or U11412 (N_11412,N_11275,N_11285);
and U11413 (N_11413,N_11355,N_11250);
or U11414 (N_11414,N_11336,N_11298);
or U11415 (N_11415,N_11316,N_11276);
or U11416 (N_11416,N_11348,N_11335);
xnor U11417 (N_11417,N_11295,N_11306);
and U11418 (N_11418,N_11363,N_11297);
nor U11419 (N_11419,N_11300,N_11252);
nor U11420 (N_11420,N_11251,N_11368);
and U11421 (N_11421,N_11334,N_11344);
and U11422 (N_11422,N_11269,N_11283);
nand U11423 (N_11423,N_11299,N_11352);
nor U11424 (N_11424,N_11319,N_11322);
and U11425 (N_11425,N_11288,N_11310);
and U11426 (N_11426,N_11284,N_11263);
nor U11427 (N_11427,N_11294,N_11311);
and U11428 (N_11428,N_11256,N_11325);
xor U11429 (N_11429,N_11258,N_11303);
or U11430 (N_11430,N_11370,N_11347);
nand U11431 (N_11431,N_11328,N_11277);
xnor U11432 (N_11432,N_11268,N_11360);
and U11433 (N_11433,N_11291,N_11342);
xor U11434 (N_11434,N_11259,N_11374);
or U11435 (N_11435,N_11264,N_11307);
nor U11436 (N_11436,N_11337,N_11293);
and U11437 (N_11437,N_11266,N_11310);
nor U11438 (N_11438,N_11359,N_11326);
nor U11439 (N_11439,N_11296,N_11291);
xor U11440 (N_11440,N_11363,N_11337);
or U11441 (N_11441,N_11266,N_11320);
xnor U11442 (N_11442,N_11285,N_11373);
or U11443 (N_11443,N_11284,N_11365);
nand U11444 (N_11444,N_11262,N_11276);
nor U11445 (N_11445,N_11305,N_11288);
and U11446 (N_11446,N_11302,N_11326);
and U11447 (N_11447,N_11331,N_11316);
and U11448 (N_11448,N_11297,N_11277);
nor U11449 (N_11449,N_11360,N_11372);
nand U11450 (N_11450,N_11298,N_11332);
nand U11451 (N_11451,N_11347,N_11373);
and U11452 (N_11452,N_11297,N_11319);
xnor U11453 (N_11453,N_11313,N_11285);
or U11454 (N_11454,N_11359,N_11337);
xor U11455 (N_11455,N_11295,N_11272);
and U11456 (N_11456,N_11250,N_11276);
or U11457 (N_11457,N_11305,N_11315);
nand U11458 (N_11458,N_11336,N_11303);
and U11459 (N_11459,N_11265,N_11322);
nand U11460 (N_11460,N_11338,N_11257);
and U11461 (N_11461,N_11350,N_11279);
nor U11462 (N_11462,N_11267,N_11340);
xor U11463 (N_11463,N_11255,N_11310);
nor U11464 (N_11464,N_11293,N_11343);
nor U11465 (N_11465,N_11338,N_11316);
xor U11466 (N_11466,N_11306,N_11250);
and U11467 (N_11467,N_11370,N_11280);
nor U11468 (N_11468,N_11316,N_11368);
or U11469 (N_11469,N_11314,N_11286);
nand U11470 (N_11470,N_11331,N_11271);
nand U11471 (N_11471,N_11276,N_11365);
and U11472 (N_11472,N_11304,N_11296);
or U11473 (N_11473,N_11359,N_11339);
xor U11474 (N_11474,N_11269,N_11268);
nor U11475 (N_11475,N_11318,N_11367);
and U11476 (N_11476,N_11342,N_11325);
nor U11477 (N_11477,N_11372,N_11370);
or U11478 (N_11478,N_11282,N_11361);
or U11479 (N_11479,N_11365,N_11302);
nand U11480 (N_11480,N_11306,N_11270);
and U11481 (N_11481,N_11319,N_11309);
nor U11482 (N_11482,N_11287,N_11289);
nand U11483 (N_11483,N_11308,N_11304);
and U11484 (N_11484,N_11323,N_11296);
or U11485 (N_11485,N_11328,N_11336);
and U11486 (N_11486,N_11260,N_11373);
nor U11487 (N_11487,N_11346,N_11274);
or U11488 (N_11488,N_11251,N_11292);
and U11489 (N_11489,N_11308,N_11334);
nand U11490 (N_11490,N_11371,N_11286);
xnor U11491 (N_11491,N_11293,N_11275);
xor U11492 (N_11492,N_11327,N_11318);
xnor U11493 (N_11493,N_11275,N_11353);
or U11494 (N_11494,N_11347,N_11356);
xnor U11495 (N_11495,N_11267,N_11352);
or U11496 (N_11496,N_11370,N_11312);
or U11497 (N_11497,N_11351,N_11263);
xor U11498 (N_11498,N_11362,N_11351);
and U11499 (N_11499,N_11271,N_11267);
or U11500 (N_11500,N_11457,N_11476);
xor U11501 (N_11501,N_11430,N_11408);
xnor U11502 (N_11502,N_11467,N_11394);
xnor U11503 (N_11503,N_11407,N_11490);
nand U11504 (N_11504,N_11381,N_11427);
nand U11505 (N_11505,N_11429,N_11482);
xnor U11506 (N_11506,N_11413,N_11480);
and U11507 (N_11507,N_11387,N_11449);
xnor U11508 (N_11508,N_11473,N_11399);
nor U11509 (N_11509,N_11410,N_11425);
nor U11510 (N_11510,N_11405,N_11441);
or U11511 (N_11511,N_11419,N_11404);
xor U11512 (N_11512,N_11483,N_11389);
nor U11513 (N_11513,N_11395,N_11421);
nand U11514 (N_11514,N_11448,N_11468);
nor U11515 (N_11515,N_11420,N_11378);
nor U11516 (N_11516,N_11401,N_11451);
and U11517 (N_11517,N_11495,N_11440);
nor U11518 (N_11518,N_11388,N_11385);
xnor U11519 (N_11519,N_11475,N_11426);
nand U11520 (N_11520,N_11443,N_11431);
and U11521 (N_11521,N_11479,N_11498);
xnor U11522 (N_11522,N_11390,N_11439);
nand U11523 (N_11523,N_11391,N_11481);
and U11524 (N_11524,N_11403,N_11424);
or U11525 (N_11525,N_11469,N_11492);
and U11526 (N_11526,N_11471,N_11465);
nor U11527 (N_11527,N_11438,N_11422);
nor U11528 (N_11528,N_11459,N_11461);
nor U11529 (N_11529,N_11485,N_11428);
xnor U11530 (N_11530,N_11484,N_11411);
xor U11531 (N_11531,N_11392,N_11382);
or U11532 (N_11532,N_11463,N_11446);
nand U11533 (N_11533,N_11418,N_11460);
nor U11534 (N_11534,N_11400,N_11486);
nor U11535 (N_11535,N_11496,N_11435);
and U11536 (N_11536,N_11377,N_11452);
nor U11537 (N_11537,N_11489,N_11383);
and U11538 (N_11538,N_11445,N_11409);
nand U11539 (N_11539,N_11444,N_11432);
nor U11540 (N_11540,N_11380,N_11393);
xor U11541 (N_11541,N_11375,N_11499);
xnor U11542 (N_11542,N_11474,N_11453);
or U11543 (N_11543,N_11470,N_11493);
or U11544 (N_11544,N_11491,N_11433);
or U11545 (N_11545,N_11472,N_11488);
nor U11546 (N_11546,N_11466,N_11376);
xor U11547 (N_11547,N_11417,N_11406);
and U11548 (N_11548,N_11436,N_11462);
or U11549 (N_11549,N_11416,N_11398);
and U11550 (N_11550,N_11497,N_11379);
xor U11551 (N_11551,N_11384,N_11478);
xor U11552 (N_11552,N_11414,N_11396);
or U11553 (N_11553,N_11455,N_11477);
or U11554 (N_11554,N_11412,N_11464);
nand U11555 (N_11555,N_11487,N_11397);
xor U11556 (N_11556,N_11458,N_11386);
and U11557 (N_11557,N_11447,N_11442);
xor U11558 (N_11558,N_11402,N_11454);
and U11559 (N_11559,N_11494,N_11437);
or U11560 (N_11560,N_11423,N_11456);
nor U11561 (N_11561,N_11434,N_11415);
nand U11562 (N_11562,N_11450,N_11481);
or U11563 (N_11563,N_11463,N_11455);
or U11564 (N_11564,N_11456,N_11436);
and U11565 (N_11565,N_11399,N_11430);
xor U11566 (N_11566,N_11402,N_11484);
or U11567 (N_11567,N_11441,N_11427);
nand U11568 (N_11568,N_11495,N_11466);
or U11569 (N_11569,N_11434,N_11451);
nand U11570 (N_11570,N_11445,N_11382);
nor U11571 (N_11571,N_11477,N_11472);
nor U11572 (N_11572,N_11488,N_11381);
xor U11573 (N_11573,N_11479,N_11397);
nor U11574 (N_11574,N_11414,N_11446);
nand U11575 (N_11575,N_11392,N_11404);
nand U11576 (N_11576,N_11461,N_11450);
and U11577 (N_11577,N_11444,N_11410);
or U11578 (N_11578,N_11468,N_11455);
xor U11579 (N_11579,N_11387,N_11441);
or U11580 (N_11580,N_11461,N_11464);
or U11581 (N_11581,N_11479,N_11379);
or U11582 (N_11582,N_11421,N_11410);
xnor U11583 (N_11583,N_11482,N_11395);
or U11584 (N_11584,N_11393,N_11428);
nor U11585 (N_11585,N_11492,N_11408);
or U11586 (N_11586,N_11384,N_11472);
and U11587 (N_11587,N_11409,N_11488);
nand U11588 (N_11588,N_11489,N_11455);
nor U11589 (N_11589,N_11381,N_11491);
and U11590 (N_11590,N_11388,N_11468);
nor U11591 (N_11591,N_11486,N_11423);
xnor U11592 (N_11592,N_11422,N_11433);
nand U11593 (N_11593,N_11441,N_11481);
nand U11594 (N_11594,N_11394,N_11456);
xor U11595 (N_11595,N_11459,N_11409);
or U11596 (N_11596,N_11476,N_11492);
xor U11597 (N_11597,N_11457,N_11438);
and U11598 (N_11598,N_11430,N_11415);
nand U11599 (N_11599,N_11451,N_11380);
xor U11600 (N_11600,N_11395,N_11397);
and U11601 (N_11601,N_11490,N_11421);
and U11602 (N_11602,N_11430,N_11392);
or U11603 (N_11603,N_11423,N_11412);
or U11604 (N_11604,N_11391,N_11392);
and U11605 (N_11605,N_11472,N_11412);
nand U11606 (N_11606,N_11378,N_11485);
and U11607 (N_11607,N_11408,N_11415);
and U11608 (N_11608,N_11382,N_11487);
nor U11609 (N_11609,N_11402,N_11476);
xnor U11610 (N_11610,N_11483,N_11482);
nand U11611 (N_11611,N_11400,N_11454);
or U11612 (N_11612,N_11465,N_11415);
xor U11613 (N_11613,N_11463,N_11403);
or U11614 (N_11614,N_11442,N_11396);
or U11615 (N_11615,N_11451,N_11449);
nand U11616 (N_11616,N_11384,N_11439);
nand U11617 (N_11617,N_11381,N_11470);
nand U11618 (N_11618,N_11490,N_11420);
or U11619 (N_11619,N_11439,N_11397);
nor U11620 (N_11620,N_11456,N_11478);
and U11621 (N_11621,N_11379,N_11413);
xor U11622 (N_11622,N_11376,N_11442);
or U11623 (N_11623,N_11406,N_11424);
or U11624 (N_11624,N_11426,N_11413);
nand U11625 (N_11625,N_11564,N_11535);
nand U11626 (N_11626,N_11549,N_11604);
nand U11627 (N_11627,N_11586,N_11510);
or U11628 (N_11628,N_11527,N_11515);
nand U11629 (N_11629,N_11565,N_11605);
or U11630 (N_11630,N_11598,N_11542);
and U11631 (N_11631,N_11618,N_11592);
and U11632 (N_11632,N_11533,N_11546);
and U11633 (N_11633,N_11566,N_11610);
or U11634 (N_11634,N_11556,N_11525);
nand U11635 (N_11635,N_11537,N_11583);
and U11636 (N_11636,N_11591,N_11579);
xnor U11637 (N_11637,N_11528,N_11555);
nor U11638 (N_11638,N_11519,N_11585);
nor U11639 (N_11639,N_11589,N_11558);
or U11640 (N_11640,N_11569,N_11516);
nand U11641 (N_11641,N_11616,N_11547);
nand U11642 (N_11642,N_11577,N_11545);
nand U11643 (N_11643,N_11553,N_11521);
and U11644 (N_11644,N_11524,N_11582);
nor U11645 (N_11645,N_11600,N_11563);
xor U11646 (N_11646,N_11503,N_11595);
nor U11647 (N_11647,N_11580,N_11620);
nor U11648 (N_11648,N_11544,N_11619);
and U11649 (N_11649,N_11505,N_11613);
or U11650 (N_11650,N_11594,N_11504);
or U11651 (N_11651,N_11559,N_11514);
xnor U11652 (N_11652,N_11573,N_11506);
and U11653 (N_11653,N_11507,N_11623);
xnor U11654 (N_11654,N_11572,N_11614);
nor U11655 (N_11655,N_11590,N_11513);
nand U11656 (N_11656,N_11551,N_11540);
or U11657 (N_11657,N_11576,N_11612);
or U11658 (N_11658,N_11522,N_11541);
and U11659 (N_11659,N_11530,N_11509);
or U11660 (N_11660,N_11523,N_11607);
or U11661 (N_11661,N_11601,N_11529);
nand U11662 (N_11662,N_11539,N_11622);
nor U11663 (N_11663,N_11512,N_11532);
nand U11664 (N_11664,N_11603,N_11543);
nand U11665 (N_11665,N_11615,N_11575);
nor U11666 (N_11666,N_11606,N_11561);
or U11667 (N_11667,N_11560,N_11588);
and U11668 (N_11668,N_11526,N_11578);
nor U11669 (N_11669,N_11552,N_11520);
or U11670 (N_11670,N_11534,N_11584);
or U11671 (N_11671,N_11570,N_11557);
nand U11672 (N_11672,N_11502,N_11568);
or U11673 (N_11673,N_11596,N_11611);
and U11674 (N_11674,N_11593,N_11538);
nor U11675 (N_11675,N_11608,N_11500);
xor U11676 (N_11676,N_11562,N_11587);
nor U11677 (N_11677,N_11574,N_11531);
nor U11678 (N_11678,N_11581,N_11517);
nor U11679 (N_11679,N_11624,N_11599);
or U11680 (N_11680,N_11617,N_11501);
nand U11681 (N_11681,N_11554,N_11508);
or U11682 (N_11682,N_11550,N_11548);
nand U11683 (N_11683,N_11597,N_11518);
nand U11684 (N_11684,N_11536,N_11567);
xnor U11685 (N_11685,N_11511,N_11602);
and U11686 (N_11686,N_11571,N_11609);
nand U11687 (N_11687,N_11621,N_11575);
nor U11688 (N_11688,N_11535,N_11563);
xor U11689 (N_11689,N_11525,N_11521);
nand U11690 (N_11690,N_11615,N_11534);
and U11691 (N_11691,N_11566,N_11620);
xnor U11692 (N_11692,N_11546,N_11513);
or U11693 (N_11693,N_11530,N_11588);
nor U11694 (N_11694,N_11604,N_11509);
and U11695 (N_11695,N_11565,N_11578);
nand U11696 (N_11696,N_11610,N_11558);
and U11697 (N_11697,N_11609,N_11586);
or U11698 (N_11698,N_11511,N_11618);
and U11699 (N_11699,N_11565,N_11624);
or U11700 (N_11700,N_11610,N_11556);
xor U11701 (N_11701,N_11508,N_11556);
and U11702 (N_11702,N_11577,N_11519);
nor U11703 (N_11703,N_11615,N_11590);
and U11704 (N_11704,N_11506,N_11622);
or U11705 (N_11705,N_11605,N_11615);
nand U11706 (N_11706,N_11547,N_11600);
xor U11707 (N_11707,N_11573,N_11610);
xnor U11708 (N_11708,N_11551,N_11610);
nor U11709 (N_11709,N_11548,N_11552);
and U11710 (N_11710,N_11570,N_11599);
nor U11711 (N_11711,N_11619,N_11511);
nand U11712 (N_11712,N_11519,N_11588);
xor U11713 (N_11713,N_11610,N_11622);
and U11714 (N_11714,N_11582,N_11567);
nor U11715 (N_11715,N_11612,N_11611);
and U11716 (N_11716,N_11550,N_11606);
xnor U11717 (N_11717,N_11571,N_11573);
nor U11718 (N_11718,N_11570,N_11584);
xnor U11719 (N_11719,N_11551,N_11575);
and U11720 (N_11720,N_11551,N_11556);
xor U11721 (N_11721,N_11562,N_11620);
or U11722 (N_11722,N_11606,N_11526);
and U11723 (N_11723,N_11587,N_11577);
or U11724 (N_11724,N_11589,N_11504);
or U11725 (N_11725,N_11551,N_11509);
nand U11726 (N_11726,N_11521,N_11528);
or U11727 (N_11727,N_11513,N_11562);
and U11728 (N_11728,N_11511,N_11521);
xor U11729 (N_11729,N_11608,N_11577);
or U11730 (N_11730,N_11531,N_11560);
nor U11731 (N_11731,N_11559,N_11602);
nand U11732 (N_11732,N_11524,N_11601);
nand U11733 (N_11733,N_11549,N_11540);
and U11734 (N_11734,N_11578,N_11527);
nor U11735 (N_11735,N_11574,N_11509);
nand U11736 (N_11736,N_11589,N_11530);
nor U11737 (N_11737,N_11615,N_11608);
and U11738 (N_11738,N_11540,N_11501);
and U11739 (N_11739,N_11594,N_11542);
and U11740 (N_11740,N_11571,N_11506);
nor U11741 (N_11741,N_11514,N_11528);
nor U11742 (N_11742,N_11568,N_11540);
nor U11743 (N_11743,N_11554,N_11536);
xor U11744 (N_11744,N_11568,N_11590);
and U11745 (N_11745,N_11531,N_11514);
nor U11746 (N_11746,N_11548,N_11600);
or U11747 (N_11747,N_11565,N_11556);
nand U11748 (N_11748,N_11605,N_11555);
xor U11749 (N_11749,N_11538,N_11604);
xnor U11750 (N_11750,N_11729,N_11712);
nand U11751 (N_11751,N_11746,N_11747);
xnor U11752 (N_11752,N_11690,N_11658);
and U11753 (N_11753,N_11656,N_11680);
nor U11754 (N_11754,N_11643,N_11650);
nor U11755 (N_11755,N_11679,N_11719);
nor U11756 (N_11756,N_11738,N_11670);
and U11757 (N_11757,N_11718,N_11691);
or U11758 (N_11758,N_11635,N_11708);
nand U11759 (N_11759,N_11742,N_11701);
and U11760 (N_11760,N_11674,N_11709);
nand U11761 (N_11761,N_11706,N_11702);
or U11762 (N_11762,N_11672,N_11734);
and U11763 (N_11763,N_11713,N_11721);
nor U11764 (N_11764,N_11653,N_11654);
nand U11765 (N_11765,N_11710,N_11657);
or U11766 (N_11766,N_11722,N_11740);
and U11767 (N_11767,N_11660,N_11749);
and U11768 (N_11768,N_11639,N_11678);
nor U11769 (N_11769,N_11732,N_11724);
nand U11770 (N_11770,N_11663,N_11673);
nand U11771 (N_11771,N_11677,N_11666);
and U11772 (N_11772,N_11667,N_11627);
nand U11773 (N_11773,N_11685,N_11700);
nor U11774 (N_11774,N_11693,N_11739);
and U11775 (N_11775,N_11748,N_11726);
xor U11776 (N_11776,N_11687,N_11717);
xnor U11777 (N_11777,N_11647,N_11651);
and U11778 (N_11778,N_11634,N_11629);
or U11779 (N_11779,N_11645,N_11697);
xnor U11780 (N_11780,N_11707,N_11630);
nor U11781 (N_11781,N_11731,N_11744);
nand U11782 (N_11782,N_11728,N_11641);
xnor U11783 (N_11783,N_11684,N_11699);
xor U11784 (N_11784,N_11704,N_11652);
or U11785 (N_11785,N_11671,N_11665);
and U11786 (N_11786,N_11703,N_11727);
or U11787 (N_11787,N_11625,N_11648);
nand U11788 (N_11788,N_11694,N_11633);
and U11789 (N_11789,N_11733,N_11675);
and U11790 (N_11790,N_11730,N_11705);
nand U11791 (N_11791,N_11725,N_11716);
xor U11792 (N_11792,N_11638,N_11655);
and U11793 (N_11793,N_11682,N_11668);
xor U11794 (N_11794,N_11720,N_11695);
nand U11795 (N_11795,N_11737,N_11689);
nand U11796 (N_11796,N_11676,N_11715);
and U11797 (N_11797,N_11646,N_11714);
nor U11798 (N_11798,N_11735,N_11669);
nand U11799 (N_11799,N_11696,N_11664);
nand U11800 (N_11800,N_11659,N_11692);
xor U11801 (N_11801,N_11745,N_11631);
or U11802 (N_11802,N_11736,N_11681);
nor U11803 (N_11803,N_11644,N_11743);
nor U11804 (N_11804,N_11642,N_11626);
or U11805 (N_11805,N_11686,N_11628);
xor U11806 (N_11806,N_11632,N_11698);
nor U11807 (N_11807,N_11640,N_11741);
xnor U11808 (N_11808,N_11688,N_11711);
or U11809 (N_11809,N_11637,N_11661);
or U11810 (N_11810,N_11723,N_11662);
nor U11811 (N_11811,N_11636,N_11649);
nor U11812 (N_11812,N_11683,N_11721);
nor U11813 (N_11813,N_11651,N_11627);
nand U11814 (N_11814,N_11706,N_11640);
or U11815 (N_11815,N_11727,N_11630);
xnor U11816 (N_11816,N_11679,N_11682);
xor U11817 (N_11817,N_11669,N_11729);
or U11818 (N_11818,N_11705,N_11703);
or U11819 (N_11819,N_11654,N_11666);
nand U11820 (N_11820,N_11727,N_11645);
nor U11821 (N_11821,N_11695,N_11696);
and U11822 (N_11822,N_11631,N_11736);
xor U11823 (N_11823,N_11674,N_11634);
nand U11824 (N_11824,N_11685,N_11688);
nor U11825 (N_11825,N_11692,N_11669);
nor U11826 (N_11826,N_11683,N_11667);
xor U11827 (N_11827,N_11645,N_11637);
xnor U11828 (N_11828,N_11748,N_11696);
xor U11829 (N_11829,N_11655,N_11748);
or U11830 (N_11830,N_11679,N_11717);
nand U11831 (N_11831,N_11738,N_11642);
and U11832 (N_11832,N_11743,N_11681);
nand U11833 (N_11833,N_11743,N_11669);
or U11834 (N_11834,N_11676,N_11654);
xor U11835 (N_11835,N_11647,N_11682);
or U11836 (N_11836,N_11643,N_11690);
and U11837 (N_11837,N_11635,N_11749);
xnor U11838 (N_11838,N_11666,N_11683);
nand U11839 (N_11839,N_11669,N_11660);
or U11840 (N_11840,N_11688,N_11700);
nor U11841 (N_11841,N_11682,N_11654);
nor U11842 (N_11842,N_11685,N_11721);
or U11843 (N_11843,N_11745,N_11647);
or U11844 (N_11844,N_11717,N_11739);
or U11845 (N_11845,N_11728,N_11724);
nor U11846 (N_11846,N_11689,N_11704);
nand U11847 (N_11847,N_11634,N_11657);
xor U11848 (N_11848,N_11674,N_11647);
nor U11849 (N_11849,N_11671,N_11702);
nor U11850 (N_11850,N_11644,N_11691);
nor U11851 (N_11851,N_11644,N_11748);
xor U11852 (N_11852,N_11686,N_11678);
or U11853 (N_11853,N_11630,N_11717);
and U11854 (N_11854,N_11700,N_11632);
and U11855 (N_11855,N_11649,N_11664);
xor U11856 (N_11856,N_11636,N_11746);
xor U11857 (N_11857,N_11719,N_11654);
nor U11858 (N_11858,N_11683,N_11685);
xor U11859 (N_11859,N_11714,N_11730);
nand U11860 (N_11860,N_11710,N_11697);
nor U11861 (N_11861,N_11644,N_11637);
nor U11862 (N_11862,N_11706,N_11726);
and U11863 (N_11863,N_11666,N_11625);
xnor U11864 (N_11864,N_11700,N_11650);
and U11865 (N_11865,N_11681,N_11749);
xnor U11866 (N_11866,N_11641,N_11637);
nor U11867 (N_11867,N_11648,N_11703);
xnor U11868 (N_11868,N_11655,N_11648);
and U11869 (N_11869,N_11705,N_11740);
or U11870 (N_11870,N_11657,N_11685);
and U11871 (N_11871,N_11690,N_11662);
xnor U11872 (N_11872,N_11629,N_11628);
nand U11873 (N_11873,N_11632,N_11646);
and U11874 (N_11874,N_11709,N_11717);
nor U11875 (N_11875,N_11856,N_11752);
nand U11876 (N_11876,N_11789,N_11842);
nor U11877 (N_11877,N_11860,N_11810);
nor U11878 (N_11878,N_11769,N_11869);
nand U11879 (N_11879,N_11773,N_11803);
xor U11880 (N_11880,N_11854,N_11799);
and U11881 (N_11881,N_11852,N_11781);
and U11882 (N_11882,N_11758,N_11825);
nand U11883 (N_11883,N_11840,N_11820);
nand U11884 (N_11884,N_11816,N_11753);
and U11885 (N_11885,N_11826,N_11843);
nor U11886 (N_11886,N_11839,N_11834);
nand U11887 (N_11887,N_11791,N_11829);
or U11888 (N_11888,N_11750,N_11755);
xor U11889 (N_11889,N_11859,N_11778);
nor U11890 (N_11890,N_11832,N_11867);
or U11891 (N_11891,N_11831,N_11845);
xor U11892 (N_11892,N_11756,N_11836);
nor U11893 (N_11893,N_11811,N_11817);
xnor U11894 (N_11894,N_11823,N_11827);
and U11895 (N_11895,N_11783,N_11777);
nor U11896 (N_11896,N_11762,N_11807);
or U11897 (N_11897,N_11848,N_11855);
nor U11898 (N_11898,N_11800,N_11768);
nor U11899 (N_11899,N_11779,N_11873);
nor U11900 (N_11900,N_11857,N_11851);
and U11901 (N_11901,N_11770,N_11797);
nor U11902 (N_11902,N_11794,N_11819);
or U11903 (N_11903,N_11761,N_11864);
nand U11904 (N_11904,N_11862,N_11815);
xnor U11905 (N_11905,N_11786,N_11784);
xnor U11906 (N_11906,N_11837,N_11798);
xor U11907 (N_11907,N_11813,N_11765);
nand U11908 (N_11908,N_11796,N_11835);
or U11909 (N_11909,N_11841,N_11838);
nor U11910 (N_11910,N_11874,N_11866);
xnor U11911 (N_11911,N_11805,N_11788);
nor U11912 (N_11912,N_11792,N_11846);
nor U11913 (N_11913,N_11871,N_11847);
xnor U11914 (N_11914,N_11833,N_11812);
nand U11915 (N_11915,N_11772,N_11766);
or U11916 (N_11916,N_11849,N_11780);
or U11917 (N_11917,N_11775,N_11763);
or U11918 (N_11918,N_11821,N_11764);
and U11919 (N_11919,N_11759,N_11787);
nor U11920 (N_11920,N_11801,N_11850);
nor U11921 (N_11921,N_11861,N_11865);
or U11922 (N_11922,N_11870,N_11830);
or U11923 (N_11923,N_11793,N_11771);
xnor U11924 (N_11924,N_11853,N_11790);
xnor U11925 (N_11925,N_11804,N_11776);
nor U11926 (N_11926,N_11808,N_11760);
xor U11927 (N_11927,N_11863,N_11802);
nor U11928 (N_11928,N_11814,N_11818);
nor U11929 (N_11929,N_11809,N_11767);
xnor U11930 (N_11930,N_11858,N_11824);
xnor U11931 (N_11931,N_11751,N_11774);
xnor U11932 (N_11932,N_11868,N_11828);
and U11933 (N_11933,N_11795,N_11844);
nand U11934 (N_11934,N_11757,N_11782);
and U11935 (N_11935,N_11806,N_11754);
or U11936 (N_11936,N_11822,N_11785);
and U11937 (N_11937,N_11872,N_11799);
xnor U11938 (N_11938,N_11866,N_11841);
and U11939 (N_11939,N_11789,N_11775);
or U11940 (N_11940,N_11788,N_11776);
nand U11941 (N_11941,N_11756,N_11779);
or U11942 (N_11942,N_11846,N_11800);
nand U11943 (N_11943,N_11778,N_11800);
or U11944 (N_11944,N_11822,N_11754);
nand U11945 (N_11945,N_11762,N_11776);
nand U11946 (N_11946,N_11852,N_11838);
nand U11947 (N_11947,N_11826,N_11785);
xor U11948 (N_11948,N_11846,N_11757);
nand U11949 (N_11949,N_11815,N_11799);
nand U11950 (N_11950,N_11779,N_11831);
and U11951 (N_11951,N_11759,N_11795);
nor U11952 (N_11952,N_11808,N_11856);
nand U11953 (N_11953,N_11820,N_11854);
and U11954 (N_11954,N_11873,N_11802);
xor U11955 (N_11955,N_11798,N_11846);
nor U11956 (N_11956,N_11871,N_11806);
xor U11957 (N_11957,N_11849,N_11832);
nand U11958 (N_11958,N_11802,N_11783);
xnor U11959 (N_11959,N_11757,N_11796);
xnor U11960 (N_11960,N_11852,N_11844);
and U11961 (N_11961,N_11850,N_11797);
nand U11962 (N_11962,N_11786,N_11751);
nand U11963 (N_11963,N_11757,N_11794);
xnor U11964 (N_11964,N_11853,N_11776);
xnor U11965 (N_11965,N_11869,N_11861);
nand U11966 (N_11966,N_11791,N_11830);
or U11967 (N_11967,N_11842,N_11874);
nand U11968 (N_11968,N_11870,N_11798);
nand U11969 (N_11969,N_11810,N_11812);
xor U11970 (N_11970,N_11752,N_11750);
and U11971 (N_11971,N_11826,N_11817);
and U11972 (N_11972,N_11797,N_11827);
nand U11973 (N_11973,N_11811,N_11777);
nand U11974 (N_11974,N_11823,N_11844);
nand U11975 (N_11975,N_11777,N_11850);
and U11976 (N_11976,N_11766,N_11818);
xnor U11977 (N_11977,N_11813,N_11817);
nor U11978 (N_11978,N_11761,N_11862);
nor U11979 (N_11979,N_11854,N_11863);
and U11980 (N_11980,N_11828,N_11800);
nor U11981 (N_11981,N_11776,N_11838);
and U11982 (N_11982,N_11751,N_11780);
xnor U11983 (N_11983,N_11848,N_11754);
xor U11984 (N_11984,N_11841,N_11861);
nor U11985 (N_11985,N_11826,N_11855);
and U11986 (N_11986,N_11850,N_11772);
xnor U11987 (N_11987,N_11771,N_11751);
or U11988 (N_11988,N_11813,N_11834);
or U11989 (N_11989,N_11770,N_11822);
or U11990 (N_11990,N_11867,N_11853);
nand U11991 (N_11991,N_11847,N_11808);
or U11992 (N_11992,N_11832,N_11873);
nor U11993 (N_11993,N_11759,N_11821);
nand U11994 (N_11994,N_11774,N_11772);
xor U11995 (N_11995,N_11865,N_11868);
or U11996 (N_11996,N_11861,N_11807);
and U11997 (N_11997,N_11757,N_11835);
nor U11998 (N_11998,N_11782,N_11779);
or U11999 (N_11999,N_11763,N_11819);
and U12000 (N_12000,N_11932,N_11888);
or U12001 (N_12001,N_11875,N_11984);
and U12002 (N_12002,N_11972,N_11930);
nor U12003 (N_12003,N_11985,N_11977);
nor U12004 (N_12004,N_11904,N_11881);
or U12005 (N_12005,N_11942,N_11966);
xor U12006 (N_12006,N_11902,N_11919);
or U12007 (N_12007,N_11974,N_11961);
or U12008 (N_12008,N_11951,N_11983);
xor U12009 (N_12009,N_11973,N_11933);
nor U12010 (N_12010,N_11915,N_11990);
xnor U12011 (N_12011,N_11978,N_11912);
nand U12012 (N_12012,N_11994,N_11906);
nor U12013 (N_12013,N_11939,N_11878);
nor U12014 (N_12014,N_11903,N_11914);
nand U12015 (N_12015,N_11900,N_11889);
or U12016 (N_12016,N_11975,N_11876);
nand U12017 (N_12017,N_11964,N_11879);
and U12018 (N_12018,N_11954,N_11884);
or U12019 (N_12019,N_11922,N_11894);
xor U12020 (N_12020,N_11963,N_11950);
or U12021 (N_12021,N_11946,N_11941);
nand U12022 (N_12022,N_11993,N_11913);
nor U12023 (N_12023,N_11956,N_11907);
or U12024 (N_12024,N_11926,N_11971);
or U12025 (N_12025,N_11901,N_11885);
xnor U12026 (N_12026,N_11976,N_11988);
nand U12027 (N_12027,N_11991,N_11945);
nand U12028 (N_12028,N_11938,N_11899);
nor U12029 (N_12029,N_11920,N_11935);
or U12030 (N_12030,N_11996,N_11980);
nor U12031 (N_12031,N_11955,N_11970);
nor U12032 (N_12032,N_11949,N_11931);
and U12033 (N_12033,N_11999,N_11886);
and U12034 (N_12034,N_11998,N_11921);
nand U12035 (N_12035,N_11995,N_11986);
xnor U12036 (N_12036,N_11896,N_11962);
nand U12037 (N_12037,N_11957,N_11887);
nor U12038 (N_12038,N_11897,N_11965);
xor U12039 (N_12039,N_11987,N_11893);
xnor U12040 (N_12040,N_11936,N_11982);
xnor U12041 (N_12041,N_11960,N_11916);
nor U12042 (N_12042,N_11953,N_11937);
nand U12043 (N_12043,N_11923,N_11890);
nor U12044 (N_12044,N_11943,N_11934);
or U12045 (N_12045,N_11989,N_11877);
and U12046 (N_12046,N_11968,N_11925);
or U12047 (N_12047,N_11952,N_11898);
and U12048 (N_12048,N_11882,N_11895);
or U12049 (N_12049,N_11911,N_11958);
nand U12050 (N_12050,N_11940,N_11880);
nor U12051 (N_12051,N_11967,N_11948);
nand U12052 (N_12052,N_11979,N_11947);
xnor U12053 (N_12053,N_11908,N_11992);
and U12054 (N_12054,N_11944,N_11891);
or U12055 (N_12055,N_11883,N_11892);
nor U12056 (N_12056,N_11924,N_11969);
nand U12057 (N_12057,N_11909,N_11918);
nor U12058 (N_12058,N_11981,N_11929);
xnor U12059 (N_12059,N_11927,N_11959);
or U12060 (N_12060,N_11928,N_11997);
and U12061 (N_12061,N_11917,N_11905);
nor U12062 (N_12062,N_11910,N_11912);
xor U12063 (N_12063,N_11976,N_11949);
or U12064 (N_12064,N_11925,N_11985);
nor U12065 (N_12065,N_11939,N_11992);
nand U12066 (N_12066,N_11938,N_11990);
or U12067 (N_12067,N_11915,N_11992);
and U12068 (N_12068,N_11970,N_11969);
or U12069 (N_12069,N_11908,N_11983);
or U12070 (N_12070,N_11904,N_11985);
nor U12071 (N_12071,N_11905,N_11969);
xor U12072 (N_12072,N_11943,N_11923);
nand U12073 (N_12073,N_11895,N_11916);
nand U12074 (N_12074,N_11983,N_11986);
xnor U12075 (N_12075,N_11924,N_11883);
and U12076 (N_12076,N_11941,N_11949);
and U12077 (N_12077,N_11902,N_11951);
or U12078 (N_12078,N_11892,N_11950);
nand U12079 (N_12079,N_11994,N_11889);
nand U12080 (N_12080,N_11944,N_11931);
and U12081 (N_12081,N_11910,N_11892);
nand U12082 (N_12082,N_11973,N_11963);
nor U12083 (N_12083,N_11937,N_11990);
nor U12084 (N_12084,N_11965,N_11920);
nand U12085 (N_12085,N_11938,N_11930);
xnor U12086 (N_12086,N_11915,N_11906);
xor U12087 (N_12087,N_11987,N_11877);
xnor U12088 (N_12088,N_11893,N_11890);
nand U12089 (N_12089,N_11989,N_11887);
xor U12090 (N_12090,N_11918,N_11901);
nand U12091 (N_12091,N_11935,N_11912);
nand U12092 (N_12092,N_11884,N_11996);
nor U12093 (N_12093,N_11974,N_11995);
nor U12094 (N_12094,N_11955,N_11895);
and U12095 (N_12095,N_11916,N_11894);
nand U12096 (N_12096,N_11885,N_11896);
xnor U12097 (N_12097,N_11995,N_11944);
nand U12098 (N_12098,N_11879,N_11997);
xor U12099 (N_12099,N_11902,N_11916);
nor U12100 (N_12100,N_11962,N_11960);
nand U12101 (N_12101,N_11897,N_11976);
nand U12102 (N_12102,N_11970,N_11900);
nand U12103 (N_12103,N_11904,N_11951);
or U12104 (N_12104,N_11918,N_11936);
and U12105 (N_12105,N_11941,N_11936);
xor U12106 (N_12106,N_11927,N_11990);
and U12107 (N_12107,N_11997,N_11911);
or U12108 (N_12108,N_11921,N_11962);
nand U12109 (N_12109,N_11954,N_11935);
xnor U12110 (N_12110,N_11889,N_11961);
nand U12111 (N_12111,N_11979,N_11945);
nor U12112 (N_12112,N_11981,N_11875);
and U12113 (N_12113,N_11981,N_11987);
nand U12114 (N_12114,N_11967,N_11931);
nand U12115 (N_12115,N_11961,N_11998);
nor U12116 (N_12116,N_11885,N_11935);
or U12117 (N_12117,N_11933,N_11985);
nor U12118 (N_12118,N_11980,N_11916);
xor U12119 (N_12119,N_11966,N_11971);
xnor U12120 (N_12120,N_11961,N_11935);
or U12121 (N_12121,N_11943,N_11963);
xor U12122 (N_12122,N_11970,N_11960);
xnor U12123 (N_12123,N_11966,N_11944);
and U12124 (N_12124,N_11886,N_11989);
xor U12125 (N_12125,N_12106,N_12086);
or U12126 (N_12126,N_12032,N_12034);
nor U12127 (N_12127,N_12122,N_12039);
nand U12128 (N_12128,N_12090,N_12052);
xor U12129 (N_12129,N_12058,N_12054);
nor U12130 (N_12130,N_12010,N_12053);
and U12131 (N_12131,N_12019,N_12088);
and U12132 (N_12132,N_12091,N_12051);
nor U12133 (N_12133,N_12021,N_12023);
nand U12134 (N_12134,N_12055,N_12031);
xnor U12135 (N_12135,N_12094,N_12077);
xor U12136 (N_12136,N_12098,N_12109);
or U12137 (N_12137,N_12100,N_12089);
xor U12138 (N_12138,N_12050,N_12047);
nand U12139 (N_12139,N_12037,N_12062);
or U12140 (N_12140,N_12008,N_12120);
or U12141 (N_12141,N_12024,N_12076);
xnor U12142 (N_12142,N_12085,N_12033);
xnor U12143 (N_12143,N_12114,N_12080);
and U12144 (N_12144,N_12029,N_12009);
or U12145 (N_12145,N_12105,N_12063);
nand U12146 (N_12146,N_12061,N_12104);
xor U12147 (N_12147,N_12048,N_12038);
nand U12148 (N_12148,N_12087,N_12007);
and U12149 (N_12149,N_12017,N_12121);
nor U12150 (N_12150,N_12074,N_12118);
and U12151 (N_12151,N_12005,N_12083);
xor U12152 (N_12152,N_12107,N_12040);
xnor U12153 (N_12153,N_12079,N_12044);
and U12154 (N_12154,N_12075,N_12012);
nor U12155 (N_12155,N_12093,N_12069);
nor U12156 (N_12156,N_12045,N_12082);
or U12157 (N_12157,N_12068,N_12099);
nand U12158 (N_12158,N_12101,N_12014);
or U12159 (N_12159,N_12030,N_12064);
or U12160 (N_12160,N_12056,N_12111);
nand U12161 (N_12161,N_12041,N_12035);
nor U12162 (N_12162,N_12015,N_12066);
and U12163 (N_12163,N_12043,N_12022);
nor U12164 (N_12164,N_12020,N_12081);
or U12165 (N_12165,N_12065,N_12092);
or U12166 (N_12166,N_12000,N_12119);
nand U12167 (N_12167,N_12026,N_12003);
or U12168 (N_12168,N_12096,N_12117);
nor U12169 (N_12169,N_12078,N_12025);
xnor U12170 (N_12170,N_12060,N_12071);
and U12171 (N_12171,N_12112,N_12115);
xnor U12172 (N_12172,N_12103,N_12057);
or U12173 (N_12173,N_12004,N_12116);
nor U12174 (N_12174,N_12113,N_12095);
nand U12175 (N_12175,N_12123,N_12018);
xnor U12176 (N_12176,N_12011,N_12073);
nor U12177 (N_12177,N_12027,N_12067);
xnor U12178 (N_12178,N_12001,N_12070);
nor U12179 (N_12179,N_12072,N_12097);
nand U12180 (N_12180,N_12016,N_12036);
and U12181 (N_12181,N_12102,N_12059);
and U12182 (N_12182,N_12006,N_12084);
nand U12183 (N_12183,N_12049,N_12124);
or U12184 (N_12184,N_12110,N_12028);
nand U12185 (N_12185,N_12046,N_12042);
nor U12186 (N_12186,N_12108,N_12013);
nor U12187 (N_12187,N_12002,N_12051);
or U12188 (N_12188,N_12033,N_12002);
nand U12189 (N_12189,N_12069,N_12086);
or U12190 (N_12190,N_12120,N_12009);
xnor U12191 (N_12191,N_12098,N_12063);
xor U12192 (N_12192,N_12073,N_12077);
xnor U12193 (N_12193,N_12050,N_12048);
or U12194 (N_12194,N_12043,N_12029);
xor U12195 (N_12195,N_12076,N_12094);
nand U12196 (N_12196,N_12072,N_12101);
nor U12197 (N_12197,N_12105,N_12117);
xor U12198 (N_12198,N_12107,N_12092);
or U12199 (N_12199,N_12086,N_12013);
xor U12200 (N_12200,N_12039,N_12090);
or U12201 (N_12201,N_12078,N_12035);
or U12202 (N_12202,N_12002,N_12036);
or U12203 (N_12203,N_12004,N_12002);
and U12204 (N_12204,N_12058,N_12005);
nor U12205 (N_12205,N_12069,N_12084);
or U12206 (N_12206,N_12082,N_12115);
and U12207 (N_12207,N_12032,N_12108);
nand U12208 (N_12208,N_12030,N_12014);
xnor U12209 (N_12209,N_12010,N_12116);
nor U12210 (N_12210,N_12110,N_12119);
nor U12211 (N_12211,N_12065,N_12093);
nand U12212 (N_12212,N_12099,N_12081);
xnor U12213 (N_12213,N_12018,N_12077);
xor U12214 (N_12214,N_12036,N_12106);
xnor U12215 (N_12215,N_12058,N_12001);
xnor U12216 (N_12216,N_12023,N_12106);
or U12217 (N_12217,N_12033,N_12080);
xnor U12218 (N_12218,N_12098,N_12025);
xnor U12219 (N_12219,N_12118,N_12068);
or U12220 (N_12220,N_12001,N_12012);
nand U12221 (N_12221,N_12073,N_12123);
nor U12222 (N_12222,N_12005,N_12092);
xnor U12223 (N_12223,N_12098,N_12067);
nor U12224 (N_12224,N_12069,N_12015);
and U12225 (N_12225,N_12092,N_12074);
nand U12226 (N_12226,N_12008,N_12075);
or U12227 (N_12227,N_12124,N_12055);
nor U12228 (N_12228,N_12036,N_12079);
xor U12229 (N_12229,N_12114,N_12014);
xnor U12230 (N_12230,N_12026,N_12067);
nand U12231 (N_12231,N_12113,N_12124);
and U12232 (N_12232,N_12023,N_12096);
or U12233 (N_12233,N_12007,N_12117);
xnor U12234 (N_12234,N_12047,N_12006);
xnor U12235 (N_12235,N_12121,N_12013);
xnor U12236 (N_12236,N_12111,N_12031);
and U12237 (N_12237,N_12110,N_12062);
nor U12238 (N_12238,N_12089,N_12013);
xor U12239 (N_12239,N_12102,N_12073);
nor U12240 (N_12240,N_12028,N_12011);
nor U12241 (N_12241,N_12025,N_12083);
xnor U12242 (N_12242,N_12029,N_12036);
nand U12243 (N_12243,N_12090,N_12076);
or U12244 (N_12244,N_12124,N_12001);
or U12245 (N_12245,N_12052,N_12081);
and U12246 (N_12246,N_12065,N_12055);
nand U12247 (N_12247,N_12038,N_12079);
and U12248 (N_12248,N_12084,N_12124);
xor U12249 (N_12249,N_12070,N_12100);
or U12250 (N_12250,N_12142,N_12232);
xnor U12251 (N_12251,N_12203,N_12170);
or U12252 (N_12252,N_12133,N_12155);
nand U12253 (N_12253,N_12194,N_12176);
nor U12254 (N_12254,N_12145,N_12161);
nand U12255 (N_12255,N_12172,N_12151);
nand U12256 (N_12256,N_12178,N_12163);
nand U12257 (N_12257,N_12125,N_12204);
and U12258 (N_12258,N_12236,N_12174);
and U12259 (N_12259,N_12138,N_12200);
or U12260 (N_12260,N_12202,N_12160);
nand U12261 (N_12261,N_12215,N_12182);
xor U12262 (N_12262,N_12246,N_12201);
nor U12263 (N_12263,N_12223,N_12221);
or U12264 (N_12264,N_12220,N_12193);
or U12265 (N_12265,N_12177,N_12153);
and U12266 (N_12266,N_12234,N_12226);
nor U12267 (N_12267,N_12129,N_12211);
xnor U12268 (N_12268,N_12213,N_12179);
xor U12269 (N_12269,N_12228,N_12187);
and U12270 (N_12270,N_12217,N_12248);
xor U12271 (N_12271,N_12241,N_12141);
nand U12272 (N_12272,N_12237,N_12134);
and U12273 (N_12273,N_12249,N_12186);
or U12274 (N_12274,N_12146,N_12143);
or U12275 (N_12275,N_12185,N_12150);
nor U12276 (N_12276,N_12209,N_12227);
or U12277 (N_12277,N_12131,N_12175);
nor U12278 (N_12278,N_12162,N_12189);
nand U12279 (N_12279,N_12210,N_12166);
xor U12280 (N_12280,N_12196,N_12183);
or U12281 (N_12281,N_12197,N_12168);
and U12282 (N_12282,N_12243,N_12219);
nor U12283 (N_12283,N_12169,N_12222);
xor U12284 (N_12284,N_12191,N_12130);
and U12285 (N_12285,N_12180,N_12144);
or U12286 (N_12286,N_12136,N_12171);
or U12287 (N_12287,N_12205,N_12148);
or U12288 (N_12288,N_12154,N_12164);
nor U12289 (N_12289,N_12230,N_12233);
and U12290 (N_12290,N_12244,N_12128);
xor U12291 (N_12291,N_12152,N_12195);
xor U12292 (N_12292,N_12184,N_12192);
or U12293 (N_12293,N_12181,N_12198);
nor U12294 (N_12294,N_12127,N_12208);
and U12295 (N_12295,N_12207,N_12159);
nor U12296 (N_12296,N_12157,N_12247);
and U12297 (N_12297,N_12212,N_12167);
nor U12298 (N_12298,N_12218,N_12245);
and U12299 (N_12299,N_12231,N_12158);
nand U12300 (N_12300,N_12135,N_12229);
nor U12301 (N_12301,N_12165,N_12190);
or U12302 (N_12302,N_12188,N_12156);
nand U12303 (N_12303,N_12140,N_12137);
or U12304 (N_12304,N_12238,N_12206);
and U12305 (N_12305,N_12224,N_12216);
nand U12306 (N_12306,N_12132,N_12242);
nand U12307 (N_12307,N_12235,N_12173);
nor U12308 (N_12308,N_12126,N_12139);
nor U12309 (N_12309,N_12199,N_12239);
and U12310 (N_12310,N_12240,N_12225);
xor U12311 (N_12311,N_12149,N_12214);
xnor U12312 (N_12312,N_12147,N_12161);
and U12313 (N_12313,N_12207,N_12216);
or U12314 (N_12314,N_12228,N_12208);
nor U12315 (N_12315,N_12213,N_12191);
or U12316 (N_12316,N_12132,N_12136);
xnor U12317 (N_12317,N_12133,N_12129);
nor U12318 (N_12318,N_12142,N_12176);
and U12319 (N_12319,N_12168,N_12212);
nor U12320 (N_12320,N_12136,N_12142);
and U12321 (N_12321,N_12198,N_12224);
and U12322 (N_12322,N_12200,N_12189);
nand U12323 (N_12323,N_12215,N_12197);
and U12324 (N_12324,N_12193,N_12235);
and U12325 (N_12325,N_12145,N_12178);
nor U12326 (N_12326,N_12167,N_12156);
or U12327 (N_12327,N_12163,N_12148);
xnor U12328 (N_12328,N_12176,N_12242);
or U12329 (N_12329,N_12241,N_12235);
or U12330 (N_12330,N_12242,N_12146);
and U12331 (N_12331,N_12153,N_12212);
and U12332 (N_12332,N_12140,N_12164);
nand U12333 (N_12333,N_12245,N_12191);
nand U12334 (N_12334,N_12169,N_12239);
nand U12335 (N_12335,N_12144,N_12237);
or U12336 (N_12336,N_12184,N_12164);
or U12337 (N_12337,N_12172,N_12204);
xnor U12338 (N_12338,N_12239,N_12173);
or U12339 (N_12339,N_12231,N_12170);
or U12340 (N_12340,N_12237,N_12177);
or U12341 (N_12341,N_12195,N_12245);
and U12342 (N_12342,N_12164,N_12131);
or U12343 (N_12343,N_12162,N_12138);
nor U12344 (N_12344,N_12228,N_12146);
xor U12345 (N_12345,N_12133,N_12191);
or U12346 (N_12346,N_12171,N_12130);
or U12347 (N_12347,N_12138,N_12186);
and U12348 (N_12348,N_12169,N_12148);
nand U12349 (N_12349,N_12170,N_12227);
xor U12350 (N_12350,N_12196,N_12228);
nor U12351 (N_12351,N_12165,N_12194);
or U12352 (N_12352,N_12238,N_12212);
nand U12353 (N_12353,N_12216,N_12213);
nor U12354 (N_12354,N_12232,N_12195);
nand U12355 (N_12355,N_12194,N_12191);
nand U12356 (N_12356,N_12125,N_12181);
xnor U12357 (N_12357,N_12133,N_12147);
nor U12358 (N_12358,N_12170,N_12169);
xnor U12359 (N_12359,N_12227,N_12167);
or U12360 (N_12360,N_12155,N_12224);
nand U12361 (N_12361,N_12230,N_12142);
and U12362 (N_12362,N_12155,N_12163);
or U12363 (N_12363,N_12174,N_12135);
nand U12364 (N_12364,N_12125,N_12238);
and U12365 (N_12365,N_12185,N_12183);
xor U12366 (N_12366,N_12154,N_12161);
and U12367 (N_12367,N_12221,N_12231);
nor U12368 (N_12368,N_12219,N_12237);
xnor U12369 (N_12369,N_12138,N_12209);
xnor U12370 (N_12370,N_12147,N_12178);
and U12371 (N_12371,N_12140,N_12178);
and U12372 (N_12372,N_12182,N_12209);
xor U12373 (N_12373,N_12160,N_12198);
and U12374 (N_12374,N_12148,N_12189);
xnor U12375 (N_12375,N_12368,N_12324);
xor U12376 (N_12376,N_12319,N_12258);
or U12377 (N_12377,N_12332,N_12348);
nand U12378 (N_12378,N_12299,N_12265);
and U12379 (N_12379,N_12291,N_12325);
and U12380 (N_12380,N_12252,N_12356);
nor U12381 (N_12381,N_12371,N_12351);
xor U12382 (N_12382,N_12301,N_12269);
or U12383 (N_12383,N_12267,N_12262);
or U12384 (N_12384,N_12313,N_12253);
nand U12385 (N_12385,N_12310,N_12336);
or U12386 (N_12386,N_12339,N_12345);
and U12387 (N_12387,N_12302,N_12349);
and U12388 (N_12388,N_12327,N_12353);
xnor U12389 (N_12389,N_12273,N_12285);
or U12390 (N_12390,N_12329,N_12333);
xor U12391 (N_12391,N_12350,N_12365);
or U12392 (N_12392,N_12303,N_12320);
or U12393 (N_12393,N_12309,N_12362);
nor U12394 (N_12394,N_12268,N_12366);
and U12395 (N_12395,N_12283,N_12275);
xor U12396 (N_12396,N_12359,N_12335);
and U12397 (N_12397,N_12355,N_12314);
xnor U12398 (N_12398,N_12292,N_12360);
xnor U12399 (N_12399,N_12343,N_12297);
xnor U12400 (N_12400,N_12300,N_12305);
xor U12401 (N_12401,N_12276,N_12316);
nand U12402 (N_12402,N_12271,N_12255);
nand U12403 (N_12403,N_12260,N_12337);
or U12404 (N_12404,N_12318,N_12294);
and U12405 (N_12405,N_12295,N_12270);
and U12406 (N_12406,N_12308,N_12341);
nand U12407 (N_12407,N_12298,N_12278);
nor U12408 (N_12408,N_12330,N_12373);
nand U12409 (N_12409,N_12334,N_12372);
and U12410 (N_12410,N_12340,N_12363);
or U12411 (N_12411,N_12274,N_12287);
and U12412 (N_12412,N_12374,N_12256);
or U12413 (N_12413,N_12281,N_12364);
xor U12414 (N_12414,N_12370,N_12306);
and U12415 (N_12415,N_12272,N_12338);
xor U12416 (N_12416,N_12311,N_12293);
nor U12417 (N_12417,N_12344,N_12257);
or U12418 (N_12418,N_12367,N_12361);
and U12419 (N_12419,N_12259,N_12326);
xor U12420 (N_12420,N_12307,N_12331);
xor U12421 (N_12421,N_12357,N_12254);
nand U12422 (N_12422,N_12277,N_12261);
nand U12423 (N_12423,N_12288,N_12250);
and U12424 (N_12424,N_12289,N_12251);
or U12425 (N_12425,N_12264,N_12312);
and U12426 (N_12426,N_12263,N_12347);
and U12427 (N_12427,N_12266,N_12280);
xnor U12428 (N_12428,N_12279,N_12342);
nand U12429 (N_12429,N_12354,N_12358);
or U12430 (N_12430,N_12282,N_12322);
xnor U12431 (N_12431,N_12321,N_12290);
nor U12432 (N_12432,N_12315,N_12296);
nand U12433 (N_12433,N_12352,N_12369);
or U12434 (N_12434,N_12346,N_12304);
nand U12435 (N_12435,N_12323,N_12317);
xor U12436 (N_12436,N_12284,N_12286);
and U12437 (N_12437,N_12328,N_12306);
or U12438 (N_12438,N_12289,N_12308);
or U12439 (N_12439,N_12326,N_12371);
and U12440 (N_12440,N_12280,N_12291);
xor U12441 (N_12441,N_12374,N_12337);
nand U12442 (N_12442,N_12292,N_12294);
or U12443 (N_12443,N_12282,N_12308);
and U12444 (N_12444,N_12304,N_12292);
nand U12445 (N_12445,N_12374,N_12371);
or U12446 (N_12446,N_12305,N_12268);
xor U12447 (N_12447,N_12298,N_12253);
and U12448 (N_12448,N_12272,N_12276);
xnor U12449 (N_12449,N_12257,N_12334);
and U12450 (N_12450,N_12301,N_12267);
or U12451 (N_12451,N_12309,N_12299);
nor U12452 (N_12452,N_12328,N_12308);
xor U12453 (N_12453,N_12324,N_12257);
and U12454 (N_12454,N_12286,N_12273);
nor U12455 (N_12455,N_12365,N_12348);
and U12456 (N_12456,N_12300,N_12264);
or U12457 (N_12457,N_12327,N_12334);
or U12458 (N_12458,N_12317,N_12335);
or U12459 (N_12459,N_12297,N_12341);
and U12460 (N_12460,N_12337,N_12290);
nand U12461 (N_12461,N_12263,N_12374);
xnor U12462 (N_12462,N_12275,N_12292);
and U12463 (N_12463,N_12323,N_12371);
nand U12464 (N_12464,N_12319,N_12348);
and U12465 (N_12465,N_12299,N_12310);
or U12466 (N_12466,N_12372,N_12331);
nor U12467 (N_12467,N_12270,N_12335);
xor U12468 (N_12468,N_12262,N_12253);
nor U12469 (N_12469,N_12285,N_12365);
and U12470 (N_12470,N_12354,N_12336);
and U12471 (N_12471,N_12351,N_12347);
and U12472 (N_12472,N_12285,N_12334);
or U12473 (N_12473,N_12312,N_12344);
xor U12474 (N_12474,N_12312,N_12351);
or U12475 (N_12475,N_12261,N_12255);
or U12476 (N_12476,N_12321,N_12306);
nand U12477 (N_12477,N_12279,N_12269);
nand U12478 (N_12478,N_12250,N_12338);
nand U12479 (N_12479,N_12257,N_12311);
nor U12480 (N_12480,N_12269,N_12259);
xor U12481 (N_12481,N_12299,N_12296);
nand U12482 (N_12482,N_12367,N_12335);
xnor U12483 (N_12483,N_12323,N_12337);
xor U12484 (N_12484,N_12257,N_12327);
and U12485 (N_12485,N_12266,N_12283);
nor U12486 (N_12486,N_12278,N_12266);
nor U12487 (N_12487,N_12276,N_12310);
and U12488 (N_12488,N_12283,N_12291);
nor U12489 (N_12489,N_12336,N_12321);
nand U12490 (N_12490,N_12320,N_12312);
and U12491 (N_12491,N_12296,N_12302);
xor U12492 (N_12492,N_12347,N_12255);
and U12493 (N_12493,N_12298,N_12283);
and U12494 (N_12494,N_12287,N_12282);
xor U12495 (N_12495,N_12300,N_12314);
nor U12496 (N_12496,N_12305,N_12274);
and U12497 (N_12497,N_12326,N_12335);
and U12498 (N_12498,N_12315,N_12353);
or U12499 (N_12499,N_12275,N_12314);
or U12500 (N_12500,N_12411,N_12427);
and U12501 (N_12501,N_12489,N_12413);
nor U12502 (N_12502,N_12483,N_12438);
or U12503 (N_12503,N_12404,N_12454);
nand U12504 (N_12504,N_12379,N_12458);
nand U12505 (N_12505,N_12398,N_12402);
or U12506 (N_12506,N_12385,N_12416);
and U12507 (N_12507,N_12464,N_12428);
and U12508 (N_12508,N_12487,N_12447);
nand U12509 (N_12509,N_12461,N_12440);
or U12510 (N_12510,N_12459,N_12455);
xnor U12511 (N_12511,N_12495,N_12472);
nand U12512 (N_12512,N_12441,N_12377);
xor U12513 (N_12513,N_12493,N_12457);
and U12514 (N_12514,N_12467,N_12431);
xnor U12515 (N_12515,N_12499,N_12397);
xnor U12516 (N_12516,N_12442,N_12400);
nor U12517 (N_12517,N_12452,N_12490);
nor U12518 (N_12518,N_12393,N_12463);
nand U12519 (N_12519,N_12387,N_12430);
nor U12520 (N_12520,N_12450,N_12421);
and U12521 (N_12521,N_12412,N_12474);
and U12522 (N_12522,N_12380,N_12475);
or U12523 (N_12523,N_12434,N_12414);
and U12524 (N_12524,N_12382,N_12408);
nand U12525 (N_12525,N_12381,N_12498);
nand U12526 (N_12526,N_12435,N_12436);
and U12527 (N_12527,N_12392,N_12423);
or U12528 (N_12528,N_12494,N_12433);
and U12529 (N_12529,N_12496,N_12448);
nor U12530 (N_12530,N_12478,N_12406);
and U12531 (N_12531,N_12468,N_12471);
xnor U12532 (N_12532,N_12469,N_12426);
or U12533 (N_12533,N_12476,N_12444);
nand U12534 (N_12534,N_12486,N_12481);
xor U12535 (N_12535,N_12432,N_12465);
nand U12536 (N_12536,N_12482,N_12429);
nand U12537 (N_12537,N_12375,N_12451);
nor U12538 (N_12538,N_12424,N_12384);
nand U12539 (N_12539,N_12445,N_12399);
or U12540 (N_12540,N_12492,N_12466);
xor U12541 (N_12541,N_12401,N_12394);
and U12542 (N_12542,N_12409,N_12391);
nand U12543 (N_12543,N_12491,N_12419);
nor U12544 (N_12544,N_12439,N_12376);
or U12545 (N_12545,N_12415,N_12456);
nand U12546 (N_12546,N_12437,N_12383);
or U12547 (N_12547,N_12396,N_12390);
xnor U12548 (N_12548,N_12417,N_12420);
nor U12549 (N_12549,N_12462,N_12388);
or U12550 (N_12550,N_12422,N_12395);
nor U12551 (N_12551,N_12403,N_12449);
or U12552 (N_12552,N_12453,N_12378);
and U12553 (N_12553,N_12480,N_12410);
nor U12554 (N_12554,N_12479,N_12446);
nor U12555 (N_12555,N_12484,N_12477);
and U12556 (N_12556,N_12407,N_12389);
or U12557 (N_12557,N_12425,N_12386);
or U12558 (N_12558,N_12443,N_12485);
xor U12559 (N_12559,N_12488,N_12460);
xnor U12560 (N_12560,N_12405,N_12470);
or U12561 (N_12561,N_12418,N_12497);
nand U12562 (N_12562,N_12473,N_12411);
and U12563 (N_12563,N_12403,N_12480);
and U12564 (N_12564,N_12415,N_12384);
nand U12565 (N_12565,N_12468,N_12407);
nor U12566 (N_12566,N_12482,N_12381);
and U12567 (N_12567,N_12472,N_12377);
nor U12568 (N_12568,N_12402,N_12444);
nor U12569 (N_12569,N_12444,N_12397);
xor U12570 (N_12570,N_12416,N_12454);
nand U12571 (N_12571,N_12406,N_12392);
and U12572 (N_12572,N_12498,N_12427);
or U12573 (N_12573,N_12472,N_12455);
and U12574 (N_12574,N_12431,N_12385);
nor U12575 (N_12575,N_12465,N_12460);
or U12576 (N_12576,N_12486,N_12496);
and U12577 (N_12577,N_12427,N_12437);
nor U12578 (N_12578,N_12383,N_12449);
nor U12579 (N_12579,N_12398,N_12381);
nand U12580 (N_12580,N_12452,N_12415);
and U12581 (N_12581,N_12446,N_12498);
xor U12582 (N_12582,N_12442,N_12445);
nor U12583 (N_12583,N_12467,N_12468);
xor U12584 (N_12584,N_12436,N_12470);
nor U12585 (N_12585,N_12463,N_12385);
xor U12586 (N_12586,N_12447,N_12377);
and U12587 (N_12587,N_12412,N_12438);
nand U12588 (N_12588,N_12401,N_12476);
or U12589 (N_12589,N_12397,N_12450);
or U12590 (N_12590,N_12389,N_12464);
or U12591 (N_12591,N_12445,N_12446);
and U12592 (N_12592,N_12451,N_12455);
nor U12593 (N_12593,N_12448,N_12386);
or U12594 (N_12594,N_12375,N_12402);
and U12595 (N_12595,N_12428,N_12397);
and U12596 (N_12596,N_12388,N_12475);
nor U12597 (N_12597,N_12384,N_12401);
or U12598 (N_12598,N_12409,N_12444);
and U12599 (N_12599,N_12440,N_12471);
xor U12600 (N_12600,N_12380,N_12460);
and U12601 (N_12601,N_12417,N_12389);
nor U12602 (N_12602,N_12421,N_12414);
and U12603 (N_12603,N_12490,N_12448);
nor U12604 (N_12604,N_12469,N_12408);
nand U12605 (N_12605,N_12405,N_12383);
xor U12606 (N_12606,N_12463,N_12489);
xnor U12607 (N_12607,N_12461,N_12489);
nand U12608 (N_12608,N_12448,N_12455);
nor U12609 (N_12609,N_12457,N_12394);
xor U12610 (N_12610,N_12381,N_12485);
or U12611 (N_12611,N_12496,N_12418);
and U12612 (N_12612,N_12437,N_12487);
nor U12613 (N_12613,N_12470,N_12419);
xnor U12614 (N_12614,N_12477,N_12466);
xor U12615 (N_12615,N_12467,N_12479);
and U12616 (N_12616,N_12406,N_12449);
nand U12617 (N_12617,N_12419,N_12450);
nor U12618 (N_12618,N_12419,N_12402);
and U12619 (N_12619,N_12470,N_12475);
nor U12620 (N_12620,N_12409,N_12389);
xor U12621 (N_12621,N_12401,N_12380);
nor U12622 (N_12622,N_12391,N_12456);
xor U12623 (N_12623,N_12400,N_12486);
and U12624 (N_12624,N_12402,N_12389);
nor U12625 (N_12625,N_12529,N_12500);
and U12626 (N_12626,N_12592,N_12544);
xnor U12627 (N_12627,N_12528,N_12508);
nor U12628 (N_12628,N_12568,N_12538);
or U12629 (N_12629,N_12554,N_12600);
xnor U12630 (N_12630,N_12523,N_12582);
xnor U12631 (N_12631,N_12550,N_12557);
or U12632 (N_12632,N_12584,N_12506);
nand U12633 (N_12633,N_12537,N_12580);
nor U12634 (N_12634,N_12521,N_12603);
or U12635 (N_12635,N_12609,N_12572);
or U12636 (N_12636,N_12533,N_12560);
or U12637 (N_12637,N_12549,N_12514);
or U12638 (N_12638,N_12610,N_12535);
xor U12639 (N_12639,N_12594,N_12519);
xnor U12640 (N_12640,N_12595,N_12589);
nand U12641 (N_12641,N_12565,N_12545);
nand U12642 (N_12642,N_12616,N_12512);
or U12643 (N_12643,N_12558,N_12507);
nor U12644 (N_12644,N_12524,N_12505);
nor U12645 (N_12645,N_12574,N_12534);
xor U12646 (N_12646,N_12599,N_12543);
and U12647 (N_12647,N_12611,N_12620);
nand U12648 (N_12648,N_12598,N_12597);
or U12649 (N_12649,N_12564,N_12502);
nand U12650 (N_12650,N_12617,N_12612);
and U12651 (N_12651,N_12619,N_12581);
nor U12652 (N_12652,N_12590,N_12552);
nor U12653 (N_12653,N_12511,N_12621);
xnor U12654 (N_12654,N_12587,N_12532);
nand U12655 (N_12655,N_12530,N_12566);
nor U12656 (N_12656,N_12536,N_12539);
xor U12657 (N_12657,N_12571,N_12542);
or U12658 (N_12658,N_12583,N_12623);
xor U12659 (N_12659,N_12525,N_12596);
nor U12660 (N_12660,N_12562,N_12622);
and U12661 (N_12661,N_12591,N_12522);
xnor U12662 (N_12662,N_12615,N_12608);
xnor U12663 (N_12663,N_12546,N_12613);
nor U12664 (N_12664,N_12567,N_12577);
or U12665 (N_12665,N_12553,N_12556);
or U12666 (N_12666,N_12516,N_12509);
nand U12667 (N_12667,N_12614,N_12559);
nor U12668 (N_12668,N_12551,N_12555);
and U12669 (N_12669,N_12540,N_12520);
or U12670 (N_12670,N_12518,N_12547);
xor U12671 (N_12671,N_12578,N_12501);
or U12672 (N_12672,N_12576,N_12573);
nor U12673 (N_12673,N_12569,N_12563);
and U12674 (N_12674,N_12515,N_12604);
or U12675 (N_12675,N_12517,N_12585);
nand U12676 (N_12676,N_12605,N_12504);
nand U12677 (N_12677,N_12588,N_12606);
and U12678 (N_12678,N_12541,N_12607);
and U12679 (N_12679,N_12624,N_12561);
and U12680 (N_12680,N_12602,N_12527);
nand U12681 (N_12681,N_12570,N_12601);
nand U12682 (N_12682,N_12531,N_12548);
or U12683 (N_12683,N_12586,N_12510);
nand U12684 (N_12684,N_12503,N_12575);
or U12685 (N_12685,N_12579,N_12526);
nor U12686 (N_12686,N_12513,N_12593);
nor U12687 (N_12687,N_12618,N_12525);
nand U12688 (N_12688,N_12619,N_12608);
and U12689 (N_12689,N_12564,N_12603);
or U12690 (N_12690,N_12520,N_12594);
or U12691 (N_12691,N_12577,N_12525);
nand U12692 (N_12692,N_12537,N_12530);
or U12693 (N_12693,N_12558,N_12575);
and U12694 (N_12694,N_12578,N_12517);
nor U12695 (N_12695,N_12515,N_12561);
nand U12696 (N_12696,N_12583,N_12575);
xor U12697 (N_12697,N_12600,N_12582);
or U12698 (N_12698,N_12619,N_12548);
or U12699 (N_12699,N_12615,N_12534);
nand U12700 (N_12700,N_12610,N_12539);
nor U12701 (N_12701,N_12522,N_12551);
nor U12702 (N_12702,N_12542,N_12585);
nand U12703 (N_12703,N_12604,N_12582);
nor U12704 (N_12704,N_12600,N_12624);
nand U12705 (N_12705,N_12556,N_12583);
nor U12706 (N_12706,N_12583,N_12563);
and U12707 (N_12707,N_12555,N_12518);
nand U12708 (N_12708,N_12506,N_12602);
xnor U12709 (N_12709,N_12582,N_12515);
nand U12710 (N_12710,N_12588,N_12508);
xor U12711 (N_12711,N_12583,N_12548);
or U12712 (N_12712,N_12610,N_12504);
or U12713 (N_12713,N_12529,N_12579);
xnor U12714 (N_12714,N_12506,N_12519);
nand U12715 (N_12715,N_12555,N_12504);
nor U12716 (N_12716,N_12541,N_12506);
nand U12717 (N_12717,N_12574,N_12535);
and U12718 (N_12718,N_12504,N_12592);
xnor U12719 (N_12719,N_12573,N_12570);
or U12720 (N_12720,N_12521,N_12531);
nand U12721 (N_12721,N_12609,N_12556);
or U12722 (N_12722,N_12534,N_12564);
or U12723 (N_12723,N_12554,N_12522);
or U12724 (N_12724,N_12536,N_12586);
and U12725 (N_12725,N_12542,N_12616);
and U12726 (N_12726,N_12613,N_12605);
nor U12727 (N_12727,N_12555,N_12531);
nor U12728 (N_12728,N_12599,N_12586);
xnor U12729 (N_12729,N_12574,N_12584);
and U12730 (N_12730,N_12574,N_12591);
and U12731 (N_12731,N_12564,N_12588);
or U12732 (N_12732,N_12606,N_12526);
and U12733 (N_12733,N_12612,N_12614);
xnor U12734 (N_12734,N_12511,N_12595);
xnor U12735 (N_12735,N_12554,N_12581);
xor U12736 (N_12736,N_12582,N_12538);
nor U12737 (N_12737,N_12529,N_12564);
nor U12738 (N_12738,N_12560,N_12624);
nand U12739 (N_12739,N_12579,N_12573);
or U12740 (N_12740,N_12568,N_12532);
xnor U12741 (N_12741,N_12555,N_12603);
or U12742 (N_12742,N_12602,N_12563);
nor U12743 (N_12743,N_12624,N_12615);
or U12744 (N_12744,N_12527,N_12599);
and U12745 (N_12745,N_12543,N_12607);
nor U12746 (N_12746,N_12615,N_12512);
xor U12747 (N_12747,N_12572,N_12551);
nor U12748 (N_12748,N_12554,N_12610);
nand U12749 (N_12749,N_12519,N_12565);
nor U12750 (N_12750,N_12654,N_12681);
and U12751 (N_12751,N_12640,N_12691);
xor U12752 (N_12752,N_12682,N_12646);
or U12753 (N_12753,N_12678,N_12718);
or U12754 (N_12754,N_12669,N_12703);
or U12755 (N_12755,N_12627,N_12714);
or U12756 (N_12756,N_12687,N_12729);
nand U12757 (N_12757,N_12720,N_12738);
or U12758 (N_12758,N_12647,N_12696);
nor U12759 (N_12759,N_12693,N_12626);
nor U12760 (N_12760,N_12657,N_12641);
or U12761 (N_12761,N_12664,N_12659);
and U12762 (N_12762,N_12661,N_12719);
xor U12763 (N_12763,N_12629,N_12734);
nand U12764 (N_12764,N_12726,N_12683);
and U12765 (N_12765,N_12711,N_12704);
nor U12766 (N_12766,N_12630,N_12744);
xor U12767 (N_12767,N_12677,N_12737);
and U12768 (N_12768,N_12648,N_12725);
xnor U12769 (N_12769,N_12670,N_12741);
and U12770 (N_12770,N_12672,N_12739);
nor U12771 (N_12771,N_12717,N_12666);
and U12772 (N_12772,N_12685,N_12644);
or U12773 (N_12773,N_12637,N_12686);
or U12774 (N_12774,N_12690,N_12735);
and U12775 (N_12775,N_12688,N_12645);
or U12776 (N_12776,N_12715,N_12695);
or U12777 (N_12777,N_12643,N_12689);
xor U12778 (N_12778,N_12697,N_12633);
xnor U12779 (N_12779,N_12702,N_12635);
nor U12780 (N_12780,N_12746,N_12736);
xor U12781 (N_12781,N_12628,N_12673);
nor U12782 (N_12782,N_12724,N_12709);
and U12783 (N_12783,N_12649,N_12692);
nor U12784 (N_12784,N_12639,N_12638);
xnor U12785 (N_12785,N_12694,N_12652);
or U12786 (N_12786,N_12684,N_12730);
or U12787 (N_12787,N_12651,N_12721);
or U12788 (N_12788,N_12634,N_12749);
or U12789 (N_12789,N_12710,N_12658);
or U12790 (N_12790,N_12728,N_12671);
and U12791 (N_12791,N_12653,N_12676);
nand U12792 (N_12792,N_12716,N_12698);
nor U12793 (N_12793,N_12631,N_12708);
nand U12794 (N_12794,N_12712,N_12701);
nor U12795 (N_12795,N_12732,N_12707);
nand U12796 (N_12796,N_12674,N_12727);
nor U12797 (N_12797,N_12745,N_12743);
or U12798 (N_12798,N_12722,N_12625);
nor U12799 (N_12799,N_12668,N_12642);
or U12800 (N_12800,N_12705,N_12665);
xnor U12801 (N_12801,N_12700,N_12632);
or U12802 (N_12802,N_12733,N_12636);
nand U12803 (N_12803,N_12663,N_12655);
nand U12804 (N_12804,N_12660,N_12656);
nor U12805 (N_12805,N_12706,N_12679);
and U12806 (N_12806,N_12731,N_12723);
or U12807 (N_12807,N_12680,N_12699);
and U12808 (N_12808,N_12675,N_12748);
nor U12809 (N_12809,N_12742,N_12747);
and U12810 (N_12810,N_12713,N_12662);
and U12811 (N_12811,N_12740,N_12650);
or U12812 (N_12812,N_12667,N_12681);
nand U12813 (N_12813,N_12692,N_12707);
or U12814 (N_12814,N_12729,N_12627);
xnor U12815 (N_12815,N_12647,N_12717);
nand U12816 (N_12816,N_12645,N_12627);
nor U12817 (N_12817,N_12703,N_12725);
nand U12818 (N_12818,N_12657,N_12730);
or U12819 (N_12819,N_12681,N_12627);
nor U12820 (N_12820,N_12667,N_12710);
and U12821 (N_12821,N_12650,N_12632);
xor U12822 (N_12822,N_12710,N_12626);
and U12823 (N_12823,N_12707,N_12711);
or U12824 (N_12824,N_12720,N_12683);
xor U12825 (N_12825,N_12715,N_12685);
nand U12826 (N_12826,N_12699,N_12677);
and U12827 (N_12827,N_12748,N_12712);
nand U12828 (N_12828,N_12740,N_12679);
nand U12829 (N_12829,N_12632,N_12729);
or U12830 (N_12830,N_12672,N_12677);
nand U12831 (N_12831,N_12726,N_12741);
and U12832 (N_12832,N_12644,N_12745);
nand U12833 (N_12833,N_12749,N_12704);
nand U12834 (N_12834,N_12731,N_12727);
nor U12835 (N_12835,N_12653,N_12687);
xnor U12836 (N_12836,N_12687,N_12627);
xnor U12837 (N_12837,N_12672,N_12727);
and U12838 (N_12838,N_12694,N_12625);
xnor U12839 (N_12839,N_12729,N_12749);
or U12840 (N_12840,N_12699,N_12670);
xor U12841 (N_12841,N_12678,N_12693);
xor U12842 (N_12842,N_12625,N_12738);
or U12843 (N_12843,N_12742,N_12707);
xnor U12844 (N_12844,N_12636,N_12719);
and U12845 (N_12845,N_12749,N_12676);
or U12846 (N_12846,N_12653,N_12713);
xnor U12847 (N_12847,N_12677,N_12730);
and U12848 (N_12848,N_12701,N_12738);
or U12849 (N_12849,N_12713,N_12629);
nor U12850 (N_12850,N_12657,N_12637);
xor U12851 (N_12851,N_12741,N_12729);
nor U12852 (N_12852,N_12711,N_12728);
or U12853 (N_12853,N_12644,N_12666);
or U12854 (N_12854,N_12690,N_12748);
or U12855 (N_12855,N_12706,N_12737);
nor U12856 (N_12856,N_12670,N_12731);
nor U12857 (N_12857,N_12626,N_12719);
and U12858 (N_12858,N_12682,N_12714);
nor U12859 (N_12859,N_12674,N_12631);
or U12860 (N_12860,N_12726,N_12686);
and U12861 (N_12861,N_12673,N_12631);
or U12862 (N_12862,N_12686,N_12665);
nor U12863 (N_12863,N_12748,N_12646);
and U12864 (N_12864,N_12628,N_12690);
and U12865 (N_12865,N_12656,N_12731);
nand U12866 (N_12866,N_12748,N_12669);
or U12867 (N_12867,N_12694,N_12726);
nand U12868 (N_12868,N_12674,N_12718);
nor U12869 (N_12869,N_12655,N_12703);
xor U12870 (N_12870,N_12704,N_12647);
xnor U12871 (N_12871,N_12675,N_12647);
xor U12872 (N_12872,N_12680,N_12638);
nand U12873 (N_12873,N_12668,N_12706);
xor U12874 (N_12874,N_12664,N_12631);
nor U12875 (N_12875,N_12781,N_12777);
nand U12876 (N_12876,N_12788,N_12758);
nor U12877 (N_12877,N_12813,N_12847);
nor U12878 (N_12878,N_12871,N_12818);
nor U12879 (N_12879,N_12807,N_12848);
and U12880 (N_12880,N_12850,N_12787);
nor U12881 (N_12881,N_12780,N_12870);
nand U12882 (N_12882,N_12829,N_12859);
and U12883 (N_12883,N_12815,N_12796);
and U12884 (N_12884,N_12861,N_12802);
and U12885 (N_12885,N_12828,N_12779);
nor U12886 (N_12886,N_12814,N_12755);
xnor U12887 (N_12887,N_12823,N_12773);
or U12888 (N_12888,N_12805,N_12864);
nor U12889 (N_12889,N_12783,N_12754);
xnor U12890 (N_12890,N_12766,N_12769);
or U12891 (N_12891,N_12792,N_12844);
nand U12892 (N_12892,N_12866,N_12800);
nor U12893 (N_12893,N_12825,N_12830);
or U12894 (N_12894,N_12851,N_12838);
xor U12895 (N_12895,N_12854,N_12837);
nand U12896 (N_12896,N_12753,N_12757);
xnor U12897 (N_12897,N_12756,N_12832);
nor U12898 (N_12898,N_12771,N_12841);
xnor U12899 (N_12899,N_12865,N_12867);
nand U12900 (N_12900,N_12797,N_12760);
nand U12901 (N_12901,N_12786,N_12853);
and U12902 (N_12902,N_12806,N_12845);
or U12903 (N_12903,N_12826,N_12811);
xnor U12904 (N_12904,N_12764,N_12862);
or U12905 (N_12905,N_12791,N_12820);
xor U12906 (N_12906,N_12824,N_12849);
nor U12907 (N_12907,N_12839,N_12819);
nor U12908 (N_12908,N_12812,N_12803);
nor U12909 (N_12909,N_12835,N_12789);
xnor U12910 (N_12910,N_12833,N_12768);
nand U12911 (N_12911,N_12782,N_12765);
and U12912 (N_12912,N_12804,N_12860);
xnor U12913 (N_12913,N_12750,N_12775);
nor U12914 (N_12914,N_12822,N_12873);
or U12915 (N_12915,N_12834,N_12763);
xor U12916 (N_12916,N_12772,N_12817);
xor U12917 (N_12917,N_12843,N_12858);
xor U12918 (N_12918,N_12816,N_12752);
or U12919 (N_12919,N_12827,N_12776);
nor U12920 (N_12920,N_12869,N_12840);
nand U12921 (N_12921,N_12799,N_12874);
nor U12922 (N_12922,N_12793,N_12842);
and U12923 (N_12923,N_12831,N_12759);
nor U12924 (N_12924,N_12836,N_12778);
and U12925 (N_12925,N_12855,N_12762);
and U12926 (N_12926,N_12794,N_12857);
or U12927 (N_12927,N_12810,N_12809);
nand U12928 (N_12928,N_12872,N_12795);
nand U12929 (N_12929,N_12846,N_12801);
xor U12930 (N_12930,N_12821,N_12761);
or U12931 (N_12931,N_12856,N_12784);
or U12932 (N_12932,N_12770,N_12863);
nor U12933 (N_12933,N_12751,N_12774);
and U12934 (N_12934,N_12808,N_12852);
and U12935 (N_12935,N_12790,N_12798);
nand U12936 (N_12936,N_12785,N_12868);
nand U12937 (N_12937,N_12767,N_12834);
xnor U12938 (N_12938,N_12788,N_12819);
nand U12939 (N_12939,N_12756,N_12783);
or U12940 (N_12940,N_12787,N_12810);
nand U12941 (N_12941,N_12820,N_12838);
nor U12942 (N_12942,N_12864,N_12758);
or U12943 (N_12943,N_12807,N_12779);
nor U12944 (N_12944,N_12762,N_12782);
and U12945 (N_12945,N_12849,N_12810);
or U12946 (N_12946,N_12808,N_12771);
nor U12947 (N_12947,N_12857,N_12810);
xnor U12948 (N_12948,N_12821,N_12784);
nand U12949 (N_12949,N_12788,N_12834);
xnor U12950 (N_12950,N_12771,N_12849);
and U12951 (N_12951,N_12862,N_12770);
xnor U12952 (N_12952,N_12821,N_12774);
or U12953 (N_12953,N_12774,N_12831);
nor U12954 (N_12954,N_12858,N_12794);
nor U12955 (N_12955,N_12796,N_12806);
and U12956 (N_12956,N_12809,N_12838);
xor U12957 (N_12957,N_12800,N_12753);
or U12958 (N_12958,N_12872,N_12874);
nor U12959 (N_12959,N_12758,N_12838);
nand U12960 (N_12960,N_12765,N_12806);
or U12961 (N_12961,N_12865,N_12776);
and U12962 (N_12962,N_12801,N_12848);
and U12963 (N_12963,N_12873,N_12823);
and U12964 (N_12964,N_12830,N_12838);
nand U12965 (N_12965,N_12773,N_12853);
or U12966 (N_12966,N_12837,N_12873);
nand U12967 (N_12967,N_12811,N_12790);
xor U12968 (N_12968,N_12774,N_12866);
nor U12969 (N_12969,N_12755,N_12781);
xor U12970 (N_12970,N_12845,N_12798);
nor U12971 (N_12971,N_12801,N_12818);
or U12972 (N_12972,N_12810,N_12788);
or U12973 (N_12973,N_12757,N_12811);
nand U12974 (N_12974,N_12828,N_12858);
or U12975 (N_12975,N_12843,N_12798);
nand U12976 (N_12976,N_12833,N_12816);
nand U12977 (N_12977,N_12840,N_12859);
or U12978 (N_12978,N_12755,N_12851);
nor U12979 (N_12979,N_12810,N_12752);
xor U12980 (N_12980,N_12812,N_12787);
or U12981 (N_12981,N_12809,N_12807);
nor U12982 (N_12982,N_12819,N_12803);
and U12983 (N_12983,N_12787,N_12765);
or U12984 (N_12984,N_12816,N_12757);
xor U12985 (N_12985,N_12854,N_12810);
nor U12986 (N_12986,N_12797,N_12809);
or U12987 (N_12987,N_12804,N_12754);
and U12988 (N_12988,N_12848,N_12760);
nor U12989 (N_12989,N_12828,N_12773);
xnor U12990 (N_12990,N_12839,N_12805);
and U12991 (N_12991,N_12832,N_12871);
and U12992 (N_12992,N_12751,N_12795);
or U12993 (N_12993,N_12756,N_12771);
or U12994 (N_12994,N_12852,N_12844);
and U12995 (N_12995,N_12798,N_12787);
and U12996 (N_12996,N_12825,N_12759);
nand U12997 (N_12997,N_12823,N_12786);
nor U12998 (N_12998,N_12765,N_12862);
nand U12999 (N_12999,N_12767,N_12763);
nor U13000 (N_13000,N_12960,N_12944);
or U13001 (N_13001,N_12909,N_12932);
and U13002 (N_13002,N_12896,N_12913);
nor U13003 (N_13003,N_12898,N_12878);
xnor U13004 (N_13004,N_12947,N_12895);
and U13005 (N_13005,N_12936,N_12900);
nand U13006 (N_13006,N_12923,N_12964);
and U13007 (N_13007,N_12925,N_12945);
xor U13008 (N_13008,N_12980,N_12994);
or U13009 (N_13009,N_12989,N_12974);
and U13010 (N_13010,N_12986,N_12907);
and U13011 (N_13011,N_12943,N_12897);
or U13012 (N_13012,N_12877,N_12984);
and U13013 (N_13013,N_12942,N_12910);
xnor U13014 (N_13014,N_12979,N_12965);
nor U13015 (N_13015,N_12961,N_12971);
nand U13016 (N_13016,N_12953,N_12977);
and U13017 (N_13017,N_12941,N_12981);
and U13018 (N_13018,N_12882,N_12915);
xnor U13019 (N_13019,N_12887,N_12999);
or U13020 (N_13020,N_12992,N_12899);
nor U13021 (N_13021,N_12995,N_12983);
or U13022 (N_13022,N_12949,N_12991);
nand U13023 (N_13023,N_12987,N_12879);
and U13024 (N_13024,N_12888,N_12937);
or U13025 (N_13025,N_12921,N_12912);
or U13026 (N_13026,N_12884,N_12889);
nand U13027 (N_13027,N_12985,N_12876);
and U13028 (N_13028,N_12920,N_12993);
or U13029 (N_13029,N_12883,N_12973);
nor U13030 (N_13030,N_12966,N_12901);
nor U13031 (N_13031,N_12934,N_12886);
nand U13032 (N_13032,N_12962,N_12922);
or U13033 (N_13033,N_12946,N_12917);
xnor U13034 (N_13034,N_12958,N_12930);
nand U13035 (N_13035,N_12951,N_12929);
nand U13036 (N_13036,N_12892,N_12890);
nor U13037 (N_13037,N_12885,N_12963);
nand U13038 (N_13038,N_12956,N_12996);
xnor U13039 (N_13039,N_12926,N_12880);
xor U13040 (N_13040,N_12911,N_12894);
and U13041 (N_13041,N_12924,N_12957);
xor U13042 (N_13042,N_12940,N_12893);
nand U13043 (N_13043,N_12968,N_12982);
and U13044 (N_13044,N_12950,N_12904);
and U13045 (N_13045,N_12997,N_12948);
nand U13046 (N_13046,N_12969,N_12970);
or U13047 (N_13047,N_12955,N_12935);
xor U13048 (N_13048,N_12954,N_12928);
xor U13049 (N_13049,N_12988,N_12967);
nand U13050 (N_13050,N_12908,N_12972);
xnor U13051 (N_13051,N_12914,N_12903);
xnor U13052 (N_13052,N_12905,N_12939);
xnor U13053 (N_13053,N_12875,N_12919);
and U13054 (N_13054,N_12978,N_12916);
xor U13055 (N_13055,N_12931,N_12938);
and U13056 (N_13056,N_12998,N_12952);
and U13057 (N_13057,N_12902,N_12933);
xor U13058 (N_13058,N_12975,N_12906);
nor U13059 (N_13059,N_12927,N_12959);
or U13060 (N_13060,N_12918,N_12990);
nand U13061 (N_13061,N_12881,N_12891);
nand U13062 (N_13062,N_12976,N_12875);
xor U13063 (N_13063,N_12928,N_12897);
or U13064 (N_13064,N_12965,N_12967);
xor U13065 (N_13065,N_12987,N_12922);
and U13066 (N_13066,N_12906,N_12995);
or U13067 (N_13067,N_12910,N_12877);
or U13068 (N_13068,N_12978,N_12953);
or U13069 (N_13069,N_12973,N_12915);
nand U13070 (N_13070,N_12979,N_12876);
nand U13071 (N_13071,N_12941,N_12974);
nand U13072 (N_13072,N_12928,N_12995);
and U13073 (N_13073,N_12920,N_12982);
and U13074 (N_13074,N_12952,N_12875);
nand U13075 (N_13075,N_12890,N_12983);
xnor U13076 (N_13076,N_12954,N_12982);
xor U13077 (N_13077,N_12964,N_12934);
or U13078 (N_13078,N_12998,N_12900);
nor U13079 (N_13079,N_12934,N_12959);
xor U13080 (N_13080,N_12943,N_12985);
and U13081 (N_13081,N_12964,N_12997);
nor U13082 (N_13082,N_12900,N_12991);
or U13083 (N_13083,N_12975,N_12925);
xor U13084 (N_13084,N_12941,N_12979);
and U13085 (N_13085,N_12896,N_12938);
and U13086 (N_13086,N_12999,N_12928);
and U13087 (N_13087,N_12892,N_12899);
nand U13088 (N_13088,N_12938,N_12995);
nand U13089 (N_13089,N_12974,N_12895);
nor U13090 (N_13090,N_12898,N_12970);
and U13091 (N_13091,N_12888,N_12914);
and U13092 (N_13092,N_12907,N_12935);
xnor U13093 (N_13093,N_12933,N_12989);
nor U13094 (N_13094,N_12973,N_12911);
nor U13095 (N_13095,N_12885,N_12914);
nor U13096 (N_13096,N_12929,N_12976);
xor U13097 (N_13097,N_12991,N_12879);
nand U13098 (N_13098,N_12926,N_12893);
and U13099 (N_13099,N_12914,N_12878);
nand U13100 (N_13100,N_12994,N_12902);
and U13101 (N_13101,N_12903,N_12904);
xor U13102 (N_13102,N_12885,N_12902);
nand U13103 (N_13103,N_12915,N_12933);
and U13104 (N_13104,N_12980,N_12899);
or U13105 (N_13105,N_12979,N_12882);
nand U13106 (N_13106,N_12959,N_12984);
and U13107 (N_13107,N_12935,N_12977);
nand U13108 (N_13108,N_12998,N_12956);
nand U13109 (N_13109,N_12958,N_12891);
or U13110 (N_13110,N_12941,N_12946);
or U13111 (N_13111,N_12901,N_12998);
nor U13112 (N_13112,N_12891,N_12924);
nand U13113 (N_13113,N_12909,N_12904);
nand U13114 (N_13114,N_12948,N_12963);
nor U13115 (N_13115,N_12929,N_12892);
or U13116 (N_13116,N_12897,N_12965);
nor U13117 (N_13117,N_12990,N_12937);
xnor U13118 (N_13118,N_12911,N_12881);
nor U13119 (N_13119,N_12952,N_12940);
and U13120 (N_13120,N_12959,N_12971);
nand U13121 (N_13121,N_12983,N_12879);
xnor U13122 (N_13122,N_12974,N_12908);
xor U13123 (N_13123,N_12912,N_12922);
xor U13124 (N_13124,N_12933,N_12892);
nand U13125 (N_13125,N_13009,N_13004);
or U13126 (N_13126,N_13005,N_13026);
xnor U13127 (N_13127,N_13069,N_13037);
or U13128 (N_13128,N_13016,N_13036);
nand U13129 (N_13129,N_13056,N_13103);
and U13130 (N_13130,N_13003,N_13055);
or U13131 (N_13131,N_13034,N_13022);
nor U13132 (N_13132,N_13031,N_13107);
or U13133 (N_13133,N_13092,N_13000);
xor U13134 (N_13134,N_13017,N_13075);
or U13135 (N_13135,N_13020,N_13077);
nand U13136 (N_13136,N_13076,N_13095);
nand U13137 (N_13137,N_13023,N_13080);
or U13138 (N_13138,N_13096,N_13014);
nor U13139 (N_13139,N_13029,N_13085);
and U13140 (N_13140,N_13047,N_13042);
and U13141 (N_13141,N_13101,N_13082);
xor U13142 (N_13142,N_13062,N_13035);
or U13143 (N_13143,N_13119,N_13050);
nor U13144 (N_13144,N_13010,N_13118);
and U13145 (N_13145,N_13028,N_13024);
nor U13146 (N_13146,N_13064,N_13065);
or U13147 (N_13147,N_13018,N_13006);
xor U13148 (N_13148,N_13110,N_13106);
and U13149 (N_13149,N_13002,N_13094);
or U13150 (N_13150,N_13079,N_13059);
nand U13151 (N_13151,N_13097,N_13112);
and U13152 (N_13152,N_13038,N_13025);
or U13153 (N_13153,N_13051,N_13066);
or U13154 (N_13154,N_13105,N_13086);
nand U13155 (N_13155,N_13120,N_13053);
and U13156 (N_13156,N_13108,N_13088);
nor U13157 (N_13157,N_13122,N_13008);
and U13158 (N_13158,N_13007,N_13114);
and U13159 (N_13159,N_13111,N_13099);
xor U13160 (N_13160,N_13091,N_13039);
xor U13161 (N_13161,N_13058,N_13070);
nor U13162 (N_13162,N_13068,N_13063);
and U13163 (N_13163,N_13057,N_13032);
or U13164 (N_13164,N_13090,N_13087);
and U13165 (N_13165,N_13044,N_13109);
nor U13166 (N_13166,N_13041,N_13123);
or U13167 (N_13167,N_13001,N_13121);
nor U13168 (N_13168,N_13046,N_13073);
and U13169 (N_13169,N_13115,N_13012);
nor U13170 (N_13170,N_13084,N_13052);
nor U13171 (N_13171,N_13043,N_13071);
nor U13172 (N_13172,N_13093,N_13124);
xor U13173 (N_13173,N_13098,N_13104);
and U13174 (N_13174,N_13072,N_13113);
nor U13175 (N_13175,N_13054,N_13048);
and U13176 (N_13176,N_13033,N_13117);
nand U13177 (N_13177,N_13011,N_13061);
nor U13178 (N_13178,N_13083,N_13067);
nor U13179 (N_13179,N_13027,N_13102);
or U13180 (N_13180,N_13045,N_13074);
and U13181 (N_13181,N_13030,N_13100);
nand U13182 (N_13182,N_13060,N_13049);
nand U13183 (N_13183,N_13013,N_13040);
xor U13184 (N_13184,N_13116,N_13089);
nand U13185 (N_13185,N_13021,N_13019);
xor U13186 (N_13186,N_13078,N_13081);
nor U13187 (N_13187,N_13015,N_13120);
nand U13188 (N_13188,N_13102,N_13116);
nor U13189 (N_13189,N_13076,N_13006);
nand U13190 (N_13190,N_13042,N_13061);
xnor U13191 (N_13191,N_13040,N_13003);
xnor U13192 (N_13192,N_13037,N_13115);
nand U13193 (N_13193,N_13033,N_13050);
nand U13194 (N_13194,N_13099,N_13071);
nor U13195 (N_13195,N_13031,N_13095);
nor U13196 (N_13196,N_13064,N_13098);
nor U13197 (N_13197,N_13057,N_13116);
and U13198 (N_13198,N_13018,N_13015);
nand U13199 (N_13199,N_13042,N_13111);
xor U13200 (N_13200,N_13030,N_13000);
nor U13201 (N_13201,N_13123,N_13059);
nand U13202 (N_13202,N_13096,N_13078);
nand U13203 (N_13203,N_13099,N_13022);
or U13204 (N_13204,N_13087,N_13120);
and U13205 (N_13205,N_13089,N_13094);
nand U13206 (N_13206,N_13101,N_13077);
nand U13207 (N_13207,N_13011,N_13103);
or U13208 (N_13208,N_13074,N_13086);
or U13209 (N_13209,N_13101,N_13123);
and U13210 (N_13210,N_13123,N_13111);
nor U13211 (N_13211,N_13015,N_13117);
nor U13212 (N_13212,N_13120,N_13078);
nor U13213 (N_13213,N_13122,N_13073);
nor U13214 (N_13214,N_13002,N_13013);
nor U13215 (N_13215,N_13075,N_13023);
or U13216 (N_13216,N_13028,N_13110);
nor U13217 (N_13217,N_13045,N_13005);
nand U13218 (N_13218,N_13051,N_13029);
and U13219 (N_13219,N_13000,N_13122);
nand U13220 (N_13220,N_13057,N_13041);
or U13221 (N_13221,N_13034,N_13033);
nand U13222 (N_13222,N_13070,N_13090);
xnor U13223 (N_13223,N_13054,N_13075);
and U13224 (N_13224,N_13042,N_13008);
and U13225 (N_13225,N_13081,N_13107);
nor U13226 (N_13226,N_13034,N_13051);
nor U13227 (N_13227,N_13108,N_13060);
and U13228 (N_13228,N_13072,N_13067);
or U13229 (N_13229,N_13016,N_13054);
and U13230 (N_13230,N_13016,N_13005);
or U13231 (N_13231,N_13034,N_13109);
nor U13232 (N_13232,N_13028,N_13074);
and U13233 (N_13233,N_13047,N_13041);
xnor U13234 (N_13234,N_13024,N_13123);
xor U13235 (N_13235,N_13051,N_13033);
and U13236 (N_13236,N_13020,N_13047);
nand U13237 (N_13237,N_13094,N_13114);
or U13238 (N_13238,N_13120,N_13011);
and U13239 (N_13239,N_13063,N_13117);
or U13240 (N_13240,N_13112,N_13105);
nor U13241 (N_13241,N_13094,N_13101);
nor U13242 (N_13242,N_13108,N_13087);
and U13243 (N_13243,N_13058,N_13013);
nor U13244 (N_13244,N_13010,N_13001);
or U13245 (N_13245,N_13024,N_13021);
or U13246 (N_13246,N_13012,N_13093);
or U13247 (N_13247,N_13000,N_13029);
and U13248 (N_13248,N_13120,N_13092);
nand U13249 (N_13249,N_13046,N_13102);
nor U13250 (N_13250,N_13249,N_13175);
or U13251 (N_13251,N_13181,N_13177);
xnor U13252 (N_13252,N_13131,N_13176);
and U13253 (N_13253,N_13183,N_13197);
xor U13254 (N_13254,N_13165,N_13206);
and U13255 (N_13255,N_13215,N_13149);
or U13256 (N_13256,N_13129,N_13125);
and U13257 (N_13257,N_13199,N_13220);
and U13258 (N_13258,N_13133,N_13172);
xor U13259 (N_13259,N_13210,N_13229);
nand U13260 (N_13260,N_13243,N_13191);
or U13261 (N_13261,N_13167,N_13230);
or U13262 (N_13262,N_13145,N_13239);
or U13263 (N_13263,N_13188,N_13234);
xor U13264 (N_13264,N_13200,N_13150);
or U13265 (N_13265,N_13248,N_13226);
or U13266 (N_13266,N_13192,N_13238);
or U13267 (N_13267,N_13204,N_13211);
or U13268 (N_13268,N_13221,N_13178);
nand U13269 (N_13269,N_13187,N_13240);
xnor U13270 (N_13270,N_13196,N_13154);
and U13271 (N_13271,N_13143,N_13242);
nand U13272 (N_13272,N_13227,N_13193);
xnor U13273 (N_13273,N_13207,N_13155);
or U13274 (N_13274,N_13184,N_13138);
nand U13275 (N_13275,N_13169,N_13218);
and U13276 (N_13276,N_13158,N_13171);
xor U13277 (N_13277,N_13212,N_13225);
nand U13278 (N_13278,N_13194,N_13182);
nor U13279 (N_13279,N_13173,N_13130);
nand U13280 (N_13280,N_13244,N_13190);
nor U13281 (N_13281,N_13170,N_13247);
nor U13282 (N_13282,N_13128,N_13189);
and U13283 (N_13283,N_13174,N_13168);
xor U13284 (N_13284,N_13140,N_13201);
nand U13285 (N_13285,N_13160,N_13214);
or U13286 (N_13286,N_13195,N_13159);
nand U13287 (N_13287,N_13153,N_13185);
xor U13288 (N_13288,N_13245,N_13151);
nor U13289 (N_13289,N_13235,N_13186);
or U13290 (N_13290,N_13202,N_13127);
nor U13291 (N_13291,N_13142,N_13216);
and U13292 (N_13292,N_13198,N_13141);
nand U13293 (N_13293,N_13209,N_13224);
xor U13294 (N_13294,N_13236,N_13217);
xor U13295 (N_13295,N_13126,N_13232);
or U13296 (N_13296,N_13246,N_13148);
and U13297 (N_13297,N_13180,N_13147);
xor U13298 (N_13298,N_13157,N_13222);
xor U13299 (N_13299,N_13241,N_13163);
nand U13300 (N_13300,N_13144,N_13208);
nor U13301 (N_13301,N_13164,N_13139);
xnor U13302 (N_13302,N_13136,N_13219);
and U13303 (N_13303,N_13166,N_13179);
nand U13304 (N_13304,N_13233,N_13134);
xnor U13305 (N_13305,N_13228,N_13205);
or U13306 (N_13306,N_13132,N_13137);
xnor U13307 (N_13307,N_13135,N_13162);
xnor U13308 (N_13308,N_13152,N_13231);
and U13309 (N_13309,N_13213,N_13161);
and U13310 (N_13310,N_13237,N_13203);
nand U13311 (N_13311,N_13223,N_13146);
or U13312 (N_13312,N_13156,N_13133);
nor U13313 (N_13313,N_13149,N_13144);
nand U13314 (N_13314,N_13205,N_13244);
and U13315 (N_13315,N_13165,N_13200);
xor U13316 (N_13316,N_13148,N_13225);
xnor U13317 (N_13317,N_13234,N_13228);
and U13318 (N_13318,N_13227,N_13222);
and U13319 (N_13319,N_13179,N_13215);
xor U13320 (N_13320,N_13164,N_13204);
nand U13321 (N_13321,N_13140,N_13154);
nor U13322 (N_13322,N_13242,N_13168);
or U13323 (N_13323,N_13133,N_13212);
nor U13324 (N_13324,N_13179,N_13228);
nand U13325 (N_13325,N_13240,N_13154);
and U13326 (N_13326,N_13134,N_13146);
nor U13327 (N_13327,N_13193,N_13130);
xor U13328 (N_13328,N_13218,N_13154);
or U13329 (N_13329,N_13178,N_13225);
nor U13330 (N_13330,N_13193,N_13224);
nand U13331 (N_13331,N_13237,N_13222);
or U13332 (N_13332,N_13135,N_13185);
or U13333 (N_13333,N_13223,N_13142);
nor U13334 (N_13334,N_13214,N_13180);
nand U13335 (N_13335,N_13241,N_13194);
nor U13336 (N_13336,N_13217,N_13131);
and U13337 (N_13337,N_13180,N_13193);
nand U13338 (N_13338,N_13246,N_13227);
and U13339 (N_13339,N_13239,N_13201);
xor U13340 (N_13340,N_13165,N_13240);
xor U13341 (N_13341,N_13135,N_13168);
nor U13342 (N_13342,N_13198,N_13160);
nor U13343 (N_13343,N_13186,N_13188);
nor U13344 (N_13344,N_13244,N_13189);
xor U13345 (N_13345,N_13225,N_13184);
nand U13346 (N_13346,N_13132,N_13178);
nand U13347 (N_13347,N_13152,N_13222);
nor U13348 (N_13348,N_13225,N_13245);
or U13349 (N_13349,N_13221,N_13245);
or U13350 (N_13350,N_13197,N_13201);
or U13351 (N_13351,N_13240,N_13226);
or U13352 (N_13352,N_13224,N_13157);
nor U13353 (N_13353,N_13208,N_13149);
or U13354 (N_13354,N_13125,N_13239);
xnor U13355 (N_13355,N_13193,N_13150);
nand U13356 (N_13356,N_13160,N_13126);
nand U13357 (N_13357,N_13188,N_13229);
nor U13358 (N_13358,N_13179,N_13226);
xnor U13359 (N_13359,N_13200,N_13210);
xor U13360 (N_13360,N_13247,N_13128);
nand U13361 (N_13361,N_13156,N_13235);
nor U13362 (N_13362,N_13238,N_13152);
nor U13363 (N_13363,N_13151,N_13132);
and U13364 (N_13364,N_13222,N_13226);
xor U13365 (N_13365,N_13224,N_13154);
or U13366 (N_13366,N_13136,N_13234);
xor U13367 (N_13367,N_13140,N_13132);
and U13368 (N_13368,N_13135,N_13203);
nand U13369 (N_13369,N_13189,N_13134);
nand U13370 (N_13370,N_13154,N_13166);
nor U13371 (N_13371,N_13145,N_13205);
nand U13372 (N_13372,N_13138,N_13139);
and U13373 (N_13373,N_13196,N_13210);
nor U13374 (N_13374,N_13166,N_13157);
xnor U13375 (N_13375,N_13312,N_13279);
and U13376 (N_13376,N_13366,N_13303);
and U13377 (N_13377,N_13306,N_13336);
nand U13378 (N_13378,N_13372,N_13333);
nand U13379 (N_13379,N_13269,N_13369);
xnor U13380 (N_13380,N_13325,N_13344);
and U13381 (N_13381,N_13305,N_13295);
nor U13382 (N_13382,N_13322,N_13271);
xnor U13383 (N_13383,N_13256,N_13309);
or U13384 (N_13384,N_13252,N_13291);
nand U13385 (N_13385,N_13284,N_13320);
nand U13386 (N_13386,N_13308,N_13323);
xnor U13387 (N_13387,N_13259,N_13343);
or U13388 (N_13388,N_13272,N_13316);
nand U13389 (N_13389,N_13337,N_13258);
nor U13390 (N_13390,N_13365,N_13361);
and U13391 (N_13391,N_13286,N_13273);
and U13392 (N_13392,N_13265,N_13351);
nor U13393 (N_13393,N_13340,N_13281);
xnor U13394 (N_13394,N_13346,N_13353);
xor U13395 (N_13395,N_13332,N_13276);
or U13396 (N_13396,N_13318,N_13287);
nand U13397 (N_13397,N_13364,N_13302);
or U13398 (N_13398,N_13368,N_13300);
nand U13399 (N_13399,N_13297,N_13310);
xnor U13400 (N_13400,N_13301,N_13280);
nand U13401 (N_13401,N_13331,N_13373);
or U13402 (N_13402,N_13285,N_13371);
or U13403 (N_13403,N_13311,N_13277);
or U13404 (N_13404,N_13335,N_13260);
nor U13405 (N_13405,N_13367,N_13328);
nor U13406 (N_13406,N_13289,N_13267);
nand U13407 (N_13407,N_13326,N_13360);
nand U13408 (N_13408,N_13374,N_13363);
nor U13409 (N_13409,N_13356,N_13314);
nor U13410 (N_13410,N_13264,N_13266);
nor U13411 (N_13411,N_13257,N_13352);
or U13412 (N_13412,N_13370,N_13347);
or U13413 (N_13413,N_13282,N_13298);
xor U13414 (N_13414,N_13358,N_13359);
xnor U13415 (N_13415,N_13288,N_13304);
nor U13416 (N_13416,N_13299,N_13339);
nand U13417 (N_13417,N_13348,N_13254);
nor U13418 (N_13418,N_13261,N_13327);
xnor U13419 (N_13419,N_13263,N_13330);
nand U13420 (N_13420,N_13278,N_13274);
or U13421 (N_13421,N_13255,N_13268);
and U13422 (N_13422,N_13341,N_13350);
xnor U13423 (N_13423,N_13321,N_13296);
nor U13424 (N_13424,N_13334,N_13251);
nor U13425 (N_13425,N_13262,N_13283);
nor U13426 (N_13426,N_13290,N_13357);
and U13427 (N_13427,N_13349,N_13329);
or U13428 (N_13428,N_13319,N_13345);
nor U13429 (N_13429,N_13253,N_13270);
xor U13430 (N_13430,N_13294,N_13317);
xor U13431 (N_13431,N_13355,N_13362);
or U13432 (N_13432,N_13324,N_13307);
nand U13433 (N_13433,N_13354,N_13293);
nor U13434 (N_13434,N_13275,N_13342);
and U13435 (N_13435,N_13338,N_13313);
nand U13436 (N_13436,N_13250,N_13315);
nor U13437 (N_13437,N_13292,N_13256);
and U13438 (N_13438,N_13371,N_13313);
nor U13439 (N_13439,N_13277,N_13308);
xnor U13440 (N_13440,N_13354,N_13271);
and U13441 (N_13441,N_13356,N_13330);
xnor U13442 (N_13442,N_13327,N_13252);
xor U13443 (N_13443,N_13265,N_13344);
nand U13444 (N_13444,N_13340,N_13310);
and U13445 (N_13445,N_13362,N_13260);
and U13446 (N_13446,N_13315,N_13276);
and U13447 (N_13447,N_13257,N_13297);
nor U13448 (N_13448,N_13253,N_13362);
nor U13449 (N_13449,N_13320,N_13305);
nor U13450 (N_13450,N_13324,N_13293);
xor U13451 (N_13451,N_13338,N_13331);
xor U13452 (N_13452,N_13371,N_13256);
or U13453 (N_13453,N_13259,N_13263);
or U13454 (N_13454,N_13291,N_13277);
or U13455 (N_13455,N_13320,N_13358);
or U13456 (N_13456,N_13272,N_13326);
nand U13457 (N_13457,N_13353,N_13337);
nand U13458 (N_13458,N_13352,N_13363);
nand U13459 (N_13459,N_13257,N_13368);
xnor U13460 (N_13460,N_13257,N_13293);
nor U13461 (N_13461,N_13260,N_13359);
and U13462 (N_13462,N_13367,N_13290);
and U13463 (N_13463,N_13252,N_13274);
nand U13464 (N_13464,N_13263,N_13281);
or U13465 (N_13465,N_13330,N_13259);
nor U13466 (N_13466,N_13292,N_13324);
nand U13467 (N_13467,N_13341,N_13269);
nor U13468 (N_13468,N_13282,N_13374);
nor U13469 (N_13469,N_13294,N_13262);
or U13470 (N_13470,N_13279,N_13337);
nor U13471 (N_13471,N_13277,N_13346);
or U13472 (N_13472,N_13301,N_13317);
nor U13473 (N_13473,N_13323,N_13328);
and U13474 (N_13474,N_13328,N_13262);
nand U13475 (N_13475,N_13336,N_13297);
nor U13476 (N_13476,N_13318,N_13338);
nor U13477 (N_13477,N_13301,N_13296);
nor U13478 (N_13478,N_13337,N_13328);
xor U13479 (N_13479,N_13297,N_13261);
xnor U13480 (N_13480,N_13365,N_13292);
xor U13481 (N_13481,N_13279,N_13293);
xnor U13482 (N_13482,N_13372,N_13277);
and U13483 (N_13483,N_13322,N_13347);
nand U13484 (N_13484,N_13325,N_13336);
xor U13485 (N_13485,N_13345,N_13258);
or U13486 (N_13486,N_13340,N_13287);
xor U13487 (N_13487,N_13358,N_13295);
nand U13488 (N_13488,N_13261,N_13309);
nand U13489 (N_13489,N_13351,N_13270);
or U13490 (N_13490,N_13316,N_13342);
nor U13491 (N_13491,N_13330,N_13324);
or U13492 (N_13492,N_13374,N_13256);
and U13493 (N_13493,N_13345,N_13313);
nor U13494 (N_13494,N_13329,N_13325);
nand U13495 (N_13495,N_13366,N_13279);
xor U13496 (N_13496,N_13326,N_13268);
xnor U13497 (N_13497,N_13263,N_13302);
xnor U13498 (N_13498,N_13368,N_13278);
or U13499 (N_13499,N_13363,N_13280);
nand U13500 (N_13500,N_13436,N_13459);
nand U13501 (N_13501,N_13440,N_13416);
and U13502 (N_13502,N_13377,N_13441);
or U13503 (N_13503,N_13421,N_13494);
or U13504 (N_13504,N_13378,N_13375);
or U13505 (N_13505,N_13387,N_13427);
or U13506 (N_13506,N_13419,N_13493);
and U13507 (N_13507,N_13432,N_13418);
nor U13508 (N_13508,N_13452,N_13396);
xnor U13509 (N_13509,N_13398,N_13486);
or U13510 (N_13510,N_13409,N_13382);
nand U13511 (N_13511,N_13467,N_13455);
or U13512 (N_13512,N_13456,N_13420);
nor U13513 (N_13513,N_13402,N_13468);
nor U13514 (N_13514,N_13483,N_13442);
nand U13515 (N_13515,N_13497,N_13458);
nand U13516 (N_13516,N_13482,N_13488);
nand U13517 (N_13517,N_13469,N_13465);
and U13518 (N_13518,N_13412,N_13484);
nand U13519 (N_13519,N_13400,N_13471);
xnor U13520 (N_13520,N_13407,N_13414);
nor U13521 (N_13521,N_13457,N_13496);
nand U13522 (N_13522,N_13401,N_13394);
or U13523 (N_13523,N_13431,N_13434);
or U13524 (N_13524,N_13429,N_13470);
and U13525 (N_13525,N_13499,N_13472);
or U13526 (N_13526,N_13446,N_13477);
xor U13527 (N_13527,N_13395,N_13397);
or U13528 (N_13528,N_13480,N_13463);
and U13529 (N_13529,N_13390,N_13426);
nor U13530 (N_13530,N_13453,N_13481);
and U13531 (N_13531,N_13476,N_13460);
nand U13532 (N_13532,N_13491,N_13437);
and U13533 (N_13533,N_13435,N_13451);
xnor U13534 (N_13534,N_13405,N_13492);
and U13535 (N_13535,N_13381,N_13487);
nand U13536 (N_13536,N_13438,N_13423);
nor U13537 (N_13537,N_13404,N_13466);
and U13538 (N_13538,N_13391,N_13449);
and U13539 (N_13539,N_13445,N_13489);
xor U13540 (N_13540,N_13495,N_13478);
nor U13541 (N_13541,N_13474,N_13410);
nand U13542 (N_13542,N_13422,N_13450);
xnor U13543 (N_13543,N_13384,N_13464);
nand U13544 (N_13544,N_13448,N_13413);
nor U13545 (N_13545,N_13430,N_13462);
or U13546 (N_13546,N_13403,N_13399);
nand U13547 (N_13547,N_13433,N_13406);
xnor U13548 (N_13548,N_13379,N_13424);
and U13549 (N_13549,N_13386,N_13454);
nand U13550 (N_13550,N_13408,N_13415);
or U13551 (N_13551,N_13443,N_13389);
nor U13552 (N_13552,N_13417,N_13479);
xnor U13553 (N_13553,N_13439,N_13425);
or U13554 (N_13554,N_13475,N_13388);
and U13555 (N_13555,N_13490,N_13428);
xor U13556 (N_13556,N_13385,N_13383);
nor U13557 (N_13557,N_13461,N_13393);
nand U13558 (N_13558,N_13376,N_13498);
and U13559 (N_13559,N_13380,N_13411);
or U13560 (N_13560,N_13447,N_13485);
nor U13561 (N_13561,N_13473,N_13392);
xor U13562 (N_13562,N_13444,N_13450);
and U13563 (N_13563,N_13474,N_13386);
nand U13564 (N_13564,N_13402,N_13455);
or U13565 (N_13565,N_13434,N_13464);
nand U13566 (N_13566,N_13448,N_13471);
nand U13567 (N_13567,N_13437,N_13486);
nand U13568 (N_13568,N_13377,N_13485);
nor U13569 (N_13569,N_13400,N_13492);
and U13570 (N_13570,N_13389,N_13448);
nand U13571 (N_13571,N_13485,N_13483);
nor U13572 (N_13572,N_13493,N_13400);
nor U13573 (N_13573,N_13458,N_13491);
xnor U13574 (N_13574,N_13459,N_13472);
xor U13575 (N_13575,N_13377,N_13380);
nand U13576 (N_13576,N_13485,N_13495);
xnor U13577 (N_13577,N_13399,N_13378);
nor U13578 (N_13578,N_13488,N_13474);
or U13579 (N_13579,N_13424,N_13482);
nand U13580 (N_13580,N_13396,N_13429);
and U13581 (N_13581,N_13379,N_13454);
and U13582 (N_13582,N_13445,N_13448);
or U13583 (N_13583,N_13376,N_13449);
nor U13584 (N_13584,N_13409,N_13395);
or U13585 (N_13585,N_13471,N_13476);
or U13586 (N_13586,N_13379,N_13392);
nor U13587 (N_13587,N_13380,N_13449);
nor U13588 (N_13588,N_13378,N_13404);
or U13589 (N_13589,N_13453,N_13410);
and U13590 (N_13590,N_13461,N_13430);
or U13591 (N_13591,N_13478,N_13442);
and U13592 (N_13592,N_13482,N_13389);
or U13593 (N_13593,N_13474,N_13397);
or U13594 (N_13594,N_13434,N_13454);
or U13595 (N_13595,N_13386,N_13380);
nand U13596 (N_13596,N_13411,N_13494);
nand U13597 (N_13597,N_13434,N_13465);
nand U13598 (N_13598,N_13435,N_13394);
or U13599 (N_13599,N_13409,N_13444);
or U13600 (N_13600,N_13396,N_13478);
and U13601 (N_13601,N_13382,N_13427);
and U13602 (N_13602,N_13458,N_13462);
nor U13603 (N_13603,N_13441,N_13423);
xor U13604 (N_13604,N_13493,N_13418);
and U13605 (N_13605,N_13407,N_13496);
nor U13606 (N_13606,N_13498,N_13409);
or U13607 (N_13607,N_13387,N_13447);
xor U13608 (N_13608,N_13401,N_13496);
xor U13609 (N_13609,N_13425,N_13400);
nand U13610 (N_13610,N_13424,N_13473);
and U13611 (N_13611,N_13387,N_13471);
or U13612 (N_13612,N_13477,N_13380);
xor U13613 (N_13613,N_13419,N_13416);
or U13614 (N_13614,N_13489,N_13470);
or U13615 (N_13615,N_13438,N_13393);
xnor U13616 (N_13616,N_13494,N_13417);
nand U13617 (N_13617,N_13422,N_13426);
or U13618 (N_13618,N_13459,N_13409);
nand U13619 (N_13619,N_13391,N_13447);
nand U13620 (N_13620,N_13432,N_13466);
nor U13621 (N_13621,N_13407,N_13460);
xor U13622 (N_13622,N_13457,N_13462);
and U13623 (N_13623,N_13444,N_13473);
nand U13624 (N_13624,N_13488,N_13401);
or U13625 (N_13625,N_13545,N_13518);
nand U13626 (N_13626,N_13524,N_13538);
or U13627 (N_13627,N_13574,N_13584);
nand U13628 (N_13628,N_13516,N_13514);
nand U13629 (N_13629,N_13593,N_13567);
nand U13630 (N_13630,N_13531,N_13605);
or U13631 (N_13631,N_13614,N_13523);
or U13632 (N_13632,N_13562,N_13580);
nand U13633 (N_13633,N_13603,N_13501);
nor U13634 (N_13634,N_13552,N_13521);
or U13635 (N_13635,N_13513,N_13624);
nand U13636 (N_13636,N_13504,N_13543);
and U13637 (N_13637,N_13522,N_13507);
nand U13638 (N_13638,N_13575,N_13587);
nand U13639 (N_13639,N_13600,N_13578);
nor U13640 (N_13640,N_13550,N_13598);
or U13641 (N_13641,N_13559,N_13609);
and U13642 (N_13642,N_13561,N_13569);
nand U13643 (N_13643,N_13555,N_13534);
and U13644 (N_13644,N_13595,N_13613);
nor U13645 (N_13645,N_13553,N_13606);
xnor U13646 (N_13646,N_13611,N_13596);
nand U13647 (N_13647,N_13599,N_13582);
or U13648 (N_13648,N_13517,N_13558);
nand U13649 (N_13649,N_13615,N_13592);
nand U13650 (N_13650,N_13540,N_13502);
and U13651 (N_13651,N_13500,N_13512);
nor U13652 (N_13652,N_13515,N_13536);
or U13653 (N_13653,N_13589,N_13542);
xnor U13654 (N_13654,N_13594,N_13544);
nand U13655 (N_13655,N_13547,N_13588);
nand U13656 (N_13656,N_13506,N_13537);
nor U13657 (N_13657,N_13585,N_13503);
xor U13658 (N_13658,N_13530,N_13576);
and U13659 (N_13659,N_13532,N_13612);
xor U13660 (N_13660,N_13565,N_13526);
or U13661 (N_13661,N_13590,N_13556);
nand U13662 (N_13662,N_13622,N_13616);
and U13663 (N_13663,N_13551,N_13554);
or U13664 (N_13664,N_13566,N_13525);
nand U13665 (N_13665,N_13581,N_13617);
or U13666 (N_13666,N_13546,N_13623);
xor U13667 (N_13667,N_13607,N_13511);
xnor U13668 (N_13668,N_13568,N_13570);
nand U13669 (N_13669,N_13583,N_13586);
nand U13670 (N_13670,N_13535,N_13601);
xnor U13671 (N_13671,N_13597,N_13564);
or U13672 (N_13672,N_13519,N_13548);
nand U13673 (N_13673,N_13529,N_13557);
nor U13674 (N_13674,N_13508,N_13620);
nor U13675 (N_13675,N_13560,N_13563);
and U13676 (N_13676,N_13528,N_13621);
nand U13677 (N_13677,N_13610,N_13533);
or U13678 (N_13678,N_13527,N_13541);
nor U13679 (N_13679,N_13505,N_13619);
nor U13680 (N_13680,N_13579,N_13539);
xnor U13681 (N_13681,N_13549,N_13618);
xor U13682 (N_13682,N_13510,N_13572);
and U13683 (N_13683,N_13520,N_13573);
or U13684 (N_13684,N_13591,N_13602);
xnor U13685 (N_13685,N_13571,N_13608);
nor U13686 (N_13686,N_13509,N_13604);
nor U13687 (N_13687,N_13577,N_13621);
nor U13688 (N_13688,N_13624,N_13522);
and U13689 (N_13689,N_13614,N_13537);
nand U13690 (N_13690,N_13593,N_13620);
and U13691 (N_13691,N_13602,N_13562);
nand U13692 (N_13692,N_13544,N_13621);
nand U13693 (N_13693,N_13558,N_13559);
nand U13694 (N_13694,N_13545,N_13566);
and U13695 (N_13695,N_13530,N_13559);
xor U13696 (N_13696,N_13562,N_13531);
nand U13697 (N_13697,N_13533,N_13591);
and U13698 (N_13698,N_13590,N_13524);
and U13699 (N_13699,N_13623,N_13582);
or U13700 (N_13700,N_13579,N_13576);
nor U13701 (N_13701,N_13612,N_13507);
and U13702 (N_13702,N_13577,N_13531);
or U13703 (N_13703,N_13606,N_13563);
and U13704 (N_13704,N_13569,N_13522);
and U13705 (N_13705,N_13520,N_13600);
and U13706 (N_13706,N_13525,N_13545);
or U13707 (N_13707,N_13511,N_13521);
xnor U13708 (N_13708,N_13555,N_13606);
or U13709 (N_13709,N_13532,N_13595);
nand U13710 (N_13710,N_13590,N_13612);
xor U13711 (N_13711,N_13525,N_13577);
nand U13712 (N_13712,N_13535,N_13533);
xnor U13713 (N_13713,N_13501,N_13517);
and U13714 (N_13714,N_13619,N_13596);
xnor U13715 (N_13715,N_13589,N_13603);
xnor U13716 (N_13716,N_13532,N_13569);
or U13717 (N_13717,N_13607,N_13566);
xnor U13718 (N_13718,N_13599,N_13510);
and U13719 (N_13719,N_13603,N_13582);
nor U13720 (N_13720,N_13519,N_13587);
nand U13721 (N_13721,N_13609,N_13589);
xor U13722 (N_13722,N_13602,N_13577);
nand U13723 (N_13723,N_13538,N_13600);
or U13724 (N_13724,N_13531,N_13528);
nor U13725 (N_13725,N_13552,N_13525);
xnor U13726 (N_13726,N_13590,N_13593);
nor U13727 (N_13727,N_13506,N_13543);
xnor U13728 (N_13728,N_13564,N_13591);
and U13729 (N_13729,N_13525,N_13595);
or U13730 (N_13730,N_13620,N_13594);
nor U13731 (N_13731,N_13554,N_13501);
xor U13732 (N_13732,N_13566,N_13600);
nor U13733 (N_13733,N_13549,N_13595);
nor U13734 (N_13734,N_13526,N_13554);
nand U13735 (N_13735,N_13609,N_13613);
and U13736 (N_13736,N_13543,N_13607);
or U13737 (N_13737,N_13554,N_13617);
nor U13738 (N_13738,N_13529,N_13534);
or U13739 (N_13739,N_13596,N_13582);
and U13740 (N_13740,N_13621,N_13519);
or U13741 (N_13741,N_13554,N_13592);
nor U13742 (N_13742,N_13559,N_13543);
xor U13743 (N_13743,N_13570,N_13503);
xnor U13744 (N_13744,N_13515,N_13524);
nor U13745 (N_13745,N_13547,N_13517);
and U13746 (N_13746,N_13613,N_13553);
and U13747 (N_13747,N_13624,N_13610);
nand U13748 (N_13748,N_13572,N_13583);
and U13749 (N_13749,N_13615,N_13505);
nand U13750 (N_13750,N_13749,N_13643);
xnor U13751 (N_13751,N_13692,N_13679);
nand U13752 (N_13752,N_13678,N_13733);
and U13753 (N_13753,N_13668,N_13631);
nand U13754 (N_13754,N_13666,N_13675);
nand U13755 (N_13755,N_13672,N_13657);
xnor U13756 (N_13756,N_13646,N_13656);
or U13757 (N_13757,N_13735,N_13714);
and U13758 (N_13758,N_13705,N_13702);
nand U13759 (N_13759,N_13680,N_13745);
nand U13760 (N_13760,N_13698,N_13690);
or U13761 (N_13761,N_13647,N_13685);
xnor U13762 (N_13762,N_13709,N_13682);
and U13763 (N_13763,N_13642,N_13644);
and U13764 (N_13764,N_13718,N_13704);
xor U13765 (N_13765,N_13660,N_13728);
nand U13766 (N_13766,N_13628,N_13625);
nor U13767 (N_13767,N_13707,N_13694);
xor U13768 (N_13768,N_13658,N_13706);
nor U13769 (N_13769,N_13697,N_13717);
nand U13770 (N_13770,N_13730,N_13630);
or U13771 (N_13771,N_13726,N_13722);
or U13772 (N_13772,N_13742,N_13712);
nand U13773 (N_13773,N_13629,N_13673);
xnor U13774 (N_13774,N_13637,N_13648);
xor U13775 (N_13775,N_13674,N_13737);
xor U13776 (N_13776,N_13736,N_13708);
nor U13777 (N_13777,N_13710,N_13740);
xnor U13778 (N_13778,N_13744,N_13699);
and U13779 (N_13779,N_13626,N_13670);
and U13780 (N_13780,N_13663,N_13654);
and U13781 (N_13781,N_13671,N_13676);
and U13782 (N_13782,N_13633,N_13703);
nand U13783 (N_13783,N_13669,N_13721);
xnor U13784 (N_13784,N_13645,N_13711);
xor U13785 (N_13785,N_13639,N_13693);
or U13786 (N_13786,N_13677,N_13635);
nor U13787 (N_13787,N_13659,N_13667);
nand U13788 (N_13788,N_13688,N_13687);
xor U13789 (N_13789,N_13655,N_13719);
or U13790 (N_13790,N_13724,N_13634);
xor U13791 (N_13791,N_13640,N_13652);
xor U13792 (N_13792,N_13650,N_13700);
or U13793 (N_13793,N_13713,N_13743);
or U13794 (N_13794,N_13716,N_13723);
and U13795 (N_13795,N_13689,N_13732);
or U13796 (N_13796,N_13686,N_13662);
or U13797 (N_13797,N_13664,N_13649);
nor U13798 (N_13798,N_13731,N_13741);
or U13799 (N_13799,N_13651,N_13638);
nor U13800 (N_13800,N_13691,N_13746);
or U13801 (N_13801,N_13747,N_13684);
and U13802 (N_13802,N_13641,N_13683);
nor U13803 (N_13803,N_13653,N_13632);
nor U13804 (N_13804,N_13727,N_13725);
or U13805 (N_13805,N_13738,N_13695);
xnor U13806 (N_13806,N_13681,N_13636);
and U13807 (N_13807,N_13739,N_13665);
nand U13808 (N_13808,N_13734,N_13729);
nor U13809 (N_13809,N_13627,N_13661);
or U13810 (N_13810,N_13720,N_13715);
nor U13811 (N_13811,N_13701,N_13696);
nor U13812 (N_13812,N_13748,N_13661);
nor U13813 (N_13813,N_13669,N_13693);
and U13814 (N_13814,N_13703,N_13727);
or U13815 (N_13815,N_13705,N_13722);
or U13816 (N_13816,N_13746,N_13685);
and U13817 (N_13817,N_13635,N_13653);
xor U13818 (N_13818,N_13700,N_13688);
nor U13819 (N_13819,N_13733,N_13644);
and U13820 (N_13820,N_13684,N_13714);
xnor U13821 (N_13821,N_13685,N_13712);
nand U13822 (N_13822,N_13629,N_13658);
nor U13823 (N_13823,N_13679,N_13734);
nand U13824 (N_13824,N_13703,N_13688);
or U13825 (N_13825,N_13688,N_13707);
or U13826 (N_13826,N_13675,N_13690);
and U13827 (N_13827,N_13665,N_13679);
and U13828 (N_13828,N_13637,N_13740);
or U13829 (N_13829,N_13694,N_13639);
or U13830 (N_13830,N_13630,N_13664);
or U13831 (N_13831,N_13748,N_13651);
nand U13832 (N_13832,N_13669,N_13661);
nand U13833 (N_13833,N_13740,N_13742);
xor U13834 (N_13834,N_13722,N_13688);
nand U13835 (N_13835,N_13642,N_13730);
nor U13836 (N_13836,N_13747,N_13661);
nand U13837 (N_13837,N_13660,N_13719);
or U13838 (N_13838,N_13666,N_13726);
nor U13839 (N_13839,N_13717,N_13655);
xnor U13840 (N_13840,N_13635,N_13644);
nand U13841 (N_13841,N_13749,N_13639);
xnor U13842 (N_13842,N_13679,N_13691);
and U13843 (N_13843,N_13672,N_13636);
and U13844 (N_13844,N_13687,N_13721);
or U13845 (N_13845,N_13692,N_13727);
and U13846 (N_13846,N_13677,N_13746);
xnor U13847 (N_13847,N_13736,N_13682);
xnor U13848 (N_13848,N_13743,N_13653);
and U13849 (N_13849,N_13668,N_13703);
nor U13850 (N_13850,N_13633,N_13650);
xor U13851 (N_13851,N_13747,N_13660);
nand U13852 (N_13852,N_13634,N_13636);
and U13853 (N_13853,N_13745,N_13690);
nor U13854 (N_13854,N_13662,N_13692);
or U13855 (N_13855,N_13663,N_13710);
xnor U13856 (N_13856,N_13667,N_13728);
and U13857 (N_13857,N_13658,N_13647);
and U13858 (N_13858,N_13649,N_13740);
or U13859 (N_13859,N_13656,N_13674);
and U13860 (N_13860,N_13644,N_13675);
nand U13861 (N_13861,N_13693,N_13628);
xnor U13862 (N_13862,N_13719,N_13706);
and U13863 (N_13863,N_13652,N_13731);
xor U13864 (N_13864,N_13653,N_13631);
xor U13865 (N_13865,N_13650,N_13651);
nor U13866 (N_13866,N_13673,N_13714);
nor U13867 (N_13867,N_13733,N_13625);
nand U13868 (N_13868,N_13747,N_13738);
nor U13869 (N_13869,N_13636,N_13717);
or U13870 (N_13870,N_13737,N_13749);
or U13871 (N_13871,N_13724,N_13746);
xor U13872 (N_13872,N_13715,N_13730);
nor U13873 (N_13873,N_13692,N_13664);
nand U13874 (N_13874,N_13717,N_13687);
and U13875 (N_13875,N_13780,N_13765);
nor U13876 (N_13876,N_13800,N_13776);
or U13877 (N_13877,N_13769,N_13827);
nor U13878 (N_13878,N_13753,N_13775);
nand U13879 (N_13879,N_13754,N_13801);
and U13880 (N_13880,N_13802,N_13867);
xor U13881 (N_13881,N_13863,N_13858);
nor U13882 (N_13882,N_13864,N_13779);
nand U13883 (N_13883,N_13823,N_13857);
or U13884 (N_13884,N_13870,N_13830);
nor U13885 (N_13885,N_13755,N_13752);
xnor U13886 (N_13886,N_13759,N_13778);
or U13887 (N_13887,N_13847,N_13806);
xor U13888 (N_13888,N_13833,N_13836);
nand U13889 (N_13889,N_13825,N_13838);
nor U13890 (N_13890,N_13771,N_13843);
and U13891 (N_13891,N_13837,N_13839);
xnor U13892 (N_13892,N_13788,N_13868);
or U13893 (N_13893,N_13797,N_13798);
and U13894 (N_13894,N_13799,N_13766);
nand U13895 (N_13895,N_13872,N_13871);
xor U13896 (N_13896,N_13850,N_13809);
xnor U13897 (N_13897,N_13832,N_13862);
or U13898 (N_13898,N_13770,N_13835);
and U13899 (N_13899,N_13758,N_13849);
or U13900 (N_13900,N_13782,N_13790);
nor U13901 (N_13901,N_13814,N_13874);
nand U13902 (N_13902,N_13777,N_13756);
or U13903 (N_13903,N_13768,N_13810);
nand U13904 (N_13904,N_13783,N_13781);
xnor U13905 (N_13905,N_13789,N_13824);
xor U13906 (N_13906,N_13764,N_13816);
or U13907 (N_13907,N_13828,N_13831);
or U13908 (N_13908,N_13853,N_13855);
and U13909 (N_13909,N_13761,N_13873);
xor U13910 (N_13910,N_13860,N_13820);
and U13911 (N_13911,N_13851,N_13815);
nand U13912 (N_13912,N_13763,N_13865);
xnor U13913 (N_13913,N_13772,N_13787);
or U13914 (N_13914,N_13841,N_13846);
xnor U13915 (N_13915,N_13786,N_13869);
xnor U13916 (N_13916,N_13819,N_13842);
and U13917 (N_13917,N_13861,N_13762);
xor U13918 (N_13918,N_13854,N_13807);
nand U13919 (N_13919,N_13834,N_13821);
xnor U13920 (N_13920,N_13795,N_13852);
and U13921 (N_13921,N_13822,N_13848);
xnor U13922 (N_13922,N_13785,N_13773);
nor U13923 (N_13923,N_13859,N_13866);
nor U13924 (N_13924,N_13845,N_13826);
and U13925 (N_13925,N_13844,N_13811);
and U13926 (N_13926,N_13813,N_13767);
xnor U13927 (N_13927,N_13808,N_13751);
or U13928 (N_13928,N_13784,N_13818);
or U13929 (N_13929,N_13840,N_13750);
nor U13930 (N_13930,N_13757,N_13774);
and U13931 (N_13931,N_13760,N_13796);
nor U13932 (N_13932,N_13804,N_13829);
or U13933 (N_13933,N_13856,N_13812);
xnor U13934 (N_13934,N_13791,N_13817);
or U13935 (N_13935,N_13805,N_13792);
and U13936 (N_13936,N_13793,N_13794);
and U13937 (N_13937,N_13803,N_13864);
nor U13938 (N_13938,N_13758,N_13825);
xor U13939 (N_13939,N_13800,N_13862);
or U13940 (N_13940,N_13842,N_13770);
nor U13941 (N_13941,N_13773,N_13777);
or U13942 (N_13942,N_13828,N_13840);
and U13943 (N_13943,N_13845,N_13752);
xnor U13944 (N_13944,N_13808,N_13793);
or U13945 (N_13945,N_13838,N_13805);
xor U13946 (N_13946,N_13795,N_13792);
and U13947 (N_13947,N_13857,N_13777);
and U13948 (N_13948,N_13840,N_13770);
and U13949 (N_13949,N_13813,N_13843);
and U13950 (N_13950,N_13832,N_13838);
xnor U13951 (N_13951,N_13777,N_13820);
or U13952 (N_13952,N_13808,N_13759);
or U13953 (N_13953,N_13781,N_13817);
xor U13954 (N_13954,N_13801,N_13825);
or U13955 (N_13955,N_13855,N_13771);
nor U13956 (N_13956,N_13813,N_13857);
and U13957 (N_13957,N_13777,N_13776);
and U13958 (N_13958,N_13796,N_13808);
nand U13959 (N_13959,N_13789,N_13821);
nand U13960 (N_13960,N_13758,N_13767);
xnor U13961 (N_13961,N_13868,N_13866);
nor U13962 (N_13962,N_13816,N_13784);
nor U13963 (N_13963,N_13849,N_13865);
xnor U13964 (N_13964,N_13870,N_13826);
or U13965 (N_13965,N_13868,N_13803);
xnor U13966 (N_13966,N_13850,N_13776);
nand U13967 (N_13967,N_13752,N_13817);
and U13968 (N_13968,N_13767,N_13831);
xnor U13969 (N_13969,N_13804,N_13820);
nor U13970 (N_13970,N_13809,N_13858);
or U13971 (N_13971,N_13792,N_13781);
nor U13972 (N_13972,N_13837,N_13794);
or U13973 (N_13973,N_13812,N_13839);
xnor U13974 (N_13974,N_13822,N_13772);
xnor U13975 (N_13975,N_13800,N_13795);
xnor U13976 (N_13976,N_13795,N_13836);
nor U13977 (N_13977,N_13776,N_13822);
xor U13978 (N_13978,N_13853,N_13854);
nor U13979 (N_13979,N_13751,N_13810);
nor U13980 (N_13980,N_13850,N_13872);
and U13981 (N_13981,N_13837,N_13764);
nand U13982 (N_13982,N_13824,N_13751);
xor U13983 (N_13983,N_13828,N_13874);
nor U13984 (N_13984,N_13811,N_13801);
nand U13985 (N_13985,N_13820,N_13780);
nand U13986 (N_13986,N_13814,N_13818);
nor U13987 (N_13987,N_13852,N_13779);
and U13988 (N_13988,N_13751,N_13868);
or U13989 (N_13989,N_13853,N_13866);
and U13990 (N_13990,N_13842,N_13773);
and U13991 (N_13991,N_13872,N_13842);
nand U13992 (N_13992,N_13788,N_13767);
or U13993 (N_13993,N_13829,N_13818);
nor U13994 (N_13994,N_13863,N_13862);
and U13995 (N_13995,N_13820,N_13790);
or U13996 (N_13996,N_13856,N_13801);
and U13997 (N_13997,N_13852,N_13858);
nand U13998 (N_13998,N_13858,N_13865);
and U13999 (N_13999,N_13829,N_13836);
nand U14000 (N_14000,N_13945,N_13907);
xor U14001 (N_14001,N_13918,N_13940);
nor U14002 (N_14002,N_13935,N_13938);
nand U14003 (N_14003,N_13958,N_13889);
nand U14004 (N_14004,N_13875,N_13877);
or U14005 (N_14005,N_13956,N_13887);
xor U14006 (N_14006,N_13951,N_13916);
nor U14007 (N_14007,N_13969,N_13953);
or U14008 (N_14008,N_13987,N_13983);
and U14009 (N_14009,N_13927,N_13949);
nand U14010 (N_14010,N_13966,N_13891);
nor U14011 (N_14011,N_13984,N_13936);
xnor U14012 (N_14012,N_13879,N_13941);
and U14013 (N_14013,N_13962,N_13954);
nand U14014 (N_14014,N_13968,N_13931);
and U14015 (N_14015,N_13905,N_13973);
nand U14016 (N_14016,N_13970,N_13976);
nor U14017 (N_14017,N_13934,N_13921);
and U14018 (N_14018,N_13977,N_13985);
or U14019 (N_14019,N_13993,N_13997);
or U14020 (N_14020,N_13919,N_13925);
nor U14021 (N_14021,N_13960,N_13897);
and U14022 (N_14022,N_13882,N_13980);
xor U14023 (N_14023,N_13876,N_13964);
nand U14024 (N_14024,N_13986,N_13999);
and U14025 (N_14025,N_13990,N_13883);
and U14026 (N_14026,N_13937,N_13892);
nor U14027 (N_14027,N_13894,N_13996);
or U14028 (N_14028,N_13965,N_13909);
xnor U14029 (N_14029,N_13898,N_13910);
xnor U14030 (N_14030,N_13946,N_13903);
nand U14031 (N_14031,N_13886,N_13928);
and U14032 (N_14032,N_13922,N_13979);
nand U14033 (N_14033,N_13915,N_13992);
or U14034 (N_14034,N_13975,N_13971);
nor U14035 (N_14035,N_13995,N_13890);
xor U14036 (N_14036,N_13994,N_13933);
or U14037 (N_14037,N_13900,N_13989);
or U14038 (N_14038,N_13948,N_13950);
nor U14039 (N_14039,N_13906,N_13961);
xor U14040 (N_14040,N_13957,N_13944);
nor U14041 (N_14041,N_13998,N_13981);
nand U14042 (N_14042,N_13880,N_13942);
nor U14043 (N_14043,N_13884,N_13930);
nor U14044 (N_14044,N_13967,N_13878);
and U14045 (N_14045,N_13929,N_13913);
or U14046 (N_14046,N_13908,N_13881);
nor U14047 (N_14047,N_13972,N_13955);
and U14048 (N_14048,N_13896,N_13943);
nand U14049 (N_14049,N_13924,N_13952);
xor U14050 (N_14050,N_13902,N_13978);
and U14051 (N_14051,N_13974,N_13982);
and U14052 (N_14052,N_13917,N_13923);
and U14053 (N_14053,N_13893,N_13895);
or U14054 (N_14054,N_13912,N_13885);
or U14055 (N_14055,N_13932,N_13991);
xor U14056 (N_14056,N_13926,N_13939);
nand U14057 (N_14057,N_13911,N_13988);
xnor U14058 (N_14058,N_13963,N_13959);
xnor U14059 (N_14059,N_13888,N_13920);
nand U14060 (N_14060,N_13901,N_13899);
nor U14061 (N_14061,N_13914,N_13947);
xnor U14062 (N_14062,N_13904,N_13906);
or U14063 (N_14063,N_13976,N_13940);
and U14064 (N_14064,N_13971,N_13882);
nor U14065 (N_14065,N_13926,N_13987);
xnor U14066 (N_14066,N_13950,N_13936);
nor U14067 (N_14067,N_13880,N_13908);
nor U14068 (N_14068,N_13905,N_13907);
nor U14069 (N_14069,N_13921,N_13978);
xor U14070 (N_14070,N_13926,N_13877);
nand U14071 (N_14071,N_13981,N_13929);
xnor U14072 (N_14072,N_13977,N_13967);
or U14073 (N_14073,N_13910,N_13883);
xor U14074 (N_14074,N_13945,N_13876);
and U14075 (N_14075,N_13906,N_13960);
nand U14076 (N_14076,N_13884,N_13968);
nor U14077 (N_14077,N_13888,N_13904);
nand U14078 (N_14078,N_13999,N_13925);
or U14079 (N_14079,N_13945,N_13899);
xor U14080 (N_14080,N_13948,N_13890);
nand U14081 (N_14081,N_13940,N_13958);
and U14082 (N_14082,N_13938,N_13936);
nor U14083 (N_14083,N_13905,N_13920);
and U14084 (N_14084,N_13908,N_13986);
and U14085 (N_14085,N_13931,N_13877);
nand U14086 (N_14086,N_13977,N_13958);
or U14087 (N_14087,N_13992,N_13897);
and U14088 (N_14088,N_13980,N_13916);
and U14089 (N_14089,N_13990,N_13904);
or U14090 (N_14090,N_13981,N_13997);
and U14091 (N_14091,N_13971,N_13908);
nand U14092 (N_14092,N_13985,N_13978);
and U14093 (N_14093,N_13972,N_13988);
and U14094 (N_14094,N_13949,N_13885);
or U14095 (N_14095,N_13970,N_13953);
and U14096 (N_14096,N_13981,N_13887);
and U14097 (N_14097,N_13917,N_13909);
or U14098 (N_14098,N_13913,N_13936);
and U14099 (N_14099,N_13986,N_13935);
xor U14100 (N_14100,N_13922,N_13896);
nand U14101 (N_14101,N_13885,N_13922);
nand U14102 (N_14102,N_13914,N_13895);
and U14103 (N_14103,N_13907,N_13900);
nand U14104 (N_14104,N_13974,N_13994);
nand U14105 (N_14105,N_13952,N_13967);
and U14106 (N_14106,N_13996,N_13988);
and U14107 (N_14107,N_13983,N_13989);
and U14108 (N_14108,N_13883,N_13935);
or U14109 (N_14109,N_13883,N_13889);
and U14110 (N_14110,N_13940,N_13883);
and U14111 (N_14111,N_13906,N_13890);
nor U14112 (N_14112,N_13997,N_13924);
nand U14113 (N_14113,N_13924,N_13949);
nand U14114 (N_14114,N_13896,N_13898);
xor U14115 (N_14115,N_13877,N_13959);
xnor U14116 (N_14116,N_13946,N_13942);
or U14117 (N_14117,N_13909,N_13986);
and U14118 (N_14118,N_13984,N_13876);
nand U14119 (N_14119,N_13922,N_13930);
nand U14120 (N_14120,N_13976,N_13942);
nor U14121 (N_14121,N_13969,N_13922);
nor U14122 (N_14122,N_13896,N_13956);
xor U14123 (N_14123,N_13938,N_13987);
and U14124 (N_14124,N_13992,N_13922);
and U14125 (N_14125,N_14071,N_14044);
nand U14126 (N_14126,N_14119,N_14053);
or U14127 (N_14127,N_14045,N_14010);
xor U14128 (N_14128,N_14022,N_14077);
xnor U14129 (N_14129,N_14118,N_14086);
nor U14130 (N_14130,N_14042,N_14024);
nor U14131 (N_14131,N_14048,N_14103);
and U14132 (N_14132,N_14095,N_14049);
or U14133 (N_14133,N_14062,N_14081);
xnor U14134 (N_14134,N_14029,N_14093);
or U14135 (N_14135,N_14079,N_14114);
xnor U14136 (N_14136,N_14105,N_14069);
and U14137 (N_14137,N_14004,N_14087);
xnor U14138 (N_14138,N_14040,N_14099);
nor U14139 (N_14139,N_14019,N_14005);
or U14140 (N_14140,N_14089,N_14108);
and U14141 (N_14141,N_14031,N_14076);
or U14142 (N_14142,N_14111,N_14112);
xnor U14143 (N_14143,N_14039,N_14121);
and U14144 (N_14144,N_14051,N_14038);
and U14145 (N_14145,N_14014,N_14032);
or U14146 (N_14146,N_14008,N_14123);
nand U14147 (N_14147,N_14006,N_14046);
xor U14148 (N_14148,N_14015,N_14116);
or U14149 (N_14149,N_14073,N_14003);
nand U14150 (N_14150,N_14100,N_14043);
nand U14151 (N_14151,N_14059,N_14083);
nor U14152 (N_14152,N_14023,N_14020);
xnor U14153 (N_14153,N_14009,N_14109);
nor U14154 (N_14154,N_14054,N_14007);
or U14155 (N_14155,N_14011,N_14064);
nand U14156 (N_14156,N_14001,N_14021);
or U14157 (N_14157,N_14041,N_14120);
xnor U14158 (N_14158,N_14030,N_14013);
and U14159 (N_14159,N_14082,N_14058);
nand U14160 (N_14160,N_14104,N_14025);
and U14161 (N_14161,N_14052,N_14110);
nand U14162 (N_14162,N_14094,N_14122);
nor U14163 (N_14163,N_14065,N_14072);
and U14164 (N_14164,N_14060,N_14084);
nand U14165 (N_14165,N_14018,N_14092);
nor U14166 (N_14166,N_14002,N_14068);
nor U14167 (N_14167,N_14063,N_14080);
or U14168 (N_14168,N_14101,N_14124);
and U14169 (N_14169,N_14106,N_14102);
nor U14170 (N_14170,N_14061,N_14078);
nor U14171 (N_14171,N_14091,N_14012);
xnor U14172 (N_14172,N_14067,N_14037);
and U14173 (N_14173,N_14028,N_14090);
or U14174 (N_14174,N_14027,N_14075);
and U14175 (N_14175,N_14036,N_14070);
nand U14176 (N_14176,N_14026,N_14057);
and U14177 (N_14177,N_14098,N_14033);
nor U14178 (N_14178,N_14016,N_14035);
nor U14179 (N_14179,N_14066,N_14050);
or U14180 (N_14180,N_14055,N_14047);
xnor U14181 (N_14181,N_14113,N_14097);
nor U14182 (N_14182,N_14017,N_14034);
xnor U14183 (N_14183,N_14117,N_14088);
xnor U14184 (N_14184,N_14000,N_14056);
nor U14185 (N_14185,N_14107,N_14074);
and U14186 (N_14186,N_14085,N_14115);
xor U14187 (N_14187,N_14096,N_14078);
nand U14188 (N_14188,N_14028,N_14006);
or U14189 (N_14189,N_14086,N_14122);
or U14190 (N_14190,N_14084,N_14103);
nand U14191 (N_14191,N_14053,N_14026);
nor U14192 (N_14192,N_14092,N_14024);
xnor U14193 (N_14193,N_14019,N_14090);
nand U14194 (N_14194,N_14098,N_14119);
nor U14195 (N_14195,N_14013,N_14090);
xor U14196 (N_14196,N_14049,N_14027);
xnor U14197 (N_14197,N_14030,N_14056);
or U14198 (N_14198,N_14064,N_14005);
and U14199 (N_14199,N_14112,N_14099);
and U14200 (N_14200,N_14064,N_14069);
nand U14201 (N_14201,N_14026,N_14120);
and U14202 (N_14202,N_14076,N_14114);
or U14203 (N_14203,N_14091,N_14010);
nand U14204 (N_14204,N_14041,N_14106);
or U14205 (N_14205,N_14050,N_14013);
xnor U14206 (N_14206,N_14113,N_14111);
or U14207 (N_14207,N_14110,N_14039);
nand U14208 (N_14208,N_14006,N_14067);
xnor U14209 (N_14209,N_14012,N_14056);
nor U14210 (N_14210,N_14004,N_14116);
xor U14211 (N_14211,N_14033,N_14004);
nor U14212 (N_14212,N_14072,N_14062);
nor U14213 (N_14213,N_14052,N_14074);
nand U14214 (N_14214,N_14073,N_14067);
or U14215 (N_14215,N_14116,N_14075);
and U14216 (N_14216,N_14053,N_14105);
or U14217 (N_14217,N_14086,N_14121);
nand U14218 (N_14218,N_14056,N_14028);
or U14219 (N_14219,N_14098,N_14096);
nand U14220 (N_14220,N_14094,N_14099);
nor U14221 (N_14221,N_14086,N_14054);
xor U14222 (N_14222,N_14123,N_14076);
and U14223 (N_14223,N_14029,N_14085);
xor U14224 (N_14224,N_14083,N_14068);
or U14225 (N_14225,N_14033,N_14063);
xor U14226 (N_14226,N_14048,N_14040);
nor U14227 (N_14227,N_14086,N_14057);
nor U14228 (N_14228,N_14092,N_14047);
nor U14229 (N_14229,N_14027,N_14074);
or U14230 (N_14230,N_14020,N_14094);
nor U14231 (N_14231,N_14095,N_14104);
nor U14232 (N_14232,N_14084,N_14123);
nor U14233 (N_14233,N_14117,N_14051);
xnor U14234 (N_14234,N_14077,N_14054);
or U14235 (N_14235,N_14098,N_14045);
nor U14236 (N_14236,N_14081,N_14036);
xnor U14237 (N_14237,N_14048,N_14014);
or U14238 (N_14238,N_14106,N_14056);
or U14239 (N_14239,N_14090,N_14080);
and U14240 (N_14240,N_14032,N_14012);
and U14241 (N_14241,N_14104,N_14072);
nand U14242 (N_14242,N_14011,N_14031);
nor U14243 (N_14243,N_14076,N_14028);
nand U14244 (N_14244,N_14017,N_14001);
nor U14245 (N_14245,N_14094,N_14111);
nor U14246 (N_14246,N_14075,N_14055);
xor U14247 (N_14247,N_14117,N_14067);
or U14248 (N_14248,N_14041,N_14030);
nand U14249 (N_14249,N_14023,N_14069);
and U14250 (N_14250,N_14174,N_14230);
nand U14251 (N_14251,N_14248,N_14238);
or U14252 (N_14252,N_14226,N_14243);
nand U14253 (N_14253,N_14128,N_14214);
or U14254 (N_14254,N_14240,N_14170);
and U14255 (N_14255,N_14146,N_14151);
nor U14256 (N_14256,N_14159,N_14212);
nand U14257 (N_14257,N_14244,N_14184);
xor U14258 (N_14258,N_14162,N_14241);
or U14259 (N_14259,N_14153,N_14150);
nor U14260 (N_14260,N_14233,N_14136);
or U14261 (N_14261,N_14165,N_14224);
or U14262 (N_14262,N_14199,N_14196);
xnor U14263 (N_14263,N_14232,N_14158);
or U14264 (N_14264,N_14206,N_14195);
nand U14265 (N_14265,N_14247,N_14182);
or U14266 (N_14266,N_14176,N_14194);
and U14267 (N_14267,N_14205,N_14155);
nor U14268 (N_14268,N_14183,N_14142);
nand U14269 (N_14269,N_14137,N_14145);
and U14270 (N_14270,N_14148,N_14178);
nand U14271 (N_14271,N_14245,N_14185);
nor U14272 (N_14272,N_14140,N_14229);
nor U14273 (N_14273,N_14220,N_14192);
xor U14274 (N_14274,N_14227,N_14141);
nand U14275 (N_14275,N_14223,N_14197);
xor U14276 (N_14276,N_14237,N_14180);
nor U14277 (N_14277,N_14186,N_14217);
nor U14278 (N_14278,N_14173,N_14181);
or U14279 (N_14279,N_14156,N_14164);
and U14280 (N_14280,N_14131,N_14129);
nand U14281 (N_14281,N_14242,N_14149);
nor U14282 (N_14282,N_14202,N_14135);
xor U14283 (N_14283,N_14166,N_14132);
nor U14284 (N_14284,N_14147,N_14219);
and U14285 (N_14285,N_14216,N_14236);
nor U14286 (N_14286,N_14172,N_14187);
and U14287 (N_14287,N_14163,N_14130);
nand U14288 (N_14288,N_14210,N_14234);
nor U14289 (N_14289,N_14144,N_14138);
or U14290 (N_14290,N_14139,N_14177);
nor U14291 (N_14291,N_14201,N_14239);
nand U14292 (N_14292,N_14249,N_14209);
and U14293 (N_14293,N_14208,N_14157);
or U14294 (N_14294,N_14167,N_14246);
nor U14295 (N_14295,N_14160,N_14168);
xnor U14296 (N_14296,N_14133,N_14127);
nand U14297 (N_14297,N_14134,N_14189);
nand U14298 (N_14298,N_14193,N_14188);
nor U14299 (N_14299,N_14154,N_14213);
or U14300 (N_14300,N_14222,N_14235);
or U14301 (N_14301,N_14218,N_14225);
nand U14302 (N_14302,N_14175,N_14191);
nor U14303 (N_14303,N_14204,N_14231);
nor U14304 (N_14304,N_14126,N_14200);
nor U14305 (N_14305,N_14207,N_14215);
nand U14306 (N_14306,N_14152,N_14198);
or U14307 (N_14307,N_14190,N_14203);
xor U14308 (N_14308,N_14125,N_14211);
nor U14309 (N_14309,N_14143,N_14161);
nor U14310 (N_14310,N_14228,N_14179);
nand U14311 (N_14311,N_14171,N_14169);
nand U14312 (N_14312,N_14221,N_14229);
xor U14313 (N_14313,N_14154,N_14170);
xnor U14314 (N_14314,N_14243,N_14178);
nand U14315 (N_14315,N_14187,N_14132);
nor U14316 (N_14316,N_14201,N_14219);
nor U14317 (N_14317,N_14202,N_14166);
nand U14318 (N_14318,N_14194,N_14215);
or U14319 (N_14319,N_14130,N_14237);
nor U14320 (N_14320,N_14129,N_14127);
nand U14321 (N_14321,N_14154,N_14206);
nor U14322 (N_14322,N_14158,N_14201);
nand U14323 (N_14323,N_14181,N_14168);
xor U14324 (N_14324,N_14239,N_14223);
and U14325 (N_14325,N_14218,N_14148);
and U14326 (N_14326,N_14153,N_14162);
xnor U14327 (N_14327,N_14183,N_14194);
nand U14328 (N_14328,N_14207,N_14158);
xor U14329 (N_14329,N_14135,N_14178);
xnor U14330 (N_14330,N_14127,N_14197);
and U14331 (N_14331,N_14175,N_14208);
nor U14332 (N_14332,N_14203,N_14187);
and U14333 (N_14333,N_14197,N_14218);
or U14334 (N_14334,N_14163,N_14199);
nor U14335 (N_14335,N_14164,N_14217);
nand U14336 (N_14336,N_14137,N_14157);
nor U14337 (N_14337,N_14171,N_14140);
xnor U14338 (N_14338,N_14136,N_14128);
or U14339 (N_14339,N_14242,N_14227);
and U14340 (N_14340,N_14242,N_14130);
and U14341 (N_14341,N_14204,N_14233);
nand U14342 (N_14342,N_14229,N_14193);
nor U14343 (N_14343,N_14153,N_14148);
nand U14344 (N_14344,N_14172,N_14199);
xor U14345 (N_14345,N_14181,N_14207);
and U14346 (N_14346,N_14139,N_14228);
nand U14347 (N_14347,N_14182,N_14160);
xnor U14348 (N_14348,N_14172,N_14185);
and U14349 (N_14349,N_14159,N_14220);
or U14350 (N_14350,N_14219,N_14224);
or U14351 (N_14351,N_14130,N_14183);
nand U14352 (N_14352,N_14201,N_14185);
nand U14353 (N_14353,N_14171,N_14205);
or U14354 (N_14354,N_14198,N_14126);
and U14355 (N_14355,N_14134,N_14168);
nor U14356 (N_14356,N_14175,N_14230);
and U14357 (N_14357,N_14187,N_14222);
and U14358 (N_14358,N_14155,N_14186);
or U14359 (N_14359,N_14233,N_14157);
nand U14360 (N_14360,N_14178,N_14182);
nor U14361 (N_14361,N_14153,N_14177);
xor U14362 (N_14362,N_14216,N_14161);
nand U14363 (N_14363,N_14140,N_14238);
and U14364 (N_14364,N_14182,N_14229);
nor U14365 (N_14365,N_14247,N_14208);
xor U14366 (N_14366,N_14146,N_14228);
and U14367 (N_14367,N_14147,N_14161);
or U14368 (N_14368,N_14243,N_14216);
and U14369 (N_14369,N_14236,N_14196);
or U14370 (N_14370,N_14189,N_14167);
and U14371 (N_14371,N_14244,N_14194);
xor U14372 (N_14372,N_14179,N_14181);
nand U14373 (N_14373,N_14191,N_14202);
and U14374 (N_14374,N_14150,N_14159);
nor U14375 (N_14375,N_14271,N_14329);
and U14376 (N_14376,N_14265,N_14277);
and U14377 (N_14377,N_14258,N_14259);
or U14378 (N_14378,N_14348,N_14337);
or U14379 (N_14379,N_14343,N_14299);
xor U14380 (N_14380,N_14339,N_14285);
and U14381 (N_14381,N_14359,N_14342);
nand U14382 (N_14382,N_14288,N_14296);
or U14383 (N_14383,N_14330,N_14302);
nor U14384 (N_14384,N_14325,N_14282);
nor U14385 (N_14385,N_14318,N_14333);
or U14386 (N_14386,N_14292,N_14312);
xor U14387 (N_14387,N_14355,N_14297);
and U14388 (N_14388,N_14266,N_14341);
and U14389 (N_14389,N_14309,N_14373);
and U14390 (N_14390,N_14362,N_14354);
xor U14391 (N_14391,N_14327,N_14273);
or U14392 (N_14392,N_14251,N_14357);
xnor U14393 (N_14393,N_14284,N_14306);
or U14394 (N_14394,N_14254,N_14372);
or U14395 (N_14395,N_14347,N_14345);
and U14396 (N_14396,N_14334,N_14361);
nor U14397 (N_14397,N_14319,N_14349);
xnor U14398 (N_14398,N_14322,N_14311);
or U14399 (N_14399,N_14304,N_14328);
xor U14400 (N_14400,N_14351,N_14307);
xnor U14401 (N_14401,N_14321,N_14300);
nand U14402 (N_14402,N_14281,N_14367);
and U14403 (N_14403,N_14291,N_14278);
xnor U14404 (N_14404,N_14279,N_14264);
or U14405 (N_14405,N_14286,N_14298);
or U14406 (N_14406,N_14331,N_14350);
nor U14407 (N_14407,N_14314,N_14313);
or U14408 (N_14408,N_14308,N_14272);
nand U14409 (N_14409,N_14310,N_14335);
nor U14410 (N_14410,N_14276,N_14269);
or U14411 (N_14411,N_14316,N_14270);
xnor U14412 (N_14412,N_14369,N_14363);
and U14413 (N_14413,N_14356,N_14290);
and U14414 (N_14414,N_14252,N_14336);
and U14415 (N_14415,N_14368,N_14294);
nand U14416 (N_14416,N_14317,N_14364);
xor U14417 (N_14417,N_14261,N_14257);
xnor U14418 (N_14418,N_14338,N_14326);
and U14419 (N_14419,N_14287,N_14303);
xnor U14420 (N_14420,N_14293,N_14366);
nand U14421 (N_14421,N_14295,N_14256);
or U14422 (N_14422,N_14340,N_14323);
and U14423 (N_14423,N_14268,N_14332);
nor U14424 (N_14424,N_14262,N_14289);
nor U14425 (N_14425,N_14315,N_14253);
nand U14426 (N_14426,N_14371,N_14305);
xnor U14427 (N_14427,N_14301,N_14250);
nand U14428 (N_14428,N_14255,N_14263);
and U14429 (N_14429,N_14275,N_14353);
nand U14430 (N_14430,N_14324,N_14260);
xnor U14431 (N_14431,N_14370,N_14360);
nand U14432 (N_14432,N_14344,N_14358);
nand U14433 (N_14433,N_14283,N_14320);
xnor U14434 (N_14434,N_14374,N_14365);
or U14435 (N_14435,N_14280,N_14352);
and U14436 (N_14436,N_14346,N_14267);
nand U14437 (N_14437,N_14274,N_14311);
nand U14438 (N_14438,N_14311,N_14374);
nand U14439 (N_14439,N_14305,N_14361);
and U14440 (N_14440,N_14315,N_14329);
nand U14441 (N_14441,N_14367,N_14316);
or U14442 (N_14442,N_14362,N_14291);
and U14443 (N_14443,N_14312,N_14343);
nand U14444 (N_14444,N_14326,N_14340);
and U14445 (N_14445,N_14371,N_14337);
xor U14446 (N_14446,N_14349,N_14294);
xor U14447 (N_14447,N_14279,N_14356);
nor U14448 (N_14448,N_14304,N_14347);
and U14449 (N_14449,N_14315,N_14319);
nand U14450 (N_14450,N_14368,N_14371);
nand U14451 (N_14451,N_14334,N_14355);
or U14452 (N_14452,N_14257,N_14313);
xor U14453 (N_14453,N_14329,N_14319);
xnor U14454 (N_14454,N_14270,N_14345);
or U14455 (N_14455,N_14292,N_14281);
nor U14456 (N_14456,N_14279,N_14358);
xor U14457 (N_14457,N_14328,N_14270);
xor U14458 (N_14458,N_14276,N_14282);
xnor U14459 (N_14459,N_14286,N_14363);
xnor U14460 (N_14460,N_14259,N_14335);
xor U14461 (N_14461,N_14350,N_14271);
or U14462 (N_14462,N_14296,N_14370);
nand U14463 (N_14463,N_14335,N_14265);
xnor U14464 (N_14464,N_14290,N_14267);
nand U14465 (N_14465,N_14328,N_14350);
xor U14466 (N_14466,N_14346,N_14374);
xnor U14467 (N_14467,N_14356,N_14251);
nand U14468 (N_14468,N_14323,N_14296);
nor U14469 (N_14469,N_14334,N_14320);
nand U14470 (N_14470,N_14266,N_14329);
and U14471 (N_14471,N_14264,N_14288);
and U14472 (N_14472,N_14344,N_14324);
xor U14473 (N_14473,N_14356,N_14351);
or U14474 (N_14474,N_14320,N_14364);
nand U14475 (N_14475,N_14337,N_14325);
nand U14476 (N_14476,N_14254,N_14360);
and U14477 (N_14477,N_14356,N_14363);
and U14478 (N_14478,N_14270,N_14281);
or U14479 (N_14479,N_14351,N_14318);
or U14480 (N_14480,N_14267,N_14291);
xnor U14481 (N_14481,N_14259,N_14316);
nand U14482 (N_14482,N_14327,N_14323);
xor U14483 (N_14483,N_14352,N_14351);
nand U14484 (N_14484,N_14302,N_14303);
nor U14485 (N_14485,N_14362,N_14353);
nand U14486 (N_14486,N_14310,N_14320);
nor U14487 (N_14487,N_14302,N_14273);
nor U14488 (N_14488,N_14345,N_14326);
nor U14489 (N_14489,N_14271,N_14310);
or U14490 (N_14490,N_14299,N_14342);
nand U14491 (N_14491,N_14285,N_14256);
nand U14492 (N_14492,N_14260,N_14285);
xor U14493 (N_14493,N_14298,N_14260);
nand U14494 (N_14494,N_14263,N_14344);
nand U14495 (N_14495,N_14374,N_14288);
or U14496 (N_14496,N_14366,N_14262);
or U14497 (N_14497,N_14312,N_14368);
or U14498 (N_14498,N_14281,N_14291);
or U14499 (N_14499,N_14349,N_14306);
nor U14500 (N_14500,N_14415,N_14476);
or U14501 (N_14501,N_14488,N_14395);
nor U14502 (N_14502,N_14473,N_14433);
nand U14503 (N_14503,N_14379,N_14424);
and U14504 (N_14504,N_14392,N_14422);
nor U14505 (N_14505,N_14465,N_14450);
xnor U14506 (N_14506,N_14487,N_14405);
nor U14507 (N_14507,N_14404,N_14446);
xnor U14508 (N_14508,N_14377,N_14444);
nor U14509 (N_14509,N_14400,N_14471);
nor U14510 (N_14510,N_14411,N_14397);
xnor U14511 (N_14511,N_14408,N_14469);
or U14512 (N_14512,N_14457,N_14483);
or U14513 (N_14513,N_14445,N_14387);
nor U14514 (N_14514,N_14378,N_14478);
xor U14515 (N_14515,N_14456,N_14416);
nand U14516 (N_14516,N_14419,N_14493);
or U14517 (N_14517,N_14390,N_14420);
xnor U14518 (N_14518,N_14463,N_14462);
or U14519 (N_14519,N_14442,N_14423);
xnor U14520 (N_14520,N_14464,N_14459);
or U14521 (N_14521,N_14418,N_14427);
and U14522 (N_14522,N_14434,N_14421);
or U14523 (N_14523,N_14426,N_14482);
nand U14524 (N_14524,N_14468,N_14432);
nand U14525 (N_14525,N_14443,N_14399);
and U14526 (N_14526,N_14451,N_14428);
nor U14527 (N_14527,N_14477,N_14491);
nor U14528 (N_14528,N_14376,N_14466);
nand U14529 (N_14529,N_14388,N_14438);
nor U14530 (N_14530,N_14449,N_14393);
xor U14531 (N_14531,N_14435,N_14437);
nor U14532 (N_14532,N_14402,N_14474);
xnor U14533 (N_14533,N_14436,N_14475);
or U14534 (N_14534,N_14414,N_14425);
and U14535 (N_14535,N_14441,N_14375);
and U14536 (N_14536,N_14382,N_14412);
nand U14537 (N_14537,N_14458,N_14389);
nand U14538 (N_14538,N_14454,N_14460);
nand U14539 (N_14539,N_14472,N_14467);
xor U14540 (N_14540,N_14479,N_14394);
xnor U14541 (N_14541,N_14492,N_14384);
nand U14542 (N_14542,N_14431,N_14481);
xor U14543 (N_14543,N_14484,N_14499);
and U14544 (N_14544,N_14410,N_14480);
nand U14545 (N_14545,N_14498,N_14406);
and U14546 (N_14546,N_14496,N_14453);
xor U14547 (N_14547,N_14486,N_14430);
nand U14548 (N_14548,N_14495,N_14490);
and U14549 (N_14549,N_14413,N_14391);
xnor U14550 (N_14550,N_14470,N_14461);
nand U14551 (N_14551,N_14396,N_14455);
and U14552 (N_14552,N_14494,N_14386);
xor U14553 (N_14553,N_14448,N_14383);
or U14554 (N_14554,N_14429,N_14485);
nor U14555 (N_14555,N_14489,N_14401);
nor U14556 (N_14556,N_14385,N_14398);
nor U14557 (N_14557,N_14439,N_14407);
xor U14558 (N_14558,N_14447,N_14381);
and U14559 (N_14559,N_14452,N_14417);
and U14560 (N_14560,N_14440,N_14403);
and U14561 (N_14561,N_14409,N_14380);
nor U14562 (N_14562,N_14497,N_14384);
xnor U14563 (N_14563,N_14413,N_14485);
or U14564 (N_14564,N_14442,N_14472);
xor U14565 (N_14565,N_14417,N_14467);
and U14566 (N_14566,N_14412,N_14484);
or U14567 (N_14567,N_14462,N_14427);
nand U14568 (N_14568,N_14422,N_14390);
xor U14569 (N_14569,N_14402,N_14456);
nor U14570 (N_14570,N_14496,N_14414);
or U14571 (N_14571,N_14494,N_14457);
nor U14572 (N_14572,N_14447,N_14424);
nand U14573 (N_14573,N_14409,N_14420);
or U14574 (N_14574,N_14449,N_14471);
xnor U14575 (N_14575,N_14376,N_14444);
nor U14576 (N_14576,N_14381,N_14465);
nor U14577 (N_14577,N_14426,N_14394);
nor U14578 (N_14578,N_14479,N_14462);
nand U14579 (N_14579,N_14403,N_14390);
xnor U14580 (N_14580,N_14382,N_14463);
or U14581 (N_14581,N_14423,N_14393);
nor U14582 (N_14582,N_14422,N_14446);
nor U14583 (N_14583,N_14388,N_14463);
xnor U14584 (N_14584,N_14407,N_14421);
nor U14585 (N_14585,N_14481,N_14485);
and U14586 (N_14586,N_14456,N_14463);
xor U14587 (N_14587,N_14499,N_14403);
nand U14588 (N_14588,N_14476,N_14395);
nor U14589 (N_14589,N_14453,N_14422);
and U14590 (N_14590,N_14471,N_14377);
and U14591 (N_14591,N_14395,N_14443);
or U14592 (N_14592,N_14459,N_14481);
or U14593 (N_14593,N_14397,N_14498);
and U14594 (N_14594,N_14477,N_14469);
nand U14595 (N_14595,N_14464,N_14481);
nor U14596 (N_14596,N_14452,N_14445);
and U14597 (N_14597,N_14437,N_14487);
xor U14598 (N_14598,N_14443,N_14486);
nor U14599 (N_14599,N_14443,N_14465);
and U14600 (N_14600,N_14442,N_14494);
nand U14601 (N_14601,N_14395,N_14461);
nand U14602 (N_14602,N_14408,N_14399);
nor U14603 (N_14603,N_14417,N_14489);
and U14604 (N_14604,N_14430,N_14388);
and U14605 (N_14605,N_14471,N_14452);
xor U14606 (N_14606,N_14400,N_14418);
nand U14607 (N_14607,N_14450,N_14430);
nor U14608 (N_14608,N_14400,N_14444);
nor U14609 (N_14609,N_14393,N_14422);
xor U14610 (N_14610,N_14431,N_14423);
xnor U14611 (N_14611,N_14404,N_14439);
nor U14612 (N_14612,N_14418,N_14447);
and U14613 (N_14613,N_14452,N_14398);
nand U14614 (N_14614,N_14473,N_14396);
nand U14615 (N_14615,N_14418,N_14470);
or U14616 (N_14616,N_14432,N_14379);
or U14617 (N_14617,N_14436,N_14405);
and U14618 (N_14618,N_14447,N_14386);
xnor U14619 (N_14619,N_14433,N_14444);
xor U14620 (N_14620,N_14396,N_14392);
nand U14621 (N_14621,N_14463,N_14428);
nor U14622 (N_14622,N_14419,N_14436);
or U14623 (N_14623,N_14410,N_14464);
nor U14624 (N_14624,N_14439,N_14380);
and U14625 (N_14625,N_14547,N_14617);
xnor U14626 (N_14626,N_14559,N_14557);
xnor U14627 (N_14627,N_14586,N_14618);
nor U14628 (N_14628,N_14579,N_14569);
nor U14629 (N_14629,N_14575,N_14621);
and U14630 (N_14630,N_14515,N_14591);
xor U14631 (N_14631,N_14540,N_14612);
nand U14632 (N_14632,N_14514,N_14572);
xnor U14633 (N_14633,N_14597,N_14526);
nor U14634 (N_14634,N_14513,N_14520);
nand U14635 (N_14635,N_14615,N_14607);
or U14636 (N_14636,N_14545,N_14507);
and U14637 (N_14637,N_14531,N_14553);
nand U14638 (N_14638,N_14523,N_14542);
and U14639 (N_14639,N_14577,N_14604);
xnor U14640 (N_14640,N_14509,N_14528);
xnor U14641 (N_14641,N_14616,N_14587);
xor U14642 (N_14642,N_14598,N_14534);
xnor U14643 (N_14643,N_14593,N_14561);
xnor U14644 (N_14644,N_14530,N_14574);
nor U14645 (N_14645,N_14522,N_14619);
and U14646 (N_14646,N_14580,N_14608);
or U14647 (N_14647,N_14548,N_14599);
nor U14648 (N_14648,N_14573,N_14502);
or U14649 (N_14649,N_14588,N_14584);
nor U14650 (N_14650,N_14589,N_14623);
nand U14651 (N_14651,N_14512,N_14570);
xnor U14652 (N_14652,N_14571,N_14566);
or U14653 (N_14653,N_14602,N_14516);
nor U14654 (N_14654,N_14544,N_14501);
nand U14655 (N_14655,N_14549,N_14565);
nand U14656 (N_14656,N_14535,N_14564);
and U14657 (N_14657,N_14558,N_14556);
nor U14658 (N_14658,N_14620,N_14567);
or U14659 (N_14659,N_14538,N_14562);
xor U14660 (N_14660,N_14560,N_14506);
xor U14661 (N_14661,N_14581,N_14610);
xor U14662 (N_14662,N_14563,N_14536);
nand U14663 (N_14663,N_14552,N_14596);
nand U14664 (N_14664,N_14609,N_14568);
xor U14665 (N_14665,N_14624,N_14511);
nor U14666 (N_14666,N_14576,N_14527);
nor U14667 (N_14667,N_14508,N_14539);
nand U14668 (N_14668,N_14503,N_14537);
xnor U14669 (N_14669,N_14622,N_14505);
nor U14670 (N_14670,N_14605,N_14603);
nand U14671 (N_14671,N_14613,N_14532);
and U14672 (N_14672,N_14500,N_14606);
nor U14673 (N_14673,N_14543,N_14524);
nand U14674 (N_14674,N_14521,N_14529);
or U14675 (N_14675,N_14554,N_14533);
or U14676 (N_14676,N_14546,N_14594);
nand U14677 (N_14677,N_14519,N_14551);
nand U14678 (N_14678,N_14592,N_14583);
xnor U14679 (N_14679,N_14601,N_14611);
or U14680 (N_14680,N_14525,N_14585);
nor U14681 (N_14681,N_14590,N_14510);
or U14682 (N_14682,N_14582,N_14517);
nand U14683 (N_14683,N_14518,N_14600);
xor U14684 (N_14684,N_14541,N_14550);
and U14685 (N_14685,N_14595,N_14614);
xnor U14686 (N_14686,N_14555,N_14578);
xnor U14687 (N_14687,N_14504,N_14596);
nand U14688 (N_14688,N_14524,N_14594);
nor U14689 (N_14689,N_14554,N_14501);
xor U14690 (N_14690,N_14543,N_14603);
or U14691 (N_14691,N_14544,N_14553);
nand U14692 (N_14692,N_14501,N_14579);
nand U14693 (N_14693,N_14617,N_14599);
and U14694 (N_14694,N_14571,N_14530);
xor U14695 (N_14695,N_14542,N_14604);
or U14696 (N_14696,N_14509,N_14558);
nor U14697 (N_14697,N_14585,N_14562);
xor U14698 (N_14698,N_14553,N_14615);
nor U14699 (N_14699,N_14536,N_14507);
nor U14700 (N_14700,N_14529,N_14535);
xnor U14701 (N_14701,N_14619,N_14530);
and U14702 (N_14702,N_14556,N_14579);
nand U14703 (N_14703,N_14582,N_14557);
nor U14704 (N_14704,N_14616,N_14617);
xor U14705 (N_14705,N_14561,N_14540);
nor U14706 (N_14706,N_14523,N_14594);
xnor U14707 (N_14707,N_14584,N_14514);
xnor U14708 (N_14708,N_14602,N_14610);
nor U14709 (N_14709,N_14524,N_14618);
and U14710 (N_14710,N_14572,N_14618);
xor U14711 (N_14711,N_14624,N_14603);
xnor U14712 (N_14712,N_14598,N_14560);
nor U14713 (N_14713,N_14554,N_14603);
nand U14714 (N_14714,N_14518,N_14566);
or U14715 (N_14715,N_14534,N_14606);
and U14716 (N_14716,N_14577,N_14525);
xnor U14717 (N_14717,N_14548,N_14556);
nor U14718 (N_14718,N_14504,N_14562);
xor U14719 (N_14719,N_14573,N_14529);
xnor U14720 (N_14720,N_14622,N_14583);
or U14721 (N_14721,N_14582,N_14550);
and U14722 (N_14722,N_14578,N_14518);
xnor U14723 (N_14723,N_14594,N_14600);
nand U14724 (N_14724,N_14600,N_14602);
xor U14725 (N_14725,N_14609,N_14593);
nor U14726 (N_14726,N_14589,N_14543);
xor U14727 (N_14727,N_14520,N_14507);
nor U14728 (N_14728,N_14598,N_14584);
or U14729 (N_14729,N_14563,N_14531);
nor U14730 (N_14730,N_14559,N_14571);
or U14731 (N_14731,N_14623,N_14567);
and U14732 (N_14732,N_14613,N_14611);
or U14733 (N_14733,N_14509,N_14623);
and U14734 (N_14734,N_14579,N_14568);
nand U14735 (N_14735,N_14584,N_14582);
nand U14736 (N_14736,N_14523,N_14548);
or U14737 (N_14737,N_14574,N_14527);
and U14738 (N_14738,N_14622,N_14538);
nor U14739 (N_14739,N_14551,N_14552);
xor U14740 (N_14740,N_14598,N_14521);
nor U14741 (N_14741,N_14596,N_14580);
and U14742 (N_14742,N_14556,N_14617);
nand U14743 (N_14743,N_14570,N_14546);
or U14744 (N_14744,N_14564,N_14619);
nand U14745 (N_14745,N_14577,N_14523);
and U14746 (N_14746,N_14596,N_14538);
nor U14747 (N_14747,N_14533,N_14517);
xnor U14748 (N_14748,N_14503,N_14514);
and U14749 (N_14749,N_14595,N_14590);
and U14750 (N_14750,N_14702,N_14717);
or U14751 (N_14751,N_14684,N_14666);
nand U14752 (N_14752,N_14732,N_14686);
or U14753 (N_14753,N_14711,N_14748);
nor U14754 (N_14754,N_14650,N_14689);
or U14755 (N_14755,N_14628,N_14642);
xnor U14756 (N_14756,N_14724,N_14649);
nand U14757 (N_14757,N_14742,N_14705);
and U14758 (N_14758,N_14648,N_14658);
nand U14759 (N_14759,N_14638,N_14714);
nor U14760 (N_14760,N_14646,N_14693);
nor U14761 (N_14761,N_14660,N_14716);
or U14762 (N_14762,N_14675,N_14695);
and U14763 (N_14763,N_14677,N_14637);
nor U14764 (N_14764,N_14632,N_14683);
nor U14765 (N_14765,N_14630,N_14657);
nor U14766 (N_14766,N_14696,N_14691);
or U14767 (N_14767,N_14659,N_14640);
nor U14768 (N_14768,N_14727,N_14701);
nor U14769 (N_14769,N_14667,N_14625);
or U14770 (N_14770,N_14633,N_14629);
or U14771 (N_14771,N_14710,N_14698);
nand U14772 (N_14772,N_14745,N_14631);
nand U14773 (N_14773,N_14739,N_14671);
nor U14774 (N_14774,N_14713,N_14738);
nor U14775 (N_14775,N_14743,N_14703);
xnor U14776 (N_14776,N_14740,N_14749);
and U14777 (N_14777,N_14654,N_14627);
nor U14778 (N_14778,N_14662,N_14651);
nor U14779 (N_14779,N_14643,N_14719);
and U14780 (N_14780,N_14685,N_14687);
and U14781 (N_14781,N_14694,N_14700);
nand U14782 (N_14782,N_14668,N_14699);
and U14783 (N_14783,N_14726,N_14652);
xnor U14784 (N_14784,N_14725,N_14679);
and U14785 (N_14785,N_14663,N_14718);
or U14786 (N_14786,N_14731,N_14733);
nand U14787 (N_14787,N_14635,N_14708);
nand U14788 (N_14788,N_14665,N_14680);
nor U14789 (N_14789,N_14639,N_14741);
or U14790 (N_14790,N_14709,N_14747);
xor U14791 (N_14791,N_14673,N_14676);
xor U14792 (N_14792,N_14653,N_14720);
nand U14793 (N_14793,N_14730,N_14661);
nor U14794 (N_14794,N_14655,N_14674);
nor U14795 (N_14795,N_14670,N_14644);
or U14796 (N_14796,N_14647,N_14634);
or U14797 (N_14797,N_14746,N_14737);
and U14798 (N_14798,N_14681,N_14734);
or U14799 (N_14799,N_14626,N_14682);
and U14800 (N_14800,N_14736,N_14669);
nor U14801 (N_14801,N_14641,N_14645);
or U14802 (N_14802,N_14688,N_14722);
nor U14803 (N_14803,N_14690,N_14672);
xor U14804 (N_14804,N_14721,N_14664);
nor U14805 (N_14805,N_14656,N_14707);
nor U14806 (N_14806,N_14704,N_14723);
or U14807 (N_14807,N_14729,N_14712);
nor U14808 (N_14808,N_14735,N_14744);
xnor U14809 (N_14809,N_14715,N_14678);
nand U14810 (N_14810,N_14706,N_14636);
xnor U14811 (N_14811,N_14692,N_14728);
or U14812 (N_14812,N_14697,N_14627);
xnor U14813 (N_14813,N_14696,N_14665);
or U14814 (N_14814,N_14640,N_14646);
and U14815 (N_14815,N_14627,N_14725);
nand U14816 (N_14816,N_14693,N_14627);
xnor U14817 (N_14817,N_14654,N_14673);
or U14818 (N_14818,N_14687,N_14700);
nor U14819 (N_14819,N_14651,N_14721);
xnor U14820 (N_14820,N_14666,N_14707);
or U14821 (N_14821,N_14737,N_14658);
nor U14822 (N_14822,N_14687,N_14691);
nand U14823 (N_14823,N_14740,N_14723);
nand U14824 (N_14824,N_14732,N_14674);
or U14825 (N_14825,N_14684,N_14733);
and U14826 (N_14826,N_14648,N_14731);
nor U14827 (N_14827,N_14675,N_14688);
and U14828 (N_14828,N_14731,N_14674);
nand U14829 (N_14829,N_14669,N_14677);
and U14830 (N_14830,N_14703,N_14669);
nand U14831 (N_14831,N_14651,N_14732);
or U14832 (N_14832,N_14625,N_14645);
nor U14833 (N_14833,N_14710,N_14700);
nor U14834 (N_14834,N_14701,N_14704);
xnor U14835 (N_14835,N_14706,N_14645);
nand U14836 (N_14836,N_14719,N_14627);
and U14837 (N_14837,N_14638,N_14641);
or U14838 (N_14838,N_14633,N_14694);
nor U14839 (N_14839,N_14657,N_14643);
xor U14840 (N_14840,N_14712,N_14644);
nand U14841 (N_14841,N_14748,N_14713);
nor U14842 (N_14842,N_14662,N_14704);
xor U14843 (N_14843,N_14705,N_14714);
and U14844 (N_14844,N_14735,N_14687);
and U14845 (N_14845,N_14654,N_14699);
xor U14846 (N_14846,N_14677,N_14655);
nor U14847 (N_14847,N_14686,N_14733);
or U14848 (N_14848,N_14629,N_14665);
nor U14849 (N_14849,N_14673,N_14749);
nand U14850 (N_14850,N_14699,N_14650);
or U14851 (N_14851,N_14726,N_14632);
xnor U14852 (N_14852,N_14666,N_14636);
nor U14853 (N_14853,N_14746,N_14664);
or U14854 (N_14854,N_14691,N_14672);
or U14855 (N_14855,N_14634,N_14720);
or U14856 (N_14856,N_14686,N_14673);
nor U14857 (N_14857,N_14739,N_14696);
nor U14858 (N_14858,N_14747,N_14746);
nand U14859 (N_14859,N_14708,N_14625);
nand U14860 (N_14860,N_14705,N_14690);
and U14861 (N_14861,N_14652,N_14633);
or U14862 (N_14862,N_14705,N_14702);
nor U14863 (N_14863,N_14648,N_14692);
xnor U14864 (N_14864,N_14639,N_14686);
and U14865 (N_14865,N_14723,N_14674);
and U14866 (N_14866,N_14744,N_14648);
nand U14867 (N_14867,N_14678,N_14683);
or U14868 (N_14868,N_14741,N_14654);
nor U14869 (N_14869,N_14646,N_14723);
nand U14870 (N_14870,N_14677,N_14727);
and U14871 (N_14871,N_14701,N_14638);
nand U14872 (N_14872,N_14725,N_14719);
nand U14873 (N_14873,N_14686,N_14625);
and U14874 (N_14874,N_14627,N_14712);
nand U14875 (N_14875,N_14760,N_14841);
nand U14876 (N_14876,N_14790,N_14851);
nor U14877 (N_14877,N_14858,N_14798);
nand U14878 (N_14878,N_14839,N_14865);
and U14879 (N_14879,N_14804,N_14848);
or U14880 (N_14880,N_14807,N_14812);
xnor U14881 (N_14881,N_14786,N_14873);
nor U14882 (N_14882,N_14764,N_14817);
nor U14883 (N_14883,N_14831,N_14816);
or U14884 (N_14884,N_14846,N_14830);
nand U14885 (N_14885,N_14833,N_14776);
nor U14886 (N_14886,N_14832,N_14778);
nand U14887 (N_14887,N_14787,N_14752);
or U14888 (N_14888,N_14780,N_14769);
nor U14889 (N_14889,N_14801,N_14829);
xor U14890 (N_14890,N_14824,N_14826);
nor U14891 (N_14891,N_14802,N_14783);
xnor U14892 (N_14892,N_14836,N_14766);
xnor U14893 (N_14893,N_14754,N_14794);
xnor U14894 (N_14894,N_14770,N_14753);
nor U14895 (N_14895,N_14762,N_14862);
xor U14896 (N_14896,N_14768,N_14757);
nor U14897 (N_14897,N_14869,N_14874);
nor U14898 (N_14898,N_14795,N_14845);
and U14899 (N_14899,N_14864,N_14843);
and U14900 (N_14900,N_14792,N_14784);
nor U14901 (N_14901,N_14793,N_14796);
or U14902 (N_14902,N_14810,N_14823);
xnor U14903 (N_14903,N_14813,N_14808);
nand U14904 (N_14904,N_14763,N_14868);
nand U14905 (N_14905,N_14853,N_14771);
nand U14906 (N_14906,N_14756,N_14765);
or U14907 (N_14907,N_14799,N_14838);
nor U14908 (N_14908,N_14785,N_14872);
nor U14909 (N_14909,N_14779,N_14791);
xor U14910 (N_14910,N_14803,N_14759);
xnor U14911 (N_14911,N_14844,N_14772);
nor U14912 (N_14912,N_14750,N_14777);
nor U14913 (N_14913,N_14840,N_14758);
and U14914 (N_14914,N_14834,N_14855);
nand U14915 (N_14915,N_14820,N_14861);
or U14916 (N_14916,N_14818,N_14870);
and U14917 (N_14917,N_14774,N_14854);
nor U14918 (N_14918,N_14827,N_14856);
nand U14919 (N_14919,N_14809,N_14837);
and U14920 (N_14920,N_14852,N_14867);
or U14921 (N_14921,N_14773,N_14849);
nand U14922 (N_14922,N_14761,N_14767);
or U14923 (N_14923,N_14805,N_14814);
and U14924 (N_14924,N_14789,N_14782);
nand U14925 (N_14925,N_14815,N_14825);
nand U14926 (N_14926,N_14871,N_14828);
and U14927 (N_14927,N_14751,N_14797);
nor U14928 (N_14928,N_14857,N_14811);
and U14929 (N_14929,N_14775,N_14819);
and U14930 (N_14930,N_14788,N_14866);
nor U14931 (N_14931,N_14842,N_14755);
xnor U14932 (N_14932,N_14859,N_14822);
and U14933 (N_14933,N_14821,N_14781);
and U14934 (N_14934,N_14800,N_14835);
nor U14935 (N_14935,N_14863,N_14850);
nand U14936 (N_14936,N_14806,N_14860);
xnor U14937 (N_14937,N_14847,N_14766);
or U14938 (N_14938,N_14795,N_14874);
nor U14939 (N_14939,N_14864,N_14828);
nand U14940 (N_14940,N_14787,N_14852);
and U14941 (N_14941,N_14857,N_14769);
and U14942 (N_14942,N_14820,N_14809);
and U14943 (N_14943,N_14863,N_14843);
xor U14944 (N_14944,N_14855,N_14757);
and U14945 (N_14945,N_14834,N_14873);
nand U14946 (N_14946,N_14782,N_14760);
nor U14947 (N_14947,N_14759,N_14833);
nor U14948 (N_14948,N_14760,N_14865);
and U14949 (N_14949,N_14816,N_14857);
xnor U14950 (N_14950,N_14835,N_14784);
nand U14951 (N_14951,N_14802,N_14780);
xnor U14952 (N_14952,N_14803,N_14808);
nor U14953 (N_14953,N_14828,N_14862);
nor U14954 (N_14954,N_14808,N_14752);
or U14955 (N_14955,N_14758,N_14762);
xnor U14956 (N_14956,N_14781,N_14812);
nor U14957 (N_14957,N_14862,N_14756);
nand U14958 (N_14958,N_14834,N_14787);
xnor U14959 (N_14959,N_14856,N_14782);
nand U14960 (N_14960,N_14815,N_14865);
nor U14961 (N_14961,N_14768,N_14856);
nand U14962 (N_14962,N_14855,N_14818);
nand U14963 (N_14963,N_14865,N_14776);
and U14964 (N_14964,N_14814,N_14757);
or U14965 (N_14965,N_14865,N_14805);
xnor U14966 (N_14966,N_14812,N_14831);
xor U14967 (N_14967,N_14848,N_14780);
xnor U14968 (N_14968,N_14833,N_14794);
and U14969 (N_14969,N_14816,N_14751);
nor U14970 (N_14970,N_14807,N_14762);
nand U14971 (N_14971,N_14766,N_14860);
nor U14972 (N_14972,N_14851,N_14772);
or U14973 (N_14973,N_14800,N_14868);
xnor U14974 (N_14974,N_14805,N_14843);
nand U14975 (N_14975,N_14757,N_14862);
and U14976 (N_14976,N_14777,N_14859);
or U14977 (N_14977,N_14793,N_14862);
xor U14978 (N_14978,N_14874,N_14790);
xor U14979 (N_14979,N_14810,N_14872);
and U14980 (N_14980,N_14763,N_14768);
nand U14981 (N_14981,N_14764,N_14812);
xor U14982 (N_14982,N_14824,N_14774);
nor U14983 (N_14983,N_14815,N_14778);
xnor U14984 (N_14984,N_14804,N_14809);
nand U14985 (N_14985,N_14861,N_14805);
nand U14986 (N_14986,N_14857,N_14852);
and U14987 (N_14987,N_14874,N_14755);
or U14988 (N_14988,N_14859,N_14759);
or U14989 (N_14989,N_14814,N_14777);
nand U14990 (N_14990,N_14767,N_14824);
xor U14991 (N_14991,N_14753,N_14845);
nand U14992 (N_14992,N_14804,N_14871);
nand U14993 (N_14993,N_14845,N_14844);
or U14994 (N_14994,N_14835,N_14778);
nor U14995 (N_14995,N_14874,N_14791);
nor U14996 (N_14996,N_14826,N_14778);
nand U14997 (N_14997,N_14765,N_14855);
nor U14998 (N_14998,N_14759,N_14812);
nor U14999 (N_14999,N_14806,N_14827);
or UO_0 (O_0,N_14981,N_14938);
or UO_1 (O_1,N_14924,N_14950);
nor UO_2 (O_2,N_14906,N_14921);
nor UO_3 (O_3,N_14915,N_14957);
and UO_4 (O_4,N_14912,N_14956);
xor UO_5 (O_5,N_14911,N_14998);
or UO_6 (O_6,N_14885,N_14952);
and UO_7 (O_7,N_14988,N_14945);
xor UO_8 (O_8,N_14989,N_14995);
xnor UO_9 (O_9,N_14959,N_14919);
nor UO_10 (O_10,N_14933,N_14970);
nor UO_11 (O_11,N_14909,N_14999);
or UO_12 (O_12,N_14910,N_14897);
or UO_13 (O_13,N_14886,N_14980);
and UO_14 (O_14,N_14918,N_14893);
nand UO_15 (O_15,N_14943,N_14967);
and UO_16 (O_16,N_14946,N_14899);
xnor UO_17 (O_17,N_14913,N_14979);
xor UO_18 (O_18,N_14890,N_14907);
nand UO_19 (O_19,N_14982,N_14947);
or UO_20 (O_20,N_14985,N_14925);
xnor UO_21 (O_21,N_14958,N_14937);
or UO_22 (O_22,N_14978,N_14972);
nor UO_23 (O_23,N_14941,N_14926);
nor UO_24 (O_24,N_14997,N_14992);
xor UO_25 (O_25,N_14881,N_14954);
nor UO_26 (O_26,N_14887,N_14935);
nor UO_27 (O_27,N_14904,N_14892);
nor UO_28 (O_28,N_14944,N_14951);
and UO_29 (O_29,N_14964,N_14932);
nor UO_30 (O_30,N_14973,N_14891);
nor UO_31 (O_31,N_14974,N_14960);
and UO_32 (O_32,N_14898,N_14963);
xnor UO_33 (O_33,N_14968,N_14971);
nand UO_34 (O_34,N_14990,N_14940);
xnor UO_35 (O_35,N_14936,N_14894);
nor UO_36 (O_36,N_14961,N_14888);
or UO_37 (O_37,N_14942,N_14994);
and UO_38 (O_38,N_14880,N_14934);
nor UO_39 (O_39,N_14903,N_14983);
nand UO_40 (O_40,N_14975,N_14902);
and UO_41 (O_41,N_14949,N_14879);
or UO_42 (O_42,N_14931,N_14889);
nand UO_43 (O_43,N_14991,N_14883);
xor UO_44 (O_44,N_14905,N_14920);
and UO_45 (O_45,N_14928,N_14987);
nor UO_46 (O_46,N_14884,N_14895);
and UO_47 (O_47,N_14900,N_14986);
xnor UO_48 (O_48,N_14878,N_14929);
nor UO_49 (O_49,N_14976,N_14996);
xnor UO_50 (O_50,N_14916,N_14962);
nor UO_51 (O_51,N_14927,N_14955);
nand UO_52 (O_52,N_14877,N_14993);
and UO_53 (O_53,N_14917,N_14977);
nand UO_54 (O_54,N_14922,N_14875);
nand UO_55 (O_55,N_14965,N_14930);
nand UO_56 (O_56,N_14939,N_14984);
nor UO_57 (O_57,N_14901,N_14896);
nor UO_58 (O_58,N_14923,N_14948);
nor UO_59 (O_59,N_14876,N_14882);
xnor UO_60 (O_60,N_14966,N_14969);
nor UO_61 (O_61,N_14953,N_14908);
xor UO_62 (O_62,N_14914,N_14896);
nor UO_63 (O_63,N_14938,N_14893);
nand UO_64 (O_64,N_14934,N_14899);
nand UO_65 (O_65,N_14977,N_14960);
nor UO_66 (O_66,N_14911,N_14947);
or UO_67 (O_67,N_14937,N_14936);
xnor UO_68 (O_68,N_14966,N_14894);
nand UO_69 (O_69,N_14930,N_14988);
xnor UO_70 (O_70,N_14916,N_14993);
or UO_71 (O_71,N_14946,N_14965);
nand UO_72 (O_72,N_14992,N_14918);
xor UO_73 (O_73,N_14964,N_14897);
and UO_74 (O_74,N_14984,N_14970);
and UO_75 (O_75,N_14947,N_14890);
nand UO_76 (O_76,N_14900,N_14917);
or UO_77 (O_77,N_14936,N_14963);
or UO_78 (O_78,N_14876,N_14999);
nor UO_79 (O_79,N_14878,N_14951);
xnor UO_80 (O_80,N_14963,N_14911);
and UO_81 (O_81,N_14937,N_14883);
or UO_82 (O_82,N_14950,N_14969);
nor UO_83 (O_83,N_14929,N_14981);
and UO_84 (O_84,N_14896,N_14903);
or UO_85 (O_85,N_14937,N_14998);
nor UO_86 (O_86,N_14995,N_14949);
and UO_87 (O_87,N_14950,N_14889);
nand UO_88 (O_88,N_14905,N_14988);
xor UO_89 (O_89,N_14944,N_14912);
nor UO_90 (O_90,N_14998,N_14927);
and UO_91 (O_91,N_14908,N_14904);
xnor UO_92 (O_92,N_14934,N_14912);
nor UO_93 (O_93,N_14884,N_14917);
nor UO_94 (O_94,N_14894,N_14920);
nand UO_95 (O_95,N_14956,N_14957);
nor UO_96 (O_96,N_14893,N_14923);
and UO_97 (O_97,N_14882,N_14885);
xnor UO_98 (O_98,N_14948,N_14920);
xnor UO_99 (O_99,N_14955,N_14916);
or UO_100 (O_100,N_14946,N_14893);
nor UO_101 (O_101,N_14967,N_14983);
nor UO_102 (O_102,N_14989,N_14935);
or UO_103 (O_103,N_14902,N_14878);
xor UO_104 (O_104,N_14931,N_14994);
nand UO_105 (O_105,N_14924,N_14961);
or UO_106 (O_106,N_14877,N_14918);
or UO_107 (O_107,N_14936,N_14931);
and UO_108 (O_108,N_14951,N_14954);
xnor UO_109 (O_109,N_14962,N_14895);
nor UO_110 (O_110,N_14957,N_14959);
and UO_111 (O_111,N_14921,N_14968);
and UO_112 (O_112,N_14894,N_14922);
or UO_113 (O_113,N_14984,N_14978);
and UO_114 (O_114,N_14946,N_14961);
nand UO_115 (O_115,N_14886,N_14932);
xnor UO_116 (O_116,N_14953,N_14951);
and UO_117 (O_117,N_14927,N_14952);
and UO_118 (O_118,N_14906,N_14875);
xnor UO_119 (O_119,N_14956,N_14892);
nand UO_120 (O_120,N_14972,N_14914);
nor UO_121 (O_121,N_14956,N_14896);
nor UO_122 (O_122,N_14961,N_14911);
or UO_123 (O_123,N_14876,N_14997);
xor UO_124 (O_124,N_14992,N_14977);
nor UO_125 (O_125,N_14916,N_14958);
xnor UO_126 (O_126,N_14978,N_14927);
or UO_127 (O_127,N_14963,N_14950);
nor UO_128 (O_128,N_14893,N_14877);
nor UO_129 (O_129,N_14972,N_14876);
or UO_130 (O_130,N_14953,N_14956);
and UO_131 (O_131,N_14986,N_14886);
nor UO_132 (O_132,N_14897,N_14913);
and UO_133 (O_133,N_14921,N_14945);
nor UO_134 (O_134,N_14876,N_14881);
xnor UO_135 (O_135,N_14980,N_14888);
and UO_136 (O_136,N_14968,N_14989);
or UO_137 (O_137,N_14946,N_14968);
xor UO_138 (O_138,N_14925,N_14926);
nand UO_139 (O_139,N_14973,N_14980);
or UO_140 (O_140,N_14915,N_14896);
nand UO_141 (O_141,N_14929,N_14980);
xnor UO_142 (O_142,N_14969,N_14912);
nand UO_143 (O_143,N_14930,N_14985);
nand UO_144 (O_144,N_14953,N_14875);
nand UO_145 (O_145,N_14966,N_14937);
or UO_146 (O_146,N_14991,N_14919);
xor UO_147 (O_147,N_14960,N_14950);
nor UO_148 (O_148,N_14990,N_14978);
or UO_149 (O_149,N_14968,N_14904);
and UO_150 (O_150,N_14934,N_14996);
and UO_151 (O_151,N_14933,N_14983);
xor UO_152 (O_152,N_14995,N_14925);
nor UO_153 (O_153,N_14943,N_14979);
xor UO_154 (O_154,N_14940,N_14930);
nor UO_155 (O_155,N_14890,N_14975);
xnor UO_156 (O_156,N_14924,N_14963);
xor UO_157 (O_157,N_14905,N_14895);
or UO_158 (O_158,N_14898,N_14887);
and UO_159 (O_159,N_14918,N_14930);
nand UO_160 (O_160,N_14929,N_14918);
nor UO_161 (O_161,N_14997,N_14890);
xor UO_162 (O_162,N_14978,N_14959);
nor UO_163 (O_163,N_14954,N_14941);
and UO_164 (O_164,N_14958,N_14880);
and UO_165 (O_165,N_14940,N_14882);
nand UO_166 (O_166,N_14964,N_14976);
xor UO_167 (O_167,N_14990,N_14904);
nand UO_168 (O_168,N_14974,N_14923);
nand UO_169 (O_169,N_14981,N_14895);
and UO_170 (O_170,N_14885,N_14995);
or UO_171 (O_171,N_14888,N_14933);
xnor UO_172 (O_172,N_14999,N_14976);
and UO_173 (O_173,N_14907,N_14966);
and UO_174 (O_174,N_14894,N_14892);
and UO_175 (O_175,N_14888,N_14899);
and UO_176 (O_176,N_14911,N_14877);
and UO_177 (O_177,N_14877,N_14948);
nor UO_178 (O_178,N_14984,N_14944);
nor UO_179 (O_179,N_14969,N_14952);
nand UO_180 (O_180,N_14980,N_14971);
nor UO_181 (O_181,N_14944,N_14913);
nor UO_182 (O_182,N_14882,N_14884);
nand UO_183 (O_183,N_14913,N_14989);
nor UO_184 (O_184,N_14980,N_14988);
or UO_185 (O_185,N_14965,N_14973);
or UO_186 (O_186,N_14970,N_14969);
xor UO_187 (O_187,N_14932,N_14893);
xor UO_188 (O_188,N_14885,N_14943);
nor UO_189 (O_189,N_14939,N_14876);
nor UO_190 (O_190,N_14917,N_14995);
and UO_191 (O_191,N_14911,N_14996);
nand UO_192 (O_192,N_14900,N_14993);
nand UO_193 (O_193,N_14925,N_14942);
nand UO_194 (O_194,N_14880,N_14931);
xnor UO_195 (O_195,N_14943,N_14953);
or UO_196 (O_196,N_14910,N_14919);
or UO_197 (O_197,N_14913,N_14990);
nor UO_198 (O_198,N_14937,N_14953);
nor UO_199 (O_199,N_14970,N_14875);
and UO_200 (O_200,N_14926,N_14983);
nor UO_201 (O_201,N_14937,N_14990);
or UO_202 (O_202,N_14991,N_14992);
or UO_203 (O_203,N_14943,N_14968);
or UO_204 (O_204,N_14981,N_14884);
xor UO_205 (O_205,N_14962,N_14884);
xor UO_206 (O_206,N_14924,N_14959);
and UO_207 (O_207,N_14947,N_14943);
and UO_208 (O_208,N_14929,N_14922);
or UO_209 (O_209,N_14899,N_14919);
and UO_210 (O_210,N_14969,N_14913);
xnor UO_211 (O_211,N_14894,N_14918);
nand UO_212 (O_212,N_14917,N_14935);
nor UO_213 (O_213,N_14914,N_14938);
nand UO_214 (O_214,N_14931,N_14912);
nand UO_215 (O_215,N_14912,N_14973);
and UO_216 (O_216,N_14912,N_14953);
and UO_217 (O_217,N_14936,N_14960);
nand UO_218 (O_218,N_14912,N_14976);
nor UO_219 (O_219,N_14976,N_14887);
nor UO_220 (O_220,N_14965,N_14949);
or UO_221 (O_221,N_14931,N_14916);
or UO_222 (O_222,N_14908,N_14999);
xor UO_223 (O_223,N_14919,N_14900);
or UO_224 (O_224,N_14957,N_14944);
nand UO_225 (O_225,N_14957,N_14898);
nor UO_226 (O_226,N_14898,N_14913);
nor UO_227 (O_227,N_14946,N_14973);
and UO_228 (O_228,N_14909,N_14924);
or UO_229 (O_229,N_14948,N_14937);
nor UO_230 (O_230,N_14951,N_14897);
nand UO_231 (O_231,N_14918,N_14898);
or UO_232 (O_232,N_14990,N_14991);
nor UO_233 (O_233,N_14956,N_14916);
xnor UO_234 (O_234,N_14968,N_14956);
and UO_235 (O_235,N_14999,N_14933);
or UO_236 (O_236,N_14932,N_14957);
xor UO_237 (O_237,N_14962,N_14908);
nor UO_238 (O_238,N_14943,N_14994);
and UO_239 (O_239,N_14947,N_14992);
or UO_240 (O_240,N_14930,N_14891);
and UO_241 (O_241,N_14924,N_14897);
nand UO_242 (O_242,N_14958,N_14974);
or UO_243 (O_243,N_14917,N_14999);
nor UO_244 (O_244,N_14928,N_14993);
or UO_245 (O_245,N_14982,N_14924);
and UO_246 (O_246,N_14985,N_14889);
nor UO_247 (O_247,N_14967,N_14903);
xnor UO_248 (O_248,N_14909,N_14974);
nand UO_249 (O_249,N_14880,N_14904);
and UO_250 (O_250,N_14886,N_14888);
nor UO_251 (O_251,N_14993,N_14949);
nand UO_252 (O_252,N_14980,N_14909);
nor UO_253 (O_253,N_14938,N_14909);
or UO_254 (O_254,N_14987,N_14908);
nand UO_255 (O_255,N_14882,N_14936);
and UO_256 (O_256,N_14934,N_14928);
or UO_257 (O_257,N_14990,N_14910);
and UO_258 (O_258,N_14883,N_14955);
or UO_259 (O_259,N_14918,N_14952);
xor UO_260 (O_260,N_14904,N_14916);
and UO_261 (O_261,N_14961,N_14992);
or UO_262 (O_262,N_14884,N_14989);
nor UO_263 (O_263,N_14893,N_14896);
xor UO_264 (O_264,N_14958,N_14987);
nor UO_265 (O_265,N_14929,N_14966);
and UO_266 (O_266,N_14876,N_14945);
or UO_267 (O_267,N_14930,N_14916);
xnor UO_268 (O_268,N_14958,N_14934);
and UO_269 (O_269,N_14929,N_14964);
nand UO_270 (O_270,N_14875,N_14932);
nand UO_271 (O_271,N_14951,N_14903);
nand UO_272 (O_272,N_14981,N_14910);
or UO_273 (O_273,N_14969,N_14933);
nand UO_274 (O_274,N_14908,N_14966);
and UO_275 (O_275,N_14936,N_14997);
nor UO_276 (O_276,N_14973,N_14987);
or UO_277 (O_277,N_14962,N_14931);
and UO_278 (O_278,N_14949,N_14962);
nor UO_279 (O_279,N_14967,N_14971);
nor UO_280 (O_280,N_14951,N_14899);
and UO_281 (O_281,N_14979,N_14984);
and UO_282 (O_282,N_14953,N_14892);
and UO_283 (O_283,N_14997,N_14891);
nor UO_284 (O_284,N_14920,N_14972);
or UO_285 (O_285,N_14904,N_14944);
and UO_286 (O_286,N_14967,N_14946);
and UO_287 (O_287,N_14925,N_14928);
or UO_288 (O_288,N_14942,N_14951);
or UO_289 (O_289,N_14965,N_14877);
nor UO_290 (O_290,N_14974,N_14954);
nand UO_291 (O_291,N_14916,N_14889);
or UO_292 (O_292,N_14976,N_14963);
nand UO_293 (O_293,N_14901,N_14978);
xnor UO_294 (O_294,N_14954,N_14982);
xnor UO_295 (O_295,N_14895,N_14972);
nand UO_296 (O_296,N_14926,N_14875);
and UO_297 (O_297,N_14875,N_14931);
nand UO_298 (O_298,N_14963,N_14964);
xor UO_299 (O_299,N_14980,N_14950);
or UO_300 (O_300,N_14884,N_14885);
nor UO_301 (O_301,N_14882,N_14901);
nand UO_302 (O_302,N_14918,N_14885);
or UO_303 (O_303,N_14972,N_14892);
xor UO_304 (O_304,N_14996,N_14927);
nor UO_305 (O_305,N_14919,N_14984);
xor UO_306 (O_306,N_14915,N_14911);
nor UO_307 (O_307,N_14980,N_14995);
xor UO_308 (O_308,N_14948,N_14890);
nor UO_309 (O_309,N_14956,N_14911);
and UO_310 (O_310,N_14883,N_14924);
nand UO_311 (O_311,N_14908,N_14887);
and UO_312 (O_312,N_14882,N_14893);
and UO_313 (O_313,N_14877,N_14954);
nor UO_314 (O_314,N_14992,N_14913);
or UO_315 (O_315,N_14887,N_14890);
or UO_316 (O_316,N_14884,N_14933);
nor UO_317 (O_317,N_14918,N_14919);
and UO_318 (O_318,N_14984,N_14967);
nand UO_319 (O_319,N_14935,N_14970);
xor UO_320 (O_320,N_14930,N_14968);
nor UO_321 (O_321,N_14935,N_14877);
nor UO_322 (O_322,N_14945,N_14966);
nor UO_323 (O_323,N_14925,N_14915);
or UO_324 (O_324,N_14945,N_14973);
nand UO_325 (O_325,N_14988,N_14972);
xnor UO_326 (O_326,N_14896,N_14886);
nand UO_327 (O_327,N_14929,N_14880);
and UO_328 (O_328,N_14991,N_14972);
nand UO_329 (O_329,N_14878,N_14906);
and UO_330 (O_330,N_14913,N_14882);
nand UO_331 (O_331,N_14996,N_14951);
nor UO_332 (O_332,N_14954,N_14880);
or UO_333 (O_333,N_14974,N_14961);
nand UO_334 (O_334,N_14927,N_14907);
and UO_335 (O_335,N_14979,N_14892);
nand UO_336 (O_336,N_14912,N_14933);
nand UO_337 (O_337,N_14898,N_14921);
and UO_338 (O_338,N_14926,N_14956);
xnor UO_339 (O_339,N_14893,N_14953);
and UO_340 (O_340,N_14994,N_14982);
xor UO_341 (O_341,N_14938,N_14903);
xor UO_342 (O_342,N_14988,N_14912);
nand UO_343 (O_343,N_14894,N_14990);
nand UO_344 (O_344,N_14879,N_14936);
xor UO_345 (O_345,N_14999,N_14955);
nand UO_346 (O_346,N_14915,N_14967);
and UO_347 (O_347,N_14993,N_14878);
nor UO_348 (O_348,N_14962,N_14889);
xnor UO_349 (O_349,N_14888,N_14963);
nor UO_350 (O_350,N_14914,N_14994);
nor UO_351 (O_351,N_14987,N_14945);
nor UO_352 (O_352,N_14897,N_14909);
and UO_353 (O_353,N_14985,N_14950);
and UO_354 (O_354,N_14929,N_14904);
nand UO_355 (O_355,N_14876,N_14913);
nand UO_356 (O_356,N_14950,N_14964);
nor UO_357 (O_357,N_14952,N_14938);
nor UO_358 (O_358,N_14955,N_14972);
xor UO_359 (O_359,N_14921,N_14998);
nor UO_360 (O_360,N_14989,N_14955);
nor UO_361 (O_361,N_14895,N_14971);
or UO_362 (O_362,N_14920,N_14963);
and UO_363 (O_363,N_14895,N_14903);
nand UO_364 (O_364,N_14979,N_14906);
nor UO_365 (O_365,N_14932,N_14905);
and UO_366 (O_366,N_14972,N_14968);
or UO_367 (O_367,N_14945,N_14908);
or UO_368 (O_368,N_14875,N_14983);
nor UO_369 (O_369,N_14877,N_14921);
nor UO_370 (O_370,N_14920,N_14994);
nand UO_371 (O_371,N_14899,N_14909);
nand UO_372 (O_372,N_14898,N_14933);
nor UO_373 (O_373,N_14901,N_14956);
and UO_374 (O_374,N_14964,N_14945);
or UO_375 (O_375,N_14959,N_14918);
nand UO_376 (O_376,N_14879,N_14944);
nand UO_377 (O_377,N_14989,N_14883);
and UO_378 (O_378,N_14946,N_14966);
and UO_379 (O_379,N_14961,N_14994);
nand UO_380 (O_380,N_14971,N_14928);
xor UO_381 (O_381,N_14997,N_14951);
nand UO_382 (O_382,N_14923,N_14993);
nand UO_383 (O_383,N_14943,N_14955);
nand UO_384 (O_384,N_14937,N_14967);
nor UO_385 (O_385,N_14923,N_14937);
xor UO_386 (O_386,N_14944,N_14910);
nor UO_387 (O_387,N_14934,N_14889);
or UO_388 (O_388,N_14969,N_14987);
and UO_389 (O_389,N_14914,N_14901);
or UO_390 (O_390,N_14898,N_14952);
nor UO_391 (O_391,N_14936,N_14928);
xor UO_392 (O_392,N_14909,N_14908);
nand UO_393 (O_393,N_14992,N_14984);
nor UO_394 (O_394,N_14914,N_14886);
or UO_395 (O_395,N_14990,N_14966);
xnor UO_396 (O_396,N_14963,N_14886);
and UO_397 (O_397,N_14954,N_14966);
nand UO_398 (O_398,N_14947,N_14951);
and UO_399 (O_399,N_14895,N_14915);
nand UO_400 (O_400,N_14970,N_14996);
and UO_401 (O_401,N_14946,N_14882);
and UO_402 (O_402,N_14916,N_14942);
or UO_403 (O_403,N_14983,N_14964);
and UO_404 (O_404,N_14933,N_14910);
and UO_405 (O_405,N_14939,N_14924);
nand UO_406 (O_406,N_14888,N_14946);
xnor UO_407 (O_407,N_14906,N_14977);
xor UO_408 (O_408,N_14926,N_14895);
or UO_409 (O_409,N_14937,N_14969);
nand UO_410 (O_410,N_14959,N_14968);
or UO_411 (O_411,N_14951,N_14913);
or UO_412 (O_412,N_14896,N_14970);
and UO_413 (O_413,N_14909,N_14915);
or UO_414 (O_414,N_14979,N_14876);
nand UO_415 (O_415,N_14986,N_14887);
nor UO_416 (O_416,N_14934,N_14969);
and UO_417 (O_417,N_14921,N_14985);
or UO_418 (O_418,N_14992,N_14983);
xnor UO_419 (O_419,N_14911,N_14972);
nand UO_420 (O_420,N_14961,N_14881);
or UO_421 (O_421,N_14883,N_14934);
and UO_422 (O_422,N_14879,N_14937);
nand UO_423 (O_423,N_14942,N_14875);
nor UO_424 (O_424,N_14959,N_14904);
nor UO_425 (O_425,N_14888,N_14998);
or UO_426 (O_426,N_14973,N_14948);
nor UO_427 (O_427,N_14887,N_14930);
xnor UO_428 (O_428,N_14948,N_14957);
or UO_429 (O_429,N_14962,N_14971);
and UO_430 (O_430,N_14876,N_14938);
and UO_431 (O_431,N_14902,N_14992);
xor UO_432 (O_432,N_14946,N_14952);
xnor UO_433 (O_433,N_14916,N_14954);
nand UO_434 (O_434,N_14971,N_14945);
and UO_435 (O_435,N_14906,N_14975);
nand UO_436 (O_436,N_14981,N_14886);
nand UO_437 (O_437,N_14998,N_14944);
and UO_438 (O_438,N_14876,N_14919);
and UO_439 (O_439,N_14937,N_14920);
or UO_440 (O_440,N_14923,N_14978);
or UO_441 (O_441,N_14984,N_14994);
nor UO_442 (O_442,N_14875,N_14972);
nor UO_443 (O_443,N_14968,N_14899);
nor UO_444 (O_444,N_14971,N_14953);
and UO_445 (O_445,N_14948,N_14916);
and UO_446 (O_446,N_14918,N_14986);
and UO_447 (O_447,N_14904,N_14973);
nand UO_448 (O_448,N_14985,N_14875);
xnor UO_449 (O_449,N_14915,N_14927);
or UO_450 (O_450,N_14972,N_14960);
and UO_451 (O_451,N_14974,N_14919);
nand UO_452 (O_452,N_14884,N_14889);
nor UO_453 (O_453,N_14992,N_14906);
nor UO_454 (O_454,N_14912,N_14894);
xor UO_455 (O_455,N_14880,N_14887);
nand UO_456 (O_456,N_14993,N_14960);
or UO_457 (O_457,N_14966,N_14887);
and UO_458 (O_458,N_14929,N_14921);
and UO_459 (O_459,N_14908,N_14955);
nor UO_460 (O_460,N_14944,N_14942);
nor UO_461 (O_461,N_14938,N_14956);
or UO_462 (O_462,N_14886,N_14879);
and UO_463 (O_463,N_14906,N_14990);
xor UO_464 (O_464,N_14945,N_14963);
xor UO_465 (O_465,N_14909,N_14992);
and UO_466 (O_466,N_14895,N_14885);
nor UO_467 (O_467,N_14889,N_14980);
nor UO_468 (O_468,N_14894,N_14901);
and UO_469 (O_469,N_14896,N_14967);
xor UO_470 (O_470,N_14977,N_14964);
and UO_471 (O_471,N_14921,N_14909);
nand UO_472 (O_472,N_14979,N_14904);
or UO_473 (O_473,N_14997,N_14888);
nand UO_474 (O_474,N_14976,N_14919);
and UO_475 (O_475,N_14894,N_14971);
xnor UO_476 (O_476,N_14937,N_14906);
and UO_477 (O_477,N_14924,N_14925);
nand UO_478 (O_478,N_14930,N_14961);
and UO_479 (O_479,N_14960,N_14961);
xor UO_480 (O_480,N_14923,N_14967);
nor UO_481 (O_481,N_14968,N_14937);
xnor UO_482 (O_482,N_14939,N_14933);
and UO_483 (O_483,N_14881,N_14993);
or UO_484 (O_484,N_14994,N_14883);
xnor UO_485 (O_485,N_14916,N_14905);
nor UO_486 (O_486,N_14986,N_14987);
nor UO_487 (O_487,N_14984,N_14964);
and UO_488 (O_488,N_14897,N_14994);
nand UO_489 (O_489,N_14974,N_14910);
or UO_490 (O_490,N_14904,N_14963);
or UO_491 (O_491,N_14896,N_14924);
or UO_492 (O_492,N_14977,N_14887);
xnor UO_493 (O_493,N_14891,N_14985);
nand UO_494 (O_494,N_14913,N_14914);
nor UO_495 (O_495,N_14932,N_14950);
nand UO_496 (O_496,N_14898,N_14950);
nor UO_497 (O_497,N_14932,N_14954);
and UO_498 (O_498,N_14886,N_14942);
or UO_499 (O_499,N_14891,N_14944);
nor UO_500 (O_500,N_14896,N_14982);
nor UO_501 (O_501,N_14906,N_14891);
or UO_502 (O_502,N_14895,N_14909);
and UO_503 (O_503,N_14957,N_14988);
xor UO_504 (O_504,N_14954,N_14942);
xor UO_505 (O_505,N_14990,N_14982);
xor UO_506 (O_506,N_14971,N_14993);
xor UO_507 (O_507,N_14896,N_14996);
and UO_508 (O_508,N_14979,N_14879);
and UO_509 (O_509,N_14996,N_14912);
and UO_510 (O_510,N_14884,N_14954);
nor UO_511 (O_511,N_14981,N_14985);
or UO_512 (O_512,N_14923,N_14973);
nor UO_513 (O_513,N_14970,N_14940);
nand UO_514 (O_514,N_14884,N_14915);
nor UO_515 (O_515,N_14970,N_14899);
xor UO_516 (O_516,N_14978,N_14913);
nor UO_517 (O_517,N_14921,N_14903);
nor UO_518 (O_518,N_14957,N_14942);
nand UO_519 (O_519,N_14934,N_14897);
and UO_520 (O_520,N_14995,N_14982);
nand UO_521 (O_521,N_14951,N_14881);
and UO_522 (O_522,N_14955,N_14898);
nand UO_523 (O_523,N_14893,N_14897);
xnor UO_524 (O_524,N_14881,N_14975);
or UO_525 (O_525,N_14900,N_14992);
nand UO_526 (O_526,N_14904,N_14919);
nor UO_527 (O_527,N_14964,N_14999);
xor UO_528 (O_528,N_14985,N_14969);
nand UO_529 (O_529,N_14890,N_14974);
nand UO_530 (O_530,N_14972,N_14916);
and UO_531 (O_531,N_14957,N_14960);
and UO_532 (O_532,N_14950,N_14955);
and UO_533 (O_533,N_14953,N_14876);
nand UO_534 (O_534,N_14954,N_14936);
or UO_535 (O_535,N_14924,N_14907);
xnor UO_536 (O_536,N_14973,N_14895);
or UO_537 (O_537,N_14891,N_14939);
nor UO_538 (O_538,N_14961,N_14899);
nand UO_539 (O_539,N_14941,N_14887);
and UO_540 (O_540,N_14935,N_14875);
xor UO_541 (O_541,N_14985,N_14927);
and UO_542 (O_542,N_14900,N_14959);
nand UO_543 (O_543,N_14940,N_14989);
nor UO_544 (O_544,N_14954,N_14924);
nor UO_545 (O_545,N_14918,N_14887);
xnor UO_546 (O_546,N_14910,N_14999);
nand UO_547 (O_547,N_14957,N_14981);
nor UO_548 (O_548,N_14947,N_14917);
and UO_549 (O_549,N_14896,N_14977);
and UO_550 (O_550,N_14940,N_14952);
or UO_551 (O_551,N_14971,N_14950);
nor UO_552 (O_552,N_14962,N_14963);
nor UO_553 (O_553,N_14975,N_14989);
or UO_554 (O_554,N_14913,N_14895);
nand UO_555 (O_555,N_14876,N_14900);
or UO_556 (O_556,N_14884,N_14971);
xor UO_557 (O_557,N_14903,N_14888);
or UO_558 (O_558,N_14975,N_14960);
nand UO_559 (O_559,N_14962,N_14936);
and UO_560 (O_560,N_14948,N_14971);
and UO_561 (O_561,N_14900,N_14994);
or UO_562 (O_562,N_14943,N_14961);
and UO_563 (O_563,N_14897,N_14948);
and UO_564 (O_564,N_14933,N_14966);
nor UO_565 (O_565,N_14951,N_14931);
nor UO_566 (O_566,N_14926,N_14935);
nor UO_567 (O_567,N_14955,N_14978);
nor UO_568 (O_568,N_14929,N_14875);
and UO_569 (O_569,N_14984,N_14999);
and UO_570 (O_570,N_14916,N_14877);
xor UO_571 (O_571,N_14956,N_14931);
xnor UO_572 (O_572,N_14883,N_14890);
nand UO_573 (O_573,N_14959,N_14934);
xnor UO_574 (O_574,N_14977,N_14889);
nor UO_575 (O_575,N_14939,N_14937);
xor UO_576 (O_576,N_14901,N_14884);
or UO_577 (O_577,N_14918,N_14964);
and UO_578 (O_578,N_14940,N_14947);
and UO_579 (O_579,N_14945,N_14911);
nor UO_580 (O_580,N_14883,N_14979);
and UO_581 (O_581,N_14966,N_14972);
or UO_582 (O_582,N_14889,N_14902);
nor UO_583 (O_583,N_14982,N_14938);
xor UO_584 (O_584,N_14996,N_14880);
xor UO_585 (O_585,N_14894,N_14908);
nor UO_586 (O_586,N_14912,N_14921);
and UO_587 (O_587,N_14978,N_14935);
xnor UO_588 (O_588,N_14956,N_14937);
xnor UO_589 (O_589,N_14984,N_14942);
or UO_590 (O_590,N_14880,N_14896);
xnor UO_591 (O_591,N_14978,N_14894);
nor UO_592 (O_592,N_14882,N_14975);
nor UO_593 (O_593,N_14973,N_14880);
xnor UO_594 (O_594,N_14939,N_14875);
xor UO_595 (O_595,N_14974,N_14899);
and UO_596 (O_596,N_14998,N_14978);
or UO_597 (O_597,N_14928,N_14975);
and UO_598 (O_598,N_14928,N_14922);
or UO_599 (O_599,N_14878,N_14890);
and UO_600 (O_600,N_14887,N_14992);
xor UO_601 (O_601,N_14887,N_14912);
or UO_602 (O_602,N_14891,N_14958);
nand UO_603 (O_603,N_14948,N_14901);
nor UO_604 (O_604,N_14905,N_14912);
nor UO_605 (O_605,N_14959,N_14899);
xnor UO_606 (O_606,N_14920,N_14979);
and UO_607 (O_607,N_14877,N_14989);
or UO_608 (O_608,N_14910,N_14893);
or UO_609 (O_609,N_14999,N_14995);
or UO_610 (O_610,N_14918,N_14994);
nor UO_611 (O_611,N_14894,N_14943);
and UO_612 (O_612,N_14978,N_14969);
or UO_613 (O_613,N_14994,N_14964);
or UO_614 (O_614,N_14913,N_14958);
and UO_615 (O_615,N_14887,N_14878);
nand UO_616 (O_616,N_14953,N_14975);
and UO_617 (O_617,N_14932,N_14888);
nand UO_618 (O_618,N_14969,N_14995);
or UO_619 (O_619,N_14932,N_14971);
nand UO_620 (O_620,N_14963,N_14931);
nor UO_621 (O_621,N_14946,N_14980);
or UO_622 (O_622,N_14921,N_14922);
nor UO_623 (O_623,N_14937,N_14986);
nor UO_624 (O_624,N_14978,N_14985);
or UO_625 (O_625,N_14996,N_14965);
xor UO_626 (O_626,N_14917,N_14953);
nor UO_627 (O_627,N_14963,N_14965);
or UO_628 (O_628,N_14995,N_14921);
and UO_629 (O_629,N_14940,N_14949);
or UO_630 (O_630,N_14968,N_14990);
xnor UO_631 (O_631,N_14882,N_14984);
nor UO_632 (O_632,N_14930,N_14956);
or UO_633 (O_633,N_14905,N_14897);
nand UO_634 (O_634,N_14985,N_14880);
nor UO_635 (O_635,N_14876,N_14918);
xnor UO_636 (O_636,N_14942,N_14915);
nand UO_637 (O_637,N_14987,N_14972);
nor UO_638 (O_638,N_14901,N_14959);
nor UO_639 (O_639,N_14952,N_14886);
or UO_640 (O_640,N_14984,N_14927);
xnor UO_641 (O_641,N_14975,N_14998);
xor UO_642 (O_642,N_14975,N_14922);
and UO_643 (O_643,N_14903,N_14948);
nand UO_644 (O_644,N_14883,N_14919);
nor UO_645 (O_645,N_14979,N_14877);
and UO_646 (O_646,N_14954,N_14965);
nor UO_647 (O_647,N_14899,N_14883);
nand UO_648 (O_648,N_14966,N_14987);
nor UO_649 (O_649,N_14996,N_14980);
xnor UO_650 (O_650,N_14902,N_14982);
xor UO_651 (O_651,N_14882,N_14904);
nor UO_652 (O_652,N_14949,N_14899);
nand UO_653 (O_653,N_14967,N_14881);
nor UO_654 (O_654,N_14959,N_14945);
or UO_655 (O_655,N_14914,N_14966);
and UO_656 (O_656,N_14974,N_14977);
nand UO_657 (O_657,N_14906,N_14880);
and UO_658 (O_658,N_14986,N_14894);
nor UO_659 (O_659,N_14970,N_14893);
xnor UO_660 (O_660,N_14925,N_14965);
xnor UO_661 (O_661,N_14924,N_14914);
and UO_662 (O_662,N_14959,N_14894);
and UO_663 (O_663,N_14959,N_14910);
nor UO_664 (O_664,N_14915,N_14963);
xor UO_665 (O_665,N_14919,N_14928);
nand UO_666 (O_666,N_14938,N_14978);
nand UO_667 (O_667,N_14949,N_14882);
nor UO_668 (O_668,N_14945,N_14982);
xor UO_669 (O_669,N_14894,N_14942);
nor UO_670 (O_670,N_14977,N_14907);
nand UO_671 (O_671,N_14898,N_14999);
xnor UO_672 (O_672,N_14950,N_14934);
nor UO_673 (O_673,N_14950,N_14938);
xor UO_674 (O_674,N_14898,N_14884);
xnor UO_675 (O_675,N_14966,N_14911);
or UO_676 (O_676,N_14929,N_14967);
xor UO_677 (O_677,N_14916,N_14927);
nor UO_678 (O_678,N_14932,N_14914);
and UO_679 (O_679,N_14896,N_14908);
xnor UO_680 (O_680,N_14939,N_14930);
xnor UO_681 (O_681,N_14979,N_14942);
or UO_682 (O_682,N_14919,N_14939);
nand UO_683 (O_683,N_14984,N_14924);
and UO_684 (O_684,N_14972,N_14981);
and UO_685 (O_685,N_14895,N_14893);
or UO_686 (O_686,N_14936,N_14952);
nor UO_687 (O_687,N_14916,N_14891);
nand UO_688 (O_688,N_14886,N_14962);
nor UO_689 (O_689,N_14938,N_14932);
nor UO_690 (O_690,N_14875,N_14890);
or UO_691 (O_691,N_14986,N_14892);
nor UO_692 (O_692,N_14989,N_14895);
or UO_693 (O_693,N_14939,N_14956);
and UO_694 (O_694,N_14906,N_14960);
or UO_695 (O_695,N_14885,N_14920);
xor UO_696 (O_696,N_14897,N_14961);
xnor UO_697 (O_697,N_14952,N_14947);
nor UO_698 (O_698,N_14994,N_14973);
xor UO_699 (O_699,N_14990,N_14967);
or UO_700 (O_700,N_14894,N_14889);
xor UO_701 (O_701,N_14941,N_14977);
nor UO_702 (O_702,N_14907,N_14987);
nor UO_703 (O_703,N_14963,N_14903);
nand UO_704 (O_704,N_14981,N_14946);
and UO_705 (O_705,N_14969,N_14915);
and UO_706 (O_706,N_14933,N_14877);
nor UO_707 (O_707,N_14900,N_14924);
xor UO_708 (O_708,N_14956,N_14996);
or UO_709 (O_709,N_14996,N_14921);
nand UO_710 (O_710,N_14952,N_14883);
nor UO_711 (O_711,N_14888,N_14913);
nand UO_712 (O_712,N_14914,N_14909);
nand UO_713 (O_713,N_14959,N_14922);
nand UO_714 (O_714,N_14975,N_14990);
nand UO_715 (O_715,N_14954,N_14975);
nand UO_716 (O_716,N_14989,N_14904);
and UO_717 (O_717,N_14950,N_14941);
nand UO_718 (O_718,N_14973,N_14924);
or UO_719 (O_719,N_14887,N_14888);
or UO_720 (O_720,N_14921,N_14952);
nor UO_721 (O_721,N_14944,N_14994);
xnor UO_722 (O_722,N_14987,N_14926);
and UO_723 (O_723,N_14984,N_14935);
nand UO_724 (O_724,N_14886,N_14893);
nand UO_725 (O_725,N_14920,N_14936);
nand UO_726 (O_726,N_14892,N_14909);
nand UO_727 (O_727,N_14900,N_14932);
or UO_728 (O_728,N_14953,N_14886);
nand UO_729 (O_729,N_14950,N_14953);
nand UO_730 (O_730,N_14894,N_14898);
or UO_731 (O_731,N_14974,N_14906);
nand UO_732 (O_732,N_14901,N_14947);
nand UO_733 (O_733,N_14939,N_14915);
or UO_734 (O_734,N_14997,N_14929);
nor UO_735 (O_735,N_14948,N_14975);
and UO_736 (O_736,N_14931,N_14923);
or UO_737 (O_737,N_14979,N_14934);
xnor UO_738 (O_738,N_14950,N_14939);
nand UO_739 (O_739,N_14932,N_14946);
nand UO_740 (O_740,N_14916,N_14903);
xnor UO_741 (O_741,N_14929,N_14926);
nor UO_742 (O_742,N_14879,N_14940);
xor UO_743 (O_743,N_14923,N_14988);
nand UO_744 (O_744,N_14875,N_14919);
or UO_745 (O_745,N_14910,N_14935);
xor UO_746 (O_746,N_14981,N_14932);
nand UO_747 (O_747,N_14977,N_14969);
xnor UO_748 (O_748,N_14949,N_14910);
nor UO_749 (O_749,N_14963,N_14878);
nand UO_750 (O_750,N_14968,N_14912);
nand UO_751 (O_751,N_14944,N_14961);
and UO_752 (O_752,N_14916,N_14914);
and UO_753 (O_753,N_14911,N_14925);
nor UO_754 (O_754,N_14899,N_14910);
xor UO_755 (O_755,N_14979,N_14923);
nor UO_756 (O_756,N_14993,N_14940);
xnor UO_757 (O_757,N_14909,N_14950);
xor UO_758 (O_758,N_14968,N_14975);
and UO_759 (O_759,N_14965,N_14968);
nor UO_760 (O_760,N_14968,N_14949);
nand UO_761 (O_761,N_14971,N_14875);
nand UO_762 (O_762,N_14960,N_14983);
nor UO_763 (O_763,N_14917,N_14915);
nor UO_764 (O_764,N_14946,N_14919);
nor UO_765 (O_765,N_14959,N_14877);
nor UO_766 (O_766,N_14995,N_14961);
xnor UO_767 (O_767,N_14981,N_14926);
xnor UO_768 (O_768,N_14981,N_14925);
nand UO_769 (O_769,N_14888,N_14909);
and UO_770 (O_770,N_14931,N_14940);
nand UO_771 (O_771,N_14985,N_14883);
nor UO_772 (O_772,N_14940,N_14914);
or UO_773 (O_773,N_14954,N_14908);
xor UO_774 (O_774,N_14928,N_14890);
or UO_775 (O_775,N_14957,N_14995);
xor UO_776 (O_776,N_14911,N_14875);
or UO_777 (O_777,N_14956,N_14977);
nor UO_778 (O_778,N_14962,N_14919);
or UO_779 (O_779,N_14991,N_14880);
or UO_780 (O_780,N_14922,N_14953);
xor UO_781 (O_781,N_14894,N_14900);
nand UO_782 (O_782,N_14946,N_14900);
and UO_783 (O_783,N_14968,N_14935);
nand UO_784 (O_784,N_14895,N_14878);
nor UO_785 (O_785,N_14964,N_14927);
nor UO_786 (O_786,N_14952,N_14899);
nand UO_787 (O_787,N_14938,N_14922);
nor UO_788 (O_788,N_14889,N_14937);
nand UO_789 (O_789,N_14884,N_14983);
and UO_790 (O_790,N_14999,N_14967);
or UO_791 (O_791,N_14931,N_14899);
and UO_792 (O_792,N_14957,N_14992);
and UO_793 (O_793,N_14893,N_14976);
and UO_794 (O_794,N_14894,N_14946);
nor UO_795 (O_795,N_14946,N_14928);
xor UO_796 (O_796,N_14946,N_14974);
xor UO_797 (O_797,N_14887,N_14931);
and UO_798 (O_798,N_14979,N_14922);
nand UO_799 (O_799,N_14913,N_14965);
or UO_800 (O_800,N_14911,N_14991);
xnor UO_801 (O_801,N_14935,N_14997);
xnor UO_802 (O_802,N_14973,N_14974);
xnor UO_803 (O_803,N_14972,N_14976);
nand UO_804 (O_804,N_14961,N_14962);
nand UO_805 (O_805,N_14976,N_14931);
xnor UO_806 (O_806,N_14878,N_14926);
and UO_807 (O_807,N_14969,N_14910);
and UO_808 (O_808,N_14950,N_14916);
nand UO_809 (O_809,N_14914,N_14979);
xor UO_810 (O_810,N_14897,N_14922);
nor UO_811 (O_811,N_14975,N_14908);
xor UO_812 (O_812,N_14980,N_14891);
nor UO_813 (O_813,N_14934,N_14936);
xor UO_814 (O_814,N_14934,N_14900);
nor UO_815 (O_815,N_14950,N_14922);
or UO_816 (O_816,N_14911,N_14993);
xnor UO_817 (O_817,N_14900,N_14910);
or UO_818 (O_818,N_14902,N_14931);
nand UO_819 (O_819,N_14958,N_14898);
nand UO_820 (O_820,N_14921,N_14882);
and UO_821 (O_821,N_14900,N_14918);
nand UO_822 (O_822,N_14920,N_14892);
nand UO_823 (O_823,N_14933,N_14903);
or UO_824 (O_824,N_14972,N_14910);
and UO_825 (O_825,N_14896,N_14890);
and UO_826 (O_826,N_14939,N_14952);
or UO_827 (O_827,N_14894,N_14934);
or UO_828 (O_828,N_14951,N_14968);
and UO_829 (O_829,N_14899,N_14898);
xnor UO_830 (O_830,N_14978,N_14966);
nand UO_831 (O_831,N_14966,N_14952);
nand UO_832 (O_832,N_14905,N_14989);
or UO_833 (O_833,N_14949,N_14894);
nand UO_834 (O_834,N_14934,N_14981);
nor UO_835 (O_835,N_14989,N_14985);
xor UO_836 (O_836,N_14997,N_14981);
xnor UO_837 (O_837,N_14908,N_14933);
and UO_838 (O_838,N_14972,N_14904);
nand UO_839 (O_839,N_14887,N_14983);
nand UO_840 (O_840,N_14885,N_14954);
or UO_841 (O_841,N_14946,N_14940);
and UO_842 (O_842,N_14910,N_14965);
xnor UO_843 (O_843,N_14927,N_14934);
nor UO_844 (O_844,N_14958,N_14957);
and UO_845 (O_845,N_14976,N_14886);
nor UO_846 (O_846,N_14920,N_14913);
and UO_847 (O_847,N_14981,N_14991);
nor UO_848 (O_848,N_14954,N_14994);
and UO_849 (O_849,N_14950,N_14917);
xor UO_850 (O_850,N_14954,N_14959);
nand UO_851 (O_851,N_14930,N_14923);
and UO_852 (O_852,N_14991,N_14881);
or UO_853 (O_853,N_14969,N_14906);
xor UO_854 (O_854,N_14967,N_14886);
xor UO_855 (O_855,N_14956,N_14989);
nor UO_856 (O_856,N_14913,N_14907);
xor UO_857 (O_857,N_14969,N_14944);
xor UO_858 (O_858,N_14875,N_14881);
or UO_859 (O_859,N_14910,N_14939);
and UO_860 (O_860,N_14955,N_14933);
nor UO_861 (O_861,N_14893,N_14960);
xnor UO_862 (O_862,N_14977,N_14899);
or UO_863 (O_863,N_14898,N_14969);
xnor UO_864 (O_864,N_14904,N_14902);
xnor UO_865 (O_865,N_14882,N_14896);
xnor UO_866 (O_866,N_14901,N_14952);
nand UO_867 (O_867,N_14976,N_14921);
xor UO_868 (O_868,N_14897,N_14879);
nor UO_869 (O_869,N_14927,N_14995);
and UO_870 (O_870,N_14893,N_14909);
or UO_871 (O_871,N_14894,N_14921);
nor UO_872 (O_872,N_14915,N_14993);
xor UO_873 (O_873,N_14968,N_14983);
and UO_874 (O_874,N_14977,N_14953);
xnor UO_875 (O_875,N_14882,N_14919);
and UO_876 (O_876,N_14956,N_14883);
nand UO_877 (O_877,N_14930,N_14970);
xor UO_878 (O_878,N_14915,N_14968);
nand UO_879 (O_879,N_14935,N_14912);
nor UO_880 (O_880,N_14921,N_14984);
xnor UO_881 (O_881,N_14914,N_14883);
nor UO_882 (O_882,N_14933,N_14916);
nand UO_883 (O_883,N_14973,N_14884);
and UO_884 (O_884,N_14914,N_14984);
and UO_885 (O_885,N_14987,N_14999);
or UO_886 (O_886,N_14970,N_14920);
nor UO_887 (O_887,N_14958,N_14977);
xor UO_888 (O_888,N_14894,N_14914);
nand UO_889 (O_889,N_14930,N_14996);
nand UO_890 (O_890,N_14895,N_14936);
xor UO_891 (O_891,N_14960,N_14880);
nand UO_892 (O_892,N_14948,N_14913);
nand UO_893 (O_893,N_14981,N_14889);
nand UO_894 (O_894,N_14917,N_14878);
and UO_895 (O_895,N_14920,N_14922);
nor UO_896 (O_896,N_14939,N_14940);
xnor UO_897 (O_897,N_14891,N_14926);
or UO_898 (O_898,N_14920,N_14990);
or UO_899 (O_899,N_14995,N_14888);
and UO_900 (O_900,N_14928,N_14921);
and UO_901 (O_901,N_14950,N_14991);
nand UO_902 (O_902,N_14949,N_14887);
xor UO_903 (O_903,N_14914,N_14995);
nor UO_904 (O_904,N_14959,N_14992);
or UO_905 (O_905,N_14887,N_14899);
or UO_906 (O_906,N_14943,N_14896);
or UO_907 (O_907,N_14925,N_14929);
nor UO_908 (O_908,N_14891,N_14943);
xnor UO_909 (O_909,N_14949,N_14966);
xnor UO_910 (O_910,N_14937,N_14985);
and UO_911 (O_911,N_14898,N_14989);
nor UO_912 (O_912,N_14974,N_14938);
nor UO_913 (O_913,N_14975,N_14904);
or UO_914 (O_914,N_14905,N_14926);
nor UO_915 (O_915,N_14963,N_14923);
or UO_916 (O_916,N_14928,N_14909);
or UO_917 (O_917,N_14933,N_14962);
or UO_918 (O_918,N_14988,N_14889);
nand UO_919 (O_919,N_14959,N_14983);
nand UO_920 (O_920,N_14960,N_14951);
or UO_921 (O_921,N_14896,N_14965);
nor UO_922 (O_922,N_14959,N_14893);
and UO_923 (O_923,N_14924,N_14957);
nor UO_924 (O_924,N_14932,N_14961);
nand UO_925 (O_925,N_14895,N_14992);
nand UO_926 (O_926,N_14982,N_14977);
or UO_927 (O_927,N_14902,N_14943);
and UO_928 (O_928,N_14990,N_14886);
xor UO_929 (O_929,N_14891,N_14933);
nand UO_930 (O_930,N_14949,N_14952);
and UO_931 (O_931,N_14985,N_14976);
nand UO_932 (O_932,N_14979,N_14910);
or UO_933 (O_933,N_14933,N_14991);
xor UO_934 (O_934,N_14965,N_14901);
nor UO_935 (O_935,N_14897,N_14958);
nand UO_936 (O_936,N_14894,N_14909);
nor UO_937 (O_937,N_14906,N_14968);
or UO_938 (O_938,N_14913,N_14904);
and UO_939 (O_939,N_14890,N_14877);
nand UO_940 (O_940,N_14889,N_14944);
xor UO_941 (O_941,N_14953,N_14974);
and UO_942 (O_942,N_14959,N_14996);
or UO_943 (O_943,N_14892,N_14893);
or UO_944 (O_944,N_14904,N_14894);
nand UO_945 (O_945,N_14939,N_14989);
nor UO_946 (O_946,N_14968,N_14984);
nor UO_947 (O_947,N_14961,N_14894);
or UO_948 (O_948,N_14943,N_14912);
nor UO_949 (O_949,N_14888,N_14938);
xor UO_950 (O_950,N_14937,N_14982);
nor UO_951 (O_951,N_14910,N_14962);
or UO_952 (O_952,N_14889,N_14897);
or UO_953 (O_953,N_14920,N_14946);
and UO_954 (O_954,N_14973,N_14989);
and UO_955 (O_955,N_14919,N_14911);
or UO_956 (O_956,N_14993,N_14917);
or UO_957 (O_957,N_14945,N_14939);
nand UO_958 (O_958,N_14979,N_14925);
or UO_959 (O_959,N_14876,N_14996);
nand UO_960 (O_960,N_14963,N_14875);
and UO_961 (O_961,N_14941,N_14928);
nor UO_962 (O_962,N_14893,N_14919);
xor UO_963 (O_963,N_14888,N_14940);
nand UO_964 (O_964,N_14992,N_14939);
nand UO_965 (O_965,N_14885,N_14879);
nand UO_966 (O_966,N_14940,N_14933);
and UO_967 (O_967,N_14931,N_14939);
nor UO_968 (O_968,N_14922,N_14951);
or UO_969 (O_969,N_14902,N_14941);
nor UO_970 (O_970,N_14947,N_14899);
xnor UO_971 (O_971,N_14903,N_14886);
nor UO_972 (O_972,N_14918,N_14935);
and UO_973 (O_973,N_14992,N_14899);
and UO_974 (O_974,N_14936,N_14998);
nor UO_975 (O_975,N_14931,N_14924);
xnor UO_976 (O_976,N_14934,N_14921);
xor UO_977 (O_977,N_14898,N_14877);
xor UO_978 (O_978,N_14981,N_14904);
and UO_979 (O_979,N_14996,N_14923);
nor UO_980 (O_980,N_14957,N_14880);
and UO_981 (O_981,N_14962,N_14913);
xnor UO_982 (O_982,N_14947,N_14962);
xnor UO_983 (O_983,N_14970,N_14924);
and UO_984 (O_984,N_14990,N_14953);
xnor UO_985 (O_985,N_14906,N_14988);
or UO_986 (O_986,N_14983,N_14947);
and UO_987 (O_987,N_14940,N_14909);
nor UO_988 (O_988,N_14958,N_14995);
and UO_989 (O_989,N_14881,N_14988);
xnor UO_990 (O_990,N_14997,N_14886);
nor UO_991 (O_991,N_14911,N_14901);
nand UO_992 (O_992,N_14876,N_14908);
nor UO_993 (O_993,N_14947,N_14970);
or UO_994 (O_994,N_14958,N_14956);
and UO_995 (O_995,N_14905,N_14945);
nor UO_996 (O_996,N_14926,N_14923);
xor UO_997 (O_997,N_14958,N_14907);
xor UO_998 (O_998,N_14929,N_14991);
and UO_999 (O_999,N_14923,N_14900);
and UO_1000 (O_1000,N_14999,N_14925);
xnor UO_1001 (O_1001,N_14953,N_14941);
nand UO_1002 (O_1002,N_14998,N_14946);
and UO_1003 (O_1003,N_14959,N_14912);
xnor UO_1004 (O_1004,N_14966,N_14971);
or UO_1005 (O_1005,N_14970,N_14903);
nand UO_1006 (O_1006,N_14979,N_14952);
and UO_1007 (O_1007,N_14904,N_14922);
or UO_1008 (O_1008,N_14927,N_14956);
and UO_1009 (O_1009,N_14969,N_14949);
xnor UO_1010 (O_1010,N_14985,N_14971);
xor UO_1011 (O_1011,N_14876,N_14904);
or UO_1012 (O_1012,N_14956,N_14890);
nand UO_1013 (O_1013,N_14916,N_14890);
and UO_1014 (O_1014,N_14898,N_14917);
xnor UO_1015 (O_1015,N_14986,N_14881);
or UO_1016 (O_1016,N_14898,N_14991);
and UO_1017 (O_1017,N_14972,N_14959);
and UO_1018 (O_1018,N_14938,N_14954);
nor UO_1019 (O_1019,N_14905,N_14915);
nor UO_1020 (O_1020,N_14897,N_14985);
nor UO_1021 (O_1021,N_14920,N_14991);
xnor UO_1022 (O_1022,N_14995,N_14895);
or UO_1023 (O_1023,N_14935,N_14894);
nand UO_1024 (O_1024,N_14976,N_14891);
xor UO_1025 (O_1025,N_14906,N_14954);
and UO_1026 (O_1026,N_14980,N_14928);
or UO_1027 (O_1027,N_14881,N_14980);
or UO_1028 (O_1028,N_14961,N_14922);
or UO_1029 (O_1029,N_14952,N_14992);
nor UO_1030 (O_1030,N_14955,N_14980);
or UO_1031 (O_1031,N_14889,N_14881);
nor UO_1032 (O_1032,N_14945,N_14946);
and UO_1033 (O_1033,N_14888,N_14968);
nor UO_1034 (O_1034,N_14986,N_14945);
or UO_1035 (O_1035,N_14985,N_14881);
nand UO_1036 (O_1036,N_14892,N_14924);
or UO_1037 (O_1037,N_14963,N_14938);
nor UO_1038 (O_1038,N_14879,N_14983);
and UO_1039 (O_1039,N_14934,N_14987);
and UO_1040 (O_1040,N_14956,N_14910);
or UO_1041 (O_1041,N_14899,N_14938);
nor UO_1042 (O_1042,N_14940,N_14918);
nand UO_1043 (O_1043,N_14988,N_14904);
xnor UO_1044 (O_1044,N_14891,N_14881);
xnor UO_1045 (O_1045,N_14915,N_14919);
nor UO_1046 (O_1046,N_14981,N_14998);
xnor UO_1047 (O_1047,N_14879,N_14998);
or UO_1048 (O_1048,N_14917,N_14963);
nor UO_1049 (O_1049,N_14876,N_14967);
nor UO_1050 (O_1050,N_14944,N_14900);
nand UO_1051 (O_1051,N_14890,N_14901);
and UO_1052 (O_1052,N_14907,N_14996);
or UO_1053 (O_1053,N_14903,N_14908);
or UO_1054 (O_1054,N_14972,N_14990);
or UO_1055 (O_1055,N_14969,N_14892);
xnor UO_1056 (O_1056,N_14945,N_14883);
nand UO_1057 (O_1057,N_14926,N_14970);
or UO_1058 (O_1058,N_14897,N_14932);
xnor UO_1059 (O_1059,N_14920,N_14899);
or UO_1060 (O_1060,N_14927,N_14896);
xnor UO_1061 (O_1061,N_14999,N_14943);
and UO_1062 (O_1062,N_14965,N_14971);
nor UO_1063 (O_1063,N_14970,N_14982);
or UO_1064 (O_1064,N_14885,N_14901);
or UO_1065 (O_1065,N_14927,N_14945);
and UO_1066 (O_1066,N_14974,N_14898);
nand UO_1067 (O_1067,N_14924,N_14948);
nor UO_1068 (O_1068,N_14968,N_14900);
xnor UO_1069 (O_1069,N_14984,N_14915);
xor UO_1070 (O_1070,N_14958,N_14954);
and UO_1071 (O_1071,N_14877,N_14999);
xor UO_1072 (O_1072,N_14896,N_14900);
nor UO_1073 (O_1073,N_14914,N_14998);
or UO_1074 (O_1074,N_14984,N_14904);
or UO_1075 (O_1075,N_14985,N_14951);
xnor UO_1076 (O_1076,N_14955,N_14899);
nor UO_1077 (O_1077,N_14889,N_14973);
nand UO_1078 (O_1078,N_14934,N_14913);
nand UO_1079 (O_1079,N_14978,N_14933);
xnor UO_1080 (O_1080,N_14924,N_14886);
nand UO_1081 (O_1081,N_14883,N_14993);
and UO_1082 (O_1082,N_14977,N_14970);
or UO_1083 (O_1083,N_14997,N_14924);
or UO_1084 (O_1084,N_14973,N_14910);
nand UO_1085 (O_1085,N_14959,N_14977);
xnor UO_1086 (O_1086,N_14964,N_14979);
and UO_1087 (O_1087,N_14943,N_14901);
and UO_1088 (O_1088,N_14974,N_14942);
nor UO_1089 (O_1089,N_14908,N_14899);
nand UO_1090 (O_1090,N_14907,N_14933);
nor UO_1091 (O_1091,N_14915,N_14897);
nand UO_1092 (O_1092,N_14959,N_14908);
nor UO_1093 (O_1093,N_14884,N_14976);
xor UO_1094 (O_1094,N_14875,N_14977);
xor UO_1095 (O_1095,N_14954,N_14921);
nor UO_1096 (O_1096,N_14889,N_14942);
nor UO_1097 (O_1097,N_14915,N_14985);
nand UO_1098 (O_1098,N_14911,N_14937);
xnor UO_1099 (O_1099,N_14876,N_14926);
and UO_1100 (O_1100,N_14950,N_14927);
or UO_1101 (O_1101,N_14980,N_14893);
nand UO_1102 (O_1102,N_14896,N_14962);
nor UO_1103 (O_1103,N_14940,N_14985);
or UO_1104 (O_1104,N_14895,N_14988);
nand UO_1105 (O_1105,N_14976,N_14888);
or UO_1106 (O_1106,N_14978,N_14915);
nor UO_1107 (O_1107,N_14886,N_14968);
nor UO_1108 (O_1108,N_14883,N_14986);
and UO_1109 (O_1109,N_14877,N_14947);
nor UO_1110 (O_1110,N_14915,N_14973);
nor UO_1111 (O_1111,N_14932,N_14985);
and UO_1112 (O_1112,N_14914,N_14997);
or UO_1113 (O_1113,N_14984,N_14932);
nand UO_1114 (O_1114,N_14946,N_14995);
or UO_1115 (O_1115,N_14981,N_14912);
xnor UO_1116 (O_1116,N_14892,N_14910);
or UO_1117 (O_1117,N_14891,N_14940);
nor UO_1118 (O_1118,N_14977,N_14935);
and UO_1119 (O_1119,N_14957,N_14994);
nor UO_1120 (O_1120,N_14907,N_14936);
nand UO_1121 (O_1121,N_14967,N_14948);
nand UO_1122 (O_1122,N_14898,N_14972);
nand UO_1123 (O_1123,N_14925,N_14955);
and UO_1124 (O_1124,N_14993,N_14908);
and UO_1125 (O_1125,N_14952,N_14965);
nor UO_1126 (O_1126,N_14899,N_14921);
xor UO_1127 (O_1127,N_14875,N_14955);
or UO_1128 (O_1128,N_14926,N_14966);
nand UO_1129 (O_1129,N_14875,N_14958);
and UO_1130 (O_1130,N_14892,N_14990);
nor UO_1131 (O_1131,N_14927,N_14947);
and UO_1132 (O_1132,N_14894,N_14974);
xnor UO_1133 (O_1133,N_14957,N_14974);
xnor UO_1134 (O_1134,N_14954,N_14985);
or UO_1135 (O_1135,N_14952,N_14970);
and UO_1136 (O_1136,N_14989,N_14902);
nand UO_1137 (O_1137,N_14920,N_14888);
xnor UO_1138 (O_1138,N_14972,N_14964);
xnor UO_1139 (O_1139,N_14931,N_14884);
xor UO_1140 (O_1140,N_14896,N_14981);
nor UO_1141 (O_1141,N_14946,N_14907);
nor UO_1142 (O_1142,N_14919,N_14937);
and UO_1143 (O_1143,N_14919,N_14934);
nand UO_1144 (O_1144,N_14876,N_14896);
nor UO_1145 (O_1145,N_14949,N_14895);
nand UO_1146 (O_1146,N_14906,N_14938);
nand UO_1147 (O_1147,N_14977,N_14972);
or UO_1148 (O_1148,N_14881,N_14933);
or UO_1149 (O_1149,N_14988,N_14915);
nor UO_1150 (O_1150,N_14925,N_14890);
nand UO_1151 (O_1151,N_14993,N_14943);
nor UO_1152 (O_1152,N_14982,N_14876);
nand UO_1153 (O_1153,N_14876,N_14942);
and UO_1154 (O_1154,N_14923,N_14925);
nand UO_1155 (O_1155,N_14945,N_14991);
or UO_1156 (O_1156,N_14993,N_14882);
nand UO_1157 (O_1157,N_14958,N_14906);
nor UO_1158 (O_1158,N_14971,N_14964);
xnor UO_1159 (O_1159,N_14999,N_14899);
xor UO_1160 (O_1160,N_14881,N_14898);
and UO_1161 (O_1161,N_14975,N_14920);
or UO_1162 (O_1162,N_14903,N_14932);
and UO_1163 (O_1163,N_14917,N_14890);
nand UO_1164 (O_1164,N_14883,N_14916);
nand UO_1165 (O_1165,N_14928,N_14974);
nand UO_1166 (O_1166,N_14876,N_14916);
or UO_1167 (O_1167,N_14897,N_14929);
nor UO_1168 (O_1168,N_14900,N_14938);
nor UO_1169 (O_1169,N_14923,N_14888);
and UO_1170 (O_1170,N_14946,N_14889);
nor UO_1171 (O_1171,N_14968,N_14928);
nor UO_1172 (O_1172,N_14969,N_14916);
nor UO_1173 (O_1173,N_14899,N_14988);
nor UO_1174 (O_1174,N_14918,N_14993);
or UO_1175 (O_1175,N_14949,N_14886);
or UO_1176 (O_1176,N_14930,N_14929);
xor UO_1177 (O_1177,N_14930,N_14919);
and UO_1178 (O_1178,N_14993,N_14876);
xnor UO_1179 (O_1179,N_14926,N_14977);
xor UO_1180 (O_1180,N_14963,N_14913);
nor UO_1181 (O_1181,N_14973,N_14966);
or UO_1182 (O_1182,N_14896,N_14966);
nor UO_1183 (O_1183,N_14958,N_14878);
xnor UO_1184 (O_1184,N_14926,N_14944);
nand UO_1185 (O_1185,N_14908,N_14952);
nor UO_1186 (O_1186,N_14982,N_14915);
xnor UO_1187 (O_1187,N_14902,N_14954);
or UO_1188 (O_1188,N_14931,N_14997);
xnor UO_1189 (O_1189,N_14926,N_14990);
nand UO_1190 (O_1190,N_14894,N_14899);
nor UO_1191 (O_1191,N_14936,N_14956);
and UO_1192 (O_1192,N_14995,N_14950);
xnor UO_1193 (O_1193,N_14967,N_14888);
nand UO_1194 (O_1194,N_14974,N_14895);
nand UO_1195 (O_1195,N_14975,N_14927);
nor UO_1196 (O_1196,N_14983,N_14952);
and UO_1197 (O_1197,N_14982,N_14882);
nor UO_1198 (O_1198,N_14935,N_14882);
nor UO_1199 (O_1199,N_14897,N_14875);
xnor UO_1200 (O_1200,N_14932,N_14956);
nor UO_1201 (O_1201,N_14914,N_14899);
nand UO_1202 (O_1202,N_14976,N_14918);
or UO_1203 (O_1203,N_14939,N_14877);
xnor UO_1204 (O_1204,N_14900,N_14983);
or UO_1205 (O_1205,N_14984,N_14875);
and UO_1206 (O_1206,N_14974,N_14885);
and UO_1207 (O_1207,N_14978,N_14916);
and UO_1208 (O_1208,N_14998,N_14953);
or UO_1209 (O_1209,N_14932,N_14913);
xor UO_1210 (O_1210,N_14961,N_14903);
nand UO_1211 (O_1211,N_14964,N_14919);
and UO_1212 (O_1212,N_14933,N_14883);
nor UO_1213 (O_1213,N_14891,N_14929);
nor UO_1214 (O_1214,N_14923,N_14907);
or UO_1215 (O_1215,N_14932,N_14904);
xnor UO_1216 (O_1216,N_14912,N_14883);
nor UO_1217 (O_1217,N_14938,N_14917);
or UO_1218 (O_1218,N_14896,N_14979);
or UO_1219 (O_1219,N_14975,N_14961);
nand UO_1220 (O_1220,N_14901,N_14968);
or UO_1221 (O_1221,N_14906,N_14898);
or UO_1222 (O_1222,N_14910,N_14909);
xnor UO_1223 (O_1223,N_14950,N_14975);
xor UO_1224 (O_1224,N_14975,N_14977);
nor UO_1225 (O_1225,N_14910,N_14914);
nor UO_1226 (O_1226,N_14956,N_14875);
nand UO_1227 (O_1227,N_14988,N_14948);
nor UO_1228 (O_1228,N_14902,N_14906);
and UO_1229 (O_1229,N_14975,N_14932);
and UO_1230 (O_1230,N_14989,N_14963);
or UO_1231 (O_1231,N_14890,N_14991);
nand UO_1232 (O_1232,N_14931,N_14921);
nor UO_1233 (O_1233,N_14995,N_14963);
nand UO_1234 (O_1234,N_14934,N_14906);
or UO_1235 (O_1235,N_14925,N_14876);
nor UO_1236 (O_1236,N_14908,N_14977);
and UO_1237 (O_1237,N_14950,N_14900);
and UO_1238 (O_1238,N_14951,N_14974);
nor UO_1239 (O_1239,N_14892,N_14898);
xor UO_1240 (O_1240,N_14982,N_14985);
nand UO_1241 (O_1241,N_14911,N_14978);
or UO_1242 (O_1242,N_14903,N_14901);
or UO_1243 (O_1243,N_14896,N_14904);
and UO_1244 (O_1244,N_14906,N_14953);
or UO_1245 (O_1245,N_14961,N_14883);
nor UO_1246 (O_1246,N_14941,N_14878);
and UO_1247 (O_1247,N_14950,N_14944);
xor UO_1248 (O_1248,N_14968,N_14938);
nand UO_1249 (O_1249,N_14943,N_14932);
or UO_1250 (O_1250,N_14878,N_14898);
nand UO_1251 (O_1251,N_14934,N_14954);
and UO_1252 (O_1252,N_14943,N_14887);
or UO_1253 (O_1253,N_14929,N_14976);
xnor UO_1254 (O_1254,N_14912,N_14999);
and UO_1255 (O_1255,N_14990,N_14996);
xor UO_1256 (O_1256,N_14952,N_14997);
and UO_1257 (O_1257,N_14985,N_14962);
and UO_1258 (O_1258,N_14993,N_14875);
xor UO_1259 (O_1259,N_14895,N_14968);
or UO_1260 (O_1260,N_14927,N_14977);
or UO_1261 (O_1261,N_14913,N_14999);
xor UO_1262 (O_1262,N_14953,N_14994);
or UO_1263 (O_1263,N_14965,N_14944);
or UO_1264 (O_1264,N_14987,N_14929);
or UO_1265 (O_1265,N_14932,N_14924);
or UO_1266 (O_1266,N_14892,N_14937);
xnor UO_1267 (O_1267,N_14884,N_14974);
nand UO_1268 (O_1268,N_14925,N_14972);
or UO_1269 (O_1269,N_14979,N_14960);
nor UO_1270 (O_1270,N_14994,N_14905);
xnor UO_1271 (O_1271,N_14895,N_14977);
or UO_1272 (O_1272,N_14895,N_14939);
xnor UO_1273 (O_1273,N_14913,N_14991);
nand UO_1274 (O_1274,N_14882,N_14927);
xor UO_1275 (O_1275,N_14881,N_14996);
or UO_1276 (O_1276,N_14982,N_14958);
or UO_1277 (O_1277,N_14981,N_14885);
or UO_1278 (O_1278,N_14985,N_14877);
nor UO_1279 (O_1279,N_14966,N_14988);
and UO_1280 (O_1280,N_14929,N_14958);
or UO_1281 (O_1281,N_14988,N_14947);
nor UO_1282 (O_1282,N_14922,N_14932);
nand UO_1283 (O_1283,N_14910,N_14947);
xnor UO_1284 (O_1284,N_14884,N_14964);
and UO_1285 (O_1285,N_14928,N_14893);
nor UO_1286 (O_1286,N_14916,N_14959);
nand UO_1287 (O_1287,N_14954,N_14956);
nor UO_1288 (O_1288,N_14950,N_14876);
nor UO_1289 (O_1289,N_14924,N_14911);
or UO_1290 (O_1290,N_14963,N_14899);
or UO_1291 (O_1291,N_14996,N_14964);
nor UO_1292 (O_1292,N_14936,N_14945);
and UO_1293 (O_1293,N_14895,N_14900);
or UO_1294 (O_1294,N_14970,N_14993);
nor UO_1295 (O_1295,N_14909,N_14889);
nand UO_1296 (O_1296,N_14901,N_14935);
and UO_1297 (O_1297,N_14998,N_14952);
nor UO_1298 (O_1298,N_14878,N_14979);
or UO_1299 (O_1299,N_14910,N_14891);
nand UO_1300 (O_1300,N_14946,N_14960);
or UO_1301 (O_1301,N_14946,N_14957);
and UO_1302 (O_1302,N_14941,N_14879);
xor UO_1303 (O_1303,N_14986,N_14999);
nand UO_1304 (O_1304,N_14899,N_14912);
nor UO_1305 (O_1305,N_14878,N_14936);
nand UO_1306 (O_1306,N_14986,N_14903);
and UO_1307 (O_1307,N_14978,N_14973);
nand UO_1308 (O_1308,N_14920,N_14950);
nand UO_1309 (O_1309,N_14977,N_14952);
nand UO_1310 (O_1310,N_14885,N_14909);
nor UO_1311 (O_1311,N_14894,N_14988);
and UO_1312 (O_1312,N_14974,N_14989);
nand UO_1313 (O_1313,N_14983,N_14924);
xor UO_1314 (O_1314,N_14996,N_14977);
and UO_1315 (O_1315,N_14927,N_14946);
or UO_1316 (O_1316,N_14963,N_14979);
xnor UO_1317 (O_1317,N_14982,N_14986);
and UO_1318 (O_1318,N_14899,N_14978);
nand UO_1319 (O_1319,N_14967,N_14993);
and UO_1320 (O_1320,N_14942,N_14949);
nor UO_1321 (O_1321,N_14941,N_14882);
or UO_1322 (O_1322,N_14909,N_14881);
or UO_1323 (O_1323,N_14994,N_14963);
or UO_1324 (O_1324,N_14964,N_14898);
nor UO_1325 (O_1325,N_14963,N_14977);
or UO_1326 (O_1326,N_14884,N_14941);
and UO_1327 (O_1327,N_14977,N_14933);
nand UO_1328 (O_1328,N_14886,N_14954);
and UO_1329 (O_1329,N_14983,N_14999);
and UO_1330 (O_1330,N_14886,N_14972);
or UO_1331 (O_1331,N_14933,N_14976);
nor UO_1332 (O_1332,N_14926,N_14920);
and UO_1333 (O_1333,N_14988,N_14878);
nand UO_1334 (O_1334,N_14941,N_14923);
or UO_1335 (O_1335,N_14909,N_14956);
nand UO_1336 (O_1336,N_14930,N_14978);
and UO_1337 (O_1337,N_14914,N_14885);
nor UO_1338 (O_1338,N_14924,N_14916);
nand UO_1339 (O_1339,N_14946,N_14948);
or UO_1340 (O_1340,N_14981,N_14999);
nor UO_1341 (O_1341,N_14894,N_14893);
xnor UO_1342 (O_1342,N_14918,N_14980);
xor UO_1343 (O_1343,N_14991,N_14989);
or UO_1344 (O_1344,N_14996,N_14978);
or UO_1345 (O_1345,N_14890,N_14995);
xor UO_1346 (O_1346,N_14994,N_14985);
xor UO_1347 (O_1347,N_14903,N_14960);
xnor UO_1348 (O_1348,N_14899,N_14906);
xnor UO_1349 (O_1349,N_14973,N_14997);
and UO_1350 (O_1350,N_14884,N_14888);
nor UO_1351 (O_1351,N_14882,N_14894);
nand UO_1352 (O_1352,N_14885,N_14953);
nor UO_1353 (O_1353,N_14987,N_14909);
xor UO_1354 (O_1354,N_14919,N_14988);
or UO_1355 (O_1355,N_14898,N_14893);
nor UO_1356 (O_1356,N_14959,N_14931);
nand UO_1357 (O_1357,N_14994,N_14880);
nand UO_1358 (O_1358,N_14952,N_14960);
xnor UO_1359 (O_1359,N_14967,N_14928);
and UO_1360 (O_1360,N_14942,N_14961);
or UO_1361 (O_1361,N_14949,N_14947);
nand UO_1362 (O_1362,N_14915,N_14940);
and UO_1363 (O_1363,N_14959,N_14927);
xor UO_1364 (O_1364,N_14916,N_14929);
nand UO_1365 (O_1365,N_14888,N_14992);
nand UO_1366 (O_1366,N_14990,N_14992);
nor UO_1367 (O_1367,N_14879,N_14921);
and UO_1368 (O_1368,N_14999,N_14902);
nand UO_1369 (O_1369,N_14935,N_14931);
xnor UO_1370 (O_1370,N_14976,N_14879);
nor UO_1371 (O_1371,N_14983,N_14943);
or UO_1372 (O_1372,N_14891,N_14961);
nand UO_1373 (O_1373,N_14889,N_14901);
and UO_1374 (O_1374,N_14961,N_14934);
xnor UO_1375 (O_1375,N_14888,N_14988);
and UO_1376 (O_1376,N_14890,N_14960);
and UO_1377 (O_1377,N_14882,N_14914);
and UO_1378 (O_1378,N_14945,N_14880);
and UO_1379 (O_1379,N_14967,N_14902);
nor UO_1380 (O_1380,N_14916,N_14995);
or UO_1381 (O_1381,N_14907,N_14894);
nor UO_1382 (O_1382,N_14928,N_14916);
and UO_1383 (O_1383,N_14942,N_14933);
nor UO_1384 (O_1384,N_14943,N_14946);
and UO_1385 (O_1385,N_14939,N_14932);
or UO_1386 (O_1386,N_14973,N_14930);
nor UO_1387 (O_1387,N_14945,N_14917);
nor UO_1388 (O_1388,N_14942,N_14978);
nand UO_1389 (O_1389,N_14998,N_14943);
and UO_1390 (O_1390,N_14988,N_14965);
and UO_1391 (O_1391,N_14907,N_14934);
xor UO_1392 (O_1392,N_14922,N_14971);
nor UO_1393 (O_1393,N_14886,N_14960);
or UO_1394 (O_1394,N_14972,N_14909);
nand UO_1395 (O_1395,N_14911,N_14958);
nand UO_1396 (O_1396,N_14979,N_14916);
and UO_1397 (O_1397,N_14984,N_14954);
nor UO_1398 (O_1398,N_14960,N_14934);
nor UO_1399 (O_1399,N_14981,N_14892);
and UO_1400 (O_1400,N_14976,N_14875);
nor UO_1401 (O_1401,N_14925,N_14992);
or UO_1402 (O_1402,N_14912,N_14903);
xnor UO_1403 (O_1403,N_14924,N_14927);
nand UO_1404 (O_1404,N_14876,N_14917);
xnor UO_1405 (O_1405,N_14900,N_14937);
nor UO_1406 (O_1406,N_14987,N_14914);
nand UO_1407 (O_1407,N_14945,N_14947);
nand UO_1408 (O_1408,N_14936,N_14987);
nand UO_1409 (O_1409,N_14991,N_14976);
nand UO_1410 (O_1410,N_14918,N_14979);
xnor UO_1411 (O_1411,N_14984,N_14941);
nor UO_1412 (O_1412,N_14896,N_14941);
or UO_1413 (O_1413,N_14958,N_14932);
nand UO_1414 (O_1414,N_14950,N_14886);
xor UO_1415 (O_1415,N_14983,N_14942);
or UO_1416 (O_1416,N_14973,N_14909);
nor UO_1417 (O_1417,N_14973,N_14960);
nand UO_1418 (O_1418,N_14894,N_14984);
nor UO_1419 (O_1419,N_14971,N_14918);
nand UO_1420 (O_1420,N_14969,N_14877);
or UO_1421 (O_1421,N_14999,N_14926);
and UO_1422 (O_1422,N_14969,N_14881);
or UO_1423 (O_1423,N_14927,N_14982);
nand UO_1424 (O_1424,N_14907,N_14981);
nor UO_1425 (O_1425,N_14887,N_14913);
or UO_1426 (O_1426,N_14932,N_14967);
nand UO_1427 (O_1427,N_14909,N_14896);
nand UO_1428 (O_1428,N_14965,N_14960);
nand UO_1429 (O_1429,N_14962,N_14930);
nand UO_1430 (O_1430,N_14890,N_14880);
and UO_1431 (O_1431,N_14958,N_14970);
and UO_1432 (O_1432,N_14956,N_14899);
nor UO_1433 (O_1433,N_14924,N_14938);
and UO_1434 (O_1434,N_14883,N_14996);
nand UO_1435 (O_1435,N_14968,N_14907);
xnor UO_1436 (O_1436,N_14885,N_14985);
nand UO_1437 (O_1437,N_14958,N_14992);
nand UO_1438 (O_1438,N_14991,N_14952);
nor UO_1439 (O_1439,N_14976,N_14923);
or UO_1440 (O_1440,N_14936,N_14891);
nand UO_1441 (O_1441,N_14917,N_14997);
nand UO_1442 (O_1442,N_14894,N_14989);
nor UO_1443 (O_1443,N_14946,N_14934);
or UO_1444 (O_1444,N_14878,N_14894);
nor UO_1445 (O_1445,N_14920,N_14931);
nand UO_1446 (O_1446,N_14894,N_14979);
and UO_1447 (O_1447,N_14887,N_14982);
xnor UO_1448 (O_1448,N_14918,N_14962);
nor UO_1449 (O_1449,N_14988,N_14882);
and UO_1450 (O_1450,N_14946,N_14986);
xnor UO_1451 (O_1451,N_14879,N_14876);
nor UO_1452 (O_1452,N_14907,N_14955);
and UO_1453 (O_1453,N_14879,N_14899);
or UO_1454 (O_1454,N_14917,N_14902);
nor UO_1455 (O_1455,N_14997,N_14970);
nor UO_1456 (O_1456,N_14970,N_14992);
or UO_1457 (O_1457,N_14946,N_14887);
and UO_1458 (O_1458,N_14987,N_14995);
and UO_1459 (O_1459,N_14896,N_14910);
and UO_1460 (O_1460,N_14921,N_14890);
xnor UO_1461 (O_1461,N_14951,N_14908);
and UO_1462 (O_1462,N_14959,N_14980);
nor UO_1463 (O_1463,N_14936,N_14993);
and UO_1464 (O_1464,N_14879,N_14956);
nand UO_1465 (O_1465,N_14943,N_14984);
xnor UO_1466 (O_1466,N_14995,N_14935);
nor UO_1467 (O_1467,N_14970,N_14937);
nor UO_1468 (O_1468,N_14974,N_14986);
xnor UO_1469 (O_1469,N_14934,N_14876);
and UO_1470 (O_1470,N_14893,N_14933);
nor UO_1471 (O_1471,N_14999,N_14923);
nor UO_1472 (O_1472,N_14877,N_14944);
nand UO_1473 (O_1473,N_14961,N_14993);
xnor UO_1474 (O_1474,N_14907,N_14903);
nand UO_1475 (O_1475,N_14963,N_14919);
and UO_1476 (O_1476,N_14940,N_14979);
nand UO_1477 (O_1477,N_14908,N_14991);
and UO_1478 (O_1478,N_14976,N_14977);
xor UO_1479 (O_1479,N_14890,N_14888);
or UO_1480 (O_1480,N_14973,N_14979);
nand UO_1481 (O_1481,N_14955,N_14979);
or UO_1482 (O_1482,N_14982,N_14897);
or UO_1483 (O_1483,N_14931,N_14927);
nand UO_1484 (O_1484,N_14890,N_14953);
or UO_1485 (O_1485,N_14928,N_14924);
nand UO_1486 (O_1486,N_14973,N_14959);
and UO_1487 (O_1487,N_14885,N_14889);
nor UO_1488 (O_1488,N_14884,N_14939);
nand UO_1489 (O_1489,N_14897,N_14972);
nor UO_1490 (O_1490,N_14895,N_14952);
and UO_1491 (O_1491,N_14894,N_14993);
xor UO_1492 (O_1492,N_14979,N_14949);
or UO_1493 (O_1493,N_14945,N_14892);
and UO_1494 (O_1494,N_14962,N_14932);
or UO_1495 (O_1495,N_14891,N_14895);
xnor UO_1496 (O_1496,N_14979,N_14926);
and UO_1497 (O_1497,N_14950,N_14925);
xor UO_1498 (O_1498,N_14995,N_14894);
nand UO_1499 (O_1499,N_14898,N_14971);
and UO_1500 (O_1500,N_14981,N_14989);
xor UO_1501 (O_1501,N_14880,N_14933);
nand UO_1502 (O_1502,N_14901,N_14907);
xnor UO_1503 (O_1503,N_14955,N_14893);
nor UO_1504 (O_1504,N_14983,N_14998);
nand UO_1505 (O_1505,N_14986,N_14994);
nor UO_1506 (O_1506,N_14895,N_14983);
or UO_1507 (O_1507,N_14893,N_14921);
nand UO_1508 (O_1508,N_14935,N_14907);
nand UO_1509 (O_1509,N_14963,N_14937);
nand UO_1510 (O_1510,N_14947,N_14993);
or UO_1511 (O_1511,N_14955,N_14897);
xor UO_1512 (O_1512,N_14918,N_14946);
nand UO_1513 (O_1513,N_14973,N_14972);
nor UO_1514 (O_1514,N_14994,N_14917);
nand UO_1515 (O_1515,N_14974,N_14927);
and UO_1516 (O_1516,N_14970,N_14887);
nand UO_1517 (O_1517,N_14932,N_14917);
nor UO_1518 (O_1518,N_14949,N_14912);
or UO_1519 (O_1519,N_14917,N_14937);
nor UO_1520 (O_1520,N_14911,N_14935);
nand UO_1521 (O_1521,N_14944,N_14893);
nand UO_1522 (O_1522,N_14985,N_14991);
and UO_1523 (O_1523,N_14948,N_14978);
and UO_1524 (O_1524,N_14890,N_14899);
and UO_1525 (O_1525,N_14972,N_14971);
xor UO_1526 (O_1526,N_14936,N_14915);
nand UO_1527 (O_1527,N_14889,N_14948);
nand UO_1528 (O_1528,N_14968,N_14953);
nor UO_1529 (O_1529,N_14925,N_14896);
nand UO_1530 (O_1530,N_14957,N_14906);
nand UO_1531 (O_1531,N_14971,N_14963);
nand UO_1532 (O_1532,N_14971,N_14959);
xor UO_1533 (O_1533,N_14911,N_14876);
xnor UO_1534 (O_1534,N_14885,N_14975);
nor UO_1535 (O_1535,N_14964,N_14878);
nand UO_1536 (O_1536,N_14980,N_14977);
nor UO_1537 (O_1537,N_14979,N_14905);
nor UO_1538 (O_1538,N_14968,N_14889);
nand UO_1539 (O_1539,N_14895,N_14917);
or UO_1540 (O_1540,N_14973,N_14983);
nor UO_1541 (O_1541,N_14991,N_14900);
nand UO_1542 (O_1542,N_14942,N_14943);
xor UO_1543 (O_1543,N_14989,N_14875);
nand UO_1544 (O_1544,N_14939,N_14999);
xnor UO_1545 (O_1545,N_14955,N_14931);
nor UO_1546 (O_1546,N_14904,N_14900);
or UO_1547 (O_1547,N_14876,N_14990);
xor UO_1548 (O_1548,N_14965,N_14883);
nand UO_1549 (O_1549,N_14961,N_14954);
and UO_1550 (O_1550,N_14975,N_14886);
nand UO_1551 (O_1551,N_14913,N_14931);
xor UO_1552 (O_1552,N_14904,N_14950);
nand UO_1553 (O_1553,N_14981,N_14995);
or UO_1554 (O_1554,N_14929,N_14985);
nand UO_1555 (O_1555,N_14960,N_14969);
nor UO_1556 (O_1556,N_14877,N_14932);
or UO_1557 (O_1557,N_14912,N_14926);
nor UO_1558 (O_1558,N_14953,N_14926);
or UO_1559 (O_1559,N_14996,N_14998);
nor UO_1560 (O_1560,N_14956,N_14993);
nor UO_1561 (O_1561,N_14890,N_14979);
or UO_1562 (O_1562,N_14951,N_14958);
and UO_1563 (O_1563,N_14967,N_14965);
xnor UO_1564 (O_1564,N_14993,N_14913);
and UO_1565 (O_1565,N_14990,N_14890);
and UO_1566 (O_1566,N_14948,N_14959);
nor UO_1567 (O_1567,N_14996,N_14892);
nor UO_1568 (O_1568,N_14997,N_14939);
nor UO_1569 (O_1569,N_14957,N_14916);
and UO_1570 (O_1570,N_14924,N_14980);
nor UO_1571 (O_1571,N_14897,N_14894);
nor UO_1572 (O_1572,N_14959,N_14964);
and UO_1573 (O_1573,N_14966,N_14970);
xnor UO_1574 (O_1574,N_14929,N_14906);
nand UO_1575 (O_1575,N_14949,N_14904);
nor UO_1576 (O_1576,N_14943,N_14893);
or UO_1577 (O_1577,N_14988,N_14953);
xnor UO_1578 (O_1578,N_14965,N_14926);
nand UO_1579 (O_1579,N_14981,N_14911);
xor UO_1580 (O_1580,N_14967,N_14974);
nor UO_1581 (O_1581,N_14901,N_14938);
xor UO_1582 (O_1582,N_14981,N_14943);
nand UO_1583 (O_1583,N_14876,N_14936);
xnor UO_1584 (O_1584,N_14910,N_14980);
xor UO_1585 (O_1585,N_14883,N_14944);
nand UO_1586 (O_1586,N_14903,N_14996);
nand UO_1587 (O_1587,N_14952,N_14942);
nor UO_1588 (O_1588,N_14941,N_14925);
and UO_1589 (O_1589,N_14908,N_14956);
and UO_1590 (O_1590,N_14986,N_14958);
xnor UO_1591 (O_1591,N_14905,N_14955);
nand UO_1592 (O_1592,N_14947,N_14978);
xnor UO_1593 (O_1593,N_14995,N_14915);
nor UO_1594 (O_1594,N_14921,N_14979);
xnor UO_1595 (O_1595,N_14897,N_14997);
and UO_1596 (O_1596,N_14915,N_14950);
nand UO_1597 (O_1597,N_14911,N_14985);
nand UO_1598 (O_1598,N_14939,N_14973);
or UO_1599 (O_1599,N_14973,N_14882);
and UO_1600 (O_1600,N_14908,N_14946);
and UO_1601 (O_1601,N_14995,N_14907);
xnor UO_1602 (O_1602,N_14903,N_14880);
nand UO_1603 (O_1603,N_14945,N_14928);
or UO_1604 (O_1604,N_14957,N_14963);
or UO_1605 (O_1605,N_14929,N_14882);
and UO_1606 (O_1606,N_14930,N_14917);
and UO_1607 (O_1607,N_14949,N_14944);
nand UO_1608 (O_1608,N_14892,N_14907);
and UO_1609 (O_1609,N_14978,N_14881);
nor UO_1610 (O_1610,N_14935,N_14973);
nand UO_1611 (O_1611,N_14876,N_14998);
nand UO_1612 (O_1612,N_14989,N_14978);
and UO_1613 (O_1613,N_14973,N_14982);
xnor UO_1614 (O_1614,N_14891,N_14886);
nand UO_1615 (O_1615,N_14998,N_14897);
and UO_1616 (O_1616,N_14961,N_14970);
or UO_1617 (O_1617,N_14912,N_14939);
nor UO_1618 (O_1618,N_14916,N_14989);
nor UO_1619 (O_1619,N_14947,N_14900);
xnor UO_1620 (O_1620,N_14933,N_14986);
nand UO_1621 (O_1621,N_14895,N_14927);
or UO_1622 (O_1622,N_14943,N_14918);
and UO_1623 (O_1623,N_14943,N_14965);
xor UO_1624 (O_1624,N_14889,N_14905);
nand UO_1625 (O_1625,N_14975,N_14876);
xnor UO_1626 (O_1626,N_14890,N_14893);
nor UO_1627 (O_1627,N_14909,N_14900);
xor UO_1628 (O_1628,N_14922,N_14913);
and UO_1629 (O_1629,N_14987,N_14952);
or UO_1630 (O_1630,N_14960,N_14910);
xor UO_1631 (O_1631,N_14923,N_14912);
nand UO_1632 (O_1632,N_14920,N_14877);
nor UO_1633 (O_1633,N_14949,N_14984);
or UO_1634 (O_1634,N_14956,N_14981);
or UO_1635 (O_1635,N_14979,N_14959);
xnor UO_1636 (O_1636,N_14921,N_14927);
nand UO_1637 (O_1637,N_14918,N_14917);
xnor UO_1638 (O_1638,N_14918,N_14975);
and UO_1639 (O_1639,N_14885,N_14924);
nor UO_1640 (O_1640,N_14942,N_14911);
xnor UO_1641 (O_1641,N_14993,N_14996);
nor UO_1642 (O_1642,N_14989,N_14892);
nor UO_1643 (O_1643,N_14938,N_14912);
xnor UO_1644 (O_1644,N_14945,N_14968);
nor UO_1645 (O_1645,N_14918,N_14942);
xor UO_1646 (O_1646,N_14948,N_14976);
and UO_1647 (O_1647,N_14984,N_14892);
nor UO_1648 (O_1648,N_14991,N_14997);
nand UO_1649 (O_1649,N_14988,N_14877);
xor UO_1650 (O_1650,N_14889,N_14908);
or UO_1651 (O_1651,N_14908,N_14884);
and UO_1652 (O_1652,N_14883,N_14969);
and UO_1653 (O_1653,N_14916,N_14960);
or UO_1654 (O_1654,N_14987,N_14879);
xnor UO_1655 (O_1655,N_14897,N_14912);
nand UO_1656 (O_1656,N_14939,N_14944);
xor UO_1657 (O_1657,N_14986,N_14978);
or UO_1658 (O_1658,N_14975,N_14982);
nand UO_1659 (O_1659,N_14927,N_14930);
nor UO_1660 (O_1660,N_14921,N_14886);
nor UO_1661 (O_1661,N_14989,N_14911);
and UO_1662 (O_1662,N_14937,N_14955);
nor UO_1663 (O_1663,N_14922,N_14978);
nor UO_1664 (O_1664,N_14875,N_14940);
nand UO_1665 (O_1665,N_14998,N_14887);
and UO_1666 (O_1666,N_14889,N_14984);
nor UO_1667 (O_1667,N_14917,N_14891);
and UO_1668 (O_1668,N_14952,N_14923);
xnor UO_1669 (O_1669,N_14941,N_14993);
xnor UO_1670 (O_1670,N_14960,N_14892);
nand UO_1671 (O_1671,N_14895,N_14947);
nand UO_1672 (O_1672,N_14980,N_14920);
nand UO_1673 (O_1673,N_14997,N_14965);
and UO_1674 (O_1674,N_14883,N_14908);
or UO_1675 (O_1675,N_14932,N_14887);
and UO_1676 (O_1676,N_14886,N_14912);
nor UO_1677 (O_1677,N_14958,N_14941);
nand UO_1678 (O_1678,N_14985,N_14876);
xnor UO_1679 (O_1679,N_14997,N_14967);
nand UO_1680 (O_1680,N_14878,N_14907);
or UO_1681 (O_1681,N_14927,N_14883);
xor UO_1682 (O_1682,N_14879,N_14994);
or UO_1683 (O_1683,N_14966,N_14994);
or UO_1684 (O_1684,N_14929,N_14876);
nor UO_1685 (O_1685,N_14954,N_14943);
xnor UO_1686 (O_1686,N_14916,N_14986);
nor UO_1687 (O_1687,N_14981,N_14986);
nor UO_1688 (O_1688,N_14959,N_14878);
or UO_1689 (O_1689,N_14915,N_14928);
or UO_1690 (O_1690,N_14899,N_14957);
xnor UO_1691 (O_1691,N_14884,N_14922);
and UO_1692 (O_1692,N_14937,N_14875);
xor UO_1693 (O_1693,N_14963,N_14984);
nand UO_1694 (O_1694,N_14992,N_14964);
xnor UO_1695 (O_1695,N_14900,N_14914);
or UO_1696 (O_1696,N_14908,N_14891);
nand UO_1697 (O_1697,N_14904,N_14951);
xor UO_1698 (O_1698,N_14931,N_14981);
nand UO_1699 (O_1699,N_14981,N_14973);
xor UO_1700 (O_1700,N_14920,N_14908);
or UO_1701 (O_1701,N_14987,N_14896);
xnor UO_1702 (O_1702,N_14973,N_14918);
and UO_1703 (O_1703,N_14901,N_14972);
or UO_1704 (O_1704,N_14919,N_14907);
and UO_1705 (O_1705,N_14963,N_14982);
or UO_1706 (O_1706,N_14970,N_14999);
xor UO_1707 (O_1707,N_14987,N_14948);
or UO_1708 (O_1708,N_14884,N_14892);
and UO_1709 (O_1709,N_14878,N_14995);
nand UO_1710 (O_1710,N_14944,N_14943);
nand UO_1711 (O_1711,N_14896,N_14905);
xnor UO_1712 (O_1712,N_14975,N_14924);
nand UO_1713 (O_1713,N_14987,N_14980);
nor UO_1714 (O_1714,N_14929,N_14889);
nor UO_1715 (O_1715,N_14936,N_14969);
and UO_1716 (O_1716,N_14969,N_14947);
and UO_1717 (O_1717,N_14935,N_14962);
nand UO_1718 (O_1718,N_14975,N_14959);
or UO_1719 (O_1719,N_14939,N_14966);
and UO_1720 (O_1720,N_14901,N_14957);
nor UO_1721 (O_1721,N_14929,N_14893);
nand UO_1722 (O_1722,N_14880,N_14925);
nand UO_1723 (O_1723,N_14901,N_14918);
nand UO_1724 (O_1724,N_14941,N_14898);
nand UO_1725 (O_1725,N_14948,N_14999);
nor UO_1726 (O_1726,N_14884,N_14875);
and UO_1727 (O_1727,N_14885,N_14921);
nand UO_1728 (O_1728,N_14904,N_14939);
and UO_1729 (O_1729,N_14992,N_14981);
nor UO_1730 (O_1730,N_14877,N_14923);
or UO_1731 (O_1731,N_14957,N_14979);
nand UO_1732 (O_1732,N_14984,N_14938);
or UO_1733 (O_1733,N_14935,N_14987);
xnor UO_1734 (O_1734,N_14995,N_14997);
xnor UO_1735 (O_1735,N_14922,N_14933);
xor UO_1736 (O_1736,N_14959,N_14903);
xor UO_1737 (O_1737,N_14979,N_14956);
and UO_1738 (O_1738,N_14943,N_14977);
xnor UO_1739 (O_1739,N_14992,N_14912);
or UO_1740 (O_1740,N_14990,N_14889);
xor UO_1741 (O_1741,N_14925,N_14987);
or UO_1742 (O_1742,N_14911,N_14944);
nand UO_1743 (O_1743,N_14936,N_14989);
nor UO_1744 (O_1744,N_14932,N_14891);
nand UO_1745 (O_1745,N_14976,N_14925);
or UO_1746 (O_1746,N_14958,N_14902);
nand UO_1747 (O_1747,N_14989,N_14990);
and UO_1748 (O_1748,N_14999,N_14968);
nand UO_1749 (O_1749,N_14914,N_14999);
and UO_1750 (O_1750,N_14882,N_14886);
nand UO_1751 (O_1751,N_14934,N_14989);
nand UO_1752 (O_1752,N_14953,N_14991);
or UO_1753 (O_1753,N_14953,N_14887);
or UO_1754 (O_1754,N_14982,N_14996);
and UO_1755 (O_1755,N_14907,N_14988);
xor UO_1756 (O_1756,N_14998,N_14958);
and UO_1757 (O_1757,N_14901,N_14961);
nand UO_1758 (O_1758,N_14918,N_14945);
or UO_1759 (O_1759,N_14984,N_14977);
nor UO_1760 (O_1760,N_14900,N_14883);
nand UO_1761 (O_1761,N_14985,N_14997);
xor UO_1762 (O_1762,N_14914,N_14884);
or UO_1763 (O_1763,N_14981,N_14944);
nor UO_1764 (O_1764,N_14927,N_14994);
xor UO_1765 (O_1765,N_14907,N_14942);
nand UO_1766 (O_1766,N_14956,N_14971);
xnor UO_1767 (O_1767,N_14955,N_14946);
and UO_1768 (O_1768,N_14889,N_14996);
nand UO_1769 (O_1769,N_14956,N_14922);
nand UO_1770 (O_1770,N_14896,N_14976);
nor UO_1771 (O_1771,N_14883,N_14879);
and UO_1772 (O_1772,N_14906,N_14888);
xnor UO_1773 (O_1773,N_14904,N_14893);
nor UO_1774 (O_1774,N_14914,N_14956);
xnor UO_1775 (O_1775,N_14977,N_14997);
or UO_1776 (O_1776,N_14881,N_14958);
nand UO_1777 (O_1777,N_14981,N_14939);
nand UO_1778 (O_1778,N_14884,N_14894);
nand UO_1779 (O_1779,N_14880,N_14997);
nand UO_1780 (O_1780,N_14916,N_14888);
and UO_1781 (O_1781,N_14974,N_14952);
and UO_1782 (O_1782,N_14983,N_14891);
or UO_1783 (O_1783,N_14895,N_14901);
nor UO_1784 (O_1784,N_14960,N_14985);
nor UO_1785 (O_1785,N_14976,N_14984);
nand UO_1786 (O_1786,N_14932,N_14976);
nor UO_1787 (O_1787,N_14944,N_14937);
and UO_1788 (O_1788,N_14909,N_14959);
or UO_1789 (O_1789,N_14950,N_14899);
and UO_1790 (O_1790,N_14986,N_14957);
and UO_1791 (O_1791,N_14965,N_14957);
xnor UO_1792 (O_1792,N_14976,N_14915);
xnor UO_1793 (O_1793,N_14936,N_14967);
or UO_1794 (O_1794,N_14927,N_14936);
and UO_1795 (O_1795,N_14880,N_14983);
nand UO_1796 (O_1796,N_14918,N_14951);
or UO_1797 (O_1797,N_14941,N_14981);
or UO_1798 (O_1798,N_14906,N_14978);
and UO_1799 (O_1799,N_14942,N_14936);
nand UO_1800 (O_1800,N_14933,N_14899);
nand UO_1801 (O_1801,N_14989,N_14982);
and UO_1802 (O_1802,N_14960,N_14925);
or UO_1803 (O_1803,N_14907,N_14908);
xnor UO_1804 (O_1804,N_14927,N_14887);
nand UO_1805 (O_1805,N_14997,N_14998);
nor UO_1806 (O_1806,N_14923,N_14969);
xor UO_1807 (O_1807,N_14914,N_14942);
nor UO_1808 (O_1808,N_14899,N_14984);
or UO_1809 (O_1809,N_14914,N_14973);
xnor UO_1810 (O_1810,N_14945,N_14951);
xor UO_1811 (O_1811,N_14978,N_14967);
nand UO_1812 (O_1812,N_14893,N_14990);
nor UO_1813 (O_1813,N_14986,N_14921);
or UO_1814 (O_1814,N_14977,N_14987);
and UO_1815 (O_1815,N_14982,N_14884);
nor UO_1816 (O_1816,N_14974,N_14976);
nor UO_1817 (O_1817,N_14891,N_14979);
nor UO_1818 (O_1818,N_14902,N_14891);
and UO_1819 (O_1819,N_14901,N_14971);
and UO_1820 (O_1820,N_14926,N_14917);
nor UO_1821 (O_1821,N_14915,N_14938);
nor UO_1822 (O_1822,N_14920,N_14988);
or UO_1823 (O_1823,N_14973,N_14922);
xor UO_1824 (O_1824,N_14976,N_14940);
and UO_1825 (O_1825,N_14884,N_14985);
nand UO_1826 (O_1826,N_14953,N_14877);
and UO_1827 (O_1827,N_14934,N_14974);
or UO_1828 (O_1828,N_14919,N_14891);
and UO_1829 (O_1829,N_14974,N_14892);
xor UO_1830 (O_1830,N_14982,N_14907);
nor UO_1831 (O_1831,N_14979,N_14994);
nand UO_1832 (O_1832,N_14968,N_14960);
xnor UO_1833 (O_1833,N_14926,N_14991);
nor UO_1834 (O_1834,N_14924,N_14968);
or UO_1835 (O_1835,N_14894,N_14881);
nor UO_1836 (O_1836,N_14905,N_14928);
and UO_1837 (O_1837,N_14938,N_14949);
or UO_1838 (O_1838,N_14879,N_14991);
xor UO_1839 (O_1839,N_14991,N_14938);
and UO_1840 (O_1840,N_14930,N_14932);
and UO_1841 (O_1841,N_14936,N_14889);
and UO_1842 (O_1842,N_14942,N_14932);
nor UO_1843 (O_1843,N_14930,N_14947);
and UO_1844 (O_1844,N_14889,N_14974);
nor UO_1845 (O_1845,N_14965,N_14902);
nand UO_1846 (O_1846,N_14885,N_14977);
xor UO_1847 (O_1847,N_14972,N_14889);
nor UO_1848 (O_1848,N_14915,N_14992);
nor UO_1849 (O_1849,N_14942,N_14976);
and UO_1850 (O_1850,N_14948,N_14887);
nor UO_1851 (O_1851,N_14891,N_14982);
xor UO_1852 (O_1852,N_14882,N_14897);
xnor UO_1853 (O_1853,N_14961,N_14913);
or UO_1854 (O_1854,N_14926,N_14972);
nand UO_1855 (O_1855,N_14980,N_14994);
and UO_1856 (O_1856,N_14899,N_14885);
nand UO_1857 (O_1857,N_14908,N_14937);
nand UO_1858 (O_1858,N_14894,N_14910);
or UO_1859 (O_1859,N_14939,N_14922);
or UO_1860 (O_1860,N_14927,N_14892);
or UO_1861 (O_1861,N_14880,N_14897);
nand UO_1862 (O_1862,N_14972,N_14922);
xnor UO_1863 (O_1863,N_14903,N_14995);
nor UO_1864 (O_1864,N_14936,N_14892);
and UO_1865 (O_1865,N_14879,N_14901);
nor UO_1866 (O_1866,N_14987,N_14979);
or UO_1867 (O_1867,N_14992,N_14985);
or UO_1868 (O_1868,N_14902,N_14911);
or UO_1869 (O_1869,N_14964,N_14902);
or UO_1870 (O_1870,N_14924,N_14921);
nand UO_1871 (O_1871,N_14969,N_14899);
xor UO_1872 (O_1872,N_14931,N_14914);
and UO_1873 (O_1873,N_14891,N_14954);
or UO_1874 (O_1874,N_14972,N_14979);
and UO_1875 (O_1875,N_14944,N_14930);
nand UO_1876 (O_1876,N_14991,N_14955);
or UO_1877 (O_1877,N_14989,N_14951);
xor UO_1878 (O_1878,N_14915,N_14956);
xnor UO_1879 (O_1879,N_14876,N_14956);
or UO_1880 (O_1880,N_14903,N_14935);
and UO_1881 (O_1881,N_14979,N_14902);
or UO_1882 (O_1882,N_14907,N_14881);
xor UO_1883 (O_1883,N_14914,N_14961);
and UO_1884 (O_1884,N_14903,N_14891);
nor UO_1885 (O_1885,N_14941,N_14935);
xor UO_1886 (O_1886,N_14934,N_14953);
or UO_1887 (O_1887,N_14990,N_14880);
xor UO_1888 (O_1888,N_14974,N_14913);
or UO_1889 (O_1889,N_14878,N_14961);
or UO_1890 (O_1890,N_14938,N_14934);
or UO_1891 (O_1891,N_14939,N_14889);
nand UO_1892 (O_1892,N_14951,N_14970);
and UO_1893 (O_1893,N_14966,N_14974);
and UO_1894 (O_1894,N_14876,N_14880);
nand UO_1895 (O_1895,N_14950,N_14878);
nor UO_1896 (O_1896,N_14951,N_14906);
xnor UO_1897 (O_1897,N_14956,N_14983);
nand UO_1898 (O_1898,N_14936,N_14905);
or UO_1899 (O_1899,N_14875,N_14915);
and UO_1900 (O_1900,N_14877,N_14915);
xnor UO_1901 (O_1901,N_14883,N_14968);
xnor UO_1902 (O_1902,N_14931,N_14893);
xor UO_1903 (O_1903,N_14995,N_14996);
and UO_1904 (O_1904,N_14976,N_14905);
nand UO_1905 (O_1905,N_14890,N_14935);
and UO_1906 (O_1906,N_14932,N_14968);
nand UO_1907 (O_1907,N_14990,N_14983);
nor UO_1908 (O_1908,N_14974,N_14920);
nand UO_1909 (O_1909,N_14914,N_14964);
xor UO_1910 (O_1910,N_14977,N_14897);
xor UO_1911 (O_1911,N_14903,N_14934);
nand UO_1912 (O_1912,N_14934,N_14887);
and UO_1913 (O_1913,N_14909,N_14946);
and UO_1914 (O_1914,N_14928,N_14939);
or UO_1915 (O_1915,N_14965,N_14887);
xor UO_1916 (O_1916,N_14922,N_14988);
nor UO_1917 (O_1917,N_14911,N_14941);
xor UO_1918 (O_1918,N_14964,N_14888);
xnor UO_1919 (O_1919,N_14877,N_14885);
nor UO_1920 (O_1920,N_14886,N_14919);
nand UO_1921 (O_1921,N_14959,N_14928);
or UO_1922 (O_1922,N_14904,N_14920);
xor UO_1923 (O_1923,N_14946,N_14950);
and UO_1924 (O_1924,N_14959,N_14891);
nor UO_1925 (O_1925,N_14960,N_14928);
xnor UO_1926 (O_1926,N_14921,N_14973);
nand UO_1927 (O_1927,N_14953,N_14902);
nand UO_1928 (O_1928,N_14891,N_14904);
nand UO_1929 (O_1929,N_14982,N_14953);
nand UO_1930 (O_1930,N_14960,N_14986);
nand UO_1931 (O_1931,N_14928,N_14913);
nor UO_1932 (O_1932,N_14900,N_14972);
or UO_1933 (O_1933,N_14924,N_14903);
nand UO_1934 (O_1934,N_14994,N_14887);
nand UO_1935 (O_1935,N_14938,N_14995);
xor UO_1936 (O_1936,N_14998,N_14942);
or UO_1937 (O_1937,N_14938,N_14877);
or UO_1938 (O_1938,N_14898,N_14912);
xor UO_1939 (O_1939,N_14913,N_14881);
or UO_1940 (O_1940,N_14878,N_14984);
or UO_1941 (O_1941,N_14957,N_14973);
xnor UO_1942 (O_1942,N_14886,N_14929);
xor UO_1943 (O_1943,N_14945,N_14972);
and UO_1944 (O_1944,N_14995,N_14887);
nor UO_1945 (O_1945,N_14885,N_14993);
or UO_1946 (O_1946,N_14956,N_14913);
nand UO_1947 (O_1947,N_14897,N_14996);
nor UO_1948 (O_1948,N_14970,N_14941);
and UO_1949 (O_1949,N_14894,N_14970);
and UO_1950 (O_1950,N_14900,N_14878);
xor UO_1951 (O_1951,N_14926,N_14880);
nor UO_1952 (O_1952,N_14881,N_14982);
and UO_1953 (O_1953,N_14917,N_14933);
xor UO_1954 (O_1954,N_14971,N_14910);
xnor UO_1955 (O_1955,N_14935,N_14893);
or UO_1956 (O_1956,N_14877,N_14936);
xnor UO_1957 (O_1957,N_14878,N_14886);
xor UO_1958 (O_1958,N_14961,N_14906);
or UO_1959 (O_1959,N_14967,N_14894);
nand UO_1960 (O_1960,N_14921,N_14896);
xnor UO_1961 (O_1961,N_14952,N_14903);
nor UO_1962 (O_1962,N_14973,N_14917);
xnor UO_1963 (O_1963,N_14970,N_14960);
or UO_1964 (O_1964,N_14960,N_14875);
or UO_1965 (O_1965,N_14902,N_14956);
nand UO_1966 (O_1966,N_14992,N_14960);
xor UO_1967 (O_1967,N_14940,N_14937);
nor UO_1968 (O_1968,N_14956,N_14941);
nand UO_1969 (O_1969,N_14961,N_14972);
or UO_1970 (O_1970,N_14992,N_14914);
xnor UO_1971 (O_1971,N_14972,N_14894);
and UO_1972 (O_1972,N_14956,N_14886);
nand UO_1973 (O_1973,N_14889,N_14940);
xnor UO_1974 (O_1974,N_14884,N_14886);
nor UO_1975 (O_1975,N_14936,N_14944);
or UO_1976 (O_1976,N_14902,N_14978);
nor UO_1977 (O_1977,N_14993,N_14962);
or UO_1978 (O_1978,N_14936,N_14966);
nand UO_1979 (O_1979,N_14907,N_14906);
and UO_1980 (O_1980,N_14964,N_14980);
or UO_1981 (O_1981,N_14981,N_14897);
and UO_1982 (O_1982,N_14888,N_14971);
and UO_1983 (O_1983,N_14927,N_14937);
nand UO_1984 (O_1984,N_14950,N_14935);
xnor UO_1985 (O_1985,N_14905,N_14906);
nand UO_1986 (O_1986,N_14887,N_14940);
nand UO_1987 (O_1987,N_14956,N_14878);
nor UO_1988 (O_1988,N_14956,N_14999);
xor UO_1989 (O_1989,N_14920,N_14934);
xor UO_1990 (O_1990,N_14879,N_14887);
nand UO_1991 (O_1991,N_14884,N_14977);
or UO_1992 (O_1992,N_14946,N_14891);
nand UO_1993 (O_1993,N_14902,N_14884);
xor UO_1994 (O_1994,N_14966,N_14881);
or UO_1995 (O_1995,N_14913,N_14890);
nor UO_1996 (O_1996,N_14944,N_14885);
and UO_1997 (O_1997,N_14911,N_14886);
and UO_1998 (O_1998,N_14888,N_14895);
nor UO_1999 (O_1999,N_14930,N_14986);
endmodule