module basic_1500_15000_2000_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_735,In_26);
and U1 (N_1,In_1238,In_55);
nor U2 (N_2,In_1145,In_1296);
nand U3 (N_3,In_350,In_587);
and U4 (N_4,In_383,In_1229);
nand U5 (N_5,In_1192,In_1073);
nor U6 (N_6,In_1117,In_1181);
or U7 (N_7,In_1118,In_954);
and U8 (N_8,In_335,In_1363);
nand U9 (N_9,In_82,In_1388);
nand U10 (N_10,In_1412,In_4);
nor U11 (N_11,In_1271,In_1315);
nand U12 (N_12,In_1276,In_1307);
nand U13 (N_13,In_892,In_649);
or U14 (N_14,In_314,In_529);
nor U15 (N_15,In_879,In_1202);
nor U16 (N_16,In_296,In_102);
or U17 (N_17,In_536,In_949);
or U18 (N_18,In_760,In_1341);
and U19 (N_19,In_1480,In_1407);
or U20 (N_20,In_1380,In_109);
or U21 (N_21,In_840,In_280);
and U22 (N_22,In_198,In_500);
or U23 (N_23,In_885,In_347);
or U24 (N_24,In_1185,In_514);
nand U25 (N_25,In_256,In_1490);
or U26 (N_26,In_1343,In_1213);
nand U27 (N_27,In_693,In_681);
nand U28 (N_28,In_983,In_1175);
xnor U29 (N_29,In_826,In_343);
nor U30 (N_30,In_240,In_763);
nand U31 (N_31,In_39,In_20);
xor U32 (N_32,In_1066,In_37);
nand U33 (N_33,In_268,In_245);
nand U34 (N_34,In_1030,In_1089);
or U35 (N_35,In_50,In_339);
nor U36 (N_36,In_481,In_61);
or U37 (N_37,In_1329,In_1237);
and U38 (N_38,In_1045,In_1136);
nor U39 (N_39,In_848,In_601);
nor U40 (N_40,In_938,In_1186);
xor U41 (N_41,In_784,In_616);
and U42 (N_42,In_59,In_658);
nor U43 (N_43,In_83,In_535);
and U44 (N_44,In_72,In_93);
nor U45 (N_45,In_537,In_700);
and U46 (N_46,In_1312,In_521);
or U47 (N_47,In_422,In_1035);
or U48 (N_48,In_292,In_984);
and U49 (N_49,In_12,In_1413);
nor U50 (N_50,In_348,In_642);
or U51 (N_51,In_51,In_1494);
nand U52 (N_52,In_842,In_151);
nor U53 (N_53,In_270,In_837);
or U54 (N_54,In_66,In_979);
and U55 (N_55,In_1024,In_1221);
and U56 (N_56,In_701,In_1308);
nand U57 (N_57,In_413,In_1448);
and U58 (N_58,In_836,In_959);
nor U59 (N_59,In_1377,In_193);
xor U60 (N_60,In_723,In_1460);
and U61 (N_61,In_850,In_1200);
or U62 (N_62,In_1242,In_556);
xnor U63 (N_63,In_303,In_708);
and U64 (N_64,In_139,In_399);
and U65 (N_65,In_71,In_94);
and U66 (N_66,In_163,In_632);
nand U67 (N_67,In_695,In_942);
or U68 (N_68,In_756,In_1114);
nand U69 (N_69,In_77,In_369);
xor U70 (N_70,In_175,In_57);
nand U71 (N_71,In_775,In_79);
nand U72 (N_72,In_310,In_386);
or U73 (N_73,In_1195,In_778);
or U74 (N_74,In_48,In_747);
nor U75 (N_75,In_1043,In_306);
nand U76 (N_76,In_1029,In_578);
xor U77 (N_77,In_1106,In_458);
and U78 (N_78,In_1067,In_177);
nand U79 (N_79,In_1058,In_1498);
nor U80 (N_80,In_277,In_1457);
nor U81 (N_81,In_844,In_107);
or U82 (N_82,In_2,In_581);
nor U83 (N_83,In_619,In_190);
and U84 (N_84,In_418,In_319);
nor U85 (N_85,In_945,In_1027);
xnor U86 (N_86,In_1087,In_569);
xor U87 (N_87,In_1172,In_1132);
and U88 (N_88,In_243,In_185);
and U89 (N_89,In_97,In_473);
nand U90 (N_90,In_337,In_1396);
nand U91 (N_91,In_1151,In_773);
or U92 (N_92,In_871,In_1168);
nor U93 (N_93,In_1023,In_489);
and U94 (N_94,In_30,In_441);
and U95 (N_95,In_1431,In_446);
and U96 (N_96,In_751,In_1421);
nand U97 (N_97,In_611,In_122);
nand U98 (N_98,In_603,In_35);
and U99 (N_99,In_135,In_255);
nor U100 (N_100,In_986,In_889);
or U101 (N_101,In_1302,In_870);
and U102 (N_102,In_1109,In_1240);
nor U103 (N_103,In_389,In_491);
xor U104 (N_104,In_921,In_1466);
or U105 (N_105,In_15,In_668);
or U106 (N_106,In_819,In_65);
and U107 (N_107,In_1107,In_1336);
or U108 (N_108,In_1373,In_6);
and U109 (N_109,In_351,In_1096);
and U110 (N_110,In_948,In_437);
or U111 (N_111,In_503,In_325);
xnor U112 (N_112,In_430,In_798);
nand U113 (N_113,In_400,In_1228);
or U114 (N_114,In_638,In_110);
or U115 (N_115,In_972,In_1463);
or U116 (N_116,In_1046,In_880);
or U117 (N_117,In_1054,In_299);
nand U118 (N_118,In_1327,In_406);
and U119 (N_119,In_757,In_199);
nor U120 (N_120,In_1320,In_542);
nor U121 (N_121,In_652,In_762);
or U122 (N_122,In_1004,In_239);
and U123 (N_123,In_410,In_1316);
nor U124 (N_124,In_125,In_660);
nand U125 (N_125,In_1311,In_13);
or U126 (N_126,In_704,In_1454);
or U127 (N_127,In_516,In_847);
and U128 (N_128,In_1153,In_40);
nor U129 (N_129,In_706,In_165);
and U130 (N_130,In_1301,In_1386);
nor U131 (N_131,In_1447,In_1039);
and U132 (N_132,In_1275,In_1305);
nand U133 (N_133,In_1338,In_133);
and U134 (N_134,In_770,In_168);
nor U135 (N_135,In_1436,In_88);
nor U136 (N_136,In_877,In_1420);
and U137 (N_137,In_962,In_1376);
xnor U138 (N_138,In_633,In_643);
xnor U139 (N_139,In_250,In_1108);
or U140 (N_140,In_242,In_45);
and U141 (N_141,In_63,In_1155);
nand U142 (N_142,In_338,In_408);
or U143 (N_143,In_1279,In_261);
or U144 (N_144,In_235,In_1357);
and U145 (N_145,In_554,In_228);
nor U146 (N_146,In_573,In_1188);
nand U147 (N_147,In_448,In_1414);
and U148 (N_148,In_1293,In_251);
nand U149 (N_149,In_381,In_140);
or U150 (N_150,In_461,In_209);
nand U151 (N_151,In_1492,In_462);
or U152 (N_152,In_999,In_327);
and U153 (N_153,In_597,In_1263);
xnor U154 (N_154,In_1351,In_1299);
xor U155 (N_155,In_810,In_46);
nand U156 (N_156,In_1286,In_1430);
or U157 (N_157,In_951,In_1093);
or U158 (N_158,In_1283,In_526);
or U159 (N_159,In_614,In_1306);
nor U160 (N_160,In_1050,In_356);
nand U161 (N_161,In_395,In_568);
nand U162 (N_162,In_1324,In_1201);
or U163 (N_163,In_767,In_657);
and U164 (N_164,In_176,In_1481);
nor U165 (N_165,In_1167,In_1383);
nor U166 (N_166,In_1321,In_85);
and U167 (N_167,In_25,In_923);
or U168 (N_168,In_532,In_577);
or U169 (N_169,In_81,In_676);
xnor U170 (N_170,In_21,In_1261);
nor U171 (N_171,In_101,In_715);
nand U172 (N_172,In_853,In_1002);
or U173 (N_173,In_260,In_815);
or U174 (N_174,In_1170,In_953);
nor U175 (N_175,In_662,In_1297);
nand U176 (N_176,In_812,In_27);
and U177 (N_177,In_904,In_1455);
and U178 (N_178,In_147,In_1422);
and U179 (N_179,In_182,In_127);
and U180 (N_180,In_470,In_765);
nand U181 (N_181,In_645,In_987);
and U182 (N_182,In_1162,In_162);
nor U183 (N_183,In_204,In_1346);
nand U184 (N_184,In_1354,In_103);
nor U185 (N_185,In_692,In_113);
or U186 (N_186,In_709,In_307);
nor U187 (N_187,In_131,In_317);
nor U188 (N_188,In_1203,In_1469);
and U189 (N_189,In_142,In_754);
nand U190 (N_190,In_687,In_468);
nor U191 (N_191,In_1074,In_803);
and U192 (N_192,In_124,In_75);
nor U193 (N_193,In_1291,In_533);
nor U194 (N_194,In_1465,In_490);
and U195 (N_195,In_690,In_293);
or U196 (N_196,In_370,In_884);
or U197 (N_197,In_648,In_563);
or U198 (N_198,In_1482,In_1154);
or U199 (N_199,In_946,In_750);
and U200 (N_200,In_1124,In_673);
nand U201 (N_201,In_192,In_89);
or U202 (N_202,In_1269,In_346);
or U203 (N_203,In_1082,In_1216);
and U204 (N_204,In_1129,In_822);
and U205 (N_205,In_1251,In_1233);
nor U206 (N_206,In_939,In_721);
and U207 (N_207,In_1205,In_380);
and U208 (N_208,In_733,In_1125);
and U209 (N_209,In_934,In_625);
or U210 (N_210,In_1011,In_213);
and U211 (N_211,In_859,In_740);
nand U212 (N_212,In_1187,In_76);
nand U213 (N_213,In_1222,In_1049);
or U214 (N_214,In_126,In_629);
and U215 (N_215,In_864,In_119);
or U216 (N_216,In_180,In_1470);
or U217 (N_217,In_820,In_1028);
and U218 (N_218,In_19,In_1111);
nand U219 (N_219,In_1405,In_41);
nand U220 (N_220,In_404,In_206);
nor U221 (N_221,In_1253,In_1101);
nor U222 (N_222,In_1174,In_1478);
nand U223 (N_223,In_912,In_774);
nand U224 (N_224,In_1184,In_1347);
xnor U225 (N_225,In_804,In_166);
or U226 (N_226,In_1331,In_759);
or U227 (N_227,In_34,In_791);
or U228 (N_228,In_928,In_828);
or U229 (N_229,In_1178,In_605);
xor U230 (N_230,In_531,In_663);
or U231 (N_231,In_367,In_62);
nand U232 (N_232,In_752,In_910);
or U233 (N_233,In_1191,In_1404);
nand U234 (N_234,In_149,In_1435);
xor U235 (N_235,In_69,In_888);
xor U236 (N_236,In_933,In_724);
nor U237 (N_237,In_1356,In_996);
xnor U238 (N_238,In_358,In_1183);
or U239 (N_239,In_1243,In_1382);
nand U240 (N_240,In_179,In_1223);
and U241 (N_241,In_29,In_785);
and U242 (N_242,In_1057,In_506);
and U243 (N_243,In_8,In_373);
or U244 (N_244,In_699,In_186);
nor U245 (N_245,In_322,In_585);
nand U246 (N_246,In_431,In_402);
or U247 (N_247,In_513,In_445);
nor U248 (N_248,In_111,In_697);
nand U249 (N_249,In_710,In_1437);
nor U250 (N_250,In_1209,In_311);
and U251 (N_251,In_218,In_1370);
and U252 (N_252,In_78,In_716);
nor U253 (N_253,In_1393,In_5);
nand U254 (N_254,In_493,In_608);
nor U255 (N_255,In_550,In_167);
nand U256 (N_256,In_1387,In_230);
nor U257 (N_257,In_1314,In_324);
xnor U258 (N_258,In_1462,In_1163);
or U259 (N_259,In_153,In_1110);
and U260 (N_260,In_18,In_1016);
or U261 (N_261,In_839,In_510);
nand U262 (N_262,In_36,In_1353);
and U263 (N_263,In_1068,In_450);
or U264 (N_264,In_1130,In_372);
xnor U265 (N_265,In_1384,In_1197);
nand U266 (N_266,In_1339,In_301);
nor U267 (N_267,In_1403,In_128);
xnor U268 (N_268,In_492,In_1098);
and U269 (N_269,In_420,In_1337);
nand U270 (N_270,In_1070,In_595);
nor U271 (N_271,In_401,In_1031);
xnor U272 (N_272,In_416,In_435);
nor U273 (N_273,In_1411,In_686);
xnor U274 (N_274,In_618,In_141);
nand U275 (N_275,In_897,In_637);
nor U276 (N_276,In_621,In_164);
nand U277 (N_277,In_300,In_439);
nand U278 (N_278,In_225,In_1491);
and U279 (N_279,In_202,In_1428);
nand U280 (N_280,In_743,In_120);
nand U281 (N_281,In_460,In_831);
nand U282 (N_282,In_817,In_958);
nor U283 (N_283,In_1140,In_860);
xnor U284 (N_284,In_748,In_970);
nor U285 (N_285,In_985,In_591);
nand U286 (N_286,In_992,In_375);
and U287 (N_287,In_42,In_1062);
or U288 (N_288,In_308,In_1149);
nor U289 (N_289,In_411,In_1217);
or U290 (N_290,In_387,In_1059);
and U291 (N_291,In_1449,In_998);
nand U292 (N_292,In_1325,In_1450);
and U293 (N_293,In_434,In_886);
nor U294 (N_294,In_1080,In_572);
nand U295 (N_295,In_624,In_866);
or U296 (N_296,In_421,In_1257);
xor U297 (N_297,In_1126,In_630);
xor U298 (N_298,In_613,In_792);
and U299 (N_299,In_7,In_800);
nor U300 (N_300,In_466,In_366);
and U301 (N_301,In_1018,In_155);
and U302 (N_302,In_957,In_607);
nand U303 (N_303,In_1210,In_1452);
or U304 (N_304,In_43,In_1434);
or U305 (N_305,In_1289,In_1020);
or U306 (N_306,In_1441,In_916);
nand U307 (N_307,In_795,In_1378);
nor U308 (N_308,In_474,In_74);
nor U309 (N_309,In_1423,In_302);
xor U310 (N_310,In_734,In_1340);
nor U311 (N_311,In_1092,In_1485);
xor U312 (N_312,In_252,In_32);
nor U313 (N_313,In_565,In_1319);
nand U314 (N_314,In_806,In_31);
or U315 (N_315,In_644,In_797);
and U316 (N_316,In_379,In_60);
and U317 (N_317,In_53,In_1365);
or U318 (N_318,In_1123,In_736);
nand U319 (N_319,In_1268,In_719);
xnor U320 (N_320,In_671,In_1474);
nand U321 (N_321,In_249,In_11);
nand U322 (N_322,In_289,In_87);
or U323 (N_323,In_496,In_1091);
nand U324 (N_324,In_1300,In_1446);
xor U325 (N_325,In_626,In_173);
nor U326 (N_326,In_407,In_830);
and U327 (N_327,In_99,In_1352);
and U328 (N_328,In_712,In_691);
nand U329 (N_329,In_382,In_940);
nor U330 (N_330,In_849,In_392);
and U331 (N_331,In_598,In_1199);
and U332 (N_332,In_17,In_920);
or U333 (N_333,In_1310,In_1146);
and U334 (N_334,In_725,In_452);
nand U335 (N_335,In_475,In_1047);
xnor U336 (N_336,In_1052,In_323);
and U337 (N_337,In_1360,In_882);
nand U338 (N_338,In_899,In_443);
xor U339 (N_339,In_544,In_472);
nand U340 (N_340,In_1071,In_1471);
and U341 (N_341,In_1424,In_1156);
and U342 (N_342,In_856,In_620);
and U343 (N_343,In_753,In_941);
xnor U344 (N_344,In_196,In_1158);
xor U345 (N_345,In_1040,In_1194);
xnor U346 (N_346,In_248,In_1139);
or U347 (N_347,In_465,In_226);
xnor U348 (N_348,In_900,In_482);
or U349 (N_349,In_426,In_584);
and U350 (N_350,In_220,In_403);
nor U351 (N_351,In_1081,In_950);
nand U352 (N_352,In_772,In_1397);
nor U353 (N_353,In_272,In_234);
xor U354 (N_354,In_570,In_157);
nand U355 (N_355,In_1493,In_1069);
nand U356 (N_356,In_1444,In_172);
and U357 (N_357,In_1053,In_424);
nor U358 (N_358,In_203,In_1193);
xnor U359 (N_359,In_1190,In_685);
or U360 (N_360,In_639,In_227);
or U361 (N_361,In_1225,In_1484);
nor U362 (N_362,In_1204,In_610);
nand U363 (N_363,In_749,In_636);
or U364 (N_364,In_1177,In_1100);
nor U365 (N_365,In_205,In_183);
and U366 (N_366,In_484,In_276);
nand U367 (N_367,In_476,In_766);
xnor U368 (N_368,In_1165,In_508);
nor U369 (N_369,In_340,In_91);
and U370 (N_370,In_720,In_23);
and U371 (N_371,In_534,In_394);
or U372 (N_372,In_478,In_698);
xor U373 (N_373,In_1415,In_44);
nor U374 (N_374,In_653,In_786);
nand U375 (N_375,In_1406,In_485);
nand U376 (N_376,In_377,In_16);
nor U377 (N_377,In_661,In_1206);
and U378 (N_378,In_1280,In_253);
nand U379 (N_379,In_486,In_872);
or U380 (N_380,In_540,In_1473);
xnor U381 (N_381,In_927,In_852);
and U382 (N_382,In_359,In_560);
nor U383 (N_383,In_197,In_782);
and U384 (N_384,In_412,In_1281);
or U385 (N_385,In_357,In_1008);
or U386 (N_386,In_1044,In_543);
xnor U387 (N_387,In_664,In_1133);
nand U388 (N_388,In_305,In_425);
xnor U389 (N_389,In_1017,In_669);
nor U390 (N_390,In_932,In_236);
or U391 (N_391,In_1259,In_1385);
nand U392 (N_392,In_429,In_640);
and U393 (N_393,In_391,In_780);
xnor U394 (N_394,In_1247,In_841);
xor U395 (N_395,In_689,In_915);
nor U396 (N_396,In_935,In_855);
nand U397 (N_397,In_1218,In_705);
nor U398 (N_398,In_397,In_1234);
nor U399 (N_399,In_455,In_1064);
and U400 (N_400,In_237,In_1267);
nand U401 (N_401,In_918,In_924);
nand U402 (N_402,In_159,In_262);
nor U403 (N_403,In_442,In_344);
xnor U404 (N_404,In_1256,In_1230);
or U405 (N_405,In_680,In_887);
or U406 (N_406,In_1390,In_364);
and U407 (N_407,In_257,In_1105);
or U408 (N_408,In_315,In_890);
and U409 (N_409,In_114,In_136);
nand U410 (N_410,In_264,In_771);
nand U411 (N_411,In_1304,In_1400);
nand U412 (N_412,In_28,In_602);
nor U413 (N_413,In_214,In_878);
and U414 (N_414,In_1120,In_432);
nor U415 (N_415,In_744,In_738);
nand U416 (N_416,In_145,In_599);
xnor U417 (N_417,In_1147,In_741);
xor U418 (N_418,In_487,In_854);
nand U419 (N_419,In_862,In_453);
nor U420 (N_420,In_1119,In_558);
and U421 (N_421,In_1032,In_1014);
or U422 (N_422,In_1467,In_726);
and U423 (N_423,In_1115,In_1138);
or U424 (N_424,In_594,In_1274);
nand U425 (N_425,In_1468,In_769);
or U426 (N_426,In_201,In_1313);
nor U427 (N_427,In_298,In_143);
nand U428 (N_428,In_283,In_994);
nand U429 (N_429,In_3,In_524);
nand U430 (N_430,In_318,In_952);
or U431 (N_431,In_1323,In_330);
and U432 (N_432,In_582,In_717);
nand U433 (N_433,In_419,In_118);
nor U434 (N_434,In_1292,In_758);
nand U435 (N_435,In_409,In_1401);
nor U436 (N_436,In_1497,In_1128);
nor U437 (N_437,In_378,In_520);
and U438 (N_438,In_1359,In_90);
nor U439 (N_439,In_64,In_851);
nor U440 (N_440,In_1037,In_336);
and U441 (N_441,In_352,In_1322);
nor U442 (N_442,In_857,In_805);
and U443 (N_443,In_1159,In_263);
nand U444 (N_444,In_1246,In_95);
nand U445 (N_445,In_231,In_1161);
or U446 (N_446,In_223,In_0);
xor U447 (N_447,In_682,In_1427);
or U448 (N_448,In_808,In_522);
and U449 (N_449,In_907,In_278);
nor U450 (N_450,In_471,In_108);
nor U451 (N_451,In_233,In_84);
and U452 (N_452,In_1451,In_1318);
and U453 (N_453,In_615,In_788);
and U454 (N_454,In_802,In_654);
xor U455 (N_455,In_1013,In_789);
nor U456 (N_456,In_1344,In_567);
and U457 (N_457,In_909,In_216);
nand U458 (N_458,In_1285,In_1094);
nand U459 (N_459,In_1355,In_33);
nand U460 (N_460,In_703,In_1425);
nand U461 (N_461,In_829,In_1226);
and U462 (N_462,In_247,In_144);
nand U463 (N_463,In_670,In_221);
xor U464 (N_464,In_1076,In_894);
and U465 (N_465,In_1127,In_282);
xnor U466 (N_466,In_1372,In_1489);
nand U467 (N_467,In_553,In_666);
nor U468 (N_468,In_254,In_683);
and U469 (N_469,In_1260,In_345);
nand U470 (N_470,In_1438,In_1394);
nor U471 (N_471,In_92,In_755);
or U472 (N_472,In_641,In_447);
and U473 (N_473,In_1368,In_169);
and U474 (N_474,In_1248,In_415);
or U475 (N_475,In_963,In_1214);
nand U476 (N_476,In_547,In_729);
and U477 (N_477,In_320,In_184);
nand U478 (N_478,In_742,In_596);
or U479 (N_479,In_627,In_480);
nand U480 (N_480,In_1456,In_794);
nor U481 (N_481,In_498,In_1148);
xnor U482 (N_482,In_931,In_875);
nand U483 (N_483,In_222,In_354);
and U484 (N_484,In_969,In_1266);
and U485 (N_485,In_47,In_1345);
nor U486 (N_486,In_628,In_722);
nand U487 (N_487,In_1180,In_188);
and U488 (N_488,In_1409,In_1171);
nand U489 (N_489,In_174,In_655);
and U490 (N_490,In_288,In_1298);
and U491 (N_491,In_604,In_647);
nor U492 (N_492,In_811,In_1398);
nand U493 (N_493,In_1121,In_1141);
nor U494 (N_494,In_210,In_1088);
or U495 (N_495,In_1055,In_291);
nor U496 (N_496,In_1348,In_1065);
nor U497 (N_497,In_355,In_1410);
and U498 (N_498,In_809,In_1288);
or U499 (N_499,In_943,In_1164);
xnor U500 (N_500,In_1330,In_1399);
nand U501 (N_501,In_1075,In_694);
and U502 (N_502,In_363,In_1479);
and U503 (N_503,In_1056,In_1290);
nor U504 (N_504,In_1264,In_956);
xor U505 (N_505,In_1418,In_814);
nor U506 (N_506,In_1294,In_49);
nor U507 (N_507,In_1116,In_1231);
and U508 (N_508,In_799,In_86);
nor U509 (N_509,In_600,In_371);
and U510 (N_510,In_714,In_617);
xor U511 (N_511,In_813,In_267);
nor U512 (N_512,In_1025,In_341);
nand U513 (N_513,In_398,In_665);
and U514 (N_514,In_589,In_549);
xor U515 (N_515,In_1371,In_718);
nor U516 (N_516,In_846,In_982);
and U517 (N_517,In_1287,In_361);
or U518 (N_518,In_1440,In_1085);
nand U519 (N_519,In_152,In_971);
nor U520 (N_520,In_1072,In_181);
and U521 (N_521,In_1102,In_1235);
and U522 (N_522,In_1278,In_509);
and U523 (N_523,In_1332,In_459);
xnor U524 (N_524,In_967,In_1113);
nor U525 (N_525,In_316,In_1254);
nand U526 (N_526,In_362,In_1000);
or U527 (N_527,In_1367,In_1015);
nand U528 (N_528,In_388,In_961);
or U529 (N_529,In_279,In_1169);
nand U530 (N_530,In_538,In_977);
nand U531 (N_531,In_739,In_1220);
nor U532 (N_532,In_672,In_883);
nor U533 (N_533,In_779,In_494);
and U534 (N_534,In_334,In_150);
nor U535 (N_535,In_1429,In_385);
and U536 (N_536,In_1086,In_586);
xor U537 (N_537,In_469,In_936);
nand U538 (N_538,In_821,In_530);
nor U539 (N_539,In_194,In_457);
or U540 (N_540,In_874,In_833);
nor U541 (N_541,In_1084,In_414);
or U542 (N_542,In_911,In_917);
nand U543 (N_543,In_650,In_592);
or U544 (N_544,In_132,In_390);
nor U545 (N_545,In_1245,In_793);
nor U546 (N_546,In_1104,In_38);
nand U547 (N_547,In_1364,In_1142);
nor U548 (N_548,In_273,In_105);
xor U549 (N_549,In_906,In_449);
nor U550 (N_550,In_1464,In_161);
xor U551 (N_551,In_130,In_635);
or U552 (N_552,In_1137,In_552);
nor U553 (N_553,In_483,In_1361);
or U554 (N_554,In_68,In_579);
or U555 (N_555,In_464,In_304);
nor U556 (N_556,In_895,In_9);
and U557 (N_557,In_1001,In_137);
nor U558 (N_558,In_1038,In_1090);
or U559 (N_559,In_436,In_488);
nor U560 (N_560,In_104,In_259);
nor U561 (N_561,In_1476,In_965);
nand U562 (N_562,In_593,In_1157);
nor U563 (N_563,In_1282,In_1212);
or U564 (N_564,In_905,In_1144);
or U565 (N_565,In_286,In_1182);
or U566 (N_566,In_777,In_284);
or U567 (N_567,In_801,In_1442);
nand U568 (N_568,In_746,In_555);
xor U569 (N_569,In_171,In_1265);
and U570 (N_570,In_22,In_56);
nor U571 (N_571,In_1369,In_290);
or U572 (N_572,In_1374,In_768);
xnor U573 (N_573,In_903,In_1349);
nand U574 (N_574,In_713,In_67);
nor U575 (N_575,In_1006,In_1196);
nand U576 (N_576,In_1458,In_858);
nand U577 (N_577,In_745,In_24);
or U578 (N_578,In_1342,In_764);
and U579 (N_579,In_1262,In_332);
nand U580 (N_580,In_1309,In_1);
nor U581 (N_581,In_1026,In_1152);
nor U582 (N_582,In_978,In_501);
or U583 (N_583,In_1487,In_189);
or U584 (N_584,In_207,In_1009);
or U585 (N_585,In_988,In_991);
and U586 (N_586,In_269,In_148);
nor U587 (N_587,In_454,In_14);
and U588 (N_588,In_384,In_1019);
nor U589 (N_589,In_834,In_576);
and U590 (N_590,In_557,In_1475);
and U591 (N_591,In_783,In_1362);
and U592 (N_592,In_590,In_898);
nor U593 (N_593,In_134,In_1402);
xor U594 (N_594,In_1326,In_732);
nand U595 (N_595,In_559,In_981);
and U596 (N_596,In_1379,In_881);
or U597 (N_597,In_54,In_1483);
or U598 (N_598,In_326,In_1443);
and U599 (N_599,In_219,In_728);
and U600 (N_600,In_497,In_571);
and U601 (N_601,In_1303,In_365);
and U602 (N_602,In_1079,In_224);
or U603 (N_603,In_1005,In_467);
nor U604 (N_604,In_634,In_930);
nor U605 (N_605,In_1496,In_845);
nor U606 (N_606,In_274,In_1208);
nand U607 (N_607,In_376,In_511);
or U608 (N_608,In_902,In_1083);
nor U609 (N_609,In_495,In_499);
nand U610 (N_610,In_1461,In_937);
nor U611 (N_611,In_1499,In_580);
nor U612 (N_612,In_796,In_973);
and U613 (N_613,In_275,In_867);
or U614 (N_614,In_1166,In_1036);
nand U615 (N_615,In_964,In_477);
nand U616 (N_616,In_678,In_456);
or U617 (N_617,In_966,In_312);
nand U618 (N_618,In_674,In_1395);
or U619 (N_619,In_1048,In_528);
nand U620 (N_620,In_546,In_925);
or U621 (N_621,In_1003,In_423);
and U622 (N_622,In_869,In_631);
xnor U623 (N_623,In_281,In_1060);
nand U624 (N_624,In_517,In_1207);
nand U625 (N_625,In_519,In_244);
or U626 (N_626,In_1295,In_1236);
xnor U627 (N_627,In_561,In_515);
or U628 (N_628,In_1219,In_1097);
nor U629 (N_629,In_944,In_989);
or U630 (N_630,In_417,In_893);
nor U631 (N_631,In_1241,In_646);
or U632 (N_632,In_451,In_258);
nor U633 (N_633,In_328,In_1042);
nand U634 (N_634,In_707,In_1459);
nor U635 (N_635,In_1134,In_891);
nor U636 (N_636,In_1160,In_711);
and U637 (N_637,In_574,In_156);
nor U638 (N_638,In_843,In_684);
nand U639 (N_639,In_1224,In_154);
nand U640 (N_640,In_730,In_215);
and U641 (N_641,In_929,In_238);
or U642 (N_642,In_374,In_901);
nor U643 (N_643,In_1179,In_868);
and U644 (N_644,In_313,In_1333);
and U645 (N_645,In_96,In_329);
and U646 (N_646,In_1078,In_342);
nand U647 (N_647,In_727,In_1135);
nand U648 (N_648,In_865,In_1232);
nor U649 (N_649,In_1095,In_504);
xnor U650 (N_650,In_1426,In_1122);
nor U651 (N_651,In_609,In_1432);
nor U652 (N_652,In_1272,In_433);
and U653 (N_653,In_1439,In_1041);
or U654 (N_654,In_1258,In_1389);
or U655 (N_655,In_129,In_696);
nand U656 (N_656,In_525,In_1021);
nand U657 (N_657,In_1472,In_761);
nor U658 (N_658,In_1252,In_1335);
or U659 (N_659,In_502,In_158);
nor U660 (N_660,In_10,In_838);
nor U661 (N_661,In_331,In_479);
and U662 (N_662,In_117,In_1112);
nand U663 (N_663,In_675,In_980);
and U664 (N_664,In_1366,In_832);
nor U665 (N_665,In_823,In_246);
or U666 (N_666,In_566,In_438);
xnor U667 (N_667,In_138,In_776);
nor U668 (N_668,In_1255,In_679);
nand U669 (N_669,In_187,In_1010);
nand U670 (N_670,In_1244,In_1176);
and U671 (N_671,In_1103,In_1239);
and U672 (N_672,In_393,In_463);
nand U673 (N_673,In_562,In_271);
xnor U674 (N_674,In_309,In_926);
or U675 (N_675,In_115,In_995);
and U676 (N_676,In_285,In_1270);
nor U677 (N_677,In_1391,In_1150);
or U678 (N_678,In_651,In_1317);
xor U679 (N_679,In_656,In_702);
xnor U680 (N_680,In_1273,In_1334);
or U681 (N_681,In_873,In_1198);
or U682 (N_682,In_1284,In_731);
or U683 (N_683,In_922,In_1051);
and U684 (N_684,In_1417,In_688);
and U685 (N_685,In_297,In_121);
nand U686 (N_686,In_1375,In_518);
xor U687 (N_687,In_287,In_123);
and U688 (N_688,In_241,In_1350);
xor U689 (N_689,In_52,In_1381);
xnor U690 (N_690,In_781,In_1173);
or U691 (N_691,In_606,In_178);
or U692 (N_692,In_787,In_896);
and U693 (N_693,In_827,In_1034);
or U694 (N_694,In_974,In_427);
or U695 (N_695,In_170,In_232);
or U696 (N_696,In_523,In_1419);
nor U697 (N_697,In_1189,In_548);
or U698 (N_698,In_975,In_807);
nand U699 (N_699,In_1250,In_1416);
or U700 (N_700,In_211,In_824);
and U701 (N_701,In_1012,In_1143);
nand U702 (N_702,In_861,In_667);
nor U703 (N_703,In_440,In_993);
nand U704 (N_704,In_1453,In_990);
nor U705 (N_705,In_545,In_200);
nor U706 (N_706,In_321,In_208);
and U707 (N_707,In_100,In_1277);
and U708 (N_708,In_623,In_835);
nand U709 (N_709,In_1033,In_212);
or U710 (N_710,In_294,In_80);
and U711 (N_711,In_960,In_1392);
or U712 (N_712,In_405,In_1495);
or U713 (N_713,In_106,In_1433);
nand U714 (N_714,In_1061,In_876);
and U715 (N_715,In_112,In_353);
and U716 (N_716,In_70,In_444);
nor U717 (N_717,In_1063,In_1007);
nand U718 (N_718,In_1227,In_266);
and U719 (N_719,In_575,In_229);
and U720 (N_720,In_825,In_58);
nand U721 (N_721,In_659,In_913);
or U722 (N_722,In_1486,In_968);
nor U723 (N_723,In_73,In_976);
nor U724 (N_724,In_737,In_1445);
and U725 (N_725,In_583,In_98);
nor U726 (N_726,In_1477,In_541);
nand U727 (N_727,In_955,In_622);
nor U728 (N_728,In_790,In_908);
or U729 (N_729,In_914,In_1358);
and U730 (N_730,In_818,In_1131);
or U731 (N_731,In_1215,In_360);
nor U732 (N_732,In_368,In_160);
nor U733 (N_733,In_512,In_265);
or U734 (N_734,In_195,In_1408);
nor U735 (N_735,In_947,In_564);
or U736 (N_736,In_349,In_551);
nor U737 (N_737,In_1022,In_333);
nor U738 (N_738,In_1077,In_146);
xor U739 (N_739,In_505,In_191);
nand U740 (N_740,In_1488,In_1099);
nor U741 (N_741,In_527,In_816);
nand U742 (N_742,In_396,In_507);
nand U743 (N_743,In_863,In_1211);
nor U744 (N_744,In_1328,In_677);
nand U745 (N_745,In_612,In_588);
xnor U746 (N_746,In_997,In_428);
nand U747 (N_747,In_295,In_116);
and U748 (N_748,In_919,In_539);
or U749 (N_749,In_217,In_1249);
or U750 (N_750,In_1435,In_1047);
nor U751 (N_751,In_195,In_1127);
and U752 (N_752,In_449,In_1328);
and U753 (N_753,In_105,In_1374);
nand U754 (N_754,In_109,In_596);
nand U755 (N_755,In_751,In_1499);
and U756 (N_756,In_351,In_7);
and U757 (N_757,In_1085,In_381);
xor U758 (N_758,In_620,In_1063);
nand U759 (N_759,In_1248,In_1161);
and U760 (N_760,In_694,In_1485);
or U761 (N_761,In_1398,In_1304);
nand U762 (N_762,In_777,In_523);
nor U763 (N_763,In_152,In_1395);
nor U764 (N_764,In_1170,In_1380);
nor U765 (N_765,In_744,In_864);
or U766 (N_766,In_207,In_1399);
nor U767 (N_767,In_1280,In_934);
nor U768 (N_768,In_139,In_613);
or U769 (N_769,In_1373,In_1413);
nor U770 (N_770,In_1295,In_8);
and U771 (N_771,In_1322,In_1300);
xor U772 (N_772,In_1098,In_1285);
nor U773 (N_773,In_1431,In_1205);
and U774 (N_774,In_647,In_1491);
and U775 (N_775,In_986,In_1038);
nand U776 (N_776,In_995,In_1443);
or U777 (N_777,In_1498,In_389);
nor U778 (N_778,In_464,In_1261);
nand U779 (N_779,In_89,In_1028);
and U780 (N_780,In_698,In_1414);
nor U781 (N_781,In_816,In_1359);
nor U782 (N_782,In_315,In_576);
or U783 (N_783,In_1081,In_846);
and U784 (N_784,In_1129,In_1148);
and U785 (N_785,In_329,In_460);
and U786 (N_786,In_945,In_566);
nand U787 (N_787,In_785,In_541);
or U788 (N_788,In_1089,In_1495);
or U789 (N_789,In_720,In_992);
and U790 (N_790,In_584,In_202);
nand U791 (N_791,In_1378,In_626);
or U792 (N_792,In_855,In_1248);
xor U793 (N_793,In_246,In_672);
nor U794 (N_794,In_71,In_1378);
nor U795 (N_795,In_1027,In_1333);
and U796 (N_796,In_626,In_1013);
or U797 (N_797,In_140,In_789);
and U798 (N_798,In_1055,In_1168);
and U799 (N_799,In_905,In_190);
nand U800 (N_800,In_166,In_1100);
and U801 (N_801,In_1388,In_661);
nor U802 (N_802,In_610,In_505);
and U803 (N_803,In_236,In_231);
nand U804 (N_804,In_903,In_1226);
and U805 (N_805,In_47,In_751);
nand U806 (N_806,In_1020,In_793);
nand U807 (N_807,In_380,In_750);
or U808 (N_808,In_822,In_229);
nand U809 (N_809,In_914,In_136);
and U810 (N_810,In_239,In_1145);
nor U811 (N_811,In_342,In_78);
and U812 (N_812,In_442,In_261);
nand U813 (N_813,In_869,In_1476);
and U814 (N_814,In_1426,In_1006);
nor U815 (N_815,In_845,In_833);
or U816 (N_816,In_1401,In_542);
or U817 (N_817,In_957,In_195);
or U818 (N_818,In_197,In_429);
nor U819 (N_819,In_1369,In_139);
or U820 (N_820,In_342,In_8);
or U821 (N_821,In_1394,In_15);
or U822 (N_822,In_465,In_801);
or U823 (N_823,In_246,In_1134);
or U824 (N_824,In_913,In_210);
xor U825 (N_825,In_502,In_125);
and U826 (N_826,In_1318,In_962);
nor U827 (N_827,In_52,In_681);
or U828 (N_828,In_736,In_775);
nor U829 (N_829,In_1362,In_270);
xnor U830 (N_830,In_488,In_905);
and U831 (N_831,In_508,In_833);
nor U832 (N_832,In_1019,In_186);
or U833 (N_833,In_882,In_435);
and U834 (N_834,In_867,In_315);
nor U835 (N_835,In_1438,In_749);
and U836 (N_836,In_948,In_432);
nand U837 (N_837,In_188,In_1240);
nand U838 (N_838,In_1437,In_313);
nand U839 (N_839,In_1208,In_327);
nand U840 (N_840,In_154,In_258);
and U841 (N_841,In_219,In_425);
or U842 (N_842,In_1326,In_755);
or U843 (N_843,In_719,In_352);
or U844 (N_844,In_447,In_704);
and U845 (N_845,In_1065,In_1112);
nor U846 (N_846,In_116,In_158);
or U847 (N_847,In_1126,In_700);
nand U848 (N_848,In_945,In_723);
or U849 (N_849,In_1040,In_945);
or U850 (N_850,In_1197,In_783);
nand U851 (N_851,In_379,In_1348);
nor U852 (N_852,In_1446,In_693);
xnor U853 (N_853,In_902,In_345);
or U854 (N_854,In_460,In_415);
and U855 (N_855,In_1396,In_861);
nor U856 (N_856,In_1133,In_804);
and U857 (N_857,In_722,In_839);
nor U858 (N_858,In_679,In_401);
nand U859 (N_859,In_23,In_786);
nand U860 (N_860,In_1110,In_1198);
nor U861 (N_861,In_635,In_46);
xnor U862 (N_862,In_518,In_177);
and U863 (N_863,In_1100,In_349);
or U864 (N_864,In_1306,In_165);
and U865 (N_865,In_1270,In_615);
or U866 (N_866,In_1258,In_661);
or U867 (N_867,In_387,In_191);
nand U868 (N_868,In_1103,In_880);
nand U869 (N_869,In_701,In_865);
and U870 (N_870,In_1153,In_890);
or U871 (N_871,In_881,In_235);
nor U872 (N_872,In_1448,In_455);
nand U873 (N_873,In_836,In_436);
nand U874 (N_874,In_287,In_733);
or U875 (N_875,In_1119,In_710);
and U876 (N_876,In_1491,In_16);
or U877 (N_877,In_1402,In_1441);
xnor U878 (N_878,In_260,In_117);
and U879 (N_879,In_611,In_152);
nor U880 (N_880,In_925,In_1313);
xor U881 (N_881,In_1449,In_771);
nand U882 (N_882,In_550,In_169);
or U883 (N_883,In_143,In_189);
or U884 (N_884,In_1174,In_809);
or U885 (N_885,In_1067,In_305);
nor U886 (N_886,In_771,In_552);
nand U887 (N_887,In_167,In_1017);
or U888 (N_888,In_44,In_885);
or U889 (N_889,In_305,In_1107);
xnor U890 (N_890,In_643,In_648);
or U891 (N_891,In_1233,In_661);
and U892 (N_892,In_460,In_724);
nor U893 (N_893,In_1255,In_153);
or U894 (N_894,In_170,In_213);
nor U895 (N_895,In_156,In_515);
and U896 (N_896,In_409,In_370);
xnor U897 (N_897,In_540,In_58);
or U898 (N_898,In_731,In_155);
and U899 (N_899,In_1012,In_407);
xnor U900 (N_900,In_1038,In_31);
xnor U901 (N_901,In_757,In_860);
xnor U902 (N_902,In_1150,In_1340);
nor U903 (N_903,In_460,In_1497);
nand U904 (N_904,In_396,In_586);
xor U905 (N_905,In_697,In_1324);
and U906 (N_906,In_688,In_1406);
or U907 (N_907,In_57,In_174);
xnor U908 (N_908,In_32,In_77);
and U909 (N_909,In_647,In_537);
or U910 (N_910,In_94,In_1198);
nand U911 (N_911,In_139,In_465);
nor U912 (N_912,In_955,In_329);
and U913 (N_913,In_1019,In_382);
nor U914 (N_914,In_417,In_1413);
nand U915 (N_915,In_1205,In_80);
or U916 (N_916,In_1322,In_696);
and U917 (N_917,In_1037,In_1190);
and U918 (N_918,In_1406,In_174);
nand U919 (N_919,In_382,In_1161);
xor U920 (N_920,In_1117,In_276);
and U921 (N_921,In_327,In_660);
nand U922 (N_922,In_588,In_966);
and U923 (N_923,In_246,In_1063);
nand U924 (N_924,In_1429,In_1007);
and U925 (N_925,In_881,In_840);
and U926 (N_926,In_516,In_1142);
nor U927 (N_927,In_1378,In_476);
and U928 (N_928,In_61,In_80);
nor U929 (N_929,In_1000,In_1103);
nand U930 (N_930,In_1451,In_1154);
and U931 (N_931,In_1061,In_1179);
nand U932 (N_932,In_1213,In_350);
nor U933 (N_933,In_1449,In_326);
or U934 (N_934,In_70,In_75);
xnor U935 (N_935,In_1420,In_846);
nand U936 (N_936,In_173,In_82);
or U937 (N_937,In_813,In_1240);
and U938 (N_938,In_297,In_561);
and U939 (N_939,In_694,In_1060);
and U940 (N_940,In_26,In_1352);
nand U941 (N_941,In_228,In_567);
nor U942 (N_942,In_1009,In_383);
and U943 (N_943,In_524,In_49);
and U944 (N_944,In_469,In_1084);
or U945 (N_945,In_1239,In_1175);
nand U946 (N_946,In_703,In_667);
xor U947 (N_947,In_894,In_677);
and U948 (N_948,In_1468,In_22);
or U949 (N_949,In_876,In_136);
nor U950 (N_950,In_92,In_36);
nor U951 (N_951,In_1431,In_776);
xnor U952 (N_952,In_1090,In_119);
or U953 (N_953,In_1174,In_1167);
and U954 (N_954,In_366,In_911);
or U955 (N_955,In_1249,In_0);
xnor U956 (N_956,In_772,In_1203);
nor U957 (N_957,In_25,In_194);
xor U958 (N_958,In_1406,In_527);
and U959 (N_959,In_887,In_974);
and U960 (N_960,In_489,In_1321);
and U961 (N_961,In_1319,In_783);
nor U962 (N_962,In_301,In_617);
or U963 (N_963,In_868,In_1488);
nor U964 (N_964,In_1455,In_1484);
nor U965 (N_965,In_913,In_1219);
nor U966 (N_966,In_1323,In_75);
nand U967 (N_967,In_519,In_1225);
xor U968 (N_968,In_1336,In_86);
nor U969 (N_969,In_1420,In_803);
nand U970 (N_970,In_876,In_814);
or U971 (N_971,In_527,In_1314);
and U972 (N_972,In_1102,In_839);
or U973 (N_973,In_1261,In_705);
nor U974 (N_974,In_118,In_1174);
nand U975 (N_975,In_541,In_460);
and U976 (N_976,In_1361,In_493);
nand U977 (N_977,In_1003,In_428);
nor U978 (N_978,In_1325,In_134);
or U979 (N_979,In_1189,In_1261);
or U980 (N_980,In_734,In_363);
and U981 (N_981,In_242,In_223);
nor U982 (N_982,In_909,In_832);
or U983 (N_983,In_112,In_315);
nand U984 (N_984,In_1072,In_422);
nand U985 (N_985,In_77,In_1251);
or U986 (N_986,In_1398,In_81);
xor U987 (N_987,In_589,In_1052);
nand U988 (N_988,In_1271,In_461);
nand U989 (N_989,In_387,In_1140);
and U990 (N_990,In_195,In_1226);
and U991 (N_991,In_652,In_1410);
xor U992 (N_992,In_1498,In_1440);
or U993 (N_993,In_1088,In_599);
and U994 (N_994,In_1217,In_527);
nand U995 (N_995,In_1208,In_470);
and U996 (N_996,In_349,In_454);
nand U997 (N_997,In_273,In_1400);
and U998 (N_998,In_1138,In_177);
or U999 (N_999,In_760,In_1093);
and U1000 (N_1000,In_702,In_1402);
nand U1001 (N_1001,In_883,In_170);
xor U1002 (N_1002,In_197,In_219);
nand U1003 (N_1003,In_492,In_322);
and U1004 (N_1004,In_1326,In_842);
or U1005 (N_1005,In_499,In_781);
or U1006 (N_1006,In_1491,In_589);
nor U1007 (N_1007,In_785,In_1004);
or U1008 (N_1008,In_338,In_677);
and U1009 (N_1009,In_981,In_1231);
nand U1010 (N_1010,In_1159,In_641);
and U1011 (N_1011,In_1382,In_1206);
or U1012 (N_1012,In_705,In_681);
nand U1013 (N_1013,In_1149,In_52);
nand U1014 (N_1014,In_216,In_297);
or U1015 (N_1015,In_1441,In_406);
and U1016 (N_1016,In_681,In_216);
nor U1017 (N_1017,In_1260,In_1408);
nor U1018 (N_1018,In_1082,In_256);
and U1019 (N_1019,In_482,In_1187);
or U1020 (N_1020,In_1021,In_623);
xnor U1021 (N_1021,In_929,In_819);
nor U1022 (N_1022,In_933,In_194);
nor U1023 (N_1023,In_139,In_161);
or U1024 (N_1024,In_369,In_842);
nor U1025 (N_1025,In_247,In_1259);
xor U1026 (N_1026,In_238,In_861);
or U1027 (N_1027,In_866,In_653);
nand U1028 (N_1028,In_858,In_622);
nor U1029 (N_1029,In_1059,In_960);
and U1030 (N_1030,In_592,In_969);
nand U1031 (N_1031,In_523,In_603);
and U1032 (N_1032,In_848,In_725);
nor U1033 (N_1033,In_703,In_400);
xnor U1034 (N_1034,In_1385,In_1192);
nor U1035 (N_1035,In_1207,In_959);
xnor U1036 (N_1036,In_878,In_357);
nand U1037 (N_1037,In_265,In_279);
xnor U1038 (N_1038,In_1037,In_1373);
or U1039 (N_1039,In_411,In_582);
or U1040 (N_1040,In_439,In_620);
or U1041 (N_1041,In_274,In_65);
or U1042 (N_1042,In_1274,In_894);
nor U1043 (N_1043,In_1086,In_381);
xnor U1044 (N_1044,In_103,In_1288);
or U1045 (N_1045,In_1047,In_713);
or U1046 (N_1046,In_1460,In_775);
and U1047 (N_1047,In_573,In_1178);
or U1048 (N_1048,In_1358,In_736);
nand U1049 (N_1049,In_85,In_226);
and U1050 (N_1050,In_11,In_1472);
nand U1051 (N_1051,In_1216,In_269);
and U1052 (N_1052,In_1209,In_1216);
nand U1053 (N_1053,In_559,In_448);
nor U1054 (N_1054,In_768,In_577);
nor U1055 (N_1055,In_62,In_1134);
xor U1056 (N_1056,In_790,In_256);
or U1057 (N_1057,In_241,In_1362);
nand U1058 (N_1058,In_231,In_49);
xnor U1059 (N_1059,In_918,In_913);
nand U1060 (N_1060,In_276,In_1321);
and U1061 (N_1061,In_593,In_483);
nand U1062 (N_1062,In_235,In_116);
nor U1063 (N_1063,In_194,In_145);
or U1064 (N_1064,In_323,In_1307);
nor U1065 (N_1065,In_1404,In_883);
or U1066 (N_1066,In_16,In_1240);
and U1067 (N_1067,In_160,In_1034);
xnor U1068 (N_1068,In_794,In_275);
nand U1069 (N_1069,In_562,In_69);
nand U1070 (N_1070,In_52,In_259);
nor U1071 (N_1071,In_347,In_322);
nor U1072 (N_1072,In_198,In_331);
xor U1073 (N_1073,In_94,In_893);
nand U1074 (N_1074,In_718,In_967);
nor U1075 (N_1075,In_1027,In_30);
nand U1076 (N_1076,In_1127,In_1405);
nand U1077 (N_1077,In_95,In_350);
xor U1078 (N_1078,In_52,In_1030);
xor U1079 (N_1079,In_791,In_166);
xnor U1080 (N_1080,In_11,In_577);
or U1081 (N_1081,In_885,In_669);
and U1082 (N_1082,In_8,In_457);
or U1083 (N_1083,In_1192,In_407);
or U1084 (N_1084,In_918,In_787);
and U1085 (N_1085,In_512,In_1411);
and U1086 (N_1086,In_1493,In_493);
or U1087 (N_1087,In_1382,In_631);
nand U1088 (N_1088,In_1219,In_1197);
nor U1089 (N_1089,In_155,In_32);
or U1090 (N_1090,In_594,In_709);
nor U1091 (N_1091,In_500,In_1393);
or U1092 (N_1092,In_1311,In_797);
and U1093 (N_1093,In_1404,In_1422);
or U1094 (N_1094,In_218,In_1009);
nand U1095 (N_1095,In_118,In_1285);
nor U1096 (N_1096,In_397,In_1038);
or U1097 (N_1097,In_1423,In_928);
nor U1098 (N_1098,In_723,In_932);
nand U1099 (N_1099,In_758,In_263);
or U1100 (N_1100,In_955,In_875);
and U1101 (N_1101,In_155,In_978);
nor U1102 (N_1102,In_673,In_312);
and U1103 (N_1103,In_1238,In_909);
and U1104 (N_1104,In_189,In_300);
nand U1105 (N_1105,In_1290,In_1181);
nand U1106 (N_1106,In_1136,In_1223);
nor U1107 (N_1107,In_238,In_634);
and U1108 (N_1108,In_647,In_737);
nor U1109 (N_1109,In_1261,In_360);
nand U1110 (N_1110,In_918,In_223);
and U1111 (N_1111,In_1321,In_1202);
and U1112 (N_1112,In_385,In_1069);
or U1113 (N_1113,In_427,In_843);
or U1114 (N_1114,In_550,In_1425);
nor U1115 (N_1115,In_1190,In_1007);
and U1116 (N_1116,In_302,In_249);
nor U1117 (N_1117,In_1447,In_1105);
nand U1118 (N_1118,In_432,In_1336);
and U1119 (N_1119,In_352,In_1224);
xor U1120 (N_1120,In_16,In_473);
or U1121 (N_1121,In_670,In_433);
and U1122 (N_1122,In_948,In_690);
or U1123 (N_1123,In_766,In_1373);
nor U1124 (N_1124,In_1270,In_1395);
and U1125 (N_1125,In_763,In_653);
xor U1126 (N_1126,In_908,In_329);
nor U1127 (N_1127,In_1331,In_607);
and U1128 (N_1128,In_777,In_131);
nor U1129 (N_1129,In_37,In_1221);
xor U1130 (N_1130,In_1138,In_1239);
or U1131 (N_1131,In_200,In_626);
and U1132 (N_1132,In_1455,In_534);
nand U1133 (N_1133,In_1153,In_896);
and U1134 (N_1134,In_1055,In_1442);
nand U1135 (N_1135,In_74,In_65);
or U1136 (N_1136,In_1453,In_374);
and U1137 (N_1137,In_1000,In_1460);
and U1138 (N_1138,In_302,In_952);
and U1139 (N_1139,In_907,In_1302);
nand U1140 (N_1140,In_1152,In_325);
or U1141 (N_1141,In_1088,In_10);
nor U1142 (N_1142,In_1101,In_692);
nand U1143 (N_1143,In_466,In_825);
or U1144 (N_1144,In_1336,In_1298);
nor U1145 (N_1145,In_328,In_448);
and U1146 (N_1146,In_570,In_473);
nor U1147 (N_1147,In_440,In_879);
xnor U1148 (N_1148,In_831,In_865);
nand U1149 (N_1149,In_1,In_1139);
nand U1150 (N_1150,In_1150,In_217);
and U1151 (N_1151,In_732,In_73);
nand U1152 (N_1152,In_283,In_974);
nor U1153 (N_1153,In_944,In_1040);
and U1154 (N_1154,In_1173,In_597);
and U1155 (N_1155,In_1341,In_1267);
nor U1156 (N_1156,In_285,In_835);
nor U1157 (N_1157,In_1418,In_470);
nor U1158 (N_1158,In_120,In_696);
nand U1159 (N_1159,In_653,In_229);
nand U1160 (N_1160,In_821,In_135);
or U1161 (N_1161,In_1192,In_1159);
nand U1162 (N_1162,In_353,In_578);
xnor U1163 (N_1163,In_319,In_448);
and U1164 (N_1164,In_539,In_530);
or U1165 (N_1165,In_478,In_926);
or U1166 (N_1166,In_530,In_500);
or U1167 (N_1167,In_1170,In_1327);
nand U1168 (N_1168,In_1017,In_593);
nor U1169 (N_1169,In_62,In_189);
or U1170 (N_1170,In_1462,In_736);
xor U1171 (N_1171,In_768,In_197);
nor U1172 (N_1172,In_1298,In_1332);
or U1173 (N_1173,In_387,In_1447);
xor U1174 (N_1174,In_146,In_640);
nor U1175 (N_1175,In_1179,In_1030);
nor U1176 (N_1176,In_474,In_1050);
nand U1177 (N_1177,In_1307,In_1283);
nand U1178 (N_1178,In_1244,In_866);
nand U1179 (N_1179,In_1204,In_1256);
nor U1180 (N_1180,In_607,In_859);
and U1181 (N_1181,In_812,In_1454);
nor U1182 (N_1182,In_1091,In_1154);
nor U1183 (N_1183,In_315,In_733);
nor U1184 (N_1184,In_1104,In_1349);
nand U1185 (N_1185,In_796,In_1252);
and U1186 (N_1186,In_533,In_636);
and U1187 (N_1187,In_1466,In_731);
or U1188 (N_1188,In_273,In_2);
or U1189 (N_1189,In_1024,In_628);
nand U1190 (N_1190,In_453,In_540);
xor U1191 (N_1191,In_1127,In_363);
nor U1192 (N_1192,In_6,In_659);
nor U1193 (N_1193,In_1428,In_375);
nor U1194 (N_1194,In_250,In_1159);
and U1195 (N_1195,In_1444,In_724);
and U1196 (N_1196,In_789,In_1087);
nand U1197 (N_1197,In_520,In_765);
or U1198 (N_1198,In_1362,In_1223);
or U1199 (N_1199,In_1194,In_1016);
nor U1200 (N_1200,In_890,In_568);
and U1201 (N_1201,In_815,In_539);
or U1202 (N_1202,In_1262,In_564);
and U1203 (N_1203,In_424,In_818);
and U1204 (N_1204,In_1284,In_580);
and U1205 (N_1205,In_971,In_1255);
nand U1206 (N_1206,In_1295,In_649);
or U1207 (N_1207,In_1113,In_1028);
xor U1208 (N_1208,In_979,In_1175);
or U1209 (N_1209,In_837,In_496);
or U1210 (N_1210,In_252,In_976);
and U1211 (N_1211,In_19,In_1371);
and U1212 (N_1212,In_996,In_687);
xnor U1213 (N_1213,In_1072,In_1489);
nand U1214 (N_1214,In_745,In_546);
xnor U1215 (N_1215,In_133,In_149);
and U1216 (N_1216,In_360,In_293);
nor U1217 (N_1217,In_350,In_852);
nor U1218 (N_1218,In_825,In_1388);
xor U1219 (N_1219,In_1418,In_527);
nor U1220 (N_1220,In_1246,In_395);
and U1221 (N_1221,In_509,In_595);
or U1222 (N_1222,In_1160,In_376);
or U1223 (N_1223,In_1206,In_712);
nand U1224 (N_1224,In_460,In_120);
nor U1225 (N_1225,In_1193,In_1363);
nand U1226 (N_1226,In_612,In_1172);
nor U1227 (N_1227,In_500,In_408);
and U1228 (N_1228,In_471,In_1232);
xnor U1229 (N_1229,In_1041,In_240);
nor U1230 (N_1230,In_1117,In_1295);
or U1231 (N_1231,In_978,In_1177);
and U1232 (N_1232,In_1305,In_317);
and U1233 (N_1233,In_537,In_1096);
nor U1234 (N_1234,In_1116,In_1496);
or U1235 (N_1235,In_136,In_595);
and U1236 (N_1236,In_69,In_72);
or U1237 (N_1237,In_221,In_68);
or U1238 (N_1238,In_1329,In_408);
nor U1239 (N_1239,In_166,In_1294);
nand U1240 (N_1240,In_664,In_891);
nor U1241 (N_1241,In_1183,In_445);
or U1242 (N_1242,In_1446,In_268);
nor U1243 (N_1243,In_493,In_1396);
and U1244 (N_1244,In_91,In_1467);
nor U1245 (N_1245,In_1106,In_670);
nor U1246 (N_1246,In_361,In_1195);
xor U1247 (N_1247,In_783,In_606);
nand U1248 (N_1248,In_1435,In_1398);
nor U1249 (N_1249,In_1306,In_57);
nand U1250 (N_1250,In_1228,In_1127);
nand U1251 (N_1251,In_22,In_98);
and U1252 (N_1252,In_271,In_45);
and U1253 (N_1253,In_342,In_1190);
and U1254 (N_1254,In_841,In_918);
or U1255 (N_1255,In_200,In_919);
or U1256 (N_1256,In_909,In_79);
and U1257 (N_1257,In_219,In_302);
nand U1258 (N_1258,In_511,In_359);
nor U1259 (N_1259,In_468,In_111);
or U1260 (N_1260,In_231,In_851);
and U1261 (N_1261,In_679,In_524);
nor U1262 (N_1262,In_583,In_586);
xor U1263 (N_1263,In_1100,In_1389);
xor U1264 (N_1264,In_46,In_1354);
and U1265 (N_1265,In_152,In_546);
nand U1266 (N_1266,In_878,In_506);
and U1267 (N_1267,In_1102,In_1349);
xnor U1268 (N_1268,In_599,In_166);
nand U1269 (N_1269,In_1226,In_61);
and U1270 (N_1270,In_1156,In_505);
nor U1271 (N_1271,In_1016,In_174);
or U1272 (N_1272,In_366,In_92);
or U1273 (N_1273,In_508,In_1307);
nor U1274 (N_1274,In_493,In_1286);
nand U1275 (N_1275,In_1067,In_1050);
or U1276 (N_1276,In_1319,In_1257);
nand U1277 (N_1277,In_1085,In_1229);
nand U1278 (N_1278,In_343,In_822);
nand U1279 (N_1279,In_421,In_4);
nand U1280 (N_1280,In_1343,In_755);
nor U1281 (N_1281,In_553,In_188);
or U1282 (N_1282,In_904,In_689);
and U1283 (N_1283,In_642,In_1031);
or U1284 (N_1284,In_435,In_1090);
and U1285 (N_1285,In_788,In_1404);
or U1286 (N_1286,In_1377,In_760);
nand U1287 (N_1287,In_784,In_369);
or U1288 (N_1288,In_1071,In_588);
nand U1289 (N_1289,In_823,In_221);
nand U1290 (N_1290,In_342,In_1034);
nor U1291 (N_1291,In_1412,In_327);
and U1292 (N_1292,In_831,In_1337);
and U1293 (N_1293,In_852,In_210);
nand U1294 (N_1294,In_463,In_258);
and U1295 (N_1295,In_1391,In_1483);
and U1296 (N_1296,In_1354,In_1423);
nor U1297 (N_1297,In_349,In_1489);
xnor U1298 (N_1298,In_494,In_960);
nand U1299 (N_1299,In_422,In_897);
nor U1300 (N_1300,In_182,In_661);
or U1301 (N_1301,In_1288,In_1310);
nor U1302 (N_1302,In_1059,In_844);
or U1303 (N_1303,In_990,In_1180);
nand U1304 (N_1304,In_22,In_638);
and U1305 (N_1305,In_501,In_616);
or U1306 (N_1306,In_551,In_281);
and U1307 (N_1307,In_1029,In_698);
nor U1308 (N_1308,In_774,In_209);
and U1309 (N_1309,In_218,In_780);
or U1310 (N_1310,In_1155,In_1341);
nand U1311 (N_1311,In_777,In_763);
xnor U1312 (N_1312,In_254,In_1299);
or U1313 (N_1313,In_762,In_1497);
nand U1314 (N_1314,In_407,In_876);
nor U1315 (N_1315,In_443,In_559);
or U1316 (N_1316,In_161,In_815);
nand U1317 (N_1317,In_1222,In_1131);
or U1318 (N_1318,In_944,In_529);
nand U1319 (N_1319,In_1225,In_638);
or U1320 (N_1320,In_1077,In_753);
and U1321 (N_1321,In_1435,In_626);
or U1322 (N_1322,In_1009,In_1114);
xor U1323 (N_1323,In_1001,In_322);
and U1324 (N_1324,In_152,In_361);
or U1325 (N_1325,In_422,In_231);
or U1326 (N_1326,In_97,In_61);
and U1327 (N_1327,In_339,In_1268);
and U1328 (N_1328,In_66,In_1266);
and U1329 (N_1329,In_1120,In_1152);
nor U1330 (N_1330,In_1418,In_834);
nor U1331 (N_1331,In_972,In_635);
xnor U1332 (N_1332,In_1480,In_905);
nor U1333 (N_1333,In_1024,In_1245);
xor U1334 (N_1334,In_840,In_1451);
and U1335 (N_1335,In_640,In_722);
or U1336 (N_1336,In_33,In_26);
or U1337 (N_1337,In_192,In_777);
or U1338 (N_1338,In_766,In_1244);
or U1339 (N_1339,In_1468,In_1219);
nand U1340 (N_1340,In_111,In_816);
nor U1341 (N_1341,In_1480,In_234);
or U1342 (N_1342,In_786,In_1411);
or U1343 (N_1343,In_1093,In_1269);
and U1344 (N_1344,In_571,In_1261);
or U1345 (N_1345,In_394,In_739);
nand U1346 (N_1346,In_548,In_561);
xnor U1347 (N_1347,In_139,In_676);
or U1348 (N_1348,In_1220,In_593);
and U1349 (N_1349,In_1343,In_1210);
nor U1350 (N_1350,In_174,In_699);
nor U1351 (N_1351,In_124,In_1010);
xnor U1352 (N_1352,In_292,In_151);
nor U1353 (N_1353,In_922,In_642);
and U1354 (N_1354,In_887,In_98);
nor U1355 (N_1355,In_583,In_1152);
nand U1356 (N_1356,In_1165,In_646);
nor U1357 (N_1357,In_708,In_1294);
nand U1358 (N_1358,In_54,In_934);
nor U1359 (N_1359,In_11,In_625);
or U1360 (N_1360,In_1383,In_185);
xnor U1361 (N_1361,In_890,In_515);
nand U1362 (N_1362,In_329,In_26);
and U1363 (N_1363,In_779,In_32);
nand U1364 (N_1364,In_545,In_980);
nor U1365 (N_1365,In_870,In_1021);
and U1366 (N_1366,In_381,In_1349);
and U1367 (N_1367,In_75,In_1326);
and U1368 (N_1368,In_1349,In_295);
nor U1369 (N_1369,In_1340,In_736);
xnor U1370 (N_1370,In_799,In_409);
nor U1371 (N_1371,In_936,In_1047);
and U1372 (N_1372,In_637,In_104);
nor U1373 (N_1373,In_903,In_533);
and U1374 (N_1374,In_1062,In_455);
or U1375 (N_1375,In_933,In_77);
nand U1376 (N_1376,In_480,In_702);
nand U1377 (N_1377,In_125,In_482);
nand U1378 (N_1378,In_319,In_159);
nand U1379 (N_1379,In_782,In_809);
and U1380 (N_1380,In_621,In_1179);
nor U1381 (N_1381,In_1442,In_1282);
or U1382 (N_1382,In_353,In_1464);
or U1383 (N_1383,In_777,In_1460);
or U1384 (N_1384,In_1200,In_855);
or U1385 (N_1385,In_373,In_1447);
and U1386 (N_1386,In_1185,In_5);
nand U1387 (N_1387,In_85,In_1358);
and U1388 (N_1388,In_875,In_1405);
nand U1389 (N_1389,In_79,In_1125);
nor U1390 (N_1390,In_670,In_1433);
nor U1391 (N_1391,In_1323,In_981);
and U1392 (N_1392,In_524,In_420);
xor U1393 (N_1393,In_379,In_908);
nand U1394 (N_1394,In_1137,In_982);
or U1395 (N_1395,In_1498,In_255);
or U1396 (N_1396,In_1030,In_1390);
nand U1397 (N_1397,In_533,In_536);
or U1398 (N_1398,In_808,In_786);
and U1399 (N_1399,In_886,In_603);
or U1400 (N_1400,In_725,In_1497);
nor U1401 (N_1401,In_441,In_481);
xnor U1402 (N_1402,In_744,In_154);
and U1403 (N_1403,In_1415,In_970);
xnor U1404 (N_1404,In_1163,In_662);
nand U1405 (N_1405,In_1382,In_534);
nand U1406 (N_1406,In_770,In_437);
and U1407 (N_1407,In_1494,In_550);
and U1408 (N_1408,In_288,In_318);
xor U1409 (N_1409,In_1210,In_1258);
xor U1410 (N_1410,In_1477,In_1423);
nor U1411 (N_1411,In_1093,In_1142);
nand U1412 (N_1412,In_133,In_1247);
and U1413 (N_1413,In_581,In_1410);
nand U1414 (N_1414,In_542,In_777);
nand U1415 (N_1415,In_152,In_1203);
xor U1416 (N_1416,In_91,In_756);
and U1417 (N_1417,In_1140,In_464);
nand U1418 (N_1418,In_570,In_1422);
and U1419 (N_1419,In_556,In_394);
and U1420 (N_1420,In_438,In_248);
xor U1421 (N_1421,In_261,In_290);
nand U1422 (N_1422,In_527,In_1395);
nand U1423 (N_1423,In_1448,In_1394);
nor U1424 (N_1424,In_276,In_1174);
or U1425 (N_1425,In_1499,In_1295);
or U1426 (N_1426,In_894,In_200);
nor U1427 (N_1427,In_1326,In_1160);
nor U1428 (N_1428,In_988,In_1192);
and U1429 (N_1429,In_505,In_305);
nand U1430 (N_1430,In_896,In_731);
or U1431 (N_1431,In_67,In_623);
nor U1432 (N_1432,In_174,In_1215);
nand U1433 (N_1433,In_359,In_1359);
nor U1434 (N_1434,In_424,In_561);
and U1435 (N_1435,In_1028,In_45);
or U1436 (N_1436,In_306,In_681);
nor U1437 (N_1437,In_868,In_906);
or U1438 (N_1438,In_1209,In_402);
and U1439 (N_1439,In_212,In_648);
nand U1440 (N_1440,In_1447,In_1055);
nor U1441 (N_1441,In_497,In_1486);
nor U1442 (N_1442,In_852,In_1133);
or U1443 (N_1443,In_1079,In_656);
or U1444 (N_1444,In_1345,In_1444);
nand U1445 (N_1445,In_1430,In_1272);
nor U1446 (N_1446,In_1134,In_392);
and U1447 (N_1447,In_758,In_1388);
nor U1448 (N_1448,In_679,In_191);
nand U1449 (N_1449,In_325,In_936);
and U1450 (N_1450,In_937,In_865);
and U1451 (N_1451,In_1039,In_1110);
or U1452 (N_1452,In_1338,In_770);
or U1453 (N_1453,In_659,In_827);
nor U1454 (N_1454,In_295,In_162);
nor U1455 (N_1455,In_938,In_431);
nor U1456 (N_1456,In_1176,In_354);
nor U1457 (N_1457,In_417,In_21);
nor U1458 (N_1458,In_198,In_428);
or U1459 (N_1459,In_1199,In_207);
nor U1460 (N_1460,In_1359,In_693);
nor U1461 (N_1461,In_479,In_507);
nor U1462 (N_1462,In_715,In_537);
and U1463 (N_1463,In_1347,In_1232);
or U1464 (N_1464,In_762,In_438);
and U1465 (N_1465,In_1178,In_556);
or U1466 (N_1466,In_206,In_143);
or U1467 (N_1467,In_189,In_768);
xnor U1468 (N_1468,In_1162,In_1111);
nand U1469 (N_1469,In_536,In_1114);
nor U1470 (N_1470,In_612,In_276);
nor U1471 (N_1471,In_12,In_1262);
xnor U1472 (N_1472,In_1489,In_1140);
xor U1473 (N_1473,In_676,In_214);
nor U1474 (N_1474,In_1080,In_1092);
or U1475 (N_1475,In_1060,In_911);
nor U1476 (N_1476,In_47,In_673);
xnor U1477 (N_1477,In_1239,In_59);
or U1478 (N_1478,In_473,In_1158);
xor U1479 (N_1479,In_917,In_229);
xnor U1480 (N_1480,In_1480,In_684);
or U1481 (N_1481,In_1461,In_411);
nor U1482 (N_1482,In_317,In_487);
or U1483 (N_1483,In_734,In_426);
and U1484 (N_1484,In_1313,In_501);
nand U1485 (N_1485,In_944,In_1424);
nor U1486 (N_1486,In_798,In_244);
or U1487 (N_1487,In_1215,In_9);
and U1488 (N_1488,In_1127,In_818);
and U1489 (N_1489,In_727,In_944);
nor U1490 (N_1490,In_462,In_983);
nand U1491 (N_1491,In_1403,In_739);
and U1492 (N_1492,In_1246,In_1452);
nand U1493 (N_1493,In_770,In_665);
nor U1494 (N_1494,In_1078,In_953);
nand U1495 (N_1495,In_1149,In_405);
nor U1496 (N_1496,In_333,In_208);
nand U1497 (N_1497,In_553,In_791);
nand U1498 (N_1498,In_405,In_421);
or U1499 (N_1499,In_922,In_818);
nor U1500 (N_1500,In_1279,In_949);
nand U1501 (N_1501,In_1167,In_473);
nand U1502 (N_1502,In_234,In_1081);
nor U1503 (N_1503,In_697,In_823);
and U1504 (N_1504,In_526,In_475);
nand U1505 (N_1505,In_632,In_310);
and U1506 (N_1506,In_991,In_238);
nor U1507 (N_1507,In_732,In_108);
or U1508 (N_1508,In_286,In_1227);
nand U1509 (N_1509,In_473,In_501);
or U1510 (N_1510,In_49,In_375);
nand U1511 (N_1511,In_192,In_259);
and U1512 (N_1512,In_232,In_1226);
and U1513 (N_1513,In_1275,In_394);
and U1514 (N_1514,In_1391,In_485);
nor U1515 (N_1515,In_126,In_1364);
and U1516 (N_1516,In_901,In_992);
or U1517 (N_1517,In_858,In_531);
nand U1518 (N_1518,In_516,In_592);
and U1519 (N_1519,In_308,In_1186);
or U1520 (N_1520,In_47,In_96);
nor U1521 (N_1521,In_1019,In_766);
and U1522 (N_1522,In_958,In_812);
xor U1523 (N_1523,In_388,In_611);
nand U1524 (N_1524,In_409,In_1452);
and U1525 (N_1525,In_448,In_69);
nor U1526 (N_1526,In_529,In_501);
or U1527 (N_1527,In_761,In_566);
nand U1528 (N_1528,In_511,In_471);
and U1529 (N_1529,In_551,In_393);
nand U1530 (N_1530,In_412,In_1222);
and U1531 (N_1531,In_1134,In_1498);
nand U1532 (N_1532,In_908,In_274);
or U1533 (N_1533,In_1411,In_990);
nand U1534 (N_1534,In_816,In_1387);
nand U1535 (N_1535,In_1477,In_1453);
and U1536 (N_1536,In_1438,In_799);
nand U1537 (N_1537,In_336,In_1448);
nor U1538 (N_1538,In_562,In_936);
or U1539 (N_1539,In_848,In_886);
and U1540 (N_1540,In_51,In_247);
nand U1541 (N_1541,In_1106,In_570);
nor U1542 (N_1542,In_1006,In_1014);
xnor U1543 (N_1543,In_295,In_240);
nor U1544 (N_1544,In_1498,In_427);
nor U1545 (N_1545,In_1447,In_330);
nor U1546 (N_1546,In_1177,In_1047);
or U1547 (N_1547,In_1324,In_554);
nand U1548 (N_1548,In_484,In_658);
nor U1549 (N_1549,In_161,In_862);
nor U1550 (N_1550,In_1319,In_987);
nand U1551 (N_1551,In_820,In_246);
and U1552 (N_1552,In_218,In_1352);
or U1553 (N_1553,In_1063,In_1388);
nand U1554 (N_1554,In_1204,In_199);
or U1555 (N_1555,In_288,In_1340);
and U1556 (N_1556,In_64,In_349);
or U1557 (N_1557,In_1475,In_1306);
or U1558 (N_1558,In_1015,In_696);
and U1559 (N_1559,In_791,In_1144);
nor U1560 (N_1560,In_499,In_1132);
and U1561 (N_1561,In_738,In_504);
and U1562 (N_1562,In_308,In_1473);
nand U1563 (N_1563,In_126,In_145);
nand U1564 (N_1564,In_875,In_1192);
nor U1565 (N_1565,In_155,In_980);
and U1566 (N_1566,In_1271,In_24);
and U1567 (N_1567,In_395,In_352);
nor U1568 (N_1568,In_326,In_115);
nor U1569 (N_1569,In_325,In_809);
or U1570 (N_1570,In_406,In_1026);
nand U1571 (N_1571,In_746,In_314);
nor U1572 (N_1572,In_225,In_1419);
nor U1573 (N_1573,In_328,In_213);
or U1574 (N_1574,In_128,In_618);
nand U1575 (N_1575,In_40,In_1346);
or U1576 (N_1576,In_752,In_1319);
xnor U1577 (N_1577,In_1068,In_945);
nor U1578 (N_1578,In_1199,In_266);
nand U1579 (N_1579,In_612,In_736);
and U1580 (N_1580,In_1155,In_1325);
nand U1581 (N_1581,In_1267,In_703);
nor U1582 (N_1582,In_527,In_616);
and U1583 (N_1583,In_1435,In_1498);
or U1584 (N_1584,In_171,In_1005);
nor U1585 (N_1585,In_875,In_79);
and U1586 (N_1586,In_552,In_1307);
nor U1587 (N_1587,In_329,In_1170);
xnor U1588 (N_1588,In_775,In_247);
or U1589 (N_1589,In_269,In_1080);
nand U1590 (N_1590,In_1272,In_806);
nand U1591 (N_1591,In_662,In_631);
or U1592 (N_1592,In_15,In_838);
nor U1593 (N_1593,In_1458,In_648);
or U1594 (N_1594,In_466,In_1217);
or U1595 (N_1595,In_1331,In_219);
nand U1596 (N_1596,In_1,In_1336);
or U1597 (N_1597,In_370,In_266);
nor U1598 (N_1598,In_1389,In_1337);
nor U1599 (N_1599,In_1005,In_308);
or U1600 (N_1600,In_1317,In_1119);
or U1601 (N_1601,In_781,In_776);
nor U1602 (N_1602,In_1339,In_1150);
nor U1603 (N_1603,In_352,In_855);
or U1604 (N_1604,In_1251,In_199);
and U1605 (N_1605,In_665,In_827);
nor U1606 (N_1606,In_898,In_56);
nor U1607 (N_1607,In_18,In_1297);
and U1608 (N_1608,In_208,In_1035);
and U1609 (N_1609,In_224,In_393);
nand U1610 (N_1610,In_545,In_233);
nor U1611 (N_1611,In_30,In_1099);
or U1612 (N_1612,In_329,In_1275);
and U1613 (N_1613,In_1462,In_739);
or U1614 (N_1614,In_242,In_107);
and U1615 (N_1615,In_793,In_1463);
nand U1616 (N_1616,In_1442,In_179);
nand U1617 (N_1617,In_649,In_83);
nand U1618 (N_1618,In_239,In_321);
and U1619 (N_1619,In_1029,In_1025);
nand U1620 (N_1620,In_908,In_1228);
or U1621 (N_1621,In_480,In_1001);
nand U1622 (N_1622,In_810,In_1094);
and U1623 (N_1623,In_1418,In_1085);
or U1624 (N_1624,In_493,In_1325);
and U1625 (N_1625,In_13,In_585);
nand U1626 (N_1626,In_504,In_1324);
nand U1627 (N_1627,In_1337,In_1260);
nor U1628 (N_1628,In_837,In_838);
nand U1629 (N_1629,In_359,In_1362);
or U1630 (N_1630,In_1163,In_1475);
and U1631 (N_1631,In_19,In_937);
nor U1632 (N_1632,In_1218,In_392);
xor U1633 (N_1633,In_927,In_748);
nand U1634 (N_1634,In_633,In_458);
nor U1635 (N_1635,In_382,In_632);
nand U1636 (N_1636,In_702,In_1243);
nor U1637 (N_1637,In_736,In_157);
or U1638 (N_1638,In_1479,In_792);
or U1639 (N_1639,In_1244,In_141);
nand U1640 (N_1640,In_318,In_403);
nand U1641 (N_1641,In_290,In_1439);
nand U1642 (N_1642,In_8,In_101);
and U1643 (N_1643,In_826,In_280);
nor U1644 (N_1644,In_228,In_816);
and U1645 (N_1645,In_1436,In_323);
and U1646 (N_1646,In_41,In_172);
xnor U1647 (N_1647,In_152,In_452);
nor U1648 (N_1648,In_1089,In_226);
xnor U1649 (N_1649,In_610,In_1059);
or U1650 (N_1650,In_1092,In_1224);
or U1651 (N_1651,In_177,In_960);
nor U1652 (N_1652,In_1416,In_1266);
or U1653 (N_1653,In_1475,In_827);
or U1654 (N_1654,In_1346,In_1159);
nand U1655 (N_1655,In_1218,In_650);
nand U1656 (N_1656,In_899,In_1185);
or U1657 (N_1657,In_492,In_70);
nor U1658 (N_1658,In_1099,In_260);
nand U1659 (N_1659,In_1262,In_1098);
or U1660 (N_1660,In_752,In_918);
and U1661 (N_1661,In_414,In_685);
nand U1662 (N_1662,In_1424,In_560);
or U1663 (N_1663,In_534,In_117);
nand U1664 (N_1664,In_267,In_1225);
nand U1665 (N_1665,In_1130,In_1117);
or U1666 (N_1666,In_197,In_1074);
nor U1667 (N_1667,In_863,In_1122);
xor U1668 (N_1668,In_492,In_102);
and U1669 (N_1669,In_70,In_250);
nand U1670 (N_1670,In_1156,In_312);
or U1671 (N_1671,In_1497,In_355);
and U1672 (N_1672,In_521,In_1146);
nand U1673 (N_1673,In_12,In_609);
and U1674 (N_1674,In_1197,In_1200);
nand U1675 (N_1675,In_482,In_60);
nand U1676 (N_1676,In_1115,In_1032);
and U1677 (N_1677,In_116,In_325);
nor U1678 (N_1678,In_1454,In_524);
nor U1679 (N_1679,In_895,In_674);
or U1680 (N_1680,In_769,In_1022);
or U1681 (N_1681,In_626,In_357);
or U1682 (N_1682,In_257,In_405);
and U1683 (N_1683,In_1423,In_802);
nand U1684 (N_1684,In_95,In_22);
nor U1685 (N_1685,In_185,In_862);
and U1686 (N_1686,In_1204,In_1361);
xnor U1687 (N_1687,In_598,In_873);
or U1688 (N_1688,In_1141,In_1225);
or U1689 (N_1689,In_797,In_382);
and U1690 (N_1690,In_264,In_630);
or U1691 (N_1691,In_1170,In_128);
nor U1692 (N_1692,In_179,In_713);
nand U1693 (N_1693,In_883,In_777);
or U1694 (N_1694,In_1227,In_1052);
nor U1695 (N_1695,In_667,In_280);
nand U1696 (N_1696,In_329,In_1435);
nand U1697 (N_1697,In_1457,In_1093);
xor U1698 (N_1698,In_1096,In_775);
and U1699 (N_1699,In_861,In_845);
or U1700 (N_1700,In_1334,In_145);
nand U1701 (N_1701,In_979,In_537);
xor U1702 (N_1702,In_1067,In_864);
nor U1703 (N_1703,In_1117,In_474);
or U1704 (N_1704,In_1000,In_815);
and U1705 (N_1705,In_1487,In_1461);
or U1706 (N_1706,In_1051,In_930);
and U1707 (N_1707,In_406,In_431);
xnor U1708 (N_1708,In_610,In_750);
nor U1709 (N_1709,In_661,In_63);
nand U1710 (N_1710,In_688,In_274);
xnor U1711 (N_1711,In_1069,In_1013);
and U1712 (N_1712,In_347,In_40);
nand U1713 (N_1713,In_931,In_317);
nor U1714 (N_1714,In_1029,In_933);
nor U1715 (N_1715,In_398,In_604);
or U1716 (N_1716,In_1282,In_1437);
xnor U1717 (N_1717,In_718,In_221);
nand U1718 (N_1718,In_1044,In_1351);
nand U1719 (N_1719,In_590,In_1305);
and U1720 (N_1720,In_1107,In_288);
and U1721 (N_1721,In_40,In_773);
and U1722 (N_1722,In_940,In_1191);
or U1723 (N_1723,In_414,In_566);
nor U1724 (N_1724,In_1081,In_1487);
or U1725 (N_1725,In_999,In_664);
and U1726 (N_1726,In_252,In_602);
nor U1727 (N_1727,In_436,In_606);
nand U1728 (N_1728,In_907,In_739);
or U1729 (N_1729,In_570,In_352);
nor U1730 (N_1730,In_412,In_236);
and U1731 (N_1731,In_1392,In_1152);
and U1732 (N_1732,In_507,In_211);
and U1733 (N_1733,In_571,In_1273);
nor U1734 (N_1734,In_737,In_576);
nor U1735 (N_1735,In_1481,In_678);
or U1736 (N_1736,In_1087,In_1067);
and U1737 (N_1737,In_1068,In_1328);
or U1738 (N_1738,In_1011,In_373);
and U1739 (N_1739,In_889,In_1251);
nand U1740 (N_1740,In_293,In_71);
and U1741 (N_1741,In_1027,In_1096);
and U1742 (N_1742,In_1319,In_19);
or U1743 (N_1743,In_419,In_1127);
nor U1744 (N_1744,In_31,In_1167);
and U1745 (N_1745,In_1357,In_1430);
nor U1746 (N_1746,In_436,In_1051);
or U1747 (N_1747,In_1229,In_308);
nand U1748 (N_1748,In_1083,In_670);
nand U1749 (N_1749,In_896,In_900);
xnor U1750 (N_1750,In_893,In_1165);
and U1751 (N_1751,In_1373,In_615);
and U1752 (N_1752,In_506,In_136);
and U1753 (N_1753,In_1378,In_830);
nor U1754 (N_1754,In_205,In_902);
nor U1755 (N_1755,In_4,In_997);
and U1756 (N_1756,In_421,In_246);
nor U1757 (N_1757,In_1095,In_507);
or U1758 (N_1758,In_10,In_445);
and U1759 (N_1759,In_944,In_744);
or U1760 (N_1760,In_1138,In_1490);
nor U1761 (N_1761,In_302,In_373);
or U1762 (N_1762,In_869,In_1444);
or U1763 (N_1763,In_687,In_149);
or U1764 (N_1764,In_1269,In_924);
nand U1765 (N_1765,In_662,In_200);
nand U1766 (N_1766,In_31,In_880);
or U1767 (N_1767,In_1118,In_521);
nor U1768 (N_1768,In_587,In_92);
xnor U1769 (N_1769,In_1359,In_1250);
and U1770 (N_1770,In_423,In_1128);
or U1771 (N_1771,In_219,In_533);
nand U1772 (N_1772,In_1431,In_525);
or U1773 (N_1773,In_1095,In_475);
or U1774 (N_1774,In_56,In_82);
nand U1775 (N_1775,In_1007,In_662);
nor U1776 (N_1776,In_1369,In_892);
or U1777 (N_1777,In_1442,In_321);
nor U1778 (N_1778,In_13,In_1379);
or U1779 (N_1779,In_25,In_1016);
nand U1780 (N_1780,In_1006,In_254);
and U1781 (N_1781,In_61,In_318);
nand U1782 (N_1782,In_628,In_366);
or U1783 (N_1783,In_945,In_970);
and U1784 (N_1784,In_1067,In_28);
and U1785 (N_1785,In_683,In_843);
and U1786 (N_1786,In_1282,In_498);
or U1787 (N_1787,In_1068,In_1314);
nand U1788 (N_1788,In_1460,In_396);
xnor U1789 (N_1789,In_507,In_589);
and U1790 (N_1790,In_311,In_142);
nor U1791 (N_1791,In_291,In_315);
nor U1792 (N_1792,In_1365,In_1304);
nand U1793 (N_1793,In_373,In_195);
nand U1794 (N_1794,In_1486,In_1119);
and U1795 (N_1795,In_555,In_1494);
and U1796 (N_1796,In_10,In_437);
and U1797 (N_1797,In_1182,In_674);
nor U1798 (N_1798,In_850,In_241);
xor U1799 (N_1799,In_1025,In_1412);
or U1800 (N_1800,In_462,In_312);
and U1801 (N_1801,In_719,In_1190);
and U1802 (N_1802,In_679,In_1297);
nand U1803 (N_1803,In_748,In_353);
nor U1804 (N_1804,In_899,In_120);
or U1805 (N_1805,In_837,In_1050);
and U1806 (N_1806,In_1351,In_499);
nand U1807 (N_1807,In_610,In_240);
nor U1808 (N_1808,In_88,In_1237);
nor U1809 (N_1809,In_1291,In_748);
or U1810 (N_1810,In_762,In_1407);
or U1811 (N_1811,In_1386,In_176);
and U1812 (N_1812,In_1087,In_1430);
and U1813 (N_1813,In_1236,In_693);
or U1814 (N_1814,In_1079,In_438);
xnor U1815 (N_1815,In_1362,In_654);
and U1816 (N_1816,In_634,In_657);
and U1817 (N_1817,In_379,In_1082);
and U1818 (N_1818,In_125,In_427);
nor U1819 (N_1819,In_15,In_705);
and U1820 (N_1820,In_983,In_107);
nand U1821 (N_1821,In_76,In_173);
and U1822 (N_1822,In_1303,In_394);
nor U1823 (N_1823,In_797,In_975);
nand U1824 (N_1824,In_650,In_1092);
xor U1825 (N_1825,In_554,In_883);
and U1826 (N_1826,In_633,In_121);
and U1827 (N_1827,In_648,In_458);
nor U1828 (N_1828,In_1301,In_1214);
nor U1829 (N_1829,In_368,In_541);
nor U1830 (N_1830,In_57,In_293);
nor U1831 (N_1831,In_940,In_264);
nand U1832 (N_1832,In_1399,In_334);
or U1833 (N_1833,In_986,In_1119);
and U1834 (N_1834,In_977,In_974);
or U1835 (N_1835,In_1121,In_200);
and U1836 (N_1836,In_599,In_1232);
nor U1837 (N_1837,In_1473,In_536);
nand U1838 (N_1838,In_152,In_1306);
nor U1839 (N_1839,In_774,In_315);
nand U1840 (N_1840,In_1230,In_25);
or U1841 (N_1841,In_1402,In_1128);
nor U1842 (N_1842,In_588,In_890);
nand U1843 (N_1843,In_242,In_1090);
xor U1844 (N_1844,In_1049,In_572);
and U1845 (N_1845,In_856,In_505);
nand U1846 (N_1846,In_627,In_941);
nand U1847 (N_1847,In_1043,In_530);
and U1848 (N_1848,In_823,In_1364);
or U1849 (N_1849,In_1465,In_1072);
nor U1850 (N_1850,In_917,In_1332);
or U1851 (N_1851,In_1402,In_59);
nor U1852 (N_1852,In_1012,In_904);
nand U1853 (N_1853,In_1053,In_1033);
xnor U1854 (N_1854,In_1402,In_1114);
nand U1855 (N_1855,In_860,In_149);
and U1856 (N_1856,In_1007,In_592);
nor U1857 (N_1857,In_67,In_258);
or U1858 (N_1858,In_1302,In_1021);
nand U1859 (N_1859,In_1116,In_351);
nand U1860 (N_1860,In_1489,In_557);
nand U1861 (N_1861,In_828,In_1304);
and U1862 (N_1862,In_448,In_1452);
and U1863 (N_1863,In_1391,In_404);
and U1864 (N_1864,In_983,In_149);
and U1865 (N_1865,In_1145,In_1383);
and U1866 (N_1866,In_1054,In_467);
and U1867 (N_1867,In_145,In_1110);
nor U1868 (N_1868,In_194,In_878);
nor U1869 (N_1869,In_626,In_443);
nand U1870 (N_1870,In_118,In_387);
and U1871 (N_1871,In_0,In_1210);
or U1872 (N_1872,In_891,In_958);
nor U1873 (N_1873,In_684,In_1040);
nor U1874 (N_1874,In_1465,In_856);
and U1875 (N_1875,In_558,In_560);
or U1876 (N_1876,In_999,In_617);
nand U1877 (N_1877,In_853,In_477);
or U1878 (N_1878,In_424,In_25);
nand U1879 (N_1879,In_1268,In_98);
and U1880 (N_1880,In_1432,In_582);
nand U1881 (N_1881,In_1307,In_247);
nor U1882 (N_1882,In_540,In_562);
nor U1883 (N_1883,In_670,In_568);
and U1884 (N_1884,In_462,In_1031);
and U1885 (N_1885,In_369,In_35);
and U1886 (N_1886,In_418,In_308);
or U1887 (N_1887,In_1024,In_1214);
or U1888 (N_1888,In_1297,In_44);
nand U1889 (N_1889,In_1058,In_30);
and U1890 (N_1890,In_1351,In_1400);
xnor U1891 (N_1891,In_882,In_321);
nor U1892 (N_1892,In_231,In_312);
nand U1893 (N_1893,In_588,In_1300);
or U1894 (N_1894,In_1002,In_454);
or U1895 (N_1895,In_932,In_317);
nand U1896 (N_1896,In_1181,In_687);
xor U1897 (N_1897,In_1164,In_514);
and U1898 (N_1898,In_461,In_485);
or U1899 (N_1899,In_266,In_1168);
or U1900 (N_1900,In_135,In_1348);
xor U1901 (N_1901,In_1411,In_638);
nand U1902 (N_1902,In_125,In_692);
and U1903 (N_1903,In_468,In_364);
or U1904 (N_1904,In_998,In_1452);
nand U1905 (N_1905,In_481,In_1149);
and U1906 (N_1906,In_1103,In_1256);
and U1907 (N_1907,In_422,In_935);
or U1908 (N_1908,In_1451,In_366);
and U1909 (N_1909,In_1351,In_1468);
nor U1910 (N_1910,In_977,In_875);
nand U1911 (N_1911,In_749,In_930);
or U1912 (N_1912,In_743,In_1339);
xor U1913 (N_1913,In_254,In_1169);
or U1914 (N_1914,In_342,In_1027);
xor U1915 (N_1915,In_710,In_1154);
nand U1916 (N_1916,In_478,In_1405);
nand U1917 (N_1917,In_1456,In_498);
nor U1918 (N_1918,In_746,In_123);
nor U1919 (N_1919,In_984,In_1257);
nor U1920 (N_1920,In_325,In_661);
nor U1921 (N_1921,In_235,In_1466);
nand U1922 (N_1922,In_112,In_208);
xor U1923 (N_1923,In_1109,In_905);
and U1924 (N_1924,In_226,In_345);
or U1925 (N_1925,In_548,In_929);
nor U1926 (N_1926,In_1245,In_1194);
and U1927 (N_1927,In_195,In_196);
nor U1928 (N_1928,In_1179,In_17);
nor U1929 (N_1929,In_1107,In_188);
or U1930 (N_1930,In_888,In_68);
or U1931 (N_1931,In_1176,In_836);
xnor U1932 (N_1932,In_1016,In_182);
nor U1933 (N_1933,In_310,In_491);
and U1934 (N_1934,In_1009,In_513);
and U1935 (N_1935,In_14,In_53);
nor U1936 (N_1936,In_579,In_430);
and U1937 (N_1937,In_1212,In_391);
and U1938 (N_1938,In_660,In_1297);
or U1939 (N_1939,In_1480,In_1131);
and U1940 (N_1940,In_1371,In_951);
and U1941 (N_1941,In_770,In_988);
xor U1942 (N_1942,In_153,In_1240);
nand U1943 (N_1943,In_47,In_852);
nand U1944 (N_1944,In_895,In_1457);
or U1945 (N_1945,In_1428,In_1055);
nand U1946 (N_1946,In_1487,In_592);
nor U1947 (N_1947,In_942,In_204);
or U1948 (N_1948,In_573,In_460);
nand U1949 (N_1949,In_831,In_1088);
and U1950 (N_1950,In_1045,In_397);
xnor U1951 (N_1951,In_415,In_127);
nand U1952 (N_1952,In_1149,In_86);
xnor U1953 (N_1953,In_524,In_458);
or U1954 (N_1954,In_824,In_550);
nor U1955 (N_1955,In_771,In_377);
or U1956 (N_1956,In_1403,In_749);
and U1957 (N_1957,In_799,In_206);
nand U1958 (N_1958,In_970,In_766);
or U1959 (N_1959,In_172,In_934);
or U1960 (N_1960,In_634,In_1236);
and U1961 (N_1961,In_1223,In_1131);
or U1962 (N_1962,In_1149,In_303);
or U1963 (N_1963,In_427,In_353);
or U1964 (N_1964,In_874,In_1416);
nor U1965 (N_1965,In_168,In_520);
nand U1966 (N_1966,In_1107,In_495);
nor U1967 (N_1967,In_1002,In_569);
nand U1968 (N_1968,In_975,In_525);
or U1969 (N_1969,In_541,In_1213);
nand U1970 (N_1970,In_1128,In_577);
nand U1971 (N_1971,In_857,In_1477);
nor U1972 (N_1972,In_780,In_1247);
or U1973 (N_1973,In_1371,In_317);
nor U1974 (N_1974,In_582,In_681);
nor U1975 (N_1975,In_1241,In_338);
nor U1976 (N_1976,In_770,In_1324);
nor U1977 (N_1977,In_795,In_334);
nor U1978 (N_1978,In_454,In_1110);
nand U1979 (N_1979,In_1379,In_1056);
xnor U1980 (N_1980,In_1311,In_1400);
or U1981 (N_1981,In_775,In_432);
or U1982 (N_1982,In_913,In_301);
nor U1983 (N_1983,In_802,In_733);
xor U1984 (N_1984,In_76,In_1005);
or U1985 (N_1985,In_27,In_1376);
and U1986 (N_1986,In_183,In_1222);
nand U1987 (N_1987,In_1360,In_249);
nor U1988 (N_1988,In_215,In_626);
nand U1989 (N_1989,In_1355,In_1029);
or U1990 (N_1990,In_387,In_920);
or U1991 (N_1991,In_744,In_692);
nor U1992 (N_1992,In_501,In_283);
or U1993 (N_1993,In_378,In_852);
or U1994 (N_1994,In_996,In_880);
and U1995 (N_1995,In_947,In_773);
nand U1996 (N_1996,In_319,In_1190);
nand U1997 (N_1997,In_415,In_20);
and U1998 (N_1998,In_987,In_1094);
nor U1999 (N_1999,In_368,In_173);
nor U2000 (N_2000,In_786,In_79);
nand U2001 (N_2001,In_808,In_877);
nand U2002 (N_2002,In_878,In_1439);
nand U2003 (N_2003,In_78,In_901);
nand U2004 (N_2004,In_710,In_618);
nor U2005 (N_2005,In_1431,In_1469);
nand U2006 (N_2006,In_1266,In_1281);
nor U2007 (N_2007,In_1480,In_1203);
nand U2008 (N_2008,In_521,In_327);
xnor U2009 (N_2009,In_893,In_251);
and U2010 (N_2010,In_86,In_301);
and U2011 (N_2011,In_694,In_1273);
or U2012 (N_2012,In_1450,In_1219);
or U2013 (N_2013,In_358,In_221);
or U2014 (N_2014,In_365,In_1271);
nand U2015 (N_2015,In_1306,In_288);
nand U2016 (N_2016,In_1128,In_1261);
or U2017 (N_2017,In_710,In_215);
nor U2018 (N_2018,In_482,In_264);
nand U2019 (N_2019,In_1031,In_243);
nor U2020 (N_2020,In_309,In_1064);
or U2021 (N_2021,In_1057,In_19);
nor U2022 (N_2022,In_146,In_1132);
and U2023 (N_2023,In_498,In_110);
nand U2024 (N_2024,In_1202,In_1208);
and U2025 (N_2025,In_227,In_183);
xor U2026 (N_2026,In_498,In_887);
xor U2027 (N_2027,In_303,In_992);
xnor U2028 (N_2028,In_1434,In_232);
or U2029 (N_2029,In_859,In_639);
and U2030 (N_2030,In_887,In_649);
or U2031 (N_2031,In_190,In_104);
or U2032 (N_2032,In_816,In_926);
nand U2033 (N_2033,In_677,In_70);
and U2034 (N_2034,In_524,In_964);
nand U2035 (N_2035,In_128,In_1253);
and U2036 (N_2036,In_931,In_177);
and U2037 (N_2037,In_72,In_603);
nand U2038 (N_2038,In_285,In_63);
xnor U2039 (N_2039,In_1475,In_1464);
nand U2040 (N_2040,In_1007,In_717);
and U2041 (N_2041,In_278,In_1209);
xnor U2042 (N_2042,In_739,In_371);
nand U2043 (N_2043,In_579,In_764);
nand U2044 (N_2044,In_285,In_148);
xnor U2045 (N_2045,In_820,In_901);
and U2046 (N_2046,In_935,In_1442);
nor U2047 (N_2047,In_212,In_853);
and U2048 (N_2048,In_803,In_1251);
and U2049 (N_2049,In_212,In_1121);
nand U2050 (N_2050,In_1069,In_305);
nand U2051 (N_2051,In_571,In_1021);
and U2052 (N_2052,In_1090,In_25);
nand U2053 (N_2053,In_1294,In_389);
nand U2054 (N_2054,In_300,In_481);
xnor U2055 (N_2055,In_702,In_65);
nand U2056 (N_2056,In_346,In_170);
nand U2057 (N_2057,In_678,In_179);
nor U2058 (N_2058,In_1054,In_1157);
or U2059 (N_2059,In_892,In_258);
nor U2060 (N_2060,In_1419,In_682);
and U2061 (N_2061,In_520,In_679);
xor U2062 (N_2062,In_1344,In_1127);
and U2063 (N_2063,In_381,In_54);
nor U2064 (N_2064,In_925,In_508);
nor U2065 (N_2065,In_942,In_362);
and U2066 (N_2066,In_1240,In_1412);
and U2067 (N_2067,In_823,In_905);
nand U2068 (N_2068,In_1211,In_286);
nor U2069 (N_2069,In_912,In_1475);
nor U2070 (N_2070,In_1057,In_437);
nor U2071 (N_2071,In_581,In_134);
and U2072 (N_2072,In_652,In_1030);
and U2073 (N_2073,In_788,In_292);
and U2074 (N_2074,In_790,In_126);
xnor U2075 (N_2075,In_532,In_1343);
or U2076 (N_2076,In_13,In_66);
or U2077 (N_2077,In_790,In_753);
nand U2078 (N_2078,In_670,In_476);
nand U2079 (N_2079,In_1326,In_354);
or U2080 (N_2080,In_1119,In_1051);
and U2081 (N_2081,In_1374,In_196);
nand U2082 (N_2082,In_41,In_1249);
or U2083 (N_2083,In_625,In_621);
and U2084 (N_2084,In_1257,In_1119);
nand U2085 (N_2085,In_44,In_165);
and U2086 (N_2086,In_1354,In_1466);
or U2087 (N_2087,In_353,In_1000);
and U2088 (N_2088,In_1459,In_631);
nand U2089 (N_2089,In_1123,In_607);
and U2090 (N_2090,In_1097,In_180);
nand U2091 (N_2091,In_632,In_104);
nor U2092 (N_2092,In_351,In_538);
and U2093 (N_2093,In_34,In_1217);
and U2094 (N_2094,In_612,In_888);
and U2095 (N_2095,In_615,In_423);
and U2096 (N_2096,In_467,In_846);
nand U2097 (N_2097,In_496,In_1309);
nand U2098 (N_2098,In_1044,In_1072);
and U2099 (N_2099,In_296,In_1353);
and U2100 (N_2100,In_1323,In_540);
xnor U2101 (N_2101,In_480,In_1068);
nand U2102 (N_2102,In_1296,In_545);
nor U2103 (N_2103,In_924,In_171);
or U2104 (N_2104,In_1451,In_152);
or U2105 (N_2105,In_59,In_100);
nor U2106 (N_2106,In_645,In_1072);
or U2107 (N_2107,In_761,In_881);
nor U2108 (N_2108,In_52,In_743);
or U2109 (N_2109,In_925,In_119);
and U2110 (N_2110,In_1167,In_671);
nand U2111 (N_2111,In_1475,In_874);
and U2112 (N_2112,In_1080,In_693);
nor U2113 (N_2113,In_560,In_638);
xnor U2114 (N_2114,In_977,In_322);
xnor U2115 (N_2115,In_892,In_1125);
or U2116 (N_2116,In_1020,In_200);
xor U2117 (N_2117,In_1168,In_733);
or U2118 (N_2118,In_1443,In_1316);
xor U2119 (N_2119,In_297,In_1100);
nand U2120 (N_2120,In_349,In_1145);
xnor U2121 (N_2121,In_1119,In_1456);
or U2122 (N_2122,In_836,In_291);
and U2123 (N_2123,In_730,In_760);
nor U2124 (N_2124,In_136,In_1146);
nand U2125 (N_2125,In_609,In_1084);
and U2126 (N_2126,In_914,In_963);
or U2127 (N_2127,In_1341,In_505);
or U2128 (N_2128,In_1233,In_572);
nor U2129 (N_2129,In_195,In_329);
and U2130 (N_2130,In_1220,In_269);
nand U2131 (N_2131,In_1182,In_411);
or U2132 (N_2132,In_9,In_1465);
nor U2133 (N_2133,In_475,In_1041);
or U2134 (N_2134,In_928,In_474);
nand U2135 (N_2135,In_1487,In_885);
nand U2136 (N_2136,In_1160,In_643);
nand U2137 (N_2137,In_605,In_299);
nand U2138 (N_2138,In_891,In_550);
nor U2139 (N_2139,In_558,In_1008);
nand U2140 (N_2140,In_365,In_491);
and U2141 (N_2141,In_727,In_423);
nor U2142 (N_2142,In_685,In_123);
nand U2143 (N_2143,In_221,In_263);
and U2144 (N_2144,In_3,In_1221);
or U2145 (N_2145,In_409,In_639);
or U2146 (N_2146,In_1198,In_1290);
nand U2147 (N_2147,In_1104,In_205);
nor U2148 (N_2148,In_515,In_151);
nand U2149 (N_2149,In_1055,In_1199);
or U2150 (N_2150,In_306,In_471);
or U2151 (N_2151,In_605,In_792);
nand U2152 (N_2152,In_1069,In_1036);
or U2153 (N_2153,In_1040,In_362);
xnor U2154 (N_2154,In_1117,In_1004);
or U2155 (N_2155,In_1212,In_1421);
and U2156 (N_2156,In_767,In_534);
and U2157 (N_2157,In_113,In_1162);
and U2158 (N_2158,In_1440,In_622);
nand U2159 (N_2159,In_535,In_1244);
and U2160 (N_2160,In_1235,In_257);
and U2161 (N_2161,In_743,In_1388);
or U2162 (N_2162,In_1240,In_470);
and U2163 (N_2163,In_1105,In_306);
nand U2164 (N_2164,In_1133,In_757);
and U2165 (N_2165,In_1062,In_21);
nor U2166 (N_2166,In_706,In_1216);
and U2167 (N_2167,In_1127,In_109);
or U2168 (N_2168,In_1161,In_1186);
xnor U2169 (N_2169,In_180,In_1443);
nor U2170 (N_2170,In_1270,In_965);
and U2171 (N_2171,In_682,In_157);
and U2172 (N_2172,In_1476,In_1006);
nor U2173 (N_2173,In_145,In_877);
xnor U2174 (N_2174,In_1350,In_307);
xnor U2175 (N_2175,In_232,In_1255);
xor U2176 (N_2176,In_177,In_695);
or U2177 (N_2177,In_817,In_47);
and U2178 (N_2178,In_1145,In_1318);
nand U2179 (N_2179,In_1192,In_104);
and U2180 (N_2180,In_91,In_1354);
nor U2181 (N_2181,In_1230,In_1414);
xnor U2182 (N_2182,In_316,In_918);
xor U2183 (N_2183,In_1021,In_348);
nor U2184 (N_2184,In_413,In_1308);
nand U2185 (N_2185,In_605,In_624);
nand U2186 (N_2186,In_802,In_172);
and U2187 (N_2187,In_1341,In_1105);
or U2188 (N_2188,In_92,In_112);
xor U2189 (N_2189,In_624,In_950);
and U2190 (N_2190,In_1183,In_101);
xnor U2191 (N_2191,In_82,In_890);
nand U2192 (N_2192,In_598,In_490);
or U2193 (N_2193,In_680,In_676);
nand U2194 (N_2194,In_459,In_192);
or U2195 (N_2195,In_201,In_1022);
nor U2196 (N_2196,In_663,In_419);
or U2197 (N_2197,In_692,In_748);
or U2198 (N_2198,In_36,In_454);
nor U2199 (N_2199,In_789,In_1092);
nor U2200 (N_2200,In_1472,In_1298);
or U2201 (N_2201,In_76,In_1136);
nor U2202 (N_2202,In_450,In_521);
or U2203 (N_2203,In_943,In_944);
nor U2204 (N_2204,In_7,In_1322);
or U2205 (N_2205,In_884,In_1419);
and U2206 (N_2206,In_204,In_151);
or U2207 (N_2207,In_305,In_1456);
and U2208 (N_2208,In_956,In_214);
and U2209 (N_2209,In_1113,In_114);
nand U2210 (N_2210,In_259,In_957);
nor U2211 (N_2211,In_591,In_167);
nand U2212 (N_2212,In_1293,In_465);
nor U2213 (N_2213,In_1251,In_122);
and U2214 (N_2214,In_1249,In_1497);
nor U2215 (N_2215,In_668,In_86);
or U2216 (N_2216,In_1387,In_984);
nand U2217 (N_2217,In_1214,In_1381);
or U2218 (N_2218,In_239,In_639);
nor U2219 (N_2219,In_814,In_618);
nor U2220 (N_2220,In_839,In_807);
nand U2221 (N_2221,In_1127,In_590);
or U2222 (N_2222,In_1439,In_303);
nand U2223 (N_2223,In_1380,In_1335);
and U2224 (N_2224,In_886,In_1134);
and U2225 (N_2225,In_252,In_985);
and U2226 (N_2226,In_22,In_328);
or U2227 (N_2227,In_417,In_1034);
and U2228 (N_2228,In_537,In_661);
nand U2229 (N_2229,In_507,In_497);
nand U2230 (N_2230,In_1079,In_805);
nand U2231 (N_2231,In_787,In_461);
or U2232 (N_2232,In_1394,In_561);
or U2233 (N_2233,In_942,In_659);
nand U2234 (N_2234,In_22,In_599);
and U2235 (N_2235,In_1173,In_297);
nand U2236 (N_2236,In_246,In_396);
nor U2237 (N_2237,In_1186,In_287);
xor U2238 (N_2238,In_280,In_1462);
and U2239 (N_2239,In_1435,In_979);
xnor U2240 (N_2240,In_1086,In_1095);
nand U2241 (N_2241,In_718,In_350);
and U2242 (N_2242,In_891,In_1023);
nor U2243 (N_2243,In_468,In_1290);
or U2244 (N_2244,In_338,In_1318);
nor U2245 (N_2245,In_1448,In_650);
and U2246 (N_2246,In_1226,In_86);
nor U2247 (N_2247,In_898,In_782);
nor U2248 (N_2248,In_818,In_581);
nand U2249 (N_2249,In_1054,In_1384);
nor U2250 (N_2250,In_1066,In_811);
or U2251 (N_2251,In_135,In_404);
and U2252 (N_2252,In_815,In_1199);
or U2253 (N_2253,In_705,In_1246);
and U2254 (N_2254,In_195,In_1251);
nor U2255 (N_2255,In_827,In_74);
nand U2256 (N_2256,In_888,In_568);
xnor U2257 (N_2257,In_1290,In_618);
xnor U2258 (N_2258,In_1364,In_1425);
and U2259 (N_2259,In_1205,In_658);
or U2260 (N_2260,In_517,In_763);
nor U2261 (N_2261,In_2,In_262);
nand U2262 (N_2262,In_1023,In_1429);
or U2263 (N_2263,In_696,In_1375);
or U2264 (N_2264,In_799,In_1130);
nor U2265 (N_2265,In_1224,In_536);
and U2266 (N_2266,In_1479,In_513);
xnor U2267 (N_2267,In_807,In_1170);
nor U2268 (N_2268,In_1278,In_677);
xnor U2269 (N_2269,In_311,In_138);
nand U2270 (N_2270,In_1036,In_80);
xnor U2271 (N_2271,In_451,In_1272);
or U2272 (N_2272,In_625,In_372);
and U2273 (N_2273,In_73,In_859);
nand U2274 (N_2274,In_1458,In_1442);
nor U2275 (N_2275,In_868,In_303);
and U2276 (N_2276,In_1095,In_1317);
and U2277 (N_2277,In_1221,In_297);
nor U2278 (N_2278,In_1431,In_1412);
and U2279 (N_2279,In_812,In_906);
nor U2280 (N_2280,In_1127,In_449);
and U2281 (N_2281,In_707,In_792);
nand U2282 (N_2282,In_661,In_849);
or U2283 (N_2283,In_1424,In_1098);
nand U2284 (N_2284,In_809,In_1453);
or U2285 (N_2285,In_60,In_345);
or U2286 (N_2286,In_131,In_1065);
and U2287 (N_2287,In_207,In_839);
or U2288 (N_2288,In_818,In_921);
and U2289 (N_2289,In_1446,In_368);
nand U2290 (N_2290,In_1000,In_747);
nor U2291 (N_2291,In_1444,In_1225);
nor U2292 (N_2292,In_910,In_992);
nor U2293 (N_2293,In_882,In_203);
and U2294 (N_2294,In_1261,In_95);
nor U2295 (N_2295,In_721,In_613);
or U2296 (N_2296,In_689,In_1340);
or U2297 (N_2297,In_1079,In_818);
and U2298 (N_2298,In_1405,In_1315);
nor U2299 (N_2299,In_938,In_144);
and U2300 (N_2300,In_22,In_661);
nand U2301 (N_2301,In_85,In_653);
nand U2302 (N_2302,In_619,In_1387);
or U2303 (N_2303,In_600,In_975);
and U2304 (N_2304,In_570,In_215);
xnor U2305 (N_2305,In_492,In_582);
or U2306 (N_2306,In_432,In_286);
nand U2307 (N_2307,In_841,In_292);
and U2308 (N_2308,In_49,In_407);
or U2309 (N_2309,In_182,In_887);
or U2310 (N_2310,In_213,In_798);
nand U2311 (N_2311,In_585,In_670);
nand U2312 (N_2312,In_399,In_339);
or U2313 (N_2313,In_383,In_1051);
and U2314 (N_2314,In_839,In_1339);
xor U2315 (N_2315,In_1117,In_1015);
nand U2316 (N_2316,In_1393,In_1112);
and U2317 (N_2317,In_421,In_236);
xnor U2318 (N_2318,In_1217,In_754);
nor U2319 (N_2319,In_650,In_505);
nor U2320 (N_2320,In_1178,In_756);
nand U2321 (N_2321,In_378,In_996);
nor U2322 (N_2322,In_1271,In_644);
xor U2323 (N_2323,In_372,In_1385);
nor U2324 (N_2324,In_266,In_17);
or U2325 (N_2325,In_1271,In_702);
and U2326 (N_2326,In_541,In_287);
nand U2327 (N_2327,In_657,In_1002);
or U2328 (N_2328,In_1320,In_111);
nor U2329 (N_2329,In_364,In_1148);
nor U2330 (N_2330,In_1361,In_1313);
and U2331 (N_2331,In_917,In_826);
nor U2332 (N_2332,In_1201,In_361);
and U2333 (N_2333,In_1107,In_1395);
nand U2334 (N_2334,In_486,In_1392);
or U2335 (N_2335,In_1250,In_413);
nor U2336 (N_2336,In_636,In_305);
nor U2337 (N_2337,In_247,In_117);
nand U2338 (N_2338,In_1363,In_879);
and U2339 (N_2339,In_106,In_1);
nor U2340 (N_2340,In_706,In_1289);
or U2341 (N_2341,In_1429,In_325);
nor U2342 (N_2342,In_540,In_1374);
or U2343 (N_2343,In_929,In_226);
and U2344 (N_2344,In_327,In_1491);
nor U2345 (N_2345,In_417,In_804);
and U2346 (N_2346,In_1304,In_5);
nor U2347 (N_2347,In_1189,In_438);
xnor U2348 (N_2348,In_237,In_928);
nor U2349 (N_2349,In_648,In_524);
or U2350 (N_2350,In_530,In_567);
or U2351 (N_2351,In_1284,In_1123);
nor U2352 (N_2352,In_550,In_1235);
nor U2353 (N_2353,In_184,In_562);
or U2354 (N_2354,In_590,In_1477);
nor U2355 (N_2355,In_1104,In_761);
and U2356 (N_2356,In_1430,In_912);
nand U2357 (N_2357,In_5,In_1085);
or U2358 (N_2358,In_702,In_669);
and U2359 (N_2359,In_849,In_156);
nor U2360 (N_2360,In_364,In_1431);
and U2361 (N_2361,In_121,In_543);
nand U2362 (N_2362,In_359,In_1010);
and U2363 (N_2363,In_1195,In_259);
xnor U2364 (N_2364,In_1450,In_491);
and U2365 (N_2365,In_687,In_412);
nor U2366 (N_2366,In_1213,In_998);
or U2367 (N_2367,In_962,In_153);
nand U2368 (N_2368,In_939,In_785);
nand U2369 (N_2369,In_384,In_516);
nor U2370 (N_2370,In_1346,In_1048);
and U2371 (N_2371,In_855,In_14);
and U2372 (N_2372,In_370,In_815);
nor U2373 (N_2373,In_215,In_1281);
or U2374 (N_2374,In_1196,In_1191);
or U2375 (N_2375,In_565,In_176);
nand U2376 (N_2376,In_1256,In_1333);
nor U2377 (N_2377,In_827,In_580);
nand U2378 (N_2378,In_1367,In_783);
or U2379 (N_2379,In_1134,In_910);
or U2380 (N_2380,In_874,In_495);
or U2381 (N_2381,In_7,In_27);
or U2382 (N_2382,In_567,In_848);
or U2383 (N_2383,In_1398,In_955);
nor U2384 (N_2384,In_135,In_599);
or U2385 (N_2385,In_877,In_652);
or U2386 (N_2386,In_719,In_1257);
nor U2387 (N_2387,In_1406,In_203);
or U2388 (N_2388,In_880,In_1006);
and U2389 (N_2389,In_1463,In_119);
nor U2390 (N_2390,In_1462,In_616);
xnor U2391 (N_2391,In_194,In_722);
and U2392 (N_2392,In_580,In_78);
and U2393 (N_2393,In_630,In_1261);
and U2394 (N_2394,In_306,In_728);
nor U2395 (N_2395,In_1498,In_452);
and U2396 (N_2396,In_436,In_248);
nor U2397 (N_2397,In_1074,In_973);
and U2398 (N_2398,In_931,In_1344);
nor U2399 (N_2399,In_60,In_599);
and U2400 (N_2400,In_1116,In_693);
nand U2401 (N_2401,In_1161,In_162);
and U2402 (N_2402,In_1040,In_326);
nor U2403 (N_2403,In_1223,In_598);
xor U2404 (N_2404,In_991,In_1457);
or U2405 (N_2405,In_384,In_394);
nor U2406 (N_2406,In_272,In_1374);
and U2407 (N_2407,In_1416,In_870);
xnor U2408 (N_2408,In_145,In_1302);
or U2409 (N_2409,In_202,In_461);
or U2410 (N_2410,In_1478,In_1025);
nand U2411 (N_2411,In_845,In_1156);
nor U2412 (N_2412,In_957,In_309);
xnor U2413 (N_2413,In_403,In_1346);
or U2414 (N_2414,In_1079,In_373);
xnor U2415 (N_2415,In_992,In_405);
nor U2416 (N_2416,In_565,In_42);
nor U2417 (N_2417,In_336,In_948);
or U2418 (N_2418,In_905,In_997);
and U2419 (N_2419,In_1107,In_496);
xnor U2420 (N_2420,In_1106,In_1406);
and U2421 (N_2421,In_418,In_323);
nand U2422 (N_2422,In_569,In_119);
and U2423 (N_2423,In_138,In_102);
nor U2424 (N_2424,In_600,In_683);
nand U2425 (N_2425,In_1204,In_607);
nand U2426 (N_2426,In_1040,In_1162);
nor U2427 (N_2427,In_353,In_620);
and U2428 (N_2428,In_637,In_358);
and U2429 (N_2429,In_1499,In_602);
nand U2430 (N_2430,In_1132,In_1076);
nand U2431 (N_2431,In_934,In_1011);
nor U2432 (N_2432,In_1028,In_505);
nand U2433 (N_2433,In_1228,In_282);
nand U2434 (N_2434,In_361,In_1115);
nor U2435 (N_2435,In_1087,In_542);
and U2436 (N_2436,In_767,In_471);
or U2437 (N_2437,In_572,In_576);
and U2438 (N_2438,In_1220,In_853);
and U2439 (N_2439,In_784,In_1087);
nor U2440 (N_2440,In_670,In_319);
nand U2441 (N_2441,In_885,In_1111);
nand U2442 (N_2442,In_1240,In_1493);
nand U2443 (N_2443,In_1438,In_979);
or U2444 (N_2444,In_1315,In_1303);
nor U2445 (N_2445,In_804,In_504);
or U2446 (N_2446,In_1457,In_363);
nor U2447 (N_2447,In_1372,In_1094);
and U2448 (N_2448,In_1404,In_382);
nand U2449 (N_2449,In_1202,In_1408);
and U2450 (N_2450,In_1309,In_694);
nor U2451 (N_2451,In_1178,In_77);
and U2452 (N_2452,In_368,In_187);
nand U2453 (N_2453,In_187,In_992);
nor U2454 (N_2454,In_1336,In_744);
or U2455 (N_2455,In_907,In_1212);
or U2456 (N_2456,In_1170,In_875);
and U2457 (N_2457,In_1380,In_895);
xor U2458 (N_2458,In_47,In_378);
nand U2459 (N_2459,In_1221,In_699);
nand U2460 (N_2460,In_899,In_915);
nand U2461 (N_2461,In_1262,In_1160);
and U2462 (N_2462,In_942,In_1176);
or U2463 (N_2463,In_1227,In_394);
nand U2464 (N_2464,In_1338,In_478);
nor U2465 (N_2465,In_320,In_794);
or U2466 (N_2466,In_1069,In_828);
and U2467 (N_2467,In_1376,In_801);
and U2468 (N_2468,In_1354,In_68);
or U2469 (N_2469,In_797,In_244);
nor U2470 (N_2470,In_768,In_1102);
xnor U2471 (N_2471,In_1206,In_724);
nand U2472 (N_2472,In_83,In_1143);
nand U2473 (N_2473,In_1019,In_959);
and U2474 (N_2474,In_81,In_446);
nor U2475 (N_2475,In_1372,In_1379);
xor U2476 (N_2476,In_961,In_847);
or U2477 (N_2477,In_477,In_78);
or U2478 (N_2478,In_210,In_1172);
nand U2479 (N_2479,In_1384,In_919);
or U2480 (N_2480,In_326,In_559);
nand U2481 (N_2481,In_637,In_1106);
nor U2482 (N_2482,In_1063,In_105);
and U2483 (N_2483,In_431,In_244);
nand U2484 (N_2484,In_281,In_1029);
nand U2485 (N_2485,In_948,In_815);
or U2486 (N_2486,In_904,In_1207);
xor U2487 (N_2487,In_479,In_14);
and U2488 (N_2488,In_641,In_609);
or U2489 (N_2489,In_1488,In_117);
xnor U2490 (N_2490,In_803,In_1201);
nor U2491 (N_2491,In_1185,In_625);
nor U2492 (N_2492,In_1100,In_1122);
nand U2493 (N_2493,In_550,In_438);
nor U2494 (N_2494,In_888,In_1418);
and U2495 (N_2495,In_405,In_1470);
and U2496 (N_2496,In_294,In_603);
nor U2497 (N_2497,In_49,In_1109);
nor U2498 (N_2498,In_206,In_287);
and U2499 (N_2499,In_1157,In_910);
nand U2500 (N_2500,In_5,In_1083);
xnor U2501 (N_2501,In_1001,In_813);
nor U2502 (N_2502,In_690,In_1221);
and U2503 (N_2503,In_1417,In_1276);
xnor U2504 (N_2504,In_355,In_1002);
nand U2505 (N_2505,In_1104,In_241);
or U2506 (N_2506,In_389,In_654);
nor U2507 (N_2507,In_1045,In_10);
xnor U2508 (N_2508,In_727,In_1450);
and U2509 (N_2509,In_1330,In_495);
and U2510 (N_2510,In_1362,In_263);
or U2511 (N_2511,In_395,In_261);
or U2512 (N_2512,In_164,In_1316);
nor U2513 (N_2513,In_270,In_724);
nand U2514 (N_2514,In_1010,In_1303);
nand U2515 (N_2515,In_216,In_1079);
nor U2516 (N_2516,In_738,In_304);
nor U2517 (N_2517,In_706,In_417);
nor U2518 (N_2518,In_673,In_513);
or U2519 (N_2519,In_1130,In_469);
nor U2520 (N_2520,In_646,In_650);
xor U2521 (N_2521,In_1307,In_1341);
nor U2522 (N_2522,In_1403,In_993);
xnor U2523 (N_2523,In_1053,In_1320);
and U2524 (N_2524,In_1435,In_632);
or U2525 (N_2525,In_756,In_807);
nor U2526 (N_2526,In_1067,In_1449);
or U2527 (N_2527,In_98,In_642);
nand U2528 (N_2528,In_1230,In_1282);
or U2529 (N_2529,In_449,In_1317);
and U2530 (N_2530,In_141,In_480);
or U2531 (N_2531,In_1458,In_335);
and U2532 (N_2532,In_1368,In_335);
and U2533 (N_2533,In_1047,In_1139);
and U2534 (N_2534,In_1346,In_1405);
nand U2535 (N_2535,In_963,In_171);
nand U2536 (N_2536,In_1296,In_864);
nand U2537 (N_2537,In_185,In_1078);
nand U2538 (N_2538,In_1122,In_1281);
and U2539 (N_2539,In_61,In_1142);
nand U2540 (N_2540,In_165,In_87);
and U2541 (N_2541,In_1423,In_652);
and U2542 (N_2542,In_175,In_278);
nor U2543 (N_2543,In_748,In_787);
nand U2544 (N_2544,In_1279,In_1058);
nor U2545 (N_2545,In_597,In_21);
nand U2546 (N_2546,In_69,In_991);
or U2547 (N_2547,In_1474,In_1000);
nand U2548 (N_2548,In_772,In_290);
nand U2549 (N_2549,In_690,In_1467);
and U2550 (N_2550,In_272,In_1010);
nor U2551 (N_2551,In_168,In_496);
and U2552 (N_2552,In_878,In_75);
nor U2553 (N_2553,In_939,In_1433);
and U2554 (N_2554,In_736,In_1313);
xnor U2555 (N_2555,In_884,In_272);
and U2556 (N_2556,In_319,In_202);
nand U2557 (N_2557,In_239,In_694);
nor U2558 (N_2558,In_1465,In_673);
nand U2559 (N_2559,In_1262,In_396);
nor U2560 (N_2560,In_472,In_458);
or U2561 (N_2561,In_1283,In_1291);
xor U2562 (N_2562,In_514,In_325);
or U2563 (N_2563,In_883,In_595);
nor U2564 (N_2564,In_1163,In_708);
or U2565 (N_2565,In_1116,In_929);
nor U2566 (N_2566,In_1070,In_8);
or U2567 (N_2567,In_348,In_160);
or U2568 (N_2568,In_284,In_320);
nand U2569 (N_2569,In_110,In_1091);
nor U2570 (N_2570,In_955,In_620);
and U2571 (N_2571,In_699,In_406);
and U2572 (N_2572,In_293,In_351);
nand U2573 (N_2573,In_831,In_1062);
and U2574 (N_2574,In_1358,In_636);
nor U2575 (N_2575,In_172,In_623);
nor U2576 (N_2576,In_1264,In_381);
or U2577 (N_2577,In_25,In_381);
nand U2578 (N_2578,In_363,In_1415);
nor U2579 (N_2579,In_662,In_974);
nor U2580 (N_2580,In_1331,In_327);
xor U2581 (N_2581,In_962,In_1473);
xor U2582 (N_2582,In_932,In_1399);
and U2583 (N_2583,In_906,In_1030);
xor U2584 (N_2584,In_434,In_1438);
and U2585 (N_2585,In_1351,In_42);
and U2586 (N_2586,In_715,In_1209);
or U2587 (N_2587,In_810,In_1052);
and U2588 (N_2588,In_1267,In_1101);
xnor U2589 (N_2589,In_592,In_1110);
and U2590 (N_2590,In_732,In_201);
or U2591 (N_2591,In_454,In_1331);
or U2592 (N_2592,In_217,In_652);
or U2593 (N_2593,In_1337,In_693);
or U2594 (N_2594,In_1241,In_1344);
and U2595 (N_2595,In_411,In_583);
nor U2596 (N_2596,In_782,In_1115);
nand U2597 (N_2597,In_920,In_472);
or U2598 (N_2598,In_925,In_1059);
and U2599 (N_2599,In_46,In_536);
nand U2600 (N_2600,In_1047,In_1430);
and U2601 (N_2601,In_1006,In_22);
nand U2602 (N_2602,In_724,In_966);
nand U2603 (N_2603,In_167,In_977);
xnor U2604 (N_2604,In_313,In_650);
and U2605 (N_2605,In_841,In_752);
nand U2606 (N_2606,In_1371,In_43);
nor U2607 (N_2607,In_984,In_985);
nand U2608 (N_2608,In_875,In_138);
or U2609 (N_2609,In_503,In_1180);
or U2610 (N_2610,In_1397,In_436);
or U2611 (N_2611,In_816,In_188);
xnor U2612 (N_2612,In_899,In_352);
nor U2613 (N_2613,In_338,In_1414);
nor U2614 (N_2614,In_736,In_1302);
and U2615 (N_2615,In_238,In_282);
nor U2616 (N_2616,In_720,In_880);
or U2617 (N_2617,In_583,In_492);
and U2618 (N_2618,In_304,In_363);
nand U2619 (N_2619,In_541,In_1031);
nand U2620 (N_2620,In_719,In_1460);
nor U2621 (N_2621,In_62,In_503);
or U2622 (N_2622,In_221,In_1272);
nor U2623 (N_2623,In_988,In_990);
nand U2624 (N_2624,In_756,In_660);
nand U2625 (N_2625,In_636,In_1112);
nor U2626 (N_2626,In_1313,In_1108);
nand U2627 (N_2627,In_1107,In_1375);
nand U2628 (N_2628,In_1329,In_780);
or U2629 (N_2629,In_976,In_1281);
nor U2630 (N_2630,In_878,In_320);
and U2631 (N_2631,In_433,In_1058);
and U2632 (N_2632,In_382,In_585);
or U2633 (N_2633,In_1401,In_579);
and U2634 (N_2634,In_206,In_1056);
nor U2635 (N_2635,In_1273,In_33);
nand U2636 (N_2636,In_97,In_750);
nor U2637 (N_2637,In_421,In_1060);
nand U2638 (N_2638,In_972,In_936);
nand U2639 (N_2639,In_518,In_450);
and U2640 (N_2640,In_56,In_937);
nor U2641 (N_2641,In_943,In_366);
xor U2642 (N_2642,In_8,In_614);
and U2643 (N_2643,In_359,In_430);
nand U2644 (N_2644,In_1208,In_294);
nand U2645 (N_2645,In_1117,In_205);
or U2646 (N_2646,In_1018,In_205);
or U2647 (N_2647,In_1480,In_286);
nand U2648 (N_2648,In_1376,In_1391);
nand U2649 (N_2649,In_733,In_467);
and U2650 (N_2650,In_1322,In_482);
nand U2651 (N_2651,In_574,In_277);
nand U2652 (N_2652,In_1177,In_93);
and U2653 (N_2653,In_1169,In_270);
nor U2654 (N_2654,In_1169,In_249);
xor U2655 (N_2655,In_1418,In_785);
nor U2656 (N_2656,In_248,In_937);
or U2657 (N_2657,In_849,In_1189);
xor U2658 (N_2658,In_1071,In_434);
nor U2659 (N_2659,In_996,In_16);
and U2660 (N_2660,In_150,In_759);
nand U2661 (N_2661,In_855,In_131);
nand U2662 (N_2662,In_321,In_976);
xor U2663 (N_2663,In_1381,In_755);
xnor U2664 (N_2664,In_536,In_1032);
xnor U2665 (N_2665,In_1430,In_217);
nand U2666 (N_2666,In_362,In_816);
nor U2667 (N_2667,In_330,In_1319);
nor U2668 (N_2668,In_177,In_1443);
nor U2669 (N_2669,In_613,In_1325);
or U2670 (N_2670,In_1474,In_830);
or U2671 (N_2671,In_124,In_313);
nor U2672 (N_2672,In_973,In_212);
and U2673 (N_2673,In_146,In_303);
or U2674 (N_2674,In_1427,In_729);
nand U2675 (N_2675,In_1191,In_508);
xor U2676 (N_2676,In_1461,In_355);
and U2677 (N_2677,In_1141,In_75);
nor U2678 (N_2678,In_1032,In_1416);
or U2679 (N_2679,In_987,In_474);
xnor U2680 (N_2680,In_678,In_326);
nand U2681 (N_2681,In_507,In_216);
and U2682 (N_2682,In_1154,In_891);
or U2683 (N_2683,In_1308,In_294);
nor U2684 (N_2684,In_1264,In_1381);
nor U2685 (N_2685,In_856,In_396);
nor U2686 (N_2686,In_583,In_1086);
nor U2687 (N_2687,In_1053,In_607);
or U2688 (N_2688,In_572,In_1252);
nand U2689 (N_2689,In_978,In_328);
nand U2690 (N_2690,In_242,In_1428);
or U2691 (N_2691,In_468,In_218);
or U2692 (N_2692,In_941,In_1157);
nor U2693 (N_2693,In_638,In_668);
nand U2694 (N_2694,In_1122,In_606);
nand U2695 (N_2695,In_1215,In_955);
or U2696 (N_2696,In_801,In_276);
nor U2697 (N_2697,In_1320,In_989);
and U2698 (N_2698,In_813,In_745);
and U2699 (N_2699,In_376,In_433);
nor U2700 (N_2700,In_1322,In_1186);
nand U2701 (N_2701,In_855,In_1267);
and U2702 (N_2702,In_643,In_392);
nor U2703 (N_2703,In_1368,In_1107);
nor U2704 (N_2704,In_615,In_1368);
nand U2705 (N_2705,In_1448,In_1322);
and U2706 (N_2706,In_266,In_53);
and U2707 (N_2707,In_1428,In_1225);
or U2708 (N_2708,In_450,In_1002);
nand U2709 (N_2709,In_1077,In_778);
or U2710 (N_2710,In_1343,In_84);
and U2711 (N_2711,In_1083,In_691);
nor U2712 (N_2712,In_1247,In_434);
nand U2713 (N_2713,In_257,In_1418);
xnor U2714 (N_2714,In_1086,In_87);
nand U2715 (N_2715,In_850,In_1235);
and U2716 (N_2716,In_334,In_425);
and U2717 (N_2717,In_1298,In_287);
nor U2718 (N_2718,In_698,In_1449);
nand U2719 (N_2719,In_271,In_893);
and U2720 (N_2720,In_1289,In_471);
or U2721 (N_2721,In_778,In_29);
nor U2722 (N_2722,In_1077,In_1055);
nor U2723 (N_2723,In_520,In_848);
or U2724 (N_2724,In_671,In_1188);
nor U2725 (N_2725,In_367,In_1226);
and U2726 (N_2726,In_512,In_1338);
nor U2727 (N_2727,In_663,In_166);
and U2728 (N_2728,In_1011,In_615);
nand U2729 (N_2729,In_1118,In_1389);
nand U2730 (N_2730,In_1415,In_334);
xnor U2731 (N_2731,In_595,In_312);
xor U2732 (N_2732,In_1154,In_511);
xor U2733 (N_2733,In_1187,In_692);
nand U2734 (N_2734,In_709,In_1064);
and U2735 (N_2735,In_858,In_1425);
and U2736 (N_2736,In_205,In_963);
nor U2737 (N_2737,In_406,In_65);
or U2738 (N_2738,In_1469,In_289);
or U2739 (N_2739,In_308,In_585);
nor U2740 (N_2740,In_471,In_880);
nand U2741 (N_2741,In_429,In_167);
and U2742 (N_2742,In_782,In_588);
nand U2743 (N_2743,In_385,In_80);
nand U2744 (N_2744,In_245,In_1275);
xor U2745 (N_2745,In_914,In_784);
or U2746 (N_2746,In_281,In_881);
and U2747 (N_2747,In_477,In_1254);
or U2748 (N_2748,In_989,In_187);
xor U2749 (N_2749,In_448,In_386);
xor U2750 (N_2750,In_918,In_29);
nand U2751 (N_2751,In_423,In_318);
xor U2752 (N_2752,In_950,In_401);
and U2753 (N_2753,In_218,In_1424);
nand U2754 (N_2754,In_839,In_799);
and U2755 (N_2755,In_427,In_908);
nand U2756 (N_2756,In_601,In_67);
nand U2757 (N_2757,In_380,In_435);
and U2758 (N_2758,In_1145,In_846);
or U2759 (N_2759,In_1256,In_629);
or U2760 (N_2760,In_1199,In_908);
or U2761 (N_2761,In_1264,In_586);
or U2762 (N_2762,In_246,In_570);
nand U2763 (N_2763,In_703,In_698);
and U2764 (N_2764,In_409,In_693);
or U2765 (N_2765,In_1000,In_1441);
and U2766 (N_2766,In_718,In_896);
nand U2767 (N_2767,In_944,In_897);
xnor U2768 (N_2768,In_1205,In_284);
nand U2769 (N_2769,In_1250,In_1496);
nand U2770 (N_2770,In_698,In_679);
xor U2771 (N_2771,In_854,In_184);
or U2772 (N_2772,In_105,In_1412);
nand U2773 (N_2773,In_608,In_823);
nor U2774 (N_2774,In_423,In_519);
or U2775 (N_2775,In_1395,In_915);
or U2776 (N_2776,In_438,In_426);
or U2777 (N_2777,In_218,In_1405);
and U2778 (N_2778,In_518,In_1496);
nand U2779 (N_2779,In_388,In_1053);
nor U2780 (N_2780,In_1091,In_317);
nor U2781 (N_2781,In_205,In_273);
xor U2782 (N_2782,In_767,In_1391);
nand U2783 (N_2783,In_300,In_1262);
nor U2784 (N_2784,In_1103,In_1397);
nand U2785 (N_2785,In_158,In_1495);
nand U2786 (N_2786,In_8,In_1411);
or U2787 (N_2787,In_603,In_282);
and U2788 (N_2788,In_1018,In_576);
nor U2789 (N_2789,In_898,In_729);
or U2790 (N_2790,In_502,In_334);
nand U2791 (N_2791,In_70,In_49);
nor U2792 (N_2792,In_570,In_319);
nor U2793 (N_2793,In_1332,In_1215);
or U2794 (N_2794,In_874,In_1455);
or U2795 (N_2795,In_617,In_1415);
or U2796 (N_2796,In_277,In_42);
nor U2797 (N_2797,In_24,In_252);
nor U2798 (N_2798,In_181,In_346);
nand U2799 (N_2799,In_240,In_86);
and U2800 (N_2800,In_684,In_297);
or U2801 (N_2801,In_1266,In_166);
nand U2802 (N_2802,In_1481,In_859);
nand U2803 (N_2803,In_1050,In_168);
and U2804 (N_2804,In_302,In_1314);
nor U2805 (N_2805,In_966,In_494);
nor U2806 (N_2806,In_975,In_1021);
or U2807 (N_2807,In_854,In_1277);
xnor U2808 (N_2808,In_1027,In_706);
or U2809 (N_2809,In_1069,In_1200);
and U2810 (N_2810,In_665,In_427);
or U2811 (N_2811,In_111,In_739);
and U2812 (N_2812,In_1321,In_51);
and U2813 (N_2813,In_404,In_666);
nor U2814 (N_2814,In_1051,In_782);
xor U2815 (N_2815,In_524,In_662);
nand U2816 (N_2816,In_1311,In_192);
nand U2817 (N_2817,In_3,In_557);
and U2818 (N_2818,In_59,In_1479);
nor U2819 (N_2819,In_600,In_982);
nor U2820 (N_2820,In_1350,In_678);
nand U2821 (N_2821,In_179,In_1479);
and U2822 (N_2822,In_343,In_254);
nand U2823 (N_2823,In_1321,In_716);
xor U2824 (N_2824,In_163,In_435);
nand U2825 (N_2825,In_1475,In_1378);
xor U2826 (N_2826,In_1265,In_647);
nor U2827 (N_2827,In_1107,In_1000);
nor U2828 (N_2828,In_489,In_266);
or U2829 (N_2829,In_453,In_1373);
and U2830 (N_2830,In_1001,In_1170);
or U2831 (N_2831,In_1379,In_259);
or U2832 (N_2832,In_1236,In_388);
nor U2833 (N_2833,In_937,In_382);
or U2834 (N_2834,In_1024,In_1116);
and U2835 (N_2835,In_1022,In_1491);
xnor U2836 (N_2836,In_918,In_374);
nand U2837 (N_2837,In_337,In_1413);
nand U2838 (N_2838,In_999,In_417);
or U2839 (N_2839,In_584,In_543);
nor U2840 (N_2840,In_168,In_489);
xnor U2841 (N_2841,In_598,In_574);
nand U2842 (N_2842,In_298,In_509);
or U2843 (N_2843,In_690,In_747);
and U2844 (N_2844,In_69,In_1431);
nand U2845 (N_2845,In_105,In_320);
or U2846 (N_2846,In_693,In_1338);
xnor U2847 (N_2847,In_312,In_445);
and U2848 (N_2848,In_379,In_810);
and U2849 (N_2849,In_420,In_1113);
or U2850 (N_2850,In_732,In_886);
and U2851 (N_2851,In_356,In_1252);
or U2852 (N_2852,In_624,In_1197);
and U2853 (N_2853,In_1277,In_1075);
nor U2854 (N_2854,In_802,In_1094);
nor U2855 (N_2855,In_134,In_442);
nand U2856 (N_2856,In_700,In_110);
or U2857 (N_2857,In_622,In_983);
and U2858 (N_2858,In_1051,In_420);
xor U2859 (N_2859,In_1456,In_514);
nand U2860 (N_2860,In_561,In_583);
and U2861 (N_2861,In_1123,In_1323);
and U2862 (N_2862,In_317,In_817);
nand U2863 (N_2863,In_1359,In_1209);
nor U2864 (N_2864,In_390,In_1159);
xnor U2865 (N_2865,In_1276,In_236);
nor U2866 (N_2866,In_1067,In_951);
and U2867 (N_2867,In_512,In_471);
or U2868 (N_2868,In_733,In_1128);
nor U2869 (N_2869,In_946,In_384);
nor U2870 (N_2870,In_1305,In_673);
nand U2871 (N_2871,In_1408,In_212);
xnor U2872 (N_2872,In_974,In_1354);
or U2873 (N_2873,In_662,In_837);
or U2874 (N_2874,In_1394,In_1195);
nor U2875 (N_2875,In_507,In_162);
or U2876 (N_2876,In_719,In_833);
and U2877 (N_2877,In_141,In_305);
and U2878 (N_2878,In_889,In_529);
xor U2879 (N_2879,In_718,In_1152);
and U2880 (N_2880,In_1081,In_81);
or U2881 (N_2881,In_889,In_1326);
nor U2882 (N_2882,In_1270,In_360);
or U2883 (N_2883,In_1443,In_1291);
nand U2884 (N_2884,In_213,In_484);
nor U2885 (N_2885,In_435,In_796);
nand U2886 (N_2886,In_1180,In_684);
nor U2887 (N_2887,In_227,In_1183);
or U2888 (N_2888,In_81,In_504);
nand U2889 (N_2889,In_379,In_444);
xor U2890 (N_2890,In_1024,In_1039);
nand U2891 (N_2891,In_1417,In_999);
or U2892 (N_2892,In_684,In_22);
nor U2893 (N_2893,In_726,In_81);
and U2894 (N_2894,In_365,In_194);
nand U2895 (N_2895,In_31,In_516);
or U2896 (N_2896,In_1413,In_906);
or U2897 (N_2897,In_477,In_944);
nand U2898 (N_2898,In_1341,In_681);
xnor U2899 (N_2899,In_921,In_374);
nor U2900 (N_2900,In_1286,In_169);
or U2901 (N_2901,In_434,In_154);
xor U2902 (N_2902,In_1014,In_911);
and U2903 (N_2903,In_309,In_398);
nor U2904 (N_2904,In_1084,In_497);
nor U2905 (N_2905,In_979,In_1441);
or U2906 (N_2906,In_905,In_1316);
or U2907 (N_2907,In_310,In_883);
nand U2908 (N_2908,In_388,In_95);
or U2909 (N_2909,In_1185,In_132);
or U2910 (N_2910,In_423,In_322);
and U2911 (N_2911,In_889,In_431);
and U2912 (N_2912,In_1305,In_947);
xnor U2913 (N_2913,In_731,In_1003);
nand U2914 (N_2914,In_463,In_245);
nor U2915 (N_2915,In_186,In_577);
nor U2916 (N_2916,In_1079,In_427);
or U2917 (N_2917,In_1054,In_499);
xnor U2918 (N_2918,In_77,In_107);
nor U2919 (N_2919,In_1489,In_1223);
and U2920 (N_2920,In_30,In_422);
or U2921 (N_2921,In_1318,In_864);
xor U2922 (N_2922,In_629,In_740);
and U2923 (N_2923,In_968,In_1382);
and U2924 (N_2924,In_1390,In_758);
nand U2925 (N_2925,In_618,In_827);
nor U2926 (N_2926,In_1023,In_208);
and U2927 (N_2927,In_1376,In_1344);
or U2928 (N_2928,In_1359,In_620);
nand U2929 (N_2929,In_1150,In_1496);
nor U2930 (N_2930,In_19,In_1122);
nand U2931 (N_2931,In_653,In_158);
and U2932 (N_2932,In_644,In_957);
nor U2933 (N_2933,In_754,In_277);
nor U2934 (N_2934,In_485,In_166);
xnor U2935 (N_2935,In_623,In_1438);
and U2936 (N_2936,In_237,In_1148);
and U2937 (N_2937,In_555,In_42);
nand U2938 (N_2938,In_698,In_1153);
or U2939 (N_2939,In_34,In_1);
nand U2940 (N_2940,In_393,In_1294);
and U2941 (N_2941,In_600,In_482);
or U2942 (N_2942,In_1317,In_1278);
or U2943 (N_2943,In_957,In_1123);
and U2944 (N_2944,In_970,In_754);
nand U2945 (N_2945,In_1128,In_693);
or U2946 (N_2946,In_612,In_1313);
nor U2947 (N_2947,In_815,In_868);
and U2948 (N_2948,In_536,In_224);
and U2949 (N_2949,In_1269,In_681);
nand U2950 (N_2950,In_11,In_803);
xor U2951 (N_2951,In_193,In_1273);
nor U2952 (N_2952,In_1432,In_762);
nor U2953 (N_2953,In_276,In_93);
nor U2954 (N_2954,In_323,In_827);
or U2955 (N_2955,In_73,In_358);
and U2956 (N_2956,In_1115,In_1281);
or U2957 (N_2957,In_334,In_596);
or U2958 (N_2958,In_1262,In_367);
nor U2959 (N_2959,In_1080,In_1063);
xnor U2960 (N_2960,In_348,In_1401);
and U2961 (N_2961,In_668,In_1293);
or U2962 (N_2962,In_1301,In_167);
or U2963 (N_2963,In_1394,In_1254);
nor U2964 (N_2964,In_1418,In_1256);
nor U2965 (N_2965,In_136,In_972);
nand U2966 (N_2966,In_1032,In_300);
nor U2967 (N_2967,In_901,In_347);
or U2968 (N_2968,In_791,In_726);
nor U2969 (N_2969,In_59,In_1208);
nand U2970 (N_2970,In_331,In_68);
nand U2971 (N_2971,In_951,In_978);
or U2972 (N_2972,In_835,In_1174);
nand U2973 (N_2973,In_426,In_362);
nand U2974 (N_2974,In_1164,In_1107);
nor U2975 (N_2975,In_280,In_249);
or U2976 (N_2976,In_357,In_40);
nor U2977 (N_2977,In_876,In_831);
xor U2978 (N_2978,In_697,In_98);
or U2979 (N_2979,In_270,In_60);
nor U2980 (N_2980,In_433,In_773);
or U2981 (N_2981,In_1026,In_1354);
nand U2982 (N_2982,In_50,In_965);
nand U2983 (N_2983,In_234,In_883);
nor U2984 (N_2984,In_394,In_105);
nand U2985 (N_2985,In_1230,In_1381);
nor U2986 (N_2986,In_98,In_852);
nand U2987 (N_2987,In_455,In_916);
nand U2988 (N_2988,In_130,In_61);
nor U2989 (N_2989,In_548,In_1329);
nand U2990 (N_2990,In_105,In_484);
nand U2991 (N_2991,In_1295,In_149);
and U2992 (N_2992,In_1084,In_212);
nand U2993 (N_2993,In_431,In_73);
or U2994 (N_2994,In_228,In_1017);
nor U2995 (N_2995,In_741,In_101);
xor U2996 (N_2996,In_861,In_506);
nand U2997 (N_2997,In_1381,In_1139);
or U2998 (N_2998,In_448,In_1119);
nor U2999 (N_2999,In_1130,In_867);
and U3000 (N_3000,N_1609,N_435);
nor U3001 (N_3001,N_1151,N_1107);
and U3002 (N_3002,N_2673,N_2722);
or U3003 (N_3003,N_1549,N_596);
or U3004 (N_3004,N_2190,N_1538);
nand U3005 (N_3005,N_1989,N_469);
and U3006 (N_3006,N_2697,N_1472);
and U3007 (N_3007,N_514,N_2321);
and U3008 (N_3008,N_350,N_2093);
and U3009 (N_3009,N_221,N_329);
and U3010 (N_3010,N_531,N_2913);
and U3011 (N_3011,N_1813,N_1500);
nor U3012 (N_3012,N_2266,N_1290);
nand U3013 (N_3013,N_1794,N_2268);
nor U3014 (N_3014,N_1228,N_2768);
or U3015 (N_3015,N_1351,N_838);
or U3016 (N_3016,N_2307,N_313);
and U3017 (N_3017,N_2134,N_1824);
nand U3018 (N_3018,N_374,N_780);
xor U3019 (N_3019,N_2685,N_1735);
and U3020 (N_3020,N_2483,N_163);
and U3021 (N_3021,N_819,N_252);
nor U3022 (N_3022,N_2285,N_226);
or U3023 (N_3023,N_671,N_2787);
or U3024 (N_3024,N_978,N_7);
and U3025 (N_3025,N_2569,N_2009);
and U3026 (N_3026,N_1900,N_2176);
or U3027 (N_3027,N_308,N_1099);
and U3028 (N_3028,N_88,N_1411);
xnor U3029 (N_3029,N_2156,N_1865);
and U3030 (N_3030,N_326,N_2962);
nor U3031 (N_3031,N_773,N_1035);
nand U3032 (N_3032,N_537,N_2919);
or U3033 (N_3033,N_2874,N_1977);
and U3034 (N_3034,N_1763,N_383);
nor U3035 (N_3035,N_1819,N_730);
xnor U3036 (N_3036,N_896,N_304);
nor U3037 (N_3037,N_2477,N_2090);
and U3038 (N_3038,N_2794,N_2803);
nand U3039 (N_3039,N_406,N_1384);
nand U3040 (N_3040,N_1670,N_2661);
nand U3041 (N_3041,N_344,N_867);
or U3042 (N_3042,N_607,N_684);
nand U3043 (N_3043,N_1967,N_1124);
or U3044 (N_3044,N_764,N_795);
nand U3045 (N_3045,N_1869,N_1523);
and U3046 (N_3046,N_2601,N_822);
and U3047 (N_3047,N_2409,N_915);
xor U3048 (N_3048,N_327,N_2716);
nor U3049 (N_3049,N_2884,N_11);
or U3050 (N_3050,N_1381,N_1329);
and U3051 (N_3051,N_999,N_1349);
nand U3052 (N_3052,N_2870,N_1374);
and U3053 (N_3053,N_1123,N_480);
xnor U3054 (N_3054,N_2905,N_2756);
and U3055 (N_3055,N_1898,N_488);
and U3056 (N_3056,N_2765,N_248);
and U3057 (N_3057,N_2588,N_376);
and U3058 (N_3058,N_934,N_1271);
nand U3059 (N_3059,N_2337,N_1651);
or U3060 (N_3060,N_891,N_301);
or U3061 (N_3061,N_2043,N_1076);
nand U3062 (N_3062,N_2796,N_1119);
or U3063 (N_3063,N_2968,N_1547);
and U3064 (N_3064,N_1449,N_1702);
or U3065 (N_3065,N_119,N_629);
nand U3066 (N_3066,N_260,N_2986);
or U3067 (N_3067,N_2762,N_1964);
nand U3068 (N_3068,N_1048,N_2993);
nor U3069 (N_3069,N_1542,N_1568);
nand U3070 (N_3070,N_2877,N_62);
and U3071 (N_3071,N_524,N_2378);
nor U3072 (N_3072,N_1879,N_1178);
nor U3073 (N_3073,N_2540,N_2581);
nor U3074 (N_3074,N_584,N_2853);
and U3075 (N_3075,N_649,N_1953);
or U3076 (N_3076,N_887,N_1682);
nand U3077 (N_3077,N_2000,N_2451);
nand U3078 (N_3078,N_2450,N_2008);
or U3079 (N_3079,N_1460,N_1180);
and U3080 (N_3080,N_2362,N_2245);
or U3081 (N_3081,N_2290,N_1826);
or U3082 (N_3082,N_1213,N_839);
nor U3083 (N_3083,N_1526,N_2772);
xnor U3084 (N_3084,N_1424,N_2433);
or U3085 (N_3085,N_844,N_1017);
and U3086 (N_3086,N_246,N_2767);
nand U3087 (N_3087,N_530,N_557);
and U3088 (N_3088,N_1278,N_983);
nor U3089 (N_3089,N_1173,N_2500);
xor U3090 (N_3090,N_2791,N_1969);
nand U3091 (N_3091,N_2092,N_2432);
nand U3092 (N_3092,N_2445,N_2388);
or U3093 (N_3093,N_755,N_402);
nor U3094 (N_3094,N_1172,N_526);
nand U3095 (N_3095,N_1970,N_2980);
or U3096 (N_3096,N_2827,N_13);
and U3097 (N_3097,N_1184,N_2749);
xor U3098 (N_3098,N_2658,N_2502);
or U3099 (N_3099,N_2162,N_1577);
nor U3100 (N_3100,N_2833,N_306);
and U3101 (N_3101,N_456,N_1186);
or U3102 (N_3102,N_620,N_728);
nor U3103 (N_3103,N_2955,N_2634);
or U3104 (N_3104,N_1498,N_1372);
or U3105 (N_3105,N_2194,N_141);
nor U3106 (N_3106,N_2954,N_2068);
and U3107 (N_3107,N_170,N_1612);
or U3108 (N_3108,N_2314,N_2900);
or U3109 (N_3109,N_388,N_1355);
or U3110 (N_3110,N_1164,N_1642);
xnor U3111 (N_3111,N_664,N_815);
or U3112 (N_3112,N_1646,N_2299);
nor U3113 (N_3113,N_338,N_630);
and U3114 (N_3114,N_2776,N_2503);
nor U3115 (N_3115,N_157,N_2505);
nor U3116 (N_3116,N_2754,N_1641);
nor U3117 (N_3117,N_1821,N_2088);
or U3118 (N_3118,N_840,N_552);
or U3119 (N_3119,N_1757,N_475);
or U3120 (N_3120,N_827,N_2029);
nand U3121 (N_3121,N_903,N_1730);
and U3122 (N_3122,N_1886,N_250);
nand U3123 (N_3123,N_1947,N_511);
nor U3124 (N_3124,N_2849,N_466);
nor U3125 (N_3125,N_1044,N_1979);
and U3126 (N_3126,N_359,N_1464);
nand U3127 (N_3127,N_1098,N_605);
or U3128 (N_3128,N_2950,N_53);
nor U3129 (N_3129,N_1331,N_2626);
nand U3130 (N_3130,N_333,N_953);
nand U3131 (N_3131,N_1811,N_2840);
nand U3132 (N_3132,N_577,N_1181);
nor U3133 (N_3133,N_386,N_225);
nor U3134 (N_3134,N_105,N_461);
nor U3135 (N_3135,N_2751,N_2340);
and U3136 (N_3136,N_416,N_2216);
xnor U3137 (N_3137,N_2017,N_2128);
nor U3138 (N_3138,N_984,N_1313);
nand U3139 (N_3139,N_472,N_1574);
nor U3140 (N_3140,N_124,N_2837);
nor U3141 (N_3141,N_1850,N_1761);
nor U3142 (N_3142,N_2535,N_2967);
and U3143 (N_3143,N_1956,N_2238);
and U3144 (N_3144,N_2724,N_880);
and U3145 (N_3145,N_1972,N_112);
nor U3146 (N_3146,N_2552,N_693);
nand U3147 (N_3147,N_2683,N_1981);
nor U3148 (N_3148,N_1852,N_1796);
or U3149 (N_3149,N_2616,N_1668);
and U3150 (N_3150,N_130,N_2107);
and U3151 (N_3151,N_1766,N_2899);
and U3152 (N_3152,N_291,N_1159);
or U3153 (N_3153,N_1634,N_2773);
and U3154 (N_3154,N_2995,N_1685);
nand U3155 (N_3155,N_2777,N_1418);
and U3156 (N_3156,N_1725,N_271);
or U3157 (N_3157,N_44,N_351);
nor U3158 (N_3158,N_169,N_2901);
or U3159 (N_3159,N_2060,N_1717);
and U3160 (N_3160,N_1769,N_973);
or U3161 (N_3161,N_847,N_733);
nand U3162 (N_3162,N_2147,N_1513);
nor U3163 (N_3163,N_192,N_1262);
nand U3164 (N_3164,N_1803,N_1308);
nor U3165 (N_3165,N_1104,N_1400);
or U3166 (N_3166,N_2880,N_851);
xor U3167 (N_3167,N_1416,N_2416);
xnor U3168 (N_3168,N_2202,N_2381);
nand U3169 (N_3169,N_1705,N_771);
and U3170 (N_3170,N_2100,N_143);
or U3171 (N_3171,N_2769,N_161);
xor U3172 (N_3172,N_1169,N_1784);
nand U3173 (N_3173,N_1556,N_240);
nor U3174 (N_3174,N_2452,N_2318);
nand U3175 (N_3175,N_750,N_614);
nor U3176 (N_3176,N_2077,N_1320);
nand U3177 (N_3177,N_2851,N_2753);
nor U3178 (N_3178,N_1322,N_2983);
nand U3179 (N_3179,N_1710,N_280);
or U3180 (N_3180,N_2517,N_2462);
or U3181 (N_3181,N_1842,N_970);
nor U3182 (N_3182,N_486,N_251);
or U3183 (N_3183,N_1663,N_1254);
nor U3184 (N_3184,N_2620,N_1699);
xnor U3185 (N_3185,N_2225,N_2957);
or U3186 (N_3186,N_126,N_1368);
nand U3187 (N_3187,N_167,N_566);
nand U3188 (N_3188,N_615,N_591);
or U3189 (N_3189,N_2869,N_946);
and U3190 (N_3190,N_423,N_61);
and U3191 (N_3191,N_2960,N_942);
nand U3192 (N_3192,N_2752,N_1031);
or U3193 (N_3193,N_2028,N_397);
or U3194 (N_3194,N_238,N_289);
and U3195 (N_3195,N_2389,N_2138);
nand U3196 (N_3196,N_2089,N_1108);
or U3197 (N_3197,N_535,N_2165);
or U3198 (N_3198,N_1752,N_110);
nand U3199 (N_3199,N_2132,N_1480);
nor U3200 (N_3200,N_1442,N_2873);
nand U3201 (N_3201,N_1974,N_463);
nand U3202 (N_3202,N_465,N_2774);
nand U3203 (N_3203,N_1350,N_180);
xnor U3204 (N_3204,N_917,N_1288);
nand U3205 (N_3205,N_2526,N_2660);
nand U3206 (N_3206,N_2990,N_1863);
xor U3207 (N_3207,N_1873,N_66);
and U3208 (N_3208,N_742,N_231);
and U3209 (N_3209,N_1045,N_2484);
nor U3210 (N_3210,N_1890,N_1265);
or U3211 (N_3211,N_1903,N_2338);
and U3212 (N_3212,N_1335,N_705);
or U3213 (N_3213,N_749,N_2615);
and U3214 (N_3214,N_1330,N_1176);
nor U3215 (N_3215,N_718,N_1287);
nand U3216 (N_3216,N_2631,N_27);
nand U3217 (N_3217,N_1062,N_223);
and U3218 (N_3218,N_1716,N_1370);
nand U3219 (N_3219,N_0,N_2254);
or U3220 (N_3220,N_608,N_547);
and U3221 (N_3221,N_434,N_2710);
nor U3222 (N_3222,N_1633,N_85);
or U3223 (N_3223,N_299,N_2487);
and U3224 (N_3224,N_644,N_1469);
nand U3225 (N_3225,N_1025,N_2065);
and U3226 (N_3226,N_1445,N_735);
and U3227 (N_3227,N_2675,N_94);
and U3228 (N_3228,N_1301,N_2013);
or U3229 (N_3229,N_310,N_2326);
nor U3230 (N_3230,N_366,N_1519);
or U3231 (N_3231,N_462,N_1948);
nor U3232 (N_3232,N_2953,N_1489);
or U3233 (N_3233,N_636,N_1130);
or U3234 (N_3234,N_297,N_508);
or U3235 (N_3235,N_1626,N_2582);
nor U3236 (N_3236,N_334,N_2044);
or U3237 (N_3237,N_1314,N_2053);
nor U3238 (N_3238,N_2702,N_1874);
and U3239 (N_3239,N_1249,N_325);
or U3240 (N_3240,N_660,N_854);
nand U3241 (N_3241,N_2779,N_2363);
nor U3242 (N_3242,N_2372,N_1615);
and U3243 (N_3243,N_943,N_30);
nand U3244 (N_3244,N_2654,N_135);
nand U3245 (N_3245,N_2403,N_1667);
xor U3246 (N_3246,N_89,N_675);
xnor U3247 (N_3247,N_950,N_710);
and U3248 (N_3248,N_2510,N_1334);
or U3249 (N_3249,N_1153,N_2126);
and U3250 (N_3250,N_2666,N_2830);
nand U3251 (N_3251,N_2521,N_2206);
nor U3252 (N_3252,N_2463,N_72);
nand U3253 (N_3253,N_2408,N_1866);
or U3254 (N_3254,N_74,N_1448);
nand U3255 (N_3255,N_2259,N_2533);
and U3256 (N_3256,N_1860,N_1738);
nand U3257 (N_3257,N_1917,N_2831);
and U3258 (N_3258,N_1244,N_335);
xor U3259 (N_3259,N_2942,N_2230);
or U3260 (N_3260,N_1291,N_1027);
nor U3261 (N_3261,N_1503,N_1407);
and U3262 (N_3262,N_2708,N_2458);
and U3263 (N_3263,N_1120,N_1918);
nand U3264 (N_3264,N_1736,N_1441);
nor U3265 (N_3265,N_2972,N_2229);
or U3266 (N_3266,N_268,N_1430);
or U3267 (N_3267,N_479,N_2410);
nor U3268 (N_3268,N_2113,N_269);
xor U3269 (N_3269,N_1586,N_505);
nand U3270 (N_3270,N_2010,N_1317);
and U3271 (N_3271,N_2367,N_952);
or U3272 (N_3272,N_1200,N_497);
and U3273 (N_3273,N_1148,N_1812);
or U3274 (N_3274,N_162,N_1516);
nand U3275 (N_3275,N_974,N_2041);
nand U3276 (N_3276,N_1101,N_1353);
nor U3277 (N_3277,N_1601,N_2427);
and U3278 (N_3278,N_1457,N_2319);
or U3279 (N_3279,N_1872,N_1459);
nor U3280 (N_3280,N_1206,N_1100);
nand U3281 (N_3281,N_1895,N_1427);
or U3282 (N_3282,N_2214,N_2878);
and U3283 (N_3283,N_1305,N_2342);
and U3284 (N_3284,N_230,N_1052);
xnor U3285 (N_3285,N_1655,N_426);
and U3286 (N_3286,N_1715,N_2261);
nand U3287 (N_3287,N_2886,N_2574);
or U3288 (N_3288,N_75,N_1337);
or U3289 (N_3289,N_1083,N_154);
nand U3290 (N_3290,N_808,N_1389);
or U3291 (N_3291,N_885,N_1671);
xnor U3292 (N_3292,N_139,N_133);
nand U3293 (N_3293,N_2102,N_570);
xnor U3294 (N_3294,N_2212,N_2829);
and U3295 (N_3295,N_302,N_1491);
nand U3296 (N_3296,N_681,N_1079);
xnor U3297 (N_3297,N_290,N_1767);
xnor U3298 (N_3298,N_1401,N_2048);
and U3299 (N_3299,N_147,N_1396);
nand U3300 (N_3300,N_929,N_2580);
and U3301 (N_3301,N_2490,N_2527);
nor U3302 (N_3302,N_1701,N_1289);
nand U3303 (N_3303,N_1438,N_1406);
and U3304 (N_3304,N_2932,N_1672);
nand U3305 (N_3305,N_1229,N_2543);
or U3306 (N_3306,N_588,N_179);
and U3307 (N_3307,N_1256,N_56);
or U3308 (N_3308,N_1889,N_2124);
or U3309 (N_3309,N_1201,N_2965);
nor U3310 (N_3310,N_540,N_1906);
or U3311 (N_3311,N_708,N_2744);
xor U3312 (N_3312,N_35,N_29);
nand U3313 (N_3313,N_2439,N_2975);
nor U3314 (N_3314,N_1167,N_320);
nor U3315 (N_3315,N_853,N_825);
or U3316 (N_3316,N_2051,N_2584);
nand U3317 (N_3317,N_2241,N_204);
nor U3318 (N_3318,N_2365,N_648);
or U3319 (N_3319,N_2903,N_1203);
or U3320 (N_3320,N_1829,N_2320);
and U3321 (N_3321,N_2867,N_1046);
or U3322 (N_3322,N_275,N_2233);
or U3323 (N_3323,N_600,N_2413);
nor U3324 (N_3324,N_1771,N_477);
and U3325 (N_3325,N_1481,N_1770);
nand U3326 (N_3326,N_28,N_2308);
nor U3327 (N_3327,N_372,N_496);
or U3328 (N_3328,N_2536,N_1094);
and U3329 (N_3329,N_2676,N_1611);
nand U3330 (N_3330,N_2024,N_975);
xnor U3331 (N_3331,N_2080,N_429);
and U3332 (N_3332,N_1490,N_83);
nor U3333 (N_3333,N_243,N_2862);
and U3334 (N_3334,N_1792,N_1728);
or U3335 (N_3335,N_525,N_2264);
or U3336 (N_3336,N_1983,N_2551);
nor U3337 (N_3337,N_1199,N_1437);
xnor U3338 (N_3338,N_993,N_1085);
or U3339 (N_3339,N_2313,N_2558);
or U3340 (N_3340,N_2579,N_1482);
and U3341 (N_3341,N_2600,N_912);
and U3342 (N_3342,N_2511,N_1117);
nand U3343 (N_3343,N_1224,N_609);
nor U3344 (N_3344,N_1485,N_713);
or U3345 (N_3345,N_2087,N_210);
or U3346 (N_3346,N_1864,N_1570);
and U3347 (N_3347,N_997,N_2461);
nor U3348 (N_3348,N_2366,N_2197);
and U3349 (N_3349,N_964,N_2406);
nand U3350 (N_3350,N_726,N_990);
nand U3351 (N_3351,N_54,N_185);
nor U3352 (N_3352,N_2509,N_57);
xnor U3353 (N_3353,N_449,N_1319);
or U3354 (N_3354,N_2783,N_1986);
xor U3355 (N_3355,N_2652,N_581);
and U3356 (N_3356,N_1261,N_128);
and U3357 (N_3357,N_940,N_1116);
nor U3358 (N_3358,N_836,N_1569);
nor U3359 (N_3359,N_2547,N_1300);
and U3360 (N_3360,N_1049,N_120);
or U3361 (N_3361,N_559,N_2653);
nor U3362 (N_3362,N_2262,N_1799);
nor U3363 (N_3363,N_1060,N_1476);
nor U3364 (N_3364,N_611,N_2707);
nor U3365 (N_3365,N_818,N_968);
nor U3366 (N_3366,N_910,N_2935);
or U3367 (N_3367,N_1992,N_2723);
and U3368 (N_3368,N_2917,N_1923);
or U3369 (N_3369,N_981,N_2154);
nor U3370 (N_3370,N_2619,N_2192);
or U3371 (N_3371,N_639,N_645);
nand U3372 (N_3372,N_923,N_937);
nand U3373 (N_3373,N_663,N_2042);
and U3374 (N_3374,N_1077,N_1961);
nor U3375 (N_3375,N_2944,N_417);
nor U3376 (N_3376,N_1061,N_2136);
nand U3377 (N_3377,N_2207,N_1158);
nor U3378 (N_3378,N_216,N_1346);
nand U3379 (N_3379,N_1662,N_2160);
and U3380 (N_3380,N_474,N_2066);
nand U3381 (N_3381,N_2014,N_258);
nand U3382 (N_3382,N_1748,N_2866);
xnor U3383 (N_3383,N_403,N_1383);
nand U3384 (N_3384,N_1036,N_321);
nand U3385 (N_3385,N_1598,N_1576);
or U3386 (N_3386,N_895,N_916);
xnor U3387 (N_3387,N_876,N_274);
or U3388 (N_3388,N_834,N_1470);
nand U3389 (N_3389,N_1940,N_947);
and U3390 (N_3390,N_843,N_2603);
xor U3391 (N_3391,N_2145,N_471);
nor U3392 (N_3392,N_342,N_2795);
nor U3393 (N_3393,N_2692,N_1388);
and U3394 (N_3394,N_2115,N_6);
nand U3395 (N_3395,N_602,N_1128);
or U3396 (N_3396,N_2164,N_2798);
or U3397 (N_3397,N_1660,N_2453);
and U3398 (N_3398,N_267,N_1461);
nand U3399 (N_3399,N_1694,N_2758);
and U3400 (N_3400,N_2098,N_622);
and U3401 (N_3401,N_988,N_115);
or U3402 (N_3402,N_1674,N_2076);
nand U3403 (N_3403,N_1902,N_652);
or U3404 (N_3404,N_431,N_2251);
or U3405 (N_3405,N_1250,N_300);
and U3406 (N_3406,N_2385,N_509);
nand U3407 (N_3407,N_1434,N_2397);
nor U3408 (N_3408,N_899,N_193);
xnor U3409 (N_3409,N_786,N_1585);
and U3410 (N_3410,N_2546,N_814);
nand U3411 (N_3411,N_2741,N_1087);
nand U3412 (N_3412,N_1654,N_279);
or U3413 (N_3413,N_1357,N_613);
or U3414 (N_3414,N_1629,N_2889);
nor U3415 (N_3415,N_1645,N_1058);
xnor U3416 (N_3416,N_911,N_945);
nand U3417 (N_3417,N_58,N_1971);
nand U3418 (N_3418,N_1285,N_1772);
or U3419 (N_3419,N_2,N_2725);
xor U3420 (N_3420,N_2875,N_2393);
nand U3421 (N_3421,N_938,N_585);
nand U3422 (N_3422,N_2971,N_1935);
nor U3423 (N_3423,N_176,N_2181);
nor U3424 (N_3424,N_2236,N_965);
nand U3425 (N_3425,N_1666,N_2784);
xnor U3426 (N_3426,N_580,N_1592);
nor U3427 (N_3427,N_2936,N_504);
nor U3428 (N_3428,N_2717,N_1073);
nor U3429 (N_3429,N_2655,N_716);
xor U3430 (N_3430,N_1754,N_2428);
nand U3431 (N_3431,N_2857,N_194);
and U3432 (N_3432,N_2470,N_2946);
nand U3433 (N_3433,N_941,N_720);
or U3434 (N_3434,N_1571,N_2438);
and U3435 (N_3435,N_1911,N_2742);
or U3436 (N_3436,N_1550,N_1403);
nor U3437 (N_3437,N_1871,N_17);
or U3438 (N_3438,N_2221,N_2222);
nand U3439 (N_3439,N_2444,N_1659);
nor U3440 (N_3440,N_2291,N_761);
nor U3441 (N_3441,N_217,N_1032);
nor U3442 (N_3442,N_458,N_2846);
nand U3443 (N_3443,N_2992,N_1390);
and U3444 (N_3444,N_2498,N_548);
or U3445 (N_3445,N_2820,N_341);
nand U3446 (N_3446,N_659,N_2185);
and U3447 (N_3447,N_2914,N_2419);
nand U3448 (N_3448,N_2549,N_319);
nand U3449 (N_3449,N_685,N_883);
nand U3450 (N_3450,N_331,N_1764);
nor U3451 (N_3451,N_1950,N_758);
nand U3452 (N_3452,N_273,N_1194);
or U3453 (N_3453,N_751,N_2390);
and U3454 (N_3454,N_2376,N_1541);
or U3455 (N_3455,N_420,N_2638);
or U3456 (N_3456,N_1653,N_2057);
nand U3457 (N_3457,N_2883,N_184);
and U3458 (N_3458,N_318,N_1183);
nor U3459 (N_3459,N_1277,N_906);
and U3460 (N_3460,N_1591,N_2283);
and U3461 (N_3461,N_2231,N_2246);
nor U3462 (N_3462,N_1606,N_1259);
nand U3463 (N_3463,N_856,N_2641);
and U3464 (N_3464,N_1880,N_2679);
and U3465 (N_3465,N_1299,N_122);
nor U3466 (N_3466,N_935,N_2276);
xnor U3467 (N_3467,N_1931,N_1580);
and U3468 (N_3468,N_1417,N_1925);
or U3469 (N_3469,N_2850,N_424);
nand U3470 (N_3470,N_2471,N_1643);
nor U3471 (N_3471,N_489,N_400);
nand U3472 (N_3472,N_1878,N_2407);
nor U3473 (N_3473,N_2730,N_1024);
and U3474 (N_3474,N_1209,N_1775);
or U3475 (N_3475,N_2071,N_365);
nand U3476 (N_3476,N_1281,N_200);
and U3477 (N_3477,N_2607,N_740);
or U3478 (N_3478,N_1946,N_1790);
or U3479 (N_3479,N_202,N_1110);
and U3480 (N_3480,N_81,N_1729);
xor U3481 (N_3481,N_1144,N_218);
and U3482 (N_3482,N_1292,N_1905);
or U3483 (N_3483,N_985,N_2865);
nor U3484 (N_3484,N_1360,N_709);
xor U3485 (N_3485,N_2361,N_2354);
xnor U3486 (N_3486,N_2485,N_1637);
or U3487 (N_3487,N_1487,N_2374);
nand U3488 (N_3488,N_2688,N_1078);
or U3489 (N_3489,N_2636,N_1376);
nand U3490 (N_3490,N_3,N_2260);
xor U3491 (N_3491,N_1356,N_1837);
nand U3492 (N_3492,N_2548,N_2091);
or U3493 (N_3493,N_385,N_206);
and U3494 (N_3494,N_1326,N_2150);
nand U3495 (N_3495,N_1001,N_2034);
nand U3496 (N_3496,N_987,N_413);
or U3497 (N_3497,N_545,N_1325);
nand U3498 (N_3498,N_2994,N_1091);
nor U3499 (N_3499,N_2210,N_2278);
or U3500 (N_3500,N_2520,N_837);
and U3501 (N_3501,N_977,N_2910);
nor U3502 (N_3502,N_1162,N_476);
or U3503 (N_3503,N_1720,N_634);
or U3504 (N_3504,N_2882,N_1707);
nor U3505 (N_3505,N_1304,N_1926);
xor U3506 (N_3506,N_2933,N_2027);
nand U3507 (N_3507,N_2728,N_731);
or U3508 (N_3508,N_2064,N_389);
and U3509 (N_3509,N_2988,N_2970);
nor U3510 (N_3510,N_1409,N_1088);
xor U3511 (N_3511,N_2847,N_2764);
nor U3512 (N_3512,N_1963,N_2622);
nor U3513 (N_3513,N_2384,N_1594);
xor U3514 (N_3514,N_918,N_1019);
nor U3515 (N_3515,N_1251,N_263);
nor U3516 (N_3516,N_1207,N_991);
nand U3517 (N_3517,N_440,N_2755);
nor U3518 (N_3518,N_732,N_1944);
and U3519 (N_3519,N_1005,N_872);
and U3520 (N_3520,N_286,N_1582);
and U3521 (N_3521,N_2550,N_2211);
or U3522 (N_3522,N_2242,N_597);
nand U3523 (N_3523,N_2140,N_205);
xnor U3524 (N_3524,N_2854,N_483);
nor U3525 (N_3525,N_2345,N_901);
nand U3526 (N_3526,N_2525,N_2371);
or U3527 (N_3527,N_2943,N_2825);
or U3528 (N_3528,N_2659,N_1597);
xor U3529 (N_3529,N_1844,N_168);
and U3530 (N_3530,N_1136,N_443);
and U3531 (N_3531,N_396,N_513);
and U3532 (N_3532,N_1613,N_2311);
or U3533 (N_3533,N_752,N_2003);
and U3534 (N_3534,N_610,N_797);
nand U3535 (N_3535,N_1377,N_1068);
or U3536 (N_3536,N_1632,N_1815);
nand U3537 (N_3537,N_765,N_1810);
xor U3538 (N_3538,N_414,N_2171);
or U3539 (N_3539,N_2949,N_1765);
and U3540 (N_3540,N_242,N_2049);
or U3541 (N_3541,N_2610,N_1678);
nor U3542 (N_3542,N_1071,N_1912);
and U3543 (N_3543,N_2443,N_712);
or U3544 (N_3544,N_1836,N_2208);
nor U3545 (N_3545,N_1584,N_812);
and U3546 (N_3546,N_1354,N_1191);
and U3547 (N_3547,N_2838,N_1901);
nor U3548 (N_3548,N_1524,N_1808);
and U3549 (N_3549,N_971,N_672);
or U3550 (N_3550,N_2868,N_2951);
nor U3551 (N_3551,N_1298,N_779);
and U3552 (N_3552,N_1945,N_485);
nor U3553 (N_3553,N_1283,N_361);
or U3554 (N_3554,N_1341,N_1090);
and U3555 (N_3555,N_1846,N_1089);
nand U3556 (N_3556,N_1006,N_188);
or U3557 (N_3557,N_2894,N_961);
xor U3558 (N_3558,N_1092,N_278);
nand U3559 (N_3559,N_2672,N_723);
nand U3560 (N_3560,N_2821,N_703);
and U3561 (N_3561,N_2357,N_1822);
and U3562 (N_3562,N_2052,N_1868);
nand U3563 (N_3563,N_2200,N_2189);
and U3564 (N_3564,N_879,N_1976);
xor U3565 (N_3565,N_2948,N_2814);
and U3566 (N_3566,N_520,N_2059);
nor U3567 (N_3567,N_2824,N_276);
nand U3568 (N_3568,N_1973,N_1908);
nor U3569 (N_3569,N_347,N_798);
xor U3570 (N_3570,N_1002,N_41);
nand U3571 (N_3571,N_775,N_567);
nor U3572 (N_3572,N_2130,N_2323);
nor U3573 (N_3573,N_909,N_2184);
nand U3574 (N_3574,N_1665,N_2306);
nor U3575 (N_3575,N_2789,N_650);
nor U3576 (N_3576,N_2495,N_387);
and U3577 (N_3577,N_2476,N_1378);
nand U3578 (N_3578,N_1129,N_1332);
nand U3579 (N_3579,N_237,N_482);
or U3580 (N_3580,N_2645,N_1567);
nor U3581 (N_3581,N_2544,N_2627);
nor U3582 (N_3582,N_2478,N_2835);
and U3583 (N_3583,N_2203,N_2213);
and U3584 (N_3584,N_2559,N_2508);
nand U3585 (N_3585,N_1056,N_1952);
nor U3586 (N_3586,N_1463,N_1382);
or U3587 (N_3587,N_239,N_2360);
nor U3588 (N_3588,N_228,N_2274);
and U3589 (N_3589,N_1897,N_9);
nand U3590 (N_3590,N_857,N_1233);
or U3591 (N_3591,N_2974,N_2651);
or U3592 (N_3592,N_1504,N_875);
xor U3593 (N_3593,N_2173,N_1276);
and U3594 (N_3594,N_939,N_2999);
or U3595 (N_3595,N_1057,N_2328);
nor U3596 (N_3596,N_1252,N_2127);
and U3597 (N_3597,N_802,N_24);
and U3598 (N_3598,N_2670,N_2897);
xor U3599 (N_3599,N_1861,N_433);
nand U3600 (N_3600,N_398,N_1140);
and U3601 (N_3601,N_2033,N_287);
nor U3602 (N_3602,N_224,N_930);
or U3603 (N_3603,N_667,N_2497);
and U3604 (N_3604,N_59,N_2583);
nand U3605 (N_3605,N_1333,N_2105);
or U3606 (N_3606,N_353,N_1525);
and U3607 (N_3607,N_117,N_826);
xnor U3608 (N_3608,N_255,N_2015);
nand U3609 (N_3609,N_957,N_2761);
nor U3610 (N_3610,N_1474,N_763);
and U3611 (N_3611,N_145,N_1497);
nand U3612 (N_3612,N_852,N_1559);
xor U3613 (N_3613,N_235,N_295);
xnor U3614 (N_3614,N_266,N_1640);
or U3615 (N_3615,N_776,N_467);
or U3616 (N_3616,N_93,N_78);
or U3617 (N_3617,N_858,N_2668);
xor U3618 (N_3618,N_2896,N_2472);
nand U3619 (N_3619,N_384,N_1236);
and U3620 (N_3620,N_1853,N_572);
or U3621 (N_3621,N_1323,N_156);
or U3622 (N_3622,N_860,N_91);
or U3623 (N_3623,N_236,N_2604);
or U3624 (N_3624,N_1521,N_2907);
nand U3625 (N_3625,N_1084,N_788);
and U3626 (N_3626,N_980,N_2398);
nor U3627 (N_3627,N_696,N_654);
nor U3628 (N_3628,N_108,N_2247);
nand U3629 (N_3629,N_1949,N_1834);
nor U3630 (N_3630,N_2488,N_2158);
and U3631 (N_3631,N_79,N_354);
and U3632 (N_3632,N_1820,N_2038);
or U3633 (N_3633,N_1700,N_624);
nand U3634 (N_3634,N_2125,N_1157);
or U3635 (N_3635,N_1444,N_828);
and U3636 (N_3636,N_691,N_2330);
nand U3637 (N_3637,N_1788,N_1484);
xnor U3638 (N_3638,N_1398,N_972);
nor U3639 (N_3639,N_803,N_2386);
nor U3640 (N_3640,N_2843,N_2909);
or U3641 (N_3641,N_1913,N_2177);
xor U3642 (N_3642,N_2733,N_1698);
nand U3643 (N_3643,N_1888,N_97);
nand U3644 (N_3644,N_2632,N_1561);
nand U3645 (N_3645,N_2499,N_2350);
or U3646 (N_3646,N_2782,N_447);
nor U3647 (N_3647,N_913,N_2074);
or U3648 (N_3648,N_43,N_2423);
nand U3649 (N_3649,N_2396,N_515);
or U3650 (N_3650,N_183,N_339);
or U3651 (N_3651,N_551,N_982);
or U3652 (N_3652,N_665,N_1737);
nor U3653 (N_3653,N_544,N_1146);
nor U3654 (N_3654,N_2287,N_594);
or U3655 (N_3655,N_1358,N_850);
and U3656 (N_3656,N_2081,N_2507);
and U3657 (N_3657,N_2842,N_1938);
and U3658 (N_3658,N_503,N_2709);
nand U3659 (N_3659,N_1741,N_2947);
xnor U3660 (N_3660,N_2465,N_2863);
nor U3661 (N_3661,N_357,N_2845);
and U3662 (N_3662,N_499,N_1065);
xnor U3663 (N_3663,N_1638,N_2669);
or U3664 (N_3664,N_2586,N_1450);
or U3665 (N_3665,N_2922,N_2613);
xor U3666 (N_3666,N_2792,N_2421);
nor U3667 (N_3667,N_2475,N_358);
and U3668 (N_3668,N_894,N_1630);
or U3669 (N_3669,N_2958,N_1026);
nor U3670 (N_3670,N_811,N_2186);
nor U3671 (N_3671,N_1978,N_1165);
or U3672 (N_3672,N_2713,N_823);
xnor U3673 (N_3673,N_285,N_1221);
nor U3674 (N_3674,N_2991,N_1473);
xor U3675 (N_3675,N_2491,N_109);
and U3676 (N_3676,N_1023,N_446);
nand U3677 (N_3677,N_647,N_689);
and U3678 (N_3678,N_2305,N_2567);
nor U3679 (N_3679,N_178,N_897);
and U3680 (N_3680,N_1137,N_65);
nor U3681 (N_3681,N_2832,N_2353);
or U3682 (N_3682,N_2111,N_704);
nor U3683 (N_3683,N_2152,N_2680);
or U3684 (N_3684,N_152,N_360);
nand U3685 (N_3685,N_741,N_2888);
and U3686 (N_3686,N_956,N_2629);
nand U3687 (N_3687,N_960,N_1627);
and U3688 (N_3688,N_1689,N_1067);
xor U3689 (N_3689,N_612,N_2025);
or U3690 (N_3690,N_2885,N_534);
or U3691 (N_3691,N_1778,N_2179);
xor U3692 (N_3692,N_19,N_2431);
nor U3693 (N_3693,N_2468,N_2539);
or U3694 (N_3694,N_47,N_1578);
xor U3695 (N_3695,N_2123,N_963);
or U3696 (N_3696,N_2045,N_2524);
and U3697 (N_3697,N_71,N_1081);
nand U3698 (N_3698,N_1614,N_270);
nand U3699 (N_3699,N_1939,N_1515);
nor U3700 (N_3700,N_766,N_1804);
nor U3701 (N_3701,N_322,N_2235);
nand U3702 (N_3702,N_679,N_1534);
or U3703 (N_3703,N_2435,N_1875);
xor U3704 (N_3704,N_2117,N_491);
and U3705 (N_3705,N_1691,N_1608);
nand U3706 (N_3706,N_1652,N_1588);
nand U3707 (N_3707,N_996,N_1697);
and U3708 (N_3708,N_405,N_1505);
or U3709 (N_3709,N_454,N_2978);
nor U3710 (N_3710,N_662,N_2589);
and U3711 (N_3711,N_2454,N_2678);
xnor U3712 (N_3712,N_2879,N_2858);
xnor U3713 (N_3713,N_101,N_1514);
nand U3714 (N_3714,N_2016,N_1798);
nor U3715 (N_3715,N_307,N_2402);
xor U3716 (N_3716,N_1554,N_1152);
nand U3717 (N_3717,N_919,N_2019);
nand U3718 (N_3718,N_2104,N_234);
nor U3719 (N_3719,N_1628,N_770);
nand U3720 (N_3720,N_2743,N_1639);
or U3721 (N_3721,N_478,N_1839);
nand U3722 (N_3722,N_1041,N_2848);
nor U3723 (N_3723,N_32,N_1795);
nand U3724 (N_3724,N_589,N_2802);
or U3725 (N_3725,N_617,N_1877);
and U3726 (N_3726,N_2599,N_259);
and U3727 (N_3727,N_2001,N_492);
nor U3728 (N_3728,N_208,N_1711);
xor U3729 (N_3729,N_64,N_1566);
or U3730 (N_3730,N_428,N_2963);
nand U3731 (N_3731,N_1096,N_2577);
nand U3732 (N_3732,N_1532,N_1127);
and U3733 (N_3733,N_2252,N_998);
and U3734 (N_3734,N_1011,N_442);
nand U3735 (N_3735,N_1,N_419);
or U3736 (N_3736,N_1817,N_1132);
nor U3737 (N_3737,N_2931,N_1142);
nand U3738 (N_3738,N_2534,N_2542);
and U3739 (N_3739,N_2934,N_1602);
nand U3740 (N_3740,N_2249,N_2997);
nor U3741 (N_3741,N_2082,N_1222);
and U3742 (N_3742,N_1205,N_2480);
and U3743 (N_3743,N_2030,N_2801);
nand U3744 (N_3744,N_719,N_1712);
and U3745 (N_3745,N_717,N_1193);
nor U3746 (N_3746,N_1404,N_121);
nor U3747 (N_3747,N_2187,N_2217);
nor U3748 (N_3748,N_1243,N_2817);
or U3749 (N_3749,N_835,N_2703);
or U3750 (N_3750,N_682,N_2637);
and U3751 (N_3751,N_2141,N_2139);
or U3752 (N_3752,N_1264,N_2172);
nand U3753 (N_3753,N_2530,N_1366);
nand U3754 (N_3754,N_1053,N_2295);
nand U3755 (N_3755,N_688,N_1451);
or U3756 (N_3756,N_2568,N_1230);
or U3757 (N_3757,N_1275,N_1018);
xor U3758 (N_3758,N_1217,N_1150);
and U3759 (N_3759,N_1246,N_1013);
and U3760 (N_3760,N_925,N_1517);
or U3761 (N_3761,N_288,N_1212);
nor U3762 (N_3762,N_190,N_2518);
nand U3763 (N_3763,N_1227,N_2504);
nand U3764 (N_3764,N_2859,N_1361);
or U3765 (N_3765,N_409,N_2623);
nor U3766 (N_3766,N_363,N_951);
nor U3767 (N_3767,N_2872,N_2344);
nor U3768 (N_3768,N_2572,N_1675);
or U3769 (N_3769,N_1467,N_2704);
nand U3770 (N_3770,N_1835,N_1155);
nand U3771 (N_3771,N_175,N_1744);
nor U3772 (N_3772,N_2731,N_1258);
xnor U3773 (N_3773,N_2852,N_959);
and U3774 (N_3774,N_783,N_1362);
nand U3775 (N_3775,N_1951,N_1783);
nor U3776 (N_3776,N_2425,N_1531);
xnor U3777 (N_3777,N_144,N_2770);
or U3778 (N_3778,N_1980,N_2694);
and U3779 (N_3779,N_1270,N_2188);
nand U3780 (N_3780,N_1443,N_2078);
xor U3781 (N_3781,N_1395,N_638);
or U3782 (N_3782,N_1174,N_1870);
or U3783 (N_3783,N_1619,N_592);
nand U3784 (N_3784,N_2144,N_2775);
nand U3785 (N_3785,N_1843,N_2004);
and U3786 (N_3786,N_1219,N_1296);
nand U3787 (N_3787,N_1693,N_1789);
nor U3788 (N_3788,N_2516,N_2807);
and U3789 (N_3789,N_2496,N_2771);
nor U3790 (N_3790,N_2952,N_1904);
and U3791 (N_3791,N_517,N_921);
or U3792 (N_3792,N_1241,N_2911);
and U3793 (N_3793,N_305,N_2804);
or U3794 (N_3794,N_969,N_468);
xnor U3795 (N_3795,N_16,N_1527);
nor U3796 (N_3796,N_127,N_1610);
nor U3797 (N_3797,N_2964,N_1631);
or U3798 (N_3798,N_2812,N_738);
and U3799 (N_3799,N_1138,N_800);
and U3800 (N_3800,N_1625,N_692);
nand U3801 (N_3801,N_315,N_1232);
nand U3802 (N_3802,N_283,N_2279);
and U3803 (N_3803,N_484,N_14);
and U3804 (N_3804,N_292,N_23);
or U3805 (N_3805,N_229,N_725);
or U3806 (N_3806,N_76,N_1985);
or U3807 (N_3807,N_2738,N_1273);
nand U3808 (N_3808,N_1664,N_1581);
or U3809 (N_3809,N_2561,N_1235);
and U3810 (N_3810,N_632,N_2640);
nand U3811 (N_3811,N_1805,N_2284);
and U3812 (N_3812,N_1551,N_317);
or U3813 (N_3813,N_787,N_1858);
and U3814 (N_3814,N_2294,N_38);
or U3815 (N_3815,N_1455,N_2712);
and U3816 (N_3816,N_1105,N_262);
nand U3817 (N_3817,N_1010,N_2826);
nand U3818 (N_3818,N_1122,N_976);
nor U3819 (N_3819,N_181,N_2734);
nand U3820 (N_3820,N_2575,N_408);
or U3821 (N_3821,N_842,N_1762);
xor U3822 (N_3822,N_2298,N_2562);
or U3823 (N_3823,N_2895,N_1003);
nor U3824 (N_3824,N_700,N_1082);
nand U3825 (N_3825,N_1579,N_362);
nor U3826 (N_3826,N_874,N_2977);
nand U3827 (N_3827,N_1245,N_1502);
nand U3828 (N_3828,N_2639,N_1315);
xor U3829 (N_3829,N_1030,N_1439);
and U3830 (N_3830,N_2170,N_2368);
nor U3831 (N_3831,N_1607,N_2441);
nand U3832 (N_3832,N_2063,N_379);
nand U3833 (N_3833,N_521,N_2925);
nand U3834 (N_3834,N_502,N_1511);
or U3835 (N_3835,N_1929,N_2258);
and U3836 (N_3836,N_1548,N_701);
nor U3837 (N_3837,N_861,N_2466);
nor U3838 (N_3838,N_2915,N_2570);
xnor U3839 (N_3839,N_1421,N_312);
or U3840 (N_3840,N_2253,N_77);
nand U3841 (N_3841,N_2412,N_1988);
or U3842 (N_3842,N_2557,N_2011);
and U3843 (N_3843,N_118,N_995);
or U3844 (N_3844,N_1854,N_31);
nor U3845 (N_3845,N_715,N_203);
nand U3846 (N_3846,N_845,N_1197);
nor U3847 (N_3847,N_104,N_626);
nor U3848 (N_3848,N_395,N_455);
and U3849 (N_3849,N_103,N_1830);
xnor U3850 (N_3850,N_2781,N_1238);
nand U3851 (N_3851,N_1593,N_1996);
nand U3852 (N_3852,N_1814,N_1080);
or U3853 (N_3853,N_2369,N_1862);
nor U3854 (N_3854,N_412,N_219);
and U3855 (N_3855,N_1309,N_1896);
or U3856 (N_3856,N_2621,N_2227);
nand U3857 (N_3857,N_706,N_1924);
or U3858 (N_3858,N_106,N_674);
nand U3859 (N_3859,N_1293,N_1280);
or U3860 (N_3860,N_172,N_1436);
nor U3861 (N_3861,N_760,N_1537);
nand U3862 (N_3862,N_528,N_542);
nor U3863 (N_3863,N_1477,N_438);
or U3864 (N_3864,N_2513,N_1673);
nand U3865 (N_3865,N_2856,N_1780);
nand U3866 (N_3866,N_2286,N_1125);
nor U3867 (N_3867,N_2630,N_668);
and U3868 (N_3868,N_1070,N_2288);
nand U3869 (N_3869,N_1522,N_1508);
nor U3870 (N_3870,N_1471,N_1848);
or U3871 (N_3871,N_1635,N_2257);
or U3872 (N_3872,N_1960,N_841);
or U3873 (N_3873,N_2316,N_2223);
nand U3874 (N_3874,N_1742,N_744);
nand U3875 (N_3875,N_1734,N_1832);
or U3876 (N_3876,N_1000,N_2272);
or U3877 (N_3877,N_2727,N_1462);
nand U3878 (N_3878,N_1386,N_1022);
xor U3879 (N_3879,N_1161,N_2058);
nor U3880 (N_3880,N_399,N_576);
and U3881 (N_3881,N_1216,N_2908);
and U3882 (N_3882,N_323,N_2243);
or U3883 (N_3883,N_1575,N_1114);
nand U3884 (N_3884,N_1223,N_2492);
xor U3885 (N_3885,N_2839,N_627);
or U3886 (N_3886,N_1528,N_2793);
and U3887 (N_3887,N_809,N_2012);
or U3888 (N_3888,N_1573,N_1791);
xor U3889 (N_3889,N_1267,N_1746);
xor U3890 (N_3890,N_2195,N_506);
and U3891 (N_3891,N_1719,N_601);
nor U3892 (N_3892,N_2785,N_1428);
nand U3893 (N_3893,N_1658,N_1797);
and U3894 (N_3894,N_2341,N_2039);
and U3895 (N_3895,N_554,N_2167);
xnor U3896 (N_3896,N_2329,N_123);
or U3897 (N_3897,N_1156,N_1188);
or U3898 (N_3898,N_2720,N_642);
nand U3899 (N_3899,N_102,N_1133);
and U3900 (N_3900,N_623,N_892);
or U3901 (N_3901,N_2032,N_2220);
and U3902 (N_3902,N_2121,N_1111);
and U3903 (N_3903,N_724,N_1493);
nor U3904 (N_3904,N_1097,N_1393);
nand U3905 (N_3905,N_2459,N_519);
nand U3906 (N_3906,N_1589,N_1644);
nand U3907 (N_3907,N_2180,N_2161);
nor U3908 (N_3908,N_1932,N_2573);
nor U3909 (N_3909,N_1553,N_2664);
and U3910 (N_3910,N_1683,N_2168);
and U3911 (N_3911,N_1680,N_2818);
nand U3912 (N_3912,N_249,N_1990);
nand U3913 (N_3913,N_2493,N_272);
nor U3914 (N_3914,N_1758,N_657);
xnor U3915 (N_3915,N_2442,N_862);
nand U3916 (N_3916,N_1072,N_1943);
or U3917 (N_3917,N_2022,N_2663);
or U3918 (N_3918,N_1338,N_2336);
or U3919 (N_3919,N_792,N_2587);
and U3920 (N_3920,N_533,N_1109);
nand U3921 (N_3921,N_1279,N_907);
and U3922 (N_3922,N_979,N_196);
xnor U3923 (N_3923,N_436,N_562);
or U3924 (N_3924,N_487,N_2649);
or U3925 (N_3925,N_2564,N_593);
and U3926 (N_3926,N_1600,N_352);
and U3927 (N_3927,N_2602,N_20);
and U3928 (N_3928,N_1458,N_829);
xnor U3929 (N_3929,N_1312,N_1043);
nor U3930 (N_3930,N_1696,N_2921);
or U3931 (N_3931,N_1776,N_1499);
nor U3932 (N_3932,N_1328,N_1968);
xor U3933 (N_3933,N_2592,N_96);
or U3934 (N_3934,N_2556,N_2312);
xnor U3935 (N_3935,N_558,N_116);
and U3936 (N_3936,N_927,N_2226);
nand U3937 (N_3937,N_866,N_34);
and U3938 (N_3938,N_2701,N_2292);
nand U3939 (N_3939,N_84,N_1740);
and U3940 (N_3940,N_2790,N_2447);
nand U3941 (N_3941,N_2819,N_2457);
or U3942 (N_3942,N_563,N_2346);
nand U3943 (N_3943,N_2698,N_1336);
nand U3944 (N_3944,N_244,N_1688);
or U3945 (N_3945,N_42,N_1134);
nor U3946 (N_3946,N_1012,N_450);
or U3947 (N_3947,N_1345,N_804);
and U3948 (N_3948,N_646,N_2420);
nor U3949 (N_3949,N_603,N_578);
nor U3950 (N_3950,N_1303,N_1828);
nor U3951 (N_3951,N_1195,N_2780);
nor U3952 (N_3952,N_2228,N_481);
nand U3953 (N_3953,N_233,N_2352);
and U3954 (N_3954,N_1465,N_2335);
nor U3955 (N_3955,N_146,N_676);
xnor U3956 (N_3956,N_1825,N_855);
and U3957 (N_3957,N_2373,N_2037);
nand U3958 (N_3958,N_1225,N_1572);
nor U3959 (N_3959,N_2881,N_2424);
nand U3960 (N_3960,N_1530,N_575);
or U3961 (N_3961,N_356,N_1269);
nand U3962 (N_3962,N_1086,N_52);
nand U3963 (N_3963,N_2924,N_1552);
or U3964 (N_3964,N_1379,N_2129);
and U3965 (N_3965,N_348,N_966);
and U3966 (N_3966,N_355,N_2256);
nand U3967 (N_3967,N_618,N_371);
xor U3968 (N_3968,N_2193,N_1446);
nand U3969 (N_3969,N_869,N_633);
and U3970 (N_3970,N_1112,N_2302);
or U3971 (N_3971,N_2700,N_1726);
xnor U3972 (N_3972,N_2205,N_2927);
and U3973 (N_3973,N_2201,N_2998);
nand U3974 (N_3974,N_871,N_859);
and U3975 (N_3975,N_2635,N_1306);
or U3976 (N_3976,N_2532,N_1982);
and U3977 (N_3977,N_1894,N_2766);
nand U3978 (N_3978,N_2358,N_1352);
or U3979 (N_3979,N_2945,N_656);
nand U3980 (N_3980,N_1371,N_2763);
nand U3981 (N_3981,N_518,N_107);
nand U3982 (N_3982,N_994,N_949);
xnor U3983 (N_3983,N_2112,N_2898);
nand U3984 (N_3984,N_1885,N_1240);
and U3985 (N_3985,N_1704,N_538);
and U3986 (N_3986,N_314,N_1849);
or U3987 (N_3987,N_1135,N_1297);
or U3988 (N_3988,N_2163,N_369);
and U3989 (N_3989,N_807,N_2593);
nand U3990 (N_3990,N_296,N_2315);
or U3991 (N_3991,N_678,N_697);
and U3992 (N_3992,N_393,N_1166);
nand U3993 (N_3993,N_340,N_2695);
or U3994 (N_3994,N_245,N_873);
nand U3995 (N_3995,N_1768,N_303);
xor U3996 (N_3996,N_1038,N_1544);
and U3997 (N_3997,N_931,N_1536);
nand U3998 (N_3998,N_137,N_1008);
and U3999 (N_3999,N_2904,N_2380);
nand U4000 (N_4000,N_1050,N_2667);
or U4001 (N_4001,N_2811,N_796);
nor U4002 (N_4002,N_877,N_914);
nand U4003 (N_4003,N_1806,N_1239);
nand U4004 (N_4004,N_373,N_2430);
nor U4005 (N_4005,N_2560,N_2411);
and U4006 (N_4006,N_2069,N_777);
or U4007 (N_4007,N_349,N_87);
and U4008 (N_4008,N_2436,N_2392);
nand U4009 (N_4009,N_2686,N_2809);
nand U4010 (N_4010,N_2711,N_2325);
or U4011 (N_4011,N_2810,N_2183);
and U4012 (N_4012,N_2778,N_2114);
nand U4013 (N_4013,N_2417,N_1749);
nand U4014 (N_4014,N_848,N_2095);
nor U4015 (N_4015,N_2628,N_2813);
nor U4016 (N_4016,N_756,N_2429);
nor U4017 (N_4017,N_2941,N_686);
or U4018 (N_4018,N_2297,N_543);
or U4019 (N_4019,N_1042,N_881);
nand U4020 (N_4020,N_2334,N_391);
nor U4021 (N_4021,N_1722,N_90);
nand U4022 (N_4022,N_661,N_2379);
or U4023 (N_4023,N_1414,N_1196);
nor U4024 (N_4024,N_201,N_680);
nand U4025 (N_4025,N_2036,N_926);
xnor U4026 (N_4026,N_2108,N_1957);
and U4027 (N_4027,N_1468,N_821);
nand U4028 (N_4028,N_1708,N_1747);
xnor U4029 (N_4029,N_791,N_1959);
nand U4030 (N_4030,N_22,N_2937);
nand U4031 (N_4031,N_790,N_1899);
or U4032 (N_4032,N_1339,N_2735);
and U4033 (N_4033,N_2289,N_561);
nor U4034 (N_4034,N_1855,N_1295);
nand U4035 (N_4035,N_1014,N_1750);
or U4036 (N_4036,N_2175,N_1718);
nor U4037 (N_4037,N_583,N_569);
and U4038 (N_4038,N_1840,N_343);
and U4039 (N_4039,N_284,N_1518);
xor U4040 (N_4040,N_345,N_311);
and U4041 (N_4041,N_444,N_2841);
nor U4042 (N_4042,N_2094,N_1927);
and U4043 (N_4043,N_2401,N_149);
nor U4044 (N_4044,N_2519,N_1454);
or U4045 (N_4045,N_769,N_1753);
or U4046 (N_4046,N_2719,N_666);
nor U4047 (N_4047,N_2067,N_579);
nor U4048 (N_4048,N_2706,N_1677);
xnor U4049 (N_4049,N_2031,N_1845);
or U4050 (N_4050,N_2864,N_590);
xor U4051 (N_4051,N_1995,N_281);
and U4052 (N_4052,N_2083,N_1037);
xnor U4053 (N_4053,N_2110,N_2333);
nand U4054 (N_4054,N_1198,N_378);
nand U4055 (N_4055,N_2625,N_2317);
nor U4056 (N_4056,N_772,N_1040);
and U4057 (N_4057,N_2303,N_2501);
and U4058 (N_4058,N_1220,N_370);
nand U4059 (N_4059,N_2674,N_1543);
or U4060 (N_4060,N_324,N_655);
and U4061 (N_4061,N_473,N_150);
xor U4062 (N_4062,N_1859,N_546);
xnor U4063 (N_4063,N_1126,N_1054);
xnor U4064 (N_4064,N_1435,N_1075);
nor U4065 (N_4065,N_727,N_1684);
or U4066 (N_4066,N_2959,N_595);
and U4067 (N_4067,N_1294,N_2693);
or U4068 (N_4068,N_863,N_1456);
nand U4069 (N_4069,N_1408,N_1816);
nand U4070 (N_4070,N_549,N_493);
nor U4071 (N_4071,N_2747,N_2611);
or U4072 (N_4072,N_1604,N_1622);
nand U4073 (N_4073,N_2482,N_213);
and U4074 (N_4074,N_1318,N_1154);
xor U4075 (N_4075,N_1286,N_1507);
xnor U4076 (N_4076,N_131,N_1380);
xor U4077 (N_4077,N_437,N_2822);
or U4078 (N_4078,N_160,N_1891);
and U4079 (N_4079,N_1047,N_2455);
and U4080 (N_4080,N_1425,N_174);
nand U4081 (N_4081,N_1703,N_2860);
nand U4082 (N_4082,N_1284,N_1595);
or U4083 (N_4083,N_1215,N_95);
xor U4084 (N_4084,N_186,N_257);
xor U4085 (N_4085,N_889,N_2101);
and U4086 (N_4086,N_1143,N_1987);
and U4087 (N_4087,N_1095,N_1681);
xor U4088 (N_4088,N_1015,N_962);
or U4089 (N_4089,N_2912,N_1214);
nand U4090 (N_4090,N_2523,N_2537);
xor U4091 (N_4091,N_1546,N_2347);
nand U4092 (N_4092,N_2293,N_2196);
or U4093 (N_4093,N_125,N_153);
nor U4094 (N_4094,N_191,N_2079);
nand U4095 (N_4095,N_1603,N_2460);
nand U4096 (N_4096,N_212,N_1564);
nor U4097 (N_4097,N_1160,N_2940);
or U4098 (N_4098,N_2578,N_1751);
or U4099 (N_4099,N_457,N_70);
nor U4100 (N_4100,N_2035,N_817);
nand U4101 (N_4101,N_722,N_498);
or U4102 (N_4102,N_1248,N_2805);
or U4103 (N_4103,N_2739,N_1774);
and U4104 (N_4104,N_1359,N_510);
and U4105 (N_4105,N_1623,N_1755);
or U4106 (N_4106,N_332,N_1686);
nand U4107 (N_4107,N_2414,N_958);
nand U4108 (N_4108,N_132,N_2596);
nand U4109 (N_4109,N_1478,N_2799);
nand U4110 (N_4110,N_1145,N_1616);
nand U4111 (N_4111,N_2920,N_2215);
xor U4112 (N_4112,N_2671,N_2918);
and U4113 (N_4113,N_2116,N_15);
and U4114 (N_4114,N_1412,N_2449);
and U4115 (N_4115,N_1190,N_2969);
and U4116 (N_4116,N_2248,N_2786);
nand U4117 (N_4117,N_1302,N_1841);
nand U4118 (N_4118,N_2715,N_415);
xnor U4119 (N_4119,N_1496,N_2893);
nor U4120 (N_4120,N_1342,N_898);
xnor U4121 (N_4121,N_846,N_1857);
nand U4122 (N_4122,N_2729,N_1324);
nand U4123 (N_4123,N_793,N_2696);
and U4124 (N_4124,N_1838,N_2218);
nor U4125 (N_4125,N_2760,N_113);
or U4126 (N_4126,N_410,N_1650);
nand U4127 (N_4127,N_2996,N_922);
xnor U4128 (N_4128,N_2479,N_2684);
and U4129 (N_4129,N_1029,N_2349);
or U4130 (N_4130,N_407,N_536);
xnor U4131 (N_4131,N_253,N_944);
or U4132 (N_4132,N_574,N_159);
and U4133 (N_4133,N_1993,N_1034);
or U4134 (N_4134,N_1618,N_695);
nor U4135 (N_4135,N_690,N_1226);
nand U4136 (N_4136,N_134,N_2612);
xnor U4137 (N_4137,N_824,N_1887);
nor U4138 (N_4138,N_882,N_2391);
nand U4139 (N_4139,N_868,N_2007);
or U4140 (N_4140,N_1733,N_2871);
nor U4141 (N_4141,N_902,N_189);
or U4142 (N_4142,N_368,N_1596);
or U4143 (N_4143,N_148,N_2566);
or U4144 (N_4144,N_1051,N_2757);
and U4145 (N_4145,N_2348,N_2816);
xnor U4146 (N_4146,N_2120,N_470);
nor U4147 (N_4147,N_2209,N_1131);
and U4148 (N_4148,N_2981,N_687);
or U4149 (N_4149,N_2554,N_86);
xor U4150 (N_4150,N_1709,N_2538);
or U4151 (N_4151,N_2244,N_220);
or U4152 (N_4152,N_2086,N_1059);
and U4153 (N_4153,N_1492,N_1621);
xnor U4154 (N_4154,N_1410,N_2681);
nand U4155 (N_4155,N_1192,N_211);
nor U4156 (N_4156,N_565,N_256);
nor U4157 (N_4157,N_1565,N_195);
nor U4158 (N_4158,N_1599,N_507);
or U4159 (N_4159,N_39,N_2976);
and U4160 (N_4160,N_1387,N_2989);
and U4161 (N_4161,N_799,N_1419);
and U4162 (N_4162,N_729,N_2085);
nand U4163 (N_4163,N_516,N_1268);
nor U4164 (N_4164,N_277,N_36);
nor U4165 (N_4165,N_1168,N_2143);
xor U4166 (N_4166,N_598,N_2239);
or U4167 (N_4167,N_2563,N_2050);
and U4168 (N_4168,N_560,N_264);
nand U4169 (N_4169,N_1185,N_1385);
xnor U4170 (N_4170,N_2399,N_1340);
or U4171 (N_4171,N_1661,N_2327);
or U4172 (N_4172,N_411,N_21);
or U4173 (N_4173,N_421,N_2923);
or U4174 (N_4174,N_490,N_813);
or U4175 (N_4175,N_2119,N_1210);
and U4176 (N_4176,N_2647,N_390);
xor U4177 (N_4177,N_707,N_529);
nand U4178 (N_4178,N_261,N_48);
nand U4179 (N_4179,N_1373,N_2280);
or U4180 (N_4180,N_199,N_564);
or U4181 (N_4181,N_2364,N_2382);
nand U4182 (N_4182,N_587,N_138);
and U4183 (N_4183,N_1676,N_2157);
nand U4184 (N_4184,N_784,N_1202);
and U4185 (N_4185,N_1975,N_1149);
or U4186 (N_4186,N_1884,N_1367);
or U4187 (N_4187,N_1234,N_2099);
and U4188 (N_4188,N_2426,N_2118);
nand U4189 (N_4189,N_187,N_2985);
nand U4190 (N_4190,N_2644,N_2808);
nand U4191 (N_4191,N_2040,N_737);
and U4192 (N_4192,N_1253,N_1636);
or U4193 (N_4193,N_1375,N_1991);
nand U4194 (N_4194,N_1066,N_2146);
nor U4195 (N_4195,N_1800,N_1520);
nor U4196 (N_4196,N_1679,N_757);
or U4197 (N_4197,N_1649,N_1115);
nor U4198 (N_4198,N_628,N_2351);
nand U4199 (N_4199,N_967,N_1423);
nand U4200 (N_4200,N_806,N_2887);
or U4201 (N_4201,N_98,N_2122);
nand U4202 (N_4202,N_1997,N_904);
and U4203 (N_4203,N_1074,N_2267);
xor U4204 (N_4204,N_2404,N_100);
or U4205 (N_4205,N_1175,N_1139);
and U4206 (N_4206,N_1882,N_2855);
and U4207 (N_4207,N_653,N_1713);
nand U4208 (N_4208,N_380,N_1327);
nand U4209 (N_4209,N_282,N_1721);
and U4210 (N_4210,N_1954,N_2736);
nor U4211 (N_4211,N_1257,N_2590);
nor U4212 (N_4212,N_1910,N_2928);
nor U4213 (N_4213,N_2434,N_2377);
nand U4214 (N_4214,N_1809,N_2159);
and U4215 (N_4215,N_1187,N_2047);
xnor U4216 (N_4216,N_394,N_2054);
or U4217 (N_4217,N_2437,N_2687);
or U4218 (N_4218,N_1415,N_2467);
and U4219 (N_4219,N_736,N_2023);
nand U4220 (N_4220,N_1321,N_1624);
nand U4221 (N_4221,N_1545,N_1405);
nor U4222 (N_4222,N_2343,N_2605);
nand U4223 (N_4223,N_40,N_541);
nand U4224 (N_4224,N_2506,N_616);
xnor U4225 (N_4225,N_830,N_2474);
nand U4226 (N_4226,N_2182,N_1316);
or U4227 (N_4227,N_1909,N_948);
xor U4228 (N_4228,N_2204,N_1984);
and U4229 (N_4229,N_1802,N_2929);
nand U4230 (N_4230,N_2691,N_316);
and U4231 (N_4231,N_865,N_1937);
nand U4232 (N_4232,N_73,N_1121);
and U4233 (N_4233,N_774,N_2585);
or U4234 (N_4234,N_1009,N_573);
and U4235 (N_4235,N_382,N_2714);
nor U4236 (N_4236,N_1558,N_2633);
nand U4237 (N_4237,N_1501,N_2844);
xor U4238 (N_4238,N_747,N_459);
and U4239 (N_4239,N_753,N_1429);
and U4240 (N_4240,N_99,N_1420);
or U4241 (N_4241,N_294,N_699);
and U4242 (N_4242,N_1020,N_1392);
and U4243 (N_4243,N_1919,N_2006);
and U4244 (N_4244,N_2277,N_377);
nor U4245 (N_4245,N_2726,N_445);
nor U4246 (N_4246,N_1555,N_1773);
or U4247 (N_4247,N_2531,N_2400);
or U4248 (N_4248,N_1399,N_2553);
nand U4249 (N_4249,N_25,N_908);
nand U4250 (N_4250,N_1867,N_767);
nand U4251 (N_4251,N_1994,N_539);
nor U4252 (N_4252,N_2339,N_1732);
or U4253 (N_4253,N_870,N_2806);
xnor U4254 (N_4254,N_2699,N_1535);
and U4255 (N_4255,N_2973,N_1907);
and U4256 (N_4256,N_182,N_1692);
or U4257 (N_4257,N_1426,N_1856);
nand U4258 (N_4258,N_2234,N_222);
nand U4259 (N_4259,N_2494,N_2070);
and U4260 (N_4260,N_2109,N_453);
or U4261 (N_4261,N_2745,N_721);
nor U4262 (N_4262,N_920,N_2737);
and U4263 (N_4263,N_166,N_512);
xor U4264 (N_4264,N_464,N_1211);
nand U4265 (N_4265,N_1539,N_1179);
nand U4266 (N_4266,N_2721,N_2732);
nand U4267 (N_4267,N_748,N_1510);
nor U4268 (N_4268,N_553,N_2916);
nor U4269 (N_4269,N_164,N_2690);
nor U4270 (N_4270,N_2545,N_1695);
nand U4271 (N_4271,N_2597,N_1617);
and U4272 (N_4272,N_1583,N_2097);
nand U4273 (N_4273,N_884,N_739);
nand U4274 (N_4274,N_1785,N_2489);
xor U4275 (N_4275,N_330,N_1266);
xor U4276 (N_4276,N_2823,N_1237);
and U4277 (N_4277,N_669,N_781);
or U4278 (N_4278,N_1965,N_1723);
and U4279 (N_4279,N_523,N_2263);
nand U4280 (N_4280,N_198,N_606);
nor U4281 (N_4281,N_2987,N_2133);
or U4282 (N_4282,N_673,N_932);
nand U4283 (N_4283,N_2135,N_2797);
and U4284 (N_4284,N_60,N_2961);
nand U4285 (N_4285,N_451,N_1307);
nor U4286 (N_4286,N_68,N_2018);
or U4287 (N_4287,N_1069,N_2740);
nand U4288 (N_4288,N_136,N_1928);
and U4289 (N_4289,N_1782,N_2446);
or U4290 (N_4290,N_833,N_864);
nor U4291 (N_4291,N_1781,N_1063);
and U4292 (N_4292,N_392,N_2073);
and U4293 (N_4293,N_2657,N_1921);
or U4294 (N_4294,N_1529,N_2296);
nand U4295 (N_4295,N_571,N_1562);
or U4296 (N_4296,N_2046,N_1999);
and U4297 (N_4297,N_309,N_550);
nor U4298 (N_4298,N_1851,N_2148);
and U4299 (N_4299,N_1724,N_2515);
or U4300 (N_4300,N_1218,N_2718);
and U4301 (N_4301,N_2834,N_1958);
xor U4302 (N_4302,N_1690,N_1433);
nand U4303 (N_4303,N_63,N_2836);
xnor U4304 (N_4304,N_55,N_2464);
or U4305 (N_4305,N_2166,N_265);
nor U4306 (N_4306,N_2304,N_2473);
nor U4307 (N_4307,N_45,N_49);
xnor U4308 (N_4308,N_1182,N_418);
or U4309 (N_4309,N_1004,N_2072);
nor U4310 (N_4310,N_2324,N_631);
and U4311 (N_4311,N_2890,N_532);
xor U4312 (N_4312,N_1687,N_1727);
nor U4313 (N_4313,N_801,N_1440);
xnor U4314 (N_4314,N_778,N_582);
or U4315 (N_4315,N_2906,N_1118);
nor U4316 (N_4316,N_702,N_2456);
xor U4317 (N_4317,N_1431,N_2151);
nand U4318 (N_4318,N_1163,N_1801);
nor U4319 (N_4319,N_1941,N_1231);
nor U4320 (N_4320,N_936,N_500);
or U4321 (N_4321,N_2966,N_556);
and U4322 (N_4322,N_67,N_986);
or U4323 (N_4323,N_759,N_568);
and U4324 (N_4324,N_2055,N_2198);
or U4325 (N_4325,N_2322,N_625);
nor U4326 (N_4326,N_2332,N_933);
nand U4327 (N_4327,N_1759,N_1453);
nor U4328 (N_4328,N_2355,N_1364);
nor U4329 (N_4329,N_2591,N_2075);
and U4330 (N_4330,N_2656,N_92);
and U4331 (N_4331,N_1189,N_8);
xor U4332 (N_4332,N_2331,N_1930);
and U4333 (N_4333,N_599,N_1007);
or U4334 (N_4334,N_1714,N_494);
xor U4335 (N_4335,N_12,N_177);
nand U4336 (N_4336,N_1093,N_1540);
or U4337 (N_4337,N_924,N_2240);
nor U4338 (N_4338,N_1171,N_810);
or U4339 (N_4339,N_2926,N_1432);
nand U4340 (N_4340,N_1113,N_1263);
and U4341 (N_4341,N_1274,N_1793);
or U4342 (N_4342,N_2565,N_2418);
or U4343 (N_4343,N_1506,N_1942);
or U4344 (N_4344,N_495,N_337);
nor U4345 (N_4345,N_50,N_375);
nand U4346 (N_4346,N_2178,N_2281);
nand U4347 (N_4347,N_33,N_1760);
nor U4348 (N_4348,N_140,N_905);
and U4349 (N_4349,N_2646,N_2677);
and U4350 (N_4350,N_640,N_460);
and U4351 (N_4351,N_1563,N_989);
nor U4352 (N_4352,N_2606,N_2026);
and U4353 (N_4353,N_1892,N_1881);
nand U4354 (N_4354,N_1915,N_5);
xnor U4355 (N_4355,N_2555,N_1743);
nor U4356 (N_4356,N_2275,N_637);
and U4357 (N_4357,N_670,N_298);
and U4358 (N_4358,N_2642,N_2265);
or U4359 (N_4359,N_2255,N_2448);
nor U4360 (N_4360,N_404,N_1779);
xor U4361 (N_4361,N_2199,N_1348);
nor U4362 (N_4362,N_694,N_2273);
and U4363 (N_4363,N_1260,N_422);
nor U4364 (N_4364,N_1495,N_2174);
nand U4365 (N_4365,N_1876,N_2608);
nand U4366 (N_4366,N_1016,N_1466);
nor U4367 (N_4367,N_293,N_886);
nand U4368 (N_4368,N_1955,N_2269);
or U4369 (N_4369,N_890,N_2142);
nor U4370 (N_4370,N_2375,N_1787);
and U4371 (N_4371,N_1033,N_2062);
nor U4372 (N_4372,N_1731,N_1447);
and U4373 (N_4373,N_2982,N_2169);
or U4374 (N_4374,N_900,N_1833);
xnor U4375 (N_4375,N_501,N_1391);
nand U4376 (N_4376,N_2232,N_2750);
and U4377 (N_4377,N_1028,N_10);
xnor U4378 (N_4378,N_111,N_832);
and U4379 (N_4379,N_2282,N_2020);
xnor U4380 (N_4380,N_114,N_604);
nor U4381 (N_4381,N_1647,N_1177);
nand U4382 (N_4382,N_2746,N_1402);
and U4383 (N_4383,N_80,N_2383);
nor U4384 (N_4384,N_2892,N_2541);
nand U4385 (N_4385,N_367,N_2356);
or U4386 (N_4386,N_214,N_1883);
and U4387 (N_4387,N_621,N_241);
nor U4388 (N_4388,N_2595,N_2405);
nand U4389 (N_4389,N_711,N_1605);
or U4390 (N_4390,N_1590,N_1657);
nor U4391 (N_4391,N_1488,N_794);
nor U4392 (N_4392,N_2618,N_4);
or U4393 (N_4393,N_155,N_165);
and U4394 (N_4394,N_658,N_2705);
and U4395 (N_4395,N_1021,N_1363);
or U4396 (N_4396,N_643,N_2394);
nor U4397 (N_4397,N_1756,N_1311);
xor U4398 (N_4398,N_2682,N_1242);
nor U4399 (N_4399,N_2301,N_849);
nand U4400 (N_4400,N_754,N_215);
and U4401 (N_4401,N_1103,N_619);
nor U4402 (N_4402,N_2956,N_1847);
nand U4403 (N_4403,N_381,N_207);
nor U4404 (N_4404,N_651,N_2469);
and U4405 (N_4405,N_2984,N_1282);
and U4406 (N_4406,N_1344,N_2576);
nor U4407 (N_4407,N_1397,N_954);
nor U4408 (N_4408,N_768,N_2650);
nand U4409 (N_4409,N_928,N_2594);
nand U4410 (N_4410,N_677,N_2861);
or U4411 (N_4411,N_2131,N_762);
nor U4412 (N_4412,N_2224,N_247);
nor U4413 (N_4413,N_427,N_1147);
nand U4414 (N_4414,N_129,N_586);
and U4415 (N_4415,N_2370,N_831);
nor U4416 (N_4416,N_171,N_1934);
nor U4417 (N_4417,N_2155,N_2815);
nor U4418 (N_4418,N_2486,N_2002);
nand U4419 (N_4419,N_448,N_26);
nor U4420 (N_4420,N_364,N_1922);
xor U4421 (N_4421,N_1486,N_1823);
nand U4422 (N_4422,N_209,N_46);
nor U4423 (N_4423,N_527,N_2571);
nor U4424 (N_4424,N_2800,N_1706);
nand U4425 (N_4425,N_2250,N_1669);
nand U4426 (N_4426,N_2938,N_1208);
and U4427 (N_4427,N_1310,N_2415);
and U4428 (N_4428,N_1998,N_1620);
or U4429 (N_4429,N_641,N_336);
nor U4430 (N_4430,N_2624,N_51);
or U4431 (N_4431,N_2788,N_37);
nor U4432 (N_4432,N_2609,N_2598);
and U4433 (N_4433,N_2891,N_1648);
nor U4434 (N_4434,N_2191,N_1587);
nand U4435 (N_4435,N_2528,N_2748);
and U4436 (N_4436,N_2106,N_2270);
or U4437 (N_4437,N_432,N_992);
and U4438 (N_4438,N_746,N_2300);
nand U4439 (N_4439,N_1343,N_2662);
nand U4440 (N_4440,N_1920,N_2021);
nand U4441 (N_4441,N_2422,N_1807);
nor U4442 (N_4442,N_782,N_1413);
nand U4443 (N_4443,N_1272,N_2387);
nor U4444 (N_4444,N_522,N_820);
or U4445 (N_4445,N_1494,N_1962);
nor U4446 (N_4446,N_2153,N_1509);
and U4447 (N_4447,N_1064,N_2359);
nand U4448 (N_4448,N_1916,N_1512);
and U4449 (N_4449,N_635,N_439);
xor U4450 (N_4450,N_425,N_2512);
or U4451 (N_4451,N_173,N_430);
nand U4452 (N_4452,N_1827,N_1933);
or U4453 (N_4453,N_2939,N_1255);
nand U4454 (N_4454,N_2219,N_151);
nor U4455 (N_4455,N_2096,N_1533);
and U4456 (N_4456,N_2005,N_2689);
and U4457 (N_4457,N_1745,N_1055);
nand U4458 (N_4458,N_734,N_2529);
and U4459 (N_4459,N_878,N_82);
nor U4460 (N_4460,N_1893,N_888);
or U4461 (N_4461,N_1204,N_452);
and U4462 (N_4462,N_142,N_1831);
xor U4463 (N_4463,N_2522,N_2979);
and U4464 (N_4464,N_2876,N_745);
and U4465 (N_4465,N_197,N_254);
and U4466 (N_4466,N_2759,N_1247);
nand U4467 (N_4467,N_1914,N_1966);
nand U4468 (N_4468,N_1479,N_346);
or U4469 (N_4469,N_1739,N_1102);
nor U4470 (N_4470,N_893,N_1347);
nor U4471 (N_4471,N_1557,N_1452);
and U4472 (N_4472,N_441,N_1936);
xnor U4473 (N_4473,N_743,N_1475);
and U4474 (N_4474,N_2614,N_2514);
nand U4475 (N_4475,N_2310,N_1141);
nand U4476 (N_4476,N_1369,N_1394);
and U4477 (N_4477,N_1422,N_2481);
nor U4478 (N_4478,N_683,N_1483);
and U4479 (N_4479,N_555,N_2149);
and U4480 (N_4480,N_2061,N_1777);
nand U4481 (N_4481,N_2056,N_805);
nand U4482 (N_4482,N_2084,N_328);
nand U4483 (N_4483,N_232,N_158);
or U4484 (N_4484,N_2237,N_18);
nor U4485 (N_4485,N_789,N_2930);
or U4486 (N_4486,N_1170,N_1039);
nand U4487 (N_4487,N_2137,N_2902);
or U4488 (N_4488,N_2309,N_1560);
xnor U4489 (N_4489,N_2665,N_816);
or U4490 (N_4490,N_401,N_785);
nor U4491 (N_4491,N_1786,N_955);
nor U4492 (N_4492,N_1365,N_2103);
and U4493 (N_4493,N_2643,N_2617);
nor U4494 (N_4494,N_1106,N_2271);
or U4495 (N_4495,N_69,N_227);
xnor U4496 (N_4496,N_2648,N_2395);
nand U4497 (N_4497,N_714,N_1818);
and U4498 (N_4498,N_1656,N_2828);
nand U4499 (N_4499,N_698,N_2440);
and U4500 (N_4500,N_826,N_2786);
or U4501 (N_4501,N_2668,N_1727);
nand U4502 (N_4502,N_1772,N_756);
nand U4503 (N_4503,N_1649,N_253);
nor U4504 (N_4504,N_238,N_790);
or U4505 (N_4505,N_128,N_2327);
and U4506 (N_4506,N_2904,N_1619);
and U4507 (N_4507,N_1649,N_2719);
and U4508 (N_4508,N_1290,N_1450);
nor U4509 (N_4509,N_686,N_380);
nand U4510 (N_4510,N_1958,N_1413);
or U4511 (N_4511,N_1012,N_2964);
xor U4512 (N_4512,N_1592,N_366);
nand U4513 (N_4513,N_1978,N_1578);
and U4514 (N_4514,N_2630,N_1890);
and U4515 (N_4515,N_2900,N_507);
nand U4516 (N_4516,N_2706,N_1865);
nand U4517 (N_4517,N_1649,N_899);
nand U4518 (N_4518,N_2624,N_1232);
nor U4519 (N_4519,N_1749,N_1978);
xor U4520 (N_4520,N_1953,N_2890);
xor U4521 (N_4521,N_1723,N_759);
or U4522 (N_4522,N_58,N_754);
nor U4523 (N_4523,N_602,N_1284);
and U4524 (N_4524,N_997,N_162);
nor U4525 (N_4525,N_1523,N_1872);
or U4526 (N_4526,N_1438,N_712);
nand U4527 (N_4527,N_2677,N_1968);
xnor U4528 (N_4528,N_2798,N_2451);
xor U4529 (N_4529,N_2356,N_1835);
nor U4530 (N_4530,N_2566,N_444);
nand U4531 (N_4531,N_2138,N_1028);
nor U4532 (N_4532,N_835,N_862);
nor U4533 (N_4533,N_712,N_2681);
nor U4534 (N_4534,N_2014,N_1454);
and U4535 (N_4535,N_2820,N_2117);
nor U4536 (N_4536,N_1728,N_2006);
nand U4537 (N_4537,N_80,N_1204);
or U4538 (N_4538,N_2871,N_221);
and U4539 (N_4539,N_1778,N_386);
nor U4540 (N_4540,N_2340,N_1127);
or U4541 (N_4541,N_757,N_2186);
nor U4542 (N_4542,N_2382,N_1672);
or U4543 (N_4543,N_2784,N_1747);
xor U4544 (N_4544,N_2634,N_1706);
or U4545 (N_4545,N_1393,N_292);
nand U4546 (N_4546,N_287,N_101);
and U4547 (N_4547,N_2481,N_2657);
and U4548 (N_4548,N_2459,N_62);
and U4549 (N_4549,N_2227,N_2800);
and U4550 (N_4550,N_144,N_533);
or U4551 (N_4551,N_512,N_2390);
nor U4552 (N_4552,N_2285,N_1951);
nor U4553 (N_4553,N_908,N_1216);
or U4554 (N_4554,N_1155,N_460);
nor U4555 (N_4555,N_1391,N_1095);
or U4556 (N_4556,N_448,N_2234);
xnor U4557 (N_4557,N_2948,N_457);
nor U4558 (N_4558,N_2152,N_2159);
nor U4559 (N_4559,N_987,N_206);
or U4560 (N_4560,N_790,N_2055);
nand U4561 (N_4561,N_973,N_1380);
nand U4562 (N_4562,N_2963,N_1209);
and U4563 (N_4563,N_741,N_2553);
and U4564 (N_4564,N_988,N_640);
and U4565 (N_4565,N_2656,N_2253);
nand U4566 (N_4566,N_309,N_2814);
or U4567 (N_4567,N_667,N_49);
nor U4568 (N_4568,N_2251,N_1360);
and U4569 (N_4569,N_2944,N_1852);
nand U4570 (N_4570,N_763,N_1046);
and U4571 (N_4571,N_203,N_54);
nand U4572 (N_4572,N_2366,N_1831);
and U4573 (N_4573,N_1045,N_943);
nor U4574 (N_4574,N_1119,N_630);
and U4575 (N_4575,N_2625,N_345);
nand U4576 (N_4576,N_962,N_1847);
or U4577 (N_4577,N_1455,N_245);
or U4578 (N_4578,N_1805,N_1462);
and U4579 (N_4579,N_1002,N_906);
or U4580 (N_4580,N_1373,N_870);
nor U4581 (N_4581,N_640,N_1930);
and U4582 (N_4582,N_2469,N_2697);
or U4583 (N_4583,N_1710,N_104);
or U4584 (N_4584,N_1492,N_1306);
nor U4585 (N_4585,N_2774,N_810);
nor U4586 (N_4586,N_2009,N_580);
xnor U4587 (N_4587,N_2257,N_1429);
nor U4588 (N_4588,N_2592,N_454);
nor U4589 (N_4589,N_2304,N_911);
and U4590 (N_4590,N_2891,N_1529);
xor U4591 (N_4591,N_1995,N_646);
and U4592 (N_4592,N_1812,N_2252);
or U4593 (N_4593,N_613,N_1141);
or U4594 (N_4594,N_1713,N_1871);
or U4595 (N_4595,N_1747,N_467);
or U4596 (N_4596,N_1914,N_2502);
nand U4597 (N_4597,N_1118,N_599);
nand U4598 (N_4598,N_1208,N_2702);
nand U4599 (N_4599,N_2399,N_1211);
or U4600 (N_4600,N_1276,N_353);
nand U4601 (N_4601,N_1536,N_1549);
and U4602 (N_4602,N_1022,N_350);
or U4603 (N_4603,N_2937,N_2352);
xnor U4604 (N_4604,N_233,N_2259);
and U4605 (N_4605,N_510,N_1866);
nand U4606 (N_4606,N_835,N_2991);
nand U4607 (N_4607,N_105,N_2655);
or U4608 (N_4608,N_334,N_2024);
nor U4609 (N_4609,N_1213,N_2654);
nand U4610 (N_4610,N_1647,N_2553);
or U4611 (N_4611,N_1793,N_1440);
or U4612 (N_4612,N_1938,N_463);
nand U4613 (N_4613,N_921,N_194);
and U4614 (N_4614,N_1479,N_2526);
or U4615 (N_4615,N_2804,N_1912);
or U4616 (N_4616,N_2198,N_2380);
and U4617 (N_4617,N_1468,N_1520);
or U4618 (N_4618,N_1553,N_661);
nor U4619 (N_4619,N_2752,N_2858);
or U4620 (N_4620,N_409,N_2494);
or U4621 (N_4621,N_2610,N_1693);
nand U4622 (N_4622,N_912,N_2159);
or U4623 (N_4623,N_1740,N_1963);
and U4624 (N_4624,N_2555,N_75);
or U4625 (N_4625,N_564,N_268);
nand U4626 (N_4626,N_494,N_2998);
nor U4627 (N_4627,N_1328,N_2151);
nor U4628 (N_4628,N_1652,N_971);
and U4629 (N_4629,N_1269,N_39);
nor U4630 (N_4630,N_1523,N_701);
nand U4631 (N_4631,N_2351,N_13);
nand U4632 (N_4632,N_947,N_1133);
nand U4633 (N_4633,N_292,N_2238);
and U4634 (N_4634,N_757,N_2767);
or U4635 (N_4635,N_471,N_1342);
or U4636 (N_4636,N_568,N_659);
and U4637 (N_4637,N_2522,N_277);
nor U4638 (N_4638,N_1908,N_2105);
xor U4639 (N_4639,N_2372,N_2960);
nand U4640 (N_4640,N_1373,N_742);
nor U4641 (N_4641,N_1470,N_2518);
and U4642 (N_4642,N_1099,N_658);
or U4643 (N_4643,N_696,N_193);
and U4644 (N_4644,N_4,N_2503);
or U4645 (N_4645,N_1856,N_2433);
and U4646 (N_4646,N_2217,N_2764);
nand U4647 (N_4647,N_2831,N_636);
or U4648 (N_4648,N_639,N_529);
nor U4649 (N_4649,N_637,N_2658);
nor U4650 (N_4650,N_2520,N_2550);
nand U4651 (N_4651,N_343,N_986);
nand U4652 (N_4652,N_2335,N_726);
nor U4653 (N_4653,N_1509,N_2942);
and U4654 (N_4654,N_912,N_2905);
or U4655 (N_4655,N_2589,N_2259);
nor U4656 (N_4656,N_2801,N_406);
and U4657 (N_4657,N_2411,N_2654);
nand U4658 (N_4658,N_2027,N_913);
nor U4659 (N_4659,N_889,N_2640);
or U4660 (N_4660,N_1105,N_2217);
nor U4661 (N_4661,N_32,N_2177);
or U4662 (N_4662,N_1959,N_1238);
nand U4663 (N_4663,N_801,N_595);
nand U4664 (N_4664,N_2823,N_2768);
and U4665 (N_4665,N_1454,N_2579);
and U4666 (N_4666,N_531,N_2180);
or U4667 (N_4667,N_1917,N_1131);
xnor U4668 (N_4668,N_188,N_1570);
xor U4669 (N_4669,N_2261,N_2751);
nand U4670 (N_4670,N_404,N_611);
xnor U4671 (N_4671,N_155,N_69);
nand U4672 (N_4672,N_2888,N_1225);
nor U4673 (N_4673,N_345,N_2949);
and U4674 (N_4674,N_2344,N_360);
nor U4675 (N_4675,N_2041,N_2783);
or U4676 (N_4676,N_1023,N_959);
and U4677 (N_4677,N_264,N_2859);
or U4678 (N_4678,N_1759,N_1568);
and U4679 (N_4679,N_2568,N_767);
or U4680 (N_4680,N_248,N_1451);
nor U4681 (N_4681,N_762,N_2519);
or U4682 (N_4682,N_2033,N_2882);
nor U4683 (N_4683,N_2597,N_2941);
xor U4684 (N_4684,N_1759,N_2170);
nor U4685 (N_4685,N_909,N_2730);
and U4686 (N_4686,N_2563,N_2278);
nor U4687 (N_4687,N_758,N_2115);
or U4688 (N_4688,N_1153,N_268);
and U4689 (N_4689,N_285,N_667);
and U4690 (N_4690,N_2276,N_1895);
nor U4691 (N_4691,N_1626,N_2262);
nand U4692 (N_4692,N_1398,N_132);
and U4693 (N_4693,N_2605,N_1082);
and U4694 (N_4694,N_1095,N_1138);
nor U4695 (N_4695,N_1420,N_2395);
or U4696 (N_4696,N_777,N_2386);
and U4697 (N_4697,N_1834,N_1828);
or U4698 (N_4698,N_1340,N_1407);
or U4699 (N_4699,N_1508,N_1488);
nor U4700 (N_4700,N_2599,N_2587);
and U4701 (N_4701,N_1237,N_2464);
nor U4702 (N_4702,N_194,N_903);
and U4703 (N_4703,N_1712,N_1929);
nand U4704 (N_4704,N_267,N_301);
nor U4705 (N_4705,N_211,N_1099);
nor U4706 (N_4706,N_2918,N_1286);
or U4707 (N_4707,N_1859,N_1352);
and U4708 (N_4708,N_1608,N_1505);
and U4709 (N_4709,N_1131,N_2581);
nor U4710 (N_4710,N_1589,N_886);
nand U4711 (N_4711,N_2771,N_47);
nor U4712 (N_4712,N_51,N_187);
nor U4713 (N_4713,N_1954,N_313);
xnor U4714 (N_4714,N_2622,N_1249);
nor U4715 (N_4715,N_366,N_381);
xor U4716 (N_4716,N_2552,N_1272);
nor U4717 (N_4717,N_471,N_2515);
or U4718 (N_4718,N_1306,N_205);
nor U4719 (N_4719,N_2594,N_1212);
and U4720 (N_4720,N_1480,N_2310);
nor U4721 (N_4721,N_2530,N_254);
or U4722 (N_4722,N_964,N_247);
or U4723 (N_4723,N_2113,N_2267);
nor U4724 (N_4724,N_1264,N_1763);
or U4725 (N_4725,N_697,N_2308);
nor U4726 (N_4726,N_903,N_671);
and U4727 (N_4727,N_1168,N_501);
nand U4728 (N_4728,N_198,N_2220);
nor U4729 (N_4729,N_1852,N_2257);
nand U4730 (N_4730,N_619,N_782);
and U4731 (N_4731,N_1007,N_1454);
and U4732 (N_4732,N_236,N_1295);
nand U4733 (N_4733,N_1459,N_1525);
nor U4734 (N_4734,N_2773,N_1958);
nor U4735 (N_4735,N_941,N_1323);
or U4736 (N_4736,N_92,N_1069);
or U4737 (N_4737,N_1437,N_1915);
nor U4738 (N_4738,N_9,N_1926);
and U4739 (N_4739,N_1518,N_1480);
nor U4740 (N_4740,N_2386,N_1273);
and U4741 (N_4741,N_42,N_2060);
or U4742 (N_4742,N_1303,N_128);
or U4743 (N_4743,N_2338,N_1483);
nor U4744 (N_4744,N_470,N_1852);
and U4745 (N_4745,N_1187,N_1198);
or U4746 (N_4746,N_413,N_1867);
and U4747 (N_4747,N_2927,N_2287);
and U4748 (N_4748,N_1962,N_72);
xor U4749 (N_4749,N_86,N_2158);
nand U4750 (N_4750,N_1576,N_2960);
nor U4751 (N_4751,N_726,N_938);
or U4752 (N_4752,N_1167,N_1422);
nand U4753 (N_4753,N_2196,N_2136);
nand U4754 (N_4754,N_1619,N_1488);
nand U4755 (N_4755,N_473,N_2742);
nor U4756 (N_4756,N_2075,N_2028);
or U4757 (N_4757,N_2458,N_1455);
nand U4758 (N_4758,N_1289,N_2218);
nand U4759 (N_4759,N_1538,N_1758);
and U4760 (N_4760,N_908,N_1967);
nand U4761 (N_4761,N_2640,N_1461);
nand U4762 (N_4762,N_241,N_1153);
nor U4763 (N_4763,N_2797,N_2659);
xnor U4764 (N_4764,N_2213,N_2728);
or U4765 (N_4765,N_2633,N_438);
nand U4766 (N_4766,N_754,N_1023);
nor U4767 (N_4767,N_2305,N_259);
nor U4768 (N_4768,N_1833,N_1748);
or U4769 (N_4769,N_2245,N_365);
nand U4770 (N_4770,N_1147,N_765);
xor U4771 (N_4771,N_1337,N_320);
nand U4772 (N_4772,N_611,N_1416);
and U4773 (N_4773,N_2807,N_1460);
nor U4774 (N_4774,N_2002,N_879);
or U4775 (N_4775,N_1531,N_1183);
or U4776 (N_4776,N_1474,N_2893);
xnor U4777 (N_4777,N_1454,N_1677);
or U4778 (N_4778,N_2841,N_2765);
nand U4779 (N_4779,N_1213,N_353);
and U4780 (N_4780,N_1892,N_696);
xnor U4781 (N_4781,N_2886,N_1792);
or U4782 (N_4782,N_2334,N_1851);
nand U4783 (N_4783,N_574,N_167);
nor U4784 (N_4784,N_2262,N_1104);
nor U4785 (N_4785,N_2037,N_1390);
or U4786 (N_4786,N_1958,N_1165);
nand U4787 (N_4787,N_2397,N_2131);
xor U4788 (N_4788,N_2842,N_1737);
nand U4789 (N_4789,N_2450,N_2310);
and U4790 (N_4790,N_2153,N_640);
and U4791 (N_4791,N_317,N_2439);
xor U4792 (N_4792,N_1808,N_2985);
or U4793 (N_4793,N_244,N_1883);
nor U4794 (N_4794,N_268,N_2378);
xor U4795 (N_4795,N_2397,N_1262);
nor U4796 (N_4796,N_142,N_2106);
nor U4797 (N_4797,N_2212,N_603);
or U4798 (N_4798,N_2566,N_2632);
nand U4799 (N_4799,N_2697,N_2947);
or U4800 (N_4800,N_479,N_2175);
nand U4801 (N_4801,N_2850,N_134);
and U4802 (N_4802,N_2893,N_942);
nand U4803 (N_4803,N_2201,N_102);
and U4804 (N_4804,N_2567,N_2904);
nor U4805 (N_4805,N_945,N_1810);
and U4806 (N_4806,N_2703,N_1422);
xor U4807 (N_4807,N_991,N_1302);
nand U4808 (N_4808,N_1674,N_674);
nor U4809 (N_4809,N_2314,N_886);
and U4810 (N_4810,N_2065,N_1080);
or U4811 (N_4811,N_2060,N_1011);
or U4812 (N_4812,N_219,N_1913);
nor U4813 (N_4813,N_1160,N_2302);
nor U4814 (N_4814,N_2424,N_1512);
xnor U4815 (N_4815,N_1758,N_1691);
and U4816 (N_4816,N_846,N_2499);
and U4817 (N_4817,N_2945,N_1716);
nand U4818 (N_4818,N_1698,N_2711);
nand U4819 (N_4819,N_1265,N_2688);
nor U4820 (N_4820,N_2947,N_332);
nor U4821 (N_4821,N_936,N_1114);
or U4822 (N_4822,N_1825,N_1960);
and U4823 (N_4823,N_2253,N_1176);
or U4824 (N_4824,N_1750,N_1041);
nor U4825 (N_4825,N_2077,N_1702);
or U4826 (N_4826,N_449,N_586);
or U4827 (N_4827,N_1881,N_564);
nor U4828 (N_4828,N_617,N_649);
nor U4829 (N_4829,N_144,N_1018);
or U4830 (N_4830,N_2521,N_2264);
and U4831 (N_4831,N_1067,N_814);
nand U4832 (N_4832,N_2109,N_84);
or U4833 (N_4833,N_2868,N_2130);
nand U4834 (N_4834,N_2442,N_1722);
and U4835 (N_4835,N_15,N_2119);
nand U4836 (N_4836,N_486,N_2407);
and U4837 (N_4837,N_2545,N_484);
nor U4838 (N_4838,N_1875,N_968);
nor U4839 (N_4839,N_846,N_720);
nor U4840 (N_4840,N_1735,N_953);
or U4841 (N_4841,N_204,N_760);
or U4842 (N_4842,N_1612,N_79);
nor U4843 (N_4843,N_568,N_470);
or U4844 (N_4844,N_872,N_1265);
and U4845 (N_4845,N_2197,N_2558);
nor U4846 (N_4846,N_243,N_943);
nor U4847 (N_4847,N_2358,N_2965);
nor U4848 (N_4848,N_2183,N_311);
nor U4849 (N_4849,N_1266,N_1020);
and U4850 (N_4850,N_551,N_443);
or U4851 (N_4851,N_1606,N_2622);
nor U4852 (N_4852,N_2882,N_1614);
nor U4853 (N_4853,N_187,N_786);
and U4854 (N_4854,N_939,N_992);
nor U4855 (N_4855,N_872,N_1484);
nand U4856 (N_4856,N_2294,N_1147);
xor U4857 (N_4857,N_626,N_2135);
nand U4858 (N_4858,N_256,N_1084);
and U4859 (N_4859,N_2758,N_1616);
and U4860 (N_4860,N_1718,N_1291);
or U4861 (N_4861,N_2101,N_1998);
and U4862 (N_4862,N_2009,N_2638);
and U4863 (N_4863,N_764,N_2127);
nand U4864 (N_4864,N_478,N_362);
or U4865 (N_4865,N_2815,N_2878);
xnor U4866 (N_4866,N_382,N_433);
nand U4867 (N_4867,N_5,N_2385);
or U4868 (N_4868,N_1948,N_1754);
and U4869 (N_4869,N_214,N_2725);
nand U4870 (N_4870,N_505,N_710);
xor U4871 (N_4871,N_1916,N_885);
nand U4872 (N_4872,N_1295,N_1022);
or U4873 (N_4873,N_581,N_2814);
xor U4874 (N_4874,N_2924,N_238);
and U4875 (N_4875,N_2845,N_1338);
nand U4876 (N_4876,N_294,N_227);
nor U4877 (N_4877,N_594,N_460);
or U4878 (N_4878,N_341,N_1883);
nor U4879 (N_4879,N_1658,N_1012);
or U4880 (N_4880,N_2255,N_2968);
or U4881 (N_4881,N_2922,N_1461);
nor U4882 (N_4882,N_2562,N_1092);
or U4883 (N_4883,N_2533,N_1458);
xnor U4884 (N_4884,N_2793,N_2030);
xnor U4885 (N_4885,N_1544,N_1726);
and U4886 (N_4886,N_2093,N_1420);
or U4887 (N_4887,N_19,N_870);
nor U4888 (N_4888,N_2559,N_2373);
and U4889 (N_4889,N_873,N_2016);
nand U4890 (N_4890,N_2816,N_1855);
nand U4891 (N_4891,N_873,N_1224);
nand U4892 (N_4892,N_1887,N_1218);
nor U4893 (N_4893,N_2889,N_430);
nor U4894 (N_4894,N_2411,N_597);
and U4895 (N_4895,N_1704,N_1224);
xor U4896 (N_4896,N_391,N_2472);
or U4897 (N_4897,N_282,N_127);
nand U4898 (N_4898,N_797,N_2976);
or U4899 (N_4899,N_2434,N_2663);
and U4900 (N_4900,N_500,N_2269);
nand U4901 (N_4901,N_2862,N_153);
xor U4902 (N_4902,N_569,N_1023);
nor U4903 (N_4903,N_2357,N_2311);
xor U4904 (N_4904,N_553,N_174);
nor U4905 (N_4905,N_544,N_2282);
or U4906 (N_4906,N_125,N_2632);
nor U4907 (N_4907,N_414,N_2995);
and U4908 (N_4908,N_2378,N_1732);
nand U4909 (N_4909,N_1773,N_1835);
or U4910 (N_4910,N_2606,N_2379);
nor U4911 (N_4911,N_1746,N_83);
nand U4912 (N_4912,N_2601,N_526);
nand U4913 (N_4913,N_1541,N_2905);
nand U4914 (N_4914,N_2016,N_2469);
or U4915 (N_4915,N_2712,N_810);
nand U4916 (N_4916,N_221,N_1250);
or U4917 (N_4917,N_1744,N_2936);
nor U4918 (N_4918,N_143,N_12);
nand U4919 (N_4919,N_2901,N_1055);
nor U4920 (N_4920,N_595,N_401);
nand U4921 (N_4921,N_2151,N_2703);
xnor U4922 (N_4922,N_189,N_2374);
nand U4923 (N_4923,N_1860,N_1928);
nor U4924 (N_4924,N_1468,N_1099);
and U4925 (N_4925,N_2582,N_530);
xor U4926 (N_4926,N_2482,N_687);
or U4927 (N_4927,N_343,N_405);
nand U4928 (N_4928,N_2512,N_2345);
or U4929 (N_4929,N_38,N_2020);
nand U4930 (N_4930,N_2266,N_2430);
nand U4931 (N_4931,N_1858,N_1228);
nor U4932 (N_4932,N_678,N_839);
or U4933 (N_4933,N_2777,N_632);
and U4934 (N_4934,N_242,N_783);
xnor U4935 (N_4935,N_2646,N_2736);
or U4936 (N_4936,N_1678,N_1476);
nor U4937 (N_4937,N_429,N_2724);
nand U4938 (N_4938,N_2177,N_504);
nand U4939 (N_4939,N_1291,N_55);
or U4940 (N_4940,N_863,N_269);
nand U4941 (N_4941,N_2888,N_674);
and U4942 (N_4942,N_1514,N_189);
and U4943 (N_4943,N_529,N_285);
nor U4944 (N_4944,N_1554,N_1772);
xor U4945 (N_4945,N_1424,N_1242);
nand U4946 (N_4946,N_1849,N_2506);
and U4947 (N_4947,N_2860,N_2411);
and U4948 (N_4948,N_1404,N_1926);
or U4949 (N_4949,N_1841,N_2167);
nand U4950 (N_4950,N_2349,N_1762);
nand U4951 (N_4951,N_2219,N_2888);
nand U4952 (N_4952,N_1604,N_2685);
xor U4953 (N_4953,N_1702,N_1017);
and U4954 (N_4954,N_564,N_76);
and U4955 (N_4955,N_2414,N_478);
and U4956 (N_4956,N_2935,N_98);
nand U4957 (N_4957,N_2802,N_1959);
and U4958 (N_4958,N_1097,N_2581);
or U4959 (N_4959,N_203,N_1080);
nor U4960 (N_4960,N_1285,N_1242);
and U4961 (N_4961,N_487,N_1060);
nor U4962 (N_4962,N_2942,N_2645);
nand U4963 (N_4963,N_1849,N_2092);
xnor U4964 (N_4964,N_1614,N_788);
nand U4965 (N_4965,N_1483,N_823);
or U4966 (N_4966,N_1804,N_2621);
and U4967 (N_4967,N_273,N_677);
and U4968 (N_4968,N_2200,N_1585);
xnor U4969 (N_4969,N_2161,N_2129);
nand U4970 (N_4970,N_1015,N_958);
nand U4971 (N_4971,N_2799,N_2226);
and U4972 (N_4972,N_723,N_690);
and U4973 (N_4973,N_2680,N_2206);
and U4974 (N_4974,N_1231,N_1957);
or U4975 (N_4975,N_2717,N_1937);
and U4976 (N_4976,N_1174,N_1509);
and U4977 (N_4977,N_138,N_2445);
nand U4978 (N_4978,N_106,N_1513);
or U4979 (N_4979,N_2236,N_2962);
and U4980 (N_4980,N_1773,N_1770);
nor U4981 (N_4981,N_2494,N_2297);
or U4982 (N_4982,N_2509,N_1429);
nand U4983 (N_4983,N_1516,N_1582);
and U4984 (N_4984,N_2867,N_1996);
nor U4985 (N_4985,N_1285,N_1442);
or U4986 (N_4986,N_484,N_1680);
or U4987 (N_4987,N_2228,N_2706);
and U4988 (N_4988,N_2252,N_987);
xor U4989 (N_4989,N_811,N_152);
xor U4990 (N_4990,N_2693,N_1760);
xnor U4991 (N_4991,N_1574,N_843);
nor U4992 (N_4992,N_2476,N_1268);
nor U4993 (N_4993,N_2275,N_2988);
and U4994 (N_4994,N_2618,N_2426);
nand U4995 (N_4995,N_2014,N_2265);
and U4996 (N_4996,N_864,N_1265);
or U4997 (N_4997,N_2223,N_1573);
or U4998 (N_4998,N_1747,N_1878);
and U4999 (N_4999,N_1872,N_2895);
xnor U5000 (N_5000,N_2431,N_1980);
nand U5001 (N_5001,N_1621,N_1600);
and U5002 (N_5002,N_347,N_170);
nand U5003 (N_5003,N_569,N_2368);
or U5004 (N_5004,N_1449,N_1831);
and U5005 (N_5005,N_1195,N_2844);
and U5006 (N_5006,N_1009,N_1071);
and U5007 (N_5007,N_1363,N_1261);
nor U5008 (N_5008,N_2405,N_1756);
and U5009 (N_5009,N_161,N_2603);
nand U5010 (N_5010,N_1998,N_1448);
or U5011 (N_5011,N_497,N_62);
xor U5012 (N_5012,N_1989,N_938);
nor U5013 (N_5013,N_2035,N_2726);
or U5014 (N_5014,N_1706,N_2411);
nand U5015 (N_5015,N_2875,N_847);
xor U5016 (N_5016,N_291,N_2579);
nand U5017 (N_5017,N_2287,N_2439);
or U5018 (N_5018,N_1201,N_2831);
nor U5019 (N_5019,N_1610,N_126);
nand U5020 (N_5020,N_1859,N_1389);
xnor U5021 (N_5021,N_902,N_1355);
and U5022 (N_5022,N_1693,N_2838);
or U5023 (N_5023,N_2682,N_2063);
and U5024 (N_5024,N_1422,N_689);
or U5025 (N_5025,N_2340,N_1815);
nor U5026 (N_5026,N_2258,N_857);
nor U5027 (N_5027,N_2161,N_1743);
nor U5028 (N_5028,N_2286,N_1291);
or U5029 (N_5029,N_1850,N_286);
nand U5030 (N_5030,N_1616,N_1182);
nand U5031 (N_5031,N_1079,N_2582);
or U5032 (N_5032,N_1190,N_1244);
nor U5033 (N_5033,N_410,N_1791);
and U5034 (N_5034,N_1888,N_2613);
or U5035 (N_5035,N_1392,N_2277);
and U5036 (N_5036,N_519,N_1609);
xor U5037 (N_5037,N_1103,N_1782);
and U5038 (N_5038,N_1205,N_228);
nand U5039 (N_5039,N_165,N_1791);
or U5040 (N_5040,N_62,N_1872);
nor U5041 (N_5041,N_2095,N_1087);
xnor U5042 (N_5042,N_433,N_1660);
xnor U5043 (N_5043,N_1837,N_646);
xnor U5044 (N_5044,N_22,N_1286);
and U5045 (N_5045,N_2987,N_638);
and U5046 (N_5046,N_1393,N_2118);
and U5047 (N_5047,N_1843,N_1998);
or U5048 (N_5048,N_778,N_32);
nor U5049 (N_5049,N_1457,N_1320);
xor U5050 (N_5050,N_1054,N_2916);
xor U5051 (N_5051,N_2290,N_1584);
nor U5052 (N_5052,N_54,N_1581);
nand U5053 (N_5053,N_899,N_2644);
and U5054 (N_5054,N_1133,N_1490);
nor U5055 (N_5055,N_1684,N_1179);
nor U5056 (N_5056,N_505,N_2621);
and U5057 (N_5057,N_2565,N_318);
nand U5058 (N_5058,N_2400,N_920);
nor U5059 (N_5059,N_278,N_1109);
and U5060 (N_5060,N_1750,N_1834);
and U5061 (N_5061,N_676,N_1926);
nand U5062 (N_5062,N_1360,N_2724);
nand U5063 (N_5063,N_1030,N_660);
nand U5064 (N_5064,N_2055,N_2510);
and U5065 (N_5065,N_1282,N_1564);
nor U5066 (N_5066,N_1676,N_548);
nand U5067 (N_5067,N_497,N_1017);
and U5068 (N_5068,N_1434,N_1042);
or U5069 (N_5069,N_1493,N_1988);
or U5070 (N_5070,N_2396,N_258);
or U5071 (N_5071,N_2652,N_1411);
and U5072 (N_5072,N_1557,N_2642);
or U5073 (N_5073,N_1464,N_2457);
nand U5074 (N_5074,N_2949,N_1773);
or U5075 (N_5075,N_609,N_2092);
or U5076 (N_5076,N_585,N_694);
nor U5077 (N_5077,N_1785,N_2368);
nor U5078 (N_5078,N_114,N_1372);
or U5079 (N_5079,N_2731,N_2237);
or U5080 (N_5080,N_2641,N_292);
nor U5081 (N_5081,N_2524,N_664);
nor U5082 (N_5082,N_2317,N_320);
and U5083 (N_5083,N_1251,N_2531);
nor U5084 (N_5084,N_1971,N_438);
and U5085 (N_5085,N_1344,N_577);
nor U5086 (N_5086,N_395,N_911);
and U5087 (N_5087,N_1012,N_2731);
and U5088 (N_5088,N_2967,N_1662);
and U5089 (N_5089,N_590,N_1237);
and U5090 (N_5090,N_2745,N_1954);
nor U5091 (N_5091,N_1925,N_2501);
nand U5092 (N_5092,N_1923,N_283);
or U5093 (N_5093,N_2255,N_1055);
and U5094 (N_5094,N_436,N_99);
or U5095 (N_5095,N_277,N_1433);
nand U5096 (N_5096,N_2234,N_2049);
or U5097 (N_5097,N_1037,N_517);
nand U5098 (N_5098,N_1379,N_1859);
and U5099 (N_5099,N_2377,N_54);
nand U5100 (N_5100,N_484,N_1588);
nor U5101 (N_5101,N_2393,N_941);
nand U5102 (N_5102,N_2677,N_556);
or U5103 (N_5103,N_1374,N_1160);
xnor U5104 (N_5104,N_632,N_1119);
nand U5105 (N_5105,N_2512,N_1495);
and U5106 (N_5106,N_2861,N_1182);
and U5107 (N_5107,N_71,N_882);
and U5108 (N_5108,N_1837,N_1644);
and U5109 (N_5109,N_1965,N_130);
nor U5110 (N_5110,N_2002,N_56);
nor U5111 (N_5111,N_2995,N_692);
xnor U5112 (N_5112,N_459,N_449);
and U5113 (N_5113,N_2537,N_2175);
or U5114 (N_5114,N_2701,N_563);
nor U5115 (N_5115,N_2123,N_1544);
xor U5116 (N_5116,N_1948,N_1663);
nand U5117 (N_5117,N_1409,N_1453);
xor U5118 (N_5118,N_1533,N_1138);
nand U5119 (N_5119,N_1609,N_304);
or U5120 (N_5120,N_1559,N_263);
and U5121 (N_5121,N_469,N_740);
and U5122 (N_5122,N_1017,N_561);
xnor U5123 (N_5123,N_2953,N_1507);
or U5124 (N_5124,N_1171,N_671);
or U5125 (N_5125,N_715,N_1623);
or U5126 (N_5126,N_1497,N_741);
and U5127 (N_5127,N_1233,N_2547);
nand U5128 (N_5128,N_1995,N_847);
and U5129 (N_5129,N_2206,N_1374);
and U5130 (N_5130,N_1305,N_1028);
and U5131 (N_5131,N_122,N_1341);
nor U5132 (N_5132,N_955,N_1260);
nand U5133 (N_5133,N_2221,N_2565);
xnor U5134 (N_5134,N_114,N_2575);
or U5135 (N_5135,N_572,N_2572);
and U5136 (N_5136,N_2247,N_1073);
nor U5137 (N_5137,N_222,N_1289);
and U5138 (N_5138,N_2968,N_819);
and U5139 (N_5139,N_1794,N_1409);
and U5140 (N_5140,N_551,N_1299);
nand U5141 (N_5141,N_951,N_1903);
and U5142 (N_5142,N_1823,N_1579);
nand U5143 (N_5143,N_2059,N_965);
nand U5144 (N_5144,N_1361,N_2576);
nand U5145 (N_5145,N_1244,N_1817);
nor U5146 (N_5146,N_1250,N_1363);
and U5147 (N_5147,N_1473,N_911);
and U5148 (N_5148,N_131,N_944);
and U5149 (N_5149,N_2762,N_1335);
xor U5150 (N_5150,N_640,N_559);
nor U5151 (N_5151,N_1051,N_1042);
or U5152 (N_5152,N_2263,N_1004);
nand U5153 (N_5153,N_215,N_2407);
or U5154 (N_5154,N_1492,N_2488);
nor U5155 (N_5155,N_745,N_1165);
nand U5156 (N_5156,N_1523,N_2450);
nor U5157 (N_5157,N_2451,N_2979);
nor U5158 (N_5158,N_2497,N_44);
or U5159 (N_5159,N_119,N_1038);
or U5160 (N_5160,N_965,N_1976);
and U5161 (N_5161,N_493,N_1861);
or U5162 (N_5162,N_2585,N_2226);
and U5163 (N_5163,N_935,N_496);
nor U5164 (N_5164,N_1309,N_1332);
nor U5165 (N_5165,N_1514,N_227);
and U5166 (N_5166,N_612,N_2195);
and U5167 (N_5167,N_1233,N_1437);
xor U5168 (N_5168,N_880,N_2137);
nor U5169 (N_5169,N_2141,N_2192);
or U5170 (N_5170,N_2139,N_1717);
or U5171 (N_5171,N_14,N_2291);
xnor U5172 (N_5172,N_218,N_2979);
or U5173 (N_5173,N_2237,N_990);
xor U5174 (N_5174,N_885,N_2928);
nand U5175 (N_5175,N_1505,N_303);
xnor U5176 (N_5176,N_1864,N_1183);
nor U5177 (N_5177,N_1699,N_865);
or U5178 (N_5178,N_1241,N_1841);
xor U5179 (N_5179,N_2335,N_154);
or U5180 (N_5180,N_412,N_1038);
or U5181 (N_5181,N_1924,N_1098);
or U5182 (N_5182,N_1740,N_582);
and U5183 (N_5183,N_49,N_549);
nand U5184 (N_5184,N_461,N_2889);
and U5185 (N_5185,N_1174,N_594);
or U5186 (N_5186,N_2635,N_1011);
nand U5187 (N_5187,N_1238,N_1447);
nand U5188 (N_5188,N_735,N_2814);
nor U5189 (N_5189,N_1639,N_1427);
xnor U5190 (N_5190,N_2479,N_568);
or U5191 (N_5191,N_2625,N_1398);
or U5192 (N_5192,N_970,N_2511);
xor U5193 (N_5193,N_1571,N_1064);
nand U5194 (N_5194,N_2207,N_1925);
and U5195 (N_5195,N_2264,N_1978);
and U5196 (N_5196,N_334,N_1927);
or U5197 (N_5197,N_1827,N_1902);
nor U5198 (N_5198,N_1667,N_927);
nor U5199 (N_5199,N_1254,N_1485);
or U5200 (N_5200,N_640,N_1313);
and U5201 (N_5201,N_820,N_1289);
or U5202 (N_5202,N_2142,N_812);
and U5203 (N_5203,N_1834,N_1958);
nor U5204 (N_5204,N_2804,N_2820);
nor U5205 (N_5205,N_1108,N_1223);
nand U5206 (N_5206,N_2712,N_440);
and U5207 (N_5207,N_1557,N_673);
nand U5208 (N_5208,N_313,N_1853);
and U5209 (N_5209,N_2084,N_2660);
nand U5210 (N_5210,N_892,N_1822);
and U5211 (N_5211,N_92,N_2605);
nor U5212 (N_5212,N_985,N_1288);
nand U5213 (N_5213,N_606,N_174);
xor U5214 (N_5214,N_1431,N_2739);
or U5215 (N_5215,N_364,N_334);
nor U5216 (N_5216,N_1263,N_408);
or U5217 (N_5217,N_2842,N_1708);
and U5218 (N_5218,N_2756,N_2290);
nor U5219 (N_5219,N_1200,N_1797);
and U5220 (N_5220,N_1157,N_2503);
or U5221 (N_5221,N_1054,N_486);
nor U5222 (N_5222,N_1836,N_1655);
or U5223 (N_5223,N_396,N_654);
xor U5224 (N_5224,N_1641,N_1805);
and U5225 (N_5225,N_2894,N_1811);
nand U5226 (N_5226,N_2256,N_2772);
and U5227 (N_5227,N_1909,N_109);
or U5228 (N_5228,N_2904,N_431);
or U5229 (N_5229,N_525,N_2429);
nand U5230 (N_5230,N_1225,N_368);
or U5231 (N_5231,N_2613,N_533);
nor U5232 (N_5232,N_2589,N_2075);
nand U5233 (N_5233,N_547,N_2617);
nor U5234 (N_5234,N_1927,N_780);
and U5235 (N_5235,N_328,N_77);
nand U5236 (N_5236,N_1981,N_169);
nand U5237 (N_5237,N_2399,N_2087);
or U5238 (N_5238,N_2327,N_1519);
nand U5239 (N_5239,N_2450,N_654);
or U5240 (N_5240,N_573,N_1148);
nor U5241 (N_5241,N_2687,N_1153);
nand U5242 (N_5242,N_830,N_1121);
nand U5243 (N_5243,N_2141,N_2272);
and U5244 (N_5244,N_2960,N_572);
nor U5245 (N_5245,N_1441,N_1237);
xnor U5246 (N_5246,N_2427,N_1836);
nand U5247 (N_5247,N_520,N_242);
nor U5248 (N_5248,N_1765,N_2959);
nor U5249 (N_5249,N_1522,N_2115);
nand U5250 (N_5250,N_784,N_1681);
nor U5251 (N_5251,N_577,N_1195);
or U5252 (N_5252,N_2402,N_1233);
nand U5253 (N_5253,N_1202,N_2936);
nand U5254 (N_5254,N_350,N_1823);
nor U5255 (N_5255,N_1267,N_605);
nor U5256 (N_5256,N_1118,N_1790);
nor U5257 (N_5257,N_1670,N_1946);
nand U5258 (N_5258,N_2896,N_1422);
nand U5259 (N_5259,N_2172,N_747);
nand U5260 (N_5260,N_2625,N_1709);
and U5261 (N_5261,N_1368,N_66);
nand U5262 (N_5262,N_434,N_2457);
or U5263 (N_5263,N_694,N_385);
nor U5264 (N_5264,N_1875,N_2907);
nor U5265 (N_5265,N_2691,N_775);
or U5266 (N_5266,N_2633,N_2249);
or U5267 (N_5267,N_2124,N_2461);
and U5268 (N_5268,N_2258,N_1580);
and U5269 (N_5269,N_1017,N_601);
nand U5270 (N_5270,N_1926,N_1297);
nand U5271 (N_5271,N_416,N_2113);
or U5272 (N_5272,N_2492,N_1866);
nor U5273 (N_5273,N_662,N_510);
or U5274 (N_5274,N_2477,N_2061);
nand U5275 (N_5275,N_494,N_1016);
nand U5276 (N_5276,N_1982,N_896);
or U5277 (N_5277,N_786,N_206);
or U5278 (N_5278,N_1742,N_2932);
or U5279 (N_5279,N_2343,N_256);
nor U5280 (N_5280,N_2442,N_1247);
or U5281 (N_5281,N_797,N_1576);
and U5282 (N_5282,N_114,N_1516);
nor U5283 (N_5283,N_1913,N_2721);
nor U5284 (N_5284,N_428,N_1198);
and U5285 (N_5285,N_2727,N_129);
nand U5286 (N_5286,N_2735,N_1980);
nand U5287 (N_5287,N_1768,N_2825);
nor U5288 (N_5288,N_2198,N_301);
xnor U5289 (N_5289,N_228,N_806);
and U5290 (N_5290,N_2475,N_1662);
or U5291 (N_5291,N_1418,N_1803);
or U5292 (N_5292,N_664,N_781);
and U5293 (N_5293,N_2913,N_2221);
and U5294 (N_5294,N_2113,N_2265);
and U5295 (N_5295,N_2133,N_2020);
nor U5296 (N_5296,N_2802,N_1624);
nand U5297 (N_5297,N_307,N_568);
or U5298 (N_5298,N_82,N_971);
or U5299 (N_5299,N_2788,N_1369);
and U5300 (N_5300,N_1081,N_2795);
or U5301 (N_5301,N_1287,N_678);
nor U5302 (N_5302,N_832,N_2521);
xnor U5303 (N_5303,N_697,N_2241);
nor U5304 (N_5304,N_638,N_2289);
nand U5305 (N_5305,N_52,N_2030);
and U5306 (N_5306,N_1584,N_146);
and U5307 (N_5307,N_566,N_1026);
nor U5308 (N_5308,N_2696,N_576);
nand U5309 (N_5309,N_2148,N_2582);
xnor U5310 (N_5310,N_2292,N_37);
nor U5311 (N_5311,N_1526,N_652);
nand U5312 (N_5312,N_2601,N_1356);
and U5313 (N_5313,N_6,N_1838);
nor U5314 (N_5314,N_1531,N_1761);
or U5315 (N_5315,N_2448,N_1835);
and U5316 (N_5316,N_546,N_2742);
nand U5317 (N_5317,N_2331,N_1431);
nor U5318 (N_5318,N_834,N_1980);
nand U5319 (N_5319,N_1055,N_2447);
and U5320 (N_5320,N_881,N_1457);
or U5321 (N_5321,N_1384,N_2988);
nor U5322 (N_5322,N_652,N_1047);
and U5323 (N_5323,N_983,N_899);
nand U5324 (N_5324,N_1549,N_2482);
nor U5325 (N_5325,N_1958,N_740);
nand U5326 (N_5326,N_2794,N_180);
nor U5327 (N_5327,N_2625,N_1841);
or U5328 (N_5328,N_1298,N_947);
and U5329 (N_5329,N_251,N_2906);
or U5330 (N_5330,N_2346,N_1669);
and U5331 (N_5331,N_2256,N_2620);
nand U5332 (N_5332,N_450,N_2020);
and U5333 (N_5333,N_1198,N_207);
nor U5334 (N_5334,N_1162,N_422);
nor U5335 (N_5335,N_68,N_1143);
nand U5336 (N_5336,N_711,N_623);
or U5337 (N_5337,N_2824,N_1587);
and U5338 (N_5338,N_2417,N_1058);
nand U5339 (N_5339,N_2149,N_1675);
nand U5340 (N_5340,N_1866,N_2173);
and U5341 (N_5341,N_2661,N_193);
and U5342 (N_5342,N_989,N_2644);
or U5343 (N_5343,N_217,N_1509);
xor U5344 (N_5344,N_2827,N_1749);
or U5345 (N_5345,N_681,N_2800);
or U5346 (N_5346,N_2349,N_1496);
nand U5347 (N_5347,N_1276,N_487);
nor U5348 (N_5348,N_1465,N_1093);
or U5349 (N_5349,N_1723,N_2303);
or U5350 (N_5350,N_1003,N_1767);
and U5351 (N_5351,N_360,N_2479);
nor U5352 (N_5352,N_1447,N_1398);
or U5353 (N_5353,N_134,N_144);
and U5354 (N_5354,N_13,N_1975);
or U5355 (N_5355,N_1653,N_2986);
xnor U5356 (N_5356,N_268,N_1403);
nor U5357 (N_5357,N_1113,N_2266);
nor U5358 (N_5358,N_980,N_995);
nand U5359 (N_5359,N_1279,N_2787);
nand U5360 (N_5360,N_929,N_1887);
nand U5361 (N_5361,N_2653,N_1766);
or U5362 (N_5362,N_2842,N_583);
nand U5363 (N_5363,N_1752,N_1829);
and U5364 (N_5364,N_736,N_1967);
nand U5365 (N_5365,N_1036,N_1840);
nand U5366 (N_5366,N_658,N_2400);
nand U5367 (N_5367,N_726,N_2242);
nand U5368 (N_5368,N_2742,N_348);
and U5369 (N_5369,N_807,N_2271);
or U5370 (N_5370,N_1319,N_1544);
nor U5371 (N_5371,N_2065,N_1384);
or U5372 (N_5372,N_89,N_2029);
or U5373 (N_5373,N_992,N_2385);
and U5374 (N_5374,N_755,N_195);
nand U5375 (N_5375,N_498,N_651);
and U5376 (N_5376,N_2212,N_1485);
xnor U5377 (N_5377,N_2711,N_2672);
and U5378 (N_5378,N_2738,N_1362);
xnor U5379 (N_5379,N_2026,N_23);
and U5380 (N_5380,N_1473,N_658);
xor U5381 (N_5381,N_1757,N_1200);
xnor U5382 (N_5382,N_2357,N_1649);
nor U5383 (N_5383,N_2894,N_1382);
nand U5384 (N_5384,N_959,N_924);
and U5385 (N_5385,N_953,N_2039);
and U5386 (N_5386,N_1692,N_170);
nor U5387 (N_5387,N_2269,N_317);
or U5388 (N_5388,N_346,N_2721);
nor U5389 (N_5389,N_1446,N_1311);
and U5390 (N_5390,N_2276,N_58);
nor U5391 (N_5391,N_2605,N_2837);
xnor U5392 (N_5392,N_1928,N_683);
nor U5393 (N_5393,N_677,N_2835);
nand U5394 (N_5394,N_1821,N_1354);
xnor U5395 (N_5395,N_1072,N_2463);
and U5396 (N_5396,N_1075,N_1407);
or U5397 (N_5397,N_416,N_690);
xnor U5398 (N_5398,N_497,N_2801);
nor U5399 (N_5399,N_2480,N_442);
or U5400 (N_5400,N_748,N_1941);
nor U5401 (N_5401,N_1595,N_1570);
nand U5402 (N_5402,N_2995,N_2993);
or U5403 (N_5403,N_2233,N_476);
and U5404 (N_5404,N_2560,N_2064);
or U5405 (N_5405,N_1922,N_459);
and U5406 (N_5406,N_2671,N_2347);
nand U5407 (N_5407,N_72,N_1225);
and U5408 (N_5408,N_2696,N_518);
and U5409 (N_5409,N_1652,N_2676);
nor U5410 (N_5410,N_2706,N_2499);
and U5411 (N_5411,N_2567,N_1469);
nand U5412 (N_5412,N_2821,N_2772);
nor U5413 (N_5413,N_541,N_1035);
and U5414 (N_5414,N_401,N_1746);
xor U5415 (N_5415,N_1226,N_40);
and U5416 (N_5416,N_378,N_170);
and U5417 (N_5417,N_1349,N_1354);
nor U5418 (N_5418,N_477,N_939);
and U5419 (N_5419,N_551,N_1567);
and U5420 (N_5420,N_1169,N_2350);
nand U5421 (N_5421,N_2982,N_640);
nand U5422 (N_5422,N_2301,N_673);
and U5423 (N_5423,N_2599,N_1255);
or U5424 (N_5424,N_69,N_2720);
nor U5425 (N_5425,N_765,N_181);
nand U5426 (N_5426,N_2157,N_549);
or U5427 (N_5427,N_2337,N_2901);
nor U5428 (N_5428,N_749,N_1399);
and U5429 (N_5429,N_2340,N_2257);
and U5430 (N_5430,N_50,N_1759);
nand U5431 (N_5431,N_1567,N_157);
and U5432 (N_5432,N_2140,N_770);
or U5433 (N_5433,N_597,N_903);
nand U5434 (N_5434,N_634,N_278);
or U5435 (N_5435,N_65,N_2591);
nand U5436 (N_5436,N_2970,N_966);
or U5437 (N_5437,N_2829,N_2800);
or U5438 (N_5438,N_1356,N_2592);
nor U5439 (N_5439,N_1912,N_1180);
nor U5440 (N_5440,N_2197,N_2019);
or U5441 (N_5441,N_2408,N_329);
nand U5442 (N_5442,N_2226,N_2409);
or U5443 (N_5443,N_2000,N_22);
xor U5444 (N_5444,N_351,N_1142);
or U5445 (N_5445,N_1843,N_1093);
or U5446 (N_5446,N_1880,N_2299);
nor U5447 (N_5447,N_133,N_1691);
and U5448 (N_5448,N_1215,N_1718);
xnor U5449 (N_5449,N_2281,N_2382);
nand U5450 (N_5450,N_2051,N_2831);
and U5451 (N_5451,N_2213,N_2568);
nor U5452 (N_5452,N_1828,N_1576);
nand U5453 (N_5453,N_1485,N_1029);
xnor U5454 (N_5454,N_803,N_1395);
nand U5455 (N_5455,N_1332,N_2174);
nand U5456 (N_5456,N_2474,N_2712);
nor U5457 (N_5457,N_2316,N_424);
xor U5458 (N_5458,N_408,N_1458);
nor U5459 (N_5459,N_244,N_2877);
and U5460 (N_5460,N_1762,N_64);
xor U5461 (N_5461,N_625,N_980);
nand U5462 (N_5462,N_2595,N_1133);
and U5463 (N_5463,N_2389,N_768);
and U5464 (N_5464,N_2172,N_1447);
and U5465 (N_5465,N_140,N_244);
or U5466 (N_5466,N_98,N_1693);
nor U5467 (N_5467,N_2444,N_475);
and U5468 (N_5468,N_442,N_1259);
xor U5469 (N_5469,N_2235,N_2606);
xor U5470 (N_5470,N_1601,N_1286);
or U5471 (N_5471,N_2055,N_1160);
nor U5472 (N_5472,N_2290,N_2352);
xor U5473 (N_5473,N_180,N_256);
and U5474 (N_5474,N_2325,N_750);
or U5475 (N_5475,N_2511,N_156);
nor U5476 (N_5476,N_2276,N_2553);
nand U5477 (N_5477,N_1964,N_149);
and U5478 (N_5478,N_694,N_1176);
or U5479 (N_5479,N_2177,N_1663);
and U5480 (N_5480,N_786,N_1399);
or U5481 (N_5481,N_2797,N_970);
nand U5482 (N_5482,N_2702,N_558);
nor U5483 (N_5483,N_801,N_2156);
and U5484 (N_5484,N_129,N_79);
nor U5485 (N_5485,N_2075,N_1534);
nor U5486 (N_5486,N_1409,N_819);
xor U5487 (N_5487,N_719,N_1635);
or U5488 (N_5488,N_1459,N_95);
and U5489 (N_5489,N_1006,N_1907);
and U5490 (N_5490,N_1757,N_2027);
xor U5491 (N_5491,N_1285,N_217);
nand U5492 (N_5492,N_456,N_508);
and U5493 (N_5493,N_261,N_253);
nor U5494 (N_5494,N_547,N_1665);
nor U5495 (N_5495,N_1761,N_2244);
nand U5496 (N_5496,N_2030,N_1928);
and U5497 (N_5497,N_194,N_474);
and U5498 (N_5498,N_120,N_1040);
nor U5499 (N_5499,N_2837,N_2851);
or U5500 (N_5500,N_2111,N_596);
nand U5501 (N_5501,N_1887,N_1644);
xnor U5502 (N_5502,N_975,N_2189);
nand U5503 (N_5503,N_1188,N_2964);
nor U5504 (N_5504,N_1844,N_2008);
xor U5505 (N_5505,N_2753,N_1914);
nor U5506 (N_5506,N_1263,N_1848);
nand U5507 (N_5507,N_1044,N_1240);
or U5508 (N_5508,N_366,N_2405);
or U5509 (N_5509,N_2703,N_766);
and U5510 (N_5510,N_387,N_1502);
nand U5511 (N_5511,N_100,N_2190);
and U5512 (N_5512,N_1253,N_2692);
or U5513 (N_5513,N_2684,N_1654);
and U5514 (N_5514,N_1075,N_1159);
nor U5515 (N_5515,N_1377,N_495);
and U5516 (N_5516,N_2269,N_330);
or U5517 (N_5517,N_2385,N_1288);
nor U5518 (N_5518,N_1170,N_527);
nand U5519 (N_5519,N_2108,N_973);
nand U5520 (N_5520,N_1500,N_2454);
and U5521 (N_5521,N_596,N_853);
nor U5522 (N_5522,N_1049,N_2637);
or U5523 (N_5523,N_820,N_627);
and U5524 (N_5524,N_2214,N_2625);
xnor U5525 (N_5525,N_2107,N_1920);
nand U5526 (N_5526,N_1168,N_1420);
nor U5527 (N_5527,N_2339,N_2025);
and U5528 (N_5528,N_1861,N_210);
nand U5529 (N_5529,N_52,N_290);
or U5530 (N_5530,N_2816,N_1560);
or U5531 (N_5531,N_2015,N_1197);
nand U5532 (N_5532,N_2865,N_1998);
nand U5533 (N_5533,N_968,N_327);
xor U5534 (N_5534,N_2474,N_2848);
nor U5535 (N_5535,N_2853,N_144);
and U5536 (N_5536,N_1003,N_450);
nand U5537 (N_5537,N_2415,N_21);
nor U5538 (N_5538,N_2310,N_1117);
nand U5539 (N_5539,N_319,N_1821);
and U5540 (N_5540,N_854,N_2232);
nor U5541 (N_5541,N_356,N_1566);
nor U5542 (N_5542,N_974,N_1296);
and U5543 (N_5543,N_1914,N_769);
and U5544 (N_5544,N_243,N_253);
and U5545 (N_5545,N_906,N_2529);
and U5546 (N_5546,N_2072,N_379);
nor U5547 (N_5547,N_1323,N_253);
nor U5548 (N_5548,N_2436,N_722);
xor U5549 (N_5549,N_1842,N_2901);
or U5550 (N_5550,N_450,N_1912);
or U5551 (N_5551,N_2445,N_1274);
or U5552 (N_5552,N_1730,N_1161);
nor U5553 (N_5553,N_1774,N_2832);
or U5554 (N_5554,N_775,N_2321);
nand U5555 (N_5555,N_2220,N_214);
nand U5556 (N_5556,N_1854,N_2829);
or U5557 (N_5557,N_932,N_2172);
nand U5558 (N_5558,N_435,N_1830);
or U5559 (N_5559,N_1065,N_1895);
nor U5560 (N_5560,N_658,N_2307);
or U5561 (N_5561,N_2151,N_103);
and U5562 (N_5562,N_2519,N_183);
nand U5563 (N_5563,N_1095,N_278);
nor U5564 (N_5564,N_368,N_1218);
xnor U5565 (N_5565,N_2472,N_2831);
and U5566 (N_5566,N_1219,N_1212);
nor U5567 (N_5567,N_168,N_1794);
nor U5568 (N_5568,N_139,N_2241);
nand U5569 (N_5569,N_600,N_238);
and U5570 (N_5570,N_2046,N_386);
xor U5571 (N_5571,N_810,N_205);
or U5572 (N_5572,N_1609,N_2848);
or U5573 (N_5573,N_2029,N_1227);
xor U5574 (N_5574,N_1321,N_2967);
nor U5575 (N_5575,N_2829,N_1431);
and U5576 (N_5576,N_2182,N_1210);
and U5577 (N_5577,N_828,N_2694);
nor U5578 (N_5578,N_2740,N_821);
nand U5579 (N_5579,N_309,N_2104);
nand U5580 (N_5580,N_1202,N_1953);
nand U5581 (N_5581,N_2441,N_1639);
nor U5582 (N_5582,N_2503,N_1277);
and U5583 (N_5583,N_2401,N_150);
or U5584 (N_5584,N_412,N_2199);
nor U5585 (N_5585,N_764,N_2510);
and U5586 (N_5586,N_1367,N_1060);
xor U5587 (N_5587,N_2694,N_923);
or U5588 (N_5588,N_1567,N_1744);
nand U5589 (N_5589,N_1644,N_1089);
or U5590 (N_5590,N_1763,N_1704);
nor U5591 (N_5591,N_8,N_744);
or U5592 (N_5592,N_912,N_2307);
and U5593 (N_5593,N_689,N_2639);
and U5594 (N_5594,N_1682,N_314);
or U5595 (N_5595,N_449,N_2461);
or U5596 (N_5596,N_2330,N_376);
nand U5597 (N_5597,N_1723,N_1346);
nand U5598 (N_5598,N_886,N_2923);
nor U5599 (N_5599,N_766,N_750);
or U5600 (N_5600,N_2256,N_2111);
xor U5601 (N_5601,N_1110,N_1385);
nor U5602 (N_5602,N_1587,N_1837);
and U5603 (N_5603,N_694,N_1007);
nand U5604 (N_5604,N_1942,N_161);
or U5605 (N_5605,N_636,N_2434);
or U5606 (N_5606,N_1690,N_2839);
and U5607 (N_5607,N_173,N_1736);
or U5608 (N_5608,N_2869,N_1750);
and U5609 (N_5609,N_414,N_334);
or U5610 (N_5610,N_1270,N_391);
or U5611 (N_5611,N_565,N_343);
nand U5612 (N_5612,N_135,N_1433);
nor U5613 (N_5613,N_1694,N_117);
xnor U5614 (N_5614,N_2140,N_338);
and U5615 (N_5615,N_1314,N_511);
nor U5616 (N_5616,N_229,N_435);
nor U5617 (N_5617,N_1920,N_548);
nand U5618 (N_5618,N_2923,N_37);
nand U5619 (N_5619,N_2009,N_1029);
and U5620 (N_5620,N_1400,N_67);
nand U5621 (N_5621,N_2502,N_2466);
nor U5622 (N_5622,N_2699,N_1477);
or U5623 (N_5623,N_1843,N_2265);
nand U5624 (N_5624,N_432,N_2760);
and U5625 (N_5625,N_1713,N_113);
or U5626 (N_5626,N_484,N_25);
nor U5627 (N_5627,N_1414,N_2525);
or U5628 (N_5628,N_393,N_1498);
xor U5629 (N_5629,N_55,N_1168);
or U5630 (N_5630,N_1333,N_929);
or U5631 (N_5631,N_11,N_1902);
nor U5632 (N_5632,N_2307,N_231);
nand U5633 (N_5633,N_1488,N_1424);
and U5634 (N_5634,N_2694,N_826);
nand U5635 (N_5635,N_216,N_2936);
and U5636 (N_5636,N_346,N_1406);
nand U5637 (N_5637,N_2609,N_1142);
nand U5638 (N_5638,N_2504,N_259);
nor U5639 (N_5639,N_450,N_2230);
or U5640 (N_5640,N_2491,N_859);
nand U5641 (N_5641,N_1026,N_2904);
nand U5642 (N_5642,N_1706,N_75);
xor U5643 (N_5643,N_909,N_1928);
nand U5644 (N_5644,N_2801,N_868);
nor U5645 (N_5645,N_199,N_2561);
nor U5646 (N_5646,N_705,N_1638);
xor U5647 (N_5647,N_1224,N_1298);
nor U5648 (N_5648,N_1042,N_2926);
and U5649 (N_5649,N_2986,N_1136);
nand U5650 (N_5650,N_2207,N_2426);
nand U5651 (N_5651,N_2176,N_1410);
or U5652 (N_5652,N_1594,N_784);
nand U5653 (N_5653,N_2256,N_2375);
xor U5654 (N_5654,N_1428,N_1552);
or U5655 (N_5655,N_1176,N_2048);
nand U5656 (N_5656,N_2098,N_2859);
xor U5657 (N_5657,N_212,N_1231);
or U5658 (N_5658,N_1242,N_795);
or U5659 (N_5659,N_2272,N_535);
or U5660 (N_5660,N_76,N_2582);
or U5661 (N_5661,N_594,N_950);
nor U5662 (N_5662,N_2479,N_2859);
xnor U5663 (N_5663,N_2335,N_2367);
or U5664 (N_5664,N_580,N_155);
or U5665 (N_5665,N_332,N_2956);
nor U5666 (N_5666,N_32,N_1243);
or U5667 (N_5667,N_2393,N_82);
nor U5668 (N_5668,N_1591,N_1622);
and U5669 (N_5669,N_15,N_1227);
nor U5670 (N_5670,N_2994,N_2943);
nor U5671 (N_5671,N_216,N_694);
nor U5672 (N_5672,N_2400,N_2596);
and U5673 (N_5673,N_513,N_2764);
or U5674 (N_5674,N_1674,N_1577);
nand U5675 (N_5675,N_2345,N_734);
nand U5676 (N_5676,N_2128,N_983);
xnor U5677 (N_5677,N_1020,N_1719);
or U5678 (N_5678,N_1574,N_2570);
nor U5679 (N_5679,N_650,N_2925);
nor U5680 (N_5680,N_715,N_2162);
nor U5681 (N_5681,N_1321,N_355);
or U5682 (N_5682,N_1206,N_987);
nand U5683 (N_5683,N_2801,N_354);
or U5684 (N_5684,N_1069,N_62);
or U5685 (N_5685,N_2356,N_1477);
nand U5686 (N_5686,N_174,N_1071);
and U5687 (N_5687,N_881,N_927);
xor U5688 (N_5688,N_2807,N_903);
xnor U5689 (N_5689,N_2029,N_2683);
nor U5690 (N_5690,N_1002,N_2243);
nand U5691 (N_5691,N_2220,N_2702);
or U5692 (N_5692,N_2179,N_1837);
and U5693 (N_5693,N_1433,N_2666);
nor U5694 (N_5694,N_2088,N_2076);
xnor U5695 (N_5695,N_863,N_1659);
or U5696 (N_5696,N_79,N_448);
nor U5697 (N_5697,N_2999,N_2207);
or U5698 (N_5698,N_897,N_794);
or U5699 (N_5699,N_1072,N_671);
or U5700 (N_5700,N_52,N_1247);
nand U5701 (N_5701,N_1395,N_353);
and U5702 (N_5702,N_1690,N_1818);
or U5703 (N_5703,N_1339,N_1060);
and U5704 (N_5704,N_118,N_2785);
or U5705 (N_5705,N_407,N_133);
nor U5706 (N_5706,N_1995,N_16);
xor U5707 (N_5707,N_2499,N_1228);
nor U5708 (N_5708,N_2782,N_1637);
nor U5709 (N_5709,N_608,N_754);
and U5710 (N_5710,N_1703,N_985);
nor U5711 (N_5711,N_628,N_825);
and U5712 (N_5712,N_2153,N_481);
or U5713 (N_5713,N_1534,N_652);
nor U5714 (N_5714,N_2549,N_673);
nor U5715 (N_5715,N_184,N_444);
nor U5716 (N_5716,N_1984,N_1425);
and U5717 (N_5717,N_1506,N_1427);
nand U5718 (N_5718,N_207,N_1075);
xor U5719 (N_5719,N_1623,N_1697);
or U5720 (N_5720,N_191,N_2835);
and U5721 (N_5721,N_270,N_1137);
xor U5722 (N_5722,N_1307,N_2448);
and U5723 (N_5723,N_843,N_547);
nor U5724 (N_5724,N_982,N_1060);
and U5725 (N_5725,N_301,N_205);
nor U5726 (N_5726,N_365,N_1173);
and U5727 (N_5727,N_717,N_11);
and U5728 (N_5728,N_804,N_2461);
xor U5729 (N_5729,N_2836,N_24);
nand U5730 (N_5730,N_108,N_509);
nand U5731 (N_5731,N_2224,N_91);
nand U5732 (N_5732,N_2493,N_1828);
and U5733 (N_5733,N_2130,N_834);
and U5734 (N_5734,N_1369,N_715);
or U5735 (N_5735,N_378,N_1421);
nand U5736 (N_5736,N_118,N_1345);
nand U5737 (N_5737,N_985,N_2061);
xnor U5738 (N_5738,N_614,N_2626);
and U5739 (N_5739,N_1034,N_2550);
nor U5740 (N_5740,N_2687,N_2538);
or U5741 (N_5741,N_1784,N_979);
nand U5742 (N_5742,N_1006,N_2659);
nand U5743 (N_5743,N_2554,N_1259);
nor U5744 (N_5744,N_2606,N_2292);
and U5745 (N_5745,N_1114,N_171);
or U5746 (N_5746,N_147,N_849);
and U5747 (N_5747,N_1191,N_2326);
nand U5748 (N_5748,N_2156,N_1146);
nand U5749 (N_5749,N_2138,N_603);
or U5750 (N_5750,N_2610,N_2487);
nand U5751 (N_5751,N_2854,N_1407);
or U5752 (N_5752,N_460,N_2270);
nor U5753 (N_5753,N_343,N_2502);
and U5754 (N_5754,N_2589,N_63);
or U5755 (N_5755,N_1771,N_2864);
nand U5756 (N_5756,N_2489,N_2308);
xor U5757 (N_5757,N_2164,N_36);
nand U5758 (N_5758,N_1414,N_255);
nand U5759 (N_5759,N_1797,N_2841);
or U5760 (N_5760,N_383,N_117);
and U5761 (N_5761,N_1204,N_1209);
or U5762 (N_5762,N_2733,N_2422);
and U5763 (N_5763,N_1498,N_2871);
nor U5764 (N_5764,N_797,N_114);
xnor U5765 (N_5765,N_1126,N_1081);
or U5766 (N_5766,N_1249,N_2493);
and U5767 (N_5767,N_207,N_1789);
nand U5768 (N_5768,N_829,N_2786);
or U5769 (N_5769,N_32,N_907);
and U5770 (N_5770,N_2701,N_766);
and U5771 (N_5771,N_303,N_1654);
or U5772 (N_5772,N_1932,N_1320);
or U5773 (N_5773,N_14,N_2638);
or U5774 (N_5774,N_1917,N_1326);
and U5775 (N_5775,N_1898,N_1070);
or U5776 (N_5776,N_1623,N_2477);
and U5777 (N_5777,N_1794,N_2636);
nand U5778 (N_5778,N_505,N_902);
nand U5779 (N_5779,N_2078,N_74);
or U5780 (N_5780,N_346,N_1401);
nand U5781 (N_5781,N_388,N_999);
nand U5782 (N_5782,N_714,N_2566);
nand U5783 (N_5783,N_3,N_1583);
or U5784 (N_5784,N_763,N_1833);
nand U5785 (N_5785,N_1772,N_1802);
xor U5786 (N_5786,N_2229,N_2444);
nor U5787 (N_5787,N_953,N_1499);
or U5788 (N_5788,N_2815,N_525);
nand U5789 (N_5789,N_2769,N_2172);
xor U5790 (N_5790,N_472,N_2526);
nor U5791 (N_5791,N_1763,N_2418);
nor U5792 (N_5792,N_2034,N_2977);
or U5793 (N_5793,N_940,N_1178);
nor U5794 (N_5794,N_2668,N_2248);
xnor U5795 (N_5795,N_1330,N_1639);
nor U5796 (N_5796,N_819,N_1893);
and U5797 (N_5797,N_1643,N_2441);
and U5798 (N_5798,N_2180,N_359);
nand U5799 (N_5799,N_185,N_940);
nor U5800 (N_5800,N_965,N_2444);
nor U5801 (N_5801,N_480,N_1489);
nand U5802 (N_5802,N_1847,N_2969);
nor U5803 (N_5803,N_527,N_243);
nor U5804 (N_5804,N_867,N_2106);
and U5805 (N_5805,N_705,N_2039);
and U5806 (N_5806,N_350,N_67);
and U5807 (N_5807,N_303,N_2964);
and U5808 (N_5808,N_1123,N_2304);
and U5809 (N_5809,N_391,N_84);
nand U5810 (N_5810,N_1931,N_2206);
nand U5811 (N_5811,N_2209,N_2798);
and U5812 (N_5812,N_2982,N_278);
or U5813 (N_5813,N_1221,N_2999);
or U5814 (N_5814,N_412,N_2728);
nor U5815 (N_5815,N_1940,N_84);
or U5816 (N_5816,N_2125,N_128);
or U5817 (N_5817,N_384,N_2231);
nand U5818 (N_5818,N_460,N_2094);
nand U5819 (N_5819,N_1948,N_142);
or U5820 (N_5820,N_2403,N_1531);
and U5821 (N_5821,N_868,N_2659);
nor U5822 (N_5822,N_2208,N_2008);
and U5823 (N_5823,N_345,N_2572);
nand U5824 (N_5824,N_1783,N_456);
nand U5825 (N_5825,N_2121,N_1461);
nand U5826 (N_5826,N_73,N_199);
nor U5827 (N_5827,N_1482,N_1122);
xor U5828 (N_5828,N_2576,N_1802);
or U5829 (N_5829,N_2115,N_2565);
or U5830 (N_5830,N_335,N_2291);
or U5831 (N_5831,N_2494,N_2537);
nand U5832 (N_5832,N_451,N_438);
and U5833 (N_5833,N_2962,N_1571);
and U5834 (N_5834,N_821,N_2209);
nand U5835 (N_5835,N_98,N_37);
xor U5836 (N_5836,N_576,N_1346);
xor U5837 (N_5837,N_1174,N_772);
or U5838 (N_5838,N_1488,N_1940);
and U5839 (N_5839,N_2432,N_546);
xor U5840 (N_5840,N_2384,N_438);
nand U5841 (N_5841,N_1450,N_2818);
nand U5842 (N_5842,N_614,N_923);
nor U5843 (N_5843,N_1897,N_2112);
nor U5844 (N_5844,N_2429,N_461);
or U5845 (N_5845,N_395,N_964);
nand U5846 (N_5846,N_2202,N_155);
nor U5847 (N_5847,N_2429,N_2076);
nor U5848 (N_5848,N_2873,N_1938);
nand U5849 (N_5849,N_1204,N_234);
nand U5850 (N_5850,N_769,N_2451);
and U5851 (N_5851,N_958,N_2925);
and U5852 (N_5852,N_326,N_2668);
nand U5853 (N_5853,N_1302,N_91);
xor U5854 (N_5854,N_45,N_2808);
xor U5855 (N_5855,N_1974,N_1861);
xnor U5856 (N_5856,N_388,N_1833);
nor U5857 (N_5857,N_602,N_672);
nand U5858 (N_5858,N_473,N_1178);
nor U5859 (N_5859,N_2976,N_498);
nor U5860 (N_5860,N_2427,N_2949);
and U5861 (N_5861,N_1438,N_1235);
nand U5862 (N_5862,N_1220,N_2600);
or U5863 (N_5863,N_1632,N_2863);
nor U5864 (N_5864,N_2292,N_224);
and U5865 (N_5865,N_2024,N_2866);
or U5866 (N_5866,N_1720,N_1540);
and U5867 (N_5867,N_2075,N_2240);
or U5868 (N_5868,N_2919,N_598);
nor U5869 (N_5869,N_2856,N_2607);
or U5870 (N_5870,N_1776,N_2442);
nor U5871 (N_5871,N_838,N_2601);
or U5872 (N_5872,N_1296,N_1277);
and U5873 (N_5873,N_2723,N_1760);
nand U5874 (N_5874,N_2411,N_1025);
nor U5875 (N_5875,N_1063,N_2925);
nand U5876 (N_5876,N_1221,N_2565);
or U5877 (N_5877,N_1960,N_2367);
or U5878 (N_5878,N_2132,N_2402);
or U5879 (N_5879,N_154,N_1791);
nand U5880 (N_5880,N_2482,N_741);
nand U5881 (N_5881,N_462,N_2355);
and U5882 (N_5882,N_1372,N_684);
xor U5883 (N_5883,N_1389,N_112);
nor U5884 (N_5884,N_1293,N_2213);
nand U5885 (N_5885,N_1638,N_633);
nand U5886 (N_5886,N_2999,N_2869);
nor U5887 (N_5887,N_2456,N_452);
xor U5888 (N_5888,N_136,N_1003);
and U5889 (N_5889,N_2427,N_113);
nor U5890 (N_5890,N_1962,N_2359);
and U5891 (N_5891,N_1063,N_103);
nand U5892 (N_5892,N_1665,N_1352);
nand U5893 (N_5893,N_133,N_1065);
nor U5894 (N_5894,N_2706,N_1766);
or U5895 (N_5895,N_2589,N_2692);
or U5896 (N_5896,N_2383,N_2724);
or U5897 (N_5897,N_2628,N_336);
nand U5898 (N_5898,N_1289,N_1277);
and U5899 (N_5899,N_2093,N_1652);
xnor U5900 (N_5900,N_1748,N_1168);
and U5901 (N_5901,N_2258,N_1950);
nor U5902 (N_5902,N_1550,N_1777);
and U5903 (N_5903,N_2496,N_402);
and U5904 (N_5904,N_51,N_485);
and U5905 (N_5905,N_619,N_2790);
nor U5906 (N_5906,N_2308,N_2901);
nand U5907 (N_5907,N_2245,N_232);
nand U5908 (N_5908,N_2279,N_2889);
and U5909 (N_5909,N_373,N_2463);
or U5910 (N_5910,N_2163,N_264);
nor U5911 (N_5911,N_879,N_1255);
and U5912 (N_5912,N_906,N_1566);
or U5913 (N_5913,N_1104,N_2653);
nor U5914 (N_5914,N_2972,N_1551);
nand U5915 (N_5915,N_2396,N_2681);
nor U5916 (N_5916,N_1716,N_690);
nor U5917 (N_5917,N_2394,N_1497);
nor U5918 (N_5918,N_2532,N_2055);
nor U5919 (N_5919,N_2395,N_137);
nand U5920 (N_5920,N_435,N_1316);
or U5921 (N_5921,N_80,N_493);
or U5922 (N_5922,N_2192,N_310);
and U5923 (N_5923,N_1149,N_541);
or U5924 (N_5924,N_1911,N_2295);
or U5925 (N_5925,N_1845,N_2217);
nand U5926 (N_5926,N_1852,N_74);
or U5927 (N_5927,N_77,N_140);
or U5928 (N_5928,N_2584,N_937);
nor U5929 (N_5929,N_442,N_2530);
or U5930 (N_5930,N_2876,N_1624);
nand U5931 (N_5931,N_1929,N_1427);
or U5932 (N_5932,N_1110,N_1826);
nand U5933 (N_5933,N_2502,N_1728);
or U5934 (N_5934,N_92,N_2937);
nand U5935 (N_5935,N_426,N_367);
or U5936 (N_5936,N_114,N_315);
nor U5937 (N_5937,N_2971,N_1230);
or U5938 (N_5938,N_1792,N_1511);
nand U5939 (N_5939,N_1043,N_1920);
and U5940 (N_5940,N_2894,N_2092);
nor U5941 (N_5941,N_80,N_2786);
or U5942 (N_5942,N_252,N_884);
nand U5943 (N_5943,N_2890,N_1006);
nand U5944 (N_5944,N_1231,N_1233);
nor U5945 (N_5945,N_778,N_1233);
and U5946 (N_5946,N_2193,N_1037);
nor U5947 (N_5947,N_1283,N_2933);
and U5948 (N_5948,N_1919,N_474);
nor U5949 (N_5949,N_2219,N_2523);
nor U5950 (N_5950,N_1339,N_1346);
or U5951 (N_5951,N_2345,N_2992);
or U5952 (N_5952,N_2412,N_2814);
xnor U5953 (N_5953,N_489,N_1907);
and U5954 (N_5954,N_1427,N_103);
nor U5955 (N_5955,N_2500,N_2621);
nor U5956 (N_5956,N_141,N_2753);
xor U5957 (N_5957,N_111,N_870);
nand U5958 (N_5958,N_916,N_628);
nor U5959 (N_5959,N_1724,N_2535);
nand U5960 (N_5960,N_2453,N_8);
and U5961 (N_5961,N_989,N_1777);
or U5962 (N_5962,N_1257,N_2328);
or U5963 (N_5963,N_2790,N_1894);
or U5964 (N_5964,N_2157,N_2215);
or U5965 (N_5965,N_802,N_1953);
xnor U5966 (N_5966,N_4,N_1957);
or U5967 (N_5967,N_1153,N_60);
nand U5968 (N_5968,N_839,N_1562);
and U5969 (N_5969,N_1497,N_2724);
nor U5970 (N_5970,N_2986,N_282);
xnor U5971 (N_5971,N_922,N_2186);
nor U5972 (N_5972,N_2460,N_437);
or U5973 (N_5973,N_235,N_117);
and U5974 (N_5974,N_2125,N_1050);
and U5975 (N_5975,N_411,N_395);
and U5976 (N_5976,N_189,N_2529);
and U5977 (N_5977,N_1415,N_1635);
and U5978 (N_5978,N_235,N_847);
and U5979 (N_5979,N_1826,N_1413);
or U5980 (N_5980,N_780,N_1827);
and U5981 (N_5981,N_1875,N_2164);
nor U5982 (N_5982,N_932,N_1974);
nand U5983 (N_5983,N_2626,N_895);
nor U5984 (N_5984,N_1547,N_1666);
nor U5985 (N_5985,N_2706,N_2901);
nor U5986 (N_5986,N_206,N_1476);
nor U5987 (N_5987,N_2254,N_880);
or U5988 (N_5988,N_1972,N_1228);
xnor U5989 (N_5989,N_1121,N_539);
xor U5990 (N_5990,N_2657,N_1332);
or U5991 (N_5991,N_1479,N_1506);
nand U5992 (N_5992,N_2805,N_9);
nand U5993 (N_5993,N_2427,N_199);
nand U5994 (N_5994,N_292,N_706);
or U5995 (N_5995,N_2109,N_2181);
xnor U5996 (N_5996,N_1695,N_2917);
or U5997 (N_5997,N_1523,N_2290);
nand U5998 (N_5998,N_2081,N_2126);
nand U5999 (N_5999,N_2670,N_2984);
nand U6000 (N_6000,N_3592,N_4590);
xnor U6001 (N_6001,N_4563,N_5633);
xnor U6002 (N_6002,N_4468,N_4606);
and U6003 (N_6003,N_5472,N_5622);
nor U6004 (N_6004,N_3907,N_4825);
and U6005 (N_6005,N_5067,N_4026);
xnor U6006 (N_6006,N_5405,N_3777);
or U6007 (N_6007,N_4278,N_3670);
and U6008 (N_6008,N_5425,N_4764);
or U6009 (N_6009,N_3635,N_4649);
or U6010 (N_6010,N_3321,N_4495);
nand U6011 (N_6011,N_3206,N_5703);
or U6012 (N_6012,N_4667,N_5450);
and U6013 (N_6013,N_3558,N_5154);
and U6014 (N_6014,N_5048,N_3312);
or U6015 (N_6015,N_3173,N_3926);
nand U6016 (N_6016,N_4378,N_4991);
or U6017 (N_6017,N_5266,N_4286);
and U6018 (N_6018,N_3970,N_4979);
nor U6019 (N_6019,N_3031,N_4214);
nand U6020 (N_6020,N_4928,N_5915);
nand U6021 (N_6021,N_4684,N_4845);
nor U6022 (N_6022,N_3574,N_5635);
xor U6023 (N_6023,N_3955,N_5458);
nand U6024 (N_6024,N_4110,N_5618);
and U6025 (N_6025,N_4582,N_3644);
nand U6026 (N_6026,N_5174,N_3057);
or U6027 (N_6027,N_4601,N_3211);
and U6028 (N_6028,N_3660,N_3408);
or U6029 (N_6029,N_4206,N_4063);
nor U6030 (N_6030,N_4349,N_4747);
and U6031 (N_6031,N_5889,N_3210);
or U6032 (N_6032,N_4467,N_4187);
nor U6033 (N_6033,N_5570,N_4524);
or U6034 (N_6034,N_4519,N_3772);
nand U6035 (N_6035,N_5448,N_4549);
nor U6036 (N_6036,N_4847,N_3274);
nand U6037 (N_6037,N_3172,N_3717);
nand U6038 (N_6038,N_3107,N_5874);
or U6039 (N_6039,N_5393,N_3056);
nand U6040 (N_6040,N_4257,N_5701);
nor U6041 (N_6041,N_4030,N_4351);
and U6042 (N_6042,N_4821,N_3367);
nor U6043 (N_6043,N_3728,N_3766);
or U6044 (N_6044,N_4093,N_5189);
and U6045 (N_6045,N_4108,N_5877);
or U6046 (N_6046,N_5024,N_5316);
nor U6047 (N_6047,N_4053,N_5246);
or U6048 (N_6048,N_4212,N_5010);
and U6049 (N_6049,N_5379,N_4967);
or U6050 (N_6050,N_5451,N_5653);
nand U6051 (N_6051,N_4782,N_4067);
nand U6052 (N_6052,N_4952,N_4746);
or U6053 (N_6053,N_3067,N_5408);
or U6054 (N_6054,N_5518,N_3437);
and U6055 (N_6055,N_3101,N_3829);
and U6056 (N_6056,N_4267,N_4607);
or U6057 (N_6057,N_5159,N_4365);
nand U6058 (N_6058,N_5418,N_5740);
xor U6059 (N_6059,N_5881,N_5052);
nor U6060 (N_6060,N_3477,N_4587);
or U6061 (N_6061,N_5878,N_5009);
or U6062 (N_6062,N_4045,N_3231);
nand U6063 (N_6063,N_4908,N_3718);
and U6064 (N_6064,N_5815,N_3234);
or U6065 (N_6065,N_3014,N_5319);
nor U6066 (N_6066,N_5085,N_3803);
and U6067 (N_6067,N_4511,N_3878);
xnor U6068 (N_6068,N_3520,N_3809);
or U6069 (N_6069,N_5867,N_5175);
or U6070 (N_6070,N_3815,N_5593);
or U6071 (N_6071,N_5003,N_4469);
xnor U6072 (N_6072,N_5515,N_3643);
nand U6073 (N_6073,N_5152,N_3919);
or U6074 (N_6074,N_5863,N_3517);
and U6075 (N_6075,N_4299,N_5489);
or U6076 (N_6076,N_4635,N_5111);
or U6077 (N_6077,N_5193,N_5713);
nand U6078 (N_6078,N_4562,N_3988);
and U6079 (N_6079,N_3962,N_5529);
xnor U6080 (N_6080,N_4665,N_5501);
and U6081 (N_6081,N_5767,N_3058);
and U6082 (N_6082,N_3171,N_4740);
or U6083 (N_6083,N_3114,N_4828);
nand U6084 (N_6084,N_4003,N_4573);
and U6085 (N_6085,N_5865,N_4732);
nor U6086 (N_6086,N_3534,N_5870);
nor U6087 (N_6087,N_4428,N_3227);
or U6088 (N_6088,N_5372,N_5310);
nand U6089 (N_6089,N_4103,N_4497);
nand U6090 (N_6090,N_4195,N_3432);
and U6091 (N_6091,N_5809,N_3868);
nand U6092 (N_6092,N_3911,N_5018);
xnor U6093 (N_6093,N_4543,N_5721);
nor U6094 (N_6094,N_3280,N_5141);
nor U6095 (N_6095,N_3200,N_3904);
nand U6096 (N_6096,N_5422,N_4217);
xnor U6097 (N_6097,N_3469,N_3886);
nor U6098 (N_6098,N_4589,N_3597);
nand U6099 (N_6099,N_5369,N_4728);
and U6100 (N_6100,N_3522,N_4865);
or U6101 (N_6101,N_4643,N_4997);
nor U6102 (N_6102,N_3253,N_4395);
xor U6103 (N_6103,N_4144,N_3615);
nor U6104 (N_6104,N_4670,N_3009);
nand U6105 (N_6105,N_5073,N_4614);
or U6106 (N_6106,N_4560,N_4001);
nand U6107 (N_6107,N_4145,N_3475);
nor U6108 (N_6108,N_4472,N_4827);
nand U6109 (N_6109,N_3339,N_4285);
nand U6110 (N_6110,N_3915,N_3472);
or U6111 (N_6111,N_5817,N_4906);
xnor U6112 (N_6112,N_3466,N_5922);
nor U6113 (N_6113,N_4430,N_5578);
nor U6114 (N_6114,N_3162,N_5226);
nand U6115 (N_6115,N_3272,N_5015);
nor U6116 (N_6116,N_5735,N_5732);
nor U6117 (N_6117,N_3608,N_4123);
nand U6118 (N_6118,N_4211,N_4554);
or U6119 (N_6119,N_4471,N_5247);
or U6120 (N_6120,N_5825,N_5259);
xnor U6121 (N_6121,N_4180,N_4948);
nor U6122 (N_6122,N_4968,N_5967);
nand U6123 (N_6123,N_5132,N_5019);
or U6124 (N_6124,N_5202,N_4444);
and U6125 (N_6125,N_5726,N_3512);
or U6126 (N_6126,N_4151,N_4427);
and U6127 (N_6127,N_3525,N_5114);
nand U6128 (N_6128,N_5241,N_4856);
or U6129 (N_6129,N_5575,N_5959);
nand U6130 (N_6130,N_4526,N_5964);
or U6131 (N_6131,N_4938,N_4013);
or U6132 (N_6132,N_4934,N_3205);
and U6133 (N_6133,N_5758,N_4333);
xor U6134 (N_6134,N_5199,N_4808);
or U6135 (N_6135,N_4687,N_5907);
xnor U6136 (N_6136,N_5394,N_5251);
nor U6137 (N_6137,N_3407,N_5745);
xor U6138 (N_6138,N_3706,N_3243);
nor U6139 (N_6139,N_5462,N_5161);
and U6140 (N_6140,N_3952,N_4954);
or U6141 (N_6141,N_3755,N_4447);
and U6142 (N_6142,N_3276,N_5936);
nand U6143 (N_6143,N_3602,N_5325);
nor U6144 (N_6144,N_3680,N_4458);
xor U6145 (N_6145,N_3805,N_5644);
or U6146 (N_6146,N_3286,N_4335);
and U6147 (N_6147,N_3527,N_4811);
or U6148 (N_6148,N_4319,N_5312);
nand U6149 (N_6149,N_5616,N_4885);
and U6150 (N_6150,N_5585,N_5945);
nand U6151 (N_6151,N_4522,N_3149);
nor U6152 (N_6152,N_4391,N_5315);
or U6153 (N_6153,N_5492,N_5228);
and U6154 (N_6154,N_3416,N_4581);
or U6155 (N_6155,N_5549,N_4245);
xnor U6156 (N_6156,N_5314,N_5296);
nor U6157 (N_6157,N_5017,N_3427);
or U6158 (N_6158,N_3861,N_5757);
or U6159 (N_6159,N_3596,N_4750);
and U6160 (N_6160,N_4059,N_3259);
or U6161 (N_6161,N_5185,N_3618);
or U6162 (N_6162,N_5514,N_3985);
nor U6163 (N_6163,N_5170,N_4377);
xnor U6164 (N_6164,N_3600,N_5493);
nor U6165 (N_6165,N_5704,N_5594);
nor U6166 (N_6166,N_5060,N_4357);
or U6167 (N_6167,N_5960,N_4647);
xnor U6168 (N_6168,N_4233,N_5939);
xnor U6169 (N_6169,N_3213,N_5370);
and U6170 (N_6170,N_3767,N_4588);
nor U6171 (N_6171,N_5357,N_4478);
xor U6172 (N_6172,N_3987,N_5563);
nand U6173 (N_6173,N_5951,N_5295);
xor U6174 (N_6174,N_5510,N_5790);
xor U6175 (N_6175,N_4939,N_5536);
and U6176 (N_6176,N_3214,N_4350);
nand U6177 (N_6177,N_4328,N_3310);
or U6178 (N_6178,N_3325,N_4314);
or U6179 (N_6179,N_3671,N_5538);
nand U6180 (N_6180,N_3697,N_4096);
xor U6181 (N_6181,N_5475,N_3724);
nand U6182 (N_6182,N_4441,N_3871);
nor U6183 (N_6183,N_4850,N_4048);
nor U6184 (N_6184,N_4612,N_4896);
and U6185 (N_6185,N_3548,N_4602);
or U6186 (N_6186,N_4733,N_4512);
nand U6187 (N_6187,N_4345,N_3323);
nand U6188 (N_6188,N_4073,N_3943);
and U6189 (N_6189,N_3735,N_5620);
xnor U6190 (N_6190,N_5348,N_4840);
nand U6191 (N_6191,N_3867,N_4824);
xor U6192 (N_6192,N_4942,N_4548);
or U6193 (N_6193,N_5780,N_5664);
nor U6194 (N_6194,N_4773,N_5139);
or U6195 (N_6195,N_5420,N_3555);
nor U6196 (N_6196,N_3598,N_4851);
and U6197 (N_6197,N_5203,N_3355);
nand U6198 (N_6198,N_5172,N_5974);
or U6199 (N_6199,N_5988,N_5088);
nor U6200 (N_6200,N_5906,N_3403);
xor U6201 (N_6201,N_4933,N_5649);
nor U6202 (N_6202,N_3072,N_5120);
or U6203 (N_6203,N_4685,N_4136);
nor U6204 (N_6204,N_3147,N_4523);
nand U6205 (N_6205,N_5699,N_4783);
or U6206 (N_6206,N_5350,N_5797);
or U6207 (N_6207,N_3792,N_5943);
or U6208 (N_6208,N_3622,N_5129);
nand U6209 (N_6209,N_5160,N_3358);
nor U6210 (N_6210,N_3939,N_3573);
or U6211 (N_6211,N_5537,N_3267);
or U6212 (N_6212,N_4630,N_3509);
xnor U6213 (N_6213,N_5971,N_4955);
nand U6214 (N_6214,N_4655,N_3664);
or U6215 (N_6215,N_4022,N_5381);
and U6216 (N_6216,N_5102,N_4150);
or U6217 (N_6217,N_3681,N_5094);
or U6218 (N_6218,N_5720,N_3889);
and U6219 (N_6219,N_4321,N_5195);
xnor U6220 (N_6220,N_3774,N_4250);
nand U6221 (N_6221,N_3983,N_3699);
xnor U6222 (N_6222,N_5897,N_5993);
nand U6223 (N_6223,N_3738,N_5455);
and U6224 (N_6224,N_4004,N_4537);
nor U6225 (N_6225,N_5207,N_3158);
nand U6226 (N_6226,N_4221,N_4658);
and U6227 (N_6227,N_4631,N_5444);
nand U6228 (N_6228,N_5920,N_5846);
nand U6229 (N_6229,N_5268,N_3941);
nor U6230 (N_6230,N_5899,N_4674);
or U6231 (N_6231,N_5321,N_4404);
or U6232 (N_6232,N_3478,N_3316);
or U6233 (N_6233,N_5747,N_4291);
and U6234 (N_6234,N_3458,N_5068);
xnor U6235 (N_6235,N_4705,N_3492);
nor U6236 (N_6236,N_4288,N_4735);
nand U6237 (N_6237,N_3306,N_5014);
nand U6238 (N_6238,N_3081,N_3197);
xnor U6239 (N_6239,N_3219,N_5516);
or U6240 (N_6240,N_5359,N_3595);
and U6241 (N_6241,N_4817,N_4356);
nand U6242 (N_6242,N_4005,N_3693);
and U6243 (N_6243,N_3552,N_3150);
and U6244 (N_6244,N_5416,N_4722);
nor U6245 (N_6245,N_4886,N_3828);
and U6246 (N_6246,N_3011,N_4303);
xnor U6247 (N_6247,N_4717,N_4400);
or U6248 (N_6248,N_3603,N_4011);
or U6249 (N_6249,N_5368,N_5366);
nand U6250 (N_6250,N_5641,N_4198);
or U6251 (N_6251,N_5816,N_5142);
and U6252 (N_6252,N_4837,N_5566);
and U6253 (N_6253,N_3048,N_3523);
nor U6254 (N_6254,N_4055,N_4800);
nor U6255 (N_6255,N_3185,N_4504);
nand U6256 (N_6256,N_3958,N_3434);
nor U6257 (N_6257,N_4691,N_5900);
and U6258 (N_6258,N_3117,N_5932);
nor U6259 (N_6259,N_3365,N_3599);
and U6260 (N_6260,N_3570,N_5206);
xnor U6261 (N_6261,N_3584,N_4092);
nor U6262 (N_6262,N_5559,N_5064);
nor U6263 (N_6263,N_5496,N_4791);
nor U6264 (N_6264,N_4927,N_5961);
and U6265 (N_6265,N_5283,N_5684);
and U6266 (N_6266,N_4081,N_3455);
nor U6267 (N_6267,N_4429,N_5991);
and U6268 (N_6268,N_3324,N_4422);
nand U6269 (N_6269,N_5008,N_3052);
and U6270 (N_6270,N_3152,N_4442);
and U6271 (N_6271,N_4390,N_5253);
or U6272 (N_6272,N_5509,N_5613);
nor U6273 (N_6273,N_5390,N_5040);
nand U6274 (N_6274,N_3816,N_3497);
and U6275 (N_6275,N_4204,N_3183);
and U6276 (N_6276,N_4957,N_3189);
and U6277 (N_6277,N_5335,N_4381);
xor U6278 (N_6278,N_4456,N_5969);
and U6279 (N_6279,N_4290,N_3181);
nand U6280 (N_6280,N_4699,N_5269);
and U6281 (N_6281,N_4473,N_5488);
nand U6282 (N_6282,N_3730,N_5115);
nor U6283 (N_6283,N_5949,N_3649);
xnor U6284 (N_6284,N_5046,N_5364);
nor U6285 (N_6285,N_4087,N_3372);
xor U6286 (N_6286,N_4986,N_3975);
nand U6287 (N_6287,N_5069,N_5551);
or U6288 (N_6288,N_5460,N_3876);
and U6289 (N_6289,N_3033,N_5947);
and U6290 (N_6290,N_3375,N_4215);
nor U6291 (N_6291,N_4237,N_5121);
nand U6292 (N_6292,N_4348,N_4510);
nor U6293 (N_6293,N_5914,N_5354);
nand U6294 (N_6294,N_4415,N_4836);
or U6295 (N_6295,N_4985,N_3508);
or U6296 (N_6296,N_3559,N_3490);
or U6297 (N_6297,N_3337,N_3084);
or U6298 (N_6298,N_5543,N_5738);
or U6299 (N_6299,N_3529,N_3551);
or U6300 (N_6300,N_5968,N_3927);
and U6301 (N_6301,N_5568,N_3873);
and U6302 (N_6302,N_3022,N_3821);
or U6303 (N_6303,N_5667,N_4281);
and U6304 (N_6304,N_4812,N_5293);
nor U6305 (N_6305,N_5334,N_3237);
nor U6306 (N_6306,N_5693,N_5412);
or U6307 (N_6307,N_4751,N_3795);
nor U6308 (N_6308,N_3630,N_4056);
and U6309 (N_6309,N_3344,N_4173);
and U6310 (N_6310,N_5157,N_3604);
xor U6311 (N_6311,N_3505,N_3757);
nand U6312 (N_6312,N_3182,N_5326);
nor U6313 (N_6313,N_4394,N_3376);
nor U6314 (N_6314,N_4608,N_5117);
nor U6315 (N_6315,N_3141,N_3217);
and U6316 (N_6316,N_5051,N_4527);
nand U6317 (N_6317,N_4373,N_3187);
nor U6318 (N_6318,N_3661,N_4780);
or U6319 (N_6319,N_4682,N_3725);
or U6320 (N_6320,N_4871,N_3381);
or U6321 (N_6321,N_4869,N_5905);
or U6322 (N_6322,N_3361,N_4520);
or U6323 (N_6323,N_5601,N_5665);
and U6324 (N_6324,N_5727,N_3963);
nor U6325 (N_6325,N_4555,N_4709);
or U6326 (N_6326,N_3575,N_4966);
or U6327 (N_6327,N_3111,N_5112);
and U6328 (N_6328,N_4192,N_4793);
and U6329 (N_6329,N_4597,N_3743);
and U6330 (N_6330,N_4044,N_4336);
nor U6331 (N_6331,N_3746,N_3960);
and U6332 (N_6332,N_4693,N_3802);
or U6333 (N_6333,N_3108,N_4179);
xor U6334 (N_6334,N_4162,N_3252);
nand U6335 (N_6335,N_4009,N_3647);
nor U6336 (N_6336,N_4463,N_5131);
xnor U6337 (N_6337,N_5540,N_5386);
nand U6338 (N_6338,N_4010,N_4556);
and U6339 (N_6339,N_5500,N_3175);
nand U6340 (N_6340,N_4710,N_4755);
nor U6341 (N_6341,N_4553,N_4690);
nand U6342 (N_6342,N_3918,N_5805);
or U6343 (N_6343,N_4625,N_3413);
or U6344 (N_6344,N_5572,N_5119);
nor U6345 (N_6345,N_5642,N_5940);
nand U6346 (N_6346,N_5965,N_3328);
and U6347 (N_6347,N_5313,N_5191);
and U6348 (N_6348,N_4894,N_3102);
or U6349 (N_6349,N_3255,N_3190);
nor U6350 (N_6350,N_5859,N_4315);
and U6351 (N_6351,N_5486,N_4716);
and U6352 (N_6352,N_5554,N_5292);
or U6353 (N_6353,N_5985,N_4701);
nor U6354 (N_6354,N_4517,N_3160);
and U6355 (N_6355,N_5886,N_4920);
nor U6356 (N_6356,N_4953,N_5777);
or U6357 (N_6357,N_4366,N_3165);
nor U6358 (N_6358,N_3311,N_4318);
nor U6359 (N_6359,N_5151,N_4593);
or U6360 (N_6360,N_4175,N_3637);
or U6361 (N_6361,N_3675,N_3199);
and U6362 (N_6362,N_3571,N_3619);
xor U6363 (N_6363,N_4362,N_5103);
and U6364 (N_6364,N_4500,N_3068);
or U6365 (N_6365,N_4460,N_3715);
or U6366 (N_6366,N_5101,N_5983);
or U6367 (N_6367,N_3864,N_3414);
nand U6368 (N_6368,N_4646,N_4960);
and U6369 (N_6369,N_4509,N_4226);
and U6370 (N_6370,N_5996,N_4703);
nand U6371 (N_6371,N_3357,N_3156);
or U6372 (N_6372,N_4626,N_3446);
nand U6373 (N_6373,N_5049,N_3070);
nand U6374 (N_6374,N_3953,N_5007);
nor U6375 (N_6375,N_4032,N_5751);
nor U6376 (N_6376,N_5034,N_4758);
or U6377 (N_6377,N_4265,N_4421);
nor U6378 (N_6378,N_3521,N_4359);
and U6379 (N_6379,N_5477,N_3665);
nand U6380 (N_6380,N_3921,N_3236);
nand U6381 (N_6381,N_3817,N_5077);
nor U6382 (N_6382,N_4207,N_4251);
or U6383 (N_6383,N_4613,N_3650);
or U6384 (N_6384,N_5555,N_3587);
nand U6385 (N_6385,N_5360,N_4858);
or U6386 (N_6386,N_3275,N_5771);
nand U6387 (N_6387,N_3703,N_3010);
and U6388 (N_6388,N_3026,N_4989);
or U6389 (N_6389,N_3530,N_4666);
or U6390 (N_6390,N_5503,N_3007);
xnor U6391 (N_6391,N_5629,N_5508);
or U6392 (N_6392,N_5453,N_3393);
or U6393 (N_6393,N_4830,N_3928);
nor U6394 (N_6394,N_3419,N_5020);
nor U6395 (N_6395,N_3425,N_5869);
and U6396 (N_6396,N_4470,N_4323);
or U6397 (N_6397,N_5522,N_3341);
nor U6398 (N_6398,N_5090,N_4550);
nor U6399 (N_6399,N_4564,N_3966);
xor U6400 (N_6400,N_3854,N_4815);
or U6401 (N_6401,N_5238,N_4079);
nand U6402 (N_6402,N_5437,N_4756);
and U6403 (N_6403,N_3999,N_4713);
nand U6404 (N_6404,N_4901,N_4165);
nor U6405 (N_6405,N_5567,N_5628);
and U6406 (N_6406,N_5999,N_5523);
or U6407 (N_6407,N_5491,N_5668);
or U6408 (N_6408,N_4706,N_4700);
or U6409 (N_6409,N_3051,N_4477);
nand U6410 (N_6410,N_5276,N_3794);
and U6411 (N_6411,N_5768,N_5729);
nand U6412 (N_6412,N_5573,N_3557);
and U6413 (N_6413,N_5934,N_5045);
and U6414 (N_6414,N_3689,N_3184);
nor U6415 (N_6415,N_5320,N_3230);
xnor U6416 (N_6416,N_3159,N_4785);
nor U6417 (N_6417,N_5081,N_4946);
nand U6418 (N_6418,N_3502,N_4981);
and U6419 (N_6419,N_3288,N_4853);
nand U6420 (N_6420,N_4169,N_3526);
or U6421 (N_6421,N_4102,N_5162);
or U6422 (N_6422,N_3621,N_4999);
or U6423 (N_6423,N_4343,N_5339);
and U6424 (N_6424,N_4576,N_4737);
nor U6425 (N_6425,N_5957,N_3947);
and U6426 (N_6426,N_5337,N_5474);
or U6427 (N_6427,N_4132,N_5106);
or U6428 (N_6428,N_5465,N_3627);
nand U6429 (N_6429,N_5862,N_3350);
nor U6430 (N_6430,N_4141,N_5801);
or U6431 (N_6431,N_4481,N_3113);
nor U6432 (N_6432,N_5205,N_3345);
and U6433 (N_6433,N_4763,N_5798);
or U6434 (N_6434,N_3247,N_4086);
nand U6435 (N_6435,N_3279,N_3790);
and U6436 (N_6436,N_5875,N_5855);
and U6437 (N_6437,N_3956,N_3320);
nand U6438 (N_6438,N_5519,N_5868);
xor U6439 (N_6439,N_3428,N_5788);
and U6440 (N_6440,N_4459,N_3761);
xor U6441 (N_6441,N_4833,N_5431);
or U6442 (N_6442,N_4064,N_3696);
xor U6443 (N_6443,N_5227,N_5970);
nor U6444 (N_6444,N_3503,N_4124);
or U6445 (N_6445,N_5098,N_5531);
nor U6446 (N_6446,N_3859,N_4983);
and U6447 (N_6447,N_5650,N_4771);
or U6448 (N_6448,N_4829,N_5910);
and U6449 (N_6449,N_5769,N_3763);
nand U6450 (N_6450,N_4718,N_3511);
nand U6451 (N_6451,N_4197,N_3006);
nand U6452 (N_6452,N_5630,N_4544);
and U6453 (N_6453,N_3139,N_5239);
and U6454 (N_6454,N_5130,N_4654);
or U6455 (N_6455,N_3613,N_4881);
and U6456 (N_6456,N_5730,N_3883);
or U6457 (N_6457,N_4070,N_4117);
and U6458 (N_6458,N_5061,N_3099);
xor U6459 (N_6459,N_3925,N_3391);
or U6460 (N_6460,N_3385,N_5011);
or U6461 (N_6461,N_3336,N_3013);
nor U6462 (N_6462,N_4702,N_4731);
nor U6463 (N_6463,N_4772,N_3695);
and U6464 (N_6464,N_5625,N_3285);
nand U6465 (N_6465,N_3076,N_4163);
and U6466 (N_6466,N_5746,N_3196);
nor U6467 (N_6467,N_4249,N_5560);
nand U6468 (N_6468,N_5445,N_5552);
or U6469 (N_6469,N_4577,N_3305);
nand U6470 (N_6470,N_3842,N_5604);
and U6471 (N_6471,N_4534,N_5066);
and U6472 (N_6472,N_3631,N_5376);
nor U6473 (N_6473,N_5646,N_3489);
or U6474 (N_6474,N_5255,N_3969);
or U6475 (N_6475,N_4752,N_4998);
or U6476 (N_6476,N_4041,N_4903);
and U6477 (N_6477,N_3762,N_4271);
or U6478 (N_6478,N_3863,N_3374);
or U6479 (N_6479,N_5753,N_5070);
and U6480 (N_6480,N_5356,N_5224);
and U6481 (N_6481,N_5415,N_4177);
nor U6482 (N_6482,N_3096,N_5791);
or U6483 (N_6483,N_4383,N_5929);
nor U6484 (N_6484,N_5443,N_3832);
nor U6485 (N_6485,N_3784,N_5225);
or U6486 (N_6486,N_4638,N_4058);
and U6487 (N_6487,N_5062,N_4571);
or U6488 (N_6488,N_3193,N_3454);
nand U6489 (N_6489,N_3204,N_5076);
nor U6490 (N_6490,N_5404,N_3287);
or U6491 (N_6491,N_5436,N_3676);
nand U6492 (N_6492,N_5958,N_4977);
and U6493 (N_6493,N_5291,N_3115);
or U6494 (N_6494,N_3788,N_3248);
or U6495 (N_6495,N_5639,N_5728);
nand U6496 (N_6496,N_3655,N_4978);
nand U6497 (N_6497,N_4921,N_3959);
nand U6498 (N_6498,N_4516,N_5526);
nor U6499 (N_6499,N_5311,N_5158);
or U6500 (N_6500,N_5715,N_3524);
nor U6501 (N_6501,N_4742,N_4804);
nand U6502 (N_6502,N_4521,N_5832);
nor U6503 (N_6503,N_4027,N_4813);
nor U6504 (N_6504,N_5811,N_5597);
nand U6505 (N_6505,N_3764,N_5036);
nor U6506 (N_6506,N_4767,N_3968);
nand U6507 (N_6507,N_3405,N_3411);
or U6508 (N_6508,N_5478,N_3617);
and U6509 (N_6509,N_3540,N_5888);
xor U6510 (N_6510,N_3768,N_4199);
or U6511 (N_6511,N_5402,N_3594);
or U6512 (N_6512,N_5147,N_4437);
nor U6513 (N_6513,N_4583,N_5694);
xnor U6514 (N_6514,N_5822,N_4907);
nand U6515 (N_6515,N_3636,N_5651);
nor U6516 (N_6516,N_3290,N_3239);
and U6517 (N_6517,N_5710,N_3862);
and U6518 (N_6518,N_3382,N_4963);
and U6519 (N_6519,N_4883,N_4809);
or U6520 (N_6520,N_5495,N_5783);
xor U6521 (N_6521,N_3299,N_4436);
nor U6522 (N_6522,N_3747,N_5528);
nand U6523 (N_6523,N_5748,N_5397);
or U6524 (N_6524,N_3484,N_5884);
nor U6525 (N_6525,N_4020,N_5930);
nor U6526 (N_6526,N_5845,N_3877);
nor U6527 (N_6527,N_4264,N_3130);
nand U6528 (N_6528,N_4152,N_3420);
nand U6529 (N_6529,N_3168,N_5284);
or U6530 (N_6530,N_4313,N_3822);
or U6531 (N_6531,N_4317,N_3798);
nand U6532 (N_6532,N_4276,N_3704);
and U6533 (N_6533,N_5187,N_4050);
nand U6534 (N_6534,N_4448,N_5784);
nor U6535 (N_6535,N_3719,N_4476);
xor U6536 (N_6536,N_4514,N_4801);
and U6537 (N_6537,N_5355,N_4239);
nand U6538 (N_6538,N_4157,N_5184);
and U6539 (N_6539,N_4852,N_5249);
nor U6540 (N_6540,N_4068,N_3964);
xnor U6541 (N_6541,N_5485,N_4438);
xnor U6542 (N_6542,N_4229,N_4134);
or U6543 (N_6543,N_5885,N_4446);
nand U6544 (N_6544,N_4120,N_4085);
and U6545 (N_6545,N_4223,N_5499);
nor U6546 (N_6546,N_3077,N_5789);
nor U6547 (N_6547,N_3188,N_3753);
or U6548 (N_6548,N_5403,N_5761);
nand U6549 (N_6549,N_5307,N_5279);
nand U6550 (N_6550,N_4765,N_4542);
and U6551 (N_6551,N_5589,N_4639);
and U6552 (N_6552,N_5609,N_3018);
and U6553 (N_6553,N_4066,N_5371);
nand U6554 (N_6554,N_4499,N_5923);
nor U6555 (N_6555,N_4552,N_5979);
and U6556 (N_6556,N_4155,N_5047);
nor U6557 (N_6557,N_4410,N_3946);
xor U6558 (N_6558,N_3338,N_5303);
nand U6559 (N_6559,N_4399,N_3049);
nand U6560 (N_6560,N_3148,N_3008);
or U6561 (N_6561,N_3457,N_4761);
nor U6562 (N_6562,N_4680,N_5299);
and U6563 (N_6563,N_3998,N_5619);
nand U6564 (N_6564,N_4219,N_4679);
or U6565 (N_6565,N_5030,N_3054);
xor U6566 (N_6566,N_5756,N_4474);
or U6567 (N_6567,N_4924,N_4475);
and U6568 (N_6568,N_4541,N_4433);
nor U6569 (N_6569,N_3709,N_4949);
nand U6570 (N_6570,N_5733,N_3024);
xor U6571 (N_6571,N_3810,N_3770);
nand U6572 (N_6572,N_4565,N_5035);
xnor U6573 (N_6573,N_5377,N_3060);
or U6574 (N_6574,N_4243,N_3448);
and U6575 (N_6575,N_4324,N_3125);
xnor U6576 (N_6576,N_5902,N_5942);
and U6577 (N_6577,N_4419,N_3846);
or U6578 (N_6578,N_5787,N_5610);
or U6579 (N_6579,N_3899,N_3929);
nand U6580 (N_6580,N_5002,N_4258);
and U6581 (N_6581,N_4178,N_3322);
or U6582 (N_6582,N_4842,N_3882);
nand U6583 (N_6583,N_3565,N_4660);
nand U6584 (N_6584,N_3470,N_3186);
nand U6585 (N_6585,N_4872,N_4925);
or U6586 (N_6586,N_3265,N_3914);
nor U6587 (N_6587,N_5793,N_4624);
and U6588 (N_6588,N_3412,N_5954);
nand U6589 (N_6589,N_4860,N_5401);
nand U6590 (N_6590,N_5308,N_5380);
xnor U6591 (N_6591,N_4186,N_3658);
nor U6592 (N_6592,N_5762,N_5190);
nand U6593 (N_6593,N_4633,N_3221);
or U6594 (N_6594,N_5941,N_3813);
nand U6595 (N_6595,N_4382,N_4816);
and U6596 (N_6596,N_5186,N_5786);
and U6597 (N_6597,N_3027,N_5533);
nor U6598 (N_6598,N_5361,N_5517);
nand U6599 (N_6599,N_5140,N_3727);
or U6600 (N_6600,N_3435,N_4205);
nand U6601 (N_6601,N_3778,N_4692);
nor U6602 (N_6602,N_4877,N_5221);
xnor U6603 (N_6603,N_3346,N_3123);
or U6604 (N_6604,N_5956,N_4049);
xor U6605 (N_6605,N_5584,N_5084);
nand U6606 (N_6606,N_4603,N_3977);
or U6607 (N_6607,N_4533,N_5297);
and U6608 (N_6608,N_3769,N_5580);
or U6609 (N_6609,N_3388,N_3733);
nand U6610 (N_6610,N_5711,N_3289);
xnor U6611 (N_6611,N_4171,N_5723);
nand U6612 (N_6612,N_3993,N_4950);
nand U6613 (N_6613,N_3894,N_3086);
or U6614 (N_6614,N_4224,N_5074);
or U6615 (N_6615,N_5469,N_5582);
or U6616 (N_6616,N_3377,N_5244);
nand U6617 (N_6617,N_3354,N_3935);
or U6618 (N_6618,N_3097,N_4929);
xor U6619 (N_6619,N_3610,N_3304);
and U6620 (N_6620,N_4038,N_5534);
xor U6621 (N_6621,N_5016,N_5909);
nor U6622 (N_6622,N_4112,N_4502);
and U6623 (N_6623,N_4720,N_4396);
and U6624 (N_6624,N_5818,N_5346);
nand U6625 (N_6625,N_3415,N_4652);
and U6626 (N_6626,N_5146,N_5171);
xor U6627 (N_6627,N_4803,N_4642);
or U6628 (N_6628,N_5937,N_3398);
and U6629 (N_6629,N_5231,N_4200);
or U6630 (N_6630,N_5849,N_3853);
or U6631 (N_6631,N_4014,N_3811);
or U6632 (N_6632,N_5075,N_4367);
and U6633 (N_6633,N_3441,N_5079);
and U6634 (N_6634,N_4413,N_3043);
or U6635 (N_6635,N_5038,N_4518);
nor U6636 (N_6636,N_4089,N_4834);
nor U6637 (N_6637,N_4182,N_5854);
nand U6638 (N_6638,N_3218,N_3447);
or U6639 (N_6639,N_4982,N_5179);
and U6640 (N_6640,N_5200,N_5918);
nor U6641 (N_6641,N_5056,N_5569);
and U6642 (N_6642,N_3973,N_5395);
or U6643 (N_6643,N_3701,N_4861);
and U6644 (N_6644,N_4408,N_4222);
or U6645 (N_6645,N_4931,N_4806);
nor U6646 (N_6646,N_5953,N_5242);
nand U6647 (N_6647,N_3913,N_3452);
nand U6648 (N_6648,N_5271,N_5835);
nand U6649 (N_6649,N_3986,N_4420);
nand U6650 (N_6650,N_5828,N_5138);
nor U6651 (N_6651,N_4018,N_3028);
and U6652 (N_6652,N_3760,N_5736);
and U6653 (N_6653,N_5057,N_5349);
and U6654 (N_6654,N_3910,N_3167);
or U6655 (N_6655,N_3269,N_5280);
nor U6656 (N_6656,N_4984,N_5772);
nor U6657 (N_6657,N_3646,N_5384);
or U6658 (N_6658,N_4188,N_5608);
nand U6659 (N_6659,N_3166,N_3965);
or U6660 (N_6660,N_4088,N_5428);
and U6661 (N_6661,N_3088,N_3082);
and U6662 (N_6662,N_4873,N_3930);
and U6663 (N_6663,N_5133,N_5795);
or U6664 (N_6664,N_5634,N_4277);
nor U6665 (N_6665,N_4225,N_3888);
or U6666 (N_6666,N_4329,N_3742);
nor U6667 (N_6667,N_3012,N_3137);
nand U6668 (N_6668,N_4849,N_3754);
xnor U6669 (N_6669,N_5282,N_4236);
or U6670 (N_6670,N_3241,N_5483);
nor U6671 (N_6671,N_3110,N_3394);
nor U6672 (N_6672,N_4676,N_3277);
nand U6673 (N_6673,N_4297,N_5542);
nor U6674 (N_6674,N_3036,N_5136);
or U6675 (N_6675,N_5716,N_5333);
nand U6676 (N_6676,N_4487,N_3900);
and U6677 (N_6677,N_3896,N_5423);
and U6678 (N_6678,N_5663,N_4401);
nor U6679 (N_6679,N_5143,N_4961);
and U6680 (N_6680,N_3004,N_4870);
nor U6681 (N_6681,N_5351,N_3640);
nor U6682 (N_6682,N_5498,N_4790);
xnor U6683 (N_6683,N_3967,N_3363);
xnor U6684 (N_6684,N_5301,N_3154);
nor U6685 (N_6685,N_3944,N_4153);
and U6686 (N_6686,N_5541,N_3294);
xor U6687 (N_6687,N_5782,N_5879);
and U6688 (N_6688,N_5166,N_4507);
nand U6689 (N_6689,N_4936,N_3330);
xor U6690 (N_6690,N_5124,N_3368);
and U6691 (N_6691,N_3396,N_4133);
nor U6692 (N_6692,N_5164,N_4738);
or U6693 (N_6693,N_4493,N_4943);
and U6694 (N_6694,N_4839,N_3083);
or U6695 (N_6695,N_3244,N_4570);
nand U6696 (N_6696,N_3736,N_4266);
and U6697 (N_6697,N_3654,N_4914);
xnor U6698 (N_6698,N_5938,N_3633);
and U6699 (N_6699,N_3569,N_4913);
and U6700 (N_6700,N_4611,N_5265);
nor U6701 (N_6701,N_5466,N_4760);
or U6702 (N_6702,N_5342,N_3418);
or U6703 (N_6703,N_4254,N_3824);
nor U6704 (N_6704,N_3532,N_4361);
and U6705 (N_6705,N_4140,N_4300);
nor U6706 (N_6706,N_4768,N_3782);
and U6707 (N_6707,N_3677,N_5201);
nor U6708 (N_6708,N_4407,N_5926);
nand U6709 (N_6709,N_5617,N_3721);
xor U6710 (N_6710,N_5389,N_4664);
or U6711 (N_6711,N_5215,N_3645);
nor U6712 (N_6712,N_3583,N_5648);
and U6713 (N_6713,N_3937,N_3866);
xnor U6714 (N_6714,N_4370,N_3836);
nor U6715 (N_6715,N_3518,N_3995);
or U6716 (N_6716,N_5096,N_5898);
nor U6717 (N_6717,N_3669,N_4402);
or U6718 (N_6718,N_3780,N_3079);
nor U6719 (N_6719,N_3745,N_5148);
and U6720 (N_6720,N_5407,N_4130);
nand U6721 (N_6721,N_5547,N_3050);
xor U6722 (N_6722,N_3708,N_3685);
xor U6723 (N_6723,N_5666,N_4786);
nand U6724 (N_6724,N_4988,N_4031);
nor U6725 (N_6725,N_5258,N_3547);
and U6726 (N_6726,N_4574,N_4455);
xnor U6727 (N_6727,N_5300,N_3273);
or U6728 (N_6728,N_3342,N_4697);
nor U6729 (N_6729,N_5994,N_5041);
and U6730 (N_6730,N_5220,N_4868);
and U6731 (N_6731,N_4892,N_5814);
or U6732 (N_6732,N_4439,N_4558);
or U6733 (N_6733,N_4228,N_4959);
nand U6734 (N_6734,N_4805,N_4127);
and U6735 (N_6735,N_4218,N_5134);
and U6736 (N_6736,N_4726,N_3564);
or U6737 (N_6737,N_5657,N_3436);
xnor U6738 (N_6738,N_4434,N_4107);
nand U6739 (N_6739,N_5779,N_3127);
xor U6740 (N_6740,N_3625,N_3787);
or U6741 (N_6741,N_4138,N_4741);
nor U6742 (N_6742,N_5218,N_3556);
or U6743 (N_6743,N_5858,N_5741);
or U6744 (N_6744,N_4418,N_4598);
and U6745 (N_6745,N_3261,N_3546);
nand U6746 (N_6746,N_4326,N_5928);
nor U6747 (N_6747,N_5198,N_5755);
nor U6748 (N_6748,N_5217,N_5919);
and U6749 (N_6749,N_5864,N_4940);
and U6750 (N_6750,N_4076,N_5059);
nor U6751 (N_6751,N_3820,N_5841);
nand U6752 (N_6752,N_4284,N_5240);
or U6753 (N_6753,N_5302,N_3875);
nor U6754 (N_6754,N_4097,N_4887);
or U6755 (N_6755,N_3474,N_4322);
nand U6756 (N_6756,N_4792,N_4696);
nor U6757 (N_6757,N_4584,N_4262);
nand U6758 (N_6758,N_4307,N_5670);
or U6759 (N_6759,N_3586,N_3553);
nand U6760 (N_6760,N_4610,N_4101);
and U6761 (N_6761,N_4992,N_4306);
or U6762 (N_6762,N_5086,N_4453);
nand U6763 (N_6763,N_4681,N_3103);
nor U6764 (N_6764,N_3422,N_3976);
and U6765 (N_6765,N_3045,N_4566);
nor U6766 (N_6766,N_4183,N_3510);
or U6767 (N_6767,N_5776,N_5562);
or U6768 (N_6768,N_5921,N_3395);
nand U6769 (N_6769,N_4678,N_3356);
nor U6770 (N_6770,N_3626,N_5636);
or U6771 (N_6771,N_4168,N_3202);
nor U6772 (N_6772,N_3215,N_5391);
and U6773 (N_6773,N_3948,N_5270);
nand U6774 (N_6774,N_5340,N_3169);
nor U6775 (N_6775,N_4874,N_5454);
xor U6776 (N_6776,N_4591,N_5722);
nand U6777 (N_6777,N_5759,N_4776);
xor U6778 (N_6778,N_4386,N_3078);
and U6779 (N_6779,N_4976,N_5235);
and U6780 (N_6780,N_5579,N_4384);
nor U6781 (N_6781,N_4595,N_3850);
and U6782 (N_6782,N_4794,N_3431);
or U6783 (N_6783,N_3835,N_3450);
nor U6784 (N_6784,N_5257,N_5234);
or U6785 (N_6785,N_3283,N_3837);
or U6786 (N_6786,N_4668,N_5842);
or U6787 (N_6787,N_4368,N_3263);
and U6788 (N_6788,N_4725,N_3812);
or U6789 (N_6789,N_4600,N_4798);
or U6790 (N_6790,N_3922,N_4708);
nand U6791 (N_6791,N_4547,N_3430);
nor U6792 (N_6792,N_3834,N_5338);
xnor U6793 (N_6793,N_5400,N_4019);
nand U6794 (N_6794,N_5078,N_4488);
or U6795 (N_6795,N_4990,N_4917);
or U6796 (N_6796,N_3133,N_4308);
and U6797 (N_6797,N_3386,N_3260);
and U6798 (N_6798,N_5632,N_5546);
nor U6799 (N_6799,N_3192,N_5765);
nor U6800 (N_6800,N_5681,N_4166);
and U6801 (N_6801,N_4888,N_3471);
xor U6802 (N_6802,N_4406,N_4047);
nand U6803 (N_6803,N_5539,N_4358);
and U6804 (N_6804,N_4283,N_5093);
and U6805 (N_6805,N_3410,N_5605);
or U6806 (N_6806,N_5482,N_5698);
and U6807 (N_6807,N_4486,N_5487);
nand U6808 (N_6808,N_4457,N_5233);
nor U6809 (N_6809,N_4035,N_5544);
nor U6810 (N_6810,N_4332,N_3232);
xnor U6811 (N_6811,N_4298,N_5480);
or U6812 (N_6812,N_4605,N_4802);
and U6813 (N_6813,N_5260,N_4891);
nand U6814 (N_6814,N_4184,N_5434);
or U6815 (N_6815,N_4973,N_3370);
nand U6816 (N_6816,N_3445,N_3157);
and U6817 (N_6817,N_5375,N_4972);
and U6818 (N_6818,N_5216,N_3439);
or U6819 (N_6819,N_4409,N_3950);
xnor U6820 (N_6820,N_3319,N_3229);
or U6821 (N_6821,N_3945,N_3590);
or U6822 (N_6822,N_3062,N_4454);
nor U6823 (N_6823,N_5323,N_5127);
or U6824 (N_6824,N_5627,N_3424);
and U6825 (N_6825,N_5588,N_5181);
or U6826 (N_6826,N_3852,N_3690);
and U6827 (N_6827,N_5071,N_3700);
nor U6828 (N_6828,N_4393,N_3313);
or U6829 (N_6829,N_5676,N_4062);
nor U6830 (N_6830,N_4125,N_4287);
nand U6831 (N_6831,N_3838,N_3104);
nor U6832 (N_6832,N_3632,N_3002);
or U6833 (N_6833,N_3225,N_5586);
xor U6834 (N_6834,N_3544,N_5033);
or U6835 (N_6835,N_3823,N_3849);
and U6836 (N_6836,N_5638,N_3651);
nand U6837 (N_6837,N_5054,N_4292);
or U6838 (N_6838,N_4389,N_5691);
and U6839 (N_6839,N_5063,N_5532);
nand U6840 (N_6840,N_3262,N_5267);
and U6841 (N_6841,N_4848,N_4592);
nor U6842 (N_6842,N_5766,N_3481);
and U6843 (N_6843,N_3087,N_3003);
and U6844 (N_6844,N_4723,N_3519);
nor U6845 (N_6845,N_4489,N_4015);
and U6846 (N_6846,N_5309,N_4629);
nor U6847 (N_6847,N_3479,N_3001);
or U6848 (N_6848,N_3698,N_5913);
and U6849 (N_6849,N_5452,N_5109);
nand U6850 (N_6850,N_3208,N_5104);
nand U6851 (N_6851,N_4724,N_4246);
nand U6852 (N_6852,N_4208,N_3112);
and U6853 (N_6853,N_5695,N_5476);
nand U6854 (N_6854,N_4296,N_4346);
nor U6855 (N_6855,N_4355,N_3298);
or U6856 (N_6856,N_4185,N_3074);
or U6857 (N_6857,N_5982,N_4880);
xnor U6858 (N_6858,N_4074,N_5781);
nor U6859 (N_6859,N_3334,N_5687);
or U6860 (N_6860,N_5872,N_5304);
or U6861 (N_6861,N_3226,N_5352);
nor U6862 (N_6862,N_5006,N_4392);
or U6863 (N_6863,N_4937,N_3793);
nand U6864 (N_6864,N_4095,N_5535);
or U6865 (N_6865,N_3120,N_5700);
nor U6866 (N_6866,N_3201,N_5055);
nor U6867 (N_6867,N_4994,N_3163);
nand U6868 (N_6868,N_5948,N_5107);
nor U6869 (N_6869,N_3739,N_3379);
and U6870 (N_6870,N_4826,N_5065);
nand U6871 (N_6871,N_3576,N_5524);
xor U6872 (N_6872,N_3136,N_4980);
nand U6873 (N_6873,N_5388,N_5997);
or U6874 (N_6874,N_4240,N_3270);
or U6875 (N_6875,N_5053,N_4686);
nand U6876 (N_6876,N_4131,N_3331);
nor U6877 (N_6877,N_4213,N_4255);
nand U6878 (N_6878,N_5826,N_5194);
or U6879 (N_6879,N_5004,N_4657);
nor U6880 (N_6880,N_5262,N_5414);
nor U6881 (N_6881,N_3268,N_3714);
xor U6882 (N_6882,N_4675,N_3781);
and U6883 (N_6883,N_3309,N_3019);
xnor U6884 (N_6884,N_4025,N_5032);
nand U6885 (N_6885,N_5197,N_4461);
nor U6886 (N_6886,N_3752,N_4536);
nor U6887 (N_6887,N_3254,N_5792);
or U6888 (N_6888,N_5626,N_5890);
xor U6889 (N_6889,N_4884,N_3140);
nand U6890 (N_6890,N_3089,N_3606);
nand U6891 (N_6891,N_3174,N_3723);
nor U6892 (N_6892,N_5294,N_4193);
and U6893 (N_6893,N_3138,N_3614);
nor U6894 (N_6894,N_5456,N_3567);
xnor U6895 (N_6895,N_4711,N_3934);
or U6896 (N_6896,N_4196,N_5847);
or U6897 (N_6897,N_3301,N_5773);
and U6898 (N_6898,N_5871,N_5882);
nor U6899 (N_6899,N_4181,N_4353);
and U6900 (N_6900,N_3318,N_4412);
nor U6901 (N_6901,N_4485,N_4779);
nor U6902 (N_6902,N_4743,N_5521);
or U6903 (N_6903,N_3901,N_5149);
xor U6904 (N_6904,N_3098,N_3756);
nand U6905 (N_6905,N_5998,N_5449);
xor U6906 (N_6906,N_5525,N_3826);
nand U6907 (N_6907,N_5556,N_5799);
nand U6908 (N_6908,N_3463,N_4006);
or U6909 (N_6909,N_3797,N_4736);
or U6910 (N_6910,N_3819,N_4238);
nand U6911 (N_6911,N_5182,N_4496);
or U6912 (N_6912,N_3751,N_3750);
xnor U6913 (N_6913,N_5413,N_5362);
and U6914 (N_6914,N_3740,N_3371);
nand U6915 (N_6915,N_4060,N_4259);
nand U6916 (N_6916,N_5712,N_4273);
nand U6917 (N_6917,N_5511,N_3491);
nand U6918 (N_6918,N_4897,N_3456);
nand U6919 (N_6919,N_5935,N_5363);
nand U6920 (N_6920,N_3789,N_4364);
nor U6921 (N_6921,N_5324,N_4965);
and U6922 (N_6922,N_5406,N_3142);
nor U6923 (N_6923,N_5250,N_4656);
nand U6924 (N_6924,N_4241,N_3242);
or U6925 (N_6925,N_4770,N_5426);
or U6926 (N_6926,N_5912,N_4339);
nor U6927 (N_6927,N_4302,N_4159);
nand U6928 (N_6928,N_3688,N_3498);
and U6929 (N_6929,N_5435,N_5775);
and U6930 (N_6930,N_5709,N_4672);
nand U6931 (N_6931,N_3438,N_4232);
and U6932 (N_6932,N_4609,N_5724);
nor U6933 (N_6933,N_5155,N_3638);
nand U6934 (N_6934,N_3020,N_3440);
nor U6935 (N_6935,N_3538,N_4148);
nor U6936 (N_6936,N_4094,N_4712);
or U6937 (N_6937,N_3860,N_5946);
nand U6938 (N_6938,N_3807,N_4160);
and U6939 (N_6939,N_4616,N_3897);
nor U6940 (N_6940,N_5192,N_3240);
nor U6941 (N_6941,N_5277,N_4320);
nor U6942 (N_6942,N_5089,N_4342);
nand U6943 (N_6943,N_5512,N_3235);
and U6944 (N_6944,N_3984,N_5955);
or U6945 (N_6945,N_4051,N_3029);
or U6946 (N_6946,N_3566,N_5896);
and U6947 (N_6947,N_5820,N_4452);
and U6948 (N_6948,N_4757,N_5692);
nor U6949 (N_6949,N_4535,N_3765);
xnor U6950 (N_6950,N_4636,N_4118);
or U6951 (N_6951,N_3712,N_3116);
xnor U6952 (N_6952,N_4781,N_5823);
and U6953 (N_6953,N_3461,N_3153);
nor U6954 (N_6954,N_3449,N_4622);
nand U6955 (N_6955,N_3429,N_4653);
nand U6956 (N_6956,N_5341,N_4575);
or U6957 (N_6957,N_4900,N_5232);
nor U6958 (N_6958,N_4775,N_5587);
or U6959 (N_6959,N_5931,N_5332);
xor U6960 (N_6960,N_4340,N_4788);
nor U6961 (N_6961,N_3151,N_4623);
and U6962 (N_6962,N_4995,N_4854);
nand U6963 (N_6963,N_5679,N_4330);
nor U6964 (N_6964,N_4729,N_3085);
and U6965 (N_6965,N_5177,N_3528);
or U6966 (N_6966,N_4796,N_3015);
nand U6967 (N_6967,N_4648,N_5848);
nor U6968 (N_6968,N_5318,N_3317);
nor U6969 (N_6969,N_4759,N_3806);
nand U6970 (N_6970,N_3460,N_5504);
nor U6971 (N_6971,N_3591,N_5432);
xor U6972 (N_6972,N_3143,N_5497);
nor U6973 (N_6973,N_4189,N_3501);
or U6974 (N_6974,N_5927,N_4479);
nor U6975 (N_6975,N_3885,N_4426);
or U6976 (N_6976,N_4669,N_3459);
xnor U6977 (N_6977,N_4312,N_5717);
nand U6978 (N_6978,N_4113,N_3585);
nand U6979 (N_6979,N_3687,N_5330);
nor U6980 (N_6980,N_3064,N_3308);
and U6981 (N_6981,N_3180,N_3759);
nand U6982 (N_6982,N_3059,N_5204);
and U6983 (N_6983,N_4734,N_3406);
nand U6984 (N_6984,N_5145,N_5256);
nand U6985 (N_6985,N_3351,N_3384);
or U6986 (N_6986,N_3179,N_4360);
and U6987 (N_6987,N_4072,N_3804);
xor U6988 (N_6988,N_3672,N_3266);
or U6989 (N_6989,N_4579,N_4057);
or U6990 (N_6990,N_4122,N_5576);
nand U6991 (N_6991,N_5023,N_5429);
and U6992 (N_6992,N_3682,N_4075);
nor U6993 (N_6993,N_5344,N_4932);
nand U6994 (N_6994,N_3238,N_5873);
nand U6995 (N_6995,N_4077,N_3409);
nand U6996 (N_6996,N_3063,N_3578);
and U6997 (N_6997,N_4627,N_3297);
nor U6998 (N_6998,N_5647,N_5718);
or U6999 (N_6999,N_5972,N_3258);
nand U7000 (N_7000,N_4043,N_3537);
nand U7001 (N_7001,N_4644,N_3579);
nor U7002 (N_7002,N_3997,N_5658);
or U7003 (N_7003,N_5029,N_5754);
xor U7004 (N_7004,N_5484,N_5908);
nor U7005 (N_7005,N_4484,N_4190);
xnor U7006 (N_7006,N_5808,N_4191);
or U7007 (N_7007,N_4274,N_4135);
nand U7008 (N_7008,N_3025,N_3588);
nand U7009 (N_7009,N_4578,N_5039);
nand U7010 (N_7010,N_4129,N_3349);
nand U7011 (N_7011,N_4944,N_4385);
and U7012 (N_7012,N_3109,N_5513);
and U7013 (N_7013,N_3433,N_4810);
nor U7014 (N_7014,N_3282,N_4111);
nor U7015 (N_7015,N_4919,N_3741);
xor U7016 (N_7016,N_4443,N_3444);
and U7017 (N_7017,N_5305,N_3467);
or U7018 (N_7018,N_4739,N_3090);
and U7019 (N_7019,N_5688,N_3126);
nor U7020 (N_7020,N_3040,N_4119);
nand U7021 (N_7021,N_5598,N_3667);
nand U7022 (N_7022,N_3352,N_5917);
nor U7023 (N_7023,N_3624,N_4923);
nor U7024 (N_7024,N_5026,N_3657);
nand U7025 (N_7025,N_3694,N_3073);
nand U7026 (N_7026,N_4464,N_4835);
and U7027 (N_7027,N_5803,N_4529);
xnor U7028 (N_7028,N_5591,N_3783);
nand U7029 (N_7029,N_3516,N_3856);
or U7030 (N_7030,N_5082,N_3848);
or U7031 (N_7031,N_5128,N_4899);
nand U7032 (N_7032,N_3046,N_3737);
or U7033 (N_7033,N_4962,N_4337);
and U7034 (N_7034,N_4663,N_3161);
or U7035 (N_7035,N_3293,N_3833);
or U7036 (N_7036,N_5714,N_5837);
nor U7037 (N_7037,N_5374,N_5659);
nor U7038 (N_7038,N_4405,N_4369);
or U7039 (N_7039,N_3830,N_3612);
or U7040 (N_7040,N_3702,N_5705);
nor U7041 (N_7041,N_4210,N_3047);
or U7042 (N_7042,N_5654,N_5674);
nor U7043 (N_7043,N_5272,N_4832);
or U7044 (N_7044,N_4539,N_3302);
and U7045 (N_7045,N_4275,N_3972);
nand U7046 (N_7046,N_5963,N_5838);
nand U7047 (N_7047,N_5785,N_5830);
or U7048 (N_7048,N_3905,N_5682);
xnor U7049 (N_7049,N_5248,N_3364);
nor U7050 (N_7050,N_3380,N_5087);
nand U7051 (N_7051,N_3485,N_5607);
or U7052 (N_7052,N_3601,N_4719);
or U7053 (N_7053,N_4037,N_5624);
nor U7054 (N_7054,N_5459,N_3207);
and U7055 (N_7055,N_4440,N_3170);
nor U7056 (N_7056,N_3131,N_4971);
and U7057 (N_7057,N_4327,N_3390);
and U7058 (N_7058,N_4126,N_3775);
and U7059 (N_7059,N_3118,N_3224);
or U7060 (N_7060,N_5734,N_3464);
and U7061 (N_7061,N_4910,N_5037);
or U7062 (N_7062,N_3122,N_4882);
and U7063 (N_7063,N_4864,N_3931);
nor U7064 (N_7064,N_3994,N_4098);
and U7065 (N_7065,N_5952,N_5655);
or U7066 (N_7066,N_5447,N_5989);
or U7067 (N_7067,N_3620,N_4154);
or U7068 (N_7068,N_5675,N_5806);
and U7069 (N_7069,N_5962,N_5196);
and U7070 (N_7070,N_5072,N_4909);
and U7071 (N_7071,N_3679,N_3065);
and U7072 (N_7072,N_3404,N_3030);
nand U7073 (N_7073,N_5924,N_3417);
and U7074 (N_7074,N_4572,N_5058);
nand U7075 (N_7075,N_4620,N_5856);
nor U7076 (N_7076,N_4309,N_3314);
nand U7077 (N_7077,N_3731,N_4268);
nand U7078 (N_7078,N_4491,N_5188);
or U7079 (N_7079,N_4397,N_4372);
nand U7080 (N_7080,N_3233,N_4424);
nor U7081 (N_7081,N_5243,N_5438);
nor U7082 (N_7082,N_4023,N_5810);
xor U7083 (N_7083,N_5725,N_4414);
nand U7084 (N_7084,N_3791,N_5764);
nand U7085 (N_7085,N_4784,N_5461);
and U7086 (N_7086,N_3392,N_3779);
nor U7087 (N_7087,N_3195,N_5660);
and U7088 (N_7088,N_3847,N_4694);
and U7089 (N_7089,N_4862,N_3146);
and U7090 (N_7090,N_3495,N_4325);
nor U7091 (N_7091,N_5984,N_4247);
nand U7092 (N_7092,N_4930,N_4301);
nand U7093 (N_7093,N_4466,N_3212);
nand U7094 (N_7094,N_3055,N_3105);
nand U7095 (N_7095,N_4721,N_5347);
or U7096 (N_7096,N_5125,N_5236);
or U7097 (N_7097,N_3343,N_5778);
and U7098 (N_7098,N_3035,N_5861);
and U7099 (N_7099,N_5980,N_3303);
nor U7100 (N_7100,N_4483,N_3974);
nor U7101 (N_7101,N_5398,N_3773);
nor U7102 (N_7102,N_5903,N_3692);
or U7103 (N_7103,N_5317,N_4843);
or U7104 (N_7104,N_4007,N_3353);
or U7105 (N_7105,N_5615,N_5561);
nor U7106 (N_7106,N_3256,N_5000);
and U7107 (N_7107,N_5289,N_4704);
and U7108 (N_7108,N_3593,N_4918);
nand U7109 (N_7109,N_4012,N_4753);
and U7110 (N_7110,N_4744,N_5031);
nor U7111 (N_7111,N_5343,N_4099);
nor U7112 (N_7112,N_5685,N_4256);
nor U7113 (N_7113,N_3326,N_4540);
nor U7114 (N_7114,N_4363,N_5602);
nor U7115 (N_7115,N_3831,N_3362);
and U7116 (N_7116,N_5614,N_5749);
nand U7117 (N_7117,N_3094,N_4777);
and U7118 (N_7118,N_4016,N_3892);
xor U7119 (N_7119,N_5973,N_3884);
nand U7120 (N_7120,N_4270,N_5527);
nor U7121 (N_7121,N_5690,N_5092);
xor U7122 (N_7122,N_4683,N_5285);
nand U7123 (N_7123,N_4799,N_5925);
or U7124 (N_7124,N_4879,N_5396);
nand U7125 (N_7125,N_4143,N_4818);
or U7126 (N_7126,N_5409,N_3005);
nor U7127 (N_7127,N_4352,N_5209);
or U7128 (N_7128,N_3561,N_4252);
nor U7129 (N_7129,N_3300,N_4272);
nand U7130 (N_7130,N_3399,N_3785);
xor U7131 (N_7131,N_4641,N_5327);
nor U7132 (N_7132,N_5950,N_3246);
nand U7133 (N_7133,N_4615,N_3895);
or U7134 (N_7134,N_5028,N_3841);
nor U7135 (N_7135,N_5210,N_4795);
xnor U7136 (N_7136,N_3991,N_4293);
nand U7137 (N_7137,N_5689,N_5439);
or U7138 (N_7138,N_3642,N_5223);
or U7139 (N_7139,N_4202,N_4503);
and U7140 (N_7140,N_5144,N_4147);
nand U7141 (N_7141,N_4115,N_3589);
nor U7142 (N_7142,N_4814,N_4730);
nand U7143 (N_7143,N_3177,N_5479);
nand U7144 (N_7144,N_5843,N_4137);
or U7145 (N_7145,N_3749,N_3673);
nand U7146 (N_7146,N_3659,N_4975);
or U7147 (N_7147,N_5043,N_4695);
or U7148 (N_7148,N_3839,N_5123);
and U7149 (N_7149,N_5378,N_4958);
or U7150 (N_7150,N_3989,N_5892);
and U7151 (N_7151,N_4416,N_5853);
or U7152 (N_7152,N_3278,N_3542);
or U7153 (N_7153,N_4024,N_3075);
nor U7154 (N_7154,N_4234,N_5463);
and U7155 (N_7155,N_5442,N_3893);
and U7156 (N_7156,N_4450,N_4046);
nor U7157 (N_7157,N_4745,N_4889);
and U7158 (N_7158,N_4820,N_3933);
and U7159 (N_7159,N_3401,N_5866);
and U7160 (N_7160,N_5840,N_3021);
nand U7161 (N_7161,N_5977,N_3423);
nand U7162 (N_7162,N_5298,N_4838);
nor U7163 (N_7163,N_4423,N_4878);
and U7164 (N_7164,N_5122,N_4334);
nand U7165 (N_7165,N_5464,N_3543);
nand U7166 (N_7166,N_3091,N_4158);
nand U7167 (N_7167,N_3990,N_5097);
nand U7168 (N_7168,N_5857,N_3080);
or U7169 (N_7169,N_5183,N_4941);
or U7170 (N_7170,N_4248,N_4766);
xnor U7171 (N_7171,N_3451,N_5091);
or U7172 (N_7172,N_4105,N_3686);
or U7173 (N_7173,N_4167,N_4121);
and U7174 (N_7174,N_4904,N_4596);
nand U7175 (N_7175,N_3000,N_5911);
nand U7176 (N_7176,N_3129,N_5596);
and U7177 (N_7177,N_3942,N_3504);
nor U7178 (N_7178,N_4974,N_3462);
xor U7179 (N_7179,N_5545,N_5774);
nor U7180 (N_7180,N_4819,N_5481);
and U7181 (N_7181,N_4139,N_5600);
xor U7182 (N_7182,N_3329,N_4310);
nor U7183 (N_7183,N_3228,N_4715);
nand U7184 (N_7184,N_5229,N_5387);
xor U7185 (N_7185,N_3476,N_4698);
nor U7186 (N_7186,N_4714,N_4911);
or U7187 (N_7187,N_5603,N_3666);
and U7188 (N_7188,N_3100,N_5581);
xor U7189 (N_7189,N_4230,N_3951);
nor U7190 (N_7190,N_5719,N_3827);
nand U7191 (N_7191,N_5850,N_3223);
nand U7192 (N_7192,N_4823,N_3369);
nor U7193 (N_7193,N_5116,N_3178);
or U7194 (N_7194,N_5860,N_4156);
xnor U7195 (N_7195,N_5612,N_3609);
or U7196 (N_7196,N_3707,N_3683);
and U7197 (N_7197,N_4084,N_3092);
nor U7198 (N_7198,N_5800,N_4462);
and U7199 (N_7199,N_4261,N_3639);
nand U7200 (N_7200,N_5222,N_5100);
or U7201 (N_7201,N_5022,N_4034);
and U7202 (N_7202,N_3216,N_5322);
or U7203 (N_7203,N_3684,N_4673);
nor U7204 (N_7204,N_3726,N_4388);
xor U7205 (N_7205,N_5467,N_5287);
and U7206 (N_7206,N_4490,N_3144);
nor U7207 (N_7207,N_4774,N_5702);
nand U7208 (N_7208,N_4209,N_3194);
or U7209 (N_7209,N_4863,N_3536);
and U7210 (N_7210,N_4619,N_4104);
nand U7211 (N_7211,N_3800,N_4008);
nand U7212 (N_7212,N_5169,N_4417);
nand U7213 (N_7213,N_4964,N_4876);
or U7214 (N_7214,N_5844,N_5502);
nor U7215 (N_7215,N_3533,N_5025);
and U7216 (N_7216,N_3121,N_3908);
nor U7217 (N_7217,N_3843,N_5981);
or U7218 (N_7218,N_3711,N_5708);
and U7219 (N_7219,N_4231,N_5978);
nand U7220 (N_7220,N_3032,N_4380);
xor U7221 (N_7221,N_3858,N_3335);
and U7222 (N_7222,N_3577,N_3465);
xor U7223 (N_7223,N_3245,N_4707);
nor U7224 (N_7224,N_5819,N_4822);
nor U7225 (N_7225,N_5505,N_5894);
xor U7226 (N_7226,N_3734,N_5382);
nand U7227 (N_7227,N_3507,N_4091);
nand U7228 (N_7228,N_3069,N_4451);
and U7229 (N_7229,N_5595,N_3562);
nand U7230 (N_7230,N_4220,N_4688);
and U7231 (N_7231,N_4161,N_3249);
and U7232 (N_7232,N_3957,N_3940);
nor U7233 (N_7233,N_3662,N_3786);
or U7234 (N_7234,N_5707,N_3879);
nor U7235 (N_7235,N_3978,N_3037);
or U7236 (N_7236,N_3890,N_5150);
nand U7237 (N_7237,N_5743,N_3347);
or U7238 (N_7238,N_4505,N_3917);
nor U7239 (N_7239,N_3128,N_4445);
nand U7240 (N_7240,N_4970,N_4831);
nor U7241 (N_7241,N_5044,N_5669);
xnor U7242 (N_7242,N_5392,N_4912);
nand U7243 (N_7243,N_3971,N_5263);
nor U7244 (N_7244,N_5446,N_4080);
nor U7245 (N_7245,N_4260,N_5468);
or U7246 (N_7246,N_4618,N_4762);
and U7247 (N_7247,N_3442,N_3722);
or U7248 (N_7248,N_5836,N_5839);
and U7249 (N_7249,N_5986,N_3554);
nor U7250 (N_7250,N_4040,N_4480);
nor U7251 (N_7251,N_4956,N_3164);
nor U7252 (N_7252,N_5731,N_5168);
xnor U7253 (N_7253,N_3912,N_5113);
xor U7254 (N_7254,N_3042,N_5876);
or U7255 (N_7255,N_3531,N_3611);
nor U7256 (N_7256,N_5933,N_3580);
or U7257 (N_7257,N_5083,N_5656);
nand U7258 (N_7258,N_5744,N_5050);
and U7259 (N_7259,N_4116,N_3327);
and U7260 (N_7260,N_5419,N_4634);
and U7261 (N_7261,N_5126,N_3801);
or U7262 (N_7262,N_4071,N_3284);
or U7263 (N_7263,N_4170,N_5590);
nor U7264 (N_7264,N_4922,N_3982);
nor U7265 (N_7265,N_4890,N_3652);
or U7266 (N_7266,N_3656,N_5574);
xnor U7267 (N_7267,N_3628,N_3135);
and U7268 (N_7268,N_4926,N_4645);
nand U7269 (N_7269,N_5108,N_4379);
nand U7270 (N_7270,N_5763,N_4269);
nor U7271 (N_7271,N_3902,N_5329);
nor U7272 (N_7272,N_5893,N_3191);
nand U7273 (N_7273,N_3209,N_4344);
and U7274 (N_7274,N_3017,N_5001);
or U7275 (N_7275,N_5470,N_5471);
nor U7276 (N_7276,N_4017,N_3378);
nor U7277 (N_7277,N_3924,N_4727);
xnor U7278 (N_7278,N_3903,N_4969);
xor U7279 (N_7279,N_5739,N_4905);
xnor U7280 (N_7280,N_5852,N_4561);
and U7281 (N_7281,N_3981,N_4632);
nand U7282 (N_7282,N_4482,N_3360);
nand U7283 (N_7283,N_3568,N_4494);
nor U7284 (N_7284,N_4935,N_5678);
nand U7285 (N_7285,N_4586,N_5623);
nor U7286 (N_7286,N_4194,N_4530);
or U7287 (N_7287,N_4432,N_3039);
and U7288 (N_7288,N_5599,N_5550);
nor U7289 (N_7289,N_5137,N_3373);
nor U7290 (N_7290,N_3560,N_5557);
or U7291 (N_7291,N_4216,N_3678);
nor U7292 (N_7292,N_5288,N_4841);
or U7293 (N_7293,N_5661,N_5621);
or U7294 (N_7294,N_5990,N_5571);
nor U7295 (N_7295,N_5219,N_3898);
nand U7296 (N_7296,N_3281,N_3758);
nand U7297 (N_7297,N_4338,N_4376);
xnor U7298 (N_7298,N_3961,N_4754);
nor U7299 (N_7299,N_3292,N_3296);
or U7300 (N_7300,N_4797,N_4916);
and U7301 (N_7301,N_4282,N_5358);
xnor U7302 (N_7302,N_4532,N_3851);
and U7303 (N_7303,N_5824,N_5373);
and U7304 (N_7304,N_5770,N_5804);
or U7305 (N_7305,N_5807,N_5275);
and U7306 (N_7306,N_4567,N_5165);
and U7307 (N_7307,N_4585,N_5530);
and U7308 (N_7308,N_5080,N_4082);
or U7309 (N_7309,N_3251,N_5135);
nand U7310 (N_7310,N_3535,N_5592);
nor U7311 (N_7311,N_3513,N_4559);
or U7312 (N_7312,N_4515,N_4331);
nor U7313 (N_7313,N_4604,N_4875);
nor U7314 (N_7314,N_5577,N_5944);
and U7315 (N_7315,N_3034,N_4895);
nor U7316 (N_7316,N_3932,N_4387);
nand U7317 (N_7317,N_3906,N_3250);
nor U7318 (N_7318,N_5631,N_3016);
or U7319 (N_7319,N_5410,N_4545);
nand U7320 (N_7320,N_4028,N_3641);
or U7321 (N_7321,N_3980,N_5583);
nor U7322 (N_7322,N_4164,N_3496);
nor U7323 (N_7323,N_5672,N_3340);
and U7324 (N_7324,N_5851,N_4580);
and U7325 (N_7325,N_5565,N_4411);
nor U7326 (N_7326,N_3155,N_3881);
and U7327 (N_7327,N_3093,N_5105);
nor U7328 (N_7328,N_3936,N_4054);
nor U7329 (N_7329,N_5520,N_4787);
nand U7330 (N_7330,N_5281,N_4403);
or U7331 (N_7331,N_5976,N_3539);
nor U7332 (N_7332,N_5278,N_5802);
nand U7333 (N_7333,N_5680,N_3366);
and U7334 (N_7334,N_3874,N_5827);
nand U7335 (N_7335,N_5640,N_4844);
nand U7336 (N_7336,N_5652,N_4263);
nand U7337 (N_7337,N_4000,N_3383);
or U7338 (N_7338,N_3865,N_5264);
nor U7339 (N_7339,N_4289,N_4078);
and U7340 (N_7340,N_3938,N_5440);
and U7341 (N_7341,N_5441,N_4398);
nor U7342 (N_7342,N_5383,N_3668);
nor U7343 (N_7343,N_3348,N_4279);
nand U7344 (N_7344,N_4052,N_4090);
nand U7345 (N_7345,N_5411,N_3291);
nor U7346 (N_7346,N_5813,N_4557);
or U7347 (N_7347,N_4947,N_4449);
xnor U7348 (N_7348,N_5274,N_4945);
or U7349 (N_7349,N_4305,N_3716);
and U7350 (N_7350,N_3514,N_5427);
nand U7351 (N_7351,N_5834,N_4857);
and U7352 (N_7352,N_5180,N_3044);
nor U7353 (N_7353,N_4146,N_4203);
and U7354 (N_7354,N_5507,N_4061);
or U7355 (N_7355,N_3880,N_5677);
nand U7356 (N_7356,N_5490,N_3486);
nand U7357 (N_7357,N_3808,N_3387);
nand U7358 (N_7358,N_3623,N_4065);
xor U7359 (N_7359,N_4083,N_5671);
or U7360 (N_7360,N_5118,N_5995);
nand U7361 (N_7361,N_5891,N_4039);
nor U7362 (N_7362,N_5156,N_4898);
nor U7363 (N_7363,N_4807,N_5548);
and U7364 (N_7364,N_3545,N_5987);
or U7365 (N_7365,N_5110,N_4280);
nor U7366 (N_7366,N_3992,N_5966);
nand U7367 (N_7367,N_4789,N_5424);
or U7368 (N_7368,N_5027,N_4253);
nand U7369 (N_7369,N_4425,N_3710);
nor U7370 (N_7370,N_4465,N_4617);
nand U7371 (N_7371,N_5261,N_4778);
nor U7372 (N_7372,N_5637,N_3872);
nor U7373 (N_7373,N_5992,N_4304);
and U7374 (N_7374,N_3359,N_4002);
nand U7375 (N_7375,N_4375,N_5796);
or U7376 (N_7376,N_4142,N_4528);
xor U7377 (N_7377,N_3264,N_5883);
and U7378 (N_7378,N_3499,N_4637);
and U7379 (N_7379,N_3176,N_4172);
and U7380 (N_7380,N_4029,N_4354);
and U7381 (N_7381,N_5178,N_5916);
nor U7382 (N_7382,N_5696,N_3916);
xor U7383 (N_7383,N_3494,N_3066);
or U7384 (N_7384,N_4855,N_4671);
nand U7385 (N_7385,N_4501,N_4294);
and U7386 (N_7386,N_5553,N_5742);
or U7387 (N_7387,N_4176,N_3443);
or U7388 (N_7388,N_3713,N_4677);
nor U7389 (N_7389,N_3844,N_3541);
and U7390 (N_7390,N_3979,N_4128);
nor U7391 (N_7391,N_5975,N_5645);
and U7392 (N_7392,N_5153,N_3748);
or U7393 (N_7393,N_5673,N_5230);
and U7394 (N_7394,N_4149,N_4498);
nor U7395 (N_7395,N_5697,N_3923);
or U7396 (N_7396,N_5365,N_4431);
or U7397 (N_7397,N_4235,N_5706);
or U7398 (N_7398,N_5254,N_3582);
or U7399 (N_7399,N_5683,N_5821);
and U7400 (N_7400,N_3487,N_4371);
or U7401 (N_7401,N_5643,N_5606);
and U7402 (N_7402,N_5904,N_5833);
xor U7403 (N_7403,N_5005,N_3124);
nand U7404 (N_7404,N_3295,N_3198);
xnor U7405 (N_7405,N_4311,N_3203);
or U7406 (N_7406,N_3744,N_3041);
and U7407 (N_7407,N_5353,N_5012);
and U7408 (N_7408,N_3397,N_5831);
or U7409 (N_7409,N_4987,N_4347);
or U7410 (N_7410,N_3071,N_3480);
nand U7411 (N_7411,N_5457,N_3038);
or U7412 (N_7412,N_3720,N_3550);
and U7413 (N_7413,N_5385,N_5829);
nand U7414 (N_7414,N_4902,N_4689);
and U7415 (N_7415,N_3315,N_5421);
nand U7416 (N_7416,N_5176,N_3691);
xnor U7417 (N_7417,N_5306,N_3648);
nor U7418 (N_7418,N_3653,N_4662);
nand U7419 (N_7419,N_5506,N_4867);
nand U7420 (N_7420,N_3053,N_3332);
nand U7421 (N_7421,N_5013,N_5245);
nand U7422 (N_7422,N_4316,N_5212);
nand U7423 (N_7423,N_3909,N_4525);
nor U7424 (N_7424,N_3453,N_4100);
or U7425 (N_7425,N_4374,N_3426);
nor U7426 (N_7426,N_5611,N_3954);
nand U7427 (N_7427,N_4201,N_4106);
and U7428 (N_7428,N_5430,N_4599);
nand U7429 (N_7429,N_4513,N_5686);
nand U7430 (N_7430,N_5211,N_3818);
or U7431 (N_7431,N_4508,N_3483);
nand U7432 (N_7432,N_4628,N_3257);
xnor U7433 (N_7433,N_5887,N_4748);
or U7434 (N_7434,N_3402,N_5367);
nor U7435 (N_7435,N_3581,N_5252);
xor U7436 (N_7436,N_3674,N_4915);
or U7437 (N_7437,N_4506,N_4021);
and U7438 (N_7438,N_4492,N_3825);
nor U7439 (N_7439,N_3732,N_4993);
nor U7440 (N_7440,N_3421,N_5473);
or U7441 (N_7441,N_3307,N_4244);
nor U7442 (N_7442,N_3095,N_3023);
xnor U7443 (N_7443,N_4568,N_4594);
nor U7444 (N_7444,N_4174,N_5021);
and U7445 (N_7445,N_4621,N_4846);
and U7446 (N_7446,N_3134,N_5331);
or U7447 (N_7447,N_3799,N_5750);
nor U7448 (N_7448,N_4242,N_3473);
or U7449 (N_7449,N_4951,N_5328);
nand U7450 (N_7450,N_5662,N_4659);
and U7451 (N_7451,N_3663,N_4866);
nor U7452 (N_7452,N_5901,N_3549);
xnor U7453 (N_7453,N_3629,N_3771);
and U7454 (N_7454,N_4893,N_3949);
nand U7455 (N_7455,N_4651,N_4069);
xor U7456 (N_7456,N_5163,N_3400);
xor U7457 (N_7457,N_5208,N_3389);
nor U7458 (N_7458,N_3482,N_4036);
xor U7459 (N_7459,N_3468,N_4996);
xnor U7460 (N_7460,N_5273,N_5213);
and U7461 (N_7461,N_5752,N_3857);
nand U7462 (N_7462,N_5286,N_3920);
or U7463 (N_7463,N_3119,N_3605);
and U7464 (N_7464,N_4042,N_5494);
or U7465 (N_7465,N_3145,N_5737);
or U7466 (N_7466,N_4227,N_5417);
nand U7467 (N_7467,N_5760,N_4769);
nor U7468 (N_7468,N_4650,N_3488);
or U7469 (N_7469,N_3814,N_3515);
nor U7470 (N_7470,N_3729,N_3563);
or U7471 (N_7471,N_3840,N_5794);
nand U7472 (N_7472,N_3607,N_5399);
nor U7473 (N_7473,N_3500,N_4859);
or U7474 (N_7474,N_5336,N_3855);
nor U7475 (N_7475,N_5345,N_3222);
nand U7476 (N_7476,N_5167,N_5880);
or U7477 (N_7477,N_5173,N_3796);
or U7478 (N_7478,N_5564,N_4435);
xor U7479 (N_7479,N_5237,N_3132);
nor U7480 (N_7480,N_4538,N_3996);
nor U7481 (N_7481,N_5042,N_3870);
nand U7482 (N_7482,N_3333,N_4661);
and U7483 (N_7483,N_3572,N_3493);
nand U7484 (N_7484,N_4640,N_3271);
nand U7485 (N_7485,N_4033,N_5214);
xor U7486 (N_7486,N_3616,N_3061);
nor U7487 (N_7487,N_4341,N_4749);
nor U7488 (N_7488,N_4546,N_3705);
nor U7489 (N_7489,N_3220,N_5095);
or U7490 (N_7490,N_3106,N_5099);
nand U7491 (N_7491,N_3845,N_4295);
or U7492 (N_7492,N_3887,N_4531);
and U7493 (N_7493,N_5290,N_5895);
and U7494 (N_7494,N_5812,N_4109);
nor U7495 (N_7495,N_3506,N_4551);
or U7496 (N_7496,N_4569,N_3891);
nand U7497 (N_7497,N_3776,N_3634);
nor U7498 (N_7498,N_3869,N_5558);
nand U7499 (N_7499,N_5433,N_4114);
and U7500 (N_7500,N_5605,N_4359);
and U7501 (N_7501,N_5385,N_3324);
nor U7502 (N_7502,N_4575,N_4253);
or U7503 (N_7503,N_5340,N_4648);
and U7504 (N_7504,N_4566,N_3013);
nand U7505 (N_7505,N_4798,N_3339);
nor U7506 (N_7506,N_4616,N_3506);
or U7507 (N_7507,N_4015,N_3158);
and U7508 (N_7508,N_5027,N_3193);
nor U7509 (N_7509,N_4301,N_5087);
nor U7510 (N_7510,N_5279,N_3631);
nand U7511 (N_7511,N_5682,N_4946);
nand U7512 (N_7512,N_4856,N_4098);
nor U7513 (N_7513,N_5870,N_5134);
or U7514 (N_7514,N_3861,N_3689);
and U7515 (N_7515,N_5057,N_4557);
xor U7516 (N_7516,N_5992,N_4425);
or U7517 (N_7517,N_5383,N_3097);
or U7518 (N_7518,N_5666,N_4797);
xnor U7519 (N_7519,N_3652,N_4571);
or U7520 (N_7520,N_4621,N_3777);
nor U7521 (N_7521,N_4126,N_5578);
xor U7522 (N_7522,N_3724,N_3682);
nand U7523 (N_7523,N_5692,N_3220);
or U7524 (N_7524,N_5865,N_5784);
nor U7525 (N_7525,N_5508,N_4008);
or U7526 (N_7526,N_5927,N_5782);
nand U7527 (N_7527,N_4926,N_4163);
nor U7528 (N_7528,N_4678,N_5448);
xor U7529 (N_7529,N_3502,N_3059);
nand U7530 (N_7530,N_5935,N_4090);
xor U7531 (N_7531,N_5439,N_4482);
xor U7532 (N_7532,N_4920,N_5473);
nor U7533 (N_7533,N_3669,N_4128);
or U7534 (N_7534,N_5112,N_5012);
nor U7535 (N_7535,N_4149,N_3355);
xor U7536 (N_7536,N_3417,N_4669);
nor U7537 (N_7537,N_3738,N_3583);
nand U7538 (N_7538,N_4764,N_5767);
nand U7539 (N_7539,N_4564,N_4930);
nand U7540 (N_7540,N_3472,N_5712);
xnor U7541 (N_7541,N_5540,N_3167);
or U7542 (N_7542,N_5874,N_3920);
nand U7543 (N_7543,N_5363,N_3104);
and U7544 (N_7544,N_5214,N_3811);
nor U7545 (N_7545,N_3442,N_5138);
or U7546 (N_7546,N_3840,N_3979);
or U7547 (N_7547,N_5139,N_3510);
xnor U7548 (N_7548,N_5818,N_4487);
or U7549 (N_7549,N_3019,N_3033);
or U7550 (N_7550,N_5460,N_3675);
xnor U7551 (N_7551,N_4648,N_3776);
nor U7552 (N_7552,N_5286,N_5996);
or U7553 (N_7553,N_4550,N_5875);
nor U7554 (N_7554,N_3727,N_5433);
or U7555 (N_7555,N_3042,N_5088);
and U7556 (N_7556,N_3416,N_4748);
nand U7557 (N_7557,N_4513,N_4176);
nand U7558 (N_7558,N_4475,N_5831);
nand U7559 (N_7559,N_5414,N_4702);
xnor U7560 (N_7560,N_5066,N_5415);
nor U7561 (N_7561,N_5218,N_5824);
and U7562 (N_7562,N_5301,N_3159);
nand U7563 (N_7563,N_3804,N_4776);
nor U7564 (N_7564,N_5646,N_5304);
and U7565 (N_7565,N_3309,N_3803);
and U7566 (N_7566,N_5500,N_3589);
nand U7567 (N_7567,N_4053,N_5383);
nand U7568 (N_7568,N_3501,N_4436);
xor U7569 (N_7569,N_4501,N_4674);
and U7570 (N_7570,N_5526,N_4548);
or U7571 (N_7571,N_5809,N_4293);
xor U7572 (N_7572,N_3653,N_3426);
or U7573 (N_7573,N_4836,N_4766);
xor U7574 (N_7574,N_4590,N_5460);
nand U7575 (N_7575,N_5670,N_5894);
nor U7576 (N_7576,N_4855,N_5305);
and U7577 (N_7577,N_4570,N_3116);
or U7578 (N_7578,N_5516,N_5983);
nand U7579 (N_7579,N_3652,N_4266);
or U7580 (N_7580,N_5924,N_4127);
nand U7581 (N_7581,N_4968,N_3597);
nand U7582 (N_7582,N_5433,N_3513);
or U7583 (N_7583,N_3307,N_5828);
nand U7584 (N_7584,N_3787,N_5873);
or U7585 (N_7585,N_4408,N_4719);
and U7586 (N_7586,N_3093,N_5692);
nor U7587 (N_7587,N_3721,N_3298);
or U7588 (N_7588,N_4268,N_4789);
and U7589 (N_7589,N_5319,N_5438);
nand U7590 (N_7590,N_3793,N_3494);
xor U7591 (N_7591,N_5366,N_3457);
xor U7592 (N_7592,N_4538,N_5315);
or U7593 (N_7593,N_3733,N_5039);
or U7594 (N_7594,N_5378,N_4215);
and U7595 (N_7595,N_5978,N_5595);
and U7596 (N_7596,N_4696,N_3203);
or U7597 (N_7597,N_5131,N_3393);
or U7598 (N_7598,N_3279,N_5055);
nand U7599 (N_7599,N_3477,N_3341);
nand U7600 (N_7600,N_3982,N_3536);
nand U7601 (N_7601,N_5130,N_3783);
nand U7602 (N_7602,N_3648,N_3529);
nor U7603 (N_7603,N_4751,N_5508);
nand U7604 (N_7604,N_5050,N_4275);
nand U7605 (N_7605,N_5443,N_5057);
and U7606 (N_7606,N_4542,N_4442);
or U7607 (N_7607,N_5190,N_4354);
xnor U7608 (N_7608,N_3723,N_3631);
nand U7609 (N_7609,N_4837,N_3869);
nor U7610 (N_7610,N_5538,N_3461);
nor U7611 (N_7611,N_3796,N_4711);
nand U7612 (N_7612,N_3961,N_4957);
nand U7613 (N_7613,N_4093,N_4866);
or U7614 (N_7614,N_4517,N_4109);
or U7615 (N_7615,N_4192,N_4520);
or U7616 (N_7616,N_5740,N_4643);
or U7617 (N_7617,N_5167,N_3104);
nand U7618 (N_7618,N_3161,N_3518);
or U7619 (N_7619,N_4070,N_5181);
nor U7620 (N_7620,N_5728,N_4416);
or U7621 (N_7621,N_4732,N_4449);
nor U7622 (N_7622,N_3487,N_3873);
xor U7623 (N_7623,N_3591,N_3527);
and U7624 (N_7624,N_3707,N_4142);
or U7625 (N_7625,N_3290,N_4252);
nor U7626 (N_7626,N_5665,N_3931);
and U7627 (N_7627,N_3716,N_5989);
xor U7628 (N_7628,N_5932,N_4050);
nor U7629 (N_7629,N_5695,N_5356);
xnor U7630 (N_7630,N_4692,N_3674);
or U7631 (N_7631,N_3894,N_3142);
nand U7632 (N_7632,N_5555,N_3423);
or U7633 (N_7633,N_4388,N_3870);
nand U7634 (N_7634,N_5658,N_4679);
and U7635 (N_7635,N_4162,N_3881);
xnor U7636 (N_7636,N_4900,N_5227);
or U7637 (N_7637,N_3855,N_4333);
and U7638 (N_7638,N_4999,N_5610);
nand U7639 (N_7639,N_5867,N_4763);
or U7640 (N_7640,N_3030,N_5743);
nor U7641 (N_7641,N_3495,N_3224);
nand U7642 (N_7642,N_5425,N_4449);
nor U7643 (N_7643,N_4601,N_3056);
nor U7644 (N_7644,N_5132,N_4324);
nand U7645 (N_7645,N_3746,N_3905);
and U7646 (N_7646,N_5791,N_3394);
nor U7647 (N_7647,N_4331,N_3954);
and U7648 (N_7648,N_3128,N_4058);
nand U7649 (N_7649,N_3678,N_5886);
nand U7650 (N_7650,N_3962,N_4087);
nand U7651 (N_7651,N_3048,N_5177);
nor U7652 (N_7652,N_4888,N_4495);
xor U7653 (N_7653,N_5014,N_5105);
nor U7654 (N_7654,N_5099,N_5226);
nand U7655 (N_7655,N_3604,N_4632);
or U7656 (N_7656,N_3368,N_5546);
or U7657 (N_7657,N_5936,N_5878);
nand U7658 (N_7658,N_3829,N_4866);
nand U7659 (N_7659,N_3894,N_4323);
nand U7660 (N_7660,N_4943,N_4486);
nor U7661 (N_7661,N_3751,N_5834);
and U7662 (N_7662,N_5850,N_3732);
nand U7663 (N_7663,N_5767,N_5376);
nand U7664 (N_7664,N_4747,N_4293);
or U7665 (N_7665,N_3005,N_5522);
nand U7666 (N_7666,N_5551,N_5655);
nand U7667 (N_7667,N_3836,N_5708);
nor U7668 (N_7668,N_5053,N_3116);
nand U7669 (N_7669,N_5499,N_3422);
nand U7670 (N_7670,N_4788,N_4399);
nor U7671 (N_7671,N_5164,N_5741);
nor U7672 (N_7672,N_4925,N_4098);
or U7673 (N_7673,N_5418,N_4819);
nor U7674 (N_7674,N_5377,N_3746);
xor U7675 (N_7675,N_5070,N_4443);
nor U7676 (N_7676,N_5031,N_3130);
nand U7677 (N_7677,N_5864,N_4246);
nor U7678 (N_7678,N_4361,N_3410);
and U7679 (N_7679,N_3502,N_5776);
nor U7680 (N_7680,N_3596,N_3033);
nor U7681 (N_7681,N_3368,N_4942);
nor U7682 (N_7682,N_4226,N_4507);
nand U7683 (N_7683,N_3704,N_3280);
or U7684 (N_7684,N_3454,N_5390);
and U7685 (N_7685,N_4369,N_5068);
nor U7686 (N_7686,N_4359,N_5607);
nand U7687 (N_7687,N_4890,N_5750);
or U7688 (N_7688,N_5706,N_5268);
nand U7689 (N_7689,N_4046,N_3312);
nand U7690 (N_7690,N_4810,N_5846);
nor U7691 (N_7691,N_3688,N_4363);
nand U7692 (N_7692,N_4394,N_3462);
or U7693 (N_7693,N_5583,N_5192);
and U7694 (N_7694,N_4666,N_3026);
or U7695 (N_7695,N_3064,N_5412);
nor U7696 (N_7696,N_4295,N_3655);
nor U7697 (N_7697,N_4255,N_5991);
or U7698 (N_7698,N_5673,N_4118);
and U7699 (N_7699,N_5053,N_3371);
nand U7700 (N_7700,N_5637,N_5109);
and U7701 (N_7701,N_4476,N_3935);
nor U7702 (N_7702,N_4984,N_5579);
and U7703 (N_7703,N_5890,N_5571);
or U7704 (N_7704,N_4928,N_4434);
xnor U7705 (N_7705,N_4521,N_5424);
nand U7706 (N_7706,N_4335,N_5582);
xnor U7707 (N_7707,N_3325,N_3288);
and U7708 (N_7708,N_5113,N_5786);
nand U7709 (N_7709,N_5301,N_3541);
and U7710 (N_7710,N_3076,N_4337);
nor U7711 (N_7711,N_3521,N_5201);
nand U7712 (N_7712,N_5049,N_4327);
nor U7713 (N_7713,N_3508,N_3082);
and U7714 (N_7714,N_3189,N_3534);
nor U7715 (N_7715,N_3616,N_3146);
nor U7716 (N_7716,N_3080,N_5312);
or U7717 (N_7717,N_5086,N_5305);
and U7718 (N_7718,N_4810,N_3256);
or U7719 (N_7719,N_3499,N_5005);
nor U7720 (N_7720,N_4158,N_3297);
or U7721 (N_7721,N_5591,N_5800);
nor U7722 (N_7722,N_3055,N_4569);
xor U7723 (N_7723,N_3671,N_3330);
nand U7724 (N_7724,N_3338,N_5131);
and U7725 (N_7725,N_4907,N_4489);
or U7726 (N_7726,N_4392,N_4428);
nand U7727 (N_7727,N_3590,N_5233);
xor U7728 (N_7728,N_4270,N_4232);
nand U7729 (N_7729,N_5362,N_5304);
and U7730 (N_7730,N_4658,N_4000);
xor U7731 (N_7731,N_5628,N_5895);
nand U7732 (N_7732,N_5130,N_3547);
xnor U7733 (N_7733,N_5118,N_3444);
or U7734 (N_7734,N_3168,N_5109);
or U7735 (N_7735,N_4332,N_4429);
or U7736 (N_7736,N_3824,N_4853);
nor U7737 (N_7737,N_3006,N_4094);
or U7738 (N_7738,N_5641,N_4907);
and U7739 (N_7739,N_4612,N_5017);
and U7740 (N_7740,N_5206,N_3115);
and U7741 (N_7741,N_5725,N_5910);
nand U7742 (N_7742,N_3125,N_3650);
xnor U7743 (N_7743,N_3375,N_4939);
nand U7744 (N_7744,N_4116,N_4321);
xnor U7745 (N_7745,N_3982,N_4375);
nand U7746 (N_7746,N_5816,N_4996);
nor U7747 (N_7747,N_3815,N_4870);
and U7748 (N_7748,N_5033,N_3374);
nand U7749 (N_7749,N_5577,N_4094);
or U7750 (N_7750,N_4769,N_4501);
xnor U7751 (N_7751,N_4329,N_5046);
nand U7752 (N_7752,N_5546,N_5412);
nor U7753 (N_7753,N_3769,N_5050);
or U7754 (N_7754,N_4873,N_3561);
nor U7755 (N_7755,N_3508,N_4103);
or U7756 (N_7756,N_4858,N_5506);
nand U7757 (N_7757,N_5927,N_3869);
and U7758 (N_7758,N_3855,N_5536);
nor U7759 (N_7759,N_4460,N_4347);
nor U7760 (N_7760,N_4863,N_5380);
xor U7761 (N_7761,N_5342,N_5726);
xor U7762 (N_7762,N_5297,N_4469);
or U7763 (N_7763,N_5759,N_5603);
and U7764 (N_7764,N_5040,N_4907);
or U7765 (N_7765,N_3187,N_5043);
nor U7766 (N_7766,N_5707,N_3932);
nand U7767 (N_7767,N_3481,N_4463);
or U7768 (N_7768,N_4843,N_4386);
nand U7769 (N_7769,N_3113,N_5298);
xnor U7770 (N_7770,N_3533,N_3424);
nand U7771 (N_7771,N_5175,N_3629);
xnor U7772 (N_7772,N_3908,N_4877);
or U7773 (N_7773,N_4347,N_5038);
nand U7774 (N_7774,N_3314,N_3365);
nand U7775 (N_7775,N_5057,N_5681);
nand U7776 (N_7776,N_5584,N_4446);
or U7777 (N_7777,N_5465,N_4127);
nor U7778 (N_7778,N_5527,N_4726);
xnor U7779 (N_7779,N_4476,N_3645);
and U7780 (N_7780,N_5883,N_5417);
or U7781 (N_7781,N_5777,N_3944);
xnor U7782 (N_7782,N_5693,N_3383);
or U7783 (N_7783,N_3313,N_3481);
and U7784 (N_7784,N_4548,N_4714);
or U7785 (N_7785,N_4236,N_3655);
and U7786 (N_7786,N_5465,N_4082);
nor U7787 (N_7787,N_4761,N_5306);
nand U7788 (N_7788,N_5921,N_3348);
nand U7789 (N_7789,N_5782,N_4286);
and U7790 (N_7790,N_5460,N_5695);
and U7791 (N_7791,N_4421,N_3383);
or U7792 (N_7792,N_5043,N_4889);
nor U7793 (N_7793,N_4118,N_4980);
or U7794 (N_7794,N_3482,N_5754);
nand U7795 (N_7795,N_4855,N_3131);
and U7796 (N_7796,N_3363,N_3171);
nand U7797 (N_7797,N_3027,N_4360);
nor U7798 (N_7798,N_4464,N_3119);
xor U7799 (N_7799,N_3095,N_5947);
nand U7800 (N_7800,N_3223,N_4234);
xnor U7801 (N_7801,N_4532,N_5589);
and U7802 (N_7802,N_3967,N_5323);
or U7803 (N_7803,N_3607,N_3031);
and U7804 (N_7804,N_5855,N_3774);
or U7805 (N_7805,N_3731,N_4014);
nand U7806 (N_7806,N_3978,N_5726);
nand U7807 (N_7807,N_5600,N_4227);
nand U7808 (N_7808,N_3594,N_3237);
and U7809 (N_7809,N_3551,N_3067);
nor U7810 (N_7810,N_4568,N_4721);
or U7811 (N_7811,N_4556,N_3635);
xnor U7812 (N_7812,N_4130,N_5408);
and U7813 (N_7813,N_5064,N_3520);
or U7814 (N_7814,N_4972,N_5255);
nand U7815 (N_7815,N_3513,N_5274);
nor U7816 (N_7816,N_5016,N_3449);
or U7817 (N_7817,N_4769,N_4701);
nand U7818 (N_7818,N_3742,N_5219);
nand U7819 (N_7819,N_5209,N_4684);
and U7820 (N_7820,N_4122,N_4231);
nor U7821 (N_7821,N_5898,N_3543);
or U7822 (N_7822,N_3936,N_4521);
nor U7823 (N_7823,N_4084,N_5995);
nand U7824 (N_7824,N_4159,N_4721);
nand U7825 (N_7825,N_3899,N_4751);
and U7826 (N_7826,N_4486,N_3380);
nor U7827 (N_7827,N_4690,N_4018);
nor U7828 (N_7828,N_3130,N_4352);
xor U7829 (N_7829,N_3578,N_3071);
nand U7830 (N_7830,N_5982,N_3967);
nor U7831 (N_7831,N_3798,N_5784);
xnor U7832 (N_7832,N_3827,N_3620);
and U7833 (N_7833,N_5084,N_3373);
nor U7834 (N_7834,N_5858,N_4891);
nor U7835 (N_7835,N_5419,N_4428);
or U7836 (N_7836,N_5371,N_4012);
xor U7837 (N_7837,N_5913,N_4167);
nand U7838 (N_7838,N_5837,N_3184);
or U7839 (N_7839,N_5962,N_3808);
or U7840 (N_7840,N_5720,N_3243);
and U7841 (N_7841,N_3189,N_5761);
nand U7842 (N_7842,N_5606,N_3701);
nand U7843 (N_7843,N_3615,N_5127);
nand U7844 (N_7844,N_5247,N_3661);
and U7845 (N_7845,N_4567,N_3354);
nor U7846 (N_7846,N_5200,N_4459);
or U7847 (N_7847,N_3804,N_4632);
and U7848 (N_7848,N_4826,N_3311);
nand U7849 (N_7849,N_4089,N_3214);
nand U7850 (N_7850,N_5012,N_5026);
nand U7851 (N_7851,N_3022,N_3762);
xnor U7852 (N_7852,N_4803,N_3849);
or U7853 (N_7853,N_4313,N_3465);
xor U7854 (N_7854,N_4516,N_3995);
and U7855 (N_7855,N_5852,N_4753);
and U7856 (N_7856,N_5593,N_4296);
or U7857 (N_7857,N_4637,N_3590);
or U7858 (N_7858,N_5917,N_3346);
nor U7859 (N_7859,N_5255,N_4185);
nand U7860 (N_7860,N_4014,N_4576);
xnor U7861 (N_7861,N_4333,N_5633);
and U7862 (N_7862,N_4775,N_4885);
nand U7863 (N_7863,N_4367,N_3259);
or U7864 (N_7864,N_3952,N_4449);
or U7865 (N_7865,N_5093,N_3238);
nor U7866 (N_7866,N_3994,N_3566);
and U7867 (N_7867,N_3249,N_5510);
nand U7868 (N_7868,N_4404,N_3401);
and U7869 (N_7869,N_5152,N_5772);
nor U7870 (N_7870,N_5811,N_4591);
and U7871 (N_7871,N_5303,N_4246);
nor U7872 (N_7872,N_3561,N_5574);
nor U7873 (N_7873,N_4852,N_5209);
nor U7874 (N_7874,N_3285,N_3637);
xor U7875 (N_7875,N_4522,N_5824);
nor U7876 (N_7876,N_5662,N_5780);
and U7877 (N_7877,N_5997,N_4178);
nor U7878 (N_7878,N_5428,N_5342);
nand U7879 (N_7879,N_5529,N_3697);
and U7880 (N_7880,N_3188,N_4213);
nor U7881 (N_7881,N_5675,N_5927);
nor U7882 (N_7882,N_5202,N_3527);
nor U7883 (N_7883,N_3132,N_5586);
and U7884 (N_7884,N_3056,N_5240);
and U7885 (N_7885,N_4780,N_5744);
nand U7886 (N_7886,N_4567,N_3246);
nor U7887 (N_7887,N_5631,N_5475);
or U7888 (N_7888,N_3608,N_3776);
nand U7889 (N_7889,N_4415,N_5082);
and U7890 (N_7890,N_5842,N_4081);
and U7891 (N_7891,N_5773,N_4418);
nand U7892 (N_7892,N_4360,N_3103);
and U7893 (N_7893,N_3551,N_5498);
and U7894 (N_7894,N_5330,N_4486);
nor U7895 (N_7895,N_4001,N_5407);
nor U7896 (N_7896,N_4810,N_5095);
or U7897 (N_7897,N_5693,N_3712);
nor U7898 (N_7898,N_3547,N_5864);
and U7899 (N_7899,N_3714,N_5938);
nand U7900 (N_7900,N_3172,N_5583);
or U7901 (N_7901,N_3386,N_3434);
nand U7902 (N_7902,N_3381,N_5085);
nand U7903 (N_7903,N_5038,N_3180);
and U7904 (N_7904,N_4054,N_5884);
xor U7905 (N_7905,N_4877,N_3489);
nor U7906 (N_7906,N_5341,N_3036);
nor U7907 (N_7907,N_5919,N_4512);
or U7908 (N_7908,N_5331,N_5549);
and U7909 (N_7909,N_3875,N_3211);
nand U7910 (N_7910,N_4802,N_4650);
or U7911 (N_7911,N_4510,N_5274);
nor U7912 (N_7912,N_4652,N_5906);
and U7913 (N_7913,N_3401,N_3989);
and U7914 (N_7914,N_4511,N_5670);
or U7915 (N_7915,N_3128,N_3142);
nand U7916 (N_7916,N_3201,N_4104);
nor U7917 (N_7917,N_3982,N_3299);
nand U7918 (N_7918,N_3915,N_4921);
nand U7919 (N_7919,N_4997,N_4819);
and U7920 (N_7920,N_3429,N_3214);
xor U7921 (N_7921,N_4824,N_3621);
and U7922 (N_7922,N_4028,N_4522);
or U7923 (N_7923,N_5710,N_4219);
nor U7924 (N_7924,N_3006,N_4872);
and U7925 (N_7925,N_4245,N_5001);
nand U7926 (N_7926,N_5512,N_4750);
nand U7927 (N_7927,N_5116,N_3070);
nand U7928 (N_7928,N_4298,N_3077);
nor U7929 (N_7929,N_3023,N_4751);
or U7930 (N_7930,N_5085,N_3290);
xor U7931 (N_7931,N_3085,N_5627);
and U7932 (N_7932,N_3439,N_5815);
nor U7933 (N_7933,N_4658,N_3480);
nand U7934 (N_7934,N_4380,N_5560);
nand U7935 (N_7935,N_3671,N_3379);
nand U7936 (N_7936,N_5496,N_5912);
xor U7937 (N_7937,N_4525,N_4789);
nor U7938 (N_7938,N_3670,N_4330);
nor U7939 (N_7939,N_4237,N_5444);
xor U7940 (N_7940,N_3216,N_5082);
or U7941 (N_7941,N_5037,N_3224);
xor U7942 (N_7942,N_5494,N_4460);
or U7943 (N_7943,N_5724,N_4659);
nor U7944 (N_7944,N_3973,N_3947);
nor U7945 (N_7945,N_3429,N_5770);
or U7946 (N_7946,N_5145,N_3533);
nand U7947 (N_7947,N_4257,N_4861);
nand U7948 (N_7948,N_5629,N_4476);
nor U7949 (N_7949,N_5086,N_5351);
or U7950 (N_7950,N_4412,N_3023);
nor U7951 (N_7951,N_5077,N_4199);
nand U7952 (N_7952,N_3376,N_4094);
or U7953 (N_7953,N_5964,N_4939);
nand U7954 (N_7954,N_4421,N_3251);
nor U7955 (N_7955,N_5457,N_4631);
or U7956 (N_7956,N_5335,N_3798);
and U7957 (N_7957,N_3809,N_4515);
nand U7958 (N_7958,N_5406,N_3271);
nor U7959 (N_7959,N_3956,N_3695);
nor U7960 (N_7960,N_5853,N_3601);
or U7961 (N_7961,N_3342,N_3835);
or U7962 (N_7962,N_3646,N_5744);
xor U7963 (N_7963,N_3407,N_3092);
or U7964 (N_7964,N_3400,N_3660);
xnor U7965 (N_7965,N_5462,N_3996);
nand U7966 (N_7966,N_4469,N_4601);
nor U7967 (N_7967,N_4077,N_3543);
or U7968 (N_7968,N_3072,N_5233);
and U7969 (N_7969,N_3683,N_3780);
nor U7970 (N_7970,N_5076,N_5421);
or U7971 (N_7971,N_4952,N_5606);
or U7972 (N_7972,N_5167,N_3317);
or U7973 (N_7973,N_3092,N_4108);
nor U7974 (N_7974,N_4289,N_4376);
or U7975 (N_7975,N_5036,N_3556);
and U7976 (N_7976,N_5226,N_3341);
nand U7977 (N_7977,N_5500,N_5419);
nand U7978 (N_7978,N_3610,N_5884);
xnor U7979 (N_7979,N_5966,N_3384);
nor U7980 (N_7980,N_4810,N_3797);
or U7981 (N_7981,N_4328,N_4021);
or U7982 (N_7982,N_3445,N_4381);
and U7983 (N_7983,N_4504,N_4251);
nand U7984 (N_7984,N_4855,N_4626);
and U7985 (N_7985,N_5424,N_4624);
nor U7986 (N_7986,N_5688,N_5292);
and U7987 (N_7987,N_4807,N_3922);
nor U7988 (N_7988,N_3509,N_5999);
nor U7989 (N_7989,N_5299,N_4916);
and U7990 (N_7990,N_3824,N_3580);
and U7991 (N_7991,N_4344,N_5708);
xor U7992 (N_7992,N_5134,N_3493);
nand U7993 (N_7993,N_4381,N_5986);
nor U7994 (N_7994,N_4932,N_5905);
or U7995 (N_7995,N_3128,N_3348);
nor U7996 (N_7996,N_4761,N_4845);
nor U7997 (N_7997,N_3608,N_5764);
nor U7998 (N_7998,N_4429,N_3391);
or U7999 (N_7999,N_4408,N_5108);
xor U8000 (N_8000,N_4690,N_5242);
and U8001 (N_8001,N_3571,N_4093);
or U8002 (N_8002,N_4838,N_5895);
xor U8003 (N_8003,N_3812,N_3907);
nand U8004 (N_8004,N_3715,N_5082);
and U8005 (N_8005,N_4737,N_5163);
nor U8006 (N_8006,N_3249,N_4776);
nand U8007 (N_8007,N_4304,N_5806);
nor U8008 (N_8008,N_5940,N_5116);
xnor U8009 (N_8009,N_4093,N_3885);
nand U8010 (N_8010,N_3276,N_5074);
and U8011 (N_8011,N_3260,N_3375);
nor U8012 (N_8012,N_3554,N_5863);
nand U8013 (N_8013,N_5059,N_3823);
or U8014 (N_8014,N_4441,N_5373);
or U8015 (N_8015,N_5720,N_4920);
or U8016 (N_8016,N_4189,N_5010);
and U8017 (N_8017,N_5944,N_3858);
or U8018 (N_8018,N_5150,N_5215);
or U8019 (N_8019,N_4621,N_3355);
xor U8020 (N_8020,N_3136,N_4830);
xnor U8021 (N_8021,N_4483,N_3857);
nor U8022 (N_8022,N_4215,N_3038);
nand U8023 (N_8023,N_4795,N_5336);
xnor U8024 (N_8024,N_5777,N_5304);
nand U8025 (N_8025,N_4219,N_5934);
or U8026 (N_8026,N_5784,N_3487);
or U8027 (N_8027,N_3928,N_5664);
nor U8028 (N_8028,N_5725,N_4479);
and U8029 (N_8029,N_3748,N_4022);
nand U8030 (N_8030,N_5441,N_3792);
nand U8031 (N_8031,N_5876,N_5575);
nor U8032 (N_8032,N_5366,N_4613);
nor U8033 (N_8033,N_4342,N_3225);
and U8034 (N_8034,N_4815,N_4040);
nor U8035 (N_8035,N_3805,N_3474);
and U8036 (N_8036,N_5212,N_5024);
and U8037 (N_8037,N_4590,N_4148);
and U8038 (N_8038,N_5910,N_4371);
nor U8039 (N_8039,N_4327,N_3098);
nor U8040 (N_8040,N_5779,N_3316);
nor U8041 (N_8041,N_5607,N_3032);
nor U8042 (N_8042,N_3924,N_4955);
nor U8043 (N_8043,N_4395,N_4885);
or U8044 (N_8044,N_5282,N_5844);
nand U8045 (N_8045,N_4498,N_3136);
or U8046 (N_8046,N_3148,N_5548);
and U8047 (N_8047,N_3130,N_5492);
nor U8048 (N_8048,N_5429,N_3225);
or U8049 (N_8049,N_4814,N_4295);
nand U8050 (N_8050,N_3744,N_3755);
nor U8051 (N_8051,N_4210,N_3488);
nand U8052 (N_8052,N_4109,N_5546);
nand U8053 (N_8053,N_3452,N_4476);
nor U8054 (N_8054,N_5095,N_4738);
or U8055 (N_8055,N_5507,N_5218);
or U8056 (N_8056,N_4674,N_5174);
and U8057 (N_8057,N_4712,N_4885);
nor U8058 (N_8058,N_4511,N_5464);
or U8059 (N_8059,N_5598,N_3418);
or U8060 (N_8060,N_4365,N_5987);
and U8061 (N_8061,N_5340,N_5771);
or U8062 (N_8062,N_3894,N_5208);
xor U8063 (N_8063,N_5286,N_5888);
and U8064 (N_8064,N_4803,N_5105);
and U8065 (N_8065,N_4279,N_4542);
xnor U8066 (N_8066,N_4224,N_4461);
nand U8067 (N_8067,N_5910,N_4288);
nor U8068 (N_8068,N_3983,N_5677);
nor U8069 (N_8069,N_3471,N_5020);
or U8070 (N_8070,N_3361,N_5062);
xnor U8071 (N_8071,N_5648,N_4696);
and U8072 (N_8072,N_3786,N_5159);
nand U8073 (N_8073,N_4427,N_4156);
nand U8074 (N_8074,N_5118,N_5902);
nor U8075 (N_8075,N_3403,N_5158);
or U8076 (N_8076,N_3638,N_3807);
or U8077 (N_8077,N_4735,N_3057);
or U8078 (N_8078,N_4821,N_3294);
and U8079 (N_8079,N_4981,N_4463);
and U8080 (N_8080,N_3526,N_5226);
or U8081 (N_8081,N_4845,N_4443);
nand U8082 (N_8082,N_5747,N_4666);
and U8083 (N_8083,N_4652,N_5622);
or U8084 (N_8084,N_4156,N_4180);
nand U8085 (N_8085,N_3589,N_3518);
and U8086 (N_8086,N_5887,N_5879);
nand U8087 (N_8087,N_3879,N_3903);
and U8088 (N_8088,N_3379,N_3539);
and U8089 (N_8089,N_5838,N_4174);
nand U8090 (N_8090,N_5275,N_5282);
nor U8091 (N_8091,N_5892,N_3949);
and U8092 (N_8092,N_5468,N_5867);
nand U8093 (N_8093,N_3835,N_5229);
and U8094 (N_8094,N_5242,N_3042);
nand U8095 (N_8095,N_4273,N_4208);
and U8096 (N_8096,N_4944,N_4471);
nand U8097 (N_8097,N_3589,N_3519);
or U8098 (N_8098,N_4425,N_3887);
and U8099 (N_8099,N_4457,N_4975);
nand U8100 (N_8100,N_5082,N_3178);
nand U8101 (N_8101,N_5478,N_4380);
nand U8102 (N_8102,N_3174,N_5877);
nor U8103 (N_8103,N_4306,N_5422);
nor U8104 (N_8104,N_5165,N_3465);
or U8105 (N_8105,N_3816,N_3247);
nand U8106 (N_8106,N_4269,N_5161);
and U8107 (N_8107,N_5843,N_3202);
or U8108 (N_8108,N_5693,N_4334);
nor U8109 (N_8109,N_4063,N_4410);
and U8110 (N_8110,N_3227,N_5640);
and U8111 (N_8111,N_4456,N_5748);
nor U8112 (N_8112,N_5285,N_5380);
or U8113 (N_8113,N_4267,N_4317);
and U8114 (N_8114,N_3817,N_4199);
nand U8115 (N_8115,N_4485,N_3700);
nor U8116 (N_8116,N_4982,N_5037);
or U8117 (N_8117,N_4808,N_4359);
and U8118 (N_8118,N_4224,N_3658);
nor U8119 (N_8119,N_4471,N_5612);
or U8120 (N_8120,N_5155,N_3089);
nand U8121 (N_8121,N_4682,N_4584);
nand U8122 (N_8122,N_5472,N_3729);
or U8123 (N_8123,N_4413,N_3896);
nand U8124 (N_8124,N_3182,N_3772);
and U8125 (N_8125,N_4466,N_5729);
and U8126 (N_8126,N_4063,N_4430);
nand U8127 (N_8127,N_3161,N_5713);
or U8128 (N_8128,N_3607,N_3460);
and U8129 (N_8129,N_4327,N_5295);
and U8130 (N_8130,N_4778,N_4285);
nand U8131 (N_8131,N_5523,N_3179);
and U8132 (N_8132,N_3734,N_5096);
nand U8133 (N_8133,N_5388,N_3506);
nor U8134 (N_8134,N_4737,N_5038);
or U8135 (N_8135,N_3634,N_4104);
nor U8136 (N_8136,N_4943,N_5845);
or U8137 (N_8137,N_4011,N_3191);
and U8138 (N_8138,N_5930,N_3833);
nand U8139 (N_8139,N_3077,N_5551);
nor U8140 (N_8140,N_4550,N_4433);
and U8141 (N_8141,N_4071,N_4091);
and U8142 (N_8142,N_5571,N_3167);
nor U8143 (N_8143,N_3160,N_5000);
nor U8144 (N_8144,N_4075,N_4103);
nand U8145 (N_8145,N_4112,N_5327);
nand U8146 (N_8146,N_5635,N_5535);
xnor U8147 (N_8147,N_5300,N_3458);
or U8148 (N_8148,N_5956,N_5700);
or U8149 (N_8149,N_5003,N_3951);
or U8150 (N_8150,N_3347,N_5060);
or U8151 (N_8151,N_3900,N_4589);
nand U8152 (N_8152,N_4588,N_4740);
nor U8153 (N_8153,N_5686,N_3468);
nand U8154 (N_8154,N_3347,N_4379);
nand U8155 (N_8155,N_4501,N_4714);
or U8156 (N_8156,N_5204,N_4459);
nand U8157 (N_8157,N_3521,N_5511);
xnor U8158 (N_8158,N_4414,N_3458);
or U8159 (N_8159,N_4663,N_3155);
and U8160 (N_8160,N_4988,N_5457);
nor U8161 (N_8161,N_4415,N_5318);
and U8162 (N_8162,N_3466,N_3832);
and U8163 (N_8163,N_3861,N_4496);
or U8164 (N_8164,N_3870,N_3291);
nand U8165 (N_8165,N_5320,N_5641);
nand U8166 (N_8166,N_4106,N_4453);
xnor U8167 (N_8167,N_4716,N_3026);
nor U8168 (N_8168,N_3793,N_4439);
nor U8169 (N_8169,N_4474,N_4487);
nand U8170 (N_8170,N_4703,N_4073);
and U8171 (N_8171,N_5688,N_5233);
nor U8172 (N_8172,N_5952,N_3171);
and U8173 (N_8173,N_3472,N_3282);
nor U8174 (N_8174,N_3425,N_3714);
nor U8175 (N_8175,N_5637,N_5172);
and U8176 (N_8176,N_4351,N_3707);
nor U8177 (N_8177,N_3226,N_5012);
nand U8178 (N_8178,N_4720,N_5181);
or U8179 (N_8179,N_4822,N_4769);
or U8180 (N_8180,N_4010,N_5540);
and U8181 (N_8181,N_4175,N_4850);
or U8182 (N_8182,N_5831,N_4624);
xor U8183 (N_8183,N_5163,N_5113);
xor U8184 (N_8184,N_4708,N_3765);
nand U8185 (N_8185,N_5510,N_5532);
and U8186 (N_8186,N_3572,N_5340);
and U8187 (N_8187,N_3200,N_5507);
and U8188 (N_8188,N_5485,N_5290);
nand U8189 (N_8189,N_3018,N_4022);
nor U8190 (N_8190,N_4222,N_4353);
and U8191 (N_8191,N_5448,N_3932);
and U8192 (N_8192,N_5576,N_3641);
or U8193 (N_8193,N_5673,N_3673);
nand U8194 (N_8194,N_5318,N_4543);
nand U8195 (N_8195,N_3706,N_5565);
nor U8196 (N_8196,N_4075,N_5946);
or U8197 (N_8197,N_3933,N_4300);
and U8198 (N_8198,N_3415,N_5448);
and U8199 (N_8199,N_4481,N_3238);
nor U8200 (N_8200,N_5598,N_3340);
nor U8201 (N_8201,N_3042,N_4415);
and U8202 (N_8202,N_4153,N_3093);
xnor U8203 (N_8203,N_5246,N_4603);
and U8204 (N_8204,N_4497,N_5836);
or U8205 (N_8205,N_4004,N_4570);
and U8206 (N_8206,N_3301,N_5800);
or U8207 (N_8207,N_3632,N_5551);
nor U8208 (N_8208,N_4196,N_4350);
and U8209 (N_8209,N_3448,N_5371);
nor U8210 (N_8210,N_3508,N_5356);
nor U8211 (N_8211,N_4641,N_5965);
nor U8212 (N_8212,N_3576,N_3873);
nor U8213 (N_8213,N_3547,N_5845);
and U8214 (N_8214,N_5586,N_4230);
and U8215 (N_8215,N_4193,N_3158);
or U8216 (N_8216,N_5145,N_5013);
nor U8217 (N_8217,N_4522,N_4184);
nor U8218 (N_8218,N_3084,N_3896);
or U8219 (N_8219,N_5035,N_5606);
and U8220 (N_8220,N_5233,N_4601);
or U8221 (N_8221,N_3970,N_5627);
nand U8222 (N_8222,N_4509,N_3304);
xor U8223 (N_8223,N_5756,N_4811);
nor U8224 (N_8224,N_3323,N_5701);
nor U8225 (N_8225,N_5922,N_5623);
or U8226 (N_8226,N_3830,N_3634);
and U8227 (N_8227,N_5933,N_3499);
nor U8228 (N_8228,N_3763,N_5918);
nand U8229 (N_8229,N_3896,N_3643);
nor U8230 (N_8230,N_3228,N_3390);
or U8231 (N_8231,N_3240,N_5286);
xnor U8232 (N_8232,N_5293,N_4054);
nor U8233 (N_8233,N_4351,N_4278);
and U8234 (N_8234,N_3170,N_3688);
or U8235 (N_8235,N_4828,N_4670);
or U8236 (N_8236,N_3069,N_3849);
nor U8237 (N_8237,N_3180,N_3344);
nand U8238 (N_8238,N_3172,N_5561);
or U8239 (N_8239,N_4448,N_4824);
and U8240 (N_8240,N_3265,N_5984);
nor U8241 (N_8241,N_5711,N_3482);
nand U8242 (N_8242,N_5576,N_3202);
or U8243 (N_8243,N_4776,N_3853);
nand U8244 (N_8244,N_3297,N_5860);
and U8245 (N_8245,N_3322,N_4499);
nand U8246 (N_8246,N_5414,N_4626);
nor U8247 (N_8247,N_5513,N_5369);
xnor U8248 (N_8248,N_5706,N_4164);
nor U8249 (N_8249,N_3074,N_4527);
and U8250 (N_8250,N_4985,N_4607);
or U8251 (N_8251,N_4809,N_5029);
nand U8252 (N_8252,N_3215,N_3204);
nand U8253 (N_8253,N_4942,N_3033);
nor U8254 (N_8254,N_5432,N_4442);
nand U8255 (N_8255,N_4043,N_5771);
nor U8256 (N_8256,N_3876,N_4288);
nor U8257 (N_8257,N_5473,N_4856);
or U8258 (N_8258,N_4092,N_4634);
or U8259 (N_8259,N_3142,N_5588);
and U8260 (N_8260,N_3877,N_3973);
nor U8261 (N_8261,N_5522,N_5015);
xnor U8262 (N_8262,N_3260,N_4468);
nand U8263 (N_8263,N_5254,N_5003);
nor U8264 (N_8264,N_3074,N_4766);
or U8265 (N_8265,N_5939,N_3112);
and U8266 (N_8266,N_4010,N_3598);
and U8267 (N_8267,N_5481,N_4635);
and U8268 (N_8268,N_5090,N_5483);
and U8269 (N_8269,N_5144,N_3926);
and U8270 (N_8270,N_3352,N_4610);
xor U8271 (N_8271,N_5307,N_4748);
nor U8272 (N_8272,N_3825,N_5971);
nor U8273 (N_8273,N_3596,N_5572);
and U8274 (N_8274,N_5545,N_4670);
or U8275 (N_8275,N_5816,N_3975);
nor U8276 (N_8276,N_3291,N_5057);
or U8277 (N_8277,N_3045,N_5708);
or U8278 (N_8278,N_4945,N_5138);
and U8279 (N_8279,N_3965,N_5770);
nor U8280 (N_8280,N_3712,N_3206);
and U8281 (N_8281,N_4052,N_5506);
or U8282 (N_8282,N_3629,N_3164);
nand U8283 (N_8283,N_5869,N_5733);
nand U8284 (N_8284,N_3792,N_5573);
nor U8285 (N_8285,N_5101,N_5088);
or U8286 (N_8286,N_4977,N_3835);
nor U8287 (N_8287,N_3668,N_4444);
and U8288 (N_8288,N_5971,N_5005);
nand U8289 (N_8289,N_5880,N_5925);
nor U8290 (N_8290,N_5825,N_4603);
and U8291 (N_8291,N_3597,N_4794);
nor U8292 (N_8292,N_5645,N_5926);
or U8293 (N_8293,N_4032,N_5412);
or U8294 (N_8294,N_4893,N_5890);
or U8295 (N_8295,N_3208,N_3787);
and U8296 (N_8296,N_4548,N_4606);
xnor U8297 (N_8297,N_5562,N_3058);
or U8298 (N_8298,N_5461,N_3595);
nand U8299 (N_8299,N_5363,N_4734);
or U8300 (N_8300,N_5219,N_3658);
or U8301 (N_8301,N_5431,N_3528);
nor U8302 (N_8302,N_3364,N_5202);
or U8303 (N_8303,N_5772,N_5431);
nor U8304 (N_8304,N_3704,N_5801);
nand U8305 (N_8305,N_5486,N_3351);
or U8306 (N_8306,N_3111,N_5655);
or U8307 (N_8307,N_4139,N_5833);
or U8308 (N_8308,N_5965,N_4514);
nor U8309 (N_8309,N_4220,N_5584);
and U8310 (N_8310,N_5324,N_5760);
or U8311 (N_8311,N_3994,N_5343);
and U8312 (N_8312,N_3079,N_4013);
xnor U8313 (N_8313,N_4415,N_5339);
xor U8314 (N_8314,N_3095,N_3697);
nor U8315 (N_8315,N_3473,N_3092);
and U8316 (N_8316,N_3088,N_5396);
and U8317 (N_8317,N_4971,N_4434);
nor U8318 (N_8318,N_4361,N_4718);
and U8319 (N_8319,N_5132,N_4370);
and U8320 (N_8320,N_3836,N_4246);
or U8321 (N_8321,N_5637,N_4552);
nor U8322 (N_8322,N_4257,N_4733);
and U8323 (N_8323,N_4075,N_4328);
and U8324 (N_8324,N_3636,N_4137);
nor U8325 (N_8325,N_5002,N_3994);
or U8326 (N_8326,N_5444,N_4123);
and U8327 (N_8327,N_3902,N_3979);
nor U8328 (N_8328,N_5515,N_4629);
nor U8329 (N_8329,N_4918,N_5641);
or U8330 (N_8330,N_4959,N_5479);
or U8331 (N_8331,N_5841,N_4212);
or U8332 (N_8332,N_3065,N_5359);
nor U8333 (N_8333,N_5550,N_3842);
nor U8334 (N_8334,N_5828,N_3935);
nor U8335 (N_8335,N_3917,N_3690);
xnor U8336 (N_8336,N_4746,N_3687);
and U8337 (N_8337,N_5023,N_4819);
nor U8338 (N_8338,N_3524,N_4635);
and U8339 (N_8339,N_3445,N_4682);
or U8340 (N_8340,N_5836,N_5421);
nor U8341 (N_8341,N_3044,N_4279);
nor U8342 (N_8342,N_4946,N_3670);
xor U8343 (N_8343,N_5865,N_4906);
and U8344 (N_8344,N_4526,N_5676);
nand U8345 (N_8345,N_4117,N_3716);
nand U8346 (N_8346,N_5326,N_5383);
or U8347 (N_8347,N_5849,N_5626);
and U8348 (N_8348,N_3192,N_5990);
nor U8349 (N_8349,N_5772,N_4636);
and U8350 (N_8350,N_4290,N_4981);
or U8351 (N_8351,N_4084,N_3112);
and U8352 (N_8352,N_4296,N_4996);
nand U8353 (N_8353,N_4656,N_4960);
xnor U8354 (N_8354,N_3233,N_5387);
nor U8355 (N_8355,N_3135,N_3588);
nor U8356 (N_8356,N_5811,N_3058);
and U8357 (N_8357,N_3481,N_5636);
or U8358 (N_8358,N_5649,N_5758);
nor U8359 (N_8359,N_4297,N_4077);
xnor U8360 (N_8360,N_3062,N_4348);
and U8361 (N_8361,N_5348,N_3631);
nand U8362 (N_8362,N_4124,N_5264);
nand U8363 (N_8363,N_3791,N_4956);
and U8364 (N_8364,N_5181,N_3930);
and U8365 (N_8365,N_5410,N_4522);
nand U8366 (N_8366,N_4395,N_4780);
nor U8367 (N_8367,N_4632,N_4912);
nor U8368 (N_8368,N_4813,N_4864);
or U8369 (N_8369,N_4758,N_3234);
nand U8370 (N_8370,N_5606,N_5130);
nand U8371 (N_8371,N_3855,N_4985);
nor U8372 (N_8372,N_5773,N_5141);
xnor U8373 (N_8373,N_4635,N_4348);
nor U8374 (N_8374,N_3269,N_5526);
nor U8375 (N_8375,N_5758,N_5367);
nor U8376 (N_8376,N_4293,N_5797);
or U8377 (N_8377,N_5692,N_3665);
nor U8378 (N_8378,N_3264,N_3816);
and U8379 (N_8379,N_5300,N_3891);
nand U8380 (N_8380,N_5838,N_3515);
xnor U8381 (N_8381,N_4982,N_5856);
or U8382 (N_8382,N_4264,N_3045);
or U8383 (N_8383,N_4824,N_4437);
nor U8384 (N_8384,N_4538,N_3395);
or U8385 (N_8385,N_5858,N_5614);
or U8386 (N_8386,N_3324,N_4898);
or U8387 (N_8387,N_5657,N_4038);
nand U8388 (N_8388,N_5379,N_4952);
or U8389 (N_8389,N_3625,N_3188);
nor U8390 (N_8390,N_5387,N_3313);
nand U8391 (N_8391,N_4335,N_5882);
and U8392 (N_8392,N_4209,N_5906);
or U8393 (N_8393,N_3298,N_4098);
nand U8394 (N_8394,N_3699,N_5105);
nand U8395 (N_8395,N_3345,N_4849);
or U8396 (N_8396,N_5776,N_3243);
nor U8397 (N_8397,N_3597,N_4791);
and U8398 (N_8398,N_3537,N_4040);
nand U8399 (N_8399,N_4835,N_4614);
nand U8400 (N_8400,N_3619,N_5536);
or U8401 (N_8401,N_4491,N_3567);
nor U8402 (N_8402,N_5070,N_3734);
or U8403 (N_8403,N_5390,N_4302);
or U8404 (N_8404,N_5415,N_5012);
nand U8405 (N_8405,N_3819,N_4099);
xnor U8406 (N_8406,N_3299,N_5880);
xor U8407 (N_8407,N_4010,N_5532);
nor U8408 (N_8408,N_3498,N_5682);
and U8409 (N_8409,N_4963,N_3870);
nor U8410 (N_8410,N_3212,N_3387);
nand U8411 (N_8411,N_5845,N_4879);
nand U8412 (N_8412,N_3338,N_4628);
and U8413 (N_8413,N_4935,N_3876);
and U8414 (N_8414,N_4639,N_5993);
nor U8415 (N_8415,N_5282,N_3893);
xnor U8416 (N_8416,N_3826,N_5362);
and U8417 (N_8417,N_5406,N_3709);
nor U8418 (N_8418,N_3308,N_3850);
nand U8419 (N_8419,N_3951,N_5887);
or U8420 (N_8420,N_4897,N_4868);
nor U8421 (N_8421,N_4693,N_5470);
nor U8422 (N_8422,N_4590,N_5213);
or U8423 (N_8423,N_4204,N_5194);
or U8424 (N_8424,N_5934,N_3498);
nor U8425 (N_8425,N_3559,N_3506);
nand U8426 (N_8426,N_5956,N_3977);
or U8427 (N_8427,N_4673,N_5614);
and U8428 (N_8428,N_5638,N_3497);
xor U8429 (N_8429,N_3515,N_3393);
nand U8430 (N_8430,N_4871,N_4188);
nor U8431 (N_8431,N_5559,N_4962);
or U8432 (N_8432,N_5673,N_5613);
or U8433 (N_8433,N_4141,N_5324);
nor U8434 (N_8434,N_5975,N_4128);
xor U8435 (N_8435,N_5348,N_5356);
and U8436 (N_8436,N_5936,N_3330);
and U8437 (N_8437,N_4294,N_4961);
or U8438 (N_8438,N_3819,N_5280);
nand U8439 (N_8439,N_4156,N_3595);
nand U8440 (N_8440,N_5664,N_5375);
or U8441 (N_8441,N_5776,N_4802);
nor U8442 (N_8442,N_3937,N_5240);
or U8443 (N_8443,N_5256,N_3028);
or U8444 (N_8444,N_4373,N_3145);
nand U8445 (N_8445,N_4690,N_3120);
nand U8446 (N_8446,N_3715,N_4367);
nor U8447 (N_8447,N_3978,N_4007);
and U8448 (N_8448,N_4512,N_3703);
and U8449 (N_8449,N_5081,N_3561);
nand U8450 (N_8450,N_4256,N_4543);
nor U8451 (N_8451,N_5582,N_4891);
nand U8452 (N_8452,N_5968,N_4262);
nand U8453 (N_8453,N_3292,N_3987);
or U8454 (N_8454,N_3284,N_3088);
or U8455 (N_8455,N_4109,N_4001);
nand U8456 (N_8456,N_5489,N_5741);
nor U8457 (N_8457,N_5768,N_3212);
nor U8458 (N_8458,N_5025,N_5544);
and U8459 (N_8459,N_5029,N_5555);
and U8460 (N_8460,N_3720,N_4585);
and U8461 (N_8461,N_3402,N_3965);
nor U8462 (N_8462,N_4288,N_3534);
nand U8463 (N_8463,N_5492,N_5648);
and U8464 (N_8464,N_4861,N_3272);
nor U8465 (N_8465,N_4968,N_5595);
and U8466 (N_8466,N_4455,N_3267);
xnor U8467 (N_8467,N_5187,N_5997);
or U8468 (N_8468,N_5599,N_4901);
or U8469 (N_8469,N_5078,N_4055);
nor U8470 (N_8470,N_3753,N_3424);
xor U8471 (N_8471,N_3533,N_5710);
nand U8472 (N_8472,N_3411,N_5513);
nor U8473 (N_8473,N_4811,N_4179);
and U8474 (N_8474,N_3581,N_5331);
or U8475 (N_8475,N_3950,N_3100);
nand U8476 (N_8476,N_5735,N_5595);
nor U8477 (N_8477,N_5675,N_5672);
and U8478 (N_8478,N_4180,N_4336);
and U8479 (N_8479,N_4314,N_3772);
nor U8480 (N_8480,N_5072,N_4107);
nand U8481 (N_8481,N_3584,N_4491);
or U8482 (N_8482,N_5888,N_5116);
nor U8483 (N_8483,N_3020,N_3322);
nand U8484 (N_8484,N_3363,N_3615);
or U8485 (N_8485,N_4769,N_4028);
nor U8486 (N_8486,N_5439,N_4603);
and U8487 (N_8487,N_3616,N_5272);
or U8488 (N_8488,N_5113,N_5029);
or U8489 (N_8489,N_4722,N_3033);
nor U8490 (N_8490,N_5973,N_4654);
nand U8491 (N_8491,N_5708,N_4962);
and U8492 (N_8492,N_3923,N_4430);
nand U8493 (N_8493,N_4260,N_4843);
and U8494 (N_8494,N_5127,N_3306);
nand U8495 (N_8495,N_4746,N_4242);
nand U8496 (N_8496,N_5572,N_3991);
nand U8497 (N_8497,N_3163,N_4096);
xor U8498 (N_8498,N_5042,N_4569);
and U8499 (N_8499,N_4652,N_4937);
nor U8500 (N_8500,N_4639,N_3812);
and U8501 (N_8501,N_5590,N_3721);
nor U8502 (N_8502,N_4181,N_5555);
and U8503 (N_8503,N_5802,N_5887);
or U8504 (N_8504,N_4113,N_3156);
or U8505 (N_8505,N_5683,N_3646);
and U8506 (N_8506,N_3527,N_5025);
nor U8507 (N_8507,N_3783,N_5521);
or U8508 (N_8508,N_5153,N_4624);
nand U8509 (N_8509,N_4997,N_4103);
and U8510 (N_8510,N_5434,N_3872);
or U8511 (N_8511,N_3818,N_5680);
and U8512 (N_8512,N_4782,N_3246);
xnor U8513 (N_8513,N_3657,N_3804);
or U8514 (N_8514,N_3464,N_5592);
xor U8515 (N_8515,N_4247,N_4963);
nand U8516 (N_8516,N_5750,N_4101);
and U8517 (N_8517,N_5175,N_3812);
nand U8518 (N_8518,N_4725,N_3851);
nand U8519 (N_8519,N_3513,N_3789);
and U8520 (N_8520,N_5700,N_3478);
or U8521 (N_8521,N_5771,N_3240);
nand U8522 (N_8522,N_4542,N_3435);
xnor U8523 (N_8523,N_4996,N_5293);
nand U8524 (N_8524,N_5736,N_4915);
nand U8525 (N_8525,N_4063,N_5212);
nor U8526 (N_8526,N_4760,N_3339);
nand U8527 (N_8527,N_5585,N_5083);
or U8528 (N_8528,N_4088,N_4503);
nor U8529 (N_8529,N_5318,N_4628);
and U8530 (N_8530,N_4816,N_3160);
xor U8531 (N_8531,N_3457,N_4106);
nand U8532 (N_8532,N_4849,N_3500);
nand U8533 (N_8533,N_4868,N_4110);
and U8534 (N_8534,N_3849,N_5707);
nand U8535 (N_8535,N_5628,N_4961);
nand U8536 (N_8536,N_3116,N_3716);
or U8537 (N_8537,N_4090,N_4466);
nand U8538 (N_8538,N_3146,N_5807);
and U8539 (N_8539,N_5093,N_4513);
nor U8540 (N_8540,N_4332,N_5930);
and U8541 (N_8541,N_5076,N_4474);
and U8542 (N_8542,N_3531,N_4788);
nand U8543 (N_8543,N_3614,N_4172);
or U8544 (N_8544,N_5964,N_4786);
or U8545 (N_8545,N_5782,N_5297);
and U8546 (N_8546,N_5809,N_5774);
xor U8547 (N_8547,N_3236,N_4042);
nor U8548 (N_8548,N_5470,N_4429);
or U8549 (N_8549,N_5493,N_3461);
or U8550 (N_8550,N_4850,N_5293);
xnor U8551 (N_8551,N_3747,N_3188);
and U8552 (N_8552,N_3381,N_5328);
nor U8553 (N_8553,N_3795,N_4378);
nand U8554 (N_8554,N_4224,N_5369);
and U8555 (N_8555,N_4272,N_3667);
nand U8556 (N_8556,N_4867,N_3512);
and U8557 (N_8557,N_5523,N_5532);
and U8558 (N_8558,N_4004,N_5852);
xnor U8559 (N_8559,N_4664,N_5193);
or U8560 (N_8560,N_4833,N_5521);
and U8561 (N_8561,N_4961,N_3228);
and U8562 (N_8562,N_3498,N_4161);
or U8563 (N_8563,N_5764,N_5847);
and U8564 (N_8564,N_4439,N_4035);
xnor U8565 (N_8565,N_4247,N_5077);
and U8566 (N_8566,N_5841,N_5215);
and U8567 (N_8567,N_3622,N_4675);
nand U8568 (N_8568,N_3160,N_3320);
nand U8569 (N_8569,N_4855,N_5321);
nor U8570 (N_8570,N_4805,N_3896);
xnor U8571 (N_8571,N_5427,N_5054);
nand U8572 (N_8572,N_5553,N_5863);
xor U8573 (N_8573,N_5699,N_3822);
xnor U8574 (N_8574,N_4361,N_5921);
nand U8575 (N_8575,N_5370,N_3339);
nand U8576 (N_8576,N_3541,N_5319);
or U8577 (N_8577,N_3035,N_5013);
nand U8578 (N_8578,N_5938,N_4484);
or U8579 (N_8579,N_4967,N_4247);
and U8580 (N_8580,N_4215,N_5432);
nand U8581 (N_8581,N_4223,N_3856);
or U8582 (N_8582,N_4649,N_3420);
nand U8583 (N_8583,N_4452,N_3014);
nor U8584 (N_8584,N_5828,N_4178);
and U8585 (N_8585,N_4777,N_4361);
or U8586 (N_8586,N_5601,N_4206);
xnor U8587 (N_8587,N_4955,N_5779);
xor U8588 (N_8588,N_3748,N_5592);
and U8589 (N_8589,N_5832,N_4019);
and U8590 (N_8590,N_5235,N_5199);
nor U8591 (N_8591,N_5169,N_3533);
nor U8592 (N_8592,N_5185,N_4240);
nand U8593 (N_8593,N_4375,N_5164);
nor U8594 (N_8594,N_4402,N_3512);
or U8595 (N_8595,N_4747,N_5654);
nand U8596 (N_8596,N_3635,N_3889);
nor U8597 (N_8597,N_4525,N_4793);
and U8598 (N_8598,N_3985,N_4138);
or U8599 (N_8599,N_3988,N_3058);
nor U8600 (N_8600,N_5707,N_3706);
nand U8601 (N_8601,N_4478,N_5444);
and U8602 (N_8602,N_4034,N_4358);
nand U8603 (N_8603,N_5623,N_4445);
and U8604 (N_8604,N_3460,N_4872);
and U8605 (N_8605,N_3228,N_3908);
or U8606 (N_8606,N_3543,N_3443);
nand U8607 (N_8607,N_5635,N_5696);
nor U8608 (N_8608,N_3762,N_3031);
and U8609 (N_8609,N_3514,N_5487);
nand U8610 (N_8610,N_5863,N_3038);
or U8611 (N_8611,N_3587,N_4610);
nor U8612 (N_8612,N_3011,N_5304);
or U8613 (N_8613,N_3410,N_5744);
nor U8614 (N_8614,N_5634,N_4944);
nand U8615 (N_8615,N_3556,N_4856);
or U8616 (N_8616,N_5701,N_3831);
xor U8617 (N_8617,N_5181,N_3358);
and U8618 (N_8618,N_3238,N_4505);
nor U8619 (N_8619,N_5557,N_4777);
nor U8620 (N_8620,N_4790,N_3963);
nand U8621 (N_8621,N_5477,N_3782);
nor U8622 (N_8622,N_3639,N_5861);
nand U8623 (N_8623,N_3006,N_5861);
nand U8624 (N_8624,N_3320,N_3050);
nand U8625 (N_8625,N_3991,N_3126);
nand U8626 (N_8626,N_5893,N_4613);
nor U8627 (N_8627,N_4458,N_4787);
nand U8628 (N_8628,N_4223,N_5424);
nand U8629 (N_8629,N_3097,N_5361);
and U8630 (N_8630,N_3714,N_4540);
nor U8631 (N_8631,N_5088,N_5646);
nand U8632 (N_8632,N_3694,N_4165);
nor U8633 (N_8633,N_5217,N_4299);
or U8634 (N_8634,N_5713,N_5987);
or U8635 (N_8635,N_5470,N_5524);
nor U8636 (N_8636,N_5331,N_5447);
or U8637 (N_8637,N_4741,N_3202);
nor U8638 (N_8638,N_5274,N_5828);
nand U8639 (N_8639,N_5797,N_5075);
and U8640 (N_8640,N_5639,N_5311);
nand U8641 (N_8641,N_5296,N_5838);
or U8642 (N_8642,N_4476,N_3742);
or U8643 (N_8643,N_3579,N_4551);
or U8644 (N_8644,N_4811,N_5357);
or U8645 (N_8645,N_4598,N_5248);
and U8646 (N_8646,N_5294,N_3809);
nor U8647 (N_8647,N_4065,N_3039);
or U8648 (N_8648,N_3668,N_3489);
nor U8649 (N_8649,N_5162,N_3042);
xor U8650 (N_8650,N_5921,N_3091);
and U8651 (N_8651,N_5493,N_4746);
and U8652 (N_8652,N_3960,N_4413);
xnor U8653 (N_8653,N_4325,N_4415);
and U8654 (N_8654,N_5542,N_5765);
nand U8655 (N_8655,N_5186,N_4571);
nor U8656 (N_8656,N_5216,N_5311);
and U8657 (N_8657,N_5792,N_5385);
xnor U8658 (N_8658,N_4642,N_3850);
nor U8659 (N_8659,N_5962,N_3455);
nand U8660 (N_8660,N_4988,N_3916);
or U8661 (N_8661,N_4867,N_5413);
nor U8662 (N_8662,N_5710,N_4971);
nand U8663 (N_8663,N_3978,N_3017);
nor U8664 (N_8664,N_5842,N_4752);
or U8665 (N_8665,N_3781,N_5601);
or U8666 (N_8666,N_3957,N_3125);
and U8667 (N_8667,N_3174,N_4168);
or U8668 (N_8668,N_5113,N_4356);
or U8669 (N_8669,N_3116,N_5284);
nor U8670 (N_8670,N_5334,N_4932);
or U8671 (N_8671,N_5318,N_4465);
nand U8672 (N_8672,N_4682,N_4572);
or U8673 (N_8673,N_5944,N_4742);
nand U8674 (N_8674,N_3638,N_3540);
nor U8675 (N_8675,N_3044,N_5146);
nor U8676 (N_8676,N_5159,N_4693);
and U8677 (N_8677,N_5174,N_3865);
nand U8678 (N_8678,N_4111,N_3198);
or U8679 (N_8679,N_3468,N_5193);
nand U8680 (N_8680,N_4215,N_5693);
nand U8681 (N_8681,N_4731,N_5369);
nor U8682 (N_8682,N_5997,N_3658);
nor U8683 (N_8683,N_4464,N_3534);
and U8684 (N_8684,N_5117,N_3354);
or U8685 (N_8685,N_3097,N_3383);
nand U8686 (N_8686,N_3439,N_5412);
nor U8687 (N_8687,N_4584,N_3796);
nor U8688 (N_8688,N_3213,N_3920);
and U8689 (N_8689,N_3271,N_3925);
or U8690 (N_8690,N_4046,N_3718);
nand U8691 (N_8691,N_4577,N_5391);
nor U8692 (N_8692,N_3407,N_4198);
nor U8693 (N_8693,N_4173,N_3384);
nor U8694 (N_8694,N_4370,N_4124);
xor U8695 (N_8695,N_4596,N_5738);
or U8696 (N_8696,N_5951,N_3939);
or U8697 (N_8697,N_5699,N_5190);
nor U8698 (N_8698,N_4955,N_3824);
xnor U8699 (N_8699,N_4628,N_4534);
xnor U8700 (N_8700,N_3020,N_5603);
nor U8701 (N_8701,N_3225,N_5391);
nor U8702 (N_8702,N_3170,N_4929);
nor U8703 (N_8703,N_3391,N_5926);
nor U8704 (N_8704,N_4303,N_5369);
and U8705 (N_8705,N_3389,N_3074);
nand U8706 (N_8706,N_4959,N_5997);
and U8707 (N_8707,N_3719,N_4828);
and U8708 (N_8708,N_4136,N_5957);
or U8709 (N_8709,N_4146,N_3158);
xnor U8710 (N_8710,N_3694,N_4531);
nand U8711 (N_8711,N_3105,N_4375);
and U8712 (N_8712,N_5335,N_3168);
or U8713 (N_8713,N_5653,N_4931);
nor U8714 (N_8714,N_3547,N_5129);
nor U8715 (N_8715,N_4698,N_3551);
nor U8716 (N_8716,N_4765,N_5215);
nand U8717 (N_8717,N_3887,N_5553);
nand U8718 (N_8718,N_5884,N_5348);
and U8719 (N_8719,N_5933,N_4535);
and U8720 (N_8720,N_3456,N_4213);
or U8721 (N_8721,N_4744,N_4532);
nand U8722 (N_8722,N_5262,N_5068);
and U8723 (N_8723,N_4162,N_5854);
nor U8724 (N_8724,N_3263,N_3110);
nor U8725 (N_8725,N_4484,N_4663);
or U8726 (N_8726,N_3976,N_4124);
xor U8727 (N_8727,N_4116,N_5712);
nand U8728 (N_8728,N_4123,N_3810);
nor U8729 (N_8729,N_5041,N_5848);
nor U8730 (N_8730,N_5834,N_3468);
and U8731 (N_8731,N_5011,N_4225);
nand U8732 (N_8732,N_4935,N_5893);
nor U8733 (N_8733,N_5821,N_3060);
or U8734 (N_8734,N_5366,N_4169);
xnor U8735 (N_8735,N_3929,N_3049);
or U8736 (N_8736,N_5962,N_3955);
xnor U8737 (N_8737,N_4175,N_5868);
nor U8738 (N_8738,N_3926,N_4153);
and U8739 (N_8739,N_4973,N_3524);
xor U8740 (N_8740,N_3060,N_4998);
nor U8741 (N_8741,N_3398,N_3977);
nand U8742 (N_8742,N_5762,N_3124);
and U8743 (N_8743,N_4589,N_3837);
and U8744 (N_8744,N_5732,N_4055);
nand U8745 (N_8745,N_4827,N_3469);
nor U8746 (N_8746,N_4147,N_5831);
or U8747 (N_8747,N_4292,N_4358);
nand U8748 (N_8748,N_3058,N_4629);
or U8749 (N_8749,N_5082,N_3527);
or U8750 (N_8750,N_4421,N_4052);
nor U8751 (N_8751,N_3591,N_4999);
and U8752 (N_8752,N_5882,N_4780);
or U8753 (N_8753,N_5961,N_3626);
or U8754 (N_8754,N_4256,N_5754);
and U8755 (N_8755,N_5984,N_4828);
or U8756 (N_8756,N_4090,N_4422);
nand U8757 (N_8757,N_5618,N_4695);
nor U8758 (N_8758,N_3622,N_4692);
or U8759 (N_8759,N_3177,N_4569);
or U8760 (N_8760,N_4722,N_3679);
nor U8761 (N_8761,N_4518,N_3114);
and U8762 (N_8762,N_4389,N_3460);
nand U8763 (N_8763,N_4688,N_4480);
or U8764 (N_8764,N_5011,N_4312);
nor U8765 (N_8765,N_3727,N_4966);
or U8766 (N_8766,N_5309,N_4777);
nor U8767 (N_8767,N_5860,N_5558);
and U8768 (N_8768,N_3044,N_5998);
nand U8769 (N_8769,N_3467,N_4183);
nor U8770 (N_8770,N_5819,N_3877);
and U8771 (N_8771,N_3595,N_4805);
nand U8772 (N_8772,N_4412,N_5628);
nand U8773 (N_8773,N_3357,N_3291);
or U8774 (N_8774,N_4937,N_5119);
and U8775 (N_8775,N_5691,N_3099);
and U8776 (N_8776,N_4503,N_5255);
nand U8777 (N_8777,N_4206,N_5769);
nand U8778 (N_8778,N_5757,N_3954);
and U8779 (N_8779,N_5986,N_4209);
nor U8780 (N_8780,N_3284,N_3614);
nor U8781 (N_8781,N_3577,N_5936);
and U8782 (N_8782,N_3272,N_4300);
nor U8783 (N_8783,N_5729,N_4421);
nor U8784 (N_8784,N_3320,N_3243);
nor U8785 (N_8785,N_4437,N_4568);
nand U8786 (N_8786,N_5849,N_3755);
or U8787 (N_8787,N_3241,N_4618);
or U8788 (N_8788,N_3399,N_4959);
or U8789 (N_8789,N_4304,N_5878);
nand U8790 (N_8790,N_5330,N_5374);
or U8791 (N_8791,N_5428,N_3846);
or U8792 (N_8792,N_3758,N_4903);
xor U8793 (N_8793,N_4254,N_4146);
or U8794 (N_8794,N_5324,N_4407);
or U8795 (N_8795,N_5444,N_4027);
and U8796 (N_8796,N_5927,N_4367);
xnor U8797 (N_8797,N_4983,N_5912);
nand U8798 (N_8798,N_3108,N_5737);
nand U8799 (N_8799,N_3574,N_5478);
and U8800 (N_8800,N_4707,N_4263);
nand U8801 (N_8801,N_4695,N_4949);
and U8802 (N_8802,N_5764,N_3409);
and U8803 (N_8803,N_3948,N_5441);
nand U8804 (N_8804,N_5075,N_3144);
nand U8805 (N_8805,N_5463,N_5354);
nand U8806 (N_8806,N_5502,N_4418);
xor U8807 (N_8807,N_4709,N_5087);
nor U8808 (N_8808,N_3125,N_5337);
and U8809 (N_8809,N_4669,N_3995);
and U8810 (N_8810,N_4525,N_3994);
nor U8811 (N_8811,N_4283,N_5292);
xor U8812 (N_8812,N_5057,N_5913);
xor U8813 (N_8813,N_4527,N_4175);
xor U8814 (N_8814,N_3589,N_3647);
nand U8815 (N_8815,N_5784,N_3316);
nor U8816 (N_8816,N_5660,N_5590);
or U8817 (N_8817,N_3684,N_4722);
nand U8818 (N_8818,N_5076,N_3269);
nand U8819 (N_8819,N_5644,N_3694);
or U8820 (N_8820,N_5216,N_3602);
xor U8821 (N_8821,N_4183,N_5878);
xor U8822 (N_8822,N_3953,N_4940);
xor U8823 (N_8823,N_4843,N_3959);
and U8824 (N_8824,N_5943,N_4453);
nor U8825 (N_8825,N_3695,N_5909);
or U8826 (N_8826,N_5048,N_5364);
nor U8827 (N_8827,N_4208,N_3666);
or U8828 (N_8828,N_3048,N_5095);
nor U8829 (N_8829,N_5204,N_3839);
and U8830 (N_8830,N_4081,N_5880);
and U8831 (N_8831,N_5781,N_5488);
xor U8832 (N_8832,N_3416,N_3563);
and U8833 (N_8833,N_5786,N_5463);
xor U8834 (N_8834,N_5248,N_3247);
nor U8835 (N_8835,N_4939,N_5812);
or U8836 (N_8836,N_3138,N_4571);
nor U8837 (N_8837,N_3089,N_5001);
and U8838 (N_8838,N_5274,N_4329);
and U8839 (N_8839,N_4224,N_4101);
and U8840 (N_8840,N_4428,N_3066);
and U8841 (N_8841,N_5291,N_3789);
nor U8842 (N_8842,N_4362,N_5372);
or U8843 (N_8843,N_4134,N_3376);
nand U8844 (N_8844,N_4158,N_5144);
and U8845 (N_8845,N_3034,N_5268);
nor U8846 (N_8846,N_4392,N_5566);
and U8847 (N_8847,N_5750,N_5139);
nand U8848 (N_8848,N_3813,N_3257);
and U8849 (N_8849,N_4005,N_5835);
or U8850 (N_8850,N_5415,N_3406);
or U8851 (N_8851,N_5333,N_3533);
or U8852 (N_8852,N_3705,N_5049);
xor U8853 (N_8853,N_5085,N_4895);
nand U8854 (N_8854,N_5457,N_4764);
nand U8855 (N_8855,N_5985,N_5990);
and U8856 (N_8856,N_4501,N_3934);
nand U8857 (N_8857,N_4430,N_3945);
xnor U8858 (N_8858,N_5569,N_3187);
nand U8859 (N_8859,N_3725,N_4964);
nor U8860 (N_8860,N_4183,N_4212);
and U8861 (N_8861,N_5038,N_3049);
nor U8862 (N_8862,N_3838,N_5656);
and U8863 (N_8863,N_4364,N_3931);
or U8864 (N_8864,N_3278,N_5246);
or U8865 (N_8865,N_4869,N_4662);
nand U8866 (N_8866,N_4680,N_4519);
nand U8867 (N_8867,N_3389,N_5898);
and U8868 (N_8868,N_4332,N_4458);
nor U8869 (N_8869,N_3449,N_4152);
nand U8870 (N_8870,N_5790,N_5960);
and U8871 (N_8871,N_3279,N_3555);
nor U8872 (N_8872,N_3509,N_3936);
nand U8873 (N_8873,N_4824,N_4120);
and U8874 (N_8874,N_4989,N_3541);
xor U8875 (N_8875,N_3537,N_4067);
or U8876 (N_8876,N_5712,N_4591);
nand U8877 (N_8877,N_4533,N_4043);
nor U8878 (N_8878,N_5618,N_4109);
nor U8879 (N_8879,N_3837,N_4212);
nand U8880 (N_8880,N_4942,N_5563);
or U8881 (N_8881,N_3682,N_5762);
nor U8882 (N_8882,N_3842,N_4986);
nand U8883 (N_8883,N_4391,N_3146);
and U8884 (N_8884,N_5766,N_3472);
and U8885 (N_8885,N_5199,N_4766);
nor U8886 (N_8886,N_3793,N_5605);
or U8887 (N_8887,N_3980,N_5220);
xor U8888 (N_8888,N_4636,N_5533);
and U8889 (N_8889,N_5783,N_4078);
nand U8890 (N_8890,N_3182,N_4028);
and U8891 (N_8891,N_4890,N_3110);
or U8892 (N_8892,N_4062,N_4262);
nand U8893 (N_8893,N_5701,N_3650);
or U8894 (N_8894,N_5523,N_3381);
nor U8895 (N_8895,N_4077,N_5670);
nand U8896 (N_8896,N_4529,N_5226);
or U8897 (N_8897,N_4342,N_4428);
and U8898 (N_8898,N_3949,N_5919);
nor U8899 (N_8899,N_3362,N_5429);
nor U8900 (N_8900,N_5024,N_5056);
nand U8901 (N_8901,N_3258,N_5925);
or U8902 (N_8902,N_4627,N_4605);
nor U8903 (N_8903,N_4068,N_3130);
nand U8904 (N_8904,N_4464,N_3377);
and U8905 (N_8905,N_3713,N_4226);
nor U8906 (N_8906,N_4231,N_3863);
xnor U8907 (N_8907,N_5097,N_3652);
and U8908 (N_8908,N_3624,N_5621);
or U8909 (N_8909,N_4225,N_5141);
and U8910 (N_8910,N_3721,N_3818);
and U8911 (N_8911,N_4814,N_5222);
nor U8912 (N_8912,N_5856,N_4003);
nand U8913 (N_8913,N_5169,N_5781);
or U8914 (N_8914,N_5159,N_5265);
nand U8915 (N_8915,N_3113,N_3768);
xor U8916 (N_8916,N_4716,N_3345);
nand U8917 (N_8917,N_3564,N_5235);
nand U8918 (N_8918,N_4106,N_3130);
nor U8919 (N_8919,N_4627,N_5952);
and U8920 (N_8920,N_3996,N_5459);
nor U8921 (N_8921,N_5880,N_5055);
nand U8922 (N_8922,N_4170,N_5434);
and U8923 (N_8923,N_4357,N_4145);
nand U8924 (N_8924,N_4241,N_4332);
nor U8925 (N_8925,N_4006,N_5474);
nand U8926 (N_8926,N_3495,N_4121);
nor U8927 (N_8927,N_3475,N_5223);
and U8928 (N_8928,N_5153,N_4730);
nor U8929 (N_8929,N_3673,N_5997);
and U8930 (N_8930,N_3269,N_3843);
xor U8931 (N_8931,N_5139,N_4093);
nor U8932 (N_8932,N_4101,N_5367);
or U8933 (N_8933,N_4437,N_3952);
or U8934 (N_8934,N_4688,N_4128);
nor U8935 (N_8935,N_4499,N_4298);
or U8936 (N_8936,N_4767,N_5060);
nand U8937 (N_8937,N_3740,N_4588);
or U8938 (N_8938,N_5722,N_4778);
or U8939 (N_8939,N_5472,N_5298);
nor U8940 (N_8940,N_5948,N_5672);
nand U8941 (N_8941,N_4775,N_4891);
nand U8942 (N_8942,N_5572,N_3714);
nand U8943 (N_8943,N_4535,N_4503);
xnor U8944 (N_8944,N_4526,N_4040);
nor U8945 (N_8945,N_4898,N_4406);
and U8946 (N_8946,N_3950,N_3522);
nor U8947 (N_8947,N_3957,N_3622);
nand U8948 (N_8948,N_5791,N_4453);
xor U8949 (N_8949,N_3640,N_4693);
and U8950 (N_8950,N_5541,N_3357);
or U8951 (N_8951,N_3031,N_3292);
and U8952 (N_8952,N_5664,N_4196);
xor U8953 (N_8953,N_5855,N_4194);
or U8954 (N_8954,N_5036,N_5839);
nand U8955 (N_8955,N_3340,N_5156);
nor U8956 (N_8956,N_3711,N_4600);
nor U8957 (N_8957,N_3244,N_3897);
nand U8958 (N_8958,N_3037,N_4903);
and U8959 (N_8959,N_5634,N_5287);
nand U8960 (N_8960,N_3890,N_5460);
nor U8961 (N_8961,N_3147,N_5989);
xor U8962 (N_8962,N_4962,N_3118);
and U8963 (N_8963,N_4933,N_5047);
and U8964 (N_8964,N_5518,N_3497);
nand U8965 (N_8965,N_5517,N_4773);
and U8966 (N_8966,N_3059,N_5102);
or U8967 (N_8967,N_5520,N_5871);
or U8968 (N_8968,N_4899,N_3060);
and U8969 (N_8969,N_4351,N_5170);
nand U8970 (N_8970,N_5638,N_3872);
and U8971 (N_8971,N_3751,N_3910);
nand U8972 (N_8972,N_3059,N_4596);
and U8973 (N_8973,N_3838,N_4107);
nor U8974 (N_8974,N_4516,N_4173);
and U8975 (N_8975,N_5487,N_3610);
and U8976 (N_8976,N_4762,N_4025);
nor U8977 (N_8977,N_4975,N_5157);
nand U8978 (N_8978,N_4863,N_3164);
and U8979 (N_8979,N_3232,N_4821);
and U8980 (N_8980,N_4405,N_3130);
nor U8981 (N_8981,N_4891,N_5756);
nor U8982 (N_8982,N_3184,N_3878);
nor U8983 (N_8983,N_5803,N_5684);
nor U8984 (N_8984,N_3919,N_5033);
or U8985 (N_8985,N_3934,N_5295);
and U8986 (N_8986,N_4733,N_4651);
and U8987 (N_8987,N_4007,N_3147);
or U8988 (N_8988,N_4438,N_3553);
nand U8989 (N_8989,N_3240,N_3153);
xor U8990 (N_8990,N_3317,N_3748);
or U8991 (N_8991,N_4746,N_3607);
or U8992 (N_8992,N_5962,N_5986);
and U8993 (N_8993,N_5408,N_4453);
nand U8994 (N_8994,N_5400,N_3142);
nor U8995 (N_8995,N_4907,N_4015);
and U8996 (N_8996,N_3007,N_4836);
xnor U8997 (N_8997,N_3136,N_5732);
nor U8998 (N_8998,N_3661,N_5858);
and U8999 (N_8999,N_5054,N_3007);
and U9000 (N_9000,N_6802,N_7486);
nand U9001 (N_9001,N_7433,N_7931);
nand U9002 (N_9002,N_6966,N_7908);
nor U9003 (N_9003,N_6085,N_6865);
and U9004 (N_9004,N_8384,N_7422);
nor U9005 (N_9005,N_6965,N_7343);
nor U9006 (N_9006,N_6653,N_7832);
xor U9007 (N_9007,N_8622,N_6396);
or U9008 (N_9008,N_8720,N_6701);
or U9009 (N_9009,N_8824,N_8387);
nand U9010 (N_9010,N_8598,N_7163);
or U9011 (N_9011,N_8898,N_6913);
and U9012 (N_9012,N_7853,N_7362);
nand U9013 (N_9013,N_7238,N_6030);
xnor U9014 (N_9014,N_6582,N_7617);
or U9015 (N_9015,N_7881,N_7518);
or U9016 (N_9016,N_8279,N_7025);
nor U9017 (N_9017,N_7221,N_8793);
nor U9018 (N_9018,N_7594,N_8472);
and U9019 (N_9019,N_7169,N_7217);
nand U9020 (N_9020,N_6687,N_7580);
xor U9021 (N_9021,N_7072,N_7255);
nand U9022 (N_9022,N_7297,N_7212);
nand U9023 (N_9023,N_7314,N_6155);
and U9024 (N_9024,N_8670,N_7969);
xor U9025 (N_9025,N_8674,N_7267);
nor U9026 (N_9026,N_6213,N_6867);
or U9027 (N_9027,N_6325,N_8282);
nand U9028 (N_9028,N_8471,N_7143);
nor U9029 (N_9029,N_6254,N_6864);
nand U9030 (N_9030,N_8284,N_8797);
nand U9031 (N_9031,N_8229,N_6788);
nor U9032 (N_9032,N_7320,N_7423);
or U9033 (N_9033,N_6063,N_7005);
nor U9034 (N_9034,N_7389,N_8699);
xor U9035 (N_9035,N_6719,N_8066);
nand U9036 (N_9036,N_7983,N_7525);
and U9037 (N_9037,N_7904,N_7963);
or U9038 (N_9038,N_8928,N_7354);
nand U9039 (N_9039,N_6319,N_6560);
nand U9040 (N_9040,N_6496,N_7324);
nor U9041 (N_9041,N_8916,N_7364);
and U9042 (N_9042,N_6776,N_6105);
and U9043 (N_9043,N_7570,N_6287);
or U9044 (N_9044,N_7576,N_8374);
and U9045 (N_9045,N_6706,N_6708);
or U9046 (N_9046,N_6064,N_8016);
or U9047 (N_9047,N_8978,N_6925);
and U9048 (N_9048,N_6385,N_7782);
nand U9049 (N_9049,N_7698,N_8303);
nand U9050 (N_9050,N_6519,N_8905);
nand U9051 (N_9051,N_8690,N_8507);
and U9052 (N_9052,N_8707,N_7470);
or U9053 (N_9053,N_6806,N_6799);
or U9054 (N_9054,N_7935,N_6649);
nor U9055 (N_9055,N_6563,N_8032);
and U9056 (N_9056,N_7290,N_7317);
or U9057 (N_9057,N_7269,N_8923);
or U9058 (N_9058,N_8323,N_7916);
nand U9059 (N_9059,N_8798,N_7595);
or U9060 (N_9060,N_7151,N_6623);
nand U9061 (N_9061,N_8342,N_8468);
nor U9062 (N_9062,N_8260,N_7149);
xnor U9063 (N_9063,N_6239,N_8850);
nand U9064 (N_9064,N_7442,N_8606);
xor U9065 (N_9065,N_8435,N_7652);
and U9066 (N_9066,N_6795,N_8930);
nand U9067 (N_9067,N_6414,N_8148);
or U9068 (N_9068,N_8573,N_6309);
xor U9069 (N_9069,N_6497,N_7420);
and U9070 (N_9070,N_6761,N_6245);
xor U9071 (N_9071,N_7167,N_6315);
or U9072 (N_9072,N_7841,N_8790);
or U9073 (N_9073,N_7348,N_7907);
and U9074 (N_9074,N_8831,N_8034);
nor U9075 (N_9075,N_7596,N_6128);
or U9076 (N_9076,N_8580,N_7715);
nor U9077 (N_9077,N_7767,N_6310);
nor U9078 (N_9078,N_8353,N_6347);
nand U9079 (N_9079,N_6292,N_6033);
and U9080 (N_9080,N_7161,N_8003);
or U9081 (N_9081,N_8609,N_7467);
and U9082 (N_9082,N_8454,N_6022);
nand U9083 (N_9083,N_8662,N_8664);
and U9084 (N_9084,N_7224,N_6525);
and U9085 (N_9085,N_8583,N_7798);
or U9086 (N_9086,N_6513,N_8018);
and U9087 (N_9087,N_6791,N_6526);
or U9088 (N_9088,N_7184,N_7358);
and U9089 (N_9089,N_7970,N_7825);
nand U9090 (N_9090,N_7625,N_7446);
or U9091 (N_9091,N_8510,N_7207);
or U9092 (N_9092,N_6205,N_8657);
xnor U9093 (N_9093,N_8906,N_7455);
or U9094 (N_9094,N_8360,N_8095);
nand U9095 (N_9095,N_8306,N_6407);
nor U9096 (N_9096,N_7264,N_8963);
and U9097 (N_9097,N_7557,N_8946);
or U9098 (N_9098,N_7340,N_6627);
nand U9099 (N_9099,N_8421,N_8420);
nor U9100 (N_9100,N_7171,N_8896);
and U9101 (N_9101,N_8001,N_8723);
nor U9102 (N_9102,N_7061,N_6814);
nand U9103 (N_9103,N_8070,N_7794);
or U9104 (N_9104,N_8271,N_6759);
nor U9105 (N_9105,N_7023,N_8777);
and U9106 (N_9106,N_8935,N_7731);
xor U9107 (N_9107,N_7559,N_8378);
xnor U9108 (N_9108,N_6992,N_8731);
and U9109 (N_9109,N_6394,N_7887);
and U9110 (N_9110,N_7547,N_7399);
nand U9111 (N_9111,N_7771,N_7564);
nand U9112 (N_9112,N_8236,N_7646);
nand U9113 (N_9113,N_8774,N_8621);
nand U9114 (N_9114,N_6252,N_8447);
or U9115 (N_9115,N_8947,N_6147);
or U9116 (N_9116,N_7382,N_6444);
or U9117 (N_9117,N_7342,N_8814);
and U9118 (N_9118,N_6723,N_6735);
and U9119 (N_9119,N_7818,N_8127);
or U9120 (N_9120,N_8410,N_8301);
nor U9121 (N_9121,N_6968,N_7544);
and U9122 (N_9122,N_6584,N_7001);
or U9123 (N_9123,N_7016,N_7651);
and U9124 (N_9124,N_6432,N_8629);
nor U9125 (N_9125,N_6928,N_6982);
nand U9126 (N_9126,N_8542,N_8596);
and U9127 (N_9127,N_8822,N_8547);
or U9128 (N_9128,N_8105,N_7249);
nor U9129 (N_9129,N_8595,N_7676);
nand U9130 (N_9130,N_8779,N_8239);
nor U9131 (N_9131,N_6754,N_7742);
and U9132 (N_9132,N_8524,N_7502);
and U9133 (N_9133,N_7851,N_6301);
and U9134 (N_9134,N_7835,N_8626);
nor U9135 (N_9135,N_7081,N_7300);
and U9136 (N_9136,N_6467,N_8735);
nand U9137 (N_9137,N_8948,N_7632);
nor U9138 (N_9138,N_7968,N_6770);
or U9139 (N_9139,N_8285,N_7836);
xnor U9140 (N_9140,N_6400,N_6683);
and U9141 (N_9141,N_8204,N_6411);
and U9142 (N_9142,N_7303,N_7511);
nor U9143 (N_9143,N_6704,N_7624);
nand U9144 (N_9144,N_8685,N_8737);
nor U9145 (N_9145,N_7589,N_8048);
nand U9146 (N_9146,N_6995,N_6975);
and U9147 (N_9147,N_7550,N_8660);
nand U9148 (N_9148,N_7438,N_7694);
xor U9149 (N_9149,N_7110,N_6220);
nand U9150 (N_9150,N_8815,N_7093);
nand U9151 (N_9151,N_7233,N_8484);
xnor U9152 (N_9152,N_8241,N_7519);
or U9153 (N_9153,N_6569,N_6980);
nor U9154 (N_9154,N_6748,N_8897);
and U9155 (N_9155,N_6591,N_6124);
or U9156 (N_9156,N_6293,N_6388);
nand U9157 (N_9157,N_8405,N_8183);
nand U9158 (N_9158,N_6994,N_7042);
and U9159 (N_9159,N_7689,N_6577);
nand U9160 (N_9160,N_7417,N_7966);
nand U9161 (N_9161,N_6068,N_8477);
or U9162 (N_9162,N_8367,N_7156);
xor U9163 (N_9163,N_8880,N_8638);
or U9164 (N_9164,N_7280,N_7458);
or U9165 (N_9165,N_7638,N_8876);
nor U9166 (N_9166,N_8732,N_7574);
or U9167 (N_9167,N_7487,N_8529);
or U9168 (N_9168,N_6734,N_6820);
or U9169 (N_9169,N_6237,N_7478);
and U9170 (N_9170,N_6323,N_7049);
nor U9171 (N_9171,N_6466,N_7037);
and U9172 (N_9172,N_8298,N_8783);
nand U9173 (N_9173,N_8373,N_8841);
or U9174 (N_9174,N_6760,N_7736);
nor U9175 (N_9175,N_8718,N_7288);
and U9176 (N_9176,N_7507,N_8316);
nor U9177 (N_9177,N_6556,N_7601);
nand U9178 (N_9178,N_8403,N_8740);
nand U9179 (N_9179,N_8076,N_6018);
nand U9180 (N_9180,N_8543,N_6811);
and U9181 (N_9181,N_6740,N_6280);
or U9182 (N_9182,N_7755,N_6099);
and U9183 (N_9183,N_7130,N_8646);
nand U9184 (N_9184,N_6756,N_7327);
nor U9185 (N_9185,N_7359,N_6118);
xor U9186 (N_9186,N_6449,N_6565);
nand U9187 (N_9187,N_6721,N_6051);
xor U9188 (N_9188,N_8220,N_8463);
nand U9189 (N_9189,N_8188,N_6831);
xor U9190 (N_9190,N_8173,N_6720);
xnor U9191 (N_9191,N_6424,N_8912);
or U9192 (N_9192,N_7797,N_6522);
or U9193 (N_9193,N_6349,N_6674);
nor U9194 (N_9194,N_8641,N_6987);
and U9195 (N_9195,N_8321,N_8357);
and U9196 (N_9196,N_8406,N_6717);
and U9197 (N_9197,N_7418,N_8124);
or U9198 (N_9198,N_8918,N_8624);
or U9199 (N_9199,N_6613,N_7241);
and U9200 (N_9200,N_7088,N_6114);
nand U9201 (N_9201,N_7246,N_8602);
and U9202 (N_9202,N_7956,N_8952);
nand U9203 (N_9203,N_6132,N_8487);
nor U9204 (N_9204,N_7747,N_6600);
nor U9205 (N_9205,N_8027,N_8516);
and U9206 (N_9206,N_7972,N_8592);
nor U9207 (N_9207,N_7326,N_8838);
and U9208 (N_9208,N_8211,N_7822);
and U9209 (N_9209,N_6086,N_8578);
nor U9210 (N_9210,N_8676,N_7137);
nand U9211 (N_9211,N_6176,N_6264);
xor U9212 (N_9212,N_6011,N_8564);
or U9213 (N_9213,N_7136,N_7411);
nand U9214 (N_9214,N_7035,N_7769);
xnor U9215 (N_9215,N_6379,N_7410);
and U9216 (N_9216,N_6681,N_6692);
xnor U9217 (N_9217,N_8224,N_8361);
nand U9218 (N_9218,N_6651,N_7645);
and U9219 (N_9219,N_6212,N_6045);
and U9220 (N_9220,N_7391,N_8747);
and U9221 (N_9221,N_7593,N_8870);
nand U9222 (N_9222,N_7295,N_6830);
nor U9223 (N_9223,N_8225,N_7273);
or U9224 (N_9224,N_6026,N_6738);
and U9225 (N_9225,N_6890,N_7152);
or U9226 (N_9226,N_8151,N_8396);
and U9227 (N_9227,N_8545,N_7817);
and U9228 (N_9228,N_6171,N_6421);
xnor U9229 (N_9229,N_7707,N_7394);
nor U9230 (N_9230,N_6423,N_8663);
and U9231 (N_9231,N_6163,N_6278);
nor U9232 (N_9232,N_7809,N_6036);
or U9233 (N_9233,N_7346,N_7670);
nor U9234 (N_9234,N_7351,N_7223);
nor U9235 (N_9235,N_8345,N_7933);
nor U9236 (N_9236,N_6062,N_6373);
nand U9237 (N_9237,N_7393,N_6991);
nand U9238 (N_9238,N_6558,N_6112);
and U9239 (N_9239,N_6305,N_8419);
or U9240 (N_9240,N_8376,N_7902);
or U9241 (N_9241,N_7682,N_8479);
nor U9242 (N_9242,N_8203,N_8072);
nor U9243 (N_9243,N_8985,N_8615);
and U9244 (N_9244,N_8766,N_8244);
and U9245 (N_9245,N_6710,N_6328);
nor U9246 (N_9246,N_8552,N_6906);
xor U9247 (N_9247,N_7950,N_8769);
xnor U9248 (N_9248,N_7690,N_8757);
and U9249 (N_9249,N_6142,N_6611);
xnor U9250 (N_9250,N_7792,N_8894);
nor U9251 (N_9251,N_6202,N_7901);
xor U9252 (N_9252,N_8891,N_6604);
nor U9253 (N_9253,N_6946,N_6680);
nand U9254 (N_9254,N_7484,N_7180);
nand U9255 (N_9255,N_6023,N_7315);
nand U9256 (N_9256,N_7777,N_8069);
nand U9257 (N_9257,N_7134,N_7710);
and U9258 (N_9258,N_7889,N_6034);
and U9259 (N_9259,N_8845,N_7336);
xnor U9260 (N_9260,N_7367,N_8518);
nand U9261 (N_9261,N_6457,N_6886);
nor U9262 (N_9262,N_7140,N_6718);
or U9263 (N_9263,N_8304,N_7400);
or U9264 (N_9264,N_7607,N_6047);
or U9265 (N_9265,N_7059,N_7425);
and U9266 (N_9266,N_6833,N_6574);
or U9267 (N_9267,N_7662,N_6543);
and U9268 (N_9268,N_7090,N_6390);
nand U9269 (N_9269,N_8253,N_6076);
nand U9270 (N_9270,N_8625,N_7196);
xor U9271 (N_9271,N_8568,N_7802);
nand U9272 (N_9272,N_7746,N_7614);
or U9273 (N_9273,N_8953,N_8842);
nand U9274 (N_9274,N_8090,N_7347);
nor U9275 (N_9275,N_6371,N_6025);
nor U9276 (N_9276,N_6950,N_6822);
or U9277 (N_9277,N_8277,N_6620);
or U9278 (N_9278,N_6183,N_7844);
nand U9279 (N_9279,N_6339,N_6797);
or U9280 (N_9280,N_8145,N_7789);
and U9281 (N_9281,N_8425,N_8789);
or U9282 (N_9282,N_7743,N_8776);
and U9283 (N_9283,N_6387,N_6167);
xnor U9284 (N_9284,N_8551,N_6366);
xor U9285 (N_9285,N_6426,N_6534);
nand U9286 (N_9286,N_8979,N_6066);
nor U9287 (N_9287,N_7366,N_6312);
nand U9288 (N_9288,N_6358,N_6849);
or U9289 (N_9289,N_7162,N_7095);
nor U9290 (N_9290,N_7256,N_7157);
nor U9291 (N_9291,N_7248,N_8539);
or U9292 (N_9292,N_6931,N_6515);
and U9293 (N_9293,N_8871,N_6903);
and U9294 (N_9294,N_7104,N_7724);
and U9295 (N_9295,N_7258,N_6599);
nor U9296 (N_9296,N_7843,N_6859);
or U9297 (N_9297,N_7080,N_7545);
or U9298 (N_9298,N_6789,N_7172);
nor U9299 (N_9299,N_7655,N_7178);
and U9300 (N_9300,N_7074,N_7700);
or U9301 (N_9301,N_8859,N_8143);
and U9302 (N_9302,N_6286,N_7975);
nor U9303 (N_9303,N_7930,N_8724);
and U9304 (N_9304,N_8497,N_7980);
nor U9305 (N_9305,N_6967,N_8589);
and U9306 (N_9306,N_6468,N_6862);
nand U9307 (N_9307,N_8557,N_7855);
nand U9308 (N_9308,N_6383,N_8337);
nand U9309 (N_9309,N_6088,N_6750);
nand U9310 (N_9310,N_8112,N_6330);
xnor U9311 (N_9311,N_8567,N_6947);
nand U9312 (N_9312,N_7503,N_8658);
xor U9313 (N_9313,N_7261,N_8250);
and U9314 (N_9314,N_6669,N_7067);
or U9315 (N_9315,N_8168,N_6164);
and U9316 (N_9316,N_6976,N_7361);
or U9317 (N_9317,N_8288,N_6943);
and U9318 (N_9318,N_8759,N_7457);
and U9319 (N_9319,N_7365,N_8125);
nor U9320 (N_9320,N_7195,N_8009);
and U9321 (N_9321,N_7128,N_8908);
nand U9322 (N_9322,N_7277,N_7415);
or U9323 (N_9323,N_6785,N_7926);
nand U9324 (N_9324,N_8319,N_8778);
nor U9325 (N_9325,N_6356,N_7115);
nor U9326 (N_9326,N_7122,N_8054);
or U9327 (N_9327,N_6075,N_7582);
and U9328 (N_9328,N_7721,N_6634);
nor U9329 (N_9329,N_7893,N_8825);
nand U9330 (N_9330,N_7513,N_6927);
or U9331 (N_9331,N_8509,N_7461);
or U9332 (N_9332,N_7360,N_7938);
or U9333 (N_9333,N_8972,N_7448);
nor U9334 (N_9334,N_8764,N_7813);
nor U9335 (N_9335,N_7220,N_8043);
and U9336 (N_9336,N_6741,N_8678);
xor U9337 (N_9337,N_6537,N_8362);
and U9338 (N_9338,N_8170,N_6544);
and U9339 (N_9339,N_6374,N_6170);
or U9340 (N_9340,N_8645,N_8816);
and U9341 (N_9341,N_6012,N_6110);
or U9342 (N_9342,N_6889,N_7649);
nand U9343 (N_9343,N_8563,N_6794);
and U9344 (N_9344,N_8493,N_7170);
or U9345 (N_9345,N_8398,N_8619);
nor U9346 (N_9346,N_8934,N_6261);
nand U9347 (N_9347,N_7884,N_8469);
nor U9348 (N_9348,N_6529,N_8352);
and U9349 (N_9349,N_8084,N_8293);
nand U9350 (N_9350,N_7575,N_8459);
and U9351 (N_9351,N_7540,N_7636);
nor U9352 (N_9352,N_7044,N_6089);
or U9353 (N_9353,N_8553,N_7793);
and U9354 (N_9354,N_8957,N_8937);
or U9355 (N_9355,N_7066,N_8581);
and U9356 (N_9356,N_8268,N_8617);
and U9357 (N_9357,N_6617,N_6377);
nor U9358 (N_9358,N_7087,N_7039);
nand U9359 (N_9359,N_8780,N_7370);
or U9360 (N_9360,N_6199,N_7718);
nand U9361 (N_9361,N_6531,N_6905);
nand U9362 (N_9362,N_8801,N_6974);
or U9363 (N_9363,N_8940,N_8498);
nor U9364 (N_9364,N_6667,N_7378);
xor U9365 (N_9365,N_6007,N_8171);
or U9366 (N_9366,N_7020,N_7432);
and U9367 (N_9367,N_7201,N_6250);
nand U9368 (N_9368,N_7621,N_6067);
nand U9369 (N_9369,N_7641,N_6838);
nand U9370 (N_9370,N_8541,N_6002);
nor U9371 (N_9371,N_6549,N_7929);
or U9372 (N_9372,N_6178,N_7754);
and U9373 (N_9373,N_7937,N_7030);
xor U9374 (N_9374,N_7356,N_7735);
and U9375 (N_9375,N_8071,N_8700);
or U9376 (N_9376,N_8721,N_6194);
and U9377 (N_9377,N_7664,N_6032);
nand U9378 (N_9378,N_7560,N_6041);
nor U9379 (N_9379,N_8827,N_6953);
nor U9380 (N_9380,N_7027,N_8432);
and U9381 (N_9381,N_7739,N_6490);
xnor U9382 (N_9382,N_6695,N_7403);
and U9383 (N_9383,N_8393,N_8719);
or U9384 (N_9384,N_6314,N_7244);
nor U9385 (N_9385,N_8976,N_7236);
xor U9386 (N_9386,N_6470,N_7758);
nor U9387 (N_9387,N_6597,N_7052);
xnor U9388 (N_9388,N_6930,N_8917);
nand U9389 (N_9389,N_7083,N_7940);
nor U9390 (N_9390,N_6020,N_7435);
or U9391 (N_9391,N_7600,N_7471);
xnor U9392 (N_9392,N_6601,N_8892);
or U9393 (N_9393,N_7133,N_7860);
nor U9394 (N_9394,N_8730,N_8667);
or U9395 (N_9395,N_8470,N_7460);
xor U9396 (N_9396,N_6185,N_8865);
or U9397 (N_9397,N_8587,N_6907);
and U9398 (N_9398,N_7232,N_7711);
or U9399 (N_9399,N_6697,N_7637);
nor U9400 (N_9400,N_6632,N_8813);
xnor U9401 (N_9401,N_8131,N_8695);
nor U9402 (N_9402,N_7831,N_7033);
or U9403 (N_9403,N_7284,N_8669);
nand U9404 (N_9404,N_7078,N_8988);
or U9405 (N_9405,N_7079,N_6688);
nand U9406 (N_9406,N_8149,N_7615);
xnor U9407 (N_9407,N_8457,N_7786);
nand U9408 (N_9408,N_8430,N_8409);
or U9409 (N_9409,N_6472,N_8096);
nor U9410 (N_9410,N_8294,N_6957);
xor U9411 (N_9411,N_6887,N_6231);
nand U9412 (N_9412,N_8633,N_7572);
and U9413 (N_9413,N_6283,N_8270);
nor U9414 (N_9414,N_8610,N_6778);
xnor U9415 (N_9415,N_8291,N_7534);
or U9416 (N_9416,N_7823,N_8575);
nand U9417 (N_9417,N_7866,N_7973);
or U9418 (N_9418,N_7390,N_8944);
or U9419 (N_9419,N_8181,N_8412);
nand U9420 (N_9420,N_6360,N_7807);
and U9421 (N_9421,N_6494,N_8480);
and U9422 (N_9422,N_7310,N_7006);
nand U9423 (N_9423,N_6686,N_8295);
nor U9424 (N_9424,N_7165,N_7064);
or U9425 (N_9425,N_8200,N_6877);
nor U9426 (N_9426,N_8175,N_6324);
nand U9427 (N_9427,N_6475,N_8179);
nor U9428 (N_9428,N_8063,N_8237);
nor U9429 (N_9429,N_8058,N_7612);
or U9430 (N_9430,N_6450,N_6751);
nor U9431 (N_9431,N_8915,N_6342);
or U9432 (N_9432,N_8649,N_8812);
or U9433 (N_9433,N_7135,N_8061);
or U9434 (N_9434,N_8828,N_6443);
nor U9435 (N_9435,N_7556,N_7727);
and U9436 (N_9436,N_6873,N_8426);
nand U9437 (N_9437,N_8147,N_7146);
nand U9438 (N_9438,N_6476,N_6046);
xnor U9439 (N_9439,N_7979,N_8289);
or U9440 (N_9440,N_7190,N_8786);
nor U9441 (N_9441,N_7848,N_6798);
or U9442 (N_9442,N_8981,N_8004);
and U9443 (N_9443,N_8531,N_8476);
nor U9444 (N_9444,N_8372,N_7581);
nor U9445 (N_9445,N_6460,N_8166);
nand U9446 (N_9446,N_7597,N_8679);
and U9447 (N_9447,N_8002,N_8921);
or U9448 (N_9448,N_6345,N_8257);
or U9449 (N_9449,N_7820,N_7753);
nor U9450 (N_9450,N_8659,N_7286);
xor U9451 (N_9451,N_7337,N_6001);
and U9452 (N_9452,N_6902,N_6891);
nand U9453 (N_9453,N_6266,N_6869);
and U9454 (N_9454,N_6469,N_8184);
nor U9455 (N_9455,N_7604,N_8423);
nor U9456 (N_9456,N_7586,N_8579);
nand U9457 (N_9457,N_6429,N_6442);
and U9458 (N_9458,N_8222,N_8240);
and U9459 (N_9459,N_6072,N_7392);
and U9460 (N_9460,N_6731,N_8330);
and U9461 (N_9461,N_8017,N_6391);
nor U9462 (N_9462,N_8332,N_8242);
and U9463 (N_9463,N_8485,N_8849);
nand U9464 (N_9464,N_8840,N_8888);
or U9465 (N_9465,N_7021,N_6733);
or U9466 (N_9466,N_6643,N_8178);
and U9467 (N_9467,N_6103,N_6079);
nor U9468 (N_9468,N_8109,N_7858);
xor U9469 (N_9469,N_6899,N_8087);
nand U9470 (N_9470,N_8931,N_6677);
nand U9471 (N_9471,N_7543,N_8358);
nand U9472 (N_9472,N_7386,N_6042);
nand U9473 (N_9473,N_8433,N_6304);
xor U9474 (N_9474,N_6431,N_6782);
or U9475 (N_9475,N_7237,N_6017);
nand U9476 (N_9476,N_8982,N_7949);
nor U9477 (N_9477,N_7756,N_7322);
and U9478 (N_9478,N_6844,N_6875);
nand U9479 (N_9479,N_6850,N_7265);
nand U9480 (N_9480,N_6592,N_8414);
nand U9481 (N_9481,N_8689,N_7330);
and U9482 (N_9482,N_7723,N_6065);
nand U9483 (N_9483,N_8548,N_7506);
and U9484 (N_9484,N_7148,N_8893);
nand U9485 (N_9485,N_6160,N_8956);
nand U9486 (N_9486,N_6979,N_7076);
nor U9487 (N_9487,N_6948,N_8212);
or U9488 (N_9488,N_8041,N_8258);
or U9489 (N_9489,N_8141,N_7780);
xnor U9490 (N_9490,N_6826,N_8038);
or U9491 (N_9491,N_7827,N_8861);
nand U9492 (N_9492,N_8512,N_6297);
or U9493 (N_9493,N_7591,N_8377);
and U9494 (N_9494,N_6193,N_7101);
nor U9495 (N_9495,N_7229,N_8455);
nor U9496 (N_9496,N_7107,N_8245);
xnor U9497 (N_9497,N_7894,N_7176);
nand U9498 (N_9498,N_7494,N_8855);
nor U9499 (N_9499,N_6334,N_8161);
xor U9500 (N_9500,N_6668,N_6535);
nand U9501 (N_9501,N_6236,N_7650);
nand U9502 (N_9502,N_6208,N_8913);
or U9503 (N_9503,N_7186,N_7943);
nor U9504 (N_9504,N_7869,N_7092);
nand U9505 (N_9505,N_6179,N_8642);
xnor U9506 (N_9506,N_6863,N_8902);
and U9507 (N_9507,N_6074,N_8513);
nand U9508 (N_9508,N_6546,N_7882);
and U9509 (N_9509,N_7606,N_6146);
and U9510 (N_9510,N_6727,N_8417);
nand U9511 (N_9511,N_7730,N_6917);
or U9512 (N_9512,N_8320,N_6939);
nor U9513 (N_9513,N_8634,N_8152);
and U9514 (N_9514,N_7729,N_8427);
and U9515 (N_9515,N_6175,N_6126);
xnor U9516 (N_9516,N_6221,N_6841);
and U9517 (N_9517,N_8651,N_7629);
nand U9518 (N_9518,N_6428,N_7630);
and U9519 (N_9519,N_8746,N_6972);
nand U9520 (N_9520,N_6793,N_7177);
xor U9521 (N_9521,N_6548,N_7912);
nand U9522 (N_9522,N_8193,N_7608);
xnor U9523 (N_9523,N_8770,N_7877);
nor U9524 (N_9524,N_8121,N_7406);
xnor U9525 (N_9525,N_6227,N_8682);
or U9526 (N_9526,N_8554,N_8750);
nand U9527 (N_9527,N_7381,N_7395);
nand U9528 (N_9528,N_6612,N_7720);
xor U9529 (N_9529,N_8481,N_6463);
and U9530 (N_9530,N_8969,N_7944);
nor U9531 (N_9531,N_8961,N_6284);
or U9532 (N_9532,N_8068,N_6921);
nor U9533 (N_9533,N_6629,N_8273);
nor U9534 (N_9534,N_7291,N_6696);
nand U9535 (N_9535,N_6511,N_6458);
and U9536 (N_9536,N_7274,N_7047);
nand U9537 (N_9537,N_7824,N_6823);
nand U9538 (N_9538,N_8502,N_6282);
nand U9539 (N_9539,N_8226,N_6077);
nand U9540 (N_9540,N_6944,N_6187);
nand U9541 (N_9541,N_6610,N_8137);
or U9542 (N_9542,N_6916,N_6614);
or U9543 (N_9543,N_6169,N_7138);
nand U9544 (N_9544,N_7837,N_6641);
xnor U9545 (N_9545,N_6153,N_6263);
nor U9546 (N_9546,N_8052,N_6219);
nand U9547 (N_9547,N_8252,N_8460);
or U9548 (N_9548,N_8451,N_8379);
nor U9549 (N_9549,N_8208,N_6699);
nor U9550 (N_9550,N_8115,N_6352);
and U9551 (N_9551,N_8555,N_6434);
xnor U9552 (N_9552,N_7849,N_6350);
or U9553 (N_9553,N_8118,N_6378);
or U9554 (N_9554,N_7722,N_8311);
or U9555 (N_9555,N_6897,N_7728);
or U9556 (N_9556,N_8909,N_7204);
or U9557 (N_9557,N_6985,N_7760);
nor U9558 (N_9558,N_7150,N_8190);
and U9559 (N_9559,N_7429,N_8269);
nor U9560 (N_9560,N_6354,N_6329);
nand U9561 (N_9561,N_8164,N_7099);
nor U9562 (N_9562,N_6988,N_6098);
nor U9563 (N_9563,N_6180,N_8853);
nand U9564 (N_9564,N_7982,N_7821);
and U9565 (N_9565,N_7385,N_6145);
or U9566 (N_9566,N_8062,N_7541);
nand U9567 (N_9567,N_7012,N_6125);
and U9568 (N_9568,N_6027,N_8694);
nor U9569 (N_9569,N_7466,N_8799);
and U9570 (N_9570,N_6082,N_6532);
xnor U9571 (N_9571,N_8160,N_6436);
or U9572 (N_9572,N_7790,N_6553);
nand U9573 (N_9573,N_8097,N_7463);
nor U9574 (N_9574,N_8274,N_8787);
nand U9575 (N_9575,N_6945,N_6542);
nor U9576 (N_9576,N_8180,N_8247);
and U9577 (N_9577,N_8576,N_6403);
nor U9578 (N_9578,N_6644,N_8534);
nand U9579 (N_9579,N_7474,N_8429);
and U9580 (N_9580,N_6861,N_6919);
xor U9581 (N_9581,N_6878,N_6858);
and U9582 (N_9582,N_8078,N_8517);
nor U9583 (N_9583,N_8749,N_8019);
nor U9584 (N_9584,N_7257,N_7993);
xor U9585 (N_9585,N_8942,N_6996);
xnor U9586 (N_9586,N_6109,N_7911);
nand U9587 (N_9587,N_6210,N_7766);
xor U9588 (N_9588,N_8458,N_6359);
and U9589 (N_9589,N_8895,N_6936);
xnor U9590 (N_9590,N_7865,N_7663);
nor U9591 (N_9591,N_7068,N_6807);
nor U9592 (N_9592,N_8021,N_8005);
nor U9593 (N_9593,N_8612,N_6365);
nor U9594 (N_9594,N_8120,N_8566);
and U9595 (N_9595,N_7942,N_8727);
xnor U9596 (N_9596,N_6726,N_7245);
xnor U9597 (N_9597,N_6016,N_7815);
and U9598 (N_9598,N_6824,N_6915);
or U9599 (N_9599,N_6372,N_7187);
or U9600 (N_9600,N_8846,N_7407);
and U9601 (N_9601,N_8951,N_7842);
and U9602 (N_9602,N_7311,N_8308);
nor U9603 (N_9603,N_8117,N_8436);
and U9604 (N_9604,N_6698,N_8452);
xnor U9605 (N_9605,N_6435,N_6914);
or U9606 (N_9606,N_7209,N_7856);
nand U9607 (N_9607,N_6473,N_7464);
or U9608 (N_9608,N_6455,N_6240);
or U9609 (N_9609,N_6321,N_8743);
nor U9610 (N_9610,N_8739,N_7009);
nor U9611 (N_9611,N_7024,N_6078);
xor U9612 (N_9612,N_6904,N_7833);
and U9613 (N_9613,N_8307,N_8920);
and U9614 (N_9614,N_6217,N_8675);
nor U9615 (N_9615,N_7770,N_8556);
nor U9616 (N_9616,N_6840,N_7974);
and U9617 (N_9617,N_7350,N_8418);
or U9618 (N_9618,N_7666,N_6447);
nor U9619 (N_9619,N_8359,N_6425);
nand U9620 (N_9620,N_8520,N_6048);
and U9621 (N_9621,N_6302,N_7971);
or U9622 (N_9622,N_7199,N_7071);
nand U9623 (N_9623,N_8191,N_8527);
and U9624 (N_9624,N_6724,N_7775);
xnor U9625 (N_9625,N_6736,N_6765);
nand U9626 (N_9626,N_8462,N_6722);
and U9627 (N_9627,N_7109,N_8984);
nor U9628 (N_9628,N_8108,N_8856);
or U9629 (N_9629,N_7687,N_6575);
nand U9630 (N_9630,N_8010,N_8977);
nor U9631 (N_9631,N_7799,N_8826);
xnor U9632 (N_9632,N_6631,N_6464);
and U9633 (N_9633,N_6061,N_6123);
nand U9634 (N_9634,N_7281,N_7527);
and U9635 (N_9635,N_8407,N_7211);
nor U9636 (N_9636,N_8064,N_8572);
and U9637 (N_9637,N_7283,N_8221);
xnor U9638 (N_9638,N_6102,N_7452);
nand U9639 (N_9639,N_7231,N_6881);
nor U9640 (N_9640,N_7900,N_7892);
nand U9641 (N_9641,N_8050,N_7819);
nor U9642 (N_9642,N_8704,N_6941);
nor U9643 (N_9643,N_7537,N_7397);
nor U9644 (N_9644,N_8099,N_7379);
and U9645 (N_9645,N_8530,N_7387);
nor U9646 (N_9646,N_7773,N_6427);
nand U9647 (N_9647,N_8139,N_6196);
and U9648 (N_9648,N_8440,N_7644);
or U9649 (N_9649,N_7434,N_8093);
xor U9650 (N_9650,N_6729,N_8867);
and U9651 (N_9651,N_8495,N_7616);
nand U9652 (N_9652,N_6491,N_6267);
xnor U9653 (N_9653,N_6006,N_6624);
nor U9654 (N_9654,N_7371,N_6080);
nand U9655 (N_9655,N_7155,N_7840);
nand U9656 (N_9656,N_8681,N_6895);
or U9657 (N_9657,N_8300,N_7857);
xnor U9658 (N_9658,N_8051,N_6550);
and U9659 (N_9659,N_6561,N_8637);
or U9660 (N_9660,N_8706,N_8037);
and U9661 (N_9661,N_6413,N_8665);
and U9662 (N_9662,N_7905,N_8796);
nor U9663 (N_9663,N_7485,N_6910);
nor U9664 (N_9664,N_8317,N_8983);
and U9665 (N_9665,N_7501,N_8782);
or U9666 (N_9666,N_7194,N_8833);
nand U9667 (N_9667,N_8805,N_8914);
nor U9668 (N_9668,N_7160,N_8199);
and U9669 (N_9669,N_7703,N_8057);
nand U9670 (N_9670,N_8561,N_8594);
nor U9671 (N_9671,N_8369,N_7218);
nor U9672 (N_9672,N_8000,N_8333);
or U9673 (N_9673,N_8290,N_8710);
and U9674 (N_9674,N_7750,N_8701);
or U9675 (N_9675,N_6320,N_8601);
nand U9676 (N_9676,N_8980,N_8365);
and U9677 (N_9677,N_7127,N_8185);
or U9678 (N_9678,N_7213,N_8600);
xnor U9679 (N_9679,N_8315,N_7398);
and U9680 (N_9680,N_6602,N_8830);
and U9681 (N_9681,N_6783,N_6509);
or U9682 (N_9682,N_7189,N_7271);
and U9683 (N_9683,N_8733,N_8623);
nand U9684 (N_9684,N_8847,N_8754);
or U9685 (N_9685,N_6682,N_7917);
or U9686 (N_9686,N_8355,N_7363);
nand U9687 (N_9687,N_6485,N_8925);
and U9688 (N_9688,N_8883,N_6564);
nor U9689 (N_9689,N_6595,N_7959);
or U9690 (N_9690,N_8413,N_6892);
nor U9691 (N_9691,N_6281,N_6876);
nor U9692 (N_9692,N_8741,N_6230);
nand U9693 (N_9693,N_7870,N_7688);
nor U9694 (N_9694,N_6004,N_7490);
nand U9695 (N_9695,N_7699,N_6851);
nor U9696 (N_9696,N_8878,N_6445);
nor U9697 (N_9697,N_6728,N_6559);
nor U9698 (N_9698,N_6998,N_7656);
and U9699 (N_9699,N_7712,N_8113);
nand U9700 (N_9700,N_7964,N_6804);
and U9701 (N_9701,N_7495,N_8158);
or U9702 (N_9702,N_8959,N_7878);
or U9703 (N_9703,N_7779,N_8119);
or U9704 (N_9704,N_6583,N_8142);
or U9705 (N_9705,N_8040,N_8562);
nand U9706 (N_9706,N_6316,N_8404);
xnor U9707 (N_9707,N_7528,N_7622);
nand U9708 (N_9708,N_6091,N_8910);
nor U9709 (N_9709,N_7555,N_8620);
nand U9710 (N_9710,N_8255,N_8089);
or U9711 (N_9711,N_6096,N_8287);
nor U9712 (N_9712,N_8614,N_6603);
nand U9713 (N_9713,N_7481,N_7631);
or U9714 (N_9714,N_7997,N_6937);
and U9715 (N_9715,N_6214,N_6693);
and U9716 (N_9716,N_8522,N_7325);
and U9717 (N_9717,N_7384,N_6201);
or U9718 (N_9718,N_7899,N_6572);
and U9719 (N_9719,N_7492,N_8872);
xor U9720 (N_9720,N_8067,N_7714);
and U9721 (N_9721,N_8088,N_8195);
or U9722 (N_9722,N_6755,N_7522);
xnor U9723 (N_9723,N_7424,N_8761);
nor U9724 (N_9724,N_7480,N_8297);
nor U9725 (N_9725,N_6121,N_6679);
xnor U9726 (N_9726,N_6037,N_7628);
and U9727 (N_9727,N_6964,N_6417);
or U9728 (N_9728,N_8533,N_8194);
or U9729 (N_9729,N_8785,N_6083);
nand U9730 (N_9730,N_6576,N_8202);
or U9731 (N_9731,N_8186,N_6622);
and U9732 (N_9732,N_6161,N_6134);
xor U9733 (N_9733,N_6204,N_6866);
and U9734 (N_9734,N_7546,N_6580);
nor U9735 (N_9735,N_6662,N_8494);
and U9736 (N_9736,N_6389,N_7952);
or U9737 (N_9737,N_6771,N_6547);
xnor U9738 (N_9738,N_7154,N_6958);
and U9739 (N_9739,N_6557,N_7341);
and U9740 (N_9740,N_7913,N_6271);
nor U9741 (N_9741,N_8176,N_8726);
nand U9742 (N_9742,N_8126,N_8677);
and U9743 (N_9743,N_8538,N_8744);
nor U9744 (N_9744,N_8008,N_8080);
nor U9745 (N_9745,N_6308,N_6144);
nor U9746 (N_9746,N_8499,N_7234);
xor U9747 (N_9747,N_6203,N_6493);
nor U9748 (N_9748,N_6709,N_8968);
or U9749 (N_9749,N_8283,N_7440);
and U9750 (N_9750,N_7801,N_8742);
nor U9751 (N_9751,N_8715,N_6961);
or U9752 (N_9752,N_7296,N_8990);
and U9753 (N_9753,N_7734,N_7909);
nand U9754 (N_9754,N_7814,N_6246);
and U9755 (N_9755,N_6581,N_7986);
or U9756 (N_9756,N_8683,N_6639);
and U9757 (N_9757,N_6168,N_6159);
or U9758 (N_9758,N_7620,N_6081);
nand U9759 (N_9759,N_8577,N_7675);
nand U9760 (N_9760,N_7272,N_7007);
xnor U9761 (N_9761,N_7924,N_8390);
nor U9762 (N_9762,N_8234,N_7654);
or U9763 (N_9763,N_8392,N_6555);
nand U9764 (N_9764,N_6660,N_8570);
or U9765 (N_9765,N_8475,N_8994);
and U9766 (N_9766,N_7948,N_7579);
or U9767 (N_9767,N_6784,N_8795);
nor U9768 (N_9768,N_6059,N_7462);
nand U9769 (N_9769,N_6270,N_7228);
and U9770 (N_9770,N_7427,N_8364);
nor U9771 (N_9771,N_7058,N_6812);
xor U9772 (N_9772,N_8438,N_8177);
nand U9773 (N_9773,N_7483,N_6970);
or U9774 (N_9774,N_8877,N_8559);
or U9775 (N_9775,N_8022,N_6151);
or U9776 (N_9776,N_7174,N_7102);
nand U9777 (N_9777,N_8899,N_8198);
nand U9778 (N_9778,N_6439,N_7847);
or U9779 (N_9779,N_8924,N_8966);
or U9780 (N_9780,N_6712,N_8725);
or U9781 (N_9781,N_7705,N_7015);
or U9782 (N_9782,N_6843,N_6981);
nand U9783 (N_9783,N_6399,N_6725);
or U9784 (N_9784,N_7552,N_8549);
and U9785 (N_9785,N_6874,N_8085);
xor U9786 (N_9786,N_6313,N_7992);
nand U9787 (N_9787,N_8336,N_8227);
nor U9788 (N_9788,N_6607,N_6362);
nor U9789 (N_9789,N_8327,N_6277);
and U9790 (N_9790,N_7329,N_8079);
or U9791 (N_9791,N_7701,N_8525);
nand U9792 (N_9792,N_8231,N_8416);
and U9793 (N_9793,N_8347,N_7744);
or U9794 (N_9794,N_7254,N_6625);
xor U9795 (N_9795,N_7977,N_8781);
nor U9796 (N_9796,N_8705,N_8394);
nor U9797 (N_9797,N_6969,N_7738);
or U9798 (N_9798,N_7331,N_7627);
or U9799 (N_9799,N_8446,N_6392);
nand U9800 (N_9800,N_6395,N_6508);
nor U9801 (N_9801,N_8356,N_6815);
and U9802 (N_9802,N_6571,N_8380);
nor U9803 (N_9803,N_6474,N_8162);
nor U9804 (N_9804,N_6932,N_7584);
nor U9805 (N_9805,N_6415,N_6780);
and U9806 (N_9806,N_8207,N_6689);
nand U9807 (N_9807,N_7748,N_6593);
nand U9808 (N_9808,N_7680,N_8696);
and U9809 (N_9809,N_6370,N_6567);
xor U9810 (N_9810,N_6842,N_8514);
nand U9811 (N_9811,N_6586,N_8886);
nand U9812 (N_9812,N_8490,N_7953);
or U9813 (N_9813,N_7623,N_7334);
nor U9814 (N_9814,N_7145,N_8015);
nor U9815 (N_9815,N_8835,N_6757);
xnor U9816 (N_9816,N_6279,N_8262);
nand U9817 (N_9817,N_7475,N_8150);
nor U9818 (N_9818,N_7316,N_6441);
xor U9819 (N_9819,N_6656,N_6223);
and U9820 (N_9820,N_7441,N_7193);
nor U9821 (N_9821,N_7695,N_6684);
nor U9822 (N_9822,N_6024,N_8272);
or U9823 (N_9823,N_8031,N_6615);
or U9824 (N_9824,N_8466,N_6053);
nor U9825 (N_9825,N_8305,N_7019);
nor U9826 (N_9826,N_6952,N_8400);
nand U9827 (N_9827,N_8467,N_7182);
nor U9828 (N_9828,N_6386,N_7094);
or U9829 (N_9829,N_6005,N_8954);
nand U9830 (N_9830,N_7175,N_8680);
nor U9831 (N_9831,N_6685,N_7414);
and U9832 (N_9832,N_6655,N_8035);
nand U9833 (N_9833,N_7962,N_6381);
nand U9834 (N_9834,N_6596,N_7055);
nor U9835 (N_9835,N_7285,N_8745);
nor U9836 (N_9836,N_6405,N_8643);
nor U9837 (N_9837,N_8028,N_8110);
nand U9838 (N_9838,N_8292,N_8932);
nor U9839 (N_9839,N_6299,N_7214);
nor U9840 (N_9840,N_6148,N_8042);
nor U9841 (N_9841,N_7549,N_7610);
and U9842 (N_9842,N_8039,N_7338);
or U9843 (N_9843,N_8686,N_8784);
or U9844 (N_9844,N_6049,N_8450);
xor U9845 (N_9845,N_6821,N_8157);
and U9846 (N_9846,N_8264,N_8431);
nand U9847 (N_9847,N_8960,N_8174);
nand U9848 (N_9848,N_8722,N_8210);
or U9849 (N_9849,N_7004,N_8092);
nor U9850 (N_9850,N_7197,N_6195);
and U9851 (N_9851,N_7751,N_6691);
or U9852 (N_9852,N_8864,N_6298);
nand U9853 (N_9853,N_6380,N_6471);
nand U9854 (N_9854,N_6181,N_7561);
and U9855 (N_9855,N_8111,N_6664);
nor U9856 (N_9856,N_7266,N_7469);
and U9857 (N_9857,N_6855,N_6768);
or U9858 (N_9858,N_7567,N_8644);
or U9859 (N_9859,N_6773,N_7761);
nand U9860 (N_9860,N_8671,N_7499);
nand U9861 (N_9861,N_7768,N_8474);
nor U9862 (N_9862,N_6251,N_6554);
nand U9863 (N_9863,N_6249,N_6816);
nor U9864 (N_9864,N_8900,N_7599);
nand U9865 (N_9865,N_8523,N_6503);
or U9866 (N_9866,N_6355,N_7278);
and U9867 (N_9867,N_8007,N_7871);
or U9868 (N_9868,N_7696,N_8368);
and U9869 (N_9869,N_8496,N_8688);
xor U9870 (N_9870,N_8197,N_6954);
nand U9871 (N_9871,N_8586,N_7191);
nand U9872 (N_9872,N_8329,N_7111);
or U9873 (N_9873,N_6705,N_7376);
xnor U9874 (N_9874,N_6742,N_6498);
or U9875 (N_9875,N_6141,N_8875);
nand U9876 (N_9876,N_6882,N_6233);
nor U9877 (N_9877,N_7585,N_6353);
nor U9878 (N_9878,N_6507,N_8478);
nand U9879 (N_9879,N_6129,N_7210);
nand U9880 (N_9880,N_7203,N_6552);
and U9881 (N_9881,N_8630,N_6256);
nor U9882 (N_9882,N_6690,N_8030);
nand U9883 (N_9883,N_8189,N_7609);
nor U9884 (N_9884,N_8033,N_8386);
xor U9885 (N_9885,N_8339,N_7830);
and U9886 (N_9886,N_6416,N_8571);
xor U9887 (N_9887,N_7598,N_8103);
nor U9888 (N_9888,N_8044,N_8442);
nand U9889 (N_9889,N_7845,N_6215);
and U9890 (N_9890,N_7995,N_6092);
and U9891 (N_9891,N_7275,N_7114);
nand U9892 (N_9892,N_8648,N_8604);
or U9893 (N_9893,N_6448,N_6343);
or U9894 (N_9894,N_7526,N_7554);
and U9895 (N_9895,N_6010,N_8970);
and U9896 (N_9896,N_6138,N_8736);
or U9897 (N_9897,N_7569,N_6764);
or U9898 (N_9898,N_7250,N_7252);
nand U9899 (N_9899,N_7957,N_7867);
or U9900 (N_9900,N_8453,N_8312);
or U9901 (N_9901,N_7915,N_7185);
nand U9902 (N_9902,N_7812,N_6197);
and U9903 (N_9903,N_7205,N_8863);
xnor U9904 (N_9904,N_8217,N_8763);
nand U9905 (N_9905,N_8232,N_6094);
and U9906 (N_9906,N_7251,N_7895);
or U9907 (N_9907,N_7661,N_6714);
nor U9908 (N_9908,N_8219,N_8807);
and U9909 (N_9909,N_7578,N_7558);
xnor U9910 (N_9910,N_8388,N_7709);
or U9911 (N_9911,N_7961,N_8266);
xnor U9912 (N_9912,N_7022,N_7542);
xnor U9913 (N_9913,N_6654,N_6920);
nor U9914 (N_9914,N_6817,N_8869);
and U9915 (N_9915,N_7684,N_8140);
nor U9916 (N_9916,N_6346,N_7618);
and U9917 (N_9917,N_7808,N_6884);
nand U9918 (N_9918,N_8267,N_6670);
nor U9919 (N_9919,N_7377,N_7922);
nand U9920 (N_9920,N_7032,N_7313);
or U9921 (N_9921,N_6929,N_6166);
nand U9922 (N_9922,N_7774,N_8811);
nand U9923 (N_9923,N_8881,N_8036);
and U9924 (N_9924,N_8936,N_6095);
and U9925 (N_9925,N_6290,N_8691);
or U9926 (N_9926,N_7987,N_8773);
nor U9927 (N_9927,N_8020,N_6702);
or U9928 (N_9928,N_8804,N_6140);
xnor U9929 (N_9929,N_6940,N_8102);
or U9930 (N_9930,N_7301,N_8762);
or U9931 (N_9931,N_6570,N_6541);
and U9932 (N_9932,N_7733,N_8249);
and U9933 (N_9933,N_6839,N_6753);
or U9934 (N_9934,N_6322,N_8668);
nor U9935 (N_9935,N_7955,N_8574);
or U9936 (N_9936,N_7679,N_6938);
nor U9937 (N_9937,N_7057,N_8758);
nand U9938 (N_9938,N_8535,N_7879);
or U9939 (N_9939,N_8756,N_7671);
and U9940 (N_9940,N_8585,N_6226);
nor U9941 (N_9941,N_8890,N_6232);
or U9942 (N_9942,N_8823,N_7029);
nor U9943 (N_9943,N_8216,N_6671);
nand U9944 (N_9944,N_7141,N_6158);
and U9945 (N_9945,N_8887,N_6478);
nor U9946 (N_9946,N_6506,N_8182);
and U9947 (N_9947,N_7740,N_8248);
and U9948 (N_9948,N_7491,N_7985);
nor U9949 (N_9949,N_7873,N_6206);
and U9950 (N_9950,N_8169,N_8343);
and U9951 (N_9951,N_6262,N_6422);
or U9952 (N_9952,N_7538,N_6484);
nand U9953 (N_9953,N_6218,N_6327);
and U9954 (N_9954,N_7051,N_8546);
nand U9955 (N_9955,N_7605,N_7054);
and U9956 (N_9956,N_8803,N_8666);
nand U9957 (N_9957,N_8537,N_6637);
nor U9958 (N_9958,N_6870,N_7489);
nand U9959 (N_9959,N_8965,N_6527);
and U9960 (N_9960,N_6070,N_8366);
xnor U9961 (N_9961,N_6052,N_6828);
xor U9962 (N_9962,N_6853,N_7803);
or U9963 (N_9963,N_6918,N_6888);
nand U9964 (N_9964,N_7667,N_7886);
and U9965 (N_9965,N_8540,N_8215);
or U9966 (N_9966,N_7551,N_6260);
nand U9967 (N_9967,N_8006,N_7200);
or U9968 (N_9968,N_7863,N_7323);
nor U9969 (N_9969,N_6135,N_7373);
or U9970 (N_9970,N_6137,N_6749);
nor U9971 (N_9971,N_8882,N_7279);
xor U9972 (N_9972,N_7374,N_6156);
or U9973 (N_9973,N_6014,N_7512);
xor U9974 (N_9974,N_7800,N_8331);
nand U9975 (N_9975,N_7778,N_6832);
and U9976 (N_9976,N_7116,N_8672);
nor U9977 (N_9977,N_6291,N_6306);
or U9978 (N_9978,N_6040,N_8024);
and U9979 (N_9979,N_6335,N_7673);
or U9980 (N_9980,N_6951,N_6273);
or U9981 (N_9981,N_7838,N_6451);
nand U9982 (N_9982,N_6787,N_7401);
nand U9983 (N_9983,N_7897,N_7439);
xnor U9984 (N_9984,N_6716,N_6338);
or U9985 (N_9985,N_8059,N_8999);
nor U9986 (N_9986,N_6152,N_8053);
and U9987 (N_9987,N_6259,N_8172);
and U9988 (N_9988,N_8134,N_7105);
nand U9989 (N_9989,N_7643,N_6578);
nand U9990 (N_9990,N_8428,N_8263);
nor U9991 (N_9991,N_6489,N_6589);
nor U9992 (N_9992,N_6288,N_6139);
nand U9993 (N_9993,N_8238,N_6357);
nand U9994 (N_9994,N_6452,N_7681);
nor U9995 (N_9995,N_6375,N_7885);
and U9996 (N_9996,N_8395,N_6019);
or U9997 (N_9997,N_7568,N_7890);
nand U9998 (N_9998,N_7372,N_8919);
xnor U9999 (N_9999,N_6154,N_8280);
or U10000 (N_10000,N_8049,N_8639);
nand U10001 (N_10001,N_6117,N_7500);
nor U10002 (N_10002,N_7259,N_7914);
and U10003 (N_10003,N_6487,N_7921);
nor U10004 (N_10004,N_7240,N_7934);
or U10005 (N_10005,N_8950,N_7045);
and U10006 (N_10006,N_8708,N_6410);
xnor U10007 (N_10007,N_6453,N_7683);
or U10008 (N_10008,N_8964,N_6073);
xnor U10009 (N_10009,N_6935,N_7089);
nand U10010 (N_10010,N_6157,N_7772);
or U10011 (N_10011,N_6307,N_8286);
or U10012 (N_10012,N_8322,N_8504);
and U10013 (N_10013,N_8101,N_6188);
xnor U10014 (N_10014,N_8631,N_7862);
and U10015 (N_10015,N_7126,N_7419);
nor U10016 (N_10016,N_6200,N_8709);
or U10017 (N_10017,N_7118,N_7413);
and U10018 (N_10018,N_7243,N_6488);
nand U10019 (N_10019,N_7717,N_6031);
and U10020 (N_10020,N_8370,N_6598);
nor U10021 (N_10021,N_6566,N_7014);
nor U10022 (N_10022,N_7611,N_7179);
xnor U10023 (N_10023,N_7369,N_7043);
or U10024 (N_10024,N_8652,N_6894);
nor U10025 (N_10025,N_8163,N_7781);
nor U10026 (N_10026,N_7562,N_6326);
nor U10027 (N_10027,N_7668,N_8593);
nand U10028 (N_10028,N_6856,N_6562);
nor U10029 (N_10029,N_6949,N_7757);
nor U10030 (N_10030,N_6590,N_8655);
or U10031 (N_10031,N_6645,N_7678);
or U10032 (N_10032,N_8128,N_8302);
or U10033 (N_10033,N_8521,N_7686);
nor U10034 (N_10034,N_8949,N_7276);
or U10035 (N_10035,N_8692,N_6296);
and U10036 (N_10036,N_8136,N_7289);
and U10037 (N_10037,N_7344,N_6116);
xnor U10038 (N_10038,N_6732,N_6311);
nand U10039 (N_10039,N_8505,N_6647);
nand U10040 (N_10040,N_7496,N_6454);
nor U10041 (N_10041,N_7806,N_6922);
nand U10042 (N_10042,N_8156,N_6056);
and U10043 (N_10043,N_8437,N_7031);
or U10044 (N_10044,N_8590,N_7060);
and U10045 (N_10045,N_6650,N_7725);
or U10046 (N_10046,N_7805,N_7208);
nand U10047 (N_10047,N_8943,N_8256);
xnor U10048 (N_10048,N_7106,N_8318);
nor U10049 (N_10049,N_7328,N_6340);
nand U10050 (N_10050,N_6628,N_8091);
and U10051 (N_10051,N_6364,N_8821);
xor U10052 (N_10052,N_8341,N_7428);
or U10053 (N_10053,N_8138,N_6758);
or U10054 (N_10054,N_6265,N_7763);
nand U10055 (N_10055,N_8086,N_7298);
xnor U10056 (N_10056,N_6763,N_7708);
and U10057 (N_10057,N_7070,N_7826);
nand U10058 (N_10058,N_8338,N_6235);
and U10059 (N_10059,N_7498,N_6908);
or U10060 (N_10060,N_8792,N_8526);
xor U10061 (N_10061,N_6480,N_8354);
or U10062 (N_10062,N_8081,N_7339);
xnor U10063 (N_10063,N_7635,N_8926);
or U10064 (N_10064,N_8927,N_8196);
nand U10065 (N_10065,N_6955,N_6766);
nor U10066 (N_10066,N_7976,N_8397);
and U10067 (N_10067,N_6419,N_8313);
or U10068 (N_10068,N_6810,N_6275);
and U10069 (N_10069,N_8082,N_8884);
nand U10070 (N_10070,N_7529,N_6912);
and U10071 (N_10071,N_6521,N_7693);
nor U10072 (N_10072,N_6983,N_7131);
nor U10073 (N_10073,N_7634,N_6510);
xor U10074 (N_10074,N_6652,N_6638);
or U10075 (N_10075,N_8734,N_7253);
xnor U10076 (N_10076,N_6333,N_6341);
xor U10077 (N_10077,N_8025,N_7077);
xor U10078 (N_10078,N_8808,N_8011);
nand U10079 (N_10079,N_6568,N_7810);
xor U10080 (N_10080,N_7046,N_7144);
and U10081 (N_10081,N_8201,N_8768);
nor U10082 (N_10082,N_7784,N_8760);
and U10083 (N_10083,N_6971,N_7053);
nor U10084 (N_10084,N_8987,N_6715);
xnor U10085 (N_10085,N_7026,N_8399);
and U10086 (N_10086,N_6635,N_7765);
nor U10087 (N_10087,N_8837,N_7173);
or U10088 (N_10088,N_6993,N_8060);
and U10089 (N_10089,N_8265,N_6829);
nand U10090 (N_10090,N_6605,N_6295);
xor U10091 (N_10091,N_6924,N_6803);
or U10092 (N_10092,N_7764,N_6111);
xnor U10093 (N_10093,N_7038,N_6382);
or U10094 (N_10094,N_7565,N_7521);
nand U10095 (N_10095,N_8444,N_6348);
and U10096 (N_10096,N_8698,N_8996);
or U10097 (N_10097,N_6837,N_7430);
and U10098 (N_10098,N_6367,N_8159);
nand U10099 (N_10099,N_8973,N_6540);
nand U10100 (N_10100,N_8489,N_6739);
or U10101 (N_10101,N_7590,N_6393);
or U10102 (N_10102,N_7989,N_7697);
nand U10103 (N_10103,N_6009,N_6274);
xnor U10104 (N_10104,N_8628,N_8056);
xnor U10105 (N_10105,N_6536,N_6579);
or U10106 (N_10106,N_7691,N_7669);
nand U10107 (N_10107,N_8314,N_8627);
or U10108 (N_10108,N_8794,N_7910);
nor U10109 (N_10109,N_6055,N_8165);
nand U10110 (N_10110,N_8975,N_6805);
nor U10111 (N_10111,N_8144,N_6642);
nand U10112 (N_10112,N_8326,N_8635);
nor U10113 (N_10113,N_8246,N_8055);
xor U10114 (N_10114,N_7539,N_8456);
nor U10115 (N_10115,N_6289,N_8986);
or U10116 (N_10116,N_7380,N_6767);
and U10117 (N_10117,N_8501,N_6893);
or U10118 (N_10118,N_7299,N_6462);
nand U10119 (N_10119,N_8065,N_6100);
and U10120 (N_10120,N_6186,N_7444);
and U10121 (N_10121,N_7459,N_8486);
nor U10122 (N_10122,N_8375,N_7181);
nor U10123 (N_10123,N_7451,N_8788);
nand U10124 (N_10124,N_8461,N_6420);
nand U10125 (N_10125,N_8483,N_7056);
or U10126 (N_10126,N_6926,N_6224);
and U10127 (N_10127,N_7292,N_6499);
nand U10128 (N_10128,N_8866,N_7941);
nor U10129 (N_10129,N_7065,N_6101);
nand U10130 (N_10130,N_6446,N_7121);
and U10131 (N_10131,N_8904,N_6984);
and U10132 (N_10132,N_7520,N_6825);
xnor U10133 (N_10133,N_6737,N_8346);
and U10134 (N_10134,N_8862,N_6182);
nor U10135 (N_10135,N_8611,N_7129);
nand U10136 (N_10136,N_8938,N_7119);
and U10137 (N_10137,N_7776,N_7293);
nand U10138 (N_10138,N_7159,N_7517);
nand U10139 (N_10139,N_8584,N_8939);
nand U10140 (N_10140,N_8133,N_6344);
nor U10141 (N_10141,N_7139,N_8962);
nor U10142 (N_10142,N_7225,N_6276);
nand U10143 (N_10143,N_8647,N_7454);
nand U10144 (N_10144,N_8223,N_6746);
nand U10145 (N_10145,N_6621,N_7333);
and U10146 (N_10146,N_6545,N_7898);
and U10147 (N_10147,N_7548,N_7168);
and U10148 (N_10148,N_8752,N_7349);
or U10149 (N_10149,N_7888,N_8714);
nand U10150 (N_10150,N_8836,N_6868);
nor U10151 (N_10151,N_7312,N_6514);
xnor U10152 (N_10152,N_7965,N_6997);
nand U10153 (N_10153,N_8422,N_8684);
and U10154 (N_10154,N_7880,N_7996);
nor U10155 (N_10155,N_6618,N_6150);
nor U10156 (N_10156,N_7945,N_6694);
nand U10157 (N_10157,N_7713,N_6130);
xnor U10158 (N_10158,N_8729,N_8135);
nor U10159 (N_10159,N_6136,N_7473);
nand U10160 (N_10160,N_6192,N_6351);
nor U10161 (N_10161,N_8488,N_6880);
and U10162 (N_10162,N_8636,N_6836);
nand U10163 (N_10163,N_7988,N_8114);
nor U10164 (N_10164,N_6483,N_7332);
nand U10165 (N_10165,N_6923,N_7626);
or U10166 (N_10166,N_7447,N_6207);
and U10167 (N_10167,N_8441,N_6481);
nand U10168 (N_10168,N_8077,N_8775);
nor U10169 (N_10169,N_8945,N_6000);
and U10170 (N_10170,N_7091,N_7219);
nand U10171 (N_10171,N_8998,N_6573);
nor U10172 (N_10172,N_8492,N_7449);
nand U10173 (N_10173,N_7426,N_8309);
and U10174 (N_10174,N_8100,N_8132);
nor U10175 (N_10175,N_6847,N_6819);
xor U10176 (N_10176,N_7226,N_7692);
nor U10177 (N_10177,N_8349,N_6551);
and U10178 (N_10178,N_6190,N_6626);
nand U10179 (N_10179,N_6963,N_7306);
or U10180 (N_10180,N_6769,N_7749);
nor U10181 (N_10181,N_7002,N_7465);
and U10182 (N_10182,N_6285,N_8503);
nand U10183 (N_10183,N_6258,N_6003);
or U10184 (N_10184,N_6173,N_7932);
and U10185 (N_10185,N_6854,N_6456);
xnor U10186 (N_10186,N_8351,N_6228);
or U10187 (N_10187,N_6516,N_7307);
nand U10188 (N_10188,N_7939,N_7978);
nand U10189 (N_10189,N_7260,N_7308);
nand U10190 (N_10190,N_7946,N_6021);
and U10191 (N_10191,N_8519,N_8771);
or U10192 (N_10192,N_6071,N_6255);
or U10193 (N_10193,N_8955,N_8755);
nor U10194 (N_10194,N_8772,N_6404);
nor U10195 (N_10195,N_6113,N_8560);
or U10196 (N_10196,N_6104,N_8192);
xor U10197 (N_10197,N_7183,N_6465);
nor U10198 (N_10198,N_6711,N_7011);
nor U10199 (N_10199,N_6106,N_8254);
nand U10200 (N_10200,N_8713,N_8703);
or U10201 (N_10201,N_7536,N_7850);
nor U10202 (N_10202,N_8653,N_6588);
or U10203 (N_10203,N_6933,N_8500);
nor U10204 (N_10204,N_7345,N_8296);
and U10205 (N_10205,N_6752,N_6376);
and U10206 (N_10206,N_7482,N_7998);
nand U10207 (N_10207,N_8154,N_6962);
or U10208 (N_10208,N_8605,N_7302);
and U10209 (N_10209,N_6242,N_8233);
and U10210 (N_10210,N_7158,N_8971);
nor U10211 (N_10211,N_6777,N_6504);
nor U10212 (N_10212,N_8728,N_7294);
or U10213 (N_10213,N_6492,N_7097);
or U10214 (N_10214,N_6225,N_6896);
and U10215 (N_10215,N_7990,N_8153);
nor U10216 (N_10216,N_7192,N_8654);
or U10217 (N_10217,N_8408,N_6500);
and U10218 (N_10218,N_7639,N_7874);
nand U10219 (N_10219,N_6029,N_8599);
and U10220 (N_10220,N_6459,N_6745);
and U10221 (N_10221,N_7741,N_6744);
and U10222 (N_10222,N_7925,N_8094);
nand U10223 (N_10223,N_6331,N_7967);
nand U10224 (N_10224,N_8995,N_6672);
or U10225 (N_10225,N_7657,N_7408);
xnor U10226 (N_10226,N_7906,N_7431);
nand U10227 (N_10227,N_7745,N_8424);
or U10228 (N_10228,N_7216,N_6336);
xnor U10229 (N_10229,N_8911,N_7416);
nand U10230 (N_10230,N_6058,N_8335);
nor U10231 (N_10231,N_6977,N_8230);
or U10232 (N_10232,N_6879,N_8613);
nor U10233 (N_10233,N_6043,N_6959);
nand U10234 (N_10234,N_8411,N_8122);
nor U10235 (N_10235,N_6028,N_7783);
nor U10236 (N_10236,N_8276,N_7685);
or U10237 (N_10237,N_8389,N_7437);
and U10238 (N_10238,N_6845,N_6700);
and U10239 (N_10239,N_8992,N_8098);
or U10240 (N_10240,N_6433,N_6317);
nor U10241 (N_10241,N_6039,N_7305);
nor U10242 (N_10242,N_6108,N_7123);
and U10243 (N_10243,N_6479,N_7592);
xnor U10244 (N_10244,N_6678,N_6008);
and U10245 (N_10245,N_8922,N_7839);
nor U10246 (N_10246,N_7619,N_6477);
nand U10247 (N_10247,N_6406,N_8550);
nor U10248 (N_10248,N_7861,N_6846);
or U10249 (N_10249,N_6060,N_6633);
nor U10250 (N_10250,N_8717,N_8278);
xor U10251 (N_10251,N_7375,N_7704);
nand U10252 (N_10252,N_8511,N_8187);
nor U10253 (N_10253,N_7450,N_7010);
nor U10254 (N_10254,N_8800,N_7706);
nand U10255 (N_10255,N_6883,N_6222);
or U10256 (N_10256,N_8104,N_6885);
nand U10257 (N_10257,N_7493,N_7535);
and U10258 (N_10258,N_8820,N_6122);
nand U10259 (N_10259,N_6942,N_8464);
nand U10260 (N_10260,N_6661,N_7896);
or U10261 (N_10261,N_6871,N_8046);
nor U10262 (N_10262,N_6216,N_7075);
nand U10263 (N_10263,N_8829,N_8844);
nand U10264 (N_10264,N_8385,N_8434);
and U10265 (N_10265,N_8281,N_7859);
nor U10266 (N_10266,N_6189,N_6666);
nor U10267 (N_10267,N_6809,N_8348);
and U10268 (N_10268,N_8228,N_7927);
and U10269 (N_10269,N_7553,N_6398);
nand U10270 (N_10270,N_7028,N_7854);
nor U10271 (N_10271,N_8588,N_8712);
and U10272 (N_10272,N_7828,N_6606);
and U10273 (N_10273,N_8834,N_8146);
nand U10274 (N_10274,N_8765,N_8687);
and U10275 (N_10275,N_8673,N_6990);
xnor U10276 (N_10276,N_7918,N_7086);
nand U10277 (N_10277,N_8214,N_7795);
and U10278 (N_10278,N_6502,N_8013);
and U10279 (N_10279,N_6762,N_7674);
and U10280 (N_10280,N_6834,N_7443);
and U10281 (N_10281,N_8074,N_7994);
or U10282 (N_10282,N_6801,N_6209);
and U10283 (N_10283,N_7515,N_7505);
or U10284 (N_10284,N_8443,N_7262);
nand U10285 (N_10285,N_7653,N_6090);
nor U10286 (N_10286,N_6594,N_6781);
nand U10287 (N_10287,N_8536,N_8810);
and U10288 (N_10288,N_7719,N_6608);
nand U10289 (N_10289,N_7477,N_7816);
or U10290 (N_10290,N_6673,N_8656);
or U10291 (N_10291,N_7166,N_7036);
or U10292 (N_10292,N_7063,N_8693);
and U10293 (N_10293,N_6368,N_7523);
nand U10294 (N_10294,N_7270,N_7920);
nor U10295 (N_10295,N_6097,N_6409);
or U10296 (N_10296,N_6860,N_7510);
or U10297 (N_10297,N_7524,N_6131);
and U10298 (N_10298,N_6986,N_7050);
nor U10299 (N_10299,N_6143,N_7923);
nand U10300 (N_10300,N_6960,N_8989);
or U10301 (N_10301,N_6272,N_6646);
and U10302 (N_10302,N_7396,N_6198);
nor U10303 (N_10303,N_6397,N_7677);
or U10304 (N_10304,N_8340,N_6337);
nor U10305 (N_10305,N_7602,N_7958);
nor U10306 (N_10306,N_8218,N_6035);
nand U10307 (N_10307,N_6800,N_8885);
nor U10308 (N_10308,N_8843,N_8107);
nor U10309 (N_10309,N_8832,N_8491);
nand U10310 (N_10310,N_7468,N_8903);
or U10311 (N_10311,N_6835,N_8299);
xor U10312 (N_10312,N_7951,N_8045);
nand U10313 (N_10313,N_7239,N_7098);
nor U10314 (N_10314,N_7960,N_6523);
or U10315 (N_10315,N_7868,N_8993);
xnor U10316 (N_10316,N_6857,N_7040);
or U10317 (N_10317,N_6440,N_7188);
nand U10318 (N_10318,N_7247,N_6119);
or U10319 (N_10319,N_8449,N_6184);
and U10320 (N_10320,N_8933,N_7563);
nand U10321 (N_10321,N_6630,N_7648);
or U10322 (N_10322,N_7984,N_8014);
nand U10323 (N_10323,N_8767,N_7230);
nor U10324 (N_10324,N_6234,N_6730);
nand U10325 (N_10325,N_7215,N_8603);
or U10326 (N_10326,N_8275,N_8116);
and U10327 (N_10327,N_7573,N_7321);
or U10328 (N_10328,N_6361,N_7453);
and U10329 (N_10329,N_8751,N_7404);
nand U10330 (N_10330,N_7206,N_7108);
or U10331 (N_10331,N_7335,N_6238);
nor U10332 (N_10332,N_6050,N_8344);
and U10333 (N_10333,N_7013,N_6517);
xor U10334 (N_10334,N_6505,N_7532);
or U10335 (N_10335,N_7062,N_6486);
or U10336 (N_10336,N_7353,N_6911);
and U10337 (N_10337,N_8852,N_7153);
nand U10338 (N_10338,N_6244,N_6363);
or U10339 (N_10339,N_8123,N_7287);
nand U10340 (N_10340,N_7479,N_7096);
nand U10341 (N_10341,N_8806,N_7759);
nor U10342 (N_10342,N_8582,N_8640);
nor U10343 (N_10343,N_6384,N_6707);
or U10344 (N_10344,N_8235,N_8350);
nand U10345 (N_10345,N_6318,N_8997);
and U10346 (N_10346,N_8941,N_6211);
and U10347 (N_10347,N_8261,N_7125);
nand U10348 (N_10348,N_8858,N_6300);
and U10349 (N_10349,N_8259,N_8482);
and U10350 (N_10350,N_8106,N_6676);
and U10351 (N_10351,N_8402,N_8130);
xor U10352 (N_10352,N_8753,N_8167);
nor U10353 (N_10353,N_6648,N_7785);
or U10354 (N_10354,N_7787,N_8445);
xor U10355 (N_10355,N_7919,N_6482);
and U10356 (N_10356,N_8558,N_8439);
or U10357 (N_10357,N_8465,N_6054);
or U10358 (N_10358,N_6530,N_7875);
nor U10359 (N_10359,N_8528,N_7533);
or U10360 (N_10360,N_6269,N_7368);
nand U10361 (N_10361,N_8711,N_7402);
and U10362 (N_10362,N_6665,N_6898);
nor U10363 (N_10363,N_7504,N_7476);
nor U10364 (N_10364,N_7132,N_6247);
or U10365 (N_10365,N_7073,N_8873);
and U10366 (N_10366,N_8851,N_6956);
and U10367 (N_10367,N_8650,N_6412);
nor U10368 (N_10368,N_6294,N_7355);
nor U10369 (N_10369,N_6790,N_6852);
or U10370 (N_10370,N_6241,N_6501);
nand U10371 (N_10371,N_8860,N_6084);
and U10372 (N_10372,N_7124,N_7383);
nor U10373 (N_10373,N_6848,N_8607);
nor U10374 (N_10374,N_7082,N_8907);
and U10375 (N_10375,N_6524,N_7084);
and U10376 (N_10376,N_7222,N_7665);
and U10377 (N_10377,N_7516,N_7587);
or U10378 (N_10378,N_8243,N_8716);
nand U10379 (N_10379,N_7791,N_8532);
or U10380 (N_10380,N_7318,N_6616);
nor U10381 (N_10381,N_7647,N_7640);
nor U10382 (N_10382,N_6619,N_7872);
nand U10383 (N_10383,N_7445,N_8155);
nor U10384 (N_10384,N_6057,N_7981);
nand U10385 (N_10385,N_7142,N_8310);
nor U10386 (N_10386,N_7017,N_7530);
nor U10387 (N_10387,N_6779,N_7732);
or U10388 (N_10388,N_6539,N_6747);
and U10389 (N_10389,N_7762,N_8974);
nor U10390 (N_10390,N_8697,N_6713);
nor U10391 (N_10391,N_7282,N_6743);
nor U10392 (N_10392,N_7811,N_6989);
or U10393 (N_10393,N_8565,N_7514);
and U10394 (N_10394,N_7034,N_7852);
xnor U10395 (N_10395,N_6827,N_8251);
xor U10396 (N_10396,N_6973,N_8448);
or U10397 (N_10397,N_8738,N_7235);
nand U10398 (N_10398,N_6162,N_7388);
or U10399 (N_10399,N_8328,N_6303);
or U10400 (N_10400,N_7588,N_7436);
and U10401 (N_10401,N_6792,N_7000);
and U10402 (N_10402,N_8791,N_8508);
nand U10403 (N_10403,N_6796,N_8661);
nand U10404 (N_10404,N_7571,N_8083);
xnor U10405 (N_10405,N_6813,N_7352);
and U10406 (N_10406,N_7085,N_8371);
xor U10407 (N_10407,N_8401,N_8929);
nand U10408 (N_10408,N_6093,N_8591);
nor U10409 (N_10409,N_8473,N_8889);
or U10410 (N_10410,N_8213,N_8383);
xor U10411 (N_10411,N_7304,N_7796);
nand U10412 (N_10412,N_7936,N_7788);
nor U10413 (N_10413,N_8023,N_8702);
xor U10414 (N_10414,N_6659,N_7113);
nand U10415 (N_10415,N_8901,N_7659);
nand U10416 (N_10416,N_6257,N_6253);
nand U10417 (N_10417,N_6438,N_6133);
xor U10418 (N_10418,N_6772,N_7472);
nand U10419 (N_10419,N_6015,N_7497);
nor U10420 (N_10420,N_7509,N_8839);
nand U10421 (N_10421,N_8506,N_8569);
and U10422 (N_10422,N_8047,N_6044);
nor U10423 (N_10423,N_8819,N_6069);
nand U10424 (N_10424,N_7227,N_6528);
or U10425 (N_10425,N_6115,N_8874);
nor U10426 (N_10426,N_6177,N_7891);
or U10427 (N_10427,N_8618,N_7583);
and U10428 (N_10428,N_6430,N_6609);
and U10429 (N_10429,N_6703,N_8205);
nand U10430 (N_10430,N_7263,N_8325);
and U10431 (N_10431,N_8381,N_8415);
or U10432 (N_10432,N_6808,N_8857);
and U10433 (N_10433,N_6229,N_8958);
and U10434 (N_10434,N_7658,N_8868);
and U10435 (N_10435,N_7829,N_8608);
and U10436 (N_10436,N_6495,N_8129);
xnor U10437 (N_10437,N_6369,N_8817);
or U10438 (N_10438,N_6999,N_7566);
nor U10439 (N_10439,N_7309,N_8809);
or U10440 (N_10440,N_7999,N_6418);
nand U10441 (N_10441,N_7202,N_7164);
nor U10442 (N_10442,N_7120,N_7018);
nand U10443 (N_10443,N_6408,N_6901);
and U10444 (N_10444,N_7357,N_8324);
nor U10445 (N_10445,N_7508,N_8632);
and U10446 (N_10446,N_6087,N_6268);
nor U10447 (N_10447,N_8748,N_6013);
and U10448 (N_10448,N_7242,N_7726);
xnor U10449 (N_10449,N_7954,N_7883);
nand U10450 (N_10450,N_6461,N_8012);
or U10451 (N_10451,N_7117,N_6658);
or U10452 (N_10452,N_7069,N_7752);
xnor U10453 (N_10453,N_8879,N_6520);
nand U10454 (N_10454,N_6172,N_7903);
nand U10455 (N_10455,N_6512,N_8209);
or U10456 (N_10456,N_7409,N_6872);
nor U10457 (N_10457,N_7103,N_8334);
and U10458 (N_10458,N_6533,N_6663);
and U10459 (N_10459,N_8991,N_6120);
xor U10460 (N_10460,N_6332,N_6127);
and U10461 (N_10461,N_8382,N_8818);
nand U10462 (N_10462,N_7737,N_6038);
and U10463 (N_10463,N_7702,N_7319);
and U10464 (N_10464,N_6657,N_7268);
xnor U10465 (N_10465,N_7603,N_7421);
xor U10466 (N_10466,N_6518,N_7577);
and U10467 (N_10467,N_7041,N_8802);
nor U10468 (N_10468,N_6149,N_7864);
or U10469 (N_10469,N_6165,N_8206);
nor U10470 (N_10470,N_7834,N_6786);
or U10471 (N_10471,N_7456,N_6585);
nor U10472 (N_10472,N_8029,N_8597);
nand U10473 (N_10473,N_7928,N_6538);
nand U10474 (N_10474,N_8515,N_8026);
or U10475 (N_10475,N_6900,N_6909);
xnor U10476 (N_10476,N_8848,N_7008);
nand U10477 (N_10477,N_7112,N_7198);
nand U10478 (N_10478,N_6437,N_6978);
or U10479 (N_10479,N_7003,N_8073);
or U10480 (N_10480,N_8363,N_7048);
and U10481 (N_10481,N_6402,N_7846);
nand U10482 (N_10482,N_6587,N_8616);
nor U10483 (N_10483,N_7613,N_7716);
or U10484 (N_10484,N_6248,N_6243);
and U10485 (N_10485,N_7412,N_6675);
nand U10486 (N_10486,N_6775,N_6107);
and U10487 (N_10487,N_7876,N_6774);
nor U10488 (N_10488,N_7488,N_8075);
or U10489 (N_10489,N_7672,N_7991);
or U10490 (N_10490,N_6818,N_6174);
or U10491 (N_10491,N_7660,N_6636);
nand U10492 (N_10492,N_8544,N_6191);
or U10493 (N_10493,N_6401,N_7947);
nor U10494 (N_10494,N_7147,N_7531);
nand U10495 (N_10495,N_6640,N_6934);
xor U10496 (N_10496,N_8854,N_8391);
nand U10497 (N_10497,N_7100,N_7633);
nor U10498 (N_10498,N_7642,N_7405);
nor U10499 (N_10499,N_8967,N_7804);
xnor U10500 (N_10500,N_7622,N_7868);
xor U10501 (N_10501,N_8001,N_6588);
nor U10502 (N_10502,N_7264,N_8785);
or U10503 (N_10503,N_8232,N_8951);
nor U10504 (N_10504,N_7988,N_8534);
nor U10505 (N_10505,N_8324,N_7607);
and U10506 (N_10506,N_6275,N_7295);
nor U10507 (N_10507,N_7820,N_6770);
or U10508 (N_10508,N_6282,N_6005);
nor U10509 (N_10509,N_6272,N_8664);
nor U10510 (N_10510,N_8265,N_7545);
nand U10511 (N_10511,N_6535,N_6246);
or U10512 (N_10512,N_7148,N_7157);
nor U10513 (N_10513,N_8324,N_7779);
and U10514 (N_10514,N_6344,N_8768);
or U10515 (N_10515,N_7351,N_8158);
and U10516 (N_10516,N_6577,N_6121);
and U10517 (N_10517,N_8785,N_8116);
nand U10518 (N_10518,N_7591,N_8235);
nand U10519 (N_10519,N_7966,N_8472);
nand U10520 (N_10520,N_7968,N_6408);
nand U10521 (N_10521,N_6007,N_8363);
nor U10522 (N_10522,N_6666,N_6713);
xnor U10523 (N_10523,N_6910,N_7709);
nor U10524 (N_10524,N_7693,N_7760);
nand U10525 (N_10525,N_7207,N_8684);
and U10526 (N_10526,N_8769,N_6592);
and U10527 (N_10527,N_8867,N_8494);
and U10528 (N_10528,N_6903,N_7151);
and U10529 (N_10529,N_7452,N_8921);
and U10530 (N_10530,N_8681,N_8389);
and U10531 (N_10531,N_8241,N_6713);
and U10532 (N_10532,N_7639,N_8215);
or U10533 (N_10533,N_8658,N_8091);
or U10534 (N_10534,N_8754,N_6243);
or U10535 (N_10535,N_6695,N_7059);
nand U10536 (N_10536,N_6028,N_7582);
and U10537 (N_10537,N_7032,N_7474);
or U10538 (N_10538,N_8430,N_8449);
nand U10539 (N_10539,N_6022,N_8804);
or U10540 (N_10540,N_6143,N_8994);
nor U10541 (N_10541,N_8171,N_7676);
nand U10542 (N_10542,N_8681,N_6634);
nor U10543 (N_10543,N_8195,N_7457);
or U10544 (N_10544,N_7270,N_7190);
and U10545 (N_10545,N_7223,N_7137);
nor U10546 (N_10546,N_8831,N_8632);
and U10547 (N_10547,N_6681,N_8219);
nor U10548 (N_10548,N_7441,N_8018);
xor U10549 (N_10549,N_8953,N_8344);
nor U10550 (N_10550,N_7641,N_8710);
nand U10551 (N_10551,N_8689,N_6681);
nand U10552 (N_10552,N_6522,N_7751);
or U10553 (N_10553,N_7316,N_6553);
nand U10554 (N_10554,N_7437,N_7327);
xnor U10555 (N_10555,N_6384,N_8114);
nand U10556 (N_10556,N_7267,N_6209);
xnor U10557 (N_10557,N_8489,N_8538);
nor U10558 (N_10558,N_8100,N_8895);
or U10559 (N_10559,N_6846,N_7446);
nor U10560 (N_10560,N_8519,N_6621);
nand U10561 (N_10561,N_8488,N_8640);
or U10562 (N_10562,N_6972,N_7419);
nor U10563 (N_10563,N_8565,N_8138);
and U10564 (N_10564,N_8812,N_6223);
or U10565 (N_10565,N_7583,N_7863);
or U10566 (N_10566,N_7103,N_7281);
nand U10567 (N_10567,N_8013,N_7856);
xnor U10568 (N_10568,N_6372,N_7275);
nand U10569 (N_10569,N_7158,N_7188);
xnor U10570 (N_10570,N_6083,N_7942);
nand U10571 (N_10571,N_8958,N_8206);
and U10572 (N_10572,N_8374,N_7084);
nand U10573 (N_10573,N_8525,N_6871);
nor U10574 (N_10574,N_6559,N_8692);
nand U10575 (N_10575,N_6173,N_6314);
nor U10576 (N_10576,N_8396,N_7616);
or U10577 (N_10577,N_8277,N_7112);
nor U10578 (N_10578,N_6327,N_8323);
xor U10579 (N_10579,N_7987,N_6312);
or U10580 (N_10580,N_7867,N_8100);
and U10581 (N_10581,N_6413,N_7565);
nand U10582 (N_10582,N_6122,N_6844);
nand U10583 (N_10583,N_8556,N_7659);
or U10584 (N_10584,N_7267,N_7968);
or U10585 (N_10585,N_6140,N_6665);
nand U10586 (N_10586,N_6582,N_8944);
nand U10587 (N_10587,N_6322,N_7943);
nor U10588 (N_10588,N_8420,N_8099);
nor U10589 (N_10589,N_7984,N_7375);
or U10590 (N_10590,N_7534,N_6064);
and U10591 (N_10591,N_8740,N_7312);
nor U10592 (N_10592,N_7705,N_7536);
nand U10593 (N_10593,N_6067,N_8885);
or U10594 (N_10594,N_8955,N_8430);
or U10595 (N_10595,N_8138,N_8545);
nor U10596 (N_10596,N_6540,N_8236);
and U10597 (N_10597,N_6740,N_8115);
nand U10598 (N_10598,N_8525,N_7320);
or U10599 (N_10599,N_7136,N_6395);
nor U10600 (N_10600,N_6296,N_7006);
nand U10601 (N_10601,N_8168,N_6513);
or U10602 (N_10602,N_7466,N_8615);
nand U10603 (N_10603,N_8325,N_7646);
or U10604 (N_10604,N_6004,N_7985);
or U10605 (N_10605,N_6217,N_6067);
nor U10606 (N_10606,N_8339,N_7469);
nand U10607 (N_10607,N_8858,N_6446);
or U10608 (N_10608,N_7556,N_6402);
nor U10609 (N_10609,N_7133,N_8024);
nor U10610 (N_10610,N_6896,N_6025);
nor U10611 (N_10611,N_8492,N_6130);
and U10612 (N_10612,N_7616,N_6935);
xor U10613 (N_10613,N_7877,N_8874);
and U10614 (N_10614,N_6439,N_8616);
nor U10615 (N_10615,N_7242,N_7500);
and U10616 (N_10616,N_8439,N_6045);
and U10617 (N_10617,N_7115,N_6246);
and U10618 (N_10618,N_6480,N_7224);
or U10619 (N_10619,N_6437,N_7272);
nor U10620 (N_10620,N_7713,N_8134);
nor U10621 (N_10621,N_7592,N_6108);
xnor U10622 (N_10622,N_8186,N_7982);
and U10623 (N_10623,N_7983,N_6288);
nand U10624 (N_10624,N_6414,N_6350);
and U10625 (N_10625,N_7399,N_6567);
xnor U10626 (N_10626,N_6772,N_8594);
nand U10627 (N_10627,N_8046,N_6057);
nand U10628 (N_10628,N_6609,N_6623);
or U10629 (N_10629,N_7638,N_6422);
nor U10630 (N_10630,N_7617,N_6788);
nor U10631 (N_10631,N_8181,N_6541);
nand U10632 (N_10632,N_7494,N_6100);
and U10633 (N_10633,N_8111,N_8703);
nand U10634 (N_10634,N_6854,N_7501);
nor U10635 (N_10635,N_6927,N_6721);
or U10636 (N_10636,N_7775,N_7993);
and U10637 (N_10637,N_6875,N_8565);
or U10638 (N_10638,N_6262,N_6142);
nand U10639 (N_10639,N_6718,N_7317);
or U10640 (N_10640,N_8565,N_6084);
nand U10641 (N_10641,N_8529,N_8302);
nor U10642 (N_10642,N_7870,N_7837);
and U10643 (N_10643,N_6579,N_6927);
nand U10644 (N_10644,N_7314,N_8321);
nand U10645 (N_10645,N_6718,N_8085);
nand U10646 (N_10646,N_7498,N_7229);
and U10647 (N_10647,N_8326,N_8314);
and U10648 (N_10648,N_6731,N_8959);
and U10649 (N_10649,N_7944,N_8008);
and U10650 (N_10650,N_7693,N_7092);
nor U10651 (N_10651,N_8277,N_8496);
nor U10652 (N_10652,N_8936,N_6509);
or U10653 (N_10653,N_8793,N_8875);
xnor U10654 (N_10654,N_6427,N_7087);
nand U10655 (N_10655,N_8837,N_7798);
and U10656 (N_10656,N_8575,N_8586);
and U10657 (N_10657,N_8385,N_8022);
or U10658 (N_10658,N_7133,N_6566);
xnor U10659 (N_10659,N_7552,N_6849);
nand U10660 (N_10660,N_7069,N_6794);
or U10661 (N_10661,N_8503,N_8919);
nor U10662 (N_10662,N_7689,N_7571);
or U10663 (N_10663,N_7245,N_6028);
nor U10664 (N_10664,N_6274,N_8418);
nor U10665 (N_10665,N_7883,N_6879);
nand U10666 (N_10666,N_7814,N_8675);
and U10667 (N_10667,N_6824,N_6081);
or U10668 (N_10668,N_8857,N_6886);
xnor U10669 (N_10669,N_6012,N_6526);
nor U10670 (N_10670,N_7385,N_6644);
or U10671 (N_10671,N_7097,N_8915);
nor U10672 (N_10672,N_8901,N_8261);
nand U10673 (N_10673,N_8570,N_7561);
nor U10674 (N_10674,N_7828,N_7854);
and U10675 (N_10675,N_8173,N_8348);
or U10676 (N_10676,N_6054,N_6783);
and U10677 (N_10677,N_6470,N_8520);
nor U10678 (N_10678,N_7465,N_6833);
and U10679 (N_10679,N_7815,N_8471);
or U10680 (N_10680,N_7903,N_6961);
nand U10681 (N_10681,N_7881,N_6094);
or U10682 (N_10682,N_6639,N_8750);
xnor U10683 (N_10683,N_6763,N_7751);
nor U10684 (N_10684,N_6259,N_6086);
and U10685 (N_10685,N_6182,N_6407);
or U10686 (N_10686,N_6080,N_6381);
nand U10687 (N_10687,N_7452,N_6142);
nor U10688 (N_10688,N_8895,N_8279);
nor U10689 (N_10689,N_8844,N_8693);
or U10690 (N_10690,N_6474,N_8857);
nor U10691 (N_10691,N_6395,N_8138);
nor U10692 (N_10692,N_8587,N_7397);
and U10693 (N_10693,N_7584,N_7163);
or U10694 (N_10694,N_6977,N_8781);
nand U10695 (N_10695,N_7841,N_7239);
or U10696 (N_10696,N_6984,N_6002);
nand U10697 (N_10697,N_7630,N_8432);
xor U10698 (N_10698,N_7056,N_6834);
nor U10699 (N_10699,N_8738,N_8038);
nor U10700 (N_10700,N_7158,N_8761);
nand U10701 (N_10701,N_7996,N_7318);
nor U10702 (N_10702,N_6749,N_8584);
nor U10703 (N_10703,N_8171,N_6274);
nor U10704 (N_10704,N_8432,N_7707);
or U10705 (N_10705,N_6222,N_7146);
nand U10706 (N_10706,N_8756,N_8765);
nor U10707 (N_10707,N_7329,N_8503);
or U10708 (N_10708,N_8555,N_7002);
or U10709 (N_10709,N_6592,N_6456);
xnor U10710 (N_10710,N_8743,N_6044);
and U10711 (N_10711,N_7210,N_7944);
or U10712 (N_10712,N_7857,N_8406);
xor U10713 (N_10713,N_6354,N_7190);
and U10714 (N_10714,N_7288,N_7797);
or U10715 (N_10715,N_7917,N_8246);
or U10716 (N_10716,N_6190,N_6594);
and U10717 (N_10717,N_6896,N_8195);
or U10718 (N_10718,N_8693,N_8821);
and U10719 (N_10719,N_7180,N_7884);
xor U10720 (N_10720,N_8653,N_6866);
nand U10721 (N_10721,N_6768,N_7599);
nor U10722 (N_10722,N_8736,N_8444);
xor U10723 (N_10723,N_6156,N_7743);
xor U10724 (N_10724,N_7647,N_8170);
or U10725 (N_10725,N_7721,N_7371);
or U10726 (N_10726,N_6003,N_8993);
nor U10727 (N_10727,N_7771,N_7812);
or U10728 (N_10728,N_7360,N_7658);
and U10729 (N_10729,N_8240,N_8489);
or U10730 (N_10730,N_8837,N_7772);
xnor U10731 (N_10731,N_7342,N_6359);
nor U10732 (N_10732,N_8054,N_6119);
nor U10733 (N_10733,N_8853,N_7989);
nor U10734 (N_10734,N_8841,N_7105);
and U10735 (N_10735,N_6993,N_7591);
xor U10736 (N_10736,N_7663,N_7311);
nor U10737 (N_10737,N_6348,N_8482);
nand U10738 (N_10738,N_7495,N_8917);
and U10739 (N_10739,N_8528,N_6024);
and U10740 (N_10740,N_7143,N_8189);
xnor U10741 (N_10741,N_8937,N_6836);
nand U10742 (N_10742,N_6878,N_6977);
and U10743 (N_10743,N_8986,N_8684);
or U10744 (N_10744,N_6655,N_8571);
nor U10745 (N_10745,N_7254,N_7738);
nor U10746 (N_10746,N_8186,N_7988);
nor U10747 (N_10747,N_7666,N_8498);
nand U10748 (N_10748,N_8215,N_7562);
and U10749 (N_10749,N_7878,N_7798);
or U10750 (N_10750,N_6917,N_6376);
or U10751 (N_10751,N_7291,N_7879);
nor U10752 (N_10752,N_8428,N_7613);
and U10753 (N_10753,N_8783,N_8551);
nor U10754 (N_10754,N_6511,N_8752);
and U10755 (N_10755,N_7606,N_7755);
nand U10756 (N_10756,N_6315,N_8136);
or U10757 (N_10757,N_8791,N_6191);
or U10758 (N_10758,N_6103,N_7851);
or U10759 (N_10759,N_8545,N_6634);
or U10760 (N_10760,N_8421,N_7235);
and U10761 (N_10761,N_7945,N_7933);
and U10762 (N_10762,N_8479,N_7638);
xor U10763 (N_10763,N_7036,N_6785);
nand U10764 (N_10764,N_6141,N_6150);
nand U10765 (N_10765,N_6043,N_8459);
or U10766 (N_10766,N_8164,N_7570);
nor U10767 (N_10767,N_8955,N_6931);
nand U10768 (N_10768,N_6037,N_6437);
or U10769 (N_10769,N_8989,N_8008);
or U10770 (N_10770,N_7845,N_8402);
or U10771 (N_10771,N_8144,N_6492);
nand U10772 (N_10772,N_6724,N_7538);
nand U10773 (N_10773,N_7194,N_8125);
and U10774 (N_10774,N_7496,N_6093);
nor U10775 (N_10775,N_8103,N_7767);
and U10776 (N_10776,N_8410,N_8266);
nand U10777 (N_10777,N_8705,N_6633);
or U10778 (N_10778,N_6769,N_7784);
or U10779 (N_10779,N_7936,N_7241);
xnor U10780 (N_10780,N_7333,N_8188);
and U10781 (N_10781,N_7364,N_6875);
nand U10782 (N_10782,N_6613,N_7935);
nand U10783 (N_10783,N_6981,N_7865);
nor U10784 (N_10784,N_8379,N_6675);
xor U10785 (N_10785,N_6352,N_8947);
and U10786 (N_10786,N_8307,N_6957);
nand U10787 (N_10787,N_6100,N_6352);
nand U10788 (N_10788,N_7429,N_6254);
xor U10789 (N_10789,N_8898,N_8111);
or U10790 (N_10790,N_6685,N_6815);
nand U10791 (N_10791,N_8899,N_8023);
nor U10792 (N_10792,N_7897,N_7849);
and U10793 (N_10793,N_6054,N_7336);
xnor U10794 (N_10794,N_6534,N_7161);
and U10795 (N_10795,N_6716,N_7781);
or U10796 (N_10796,N_8372,N_6037);
nand U10797 (N_10797,N_7065,N_6702);
nor U10798 (N_10798,N_6692,N_7817);
or U10799 (N_10799,N_7658,N_6022);
and U10800 (N_10800,N_7532,N_6666);
and U10801 (N_10801,N_8829,N_6764);
and U10802 (N_10802,N_7719,N_8830);
and U10803 (N_10803,N_6875,N_6151);
nand U10804 (N_10804,N_7478,N_7512);
and U10805 (N_10805,N_6935,N_7634);
nand U10806 (N_10806,N_7657,N_8153);
xnor U10807 (N_10807,N_8023,N_8673);
or U10808 (N_10808,N_7055,N_8600);
or U10809 (N_10809,N_6985,N_6982);
nor U10810 (N_10810,N_8963,N_7368);
and U10811 (N_10811,N_7429,N_8970);
or U10812 (N_10812,N_6413,N_8137);
or U10813 (N_10813,N_8429,N_6365);
or U10814 (N_10814,N_7362,N_6326);
and U10815 (N_10815,N_6699,N_8712);
nor U10816 (N_10816,N_6280,N_6045);
and U10817 (N_10817,N_6541,N_8583);
or U10818 (N_10818,N_6190,N_6839);
and U10819 (N_10819,N_7514,N_7935);
xnor U10820 (N_10820,N_7199,N_7452);
and U10821 (N_10821,N_6580,N_8512);
and U10822 (N_10822,N_6183,N_7623);
nor U10823 (N_10823,N_8392,N_7830);
xnor U10824 (N_10824,N_6211,N_8346);
or U10825 (N_10825,N_7570,N_6582);
xor U10826 (N_10826,N_7584,N_7709);
or U10827 (N_10827,N_7750,N_6148);
or U10828 (N_10828,N_7098,N_8407);
nand U10829 (N_10829,N_6005,N_6545);
nor U10830 (N_10830,N_7592,N_8434);
or U10831 (N_10831,N_6008,N_8446);
or U10832 (N_10832,N_6797,N_6463);
nor U10833 (N_10833,N_8756,N_6790);
nand U10834 (N_10834,N_6448,N_8562);
nand U10835 (N_10835,N_6766,N_6237);
and U10836 (N_10836,N_6845,N_7982);
nand U10837 (N_10837,N_8317,N_6893);
or U10838 (N_10838,N_6922,N_7766);
nand U10839 (N_10839,N_8336,N_6566);
or U10840 (N_10840,N_8405,N_8233);
nor U10841 (N_10841,N_8136,N_7698);
nor U10842 (N_10842,N_8914,N_8594);
or U10843 (N_10843,N_8821,N_8652);
nor U10844 (N_10844,N_8452,N_8230);
or U10845 (N_10845,N_6550,N_6154);
nand U10846 (N_10846,N_8989,N_6652);
xnor U10847 (N_10847,N_8615,N_6050);
nor U10848 (N_10848,N_7570,N_8227);
and U10849 (N_10849,N_6546,N_8490);
nand U10850 (N_10850,N_7932,N_7945);
or U10851 (N_10851,N_7850,N_6138);
xor U10852 (N_10852,N_7227,N_7544);
xnor U10853 (N_10853,N_7620,N_7627);
and U10854 (N_10854,N_6466,N_8927);
nand U10855 (N_10855,N_7899,N_6993);
nor U10856 (N_10856,N_8862,N_6795);
and U10857 (N_10857,N_6456,N_8487);
or U10858 (N_10858,N_8306,N_8760);
or U10859 (N_10859,N_8786,N_6388);
nand U10860 (N_10860,N_7604,N_6664);
nor U10861 (N_10861,N_7273,N_7308);
or U10862 (N_10862,N_8542,N_8889);
xor U10863 (N_10863,N_7727,N_6447);
and U10864 (N_10864,N_6250,N_8556);
or U10865 (N_10865,N_6013,N_6892);
nor U10866 (N_10866,N_7297,N_8491);
nor U10867 (N_10867,N_6444,N_7261);
or U10868 (N_10868,N_8169,N_8566);
xor U10869 (N_10869,N_8364,N_6515);
and U10870 (N_10870,N_6786,N_7474);
and U10871 (N_10871,N_8374,N_6484);
or U10872 (N_10872,N_7587,N_7391);
and U10873 (N_10873,N_7903,N_6896);
or U10874 (N_10874,N_7465,N_6030);
nor U10875 (N_10875,N_7417,N_7606);
and U10876 (N_10876,N_8934,N_7008);
nand U10877 (N_10877,N_7637,N_7083);
and U10878 (N_10878,N_7579,N_8836);
or U10879 (N_10879,N_6884,N_7638);
or U10880 (N_10880,N_6415,N_8945);
nand U10881 (N_10881,N_7462,N_7806);
nand U10882 (N_10882,N_7955,N_6585);
or U10883 (N_10883,N_6024,N_8076);
nor U10884 (N_10884,N_6692,N_6274);
and U10885 (N_10885,N_8992,N_7487);
nand U10886 (N_10886,N_8677,N_8310);
or U10887 (N_10887,N_7569,N_7823);
nand U10888 (N_10888,N_6383,N_7152);
xor U10889 (N_10889,N_7803,N_6730);
nand U10890 (N_10890,N_8292,N_8518);
or U10891 (N_10891,N_6978,N_8249);
and U10892 (N_10892,N_6274,N_8040);
nor U10893 (N_10893,N_8429,N_8857);
nand U10894 (N_10894,N_8305,N_7845);
nand U10895 (N_10895,N_7671,N_6582);
nor U10896 (N_10896,N_6886,N_6330);
xnor U10897 (N_10897,N_8455,N_8669);
or U10898 (N_10898,N_8943,N_6564);
and U10899 (N_10899,N_7868,N_6627);
and U10900 (N_10900,N_6042,N_6730);
and U10901 (N_10901,N_7787,N_8602);
and U10902 (N_10902,N_7166,N_8917);
xnor U10903 (N_10903,N_6328,N_7722);
nand U10904 (N_10904,N_8520,N_6779);
or U10905 (N_10905,N_6836,N_7803);
and U10906 (N_10906,N_7214,N_6054);
nor U10907 (N_10907,N_7182,N_8770);
and U10908 (N_10908,N_7562,N_6945);
nor U10909 (N_10909,N_7663,N_6467);
nand U10910 (N_10910,N_6913,N_6117);
or U10911 (N_10911,N_7284,N_7822);
or U10912 (N_10912,N_7976,N_8023);
or U10913 (N_10913,N_8781,N_7950);
or U10914 (N_10914,N_8080,N_6800);
and U10915 (N_10915,N_8107,N_8493);
and U10916 (N_10916,N_7772,N_7747);
or U10917 (N_10917,N_8630,N_8877);
and U10918 (N_10918,N_6854,N_8581);
nand U10919 (N_10919,N_8368,N_6995);
nor U10920 (N_10920,N_7587,N_7047);
or U10921 (N_10921,N_7019,N_7549);
or U10922 (N_10922,N_7696,N_6274);
nor U10923 (N_10923,N_8787,N_6338);
or U10924 (N_10924,N_6041,N_6566);
nor U10925 (N_10925,N_7461,N_6328);
nand U10926 (N_10926,N_8355,N_8524);
xnor U10927 (N_10927,N_6865,N_8132);
and U10928 (N_10928,N_8442,N_7781);
xnor U10929 (N_10929,N_8697,N_7002);
nand U10930 (N_10930,N_8938,N_7113);
or U10931 (N_10931,N_7017,N_7427);
nand U10932 (N_10932,N_7354,N_6191);
and U10933 (N_10933,N_8429,N_8673);
and U10934 (N_10934,N_7515,N_7632);
nor U10935 (N_10935,N_6170,N_8662);
nand U10936 (N_10936,N_8610,N_6375);
xor U10937 (N_10937,N_7861,N_8384);
nand U10938 (N_10938,N_7621,N_8241);
nand U10939 (N_10939,N_7088,N_7913);
nor U10940 (N_10940,N_6419,N_7246);
nor U10941 (N_10941,N_7869,N_6805);
or U10942 (N_10942,N_8698,N_8885);
or U10943 (N_10943,N_7629,N_6988);
and U10944 (N_10944,N_6065,N_7876);
or U10945 (N_10945,N_6576,N_8186);
xor U10946 (N_10946,N_6386,N_8067);
nand U10947 (N_10947,N_7621,N_6033);
nor U10948 (N_10948,N_7057,N_8668);
xnor U10949 (N_10949,N_7024,N_6269);
and U10950 (N_10950,N_6201,N_6965);
or U10951 (N_10951,N_7668,N_7248);
and U10952 (N_10952,N_8253,N_8619);
xnor U10953 (N_10953,N_6354,N_6245);
nand U10954 (N_10954,N_7042,N_7549);
nor U10955 (N_10955,N_6141,N_8874);
and U10956 (N_10956,N_8138,N_7501);
nand U10957 (N_10957,N_7644,N_7994);
nor U10958 (N_10958,N_7747,N_6698);
nand U10959 (N_10959,N_7464,N_8971);
xor U10960 (N_10960,N_7504,N_7064);
nand U10961 (N_10961,N_7347,N_7158);
or U10962 (N_10962,N_7040,N_7025);
xor U10963 (N_10963,N_6189,N_7236);
nor U10964 (N_10964,N_6976,N_6846);
or U10965 (N_10965,N_6782,N_7315);
or U10966 (N_10966,N_7878,N_7104);
or U10967 (N_10967,N_6689,N_6280);
nand U10968 (N_10968,N_6649,N_7447);
and U10969 (N_10969,N_6983,N_6317);
nand U10970 (N_10970,N_8915,N_6674);
nand U10971 (N_10971,N_8926,N_6626);
nand U10972 (N_10972,N_8586,N_8848);
and U10973 (N_10973,N_8500,N_7661);
or U10974 (N_10974,N_7618,N_6168);
nand U10975 (N_10975,N_7219,N_6064);
or U10976 (N_10976,N_8390,N_8002);
xor U10977 (N_10977,N_7560,N_7898);
nand U10978 (N_10978,N_7873,N_6041);
and U10979 (N_10979,N_6802,N_7782);
nor U10980 (N_10980,N_6594,N_6855);
xor U10981 (N_10981,N_8399,N_8505);
nor U10982 (N_10982,N_8348,N_8668);
and U10983 (N_10983,N_7078,N_6394);
nor U10984 (N_10984,N_7660,N_6674);
and U10985 (N_10985,N_7260,N_6044);
nor U10986 (N_10986,N_8910,N_7488);
and U10987 (N_10987,N_7118,N_6235);
and U10988 (N_10988,N_7147,N_7820);
or U10989 (N_10989,N_7588,N_6411);
or U10990 (N_10990,N_8470,N_7464);
nand U10991 (N_10991,N_8671,N_7681);
nand U10992 (N_10992,N_6681,N_8158);
nand U10993 (N_10993,N_6087,N_7588);
nor U10994 (N_10994,N_6724,N_8911);
nor U10995 (N_10995,N_6917,N_7869);
nor U10996 (N_10996,N_8097,N_8957);
or U10997 (N_10997,N_8644,N_8091);
nor U10998 (N_10998,N_6657,N_8164);
and U10999 (N_10999,N_7947,N_8597);
xnor U11000 (N_11000,N_8958,N_8553);
nor U11001 (N_11001,N_6389,N_6123);
and U11002 (N_11002,N_6600,N_6940);
nand U11003 (N_11003,N_8854,N_6165);
or U11004 (N_11004,N_8869,N_6547);
xor U11005 (N_11005,N_7360,N_6218);
nand U11006 (N_11006,N_8372,N_7508);
and U11007 (N_11007,N_8742,N_6895);
nand U11008 (N_11008,N_8040,N_6391);
and U11009 (N_11009,N_8995,N_6661);
nor U11010 (N_11010,N_7112,N_6079);
and U11011 (N_11011,N_8276,N_6281);
and U11012 (N_11012,N_8253,N_7123);
nand U11013 (N_11013,N_7183,N_8856);
xnor U11014 (N_11014,N_8234,N_7148);
nand U11015 (N_11015,N_8360,N_6135);
and U11016 (N_11016,N_7285,N_6335);
nand U11017 (N_11017,N_8513,N_8458);
nand U11018 (N_11018,N_6183,N_8024);
nor U11019 (N_11019,N_8641,N_6264);
or U11020 (N_11020,N_8347,N_8995);
nor U11021 (N_11021,N_7139,N_6563);
and U11022 (N_11022,N_8611,N_6580);
nor U11023 (N_11023,N_8975,N_7376);
nor U11024 (N_11024,N_8598,N_7350);
nor U11025 (N_11025,N_7064,N_7262);
and U11026 (N_11026,N_8843,N_7165);
xor U11027 (N_11027,N_7363,N_6103);
nor U11028 (N_11028,N_6631,N_8703);
nor U11029 (N_11029,N_7402,N_6427);
or U11030 (N_11030,N_6125,N_6460);
nand U11031 (N_11031,N_7903,N_7810);
nor U11032 (N_11032,N_7930,N_8299);
nor U11033 (N_11033,N_7810,N_6856);
and U11034 (N_11034,N_7591,N_8499);
or U11035 (N_11035,N_7881,N_8141);
and U11036 (N_11036,N_6388,N_7123);
nand U11037 (N_11037,N_8959,N_6062);
nand U11038 (N_11038,N_8039,N_8464);
and U11039 (N_11039,N_7845,N_8890);
nor U11040 (N_11040,N_7039,N_6646);
nor U11041 (N_11041,N_8697,N_7712);
and U11042 (N_11042,N_8950,N_6778);
nand U11043 (N_11043,N_7166,N_6286);
and U11044 (N_11044,N_6678,N_7085);
or U11045 (N_11045,N_6015,N_7544);
or U11046 (N_11046,N_7391,N_6856);
nor U11047 (N_11047,N_7698,N_8792);
nor U11048 (N_11048,N_8837,N_6388);
nor U11049 (N_11049,N_8113,N_8121);
nand U11050 (N_11050,N_7787,N_7047);
or U11051 (N_11051,N_7776,N_7535);
nor U11052 (N_11052,N_6313,N_6019);
and U11053 (N_11053,N_6720,N_8579);
or U11054 (N_11054,N_7318,N_8648);
nor U11055 (N_11055,N_7042,N_7592);
nand U11056 (N_11056,N_7645,N_6343);
and U11057 (N_11057,N_7218,N_7313);
and U11058 (N_11058,N_8199,N_6050);
and U11059 (N_11059,N_8423,N_8995);
nand U11060 (N_11060,N_6193,N_6699);
or U11061 (N_11061,N_8991,N_6003);
or U11062 (N_11062,N_7605,N_7253);
nand U11063 (N_11063,N_8667,N_6542);
nor U11064 (N_11064,N_8099,N_8475);
xor U11065 (N_11065,N_6970,N_8482);
or U11066 (N_11066,N_8582,N_7425);
xor U11067 (N_11067,N_7174,N_7650);
xnor U11068 (N_11068,N_6318,N_8543);
nor U11069 (N_11069,N_7836,N_6680);
or U11070 (N_11070,N_8518,N_8920);
nor U11071 (N_11071,N_7125,N_8819);
and U11072 (N_11072,N_7382,N_7300);
nand U11073 (N_11073,N_7889,N_7877);
and U11074 (N_11074,N_8957,N_8338);
or U11075 (N_11075,N_7777,N_7205);
nand U11076 (N_11076,N_6279,N_7354);
or U11077 (N_11077,N_6172,N_6508);
or U11078 (N_11078,N_8766,N_8729);
nor U11079 (N_11079,N_7068,N_8822);
nand U11080 (N_11080,N_8133,N_8696);
xnor U11081 (N_11081,N_6228,N_6276);
nor U11082 (N_11082,N_8430,N_7397);
xor U11083 (N_11083,N_7079,N_6179);
and U11084 (N_11084,N_8309,N_6358);
nor U11085 (N_11085,N_8384,N_7951);
nand U11086 (N_11086,N_7339,N_8710);
and U11087 (N_11087,N_8430,N_7892);
nor U11088 (N_11088,N_7264,N_8061);
nand U11089 (N_11089,N_8401,N_7135);
or U11090 (N_11090,N_8502,N_8440);
or U11091 (N_11091,N_8091,N_6328);
nor U11092 (N_11092,N_8714,N_6069);
nand U11093 (N_11093,N_7108,N_8803);
nand U11094 (N_11094,N_8146,N_8440);
nor U11095 (N_11095,N_7682,N_7383);
nor U11096 (N_11096,N_8186,N_8960);
and U11097 (N_11097,N_6888,N_6193);
nand U11098 (N_11098,N_8624,N_8993);
nor U11099 (N_11099,N_8574,N_6187);
nor U11100 (N_11100,N_8799,N_8121);
nand U11101 (N_11101,N_7153,N_8305);
and U11102 (N_11102,N_7422,N_7391);
or U11103 (N_11103,N_6075,N_6193);
xnor U11104 (N_11104,N_7476,N_6060);
nor U11105 (N_11105,N_7189,N_7485);
nand U11106 (N_11106,N_6431,N_6605);
or U11107 (N_11107,N_6791,N_7409);
or U11108 (N_11108,N_6656,N_6976);
nor U11109 (N_11109,N_6499,N_8387);
or U11110 (N_11110,N_8443,N_8595);
xor U11111 (N_11111,N_7455,N_8638);
nor U11112 (N_11112,N_8498,N_6730);
or U11113 (N_11113,N_7516,N_6762);
or U11114 (N_11114,N_6466,N_8671);
nand U11115 (N_11115,N_7796,N_8551);
or U11116 (N_11116,N_7566,N_7282);
or U11117 (N_11117,N_7492,N_8327);
nand U11118 (N_11118,N_6328,N_6918);
or U11119 (N_11119,N_7200,N_7383);
nand U11120 (N_11120,N_8137,N_7650);
nor U11121 (N_11121,N_6916,N_6546);
nand U11122 (N_11122,N_8346,N_8849);
and U11123 (N_11123,N_6937,N_8445);
nand U11124 (N_11124,N_6781,N_6243);
or U11125 (N_11125,N_7819,N_7697);
and U11126 (N_11126,N_7058,N_8670);
and U11127 (N_11127,N_7186,N_8245);
or U11128 (N_11128,N_6126,N_6611);
or U11129 (N_11129,N_6480,N_8544);
nand U11130 (N_11130,N_7462,N_8992);
nor U11131 (N_11131,N_7076,N_8778);
and U11132 (N_11132,N_6749,N_7533);
and U11133 (N_11133,N_8636,N_8055);
nor U11134 (N_11134,N_6352,N_7163);
nand U11135 (N_11135,N_7885,N_7599);
and U11136 (N_11136,N_7254,N_7011);
or U11137 (N_11137,N_7266,N_6588);
and U11138 (N_11138,N_7251,N_6999);
and U11139 (N_11139,N_6958,N_8719);
nor U11140 (N_11140,N_8543,N_6735);
or U11141 (N_11141,N_6440,N_6578);
or U11142 (N_11142,N_7537,N_7732);
or U11143 (N_11143,N_8371,N_6967);
or U11144 (N_11144,N_7587,N_7070);
nand U11145 (N_11145,N_7733,N_8018);
or U11146 (N_11146,N_7202,N_8090);
and U11147 (N_11147,N_7691,N_6716);
and U11148 (N_11148,N_8698,N_7735);
nand U11149 (N_11149,N_6310,N_8638);
nand U11150 (N_11150,N_6881,N_6515);
nor U11151 (N_11151,N_8254,N_8322);
nand U11152 (N_11152,N_6832,N_7992);
xnor U11153 (N_11153,N_7373,N_6291);
nor U11154 (N_11154,N_6548,N_7266);
and U11155 (N_11155,N_7593,N_8631);
and U11156 (N_11156,N_6900,N_8318);
nand U11157 (N_11157,N_8755,N_7403);
or U11158 (N_11158,N_8886,N_6948);
nand U11159 (N_11159,N_7564,N_7692);
and U11160 (N_11160,N_7793,N_6250);
nor U11161 (N_11161,N_8033,N_6124);
and U11162 (N_11162,N_7834,N_6492);
and U11163 (N_11163,N_7519,N_7268);
or U11164 (N_11164,N_6177,N_7173);
xnor U11165 (N_11165,N_8706,N_8277);
nor U11166 (N_11166,N_8534,N_8392);
and U11167 (N_11167,N_6631,N_8463);
or U11168 (N_11168,N_8022,N_7750);
and U11169 (N_11169,N_8451,N_7879);
and U11170 (N_11170,N_7777,N_8123);
nand U11171 (N_11171,N_8404,N_8887);
or U11172 (N_11172,N_8809,N_6656);
nor U11173 (N_11173,N_6552,N_7452);
nor U11174 (N_11174,N_8710,N_8730);
nand U11175 (N_11175,N_7490,N_7001);
nor U11176 (N_11176,N_7294,N_6391);
nand U11177 (N_11177,N_8264,N_7587);
or U11178 (N_11178,N_8961,N_6612);
nor U11179 (N_11179,N_7850,N_8665);
and U11180 (N_11180,N_6244,N_6031);
or U11181 (N_11181,N_7647,N_6496);
and U11182 (N_11182,N_6974,N_8218);
or U11183 (N_11183,N_6420,N_8748);
or U11184 (N_11184,N_8076,N_6202);
nor U11185 (N_11185,N_8779,N_8617);
nor U11186 (N_11186,N_7490,N_8287);
or U11187 (N_11187,N_8196,N_6591);
nand U11188 (N_11188,N_6048,N_7870);
or U11189 (N_11189,N_8483,N_7856);
and U11190 (N_11190,N_8647,N_6373);
or U11191 (N_11191,N_6714,N_8895);
or U11192 (N_11192,N_7221,N_7434);
and U11193 (N_11193,N_8436,N_7541);
nor U11194 (N_11194,N_6689,N_7051);
nor U11195 (N_11195,N_8688,N_6682);
xor U11196 (N_11196,N_8940,N_7729);
and U11197 (N_11197,N_7000,N_7666);
nor U11198 (N_11198,N_6787,N_7816);
or U11199 (N_11199,N_6399,N_6339);
and U11200 (N_11200,N_7178,N_8671);
nor U11201 (N_11201,N_7694,N_7948);
or U11202 (N_11202,N_8535,N_8630);
or U11203 (N_11203,N_8622,N_6418);
nand U11204 (N_11204,N_8401,N_6945);
nor U11205 (N_11205,N_6095,N_6043);
or U11206 (N_11206,N_7753,N_7152);
and U11207 (N_11207,N_8604,N_6886);
nand U11208 (N_11208,N_7897,N_6488);
nor U11209 (N_11209,N_8641,N_8850);
or U11210 (N_11210,N_8839,N_7007);
and U11211 (N_11211,N_7246,N_8338);
xor U11212 (N_11212,N_6670,N_7129);
or U11213 (N_11213,N_7447,N_8367);
nor U11214 (N_11214,N_6636,N_8354);
nor U11215 (N_11215,N_6418,N_8429);
nor U11216 (N_11216,N_7739,N_8130);
or U11217 (N_11217,N_8687,N_6071);
or U11218 (N_11218,N_6319,N_7589);
nand U11219 (N_11219,N_7504,N_7222);
or U11220 (N_11220,N_6348,N_7515);
and U11221 (N_11221,N_7784,N_7877);
nor U11222 (N_11222,N_6438,N_6279);
or U11223 (N_11223,N_6710,N_6748);
xor U11224 (N_11224,N_6161,N_6953);
and U11225 (N_11225,N_7131,N_7297);
nand U11226 (N_11226,N_7105,N_6684);
nor U11227 (N_11227,N_8166,N_6411);
xnor U11228 (N_11228,N_8479,N_6827);
and U11229 (N_11229,N_7616,N_7009);
nand U11230 (N_11230,N_7090,N_7889);
nand U11231 (N_11231,N_6614,N_8834);
nand U11232 (N_11232,N_7782,N_8547);
nand U11233 (N_11233,N_8319,N_7901);
nor U11234 (N_11234,N_6273,N_6036);
nand U11235 (N_11235,N_8078,N_8180);
or U11236 (N_11236,N_8109,N_8036);
and U11237 (N_11237,N_7097,N_7435);
or U11238 (N_11238,N_6978,N_6359);
or U11239 (N_11239,N_7497,N_7450);
or U11240 (N_11240,N_6619,N_8357);
nand U11241 (N_11241,N_7313,N_8445);
nor U11242 (N_11242,N_7157,N_8950);
or U11243 (N_11243,N_7181,N_8905);
nand U11244 (N_11244,N_7821,N_8931);
xnor U11245 (N_11245,N_7471,N_6348);
nor U11246 (N_11246,N_6159,N_8082);
nand U11247 (N_11247,N_8035,N_7972);
and U11248 (N_11248,N_7772,N_7094);
and U11249 (N_11249,N_8998,N_6820);
nor U11250 (N_11250,N_8022,N_7474);
or U11251 (N_11251,N_8266,N_6625);
nand U11252 (N_11252,N_7822,N_8993);
and U11253 (N_11253,N_6051,N_8792);
or U11254 (N_11254,N_7082,N_7726);
or U11255 (N_11255,N_7090,N_7604);
and U11256 (N_11256,N_7403,N_7227);
and U11257 (N_11257,N_8945,N_6968);
and U11258 (N_11258,N_8850,N_7482);
nor U11259 (N_11259,N_7566,N_6624);
and U11260 (N_11260,N_6524,N_6035);
nand U11261 (N_11261,N_7744,N_6457);
and U11262 (N_11262,N_7593,N_6804);
nor U11263 (N_11263,N_8154,N_6683);
and U11264 (N_11264,N_7560,N_8325);
and U11265 (N_11265,N_6156,N_8306);
nor U11266 (N_11266,N_8858,N_6495);
and U11267 (N_11267,N_8050,N_7828);
or U11268 (N_11268,N_8292,N_7486);
nand U11269 (N_11269,N_8037,N_6319);
nor U11270 (N_11270,N_8200,N_7268);
and U11271 (N_11271,N_7165,N_8001);
and U11272 (N_11272,N_6701,N_8944);
or U11273 (N_11273,N_8778,N_6420);
nand U11274 (N_11274,N_6102,N_7902);
xnor U11275 (N_11275,N_8689,N_6013);
nor U11276 (N_11276,N_6076,N_8605);
or U11277 (N_11277,N_7591,N_7216);
or U11278 (N_11278,N_8354,N_6520);
nand U11279 (N_11279,N_8974,N_7647);
or U11280 (N_11280,N_7125,N_8507);
xor U11281 (N_11281,N_8721,N_7101);
nor U11282 (N_11282,N_8961,N_8945);
xnor U11283 (N_11283,N_8128,N_8883);
nand U11284 (N_11284,N_7405,N_6479);
nand U11285 (N_11285,N_8214,N_6777);
xnor U11286 (N_11286,N_6758,N_8377);
and U11287 (N_11287,N_6690,N_8468);
nor U11288 (N_11288,N_8459,N_8750);
and U11289 (N_11289,N_7119,N_6629);
xor U11290 (N_11290,N_8728,N_6472);
xnor U11291 (N_11291,N_8607,N_7460);
nor U11292 (N_11292,N_6171,N_7393);
and U11293 (N_11293,N_7094,N_7113);
or U11294 (N_11294,N_7898,N_8019);
nor U11295 (N_11295,N_6338,N_7628);
and U11296 (N_11296,N_7367,N_7873);
or U11297 (N_11297,N_7347,N_8009);
or U11298 (N_11298,N_8391,N_7590);
xor U11299 (N_11299,N_7078,N_7999);
nand U11300 (N_11300,N_8316,N_8730);
or U11301 (N_11301,N_7699,N_7052);
xnor U11302 (N_11302,N_7072,N_7758);
xnor U11303 (N_11303,N_8459,N_6811);
xor U11304 (N_11304,N_7501,N_7399);
nor U11305 (N_11305,N_8151,N_8484);
nor U11306 (N_11306,N_7045,N_7610);
nand U11307 (N_11307,N_6665,N_7583);
xor U11308 (N_11308,N_6256,N_8784);
and U11309 (N_11309,N_7786,N_8900);
xnor U11310 (N_11310,N_8416,N_8485);
nand U11311 (N_11311,N_6788,N_6852);
and U11312 (N_11312,N_6746,N_8623);
and U11313 (N_11313,N_7695,N_8066);
or U11314 (N_11314,N_8719,N_7604);
nor U11315 (N_11315,N_6137,N_6152);
nor U11316 (N_11316,N_6540,N_6626);
nand U11317 (N_11317,N_6146,N_7882);
or U11318 (N_11318,N_7655,N_7342);
nor U11319 (N_11319,N_6101,N_6563);
nor U11320 (N_11320,N_7870,N_7579);
and U11321 (N_11321,N_6993,N_7292);
and U11322 (N_11322,N_8205,N_7723);
nand U11323 (N_11323,N_8618,N_7188);
nand U11324 (N_11324,N_6703,N_7520);
nand U11325 (N_11325,N_6483,N_6138);
nand U11326 (N_11326,N_8733,N_6187);
or U11327 (N_11327,N_8132,N_8547);
xor U11328 (N_11328,N_6817,N_8457);
xnor U11329 (N_11329,N_8623,N_7104);
nand U11330 (N_11330,N_8747,N_8238);
xor U11331 (N_11331,N_7453,N_6040);
nand U11332 (N_11332,N_8515,N_7160);
and U11333 (N_11333,N_7735,N_6031);
or U11334 (N_11334,N_6684,N_6519);
and U11335 (N_11335,N_7685,N_6393);
nor U11336 (N_11336,N_6536,N_8812);
nor U11337 (N_11337,N_6285,N_7027);
nand U11338 (N_11338,N_7638,N_6613);
xnor U11339 (N_11339,N_6100,N_8318);
and U11340 (N_11340,N_8332,N_6377);
nor U11341 (N_11341,N_7198,N_6264);
nand U11342 (N_11342,N_8785,N_8743);
xnor U11343 (N_11343,N_8033,N_8832);
and U11344 (N_11344,N_8730,N_8340);
nor U11345 (N_11345,N_7804,N_7414);
nand U11346 (N_11346,N_7381,N_8993);
nor U11347 (N_11347,N_6320,N_8264);
nand U11348 (N_11348,N_6419,N_6076);
and U11349 (N_11349,N_8101,N_7508);
xnor U11350 (N_11350,N_7174,N_6157);
nand U11351 (N_11351,N_7957,N_6866);
and U11352 (N_11352,N_7016,N_7203);
nand U11353 (N_11353,N_7056,N_7337);
nand U11354 (N_11354,N_8392,N_6842);
xor U11355 (N_11355,N_7397,N_8936);
xnor U11356 (N_11356,N_6648,N_7552);
nand U11357 (N_11357,N_8122,N_6733);
nor U11358 (N_11358,N_6879,N_8405);
nand U11359 (N_11359,N_7694,N_8390);
xnor U11360 (N_11360,N_6621,N_6046);
xnor U11361 (N_11361,N_8349,N_7015);
or U11362 (N_11362,N_7223,N_7070);
xor U11363 (N_11363,N_8881,N_6019);
or U11364 (N_11364,N_8087,N_6582);
and U11365 (N_11365,N_6867,N_8725);
nor U11366 (N_11366,N_6697,N_8655);
or U11367 (N_11367,N_8084,N_8979);
and U11368 (N_11368,N_6672,N_7372);
nand U11369 (N_11369,N_8127,N_6203);
and U11370 (N_11370,N_6947,N_7516);
nor U11371 (N_11371,N_8711,N_7484);
nor U11372 (N_11372,N_6733,N_8401);
and U11373 (N_11373,N_6789,N_8496);
and U11374 (N_11374,N_7454,N_8349);
xnor U11375 (N_11375,N_7437,N_6733);
or U11376 (N_11376,N_6156,N_7794);
nand U11377 (N_11377,N_6281,N_7973);
and U11378 (N_11378,N_6384,N_7977);
nand U11379 (N_11379,N_6356,N_8775);
and U11380 (N_11380,N_7415,N_8106);
and U11381 (N_11381,N_8151,N_6544);
nand U11382 (N_11382,N_7147,N_8652);
nand U11383 (N_11383,N_8285,N_6155);
and U11384 (N_11384,N_7496,N_7224);
nor U11385 (N_11385,N_7365,N_8899);
nor U11386 (N_11386,N_8544,N_6460);
xor U11387 (N_11387,N_6111,N_8376);
or U11388 (N_11388,N_7499,N_8332);
nor U11389 (N_11389,N_6162,N_7015);
nand U11390 (N_11390,N_6680,N_8376);
nor U11391 (N_11391,N_8367,N_8872);
nand U11392 (N_11392,N_8342,N_8931);
or U11393 (N_11393,N_7613,N_6493);
and U11394 (N_11394,N_6210,N_7659);
nand U11395 (N_11395,N_8407,N_6556);
and U11396 (N_11396,N_8986,N_6302);
nor U11397 (N_11397,N_7685,N_6990);
and U11398 (N_11398,N_6846,N_8153);
or U11399 (N_11399,N_7423,N_6924);
or U11400 (N_11400,N_8485,N_7615);
nand U11401 (N_11401,N_7411,N_8824);
nand U11402 (N_11402,N_6963,N_8946);
and U11403 (N_11403,N_8880,N_6083);
nand U11404 (N_11404,N_6198,N_6911);
and U11405 (N_11405,N_7578,N_7898);
nand U11406 (N_11406,N_8552,N_6985);
xor U11407 (N_11407,N_7743,N_8306);
nor U11408 (N_11408,N_7804,N_6598);
and U11409 (N_11409,N_6624,N_6278);
nand U11410 (N_11410,N_7867,N_7906);
nand U11411 (N_11411,N_8432,N_8652);
nand U11412 (N_11412,N_6048,N_6905);
nand U11413 (N_11413,N_6878,N_7972);
nand U11414 (N_11414,N_7232,N_8721);
and U11415 (N_11415,N_6055,N_7182);
and U11416 (N_11416,N_8276,N_7742);
or U11417 (N_11417,N_7131,N_7935);
or U11418 (N_11418,N_7308,N_6499);
xnor U11419 (N_11419,N_7354,N_6365);
xnor U11420 (N_11420,N_7311,N_7090);
nand U11421 (N_11421,N_8055,N_7720);
and U11422 (N_11422,N_7085,N_8412);
nor U11423 (N_11423,N_7170,N_6504);
nor U11424 (N_11424,N_8746,N_7027);
nor U11425 (N_11425,N_7993,N_7122);
nand U11426 (N_11426,N_7825,N_7132);
and U11427 (N_11427,N_6572,N_8405);
xor U11428 (N_11428,N_6921,N_8669);
or U11429 (N_11429,N_8218,N_8249);
nand U11430 (N_11430,N_8523,N_8331);
and U11431 (N_11431,N_7392,N_8460);
or U11432 (N_11432,N_7130,N_7092);
and U11433 (N_11433,N_6266,N_6128);
nand U11434 (N_11434,N_7352,N_6703);
nor U11435 (N_11435,N_7702,N_8035);
xnor U11436 (N_11436,N_6893,N_6680);
or U11437 (N_11437,N_6980,N_8702);
nand U11438 (N_11438,N_7119,N_8057);
nand U11439 (N_11439,N_7190,N_8469);
or U11440 (N_11440,N_7213,N_6627);
nor U11441 (N_11441,N_8321,N_8019);
nand U11442 (N_11442,N_8494,N_6045);
and U11443 (N_11443,N_6999,N_6709);
nand U11444 (N_11444,N_7286,N_7758);
nand U11445 (N_11445,N_8503,N_8207);
nor U11446 (N_11446,N_8260,N_7864);
nand U11447 (N_11447,N_7285,N_8366);
and U11448 (N_11448,N_8966,N_7244);
nor U11449 (N_11449,N_6536,N_7582);
nor U11450 (N_11450,N_6607,N_6916);
nor U11451 (N_11451,N_7917,N_8235);
and U11452 (N_11452,N_6700,N_8322);
or U11453 (N_11453,N_6212,N_8378);
nor U11454 (N_11454,N_8792,N_6282);
and U11455 (N_11455,N_8969,N_7957);
xnor U11456 (N_11456,N_8000,N_7135);
xor U11457 (N_11457,N_6648,N_7788);
nand U11458 (N_11458,N_6632,N_6024);
or U11459 (N_11459,N_6282,N_7806);
nor U11460 (N_11460,N_8917,N_7850);
and U11461 (N_11461,N_8673,N_6139);
nor U11462 (N_11462,N_6381,N_8339);
xnor U11463 (N_11463,N_6698,N_7474);
and U11464 (N_11464,N_7722,N_7270);
nor U11465 (N_11465,N_6428,N_6080);
nand U11466 (N_11466,N_8734,N_7958);
or U11467 (N_11467,N_6852,N_6188);
or U11468 (N_11468,N_7796,N_7819);
nand U11469 (N_11469,N_7283,N_8074);
nand U11470 (N_11470,N_6229,N_6667);
nand U11471 (N_11471,N_8446,N_8532);
nand U11472 (N_11472,N_7863,N_7907);
or U11473 (N_11473,N_7891,N_6054);
nand U11474 (N_11474,N_6373,N_8904);
nor U11475 (N_11475,N_6480,N_8179);
and U11476 (N_11476,N_6215,N_8159);
nor U11477 (N_11477,N_8053,N_8502);
or U11478 (N_11478,N_7512,N_6254);
or U11479 (N_11479,N_8162,N_6759);
xor U11480 (N_11480,N_8191,N_8871);
nand U11481 (N_11481,N_8173,N_7254);
and U11482 (N_11482,N_7085,N_6089);
nor U11483 (N_11483,N_6810,N_8108);
nor U11484 (N_11484,N_8179,N_8289);
or U11485 (N_11485,N_7489,N_6033);
or U11486 (N_11486,N_7112,N_6992);
or U11487 (N_11487,N_6004,N_7646);
or U11488 (N_11488,N_6215,N_7001);
nor U11489 (N_11489,N_6006,N_6983);
or U11490 (N_11490,N_6264,N_8872);
and U11491 (N_11491,N_8562,N_6153);
or U11492 (N_11492,N_7258,N_6280);
and U11493 (N_11493,N_7958,N_6353);
nor U11494 (N_11494,N_6894,N_6950);
and U11495 (N_11495,N_7563,N_7885);
or U11496 (N_11496,N_8713,N_8027);
or U11497 (N_11497,N_6322,N_8764);
xnor U11498 (N_11498,N_8909,N_7059);
nand U11499 (N_11499,N_6607,N_8970);
nand U11500 (N_11500,N_7105,N_8292);
and U11501 (N_11501,N_6206,N_8412);
and U11502 (N_11502,N_7903,N_6476);
or U11503 (N_11503,N_8428,N_6123);
nor U11504 (N_11504,N_8551,N_8332);
and U11505 (N_11505,N_6358,N_6803);
nor U11506 (N_11506,N_8024,N_8585);
and U11507 (N_11507,N_7958,N_8454);
nor U11508 (N_11508,N_6667,N_8413);
nor U11509 (N_11509,N_7525,N_7315);
and U11510 (N_11510,N_8554,N_6132);
and U11511 (N_11511,N_6525,N_7716);
nor U11512 (N_11512,N_8835,N_7124);
xor U11513 (N_11513,N_7327,N_7398);
nand U11514 (N_11514,N_8070,N_7332);
and U11515 (N_11515,N_7184,N_7536);
nand U11516 (N_11516,N_8790,N_8299);
and U11517 (N_11517,N_8764,N_8516);
and U11518 (N_11518,N_7410,N_6834);
or U11519 (N_11519,N_7735,N_8934);
nand U11520 (N_11520,N_7934,N_7938);
xor U11521 (N_11521,N_7915,N_8889);
xnor U11522 (N_11522,N_8073,N_7006);
nor U11523 (N_11523,N_7492,N_6204);
nand U11524 (N_11524,N_8932,N_6366);
or U11525 (N_11525,N_7602,N_7304);
nand U11526 (N_11526,N_6333,N_7440);
xor U11527 (N_11527,N_6319,N_7019);
nor U11528 (N_11528,N_7577,N_7277);
nand U11529 (N_11529,N_7439,N_6595);
nor U11530 (N_11530,N_8845,N_8452);
and U11531 (N_11531,N_6161,N_6346);
and U11532 (N_11532,N_6021,N_6935);
nor U11533 (N_11533,N_8352,N_8188);
nor U11534 (N_11534,N_6498,N_6482);
xnor U11535 (N_11535,N_8294,N_7578);
nor U11536 (N_11536,N_6950,N_7938);
nor U11537 (N_11537,N_8763,N_6655);
xnor U11538 (N_11538,N_6216,N_6107);
nand U11539 (N_11539,N_6096,N_6270);
and U11540 (N_11540,N_6057,N_6378);
or U11541 (N_11541,N_7892,N_6866);
and U11542 (N_11542,N_6650,N_6280);
and U11543 (N_11543,N_8540,N_7866);
and U11544 (N_11544,N_8402,N_7990);
nand U11545 (N_11545,N_7889,N_6027);
and U11546 (N_11546,N_7768,N_7895);
and U11547 (N_11547,N_6205,N_6076);
and U11548 (N_11548,N_6655,N_6297);
and U11549 (N_11549,N_7679,N_6577);
xnor U11550 (N_11550,N_8075,N_8267);
nand U11551 (N_11551,N_6231,N_7618);
nor U11552 (N_11552,N_7653,N_6501);
or U11553 (N_11553,N_8315,N_8233);
or U11554 (N_11554,N_8563,N_7951);
nor U11555 (N_11555,N_6203,N_6447);
and U11556 (N_11556,N_8335,N_7463);
and U11557 (N_11557,N_8352,N_8245);
nor U11558 (N_11558,N_7667,N_7303);
nand U11559 (N_11559,N_6568,N_6782);
and U11560 (N_11560,N_8292,N_8035);
nor U11561 (N_11561,N_7148,N_6481);
nor U11562 (N_11562,N_6699,N_8940);
nand U11563 (N_11563,N_6117,N_8874);
and U11564 (N_11564,N_7655,N_7497);
and U11565 (N_11565,N_8546,N_6637);
and U11566 (N_11566,N_8322,N_8749);
xor U11567 (N_11567,N_7715,N_8927);
nand U11568 (N_11568,N_7231,N_8514);
or U11569 (N_11569,N_8243,N_8537);
xor U11570 (N_11570,N_6815,N_8784);
or U11571 (N_11571,N_7337,N_8995);
or U11572 (N_11572,N_7622,N_8014);
nor U11573 (N_11573,N_7047,N_7729);
or U11574 (N_11574,N_8019,N_8690);
nand U11575 (N_11575,N_7728,N_7000);
nor U11576 (N_11576,N_7714,N_6048);
nand U11577 (N_11577,N_8660,N_6525);
nand U11578 (N_11578,N_8612,N_8730);
nand U11579 (N_11579,N_6104,N_7141);
and U11580 (N_11580,N_8189,N_6451);
and U11581 (N_11581,N_7277,N_7615);
xor U11582 (N_11582,N_7686,N_7642);
and U11583 (N_11583,N_8202,N_7886);
and U11584 (N_11584,N_7934,N_7150);
and U11585 (N_11585,N_6299,N_7701);
or U11586 (N_11586,N_8714,N_7793);
xor U11587 (N_11587,N_6686,N_8603);
nand U11588 (N_11588,N_6523,N_8770);
and U11589 (N_11589,N_7925,N_6472);
or U11590 (N_11590,N_8588,N_7957);
nor U11591 (N_11591,N_8151,N_6872);
or U11592 (N_11592,N_7515,N_6660);
or U11593 (N_11593,N_7799,N_8151);
nand U11594 (N_11594,N_8066,N_8274);
nor U11595 (N_11595,N_6079,N_7364);
nor U11596 (N_11596,N_7095,N_8287);
nand U11597 (N_11597,N_6917,N_6563);
nand U11598 (N_11598,N_6571,N_6950);
nor U11599 (N_11599,N_8224,N_8334);
or U11600 (N_11600,N_8577,N_7113);
nand U11601 (N_11601,N_7029,N_6941);
nor U11602 (N_11602,N_8717,N_6987);
nand U11603 (N_11603,N_7685,N_7852);
or U11604 (N_11604,N_6019,N_6536);
xnor U11605 (N_11605,N_7804,N_6738);
nor U11606 (N_11606,N_8874,N_7693);
nor U11607 (N_11607,N_6735,N_7821);
or U11608 (N_11608,N_7009,N_8498);
and U11609 (N_11609,N_7355,N_7027);
and U11610 (N_11610,N_7094,N_8915);
and U11611 (N_11611,N_7163,N_6585);
nor U11612 (N_11612,N_7477,N_7677);
or U11613 (N_11613,N_8640,N_8528);
nor U11614 (N_11614,N_6348,N_6336);
and U11615 (N_11615,N_6173,N_7295);
and U11616 (N_11616,N_8969,N_6353);
or U11617 (N_11617,N_6977,N_6325);
nand U11618 (N_11618,N_7416,N_6658);
or U11619 (N_11619,N_6717,N_6083);
and U11620 (N_11620,N_6967,N_8475);
nor U11621 (N_11621,N_7936,N_6346);
nor U11622 (N_11622,N_6057,N_7095);
or U11623 (N_11623,N_6415,N_8037);
nand U11624 (N_11624,N_7121,N_7937);
or U11625 (N_11625,N_6570,N_6218);
nand U11626 (N_11626,N_6951,N_8374);
nand U11627 (N_11627,N_7805,N_8605);
or U11628 (N_11628,N_6352,N_8386);
nor U11629 (N_11629,N_8698,N_8950);
nor U11630 (N_11630,N_8750,N_8290);
or U11631 (N_11631,N_6695,N_7890);
and U11632 (N_11632,N_8979,N_8172);
nand U11633 (N_11633,N_8486,N_7226);
nand U11634 (N_11634,N_8043,N_7300);
xor U11635 (N_11635,N_7145,N_8495);
or U11636 (N_11636,N_6539,N_8105);
xor U11637 (N_11637,N_8853,N_8186);
nand U11638 (N_11638,N_6213,N_8653);
nor U11639 (N_11639,N_7790,N_7594);
nand U11640 (N_11640,N_7934,N_6520);
nor U11641 (N_11641,N_8015,N_6301);
and U11642 (N_11642,N_7917,N_6567);
and U11643 (N_11643,N_6810,N_7603);
nor U11644 (N_11644,N_7549,N_6152);
nand U11645 (N_11645,N_7424,N_6163);
and U11646 (N_11646,N_8029,N_6987);
nor U11647 (N_11647,N_6908,N_7329);
or U11648 (N_11648,N_6405,N_7112);
xnor U11649 (N_11649,N_8213,N_6011);
xor U11650 (N_11650,N_7003,N_6716);
and U11651 (N_11651,N_8467,N_7088);
nand U11652 (N_11652,N_7250,N_6667);
nand U11653 (N_11653,N_7228,N_7121);
or U11654 (N_11654,N_7772,N_7317);
or U11655 (N_11655,N_7561,N_6592);
and U11656 (N_11656,N_7851,N_6943);
and U11657 (N_11657,N_7489,N_8053);
and U11658 (N_11658,N_8948,N_8587);
nand U11659 (N_11659,N_6959,N_6661);
and U11660 (N_11660,N_6700,N_7849);
and U11661 (N_11661,N_6381,N_8212);
nand U11662 (N_11662,N_8505,N_7077);
and U11663 (N_11663,N_6610,N_6369);
nand U11664 (N_11664,N_7541,N_7504);
nor U11665 (N_11665,N_7081,N_6580);
and U11666 (N_11666,N_6766,N_6223);
or U11667 (N_11667,N_7112,N_7579);
and U11668 (N_11668,N_6192,N_8877);
nand U11669 (N_11669,N_7927,N_6768);
or U11670 (N_11670,N_6159,N_7044);
nor U11671 (N_11671,N_8807,N_6715);
and U11672 (N_11672,N_8728,N_7860);
xor U11673 (N_11673,N_8790,N_8110);
xnor U11674 (N_11674,N_6521,N_6955);
or U11675 (N_11675,N_6110,N_8358);
nor U11676 (N_11676,N_8882,N_6876);
nor U11677 (N_11677,N_8694,N_6906);
or U11678 (N_11678,N_8625,N_6562);
nor U11679 (N_11679,N_8277,N_6348);
nor U11680 (N_11680,N_6556,N_7007);
or U11681 (N_11681,N_7528,N_6497);
nor U11682 (N_11682,N_8810,N_7597);
or U11683 (N_11683,N_7434,N_7555);
nor U11684 (N_11684,N_6377,N_8067);
and U11685 (N_11685,N_7106,N_6447);
and U11686 (N_11686,N_6478,N_8122);
nand U11687 (N_11687,N_7949,N_8597);
nor U11688 (N_11688,N_8656,N_8970);
and U11689 (N_11689,N_8766,N_8006);
and U11690 (N_11690,N_6195,N_8012);
nor U11691 (N_11691,N_8558,N_8206);
nor U11692 (N_11692,N_7548,N_7405);
nor U11693 (N_11693,N_6830,N_8151);
or U11694 (N_11694,N_8426,N_6138);
nor U11695 (N_11695,N_7325,N_7345);
nor U11696 (N_11696,N_6620,N_6052);
nand U11697 (N_11697,N_8640,N_7514);
nor U11698 (N_11698,N_8399,N_7296);
and U11699 (N_11699,N_7228,N_6769);
xnor U11700 (N_11700,N_6695,N_7554);
or U11701 (N_11701,N_6941,N_6204);
or U11702 (N_11702,N_7231,N_8935);
xor U11703 (N_11703,N_8050,N_8336);
or U11704 (N_11704,N_6416,N_8339);
nand U11705 (N_11705,N_6641,N_6310);
or U11706 (N_11706,N_7594,N_6496);
or U11707 (N_11707,N_7312,N_8948);
nand U11708 (N_11708,N_7395,N_6534);
or U11709 (N_11709,N_6689,N_6114);
or U11710 (N_11710,N_7239,N_8668);
or U11711 (N_11711,N_7423,N_6912);
and U11712 (N_11712,N_7636,N_8954);
and U11713 (N_11713,N_7887,N_7465);
and U11714 (N_11714,N_8953,N_7445);
nor U11715 (N_11715,N_6849,N_7412);
nand U11716 (N_11716,N_6713,N_7605);
and U11717 (N_11717,N_6755,N_8057);
nand U11718 (N_11718,N_8405,N_8816);
nand U11719 (N_11719,N_7603,N_6487);
or U11720 (N_11720,N_8219,N_6856);
xnor U11721 (N_11721,N_7117,N_6176);
nor U11722 (N_11722,N_6977,N_8512);
nor U11723 (N_11723,N_7951,N_8550);
nand U11724 (N_11724,N_6547,N_8284);
and U11725 (N_11725,N_6643,N_7668);
nor U11726 (N_11726,N_6029,N_7748);
xor U11727 (N_11727,N_7980,N_7219);
and U11728 (N_11728,N_6641,N_6590);
and U11729 (N_11729,N_7703,N_6668);
nand U11730 (N_11730,N_6886,N_8322);
and U11731 (N_11731,N_8265,N_7203);
nor U11732 (N_11732,N_7583,N_6862);
or U11733 (N_11733,N_6373,N_6185);
xor U11734 (N_11734,N_6993,N_7345);
nand U11735 (N_11735,N_6230,N_7965);
nand U11736 (N_11736,N_6406,N_7783);
nand U11737 (N_11737,N_6756,N_6446);
or U11738 (N_11738,N_8960,N_8249);
nand U11739 (N_11739,N_7478,N_6256);
or U11740 (N_11740,N_6529,N_6301);
nand U11741 (N_11741,N_6454,N_8576);
or U11742 (N_11742,N_8921,N_7031);
nand U11743 (N_11743,N_7087,N_7615);
and U11744 (N_11744,N_6279,N_7064);
nor U11745 (N_11745,N_8455,N_6188);
or U11746 (N_11746,N_8244,N_7217);
xor U11747 (N_11747,N_6292,N_7434);
nor U11748 (N_11748,N_8123,N_6217);
xor U11749 (N_11749,N_8010,N_6595);
or U11750 (N_11750,N_7552,N_8237);
and U11751 (N_11751,N_6524,N_8628);
or U11752 (N_11752,N_6228,N_8265);
or U11753 (N_11753,N_6525,N_7992);
nor U11754 (N_11754,N_6584,N_8970);
and U11755 (N_11755,N_6285,N_8895);
or U11756 (N_11756,N_6843,N_8437);
nor U11757 (N_11757,N_6147,N_8516);
nand U11758 (N_11758,N_8584,N_8812);
nand U11759 (N_11759,N_6749,N_7798);
and U11760 (N_11760,N_8575,N_8363);
nor U11761 (N_11761,N_8137,N_7622);
nand U11762 (N_11762,N_7526,N_6184);
nand U11763 (N_11763,N_8120,N_7342);
nor U11764 (N_11764,N_8225,N_8236);
nor U11765 (N_11765,N_8042,N_7909);
or U11766 (N_11766,N_6806,N_6756);
nor U11767 (N_11767,N_8048,N_8719);
nor U11768 (N_11768,N_8488,N_8318);
and U11769 (N_11769,N_8537,N_7738);
or U11770 (N_11770,N_7436,N_8081);
nor U11771 (N_11771,N_8454,N_6266);
xor U11772 (N_11772,N_6522,N_8000);
nor U11773 (N_11773,N_8405,N_6717);
nand U11774 (N_11774,N_7853,N_6191);
or U11775 (N_11775,N_6130,N_7845);
nor U11776 (N_11776,N_7017,N_6074);
nand U11777 (N_11777,N_6843,N_8475);
or U11778 (N_11778,N_7139,N_7175);
nand U11779 (N_11779,N_6480,N_7829);
and U11780 (N_11780,N_6729,N_8096);
or U11781 (N_11781,N_8516,N_8074);
nor U11782 (N_11782,N_7898,N_8274);
and U11783 (N_11783,N_6970,N_7774);
xnor U11784 (N_11784,N_6801,N_6571);
or U11785 (N_11785,N_7065,N_6856);
xnor U11786 (N_11786,N_6345,N_6958);
and U11787 (N_11787,N_7439,N_7904);
nor U11788 (N_11788,N_6162,N_8413);
or U11789 (N_11789,N_7499,N_8215);
or U11790 (N_11790,N_8016,N_7786);
or U11791 (N_11791,N_7960,N_8871);
and U11792 (N_11792,N_8222,N_7465);
and U11793 (N_11793,N_7578,N_7320);
xnor U11794 (N_11794,N_6488,N_6939);
or U11795 (N_11795,N_8455,N_6161);
nor U11796 (N_11796,N_8584,N_6969);
and U11797 (N_11797,N_8907,N_7593);
nand U11798 (N_11798,N_8450,N_8790);
nand U11799 (N_11799,N_7776,N_8665);
or U11800 (N_11800,N_8380,N_6391);
nand U11801 (N_11801,N_6906,N_6677);
nand U11802 (N_11802,N_8026,N_7383);
nand U11803 (N_11803,N_7040,N_8983);
or U11804 (N_11804,N_8684,N_7051);
nor U11805 (N_11805,N_8451,N_8180);
xor U11806 (N_11806,N_6097,N_8528);
and U11807 (N_11807,N_6968,N_6455);
nor U11808 (N_11808,N_7471,N_6497);
and U11809 (N_11809,N_6401,N_6064);
or U11810 (N_11810,N_7910,N_7002);
or U11811 (N_11811,N_8500,N_6889);
nand U11812 (N_11812,N_7891,N_6953);
and U11813 (N_11813,N_7387,N_8775);
and U11814 (N_11814,N_8758,N_8137);
or U11815 (N_11815,N_7173,N_7663);
and U11816 (N_11816,N_6527,N_7458);
and U11817 (N_11817,N_8196,N_6878);
nand U11818 (N_11818,N_7501,N_7868);
nor U11819 (N_11819,N_6335,N_6875);
nand U11820 (N_11820,N_6399,N_6620);
nor U11821 (N_11821,N_8540,N_8561);
nor U11822 (N_11822,N_6203,N_7390);
nor U11823 (N_11823,N_8336,N_8610);
nor U11824 (N_11824,N_6046,N_7557);
or U11825 (N_11825,N_6222,N_6296);
and U11826 (N_11826,N_7626,N_8602);
nand U11827 (N_11827,N_8914,N_7934);
or U11828 (N_11828,N_8064,N_8454);
or U11829 (N_11829,N_6228,N_6610);
nand U11830 (N_11830,N_6337,N_8920);
nor U11831 (N_11831,N_6823,N_6278);
nor U11832 (N_11832,N_6951,N_8606);
nand U11833 (N_11833,N_6533,N_6644);
xnor U11834 (N_11834,N_6967,N_6238);
or U11835 (N_11835,N_6412,N_7831);
or U11836 (N_11836,N_6305,N_7056);
and U11837 (N_11837,N_6580,N_7413);
nand U11838 (N_11838,N_8681,N_8049);
nand U11839 (N_11839,N_8876,N_8289);
nand U11840 (N_11840,N_7512,N_6048);
xnor U11841 (N_11841,N_7521,N_6759);
or U11842 (N_11842,N_6813,N_8322);
and U11843 (N_11843,N_6942,N_7413);
and U11844 (N_11844,N_7803,N_7786);
and U11845 (N_11845,N_8503,N_7284);
nor U11846 (N_11846,N_7508,N_7162);
and U11847 (N_11847,N_8112,N_7631);
nand U11848 (N_11848,N_6424,N_6140);
and U11849 (N_11849,N_8923,N_7411);
or U11850 (N_11850,N_8531,N_7037);
nor U11851 (N_11851,N_8834,N_6858);
xnor U11852 (N_11852,N_8826,N_7908);
or U11853 (N_11853,N_8319,N_7137);
nor U11854 (N_11854,N_6413,N_7134);
and U11855 (N_11855,N_6317,N_7868);
or U11856 (N_11856,N_8006,N_8777);
nand U11857 (N_11857,N_8242,N_7676);
and U11858 (N_11858,N_6687,N_8477);
nand U11859 (N_11859,N_8117,N_8951);
nand U11860 (N_11860,N_6361,N_8624);
and U11861 (N_11861,N_6696,N_7168);
nand U11862 (N_11862,N_7274,N_6555);
nand U11863 (N_11863,N_8822,N_7087);
nand U11864 (N_11864,N_7939,N_6368);
nand U11865 (N_11865,N_7116,N_8895);
and U11866 (N_11866,N_7058,N_8640);
and U11867 (N_11867,N_6313,N_6410);
nand U11868 (N_11868,N_7517,N_7918);
nand U11869 (N_11869,N_7822,N_7636);
and U11870 (N_11870,N_7277,N_7816);
or U11871 (N_11871,N_6360,N_8367);
or U11872 (N_11872,N_7168,N_7774);
nor U11873 (N_11873,N_7729,N_7493);
xnor U11874 (N_11874,N_7483,N_6221);
nor U11875 (N_11875,N_7052,N_8541);
and U11876 (N_11876,N_6875,N_6773);
or U11877 (N_11877,N_8159,N_7610);
or U11878 (N_11878,N_7780,N_6034);
nand U11879 (N_11879,N_6153,N_6944);
nand U11880 (N_11880,N_6204,N_8140);
or U11881 (N_11881,N_8948,N_6747);
nand U11882 (N_11882,N_6689,N_7764);
nand U11883 (N_11883,N_6467,N_7866);
xor U11884 (N_11884,N_6838,N_6488);
nand U11885 (N_11885,N_6166,N_8667);
or U11886 (N_11886,N_7541,N_7796);
and U11887 (N_11887,N_7767,N_6397);
or U11888 (N_11888,N_8809,N_7243);
and U11889 (N_11889,N_6448,N_8760);
or U11890 (N_11890,N_6124,N_7307);
or U11891 (N_11891,N_8729,N_8406);
xnor U11892 (N_11892,N_6202,N_8284);
nand U11893 (N_11893,N_7412,N_8058);
nand U11894 (N_11894,N_7422,N_8678);
nor U11895 (N_11895,N_8950,N_6953);
xnor U11896 (N_11896,N_6512,N_6619);
or U11897 (N_11897,N_6689,N_6022);
nand U11898 (N_11898,N_8251,N_7158);
or U11899 (N_11899,N_7098,N_7323);
or U11900 (N_11900,N_7794,N_6987);
nor U11901 (N_11901,N_7739,N_6679);
or U11902 (N_11902,N_7913,N_7569);
or U11903 (N_11903,N_7466,N_8680);
nand U11904 (N_11904,N_8795,N_7551);
xnor U11905 (N_11905,N_7785,N_8855);
nand U11906 (N_11906,N_7483,N_8168);
or U11907 (N_11907,N_8477,N_6880);
nand U11908 (N_11908,N_7098,N_7423);
and U11909 (N_11909,N_7374,N_6064);
nand U11910 (N_11910,N_8466,N_6043);
nand U11911 (N_11911,N_7866,N_7698);
and U11912 (N_11912,N_6303,N_6651);
xnor U11913 (N_11913,N_8517,N_7434);
nand U11914 (N_11914,N_6677,N_8060);
or U11915 (N_11915,N_7907,N_6028);
or U11916 (N_11916,N_8354,N_8238);
nor U11917 (N_11917,N_7794,N_7153);
or U11918 (N_11918,N_7762,N_7114);
nand U11919 (N_11919,N_8359,N_6003);
and U11920 (N_11920,N_6518,N_6695);
xnor U11921 (N_11921,N_7508,N_8865);
or U11922 (N_11922,N_7540,N_6646);
nand U11923 (N_11923,N_8867,N_7208);
nand U11924 (N_11924,N_7389,N_8383);
and U11925 (N_11925,N_8998,N_8537);
or U11926 (N_11926,N_6108,N_8891);
nor U11927 (N_11927,N_7637,N_7929);
nand U11928 (N_11928,N_7068,N_6690);
and U11929 (N_11929,N_8039,N_8088);
nand U11930 (N_11930,N_8633,N_6568);
xor U11931 (N_11931,N_6696,N_7341);
nand U11932 (N_11932,N_8582,N_7475);
and U11933 (N_11933,N_7870,N_6382);
nand U11934 (N_11934,N_8998,N_8887);
nor U11935 (N_11935,N_7220,N_8176);
or U11936 (N_11936,N_7145,N_8867);
or U11937 (N_11937,N_7986,N_6747);
nor U11938 (N_11938,N_6357,N_7497);
or U11939 (N_11939,N_6016,N_8502);
xnor U11940 (N_11940,N_6413,N_7858);
or U11941 (N_11941,N_6216,N_6572);
or U11942 (N_11942,N_6752,N_8161);
nand U11943 (N_11943,N_6133,N_6293);
and U11944 (N_11944,N_8533,N_6779);
nand U11945 (N_11945,N_6444,N_8681);
nor U11946 (N_11946,N_8515,N_6388);
nand U11947 (N_11947,N_6503,N_6706);
and U11948 (N_11948,N_7108,N_8699);
and U11949 (N_11949,N_8224,N_7941);
and U11950 (N_11950,N_8949,N_6739);
or U11951 (N_11951,N_6899,N_6756);
nor U11952 (N_11952,N_7951,N_8161);
and U11953 (N_11953,N_6472,N_6682);
xor U11954 (N_11954,N_6792,N_7738);
nand U11955 (N_11955,N_8933,N_6162);
nor U11956 (N_11956,N_8475,N_6396);
nand U11957 (N_11957,N_7491,N_7067);
nand U11958 (N_11958,N_8214,N_6887);
xnor U11959 (N_11959,N_6100,N_6708);
nor U11960 (N_11960,N_6998,N_7908);
or U11961 (N_11961,N_7330,N_6985);
and U11962 (N_11962,N_6150,N_8158);
xor U11963 (N_11963,N_7025,N_7634);
nor U11964 (N_11964,N_6805,N_7129);
nor U11965 (N_11965,N_8020,N_6369);
or U11966 (N_11966,N_8813,N_8038);
nand U11967 (N_11967,N_6521,N_8200);
nand U11968 (N_11968,N_8575,N_7577);
or U11969 (N_11969,N_6123,N_7991);
nand U11970 (N_11970,N_6439,N_6865);
nor U11971 (N_11971,N_8374,N_6928);
nor U11972 (N_11972,N_6012,N_6837);
and U11973 (N_11973,N_8428,N_6791);
nor U11974 (N_11974,N_8350,N_8279);
and U11975 (N_11975,N_7237,N_8371);
nand U11976 (N_11976,N_8491,N_7776);
nor U11977 (N_11977,N_7600,N_6973);
and U11978 (N_11978,N_7517,N_6672);
nor U11979 (N_11979,N_8796,N_7882);
nor U11980 (N_11980,N_6773,N_8235);
nand U11981 (N_11981,N_8934,N_7033);
and U11982 (N_11982,N_8913,N_6857);
nor U11983 (N_11983,N_8584,N_6928);
nand U11984 (N_11984,N_6925,N_7352);
or U11985 (N_11985,N_7165,N_6442);
nand U11986 (N_11986,N_6905,N_6222);
nand U11987 (N_11987,N_6301,N_8392);
or U11988 (N_11988,N_8371,N_6235);
or U11989 (N_11989,N_7307,N_8476);
or U11990 (N_11990,N_6134,N_8844);
or U11991 (N_11991,N_7021,N_6196);
nand U11992 (N_11992,N_6725,N_6115);
nor U11993 (N_11993,N_8885,N_8579);
and U11994 (N_11994,N_8585,N_8365);
nand U11995 (N_11995,N_8433,N_8941);
or U11996 (N_11996,N_8501,N_8332);
or U11997 (N_11997,N_8560,N_6073);
nor U11998 (N_11998,N_8662,N_6456);
or U11999 (N_11999,N_7243,N_6739);
nor U12000 (N_12000,N_9038,N_11750);
and U12001 (N_12001,N_10028,N_9464);
nand U12002 (N_12002,N_9388,N_11287);
nand U12003 (N_12003,N_9888,N_9330);
nor U12004 (N_12004,N_11334,N_11613);
or U12005 (N_12005,N_11438,N_9911);
xnor U12006 (N_12006,N_11770,N_11077);
or U12007 (N_12007,N_11366,N_9612);
nand U12008 (N_12008,N_10820,N_9735);
nand U12009 (N_12009,N_9240,N_10739);
and U12010 (N_12010,N_11248,N_10760);
nand U12011 (N_12011,N_10159,N_9710);
nand U12012 (N_12012,N_9596,N_9780);
and U12013 (N_12013,N_9857,N_9946);
nor U12014 (N_12014,N_10615,N_10668);
and U12015 (N_12015,N_10179,N_11514);
and U12016 (N_12016,N_10768,N_10323);
or U12017 (N_12017,N_11680,N_10343);
nor U12018 (N_12018,N_9491,N_9499);
or U12019 (N_12019,N_9969,N_10680);
nand U12020 (N_12020,N_9262,N_10614);
and U12021 (N_12021,N_9691,N_11369);
and U12022 (N_12022,N_10688,N_11411);
nand U12023 (N_12023,N_11407,N_9152);
and U12024 (N_12024,N_9487,N_11188);
nor U12025 (N_12025,N_9065,N_11832);
nand U12026 (N_12026,N_11747,N_10581);
or U12027 (N_12027,N_9413,N_9938);
or U12028 (N_12028,N_9971,N_11524);
nand U12029 (N_12029,N_9353,N_9091);
nor U12030 (N_12030,N_9422,N_9712);
nand U12031 (N_12031,N_9173,N_9520);
nand U12032 (N_12032,N_10977,N_9279);
and U12033 (N_12033,N_11452,N_10289);
nand U12034 (N_12034,N_10004,N_11622);
nor U12035 (N_12035,N_10194,N_9602);
and U12036 (N_12036,N_11529,N_10859);
or U12037 (N_12037,N_10936,N_10453);
nor U12038 (N_12038,N_10539,N_11170);
nand U12039 (N_12039,N_11310,N_9160);
or U12040 (N_12040,N_10899,N_11738);
or U12041 (N_12041,N_10772,N_11006);
nor U12042 (N_12042,N_10745,N_11149);
or U12043 (N_12043,N_11111,N_9868);
and U12044 (N_12044,N_11639,N_9940);
or U12045 (N_12045,N_9733,N_10832);
and U12046 (N_12046,N_9168,N_10372);
xor U12047 (N_12047,N_10093,N_10074);
and U12048 (N_12048,N_11079,N_11228);
or U12049 (N_12049,N_11752,N_10065);
xnor U12050 (N_12050,N_11207,N_9711);
and U12051 (N_12051,N_9545,N_10340);
and U12052 (N_12052,N_10559,N_10332);
or U12053 (N_12053,N_11164,N_11692);
nand U12054 (N_12054,N_9478,N_9116);
nor U12055 (N_12055,N_9725,N_9890);
and U12056 (N_12056,N_11425,N_11018);
nand U12057 (N_12057,N_10360,N_10046);
nand U12058 (N_12058,N_10992,N_11532);
nor U12059 (N_12059,N_11621,N_9473);
nand U12060 (N_12060,N_9433,N_9933);
nor U12061 (N_12061,N_9690,N_10122);
nor U12062 (N_12062,N_9925,N_9158);
nand U12063 (N_12063,N_10035,N_10007);
nor U12064 (N_12064,N_9517,N_11444);
nand U12065 (N_12065,N_9072,N_10097);
nand U12066 (N_12066,N_11651,N_10967);
xnor U12067 (N_12067,N_9761,N_9221);
nor U12068 (N_12068,N_11501,N_10994);
nand U12069 (N_12069,N_11855,N_10841);
nand U12070 (N_12070,N_11705,N_11120);
and U12071 (N_12071,N_11488,N_11543);
xnor U12072 (N_12072,N_11424,N_10100);
nand U12073 (N_12073,N_9273,N_9189);
and U12074 (N_12074,N_11729,N_11667);
nor U12075 (N_12075,N_10068,N_10962);
and U12076 (N_12076,N_11908,N_10753);
or U12077 (N_12077,N_9106,N_11263);
nand U12078 (N_12078,N_11986,N_9174);
nor U12079 (N_12079,N_11762,N_10823);
and U12080 (N_12080,N_11527,N_9426);
nor U12081 (N_12081,N_9034,N_10444);
or U12082 (N_12082,N_11503,N_10445);
or U12083 (N_12083,N_9894,N_9172);
and U12084 (N_12084,N_10677,N_11582);
nand U12085 (N_12085,N_10866,N_10766);
nand U12086 (N_12086,N_10432,N_11174);
and U12087 (N_12087,N_9226,N_9744);
or U12088 (N_12088,N_9453,N_10512);
or U12089 (N_12089,N_10812,N_11493);
nor U12090 (N_12090,N_9755,N_9959);
nor U12091 (N_12091,N_9944,N_11222);
nor U12092 (N_12092,N_9856,N_10954);
or U12093 (N_12093,N_10346,N_9895);
or U12094 (N_12094,N_11601,N_11952);
or U12095 (N_12095,N_10361,N_9247);
nand U12096 (N_12096,N_9220,N_11447);
nand U12097 (N_12097,N_11713,N_9313);
nor U12098 (N_12098,N_9929,N_11481);
nand U12099 (N_12099,N_10722,N_11051);
xnor U12100 (N_12100,N_11735,N_10293);
nor U12101 (N_12101,N_11870,N_9992);
nand U12102 (N_12102,N_10968,N_10758);
nor U12103 (N_12103,N_11110,N_10807);
nand U12104 (N_12104,N_9885,N_11707);
nand U12105 (N_12105,N_11135,N_10240);
nor U12106 (N_12106,N_9452,N_10817);
and U12107 (N_12107,N_11001,N_11560);
xnor U12108 (N_12108,N_11666,N_11749);
and U12109 (N_12109,N_10996,N_11740);
and U12110 (N_12110,N_11399,N_11595);
and U12111 (N_12111,N_10025,N_11344);
nor U12112 (N_12112,N_10462,N_11193);
and U12113 (N_12113,N_9742,N_9652);
and U12114 (N_12114,N_9335,N_10834);
nor U12115 (N_12115,N_9627,N_11904);
and U12116 (N_12116,N_9937,N_9649);
and U12117 (N_12117,N_11247,N_11437);
nand U12118 (N_12118,N_10472,N_9859);
or U12119 (N_12119,N_9418,N_11609);
and U12120 (N_12120,N_10139,N_11069);
nor U12121 (N_12121,N_9178,N_11883);
nor U12122 (N_12122,N_10281,N_10514);
xnor U12123 (N_12123,N_10811,N_9212);
and U12124 (N_12124,N_10258,N_10019);
nand U12125 (N_12125,N_9367,N_10185);
nor U12126 (N_12126,N_10051,N_9547);
or U12127 (N_12127,N_10984,N_11333);
or U12128 (N_12128,N_9037,N_10575);
nor U12129 (N_12129,N_9722,N_11664);
or U12130 (N_12130,N_9993,N_11377);
and U12131 (N_12131,N_9290,N_11092);
nor U12132 (N_12132,N_9949,N_11649);
or U12133 (N_12133,N_9784,N_11823);
and U12134 (N_12134,N_9689,N_9489);
and U12135 (N_12135,N_10684,N_11098);
nor U12136 (N_12136,N_10489,N_9512);
nand U12137 (N_12137,N_10925,N_10211);
and U12138 (N_12138,N_9497,N_10558);
or U12139 (N_12139,N_10848,N_11237);
nor U12140 (N_12140,N_11874,N_11365);
nor U12141 (N_12141,N_11227,N_11242);
and U12142 (N_12142,N_11795,N_11321);
xnor U12143 (N_12143,N_9082,N_10325);
or U12144 (N_12144,N_9077,N_10145);
nor U12145 (N_12145,N_10588,N_11725);
and U12146 (N_12146,N_10241,N_10061);
and U12147 (N_12147,N_10413,N_9345);
nor U12148 (N_12148,N_9154,N_9011);
nor U12149 (N_12149,N_11066,N_11246);
nor U12150 (N_12150,N_11922,N_9886);
and U12151 (N_12151,N_9781,N_10013);
and U12152 (N_12152,N_11654,N_10526);
nor U12153 (N_12153,N_9257,N_10502);
and U12154 (N_12154,N_11026,N_9736);
xnor U12155 (N_12155,N_11233,N_11721);
or U12156 (N_12156,N_10550,N_9383);
and U12157 (N_12157,N_10981,N_10594);
nor U12158 (N_12158,N_10278,N_11893);
or U12159 (N_12159,N_9393,N_9145);
nor U12160 (N_12160,N_9439,N_10170);
nor U12161 (N_12161,N_9964,N_10762);
nor U12162 (N_12162,N_10063,N_11270);
nand U12163 (N_12163,N_11802,N_9915);
xor U12164 (N_12164,N_10543,N_10390);
nand U12165 (N_12165,N_9347,N_10902);
or U12166 (N_12166,N_10112,N_9440);
nand U12167 (N_12167,N_11157,N_11388);
nand U12168 (N_12168,N_10460,N_9398);
nand U12169 (N_12169,N_11583,N_11943);
nor U12170 (N_12170,N_9568,N_11045);
or U12171 (N_12171,N_10197,N_10826);
nor U12172 (N_12172,N_10394,N_11957);
nor U12173 (N_12173,N_9519,N_9527);
and U12174 (N_12174,N_10080,N_11013);
or U12175 (N_12175,N_10257,N_10307);
or U12176 (N_12176,N_10113,N_10914);
and U12177 (N_12177,N_10754,N_9905);
nand U12178 (N_12178,N_9558,N_10591);
or U12179 (N_12179,N_9076,N_11876);
nor U12180 (N_12180,N_9292,N_10710);
nor U12181 (N_12181,N_10192,N_11303);
nor U12182 (N_12182,N_11137,N_9099);
xor U12183 (N_12183,N_10647,N_9598);
nor U12184 (N_12184,N_10029,N_9556);
nand U12185 (N_12185,N_9343,N_10733);
or U12186 (N_12186,N_9067,N_11350);
or U12187 (N_12187,N_9705,N_9331);
nand U12188 (N_12188,N_9447,N_10057);
xnor U12189 (N_12189,N_11511,N_9640);
and U12190 (N_12190,N_11196,N_11746);
nor U12191 (N_12191,N_11240,N_10259);
and U12192 (N_12192,N_10813,N_11857);
xnor U12193 (N_12193,N_11487,N_10619);
nor U12194 (N_12194,N_10107,N_9291);
or U12195 (N_12195,N_11868,N_9889);
and U12196 (N_12196,N_11919,N_11146);
and U12197 (N_12197,N_9004,N_9211);
nand U12198 (N_12198,N_11895,N_10334);
or U12199 (N_12199,N_9363,N_10264);
and U12200 (N_12200,N_9719,N_9955);
nand U12201 (N_12201,N_9751,N_9770);
nor U12202 (N_12202,N_10862,N_11837);
nand U12203 (N_12203,N_11504,N_11357);
or U12204 (N_12204,N_9282,N_11508);
nand U12205 (N_12205,N_11800,N_9000);
and U12206 (N_12206,N_10429,N_10956);
nor U12207 (N_12207,N_9739,N_9919);
and U12208 (N_12208,N_11484,N_11281);
xor U12209 (N_12209,N_10528,N_10697);
nand U12210 (N_12210,N_10313,N_10180);
nand U12211 (N_12211,N_11078,N_11476);
and U12212 (N_12212,N_11858,N_10015);
and U12213 (N_12213,N_10036,N_10000);
xor U12214 (N_12214,N_10484,N_11323);
and U12215 (N_12215,N_9295,N_10976);
nand U12216 (N_12216,N_10838,N_11463);
nor U12217 (N_12217,N_9248,N_11523);
and U12218 (N_12218,N_10297,N_9385);
nand U12219 (N_12219,N_9490,N_10879);
or U12220 (N_12220,N_11700,N_9031);
or U12221 (N_12221,N_11685,N_11814);
nor U12222 (N_12222,N_10085,N_10948);
nor U12223 (N_12223,N_9968,N_9853);
or U12224 (N_12224,N_11615,N_11141);
nor U12225 (N_12225,N_9534,N_11326);
xor U12226 (N_12226,N_9530,N_11933);
or U12227 (N_12227,N_11611,N_10212);
xor U12228 (N_12228,N_9669,N_9941);
nand U12229 (N_12229,N_11181,N_11902);
or U12230 (N_12230,N_9263,N_9327);
nand U12231 (N_12231,N_11683,N_9100);
and U12232 (N_12232,N_11154,N_9636);
or U12233 (N_12233,N_11122,N_10157);
and U12234 (N_12234,N_9797,N_9175);
nor U12235 (N_12235,N_9578,N_10843);
and U12236 (N_12236,N_10928,N_9769);
or U12237 (N_12237,N_9697,N_10705);
and U12238 (N_12238,N_9169,N_11914);
nand U12239 (N_12239,N_10142,N_9504);
or U12240 (N_12240,N_9429,N_11024);
and U12241 (N_12241,N_11776,N_9581);
and U12242 (N_12242,N_10597,N_9550);
nand U12243 (N_12243,N_11982,N_10224);
nand U12244 (N_12244,N_9161,N_10917);
or U12245 (N_12245,N_11696,N_9006);
nor U12246 (N_12246,N_9579,N_11367);
nor U12247 (N_12247,N_11002,N_11040);
nand U12248 (N_12248,N_11567,N_9924);
and U12249 (N_12249,N_11056,N_11273);
nand U12250 (N_12250,N_10506,N_10407);
nor U12251 (N_12251,N_11833,N_10676);
and U12252 (N_12252,N_11179,N_11029);
nand U12253 (N_12253,N_10802,N_9671);
or U12254 (N_12254,N_9724,N_10808);
nor U12255 (N_12255,N_11606,N_10441);
nand U12256 (N_12256,N_11182,N_11549);
nor U12257 (N_12257,N_11408,N_11360);
and U12258 (N_12258,N_11891,N_10347);
nand U12259 (N_12259,N_11245,N_10064);
and U12260 (N_12260,N_10828,N_10136);
nand U12261 (N_12261,N_10108,N_10806);
or U12262 (N_12262,N_9566,N_11964);
nor U12263 (N_12263,N_9427,N_9832);
nand U12264 (N_12264,N_9210,N_10524);
nor U12265 (N_12265,N_9577,N_9023);
nand U12266 (N_12266,N_10238,N_11668);
nand U12267 (N_12267,N_10103,N_10671);
nor U12268 (N_12268,N_10290,N_10189);
and U12269 (N_12269,N_10009,N_10577);
nand U12270 (N_12270,N_10475,N_10260);
or U12271 (N_12271,N_11550,N_9228);
and U12272 (N_12272,N_9546,N_10243);
nand U12273 (N_12273,N_9514,N_10294);
nand U12274 (N_12274,N_10188,N_9907);
and U12275 (N_12275,N_9713,N_10470);
nor U12276 (N_12276,N_11505,N_10451);
xor U12277 (N_12277,N_11482,N_11307);
or U12278 (N_12278,N_11566,N_9663);
nand U12279 (N_12279,N_9498,N_10392);
or U12280 (N_12280,N_11635,N_9417);
or U12281 (N_12281,N_9644,N_10711);
or U12282 (N_12282,N_11663,N_10805);
or U12283 (N_12283,N_9167,N_9686);
or U12284 (N_12284,N_9776,N_9960);
xor U12285 (N_12285,N_11112,N_11072);
or U12286 (N_12286,N_9488,N_9648);
and U12287 (N_12287,N_11852,N_10836);
nand U12288 (N_12288,N_11008,N_11925);
or U12289 (N_12289,N_9752,N_10349);
or U12290 (N_12290,N_10079,N_9125);
xnor U12291 (N_12291,N_11854,N_9983);
nand U12292 (N_12292,N_10961,N_9320);
nor U12293 (N_12293,N_9536,N_10352);
nor U12294 (N_12294,N_10164,N_9328);
or U12295 (N_12295,N_10153,N_10427);
xor U12296 (N_12296,N_9087,N_10098);
nand U12297 (N_12297,N_10835,N_11093);
or U12298 (N_12298,N_9457,N_10355);
and U12299 (N_12299,N_11882,N_9216);
nor U12300 (N_12300,N_9013,N_10253);
or U12301 (N_12301,N_10439,N_10777);
nor U12302 (N_12302,N_11023,N_9419);
nor U12303 (N_12303,N_11299,N_11525);
nand U12304 (N_12304,N_10696,N_9700);
xnor U12305 (N_12305,N_10495,N_9537);
nand U12306 (N_12306,N_9316,N_9951);
xor U12307 (N_12307,N_10544,N_11600);
and U12308 (N_12308,N_11265,N_10242);
nand U12309 (N_12309,N_11250,N_10646);
and U12310 (N_12310,N_9591,N_9775);
and U12311 (N_12311,N_11301,N_9092);
and U12312 (N_12312,N_10350,N_11702);
nor U12313 (N_12313,N_11329,N_10568);
and U12314 (N_12314,N_9289,N_9802);
xnor U12315 (N_12315,N_11348,N_9467);
nand U12316 (N_12316,N_11537,N_9777);
xor U12317 (N_12317,N_11378,N_11198);
nor U12318 (N_12318,N_9768,N_10296);
or U12319 (N_12319,N_9151,N_9675);
xnor U12320 (N_12320,N_10341,N_9851);
or U12321 (N_12321,N_11605,N_10927);
nand U12322 (N_12322,N_11086,N_9513);
and U12323 (N_12323,N_10989,N_11998);
or U12324 (N_12324,N_10338,N_10723);
or U12325 (N_12325,N_9618,N_10482);
nor U12326 (N_12326,N_11830,N_10020);
xor U12327 (N_12327,N_9286,N_11594);
xnor U12328 (N_12328,N_9718,N_10207);
nand U12329 (N_12329,N_10148,N_11589);
nand U12330 (N_12330,N_9050,N_10778);
nand U12331 (N_12331,N_10055,N_11224);
nand U12332 (N_12332,N_10381,N_11522);
or U12333 (N_12333,N_9796,N_10269);
or U12334 (N_12334,N_11880,N_9985);
xor U12335 (N_12335,N_9156,N_10230);
nand U12336 (N_12336,N_9254,N_11404);
and U12337 (N_12337,N_11827,N_11864);
and U12338 (N_12338,N_9338,N_11088);
or U12339 (N_12339,N_11291,N_11331);
nand U12340 (N_12340,N_10542,N_9430);
nor U12341 (N_12341,N_11644,N_10727);
nor U12342 (N_12342,N_10500,N_11570);
or U12343 (N_12343,N_11542,N_11708);
xnor U12344 (N_12344,N_10239,N_10328);
nand U12345 (N_12345,N_10895,N_11819);
nand U12346 (N_12346,N_10314,N_11067);
and U12347 (N_12347,N_10573,N_9656);
or U12348 (N_12348,N_9217,N_11808);
nand U12349 (N_12349,N_11148,N_11913);
and U12350 (N_12350,N_9283,N_10104);
nor U12351 (N_12351,N_11140,N_11244);
or U12352 (N_12352,N_9348,N_9203);
nand U12353 (N_12353,N_9355,N_11199);
nand U12354 (N_12354,N_11121,N_11965);
xor U12355 (N_12355,N_10102,N_9144);
xnor U12356 (N_12356,N_11255,N_9854);
or U12357 (N_12357,N_11486,N_9296);
nand U12358 (N_12358,N_9528,N_10904);
or U12359 (N_12359,N_10686,N_9202);
and U12360 (N_12360,N_9105,N_10958);
nor U12361 (N_12361,N_11389,N_11608);
or U12362 (N_12362,N_9773,N_10531);
and U12363 (N_12363,N_11896,N_9239);
nand U12364 (N_12364,N_11576,N_11052);
nor U12365 (N_12365,N_10105,N_9753);
or U12366 (N_12366,N_9045,N_9039);
or U12367 (N_12367,N_9952,N_9935);
nand U12368 (N_12368,N_10272,N_11544);
nor U12369 (N_12369,N_11172,N_11446);
nor U12370 (N_12370,N_9576,N_9408);
nor U12371 (N_12371,N_11743,N_10375);
or U12372 (N_12372,N_11266,N_10030);
and U12373 (N_12373,N_11975,N_11726);
nor U12374 (N_12374,N_9500,N_11068);
nor U12375 (N_12375,N_10865,N_9056);
nand U12376 (N_12376,N_9410,N_10703);
nand U12377 (N_12377,N_9101,N_9871);
nor U12378 (N_12378,N_9390,N_11478);
and U12379 (N_12379,N_11551,N_9459);
nand U12380 (N_12380,N_11821,N_11144);
and U12381 (N_12381,N_10149,N_10440);
nor U12382 (N_12382,N_9564,N_10202);
or U12383 (N_12383,N_9632,N_11230);
nor U12384 (N_12384,N_9645,N_11390);
or U12385 (N_12385,N_10492,N_11796);
or U12386 (N_12386,N_11361,N_11206);
nor U12387 (N_12387,N_10856,N_10532);
or U12388 (N_12388,N_10467,N_9639);
and U12389 (N_12389,N_10576,N_9628);
or U12390 (N_12390,N_11978,N_10126);
nand U12391 (N_12391,N_11995,N_11967);
and U12392 (N_12392,N_9928,N_9437);
nor U12393 (N_12393,N_11443,N_9963);
nor U12394 (N_12394,N_10868,N_10523);
nor U12395 (N_12395,N_10561,N_9068);
xnor U12396 (N_12396,N_9807,N_10673);
nand U12397 (N_12397,N_9694,N_9232);
or U12398 (N_12398,N_10761,N_9759);
nor U12399 (N_12399,N_11989,N_9269);
and U12400 (N_12400,N_11588,N_11612);
nand U12401 (N_12401,N_11211,N_11084);
and U12402 (N_12402,N_9372,N_10210);
nor U12403 (N_12403,N_11125,N_11316);
and U12404 (N_12404,N_10311,N_9192);
and U12405 (N_12405,N_11983,N_10624);
nor U12406 (N_12406,N_11778,N_9760);
nand U12407 (N_12407,N_11736,N_10410);
nand U12408 (N_12408,N_10771,N_11229);
or U12409 (N_12409,N_11962,N_9730);
nand U12410 (N_12410,N_11768,N_10549);
nor U12411 (N_12411,N_10208,N_9134);
nand U12412 (N_12412,N_9842,N_9732);
or U12413 (N_12413,N_10553,N_11494);
nand U12414 (N_12414,N_10535,N_9839);
and U12415 (N_12415,N_11565,N_11974);
nand U12416 (N_12416,N_11368,N_9253);
or U12417 (N_12417,N_9574,N_10872);
or U12418 (N_12418,N_11131,N_10363);
or U12419 (N_12419,N_9020,N_9800);
or U12420 (N_12420,N_9609,N_11687);
xor U12421 (N_12421,N_9825,N_11364);
and U12422 (N_12422,N_9325,N_9779);
nor U12423 (N_12423,N_10950,N_11436);
or U12424 (N_12424,N_11540,N_11031);
and U12425 (N_12425,N_10096,N_11657);
nand U12426 (N_12426,N_11577,N_10088);
and U12427 (N_12427,N_11617,N_11728);
xnor U12428 (N_12428,N_10508,N_10234);
nor U12429 (N_12429,N_9967,N_10273);
and U12430 (N_12430,N_10274,N_10123);
or U12431 (N_12431,N_11183,N_9406);
nor U12432 (N_12432,N_11243,N_9672);
or U12433 (N_12433,N_11380,N_9643);
and U12434 (N_12434,N_9236,N_11760);
and U12435 (N_12435,N_11221,N_10885);
nand U12436 (N_12436,N_9979,N_9861);
nor U12437 (N_12437,N_11103,N_11528);
or U12438 (N_12438,N_10815,N_10628);
and U12439 (N_12439,N_11899,N_10504);
or U12440 (N_12440,N_11383,N_11238);
xnor U12441 (N_12441,N_11409,N_10538);
nand U12442 (N_12442,N_11994,N_11704);
xnor U12443 (N_12443,N_11355,N_11319);
xor U12444 (N_12444,N_11302,N_11960);
and U12445 (N_12445,N_9521,N_11309);
and U12446 (N_12446,N_11012,N_11027);
or U12447 (N_12447,N_10518,N_11737);
nand U12448 (N_12448,N_10437,N_11706);
nor U12449 (N_12449,N_11405,N_10486);
nand U12450 (N_12450,N_10665,N_9703);
nor U12451 (N_12451,N_9136,N_9709);
nor U12452 (N_12452,N_10450,N_11679);
or U12453 (N_12453,N_10071,N_11673);
and U12454 (N_12454,N_11690,N_11733);
or U12455 (N_12455,N_9749,N_10683);
or U12456 (N_12456,N_10829,N_11940);
or U12457 (N_12457,N_10995,N_9040);
nand U12458 (N_12458,N_11279,N_11280);
nand U12459 (N_12459,N_9191,N_9024);
nand U12460 (N_12460,N_10040,N_11173);
nand U12461 (N_12461,N_11603,N_9061);
and U12462 (N_12462,N_10428,N_11371);
and U12463 (N_12463,N_11175,N_9745);
xor U12464 (N_12464,N_9285,N_9896);
nand U12465 (N_12465,N_9199,N_9271);
nor U12466 (N_12466,N_10990,N_11153);
or U12467 (N_12467,N_11000,N_11759);
nor U12468 (N_12468,N_9492,N_10268);
nand U12469 (N_12469,N_10901,N_11987);
and U12470 (N_12470,N_9147,N_10319);
and U12471 (N_12471,N_9297,N_10803);
or U12472 (N_12472,N_11132,N_10897);
and U12473 (N_12473,N_10578,N_9009);
nand U12474 (N_12474,N_11490,N_10465);
and U12475 (N_12475,N_10005,N_10010);
or U12476 (N_12476,N_10801,N_9984);
nand U12477 (N_12477,N_11777,N_9977);
nor U12478 (N_12478,N_9458,N_9276);
or U12479 (N_12479,N_11877,N_9835);
nand U12480 (N_12480,N_10540,N_9042);
nand U12481 (N_12481,N_10499,N_11531);
nand U12482 (N_12482,N_9140,N_10271);
or U12483 (N_12483,N_10449,N_11455);
xor U12484 (N_12484,N_11694,N_11275);
nor U12485 (N_12485,N_11458,N_11354);
nor U12486 (N_12486,N_9589,N_9235);
nand U12487 (N_12487,N_10567,N_9523);
nor U12488 (N_12488,N_10534,N_9046);
nor U12489 (N_12489,N_11046,N_11948);
or U12490 (N_12490,N_10322,N_11961);
nor U12491 (N_12491,N_9683,N_10382);
or U12492 (N_12492,N_10026,N_10396);
nor U12493 (N_12493,N_9463,N_10800);
nor U12494 (N_12494,N_10659,N_9256);
nand U12495 (N_12495,N_9509,N_10704);
and U12496 (N_12496,N_9462,N_9176);
and U12497 (N_12497,N_11470,N_11672);
and U12498 (N_12498,N_10154,N_9364);
xor U12499 (N_12499,N_9163,N_10072);
and U12500 (N_12500,N_10639,N_11048);
and U12501 (N_12501,N_9631,N_10699);
nand U12502 (N_12502,N_10474,N_11906);
and U12503 (N_12503,N_9567,N_11597);
nor U12504 (N_12504,N_10191,N_11586);
or U12505 (N_12505,N_11379,N_9129);
or U12506 (N_12506,N_10417,N_10886);
and U12507 (N_12507,N_9403,N_10251);
or U12508 (N_12508,N_11100,N_11968);
nor U12509 (N_12509,N_11025,N_11641);
nor U12510 (N_12510,N_9670,N_11351);
or U12511 (N_12511,N_10235,N_11075);
nor U12512 (N_12512,N_9261,N_10226);
or U12513 (N_12513,N_10089,N_9195);
and U12514 (N_12514,N_9139,N_9058);
nand U12515 (N_12515,N_11442,N_9180);
and U12516 (N_12516,N_9950,N_11731);
nor U12517 (N_12517,N_9241,N_10110);
and U12518 (N_12518,N_11346,N_11292);
and U12519 (N_12519,N_10487,N_9019);
nor U12520 (N_12520,N_10882,N_9966);
nor U12521 (N_12521,N_11097,N_9337);
nand U12522 (N_12522,N_9373,N_11382);
and U12523 (N_12523,N_10972,N_11714);
nor U12524 (N_12524,N_9196,N_10522);
xnor U12525 (N_12525,N_10944,N_9706);
and U12526 (N_12526,N_9224,N_9765);
nand U12527 (N_12527,N_10245,N_10468);
and U12528 (N_12528,N_11363,N_9660);
nor U12529 (N_12529,N_11058,N_11912);
or U12530 (N_12530,N_11826,N_11136);
or U12531 (N_12531,N_10873,N_10718);
nor U12532 (N_12532,N_9572,N_9471);
nand U12533 (N_12533,N_10127,N_10564);
or U12534 (N_12534,N_10779,N_10075);
and U12535 (N_12535,N_11467,N_9095);
nor U12536 (N_12536,N_10461,N_11782);
xor U12537 (N_12537,N_10318,N_9131);
nand U12538 (N_12538,N_10616,N_11630);
or U12539 (N_12539,N_9953,N_11185);
or U12540 (N_12540,N_10818,N_9544);
nor U12541 (N_12541,N_11927,N_10266);
nand U12542 (N_12542,N_9494,N_9936);
or U12543 (N_12543,N_10695,N_9621);
or U12544 (N_12544,N_9947,N_9507);
nand U12545 (N_12545,N_10099,N_9493);
and U12546 (N_12546,N_11096,N_10510);
nand U12547 (N_12547,N_9810,N_10478);
nor U12548 (N_12548,N_9468,N_11681);
or U12549 (N_12549,N_10602,N_9877);
and U12550 (N_12550,N_10181,N_10713);
xnor U12551 (N_12551,N_9515,N_10633);
or U12552 (N_12552,N_10367,N_11335);
or U12553 (N_12553,N_11691,N_9586);
and U12554 (N_12554,N_9182,N_10431);
and U12555 (N_12555,N_11637,N_11277);
or U12556 (N_12556,N_11203,N_11171);
and U12557 (N_12557,N_9608,N_9665);
xor U12558 (N_12558,N_10657,N_9094);
nand U12559 (N_12559,N_9083,N_11332);
or U12560 (N_12560,N_9412,N_9214);
and U12561 (N_12561,N_11076,N_10734);
nand U12562 (N_12562,N_9786,N_10199);
nand U12563 (N_12563,N_11129,N_9573);
nor U12564 (N_12564,N_11593,N_10301);
or U12565 (N_12565,N_9307,N_9611);
nor U12566 (N_12566,N_11118,N_10609);
or U12567 (N_12567,N_10764,N_9738);
nor U12568 (N_12568,N_9599,N_10911);
nor U12569 (N_12569,N_9450,N_9481);
or U12570 (N_12570,N_11534,N_10132);
and U12571 (N_12571,N_10423,N_9392);
or U12572 (N_12572,N_9592,N_10128);
nand U12573 (N_12573,N_10923,N_11061);
and U12574 (N_12574,N_11753,N_10755);
nand U12575 (N_12575,N_11480,N_10023);
or U12576 (N_12576,N_9043,N_11370);
and U12577 (N_12577,N_10728,N_11686);
or U12578 (N_12578,N_11944,N_11842);
nor U12579 (N_12579,N_10214,N_11267);
xnor U12580 (N_12580,N_11123,N_10912);
or U12581 (N_12581,N_9107,N_11195);
and U12582 (N_12582,N_11191,N_10285);
and U12583 (N_12583,N_9183,N_11820);
or U12584 (N_12584,N_10587,N_11539);
and U12585 (N_12585,N_11201,N_9208);
or U12586 (N_12586,N_9616,N_9870);
and U12587 (N_12587,N_10321,N_10658);
nor U12588 (N_12588,N_10858,N_9909);
nand U12589 (N_12589,N_11572,N_10270);
and U12590 (N_12590,N_10837,N_11089);
or U12591 (N_12591,N_10436,N_9052);
or U12592 (N_12592,N_10625,N_11127);
and U12593 (N_12593,N_9876,N_11579);
and U12594 (N_12594,N_11495,N_11688);
xor U12595 (N_12595,N_9090,N_9329);
or U12596 (N_12596,N_10151,N_10130);
and U12597 (N_12597,N_10799,N_10579);
nor U12598 (N_12598,N_11241,N_11500);
nor U12599 (N_12599,N_10638,N_11226);
nor U12600 (N_12600,N_9010,N_11428);
nand U12601 (N_12601,N_10083,N_11128);
nand U12602 (N_12602,N_9884,N_10397);
xnor U12603 (N_12603,N_9783,N_9480);
and U12604 (N_12604,N_10947,N_10770);
xnor U12605 (N_12605,N_11599,N_10726);
nor U12606 (N_12606,N_10867,N_11392);
and U12607 (N_12607,N_10027,N_10299);
nor U12608 (N_12608,N_11828,N_11439);
and U12609 (N_12609,N_9088,N_9074);
nand U12610 (N_12610,N_11934,N_11338);
xnor U12611 (N_12611,N_11885,N_11785);
or U12612 (N_12612,N_11546,N_10471);
nor U12613 (N_12613,N_9828,N_11591);
or U12614 (N_12614,N_10580,N_10052);
nor U12615 (N_12615,N_11873,N_11448);
and U12616 (N_12616,N_9615,N_11856);
nand U12617 (N_12617,N_10687,N_11991);
nand U12618 (N_12618,N_10554,N_11412);
nand U12619 (N_12619,N_10378,N_10732);
nor U12620 (N_12620,N_10821,N_9747);
and U12621 (N_12621,N_10797,N_11722);
and U12622 (N_12622,N_9326,N_11624);
or U12623 (N_12623,N_9411,N_9532);
nand U12624 (N_12624,N_11769,N_10541);
nor U12625 (N_12625,N_9930,N_9655);
xor U12626 (N_12626,N_10946,N_11113);
or U12627 (N_12627,N_9583,N_9508);
or U12628 (N_12628,N_11711,N_9989);
and U12629 (N_12629,N_11709,N_9820);
nand U12630 (N_12630,N_11619,N_11648);
nand U12631 (N_12631,N_11483,N_11145);
or U12632 (N_12632,N_10682,N_9306);
nor U12633 (N_12633,N_9597,N_10169);
nor U12634 (N_12634,N_10304,N_11507);
and U12635 (N_12635,N_11385,N_10412);
or U12636 (N_12636,N_9734,N_9298);
nand U12637 (N_12637,N_11875,N_10780);
nand U12638 (N_12638,N_11831,N_11973);
or U12639 (N_12639,N_9614,N_11060);
nor U12640 (N_12640,N_10263,N_11553);
or U12641 (N_12641,N_10255,N_9926);
and U12642 (N_12642,N_11860,N_10735);
and U12643 (N_12643,N_10369,N_11358);
and U12644 (N_12644,N_9748,N_9674);
nor U12645 (N_12645,N_11440,N_9918);
nand U12646 (N_12646,N_10354,N_9062);
or U12647 (N_12647,N_11015,N_10138);
xor U12648 (N_12648,N_9376,N_11969);
or U12649 (N_12649,N_11812,N_10358);
or U12650 (N_12650,N_10284,N_10825);
and U12651 (N_12651,N_10003,N_9395);
nor U12652 (N_12652,N_10737,N_10001);
xnor U12653 (N_12653,N_9402,N_11921);
nor U12654 (N_12654,N_10769,N_9069);
nand U12655 (N_12655,N_10177,N_11807);
nor U12656 (N_12656,N_11931,N_11384);
or U12657 (N_12657,N_9311,N_9729);
or U12658 (N_12658,N_9423,N_11938);
and U12659 (N_12659,N_10463,N_9460);
nor U12660 (N_12660,N_11670,N_9571);
nand U12661 (N_12661,N_10076,N_9104);
or U12662 (N_12662,N_10213,N_10135);
nor U12663 (N_12663,N_11950,N_11231);
and U12664 (N_12664,N_10691,N_9396);
nor U12665 (N_12665,N_11869,N_11628);
nand U12666 (N_12666,N_10830,N_9702);
nor U12667 (N_12667,N_10608,N_9436);
and U12668 (N_12668,N_11646,N_9213);
and U12669 (N_12669,N_9866,N_11918);
nor U12670 (N_12670,N_11352,N_9415);
or U12671 (N_12671,N_11105,N_10623);
nand U12672 (N_12672,N_11014,N_10700);
xnor U12673 (N_12673,N_9932,N_9053);
nor U12674 (N_12674,N_11878,N_11180);
nand U12675 (N_12675,N_10043,N_9324);
and U12676 (N_12676,N_10336,N_10250);
nand U12677 (N_12677,N_10150,N_10655);
and U12678 (N_12678,N_9231,N_10446);
xor U12679 (N_12679,N_10892,N_10924);
nand U12680 (N_12680,N_11460,N_9819);
xnor U12681 (N_12681,N_9155,N_11419);
or U12682 (N_12682,N_10908,N_10679);
or U12683 (N_12683,N_10262,N_9225);
nand U12684 (N_12684,N_10957,N_10116);
or U12685 (N_12685,N_9873,N_10218);
or U12686 (N_12686,N_9657,N_10791);
or U12687 (N_12687,N_10846,N_11336);
nor U12688 (N_12688,N_10748,N_9561);
and U12689 (N_12689,N_10756,N_11924);
or U12690 (N_12690,N_9365,N_10971);
nor U12691 (N_12691,N_11675,N_9899);
or U12692 (N_12692,N_11214,N_9570);
and U12693 (N_12693,N_11851,N_10833);
nand U12694 (N_12694,N_10012,N_11674);
nor U12695 (N_12695,N_11142,N_9741);
or U12696 (N_12696,N_10787,N_9387);
and U12697 (N_12697,N_11715,N_10749);
nor U12698 (N_12698,N_9684,N_11661);
nor U12699 (N_12699,N_10443,N_10491);
or U12700 (N_12700,N_10488,N_11662);
and U12701 (N_12701,N_10386,N_9420);
xor U12702 (N_12702,N_9549,N_11744);
or U12703 (N_12703,N_9362,N_10876);
or U12704 (N_12704,N_9653,N_11590);
or U12705 (N_12705,N_11557,N_10247);
nor U12706 (N_12706,N_9484,N_9401);
nand U12707 (N_12707,N_10863,N_10176);
and U12708 (N_12708,N_11260,N_9912);
xnor U12709 (N_12709,N_9119,N_9594);
nand U12710 (N_12710,N_9774,N_10186);
or U12711 (N_12711,N_9035,N_11033);
nor U12712 (N_12712,N_10889,N_11829);
nand U12713 (N_12713,N_9641,N_11859);
nand U12714 (N_12714,N_11204,N_9332);
nor U12715 (N_12715,N_10850,N_10644);
and U12716 (N_12716,N_11701,N_10286);
and U12717 (N_12717,N_11610,N_11780);
xor U12718 (N_12718,N_9605,N_11953);
or U12719 (N_12719,N_9476,N_9164);
nor U12720 (N_12720,N_9518,N_9673);
nand U12721 (N_12721,N_9610,N_10124);
or U12722 (N_12722,N_10819,N_10225);
nand U12723 (N_12723,N_11839,N_9737);
and U12724 (N_12724,N_10631,N_11990);
or U12725 (N_12725,N_11259,N_10861);
or U12726 (N_12726,N_11645,N_10167);
or U12727 (N_12727,N_9193,N_9892);
nand U12728 (N_12728,N_11941,N_9448);
xor U12729 (N_12729,N_10137,N_9063);
nor U12730 (N_12730,N_9880,N_10750);
nand U12731 (N_12731,N_9342,N_10178);
or U12732 (N_12732,N_11479,N_11293);
xor U12733 (N_12733,N_9595,N_11401);
or U12734 (N_12734,N_9654,N_9126);
and U12735 (N_12735,N_9542,N_10201);
xnor U12736 (N_12736,N_9808,N_10590);
xor U12737 (N_12737,N_9864,N_9352);
and U12738 (N_12738,N_10599,N_11996);
nand U12739 (N_12739,N_10039,N_10017);
nand U12740 (N_12740,N_11053,N_9756);
nor U12741 (N_12741,N_9778,N_11863);
and U12742 (N_12742,N_10738,N_11362);
xor U12743 (N_12743,N_11239,N_11911);
and U12744 (N_12744,N_10455,N_9676);
and U12745 (N_12745,N_10870,N_10605);
nand U12746 (N_12746,N_11999,N_11258);
and U12747 (N_12747,N_9044,N_9715);
xnor U12748 (N_12748,N_9349,N_11212);
and U12749 (N_12749,N_11095,N_11035);
or U12750 (N_12750,N_11748,N_9897);
nand U12751 (N_12751,N_11928,N_9642);
or U12752 (N_12752,N_11209,N_11353);
nand U12753 (N_12753,N_9559,N_11192);
nor U12754 (N_12754,N_9369,N_9374);
and U12755 (N_12755,N_9223,N_10952);
xnor U12756 (N_12756,N_10920,N_10254);
or U12757 (N_12757,N_11888,N_10672);
and U12758 (N_12758,N_10196,N_10237);
and U12759 (N_12759,N_10643,N_11568);
xnor U12760 (N_12760,N_10844,N_11343);
or U12761 (N_12761,N_9981,N_10032);
nor U12762 (N_12762,N_10656,N_9277);
xnor U12763 (N_12763,N_10937,N_9604);
nor U12764 (N_12764,N_11489,N_10309);
nand U12765 (N_12765,N_9121,N_9901);
nor U12766 (N_12766,N_10393,N_11763);
and U12767 (N_12767,N_11861,N_9148);
xor U12768 (N_12768,N_10916,N_11429);
and U12769 (N_12769,N_9165,N_9707);
nand U12770 (N_12770,N_10366,N_10368);
nor U12771 (N_12771,N_10384,N_9962);
nand U12772 (N_12772,N_10664,N_9382);
nor U12773 (N_12773,N_10997,N_9370);
nand U12774 (N_12774,N_9018,N_10292);
or U12775 (N_12775,N_9259,N_11498);
xor U12776 (N_12776,N_10219,N_9844);
xnor U12777 (N_12777,N_11187,N_9548);
nand U12778 (N_12778,N_11091,N_10736);
nor U12779 (N_12779,N_9764,N_10303);
nand U12780 (N_12780,N_9287,N_9322);
nor U12781 (N_12781,N_9849,N_10215);
nand U12782 (N_12782,N_11653,N_9860);
nand U12783 (N_12783,N_9351,N_10249);
nand U12784 (N_12784,N_10793,N_9022);
nor U12785 (N_12785,N_10517,N_10337);
and U12786 (N_12786,N_11410,N_9442);
or U12787 (N_12787,N_9717,N_11783);
xor U12788 (N_12788,N_10454,N_10792);
nand U12789 (N_12789,N_11751,N_9354);
or U12790 (N_12790,N_10670,N_11552);
nand U12791 (N_12791,N_11472,N_10874);
nand U12792 (N_12792,N_11080,N_11109);
xor U12793 (N_12793,N_10667,N_11215);
or U12794 (N_12794,N_11671,N_10070);
or U12795 (N_12795,N_11631,N_9887);
and U12796 (N_12796,N_11381,N_10675);
or U12797 (N_12797,N_10913,N_9973);
nor U12798 (N_12798,N_9128,N_10527);
or U12799 (N_12799,N_10941,N_9243);
nor U12800 (N_12800,N_11723,N_10883);
or U12801 (N_12801,N_9782,N_11547);
nor U12802 (N_12802,N_10187,N_9033);
or U12803 (N_12803,N_9677,N_9404);
nor U12804 (N_12804,N_9075,N_10864);
nor U12805 (N_12805,N_10785,N_9524);
xor U12806 (N_12806,N_10596,N_11156);
xnor U12807 (N_12807,N_11304,N_9344);
nor U12808 (N_12808,N_9836,N_11897);
xnor U12809 (N_12809,N_10077,N_11167);
and U12810 (N_12810,N_10809,N_9872);
xnor U12811 (N_12811,N_11892,N_10049);
xnor U12812 (N_12812,N_10300,N_11824);
and U12813 (N_12813,N_9242,N_9206);
nor U12814 (N_12814,N_9204,N_9792);
nand U12815 (N_12815,N_11016,N_10501);
or U12816 (N_12816,N_10552,N_11003);
xor U12817 (N_12817,N_9997,N_9987);
nand U12818 (N_12818,N_10353,N_10849);
xnor U12819 (N_12819,N_9772,N_10008);
and U12820 (N_12820,N_10891,N_9264);
nor U12821 (N_12821,N_9317,N_10775);
or U12822 (N_12822,N_11062,N_11558);
xor U12823 (N_12823,N_9934,N_9948);
xnor U12824 (N_12824,N_10246,N_11034);
or U12825 (N_12825,N_9913,N_11724);
or U12826 (N_12826,N_10693,N_11028);
nand U12827 (N_12827,N_9274,N_9767);
xnor U12828 (N_12828,N_10184,N_9619);
nor U12829 (N_12829,N_11290,N_10890);
and U12830 (N_12830,N_10229,N_11581);
nand U12831 (N_12831,N_9159,N_11426);
and U12832 (N_12832,N_10163,N_9339);
xor U12833 (N_12833,N_11090,N_10840);
nor U12834 (N_12834,N_9007,N_11471);
nand U12835 (N_12835,N_10714,N_11767);
or U12836 (N_12836,N_9117,N_9688);
or U12837 (N_12837,N_9920,N_10115);
xor U12838 (N_12838,N_9522,N_11322);
and U12839 (N_12839,N_9434,N_9267);
nor U12840 (N_12840,N_11533,N_9454);
nor U12841 (N_12841,N_10719,N_11712);
or U12842 (N_12842,N_11468,N_9445);
nor U12843 (N_12843,N_11618,N_9438);
or U12844 (N_12844,N_9833,N_9716);
xor U12845 (N_12845,N_11274,N_10002);
nor U12846 (N_12846,N_11627,N_11269);
nor U12847 (N_12847,N_9723,N_9424);
and U12848 (N_12848,N_9879,N_10066);
nand U12849 (N_12849,N_11636,N_9555);
nor U12850 (N_12850,N_9881,N_9727);
nor U12851 (N_12851,N_10831,N_9304);
and U12852 (N_12852,N_10767,N_10744);
nor U12853 (N_12853,N_9341,N_9970);
nand U12854 (N_12854,N_10481,N_9647);
nor U12855 (N_12855,N_9073,N_9110);
nand U12856 (N_12856,N_11340,N_10430);
nor U12857 (N_12857,N_9988,N_11929);
and U12858 (N_12858,N_9667,N_10310);
xor U12859 (N_12859,N_10014,N_10464);
and U12860 (N_12860,N_11520,N_10964);
nor U12861 (N_12861,N_9157,N_9472);
nor U12862 (N_12862,N_9181,N_9961);
nor U12863 (N_12863,N_11535,N_11213);
xnor U12864 (N_12864,N_11497,N_9194);
xor U12865 (N_12865,N_10434,N_9041);
and U12866 (N_12866,N_9855,N_11638);
and U12867 (N_12867,N_9908,N_10746);
or U12868 (N_12868,N_11083,N_10198);
or U12869 (N_12869,N_9580,N_10047);
and U12870 (N_12870,N_11491,N_10765);
xor U12871 (N_12871,N_9995,N_11838);
or U12872 (N_12872,N_10327,N_9268);
nor U12873 (N_12873,N_11039,N_9638);
and U12874 (N_12874,N_11208,N_10707);
nand U12875 (N_12875,N_11791,N_11515);
nor U12876 (N_12876,N_11441,N_11815);
nor U12877 (N_12877,N_10161,N_9650);
nand U12878 (N_12878,N_11773,N_9185);
nand U12879 (N_12879,N_9903,N_10991);
xor U12880 (N_12880,N_9681,N_10877);
nand U12881 (N_12881,N_11629,N_11394);
or U12882 (N_12882,N_10216,N_10414);
or U12883 (N_12883,N_9957,N_11037);
nor U12884 (N_12884,N_9501,N_11562);
nor U12885 (N_12885,N_9386,N_9281);
or U12886 (N_12886,N_9687,N_10640);
nor U12887 (N_12887,N_10701,N_11643);
or U12888 (N_12888,N_11840,N_10551);
and U12889 (N_12889,N_11297,N_11587);
and U12890 (N_12890,N_9421,N_10690);
or U12891 (N_12891,N_11178,N_10930);
or U12892 (N_12892,N_11865,N_9617);
or U12893 (N_12893,N_11454,N_10660);
or U12894 (N_12894,N_10953,N_9956);
and U12895 (N_12895,N_9878,N_10627);
nand U12896 (N_12896,N_9334,N_11162);
nor U12897 (N_12897,N_11574,N_9562);
nor U12898 (N_12898,N_11216,N_10425);
or U12899 (N_12899,N_9483,N_10416);
and U12900 (N_12900,N_9008,N_11073);
nand U12901 (N_12901,N_10822,N_10529);
xor U12902 (N_12902,N_10715,N_11055);
xnor U12903 (N_12903,N_9787,N_11584);
and U12904 (N_12904,N_9201,N_11669);
or U12905 (N_12905,N_9869,N_10498);
xor U12906 (N_12906,N_11235,N_11138);
or U12907 (N_12907,N_9893,N_9474);
nor U12908 (N_12908,N_10773,N_10794);
or U12909 (N_12909,N_9495,N_10193);
and U12910 (N_12910,N_9469,N_11219);
nand U12911 (N_12911,N_10084,N_11081);
or U12912 (N_12912,N_11397,N_10038);
or U12913 (N_12913,N_10741,N_11496);
nor U12914 (N_12914,N_11693,N_10050);
and U12915 (N_12915,N_9815,N_9904);
nor U12916 (N_12916,N_10852,N_10060);
xnor U12917 (N_12917,N_10276,N_11330);
xor U12918 (N_12918,N_11905,N_11054);
nor U12919 (N_12919,N_11677,N_10595);
nor U12920 (N_12920,N_11548,N_11798);
nor U12921 (N_12921,N_11956,N_9954);
nand U12922 (N_12922,N_9003,N_9379);
nor U12923 (N_12923,N_10405,N_9603);
xor U12924 (N_12924,N_9754,N_11115);
and U12925 (N_12925,N_9824,N_9109);
or U12926 (N_12926,N_9917,N_10562);
nor U12927 (N_12927,N_9714,N_11393);
nor U12928 (N_12928,N_10395,N_9209);
or U12929 (N_12929,N_9563,N_10101);
and U12930 (N_12930,N_10174,N_9806);
nand U12931 (N_12931,N_11955,N_10316);
and U12932 (N_12932,N_10513,N_9906);
or U12933 (N_12933,N_9032,N_11386);
nand U12934 (N_12934,N_10221,N_10091);
and U12935 (N_12935,N_9945,N_10786);
nor U12936 (N_12936,N_11007,N_10442);
nor U12937 (N_12937,N_10330,N_9162);
xnor U12938 (N_12938,N_11958,N_11466);
and U12939 (N_12939,N_10383,N_11433);
xor U12940 (N_12940,N_9111,N_11766);
nand U12941 (N_12941,N_11923,N_11825);
and U12942 (N_12942,N_10415,N_9108);
nor U12943 (N_12943,N_11788,N_11414);
xnor U12944 (N_12944,N_11834,N_11787);
nor U12945 (N_12945,N_11971,N_9922);
nand U12946 (N_12946,N_11717,N_10652);
xnor U12947 (N_12947,N_10938,N_9114);
nor U12948 (N_12948,N_9531,N_10751);
xnor U12949 (N_12949,N_10560,N_10747);
nand U12950 (N_12950,N_10320,N_9763);
or U12951 (N_12951,N_9867,N_10589);
or U12952 (N_12952,N_11289,N_10448);
nand U12953 (N_12953,N_9245,N_9994);
nor U12954 (N_12954,N_10111,N_9535);
nor U12955 (N_12955,N_10973,N_10983);
nor U12956 (N_12956,N_9078,N_10600);
nor U12957 (N_12957,N_9882,N_10827);
or U12958 (N_12958,N_9400,N_10533);
and U12959 (N_12959,N_11254,N_9391);
or U12960 (N_12960,N_9804,N_9585);
or U12961 (N_12961,N_9661,N_11047);
or U12962 (N_12962,N_9059,N_11607);
xnor U12963 (N_12963,N_10636,N_10881);
nor U12964 (N_12964,N_10847,N_10119);
nand U12965 (N_12965,N_11764,N_9456);
nand U12966 (N_12966,N_11139,N_10090);
and U12967 (N_12967,N_9543,N_10371);
or U12968 (N_12968,N_10694,N_10171);
nand U12969 (N_12969,N_9516,N_11900);
nor U12970 (N_12970,N_9799,N_11862);
nor U12971 (N_12971,N_9293,N_10261);
nor U12972 (N_12972,N_11474,N_9428);
xnor U12973 (N_12973,N_11200,N_9237);
or U12974 (N_12974,N_11845,N_9858);
nor U12975 (N_12975,N_9187,N_9533);
nor U12976 (N_12976,N_11464,N_10650);
and U12977 (N_12977,N_10661,N_11739);
nor U12978 (N_12978,N_10143,N_10317);
or U12979 (N_12979,N_9846,N_10045);
and U12980 (N_12980,N_11312,N_10279);
xor U12981 (N_12981,N_10855,N_11966);
or U12982 (N_12982,N_9048,N_9958);
xor U12983 (N_12983,N_10507,N_11166);
nand U12984 (N_12984,N_11720,N_10387);
nand U12985 (N_12985,N_11306,N_9014);
xor U12986 (N_12986,N_10720,N_11422);
nand U12987 (N_12987,N_10810,N_11435);
and U12988 (N_12988,N_11119,N_9829);
nand U12989 (N_12989,N_9098,N_11218);
nand U12990 (N_12990,N_9803,N_10555);
nor U12991 (N_12991,N_10391,N_10183);
xor U12992 (N_12992,N_10435,N_9133);
or U12993 (N_12993,N_10087,N_10919);
or U12994 (N_12994,N_11903,N_10048);
and U12995 (N_12995,N_10621,N_10918);
or U12996 (N_12996,N_10635,N_11596);
or U12997 (N_12997,N_9066,N_11032);
nor U12998 (N_12998,N_11453,N_11057);
xnor U12999 (N_12999,N_9827,N_9900);
xor U13000 (N_13000,N_10757,N_10681);
nor U13001 (N_13001,N_11757,N_9991);
xor U13002 (N_13002,N_9444,N_11288);
nand U13003 (N_13003,N_9312,N_10702);
nand U13004 (N_13004,N_10798,N_9554);
and U13005 (N_13005,N_10662,N_9102);
nor U13006 (N_13006,N_10666,N_10689);
nand U13007 (N_13007,N_10985,N_9049);
nor U13008 (N_13008,N_9902,N_11253);
xnor U13009 (N_13009,N_9975,N_10062);
or U13010 (N_13010,N_11970,N_9565);
nor U13011 (N_13011,N_11004,N_11655);
or U13012 (N_13012,N_10329,N_11817);
or U13013 (N_13013,N_11816,N_11009);
nor U13014 (N_13014,N_9115,N_9569);
nor U13015 (N_13015,N_10632,N_9623);
nor U13016 (N_13016,N_11074,N_9186);
nor U13017 (N_13017,N_11262,N_10182);
nand U13018 (N_13018,N_11396,N_9012);
nor U13019 (N_13019,N_9435,N_9923);
nand U13020 (N_13020,N_11813,N_9375);
and U13021 (N_13021,N_10370,N_11620);
nor U13022 (N_13022,N_9646,N_11475);
and U13023 (N_13023,N_9812,N_11155);
or U13024 (N_13024,N_10880,N_11130);
nand U13025 (N_13025,N_10069,N_9505);
and U13026 (N_13026,N_10364,N_9999);
and U13027 (N_13027,N_9996,N_11050);
or U13028 (N_13028,N_9394,N_10082);
nand U13029 (N_13029,N_9005,N_10117);
xnor U13030 (N_13030,N_11416,N_10344);
nand U13031 (N_13031,N_9016,N_11465);
nor U13032 (N_13032,N_10530,N_10712);
and U13033 (N_13033,N_9233,N_10152);
and U13034 (N_13034,N_10586,N_10418);
nor U13035 (N_13035,N_9096,N_9381);
nand U13036 (N_13036,N_10204,N_9601);
and U13037 (N_13037,N_9822,N_11418);
and U13038 (N_13038,N_10943,N_9336);
nor U13039 (N_13039,N_10708,N_11124);
nor U13040 (N_13040,N_9405,N_10331);
nand U13041 (N_13041,N_11710,N_11485);
xor U13042 (N_13042,N_10287,N_9234);
nor U13043 (N_13043,N_9138,N_9238);
or U13044 (N_13044,N_11585,N_11563);
nor U13045 (N_13045,N_11402,N_11434);
xnor U13046 (N_13046,N_9972,N_9998);
nand U13047 (N_13047,N_10389,N_11161);
nor U13048 (N_13048,N_10776,N_11719);
nor U13049 (N_13049,N_9272,N_10618);
nand U13050 (N_13050,N_10380,N_9120);
nand U13051 (N_13051,N_11427,N_11461);
nand U13052 (N_13052,N_10421,N_10620);
nand U13053 (N_13053,N_10603,N_11556);
or U13054 (N_13054,N_9089,N_10993);
nand U13055 (N_13055,N_9620,N_9698);
nor U13056 (N_13056,N_11064,N_9793);
nand U13057 (N_13057,N_11809,N_11143);
or U13058 (N_13058,N_9222,N_11771);
and U13059 (N_13059,N_10725,N_11992);
and U13060 (N_13060,N_11797,N_11318);
nor U13061 (N_13061,N_9976,N_10709);
or U13062 (N_13062,N_11337,N_10521);
or U13063 (N_13063,N_11803,N_11510);
or U13064 (N_13064,N_9229,N_10729);
or U13065 (N_13065,N_11324,N_11939);
and U13066 (N_13066,N_11373,N_10970);
and U13067 (N_13067,N_9380,N_10121);
and U13068 (N_13068,N_10940,N_11457);
or U13069 (N_13069,N_9284,N_10106);
and U13070 (N_13070,N_10291,N_9137);
nand U13071 (N_13071,N_10593,N_10308);
nand U13072 (N_13072,N_9942,N_9366);
nand U13073 (N_13073,N_10845,N_10853);
nand U13074 (N_13074,N_11889,N_11315);
or U13075 (N_13075,N_9084,N_10158);
or U13076 (N_13076,N_11981,N_11308);
or U13077 (N_13077,N_9294,N_9630);
or U13078 (N_13078,N_11298,N_10377);
or U13079 (N_13079,N_9693,N_9831);
nor U13080 (N_13080,N_9280,N_11598);
or U13081 (N_13081,N_10790,N_9939);
nand U13082 (N_13082,N_10782,N_9840);
and U13083 (N_13083,N_9584,N_10195);
nand U13084 (N_13084,N_9085,N_9721);
xor U13085 (N_13085,N_11473,N_9794);
nand U13086 (N_13086,N_9321,N_9135);
nand U13087 (N_13087,N_11604,N_11847);
nand U13088 (N_13088,N_11695,N_11285);
and U13089 (N_13089,N_11972,N_9432);
and U13090 (N_13090,N_11372,N_9141);
or U13091 (N_13091,N_11021,N_11041);
and U13092 (N_13092,N_10053,N_9506);
nor U13093 (N_13093,N_9475,N_10939);
or U13094 (N_13094,N_11741,N_9197);
xnor U13095 (N_13095,N_9378,N_10351);
xor U13096 (N_13096,N_11376,N_11043);
and U13097 (N_13097,N_9805,N_11210);
xnor U13098 (N_13098,N_10626,N_9446);
xnor U13099 (N_13099,N_9397,N_9407);
nand U13100 (N_13100,N_10975,N_10949);
and U13101 (N_13101,N_11841,N_10716);
and U13102 (N_13102,N_11554,N_9552);
nor U13103 (N_13103,N_11871,N_9118);
xor U13104 (N_13104,N_10515,N_10931);
nor U13105 (N_13105,N_10217,N_9357);
nor U13106 (N_13106,N_9980,N_11147);
nor U13107 (N_13107,N_11732,N_10796);
nor U13108 (N_13108,N_11647,N_10024);
or U13109 (N_13109,N_11022,N_10884);
xor U13110 (N_13110,N_10649,N_9079);
nand U13111 (N_13111,N_11085,N_11375);
and U13112 (N_13112,N_10999,N_9359);
xor U13113 (N_13113,N_10298,N_10648);
or U13114 (N_13114,N_10869,N_10265);
nand U13115 (N_13115,N_10168,N_9540);
nor U13116 (N_13116,N_9503,N_11755);
nor U13117 (N_13117,N_9301,N_11541);
nor U13118 (N_13118,N_9190,N_9511);
or U13119 (N_13119,N_9891,N_10162);
nor U13120 (N_13120,N_11867,N_10496);
or U13121 (N_13121,N_11099,N_11190);
or U13122 (N_13122,N_10520,N_9361);
and U13123 (N_13123,N_10569,N_11313);
or U13124 (N_13124,N_9659,N_9132);
and U13125 (N_13125,N_10426,N_11602);
nor U13126 (N_13126,N_11979,N_10537);
nor U13127 (N_13127,N_11945,N_10424);
nor U13128 (N_13128,N_10900,N_9441);
or U13129 (N_13129,N_10280,N_9750);
and U13130 (N_13130,N_11614,N_11884);
and U13131 (N_13131,N_11765,N_9510);
nand U13132 (N_13132,N_9310,N_10283);
nor U13133 (N_13133,N_9015,N_9633);
nor U13134 (N_13134,N_11555,N_10305);
xnor U13135 (N_13135,N_10759,N_10606);
nand U13136 (N_13136,N_10933,N_9766);
nand U13137 (N_13137,N_11932,N_10851);
nand U13138 (N_13138,N_11569,N_9699);
nand U13139 (N_13139,N_10166,N_11374);
nor U13140 (N_13140,N_9451,N_9377);
nand U13141 (N_13141,N_10645,N_11359);
xnor U13142 (N_13142,N_9409,N_11150);
or U13143 (N_13143,N_9218,N_11794);
and U13144 (N_13144,N_9318,N_10842);
and U13145 (N_13145,N_11879,N_10651);
and U13146 (N_13146,N_11632,N_9315);
and U13147 (N_13147,N_10743,N_11806);
and U13148 (N_13148,N_10795,N_9171);
nor U13149 (N_13149,N_10081,N_11976);
and U13150 (N_13150,N_11682,N_10398);
nand U13151 (N_13151,N_10335,N_10483);
nand U13152 (N_13152,N_10312,N_9308);
nor U13153 (N_13153,N_10909,N_10409);
nand U13154 (N_13154,N_10022,N_11626);
and U13155 (N_13155,N_9443,N_9865);
or U13156 (N_13156,N_10497,N_10374);
and U13157 (N_13157,N_11890,N_10092);
nor U13158 (N_13158,N_10144,N_10339);
nand U13159 (N_13159,N_11126,N_10275);
nor U13160 (N_13160,N_9695,N_11286);
or U13161 (N_13161,N_10935,N_10477);
nand U13162 (N_13162,N_9207,N_10365);
and U13163 (N_13163,N_10685,N_11133);
nor U13164 (N_13164,N_9047,N_10155);
and U13165 (N_13165,N_10557,N_11217);
xnor U13166 (N_13166,N_10955,N_9227);
nor U13167 (N_13167,N_10669,N_9575);
nand U13168 (N_13168,N_10422,N_11502);
nand U13169 (N_13169,N_9179,N_10536);
and U13170 (N_13170,N_11469,N_9916);
and U13171 (N_13171,N_9093,N_10678);
or U13172 (N_13172,N_9539,N_9482);
xnor U13173 (N_13173,N_10342,N_11284);
nor U13174 (N_13174,N_9502,N_9149);
nor U13175 (N_13175,N_9070,N_10804);
nand U13176 (N_13176,N_11793,N_11017);
xnor U13177 (N_13177,N_9965,N_10452);
nand U13178 (N_13178,N_10326,N_10572);
xnor U13179 (N_13179,N_11347,N_11271);
or U13180 (N_13180,N_9350,N_11456);
nand U13181 (N_13181,N_11420,N_11937);
and U13182 (N_13182,N_10086,N_9613);
nand U13183 (N_13183,N_10503,N_10493);
nand U13184 (N_13184,N_9982,N_9323);
and U13185 (N_13185,N_10692,N_10479);
nand U13186 (N_13186,N_10044,N_11189);
and U13187 (N_13187,N_9112,N_9124);
and U13188 (N_13188,N_11459,N_9071);
or U13189 (N_13189,N_10906,N_9219);
or U13190 (N_13190,N_9830,N_11432);
nand U13191 (N_13191,N_11786,N_11665);
nor U13192 (N_13192,N_9921,N_11038);
and U13193 (N_13193,N_11492,N_11087);
and U13194 (N_13194,N_10871,N_11387);
and U13195 (N_13195,N_10545,N_9927);
xor U13196 (N_13196,N_9526,N_10663);
xor U13197 (N_13197,N_11849,N_10277);
or U13198 (N_13198,N_9728,N_9634);
xor U13199 (N_13199,N_9113,N_9590);
or U13200 (N_13200,N_10315,N_10987);
or U13201 (N_13201,N_10910,N_11431);
nor U13202 (N_13202,N_10582,N_9582);
and U13203 (N_13203,N_11169,N_11988);
nand U13204 (N_13204,N_10141,N_9845);
or U13205 (N_13205,N_10887,N_11252);
nand U13206 (N_13206,N_9300,N_11421);
and U13207 (N_13207,N_10563,N_11010);
nand U13208 (N_13208,N_9461,N_10228);
nor U13209 (N_13209,N_9731,N_10288);
nand U13210 (N_13210,N_11942,N_9682);
or U13211 (N_13211,N_11294,N_10223);
or U13212 (N_13212,N_11223,N_9251);
and U13213 (N_13213,N_11761,N_9358);
nor U13214 (N_13214,N_11356,N_9898);
nand U13215 (N_13215,N_10888,N_11391);
nand U13216 (N_13216,N_9340,N_11716);
or U13217 (N_13217,N_10411,N_11947);
or U13218 (N_13218,N_10574,N_11689);
or U13219 (N_13219,N_9017,N_9788);
or U13220 (N_13220,N_11165,N_10610);
nor U13221 (N_13221,N_10140,N_10457);
nand U13222 (N_13222,N_9816,N_9198);
or U13223 (N_13223,N_10966,N_9743);
nor U13224 (N_13224,N_10781,N_9153);
or U13225 (N_13225,N_11300,N_11779);
nor U13226 (N_13226,N_9666,N_10388);
or U13227 (N_13227,N_9123,N_9260);
nand U13228 (N_13228,N_10456,N_10073);
nand U13229 (N_13229,N_9600,N_11742);
or U13230 (N_13230,N_10480,N_11186);
nor U13231 (N_13231,N_10172,N_11423);
nand U13232 (N_13232,N_11205,N_9303);
nand U13233 (N_13233,N_10907,N_11036);
and U13234 (N_13234,N_10175,N_10469);
or U13235 (N_13235,N_10516,N_9184);
xor U13236 (N_13236,N_10893,N_10447);
and U13237 (N_13237,N_9449,N_11168);
nand U13238 (N_13238,N_9874,N_11341);
nor U13239 (N_13239,N_11886,N_10784);
and U13240 (N_13240,N_11656,N_10011);
and U13241 (N_13241,N_11065,N_9726);
nand U13242 (N_13242,N_11756,N_11836);
or U13243 (N_13243,N_11866,N_10854);
and U13244 (N_13244,N_10839,N_10629);
nor U13245 (N_13245,N_11804,N_9416);
nand U13246 (N_13246,N_10724,N_11985);
nor U13247 (N_13247,N_9080,N_9001);
nand U13248 (N_13248,N_11660,N_11519);
nor U13249 (N_13249,N_11413,N_9384);
or U13250 (N_13250,N_11959,N_11727);
or U13251 (N_13251,N_9057,N_9553);
nand U13252 (N_13252,N_9305,N_11151);
xnor U13253 (N_13253,N_11044,N_11114);
xor U13254 (N_13254,N_9309,N_11030);
and U13255 (N_13255,N_10570,N_11810);
nand U13256 (N_13256,N_10980,N_10147);
or U13257 (N_13257,N_11311,N_9002);
nand U13258 (N_13258,N_10565,N_10200);
nor U13259 (N_13259,N_10929,N_11398);
nand U13260 (N_13260,N_9142,N_11106);
xor U13261 (N_13261,N_9809,N_11251);
or U13262 (N_13262,N_11850,N_10706);
nand U13263 (N_13263,N_11792,N_11573);
xor U13264 (N_13264,N_10165,N_10034);
nand U13265 (N_13265,N_9028,N_11328);
nand U13266 (N_13266,N_9055,N_11509);
or U13267 (N_13267,N_10021,N_10613);
nand U13268 (N_13268,N_9205,N_10125);
and U13269 (N_13269,N_9826,N_11907);
xor U13270 (N_13270,N_9275,N_11571);
nand U13271 (N_13271,N_9356,N_9122);
xor U13272 (N_13272,N_9785,N_11305);
nand U13273 (N_13273,N_11342,N_11117);
nor U13274 (N_13274,N_10476,N_10206);
nand U13275 (N_13275,N_10634,N_9862);
and U13276 (N_13276,N_9103,N_9200);
and U13277 (N_13277,N_10466,N_11116);
and U13278 (N_13278,N_10324,N_10385);
nand U13279 (N_13279,N_11232,N_9696);
xnor U13280 (N_13280,N_10789,N_11775);
and U13281 (N_13281,N_10227,N_11517);
nor U13282 (N_13282,N_11963,N_9795);
nand U13283 (N_13283,N_9704,N_11314);
or U13284 (N_13284,N_10190,N_11901);
nand U13285 (N_13285,N_10637,N_10459);
and U13286 (N_13286,N_9250,N_10607);
xor U13287 (N_13287,N_11642,N_10814);
nand U13288 (N_13288,N_11977,N_10231);
nand U13289 (N_13289,N_11104,N_11678);
nor U13290 (N_13290,N_9166,N_11521);
nand U13291 (N_13291,N_10509,N_11997);
nor U13292 (N_13292,N_9455,N_11278);
and U13293 (N_13293,N_9255,N_11197);
nand U13294 (N_13294,N_11980,N_10041);
nand U13295 (N_13295,N_9252,N_11063);
or U13296 (N_13296,N_11449,N_11930);
and U13297 (N_13297,N_10511,N_10094);
nor U13298 (N_13298,N_11917,N_11799);
or U13299 (N_13299,N_10236,N_9025);
nor U13300 (N_13300,N_11530,N_10742);
nand U13301 (N_13301,N_9943,N_9399);
nor U13302 (N_13302,N_10485,N_10160);
or U13303 (N_13303,N_10878,N_11926);
and U13304 (N_13304,N_9150,N_11659);
nor U13305 (N_13305,N_10763,N_10934);
or U13306 (N_13306,N_10095,N_10282);
nand U13307 (N_13307,N_10345,N_10408);
or U13308 (N_13308,N_11894,N_10458);
nor U13309 (N_13309,N_9081,N_10054);
nand U13310 (N_13310,N_9302,N_9244);
and U13311 (N_13311,N_10752,N_10220);
nor U13312 (N_13312,N_9278,N_9249);
nor U13313 (N_13313,N_11781,N_10611);
xnor U13314 (N_13314,N_11108,N_11395);
nand U13315 (N_13315,N_11822,N_10376);
or U13316 (N_13316,N_9834,N_10433);
nand U13317 (N_13317,N_10926,N_11134);
nor U13318 (N_13318,N_10399,N_11417);
xor U13319 (N_13319,N_10209,N_10109);
or U13320 (N_13320,N_9701,N_9990);
or U13321 (N_13321,N_10404,N_10129);
nand U13322 (N_13322,N_10525,N_10547);
and U13323 (N_13323,N_11177,N_11070);
xor U13324 (N_13324,N_11257,N_11101);
and U13325 (N_13325,N_10146,N_9299);
nand U13326 (N_13326,N_11811,N_11774);
nor U13327 (N_13327,N_10403,N_10134);
or U13328 (N_13328,N_11071,N_9230);
nor U13329 (N_13329,N_11575,N_9658);
and U13330 (N_13330,N_11946,N_9538);
nand U13331 (N_13331,N_9986,N_10400);
or U13332 (N_13332,N_9560,N_10016);
or U13333 (N_13333,N_11578,N_10965);
and U13334 (N_13334,N_10959,N_10295);
nand U13335 (N_13335,N_10922,N_11784);
and U13336 (N_13336,N_11676,N_10419);
and U13337 (N_13337,N_11633,N_11898);
and U13338 (N_13338,N_11268,N_11652);
nor U13339 (N_13339,N_11325,N_9541);
nand U13340 (N_13340,N_11512,N_10302);
xor U13341 (N_13341,N_9791,N_9479);
or U13342 (N_13342,N_9692,N_10942);
nor U13343 (N_13343,N_10256,N_10774);
and U13344 (N_13344,N_10969,N_9850);
nand U13345 (N_13345,N_9054,N_11339);
or U13346 (N_13346,N_9746,N_10114);
and U13347 (N_13347,N_9875,N_9029);
or U13348 (N_13348,N_9368,N_10006);
nor U13349 (N_13349,N_10978,N_9811);
nand U13350 (N_13350,N_11623,N_11993);
nor U13351 (N_13351,N_9319,N_9265);
nand U13352 (N_13352,N_10963,N_10018);
nor U13353 (N_13353,N_9026,N_11011);
nor U13354 (N_13354,N_10721,N_11881);
nor U13355 (N_13355,N_11658,N_9266);
and U13356 (N_13356,N_11042,N_11951);
nand U13357 (N_13357,N_11561,N_10641);
nor U13358 (N_13358,N_9360,N_10058);
and U13359 (N_13359,N_11805,N_9215);
nand U13360 (N_13360,N_9863,N_10203);
and U13361 (N_13361,N_11194,N_11920);
nor U13362 (N_13362,N_10857,N_10438);
or U13363 (N_13363,N_10306,N_9720);
nor U13364 (N_13364,N_10120,N_11538);
xor U13365 (N_13365,N_10932,N_9910);
or U13366 (N_13366,N_10905,N_9485);
or U13367 (N_13367,N_10585,N_9841);
or U13368 (N_13368,N_9664,N_10617);
and U13369 (N_13369,N_9051,N_9021);
nand U13370 (N_13370,N_9740,N_10960);
and U13371 (N_13371,N_9974,N_11846);
nand U13372 (N_13372,N_11745,N_11564);
nand U13373 (N_13373,N_10601,N_9036);
and U13374 (N_13374,N_10986,N_11094);
xnor U13375 (N_13375,N_11592,N_10583);
or U13376 (N_13376,N_10566,N_11282);
nor U13377 (N_13377,N_9680,N_10244);
nand U13378 (N_13378,N_10731,N_9607);
xnor U13379 (N_13379,N_11853,N_10783);
nand U13380 (N_13380,N_9679,N_10903);
or U13381 (N_13381,N_9064,N_10604);
or U13382 (N_13382,N_11176,N_9593);
and U13383 (N_13383,N_11049,N_10740);
and U13384 (N_13384,N_9758,N_11430);
nor U13385 (N_13385,N_10133,N_10267);
and U13386 (N_13386,N_10362,N_9496);
nor U13387 (N_13387,N_9486,N_9557);
nand U13388 (N_13388,N_9177,N_11152);
xnor U13389 (N_13389,N_9246,N_9130);
nand U13390 (N_13390,N_10056,N_10894);
or U13391 (N_13391,N_11699,N_11936);
and U13392 (N_13392,N_11005,N_11684);
nand U13393 (N_13393,N_11916,N_11403);
or U13394 (N_13394,N_11256,N_9477);
nor U13395 (N_13395,N_9823,N_11234);
and U13396 (N_13396,N_9838,N_11320);
and U13397 (N_13397,N_10598,N_11801);
and U13398 (N_13398,N_11451,N_11163);
or U13399 (N_13399,N_10401,N_10373);
nand U13400 (N_13400,N_10653,N_11406);
or U13401 (N_13401,N_11843,N_10037);
nand U13402 (N_13402,N_9668,N_11059);
nor U13403 (N_13403,N_11295,N_9414);
or U13404 (N_13404,N_9801,N_10473);
nand U13405 (N_13405,N_11506,N_11499);
and U13406 (N_13406,N_11158,N_10592);
nor U13407 (N_13407,N_11082,N_9333);
nor U13408 (N_13408,N_9551,N_11910);
xor U13409 (N_13409,N_11818,N_11949);
or U13410 (N_13410,N_11954,N_9389);
and U13411 (N_13411,N_11202,N_9606);
or U13412 (N_13412,N_10548,N_10898);
nand U13413 (N_13413,N_9635,N_9883);
or U13414 (N_13414,N_9258,N_11327);
nand U13415 (N_13415,N_10067,N_10974);
nand U13416 (N_13416,N_9848,N_10921);
nor U13417 (N_13417,N_11415,N_11184);
and U13418 (N_13418,N_11754,N_11772);
nor U13419 (N_13419,N_10379,N_11698);
and U13420 (N_13420,N_11734,N_10979);
nor U13421 (N_13421,N_9188,N_9852);
and U13422 (N_13422,N_11518,N_10915);
and U13423 (N_13423,N_11283,N_10131);
or U13424 (N_13424,N_11345,N_10248);
and U13425 (N_13425,N_9821,N_10333);
nor U13426 (N_13426,N_11160,N_9814);
or U13427 (N_13427,N_9629,N_11462);
or U13428 (N_13428,N_11513,N_11272);
nand U13429 (N_13429,N_10816,N_11634);
nor U13430 (N_13430,N_10059,N_11616);
or U13431 (N_13431,N_10233,N_9525);
nor U13432 (N_13432,N_10982,N_11019);
and U13433 (N_13433,N_9288,N_10998);
nand U13434 (N_13434,N_10359,N_9798);
nand U13435 (N_13435,N_10232,N_10988);
or U13436 (N_13436,N_9060,N_9914);
and U13437 (N_13437,N_10698,N_10860);
and U13438 (N_13438,N_11536,N_9685);
nor U13439 (N_13439,N_9817,N_9146);
nor U13440 (N_13440,N_9346,N_10788);
and U13441 (N_13441,N_9097,N_10173);
or U13442 (N_13442,N_9626,N_11159);
or U13443 (N_13443,N_11249,N_10642);
nor U13444 (N_13444,N_11580,N_9431);
nor U13445 (N_13445,N_10205,N_11445);
or U13446 (N_13446,N_10118,N_9651);
or U13447 (N_13447,N_9529,N_10546);
and U13448 (N_13448,N_10252,N_9470);
nor U13449 (N_13449,N_10505,N_9027);
nor U13450 (N_13450,N_10078,N_9637);
nand U13451 (N_13451,N_10556,N_9931);
xor U13452 (N_13452,N_9622,N_9843);
and U13453 (N_13453,N_11264,N_11225);
and U13454 (N_13454,N_10674,N_10357);
nor U13455 (N_13455,N_9127,N_9757);
nor U13456 (N_13456,N_11984,N_9790);
nor U13457 (N_13457,N_9678,N_11107);
nor U13458 (N_13458,N_11020,N_11276);
nand U13459 (N_13459,N_11400,N_9030);
nand U13460 (N_13460,N_10420,N_11261);
nor U13461 (N_13461,N_9466,N_9587);
nor U13462 (N_13462,N_10951,N_9708);
nor U13463 (N_13463,N_11872,N_9624);
or U13464 (N_13464,N_11730,N_11935);
nand U13465 (N_13465,N_9465,N_9425);
nand U13466 (N_13466,N_11844,N_9270);
or U13467 (N_13467,N_10494,N_10042);
nand U13468 (N_13468,N_9789,N_11317);
nand U13469 (N_13469,N_9978,N_11758);
nor U13470 (N_13470,N_9086,N_11887);
or U13471 (N_13471,N_11789,N_11296);
nor U13472 (N_13472,N_11236,N_11477);
or U13473 (N_13473,N_11559,N_11790);
or U13474 (N_13474,N_10584,N_9837);
xnor U13475 (N_13475,N_10490,N_10571);
and U13476 (N_13476,N_10406,N_11703);
or U13477 (N_13477,N_11915,N_11697);
nor U13478 (N_13478,N_11718,N_10630);
and U13479 (N_13479,N_10222,N_10730);
or U13480 (N_13480,N_9314,N_9662);
nand U13481 (N_13481,N_10824,N_11848);
or U13482 (N_13482,N_11650,N_10896);
xor U13483 (N_13483,N_11450,N_9818);
or U13484 (N_13484,N_10033,N_10717);
and U13485 (N_13485,N_11349,N_9625);
nor U13486 (N_13486,N_10945,N_9813);
nor U13487 (N_13487,N_10654,N_11640);
or U13488 (N_13488,N_11102,N_9170);
nor U13489 (N_13489,N_10156,N_10612);
nor U13490 (N_13490,N_9847,N_9762);
nor U13491 (N_13491,N_10402,N_10348);
xor U13492 (N_13492,N_11625,N_11220);
or U13493 (N_13493,N_10031,N_11909);
or U13494 (N_13494,N_11545,N_9371);
and U13495 (N_13495,N_11835,N_11516);
and U13496 (N_13496,N_9771,N_10622);
nand U13497 (N_13497,N_9143,N_10519);
or U13498 (N_13498,N_10875,N_11526);
nor U13499 (N_13499,N_9588,N_10356);
nand U13500 (N_13500,N_10111,N_11764);
and U13501 (N_13501,N_10270,N_10502);
nor U13502 (N_13502,N_9917,N_9731);
nand U13503 (N_13503,N_11381,N_9618);
xor U13504 (N_13504,N_11609,N_10769);
xnor U13505 (N_13505,N_11020,N_11066);
and U13506 (N_13506,N_10838,N_9629);
and U13507 (N_13507,N_9304,N_11654);
or U13508 (N_13508,N_10421,N_10299);
and U13509 (N_13509,N_10112,N_9494);
nand U13510 (N_13510,N_10730,N_9806);
or U13511 (N_13511,N_10412,N_10752);
and U13512 (N_13512,N_11003,N_9747);
nor U13513 (N_13513,N_9769,N_11888);
nand U13514 (N_13514,N_11325,N_9630);
nor U13515 (N_13515,N_9439,N_10795);
nor U13516 (N_13516,N_11543,N_10221);
or U13517 (N_13517,N_10021,N_10995);
or U13518 (N_13518,N_9195,N_11684);
nor U13519 (N_13519,N_10870,N_9072);
or U13520 (N_13520,N_10353,N_9597);
or U13521 (N_13521,N_10197,N_11092);
nor U13522 (N_13522,N_11506,N_10387);
xnor U13523 (N_13523,N_11283,N_9546);
nor U13524 (N_13524,N_11565,N_10060);
xnor U13525 (N_13525,N_10508,N_11645);
or U13526 (N_13526,N_10291,N_9894);
nand U13527 (N_13527,N_10442,N_9411);
xor U13528 (N_13528,N_11047,N_10361);
nand U13529 (N_13529,N_9947,N_11973);
nor U13530 (N_13530,N_11614,N_9346);
nand U13531 (N_13531,N_11533,N_9506);
and U13532 (N_13532,N_10947,N_11188);
nand U13533 (N_13533,N_9679,N_11136);
nor U13534 (N_13534,N_11194,N_9380);
and U13535 (N_13535,N_10127,N_9282);
and U13536 (N_13536,N_9246,N_9490);
or U13537 (N_13537,N_9269,N_10604);
nand U13538 (N_13538,N_11195,N_9944);
xor U13539 (N_13539,N_10304,N_11006);
or U13540 (N_13540,N_9559,N_11175);
nor U13541 (N_13541,N_11740,N_10245);
nand U13542 (N_13542,N_11508,N_9425);
nand U13543 (N_13543,N_11249,N_10036);
and U13544 (N_13544,N_9237,N_11820);
xnor U13545 (N_13545,N_9926,N_11011);
and U13546 (N_13546,N_9971,N_11275);
nor U13547 (N_13547,N_10237,N_11458);
or U13548 (N_13548,N_9896,N_10961);
nand U13549 (N_13549,N_9294,N_9220);
and U13550 (N_13550,N_11344,N_10879);
nand U13551 (N_13551,N_10353,N_11240);
xnor U13552 (N_13552,N_11153,N_11985);
nand U13553 (N_13553,N_10172,N_10840);
nand U13554 (N_13554,N_9177,N_10975);
nand U13555 (N_13555,N_10807,N_9829);
nor U13556 (N_13556,N_11965,N_11052);
or U13557 (N_13557,N_10688,N_11950);
or U13558 (N_13558,N_9970,N_9520);
nand U13559 (N_13559,N_9095,N_10609);
xor U13560 (N_13560,N_11729,N_11191);
nor U13561 (N_13561,N_9870,N_9949);
or U13562 (N_13562,N_11879,N_10088);
nor U13563 (N_13563,N_9970,N_11561);
nand U13564 (N_13564,N_9938,N_10690);
nand U13565 (N_13565,N_10389,N_9627);
and U13566 (N_13566,N_11886,N_10610);
or U13567 (N_13567,N_9122,N_10470);
nand U13568 (N_13568,N_9213,N_9742);
nor U13569 (N_13569,N_9720,N_9147);
nand U13570 (N_13570,N_9865,N_10357);
or U13571 (N_13571,N_11756,N_9758);
and U13572 (N_13572,N_9342,N_10794);
nor U13573 (N_13573,N_10039,N_11171);
nor U13574 (N_13574,N_9394,N_11296);
or U13575 (N_13575,N_11386,N_11937);
and U13576 (N_13576,N_9337,N_10450);
or U13577 (N_13577,N_10857,N_11878);
nor U13578 (N_13578,N_11878,N_11396);
nor U13579 (N_13579,N_9791,N_10284);
nand U13580 (N_13580,N_11447,N_11340);
or U13581 (N_13581,N_10687,N_9044);
nand U13582 (N_13582,N_11458,N_11437);
or U13583 (N_13583,N_9556,N_9789);
or U13584 (N_13584,N_10114,N_9749);
and U13585 (N_13585,N_9394,N_11549);
nor U13586 (N_13586,N_9464,N_9628);
or U13587 (N_13587,N_10579,N_11057);
nand U13588 (N_13588,N_11939,N_9677);
and U13589 (N_13589,N_11235,N_11586);
and U13590 (N_13590,N_10872,N_9651);
nand U13591 (N_13591,N_9528,N_10297);
or U13592 (N_13592,N_10143,N_11334);
nand U13593 (N_13593,N_10539,N_10345);
nor U13594 (N_13594,N_10342,N_11232);
nand U13595 (N_13595,N_9335,N_9393);
or U13596 (N_13596,N_11859,N_9144);
nand U13597 (N_13597,N_9358,N_9433);
and U13598 (N_13598,N_11141,N_11812);
xnor U13599 (N_13599,N_9497,N_10944);
and U13600 (N_13600,N_10169,N_11661);
and U13601 (N_13601,N_10361,N_10898);
nand U13602 (N_13602,N_9915,N_9121);
or U13603 (N_13603,N_11929,N_11146);
and U13604 (N_13604,N_11613,N_9647);
or U13605 (N_13605,N_11230,N_9883);
nor U13606 (N_13606,N_11130,N_11056);
or U13607 (N_13607,N_9989,N_9881);
nor U13608 (N_13608,N_11114,N_10122);
or U13609 (N_13609,N_9955,N_11663);
or U13610 (N_13610,N_11541,N_9765);
nor U13611 (N_13611,N_10837,N_10511);
nor U13612 (N_13612,N_10755,N_10083);
and U13613 (N_13613,N_10087,N_11373);
xor U13614 (N_13614,N_9967,N_10556);
nand U13615 (N_13615,N_10169,N_9623);
and U13616 (N_13616,N_9805,N_10203);
and U13617 (N_13617,N_10473,N_10668);
or U13618 (N_13618,N_10522,N_11816);
or U13619 (N_13619,N_9885,N_9541);
nand U13620 (N_13620,N_9038,N_9681);
xor U13621 (N_13621,N_10089,N_9533);
or U13622 (N_13622,N_11709,N_9378);
xnor U13623 (N_13623,N_11071,N_11126);
nand U13624 (N_13624,N_9261,N_9251);
xor U13625 (N_13625,N_11895,N_10000);
or U13626 (N_13626,N_9837,N_9703);
or U13627 (N_13627,N_10647,N_11475);
and U13628 (N_13628,N_11781,N_11176);
nor U13629 (N_13629,N_10823,N_9192);
nor U13630 (N_13630,N_11711,N_9824);
and U13631 (N_13631,N_11668,N_9606);
or U13632 (N_13632,N_10369,N_11712);
nor U13633 (N_13633,N_10660,N_11861);
and U13634 (N_13634,N_9267,N_10828);
nand U13635 (N_13635,N_11374,N_9228);
and U13636 (N_13636,N_9838,N_10023);
nor U13637 (N_13637,N_10834,N_9473);
nand U13638 (N_13638,N_9505,N_11172);
nor U13639 (N_13639,N_10496,N_10689);
xor U13640 (N_13640,N_9251,N_11928);
nand U13641 (N_13641,N_9947,N_9333);
nand U13642 (N_13642,N_11294,N_10953);
nor U13643 (N_13643,N_9647,N_11470);
or U13644 (N_13644,N_9984,N_11546);
nor U13645 (N_13645,N_9321,N_11898);
and U13646 (N_13646,N_9823,N_10967);
and U13647 (N_13647,N_9347,N_10060);
and U13648 (N_13648,N_10978,N_10338);
or U13649 (N_13649,N_9821,N_9636);
and U13650 (N_13650,N_9140,N_11978);
xnor U13651 (N_13651,N_9010,N_11079);
nand U13652 (N_13652,N_10765,N_10256);
or U13653 (N_13653,N_9178,N_9179);
and U13654 (N_13654,N_9782,N_11894);
nand U13655 (N_13655,N_10488,N_9635);
or U13656 (N_13656,N_9459,N_9839);
nand U13657 (N_13657,N_11636,N_9386);
or U13658 (N_13658,N_10215,N_9808);
xor U13659 (N_13659,N_10770,N_9332);
nor U13660 (N_13660,N_10985,N_9799);
nor U13661 (N_13661,N_10062,N_10196);
nand U13662 (N_13662,N_9669,N_11322);
or U13663 (N_13663,N_9551,N_11606);
nor U13664 (N_13664,N_11765,N_9304);
nor U13665 (N_13665,N_11998,N_10212);
nor U13666 (N_13666,N_9538,N_11729);
or U13667 (N_13667,N_9674,N_11223);
nand U13668 (N_13668,N_10995,N_10827);
or U13669 (N_13669,N_9767,N_11184);
and U13670 (N_13670,N_11087,N_11825);
or U13671 (N_13671,N_11154,N_11347);
nor U13672 (N_13672,N_10996,N_9143);
and U13673 (N_13673,N_9626,N_10541);
or U13674 (N_13674,N_11192,N_9252);
nand U13675 (N_13675,N_9747,N_9281);
or U13676 (N_13676,N_11307,N_10790);
and U13677 (N_13677,N_10488,N_9399);
or U13678 (N_13678,N_9354,N_9034);
or U13679 (N_13679,N_11451,N_10009);
nand U13680 (N_13680,N_9383,N_11632);
nand U13681 (N_13681,N_11507,N_10845);
and U13682 (N_13682,N_11531,N_9298);
and U13683 (N_13683,N_11505,N_9024);
nor U13684 (N_13684,N_11310,N_11183);
or U13685 (N_13685,N_11328,N_10099);
nor U13686 (N_13686,N_10199,N_11833);
nor U13687 (N_13687,N_10170,N_10431);
and U13688 (N_13688,N_9089,N_10529);
or U13689 (N_13689,N_11754,N_10245);
nand U13690 (N_13690,N_11167,N_9163);
or U13691 (N_13691,N_9078,N_11707);
nor U13692 (N_13692,N_10663,N_9855);
or U13693 (N_13693,N_11734,N_9722);
nor U13694 (N_13694,N_10818,N_9862);
nor U13695 (N_13695,N_9422,N_9165);
xnor U13696 (N_13696,N_11101,N_10760);
or U13697 (N_13697,N_10038,N_9197);
nor U13698 (N_13698,N_11257,N_10221);
nand U13699 (N_13699,N_11707,N_10050);
nor U13700 (N_13700,N_11758,N_11116);
nand U13701 (N_13701,N_9010,N_10331);
nand U13702 (N_13702,N_10145,N_11506);
nor U13703 (N_13703,N_11338,N_9329);
nor U13704 (N_13704,N_10894,N_9735);
nand U13705 (N_13705,N_9415,N_10342);
nor U13706 (N_13706,N_11737,N_9655);
and U13707 (N_13707,N_9328,N_9577);
nand U13708 (N_13708,N_9864,N_11104);
nand U13709 (N_13709,N_11156,N_11778);
or U13710 (N_13710,N_11235,N_10677);
and U13711 (N_13711,N_11702,N_11310);
xnor U13712 (N_13712,N_10089,N_9712);
nand U13713 (N_13713,N_11314,N_11500);
or U13714 (N_13714,N_9375,N_9949);
and U13715 (N_13715,N_9737,N_10136);
nor U13716 (N_13716,N_9706,N_9737);
and U13717 (N_13717,N_10130,N_11387);
xnor U13718 (N_13718,N_10801,N_11737);
and U13719 (N_13719,N_9481,N_9085);
and U13720 (N_13720,N_10220,N_11457);
nor U13721 (N_13721,N_10689,N_9126);
and U13722 (N_13722,N_9567,N_9339);
nand U13723 (N_13723,N_10902,N_11403);
and U13724 (N_13724,N_9157,N_10545);
and U13725 (N_13725,N_11381,N_9854);
and U13726 (N_13726,N_10997,N_11777);
and U13727 (N_13727,N_11057,N_9349);
xnor U13728 (N_13728,N_11979,N_11953);
nor U13729 (N_13729,N_10456,N_9360);
nand U13730 (N_13730,N_9408,N_10616);
nand U13731 (N_13731,N_9167,N_10048);
xor U13732 (N_13732,N_11098,N_11550);
xnor U13733 (N_13733,N_10845,N_9753);
or U13734 (N_13734,N_9732,N_11856);
nor U13735 (N_13735,N_9536,N_10356);
nand U13736 (N_13736,N_11729,N_9974);
and U13737 (N_13737,N_9492,N_10893);
nand U13738 (N_13738,N_11680,N_9953);
or U13739 (N_13739,N_10990,N_11880);
or U13740 (N_13740,N_10602,N_10915);
nand U13741 (N_13741,N_9482,N_10270);
xor U13742 (N_13742,N_11883,N_10266);
nand U13743 (N_13743,N_11677,N_9598);
or U13744 (N_13744,N_10099,N_10361);
or U13745 (N_13745,N_10314,N_11603);
or U13746 (N_13746,N_11903,N_9230);
and U13747 (N_13747,N_10073,N_9487);
or U13748 (N_13748,N_11185,N_9873);
or U13749 (N_13749,N_10776,N_10156);
or U13750 (N_13750,N_9654,N_11061);
or U13751 (N_13751,N_9492,N_10645);
nand U13752 (N_13752,N_9750,N_9660);
nand U13753 (N_13753,N_11310,N_11505);
and U13754 (N_13754,N_10844,N_9569);
xnor U13755 (N_13755,N_11890,N_9020);
or U13756 (N_13756,N_11947,N_9055);
nor U13757 (N_13757,N_11719,N_9384);
nor U13758 (N_13758,N_9927,N_10512);
or U13759 (N_13759,N_11509,N_11539);
nor U13760 (N_13760,N_10211,N_9861);
and U13761 (N_13761,N_9796,N_10529);
nand U13762 (N_13762,N_11284,N_10229);
or U13763 (N_13763,N_11224,N_10810);
nor U13764 (N_13764,N_10573,N_10398);
nand U13765 (N_13765,N_11950,N_9312);
and U13766 (N_13766,N_11632,N_11678);
and U13767 (N_13767,N_11241,N_11799);
and U13768 (N_13768,N_9288,N_9654);
nand U13769 (N_13769,N_11071,N_9552);
xnor U13770 (N_13770,N_11866,N_9432);
xnor U13771 (N_13771,N_10671,N_11382);
nor U13772 (N_13772,N_11830,N_11853);
xor U13773 (N_13773,N_9209,N_9385);
xor U13774 (N_13774,N_9037,N_10770);
xnor U13775 (N_13775,N_10756,N_11577);
and U13776 (N_13776,N_9601,N_10808);
nor U13777 (N_13777,N_10697,N_9884);
nor U13778 (N_13778,N_9283,N_10163);
and U13779 (N_13779,N_9372,N_11948);
or U13780 (N_13780,N_9763,N_10370);
nand U13781 (N_13781,N_11612,N_11788);
or U13782 (N_13782,N_9644,N_11082);
or U13783 (N_13783,N_9238,N_9227);
and U13784 (N_13784,N_11521,N_10349);
and U13785 (N_13785,N_10243,N_10955);
nand U13786 (N_13786,N_9792,N_11071);
or U13787 (N_13787,N_10040,N_11593);
or U13788 (N_13788,N_11937,N_11057);
nand U13789 (N_13789,N_9306,N_11553);
or U13790 (N_13790,N_11211,N_11413);
nor U13791 (N_13791,N_9074,N_10459);
and U13792 (N_13792,N_10272,N_11705);
or U13793 (N_13793,N_10668,N_10152);
nand U13794 (N_13794,N_10304,N_9218);
or U13795 (N_13795,N_10149,N_11821);
and U13796 (N_13796,N_11511,N_10542);
nor U13797 (N_13797,N_11321,N_10299);
nand U13798 (N_13798,N_10774,N_11096);
or U13799 (N_13799,N_11773,N_9930);
and U13800 (N_13800,N_10908,N_11609);
nand U13801 (N_13801,N_10845,N_9212);
or U13802 (N_13802,N_11417,N_11664);
and U13803 (N_13803,N_9053,N_9564);
nor U13804 (N_13804,N_11414,N_9516);
or U13805 (N_13805,N_9687,N_10730);
and U13806 (N_13806,N_11207,N_10499);
or U13807 (N_13807,N_9905,N_9365);
xnor U13808 (N_13808,N_11697,N_10674);
nand U13809 (N_13809,N_11450,N_9924);
or U13810 (N_13810,N_11587,N_9399);
nand U13811 (N_13811,N_11203,N_10095);
nor U13812 (N_13812,N_9718,N_9609);
or U13813 (N_13813,N_10473,N_10994);
nor U13814 (N_13814,N_9598,N_10412);
or U13815 (N_13815,N_9932,N_9090);
or U13816 (N_13816,N_9403,N_11088);
nand U13817 (N_13817,N_10494,N_10898);
nor U13818 (N_13818,N_10511,N_9097);
or U13819 (N_13819,N_10288,N_9272);
or U13820 (N_13820,N_9066,N_10133);
nor U13821 (N_13821,N_9325,N_10774);
xor U13822 (N_13822,N_10583,N_9375);
nor U13823 (N_13823,N_10911,N_10465);
and U13824 (N_13824,N_11692,N_11161);
nand U13825 (N_13825,N_11234,N_11409);
xor U13826 (N_13826,N_9123,N_9968);
nor U13827 (N_13827,N_9468,N_11939);
or U13828 (N_13828,N_9539,N_9887);
or U13829 (N_13829,N_10826,N_9088);
and U13830 (N_13830,N_11852,N_11418);
or U13831 (N_13831,N_9199,N_9781);
or U13832 (N_13832,N_11538,N_9421);
nand U13833 (N_13833,N_9876,N_10986);
nand U13834 (N_13834,N_11894,N_9112);
or U13835 (N_13835,N_9584,N_10508);
nand U13836 (N_13836,N_9010,N_9054);
nor U13837 (N_13837,N_10585,N_10691);
nor U13838 (N_13838,N_10370,N_11341);
nand U13839 (N_13839,N_9329,N_11325);
nand U13840 (N_13840,N_11896,N_9523);
or U13841 (N_13841,N_10504,N_11927);
or U13842 (N_13842,N_10343,N_10635);
xor U13843 (N_13843,N_9581,N_10756);
nor U13844 (N_13844,N_11399,N_11032);
or U13845 (N_13845,N_10805,N_10576);
or U13846 (N_13846,N_10850,N_10240);
or U13847 (N_13847,N_10960,N_9862);
nor U13848 (N_13848,N_9074,N_10685);
nand U13849 (N_13849,N_10565,N_10459);
nor U13850 (N_13850,N_9512,N_11729);
or U13851 (N_13851,N_10486,N_11222);
and U13852 (N_13852,N_10449,N_9591);
nor U13853 (N_13853,N_9784,N_9583);
or U13854 (N_13854,N_10778,N_9128);
nor U13855 (N_13855,N_9710,N_11486);
nor U13856 (N_13856,N_9262,N_11410);
nand U13857 (N_13857,N_10332,N_11278);
or U13858 (N_13858,N_10916,N_11796);
nand U13859 (N_13859,N_11093,N_11199);
and U13860 (N_13860,N_10227,N_11029);
xor U13861 (N_13861,N_10303,N_10244);
nor U13862 (N_13862,N_11785,N_10461);
and U13863 (N_13863,N_9292,N_9914);
nand U13864 (N_13864,N_10477,N_11439);
and U13865 (N_13865,N_10827,N_9667);
nand U13866 (N_13866,N_10324,N_9596);
or U13867 (N_13867,N_9709,N_10812);
nor U13868 (N_13868,N_11494,N_10348);
nor U13869 (N_13869,N_9204,N_11393);
and U13870 (N_13870,N_10049,N_9604);
nand U13871 (N_13871,N_9952,N_11884);
nand U13872 (N_13872,N_11988,N_9095);
or U13873 (N_13873,N_9231,N_11588);
or U13874 (N_13874,N_11512,N_11106);
nand U13875 (N_13875,N_10326,N_10283);
or U13876 (N_13876,N_10928,N_9609);
nand U13877 (N_13877,N_10624,N_9933);
nor U13878 (N_13878,N_10670,N_11927);
nand U13879 (N_13879,N_11130,N_11729);
and U13880 (N_13880,N_11456,N_11218);
nor U13881 (N_13881,N_11162,N_10667);
or U13882 (N_13882,N_10726,N_10160);
nand U13883 (N_13883,N_10658,N_9570);
or U13884 (N_13884,N_9690,N_9981);
nand U13885 (N_13885,N_10588,N_9892);
nand U13886 (N_13886,N_10690,N_11636);
nor U13887 (N_13887,N_9292,N_10763);
or U13888 (N_13888,N_10923,N_10212);
nor U13889 (N_13889,N_9991,N_10000);
and U13890 (N_13890,N_11853,N_9840);
or U13891 (N_13891,N_11134,N_9232);
nor U13892 (N_13892,N_9630,N_9124);
or U13893 (N_13893,N_10926,N_11080);
nand U13894 (N_13894,N_9903,N_10446);
or U13895 (N_13895,N_11708,N_10745);
nor U13896 (N_13896,N_10666,N_9967);
nor U13897 (N_13897,N_9110,N_9309);
nand U13898 (N_13898,N_10276,N_10601);
xor U13899 (N_13899,N_9650,N_11245);
nand U13900 (N_13900,N_9387,N_9936);
or U13901 (N_13901,N_10980,N_10038);
nor U13902 (N_13902,N_10562,N_10034);
and U13903 (N_13903,N_11109,N_10864);
xnor U13904 (N_13904,N_11389,N_10477);
or U13905 (N_13905,N_10539,N_10742);
and U13906 (N_13906,N_10306,N_9891);
nor U13907 (N_13907,N_11080,N_9629);
and U13908 (N_13908,N_9925,N_11929);
nor U13909 (N_13909,N_9460,N_9826);
or U13910 (N_13910,N_11052,N_10511);
nand U13911 (N_13911,N_10591,N_10823);
or U13912 (N_13912,N_11939,N_9412);
nor U13913 (N_13913,N_10166,N_10936);
nor U13914 (N_13914,N_10530,N_9020);
and U13915 (N_13915,N_9879,N_11275);
xnor U13916 (N_13916,N_9674,N_11520);
nand U13917 (N_13917,N_10206,N_9528);
nand U13918 (N_13918,N_10006,N_9640);
or U13919 (N_13919,N_11364,N_9807);
and U13920 (N_13920,N_9938,N_9441);
nand U13921 (N_13921,N_9901,N_9290);
and U13922 (N_13922,N_11147,N_11396);
xor U13923 (N_13923,N_11990,N_9913);
nor U13924 (N_13924,N_9611,N_9944);
and U13925 (N_13925,N_9012,N_9008);
or U13926 (N_13926,N_10072,N_9008);
nand U13927 (N_13927,N_9440,N_10985);
or U13928 (N_13928,N_11631,N_11636);
and U13929 (N_13929,N_10615,N_10642);
nor U13930 (N_13930,N_9400,N_9175);
nor U13931 (N_13931,N_9019,N_11104);
nand U13932 (N_13932,N_10581,N_11093);
nor U13933 (N_13933,N_11100,N_10978);
xnor U13934 (N_13934,N_11155,N_11305);
and U13935 (N_13935,N_11326,N_10345);
nand U13936 (N_13936,N_11753,N_9113);
nand U13937 (N_13937,N_10083,N_9491);
and U13938 (N_13938,N_9665,N_10877);
and U13939 (N_13939,N_9989,N_9029);
or U13940 (N_13940,N_11185,N_9355);
and U13941 (N_13941,N_11350,N_9187);
nor U13942 (N_13942,N_9935,N_10230);
and U13943 (N_13943,N_9860,N_10394);
nand U13944 (N_13944,N_11390,N_10804);
nand U13945 (N_13945,N_9373,N_10047);
and U13946 (N_13946,N_9696,N_10334);
or U13947 (N_13947,N_11252,N_11886);
and U13948 (N_13948,N_11661,N_10004);
nor U13949 (N_13949,N_10833,N_10965);
and U13950 (N_13950,N_11895,N_10233);
and U13951 (N_13951,N_10713,N_11544);
and U13952 (N_13952,N_9352,N_10169);
nor U13953 (N_13953,N_11590,N_9468);
or U13954 (N_13954,N_11010,N_9205);
and U13955 (N_13955,N_9109,N_9546);
nand U13956 (N_13956,N_9579,N_9178);
or U13957 (N_13957,N_9758,N_10235);
nor U13958 (N_13958,N_9881,N_9208);
and U13959 (N_13959,N_9428,N_9273);
nor U13960 (N_13960,N_10308,N_10778);
xnor U13961 (N_13961,N_9722,N_11170);
and U13962 (N_13962,N_9737,N_10409);
nand U13963 (N_13963,N_9362,N_11712);
or U13964 (N_13964,N_11338,N_9935);
nand U13965 (N_13965,N_10182,N_9275);
nor U13966 (N_13966,N_9874,N_11630);
and U13967 (N_13967,N_9650,N_10814);
nor U13968 (N_13968,N_10204,N_9765);
and U13969 (N_13969,N_9625,N_10873);
nand U13970 (N_13970,N_10103,N_10018);
or U13971 (N_13971,N_9659,N_9357);
nor U13972 (N_13972,N_10995,N_9706);
nor U13973 (N_13973,N_11469,N_11681);
xor U13974 (N_13974,N_10251,N_9397);
nand U13975 (N_13975,N_11608,N_9327);
nor U13976 (N_13976,N_11887,N_10272);
or U13977 (N_13977,N_10614,N_11205);
xor U13978 (N_13978,N_9219,N_11373);
nor U13979 (N_13979,N_10558,N_10263);
xnor U13980 (N_13980,N_9248,N_10955);
nand U13981 (N_13981,N_10224,N_10106);
and U13982 (N_13982,N_9285,N_11410);
xnor U13983 (N_13983,N_9331,N_10326);
or U13984 (N_13984,N_11734,N_11533);
nand U13985 (N_13985,N_10249,N_11309);
and U13986 (N_13986,N_9604,N_11946);
xnor U13987 (N_13987,N_10681,N_10427);
xor U13988 (N_13988,N_11333,N_10448);
and U13989 (N_13989,N_9191,N_9793);
and U13990 (N_13990,N_11340,N_9080);
or U13991 (N_13991,N_9542,N_9710);
nor U13992 (N_13992,N_11821,N_11452);
or U13993 (N_13993,N_9548,N_10343);
xnor U13994 (N_13994,N_11009,N_10028);
nor U13995 (N_13995,N_9125,N_10208);
or U13996 (N_13996,N_11857,N_9927);
nor U13997 (N_13997,N_11515,N_10643);
and U13998 (N_13998,N_11807,N_10324);
nand U13999 (N_13999,N_10766,N_10307);
or U14000 (N_14000,N_10850,N_9562);
nand U14001 (N_14001,N_10961,N_9639);
nor U14002 (N_14002,N_9827,N_11482);
nor U14003 (N_14003,N_9930,N_10184);
and U14004 (N_14004,N_9024,N_10383);
and U14005 (N_14005,N_11567,N_9103);
or U14006 (N_14006,N_9244,N_10697);
xnor U14007 (N_14007,N_10043,N_9194);
nor U14008 (N_14008,N_10547,N_11812);
or U14009 (N_14009,N_10022,N_9292);
nor U14010 (N_14010,N_11916,N_10261);
or U14011 (N_14011,N_10807,N_11845);
and U14012 (N_14012,N_9724,N_11288);
nor U14013 (N_14013,N_9772,N_10311);
or U14014 (N_14014,N_11154,N_11247);
xnor U14015 (N_14015,N_11204,N_9434);
nand U14016 (N_14016,N_10559,N_10116);
nor U14017 (N_14017,N_11192,N_10233);
xor U14018 (N_14018,N_9300,N_9339);
nand U14019 (N_14019,N_10278,N_11319);
and U14020 (N_14020,N_9657,N_10624);
and U14021 (N_14021,N_10195,N_10601);
xor U14022 (N_14022,N_9145,N_10049);
and U14023 (N_14023,N_9243,N_11662);
or U14024 (N_14024,N_11277,N_10408);
or U14025 (N_14025,N_9962,N_10993);
nor U14026 (N_14026,N_9102,N_10648);
and U14027 (N_14027,N_10110,N_10297);
and U14028 (N_14028,N_10827,N_9834);
xnor U14029 (N_14029,N_11608,N_9924);
nor U14030 (N_14030,N_9114,N_9217);
nor U14031 (N_14031,N_9436,N_10616);
and U14032 (N_14032,N_11044,N_11824);
nand U14033 (N_14033,N_9955,N_10630);
and U14034 (N_14034,N_9933,N_11260);
and U14035 (N_14035,N_10714,N_9669);
nor U14036 (N_14036,N_10528,N_10141);
and U14037 (N_14037,N_10310,N_10652);
xnor U14038 (N_14038,N_9230,N_9833);
xnor U14039 (N_14039,N_9280,N_9597);
nand U14040 (N_14040,N_10529,N_9829);
xnor U14041 (N_14041,N_10063,N_9285);
nor U14042 (N_14042,N_11743,N_11441);
and U14043 (N_14043,N_9311,N_10051);
nor U14044 (N_14044,N_10651,N_10170);
nand U14045 (N_14045,N_10777,N_9050);
nor U14046 (N_14046,N_11319,N_10038);
nand U14047 (N_14047,N_10114,N_11752);
or U14048 (N_14048,N_11894,N_10872);
nand U14049 (N_14049,N_11541,N_10297);
nor U14050 (N_14050,N_10398,N_10854);
nand U14051 (N_14051,N_10398,N_9921);
and U14052 (N_14052,N_9909,N_9975);
nor U14053 (N_14053,N_10519,N_9265);
nand U14054 (N_14054,N_10278,N_11805);
nand U14055 (N_14055,N_10485,N_11587);
nand U14056 (N_14056,N_10896,N_11804);
and U14057 (N_14057,N_11871,N_9597);
or U14058 (N_14058,N_11843,N_11422);
xnor U14059 (N_14059,N_9757,N_10973);
nor U14060 (N_14060,N_10548,N_10976);
or U14061 (N_14061,N_11656,N_10389);
and U14062 (N_14062,N_11745,N_10898);
nor U14063 (N_14063,N_10497,N_10323);
and U14064 (N_14064,N_11702,N_11118);
and U14065 (N_14065,N_9395,N_9115);
nand U14066 (N_14066,N_9770,N_11767);
and U14067 (N_14067,N_9884,N_11343);
nor U14068 (N_14068,N_11689,N_11652);
nand U14069 (N_14069,N_10030,N_11541);
or U14070 (N_14070,N_11890,N_9292);
nor U14071 (N_14071,N_11203,N_11941);
and U14072 (N_14072,N_10317,N_9173);
or U14073 (N_14073,N_9120,N_10217);
nand U14074 (N_14074,N_10357,N_11784);
and U14075 (N_14075,N_9702,N_11407);
nand U14076 (N_14076,N_11863,N_10541);
or U14077 (N_14077,N_10530,N_9317);
nor U14078 (N_14078,N_9024,N_11994);
or U14079 (N_14079,N_10134,N_9797);
or U14080 (N_14080,N_11878,N_11110);
nand U14081 (N_14081,N_9612,N_11006);
and U14082 (N_14082,N_11790,N_10130);
and U14083 (N_14083,N_10604,N_10086);
or U14084 (N_14084,N_10896,N_11249);
nor U14085 (N_14085,N_10117,N_10750);
nor U14086 (N_14086,N_11229,N_10527);
nand U14087 (N_14087,N_9112,N_10228);
and U14088 (N_14088,N_10909,N_10552);
or U14089 (N_14089,N_9182,N_11483);
nand U14090 (N_14090,N_10512,N_11543);
nor U14091 (N_14091,N_11871,N_10287);
nor U14092 (N_14092,N_11421,N_9591);
nor U14093 (N_14093,N_11973,N_9120);
nand U14094 (N_14094,N_10720,N_11462);
nor U14095 (N_14095,N_10957,N_9842);
nand U14096 (N_14096,N_11122,N_11017);
xor U14097 (N_14097,N_9177,N_11636);
nand U14098 (N_14098,N_10849,N_9230);
or U14099 (N_14099,N_10205,N_10257);
nor U14100 (N_14100,N_11870,N_9782);
nand U14101 (N_14101,N_10722,N_11332);
and U14102 (N_14102,N_10739,N_10893);
and U14103 (N_14103,N_11567,N_10675);
or U14104 (N_14104,N_10903,N_11980);
nor U14105 (N_14105,N_9541,N_9108);
and U14106 (N_14106,N_11633,N_9264);
nand U14107 (N_14107,N_11528,N_10039);
nand U14108 (N_14108,N_9539,N_9001);
and U14109 (N_14109,N_10971,N_9879);
and U14110 (N_14110,N_11830,N_9481);
xor U14111 (N_14111,N_11157,N_10891);
nor U14112 (N_14112,N_10641,N_11001);
nand U14113 (N_14113,N_11648,N_10333);
or U14114 (N_14114,N_11029,N_11458);
nor U14115 (N_14115,N_10660,N_9495);
nand U14116 (N_14116,N_11661,N_10084);
nor U14117 (N_14117,N_10880,N_9435);
nor U14118 (N_14118,N_11206,N_10720);
and U14119 (N_14119,N_10051,N_10704);
and U14120 (N_14120,N_11672,N_10516);
nor U14121 (N_14121,N_9845,N_11284);
or U14122 (N_14122,N_10609,N_9090);
nand U14123 (N_14123,N_11528,N_10642);
or U14124 (N_14124,N_10651,N_11679);
or U14125 (N_14125,N_11164,N_9027);
or U14126 (N_14126,N_11021,N_11826);
or U14127 (N_14127,N_9096,N_10695);
xor U14128 (N_14128,N_10621,N_11915);
nand U14129 (N_14129,N_11347,N_11014);
xor U14130 (N_14130,N_9071,N_11002);
and U14131 (N_14131,N_9070,N_10364);
nor U14132 (N_14132,N_10272,N_11618);
nor U14133 (N_14133,N_9290,N_9061);
nor U14134 (N_14134,N_11968,N_9438);
nand U14135 (N_14135,N_11381,N_10361);
nand U14136 (N_14136,N_11140,N_11132);
nor U14137 (N_14137,N_11937,N_11934);
nand U14138 (N_14138,N_9154,N_10436);
nand U14139 (N_14139,N_9182,N_10299);
nor U14140 (N_14140,N_11705,N_11213);
nor U14141 (N_14141,N_10173,N_9134);
xor U14142 (N_14142,N_9510,N_9160);
nor U14143 (N_14143,N_11276,N_10571);
or U14144 (N_14144,N_11544,N_9368);
nand U14145 (N_14145,N_11148,N_9288);
and U14146 (N_14146,N_10813,N_9705);
nand U14147 (N_14147,N_9112,N_9970);
and U14148 (N_14148,N_9121,N_11797);
nand U14149 (N_14149,N_10753,N_11481);
or U14150 (N_14150,N_11229,N_11592);
and U14151 (N_14151,N_11656,N_9357);
nand U14152 (N_14152,N_11344,N_9711);
nand U14153 (N_14153,N_11190,N_10685);
or U14154 (N_14154,N_10571,N_10533);
or U14155 (N_14155,N_10291,N_9427);
nor U14156 (N_14156,N_11249,N_9112);
or U14157 (N_14157,N_10939,N_9281);
and U14158 (N_14158,N_9236,N_10950);
or U14159 (N_14159,N_9214,N_10691);
or U14160 (N_14160,N_9462,N_10152);
or U14161 (N_14161,N_11507,N_11672);
nand U14162 (N_14162,N_10259,N_10268);
and U14163 (N_14163,N_10641,N_10202);
or U14164 (N_14164,N_9746,N_11730);
xnor U14165 (N_14165,N_10229,N_10795);
xnor U14166 (N_14166,N_11786,N_10929);
or U14167 (N_14167,N_10319,N_10798);
and U14168 (N_14168,N_10774,N_9173);
and U14169 (N_14169,N_9075,N_9167);
nor U14170 (N_14170,N_9966,N_10752);
or U14171 (N_14171,N_10409,N_11539);
xor U14172 (N_14172,N_10367,N_10717);
xnor U14173 (N_14173,N_9468,N_11134);
nor U14174 (N_14174,N_10668,N_9001);
or U14175 (N_14175,N_10514,N_10272);
nand U14176 (N_14176,N_10130,N_10230);
and U14177 (N_14177,N_10567,N_11734);
nand U14178 (N_14178,N_9029,N_10073);
and U14179 (N_14179,N_11257,N_11994);
and U14180 (N_14180,N_10462,N_10899);
nor U14181 (N_14181,N_10565,N_10429);
and U14182 (N_14182,N_9942,N_11232);
and U14183 (N_14183,N_11884,N_9674);
and U14184 (N_14184,N_11721,N_11805);
nor U14185 (N_14185,N_11085,N_11486);
or U14186 (N_14186,N_11820,N_10678);
nand U14187 (N_14187,N_10103,N_11453);
or U14188 (N_14188,N_9226,N_11670);
nand U14189 (N_14189,N_9166,N_10144);
nand U14190 (N_14190,N_11469,N_9833);
xnor U14191 (N_14191,N_11923,N_11572);
nand U14192 (N_14192,N_9971,N_10866);
nor U14193 (N_14193,N_9399,N_9695);
nand U14194 (N_14194,N_9502,N_9022);
or U14195 (N_14195,N_9618,N_9481);
or U14196 (N_14196,N_9238,N_9711);
and U14197 (N_14197,N_11346,N_9167);
and U14198 (N_14198,N_10855,N_9741);
nand U14199 (N_14199,N_10059,N_11057);
or U14200 (N_14200,N_11940,N_9808);
nor U14201 (N_14201,N_11887,N_9898);
xor U14202 (N_14202,N_11297,N_11255);
or U14203 (N_14203,N_9192,N_10315);
nor U14204 (N_14204,N_11362,N_9839);
nand U14205 (N_14205,N_9141,N_11354);
nand U14206 (N_14206,N_9512,N_10937);
and U14207 (N_14207,N_10853,N_11819);
or U14208 (N_14208,N_10918,N_11058);
nand U14209 (N_14209,N_9611,N_10581);
or U14210 (N_14210,N_10752,N_10291);
and U14211 (N_14211,N_10938,N_9581);
nor U14212 (N_14212,N_9037,N_10571);
or U14213 (N_14213,N_10344,N_9929);
nor U14214 (N_14214,N_10776,N_9696);
and U14215 (N_14215,N_11635,N_9351);
nand U14216 (N_14216,N_11991,N_9963);
and U14217 (N_14217,N_11692,N_11941);
or U14218 (N_14218,N_9960,N_9246);
and U14219 (N_14219,N_9559,N_9790);
and U14220 (N_14220,N_9067,N_9872);
nor U14221 (N_14221,N_11816,N_10538);
and U14222 (N_14222,N_10038,N_9320);
nor U14223 (N_14223,N_11016,N_10775);
nand U14224 (N_14224,N_10740,N_9749);
or U14225 (N_14225,N_9208,N_10529);
and U14226 (N_14226,N_9483,N_10518);
nor U14227 (N_14227,N_10026,N_10706);
nor U14228 (N_14228,N_10505,N_10882);
nand U14229 (N_14229,N_11487,N_9833);
or U14230 (N_14230,N_11017,N_9527);
nand U14231 (N_14231,N_11995,N_10745);
or U14232 (N_14232,N_11600,N_11751);
or U14233 (N_14233,N_10258,N_10477);
and U14234 (N_14234,N_10284,N_9935);
or U14235 (N_14235,N_10097,N_10868);
nor U14236 (N_14236,N_10881,N_11121);
nand U14237 (N_14237,N_11763,N_11269);
nor U14238 (N_14238,N_11079,N_11323);
nor U14239 (N_14239,N_9884,N_10820);
and U14240 (N_14240,N_9727,N_11594);
or U14241 (N_14241,N_10800,N_11645);
nor U14242 (N_14242,N_9345,N_9449);
or U14243 (N_14243,N_11071,N_9083);
nor U14244 (N_14244,N_11973,N_10887);
or U14245 (N_14245,N_9402,N_9966);
or U14246 (N_14246,N_10141,N_10494);
xnor U14247 (N_14247,N_11996,N_9096);
and U14248 (N_14248,N_9640,N_10211);
nor U14249 (N_14249,N_10294,N_11524);
and U14250 (N_14250,N_10875,N_11063);
nand U14251 (N_14251,N_9386,N_10228);
nor U14252 (N_14252,N_9870,N_10406);
nand U14253 (N_14253,N_11126,N_11675);
nand U14254 (N_14254,N_9487,N_11868);
or U14255 (N_14255,N_9874,N_9177);
nor U14256 (N_14256,N_9632,N_9144);
or U14257 (N_14257,N_11145,N_11593);
or U14258 (N_14258,N_11119,N_9357);
nand U14259 (N_14259,N_10663,N_9807);
or U14260 (N_14260,N_9679,N_11585);
or U14261 (N_14261,N_9965,N_9154);
and U14262 (N_14262,N_10978,N_11873);
or U14263 (N_14263,N_11508,N_10143);
nand U14264 (N_14264,N_10621,N_9156);
nor U14265 (N_14265,N_9959,N_11531);
nor U14266 (N_14266,N_11815,N_11166);
and U14267 (N_14267,N_9076,N_11178);
nor U14268 (N_14268,N_10016,N_11431);
and U14269 (N_14269,N_10081,N_9092);
and U14270 (N_14270,N_9813,N_10406);
nand U14271 (N_14271,N_11178,N_9123);
nor U14272 (N_14272,N_11407,N_10747);
nor U14273 (N_14273,N_11575,N_11468);
or U14274 (N_14274,N_11942,N_11664);
and U14275 (N_14275,N_11806,N_11990);
nand U14276 (N_14276,N_11880,N_11059);
nor U14277 (N_14277,N_11408,N_10365);
nand U14278 (N_14278,N_9573,N_9323);
xnor U14279 (N_14279,N_10017,N_11446);
and U14280 (N_14280,N_11390,N_10690);
and U14281 (N_14281,N_9114,N_11845);
nand U14282 (N_14282,N_9317,N_9037);
nand U14283 (N_14283,N_11950,N_11096);
or U14284 (N_14284,N_11514,N_9820);
nand U14285 (N_14285,N_9915,N_10264);
and U14286 (N_14286,N_10292,N_11049);
and U14287 (N_14287,N_10694,N_9400);
or U14288 (N_14288,N_9040,N_10233);
or U14289 (N_14289,N_10848,N_9648);
xor U14290 (N_14290,N_11776,N_9537);
nand U14291 (N_14291,N_10316,N_10871);
nor U14292 (N_14292,N_9541,N_9908);
or U14293 (N_14293,N_9477,N_9929);
or U14294 (N_14294,N_10342,N_10998);
nand U14295 (N_14295,N_11252,N_11119);
or U14296 (N_14296,N_11231,N_10069);
or U14297 (N_14297,N_9979,N_11228);
and U14298 (N_14298,N_9189,N_10087);
and U14299 (N_14299,N_11267,N_9650);
and U14300 (N_14300,N_10140,N_9507);
and U14301 (N_14301,N_11595,N_9245);
nor U14302 (N_14302,N_11576,N_10599);
nand U14303 (N_14303,N_9546,N_10091);
nor U14304 (N_14304,N_9005,N_9290);
and U14305 (N_14305,N_10658,N_10193);
and U14306 (N_14306,N_11270,N_9614);
nand U14307 (N_14307,N_9971,N_11104);
xor U14308 (N_14308,N_11338,N_11150);
nand U14309 (N_14309,N_11849,N_10931);
and U14310 (N_14310,N_10498,N_10107);
nor U14311 (N_14311,N_11839,N_9607);
nand U14312 (N_14312,N_10614,N_9751);
nand U14313 (N_14313,N_10709,N_9511);
or U14314 (N_14314,N_10052,N_9464);
or U14315 (N_14315,N_9052,N_9455);
nor U14316 (N_14316,N_10715,N_10729);
or U14317 (N_14317,N_9999,N_10150);
nor U14318 (N_14318,N_9741,N_9187);
nor U14319 (N_14319,N_11776,N_11093);
and U14320 (N_14320,N_9826,N_9946);
or U14321 (N_14321,N_10299,N_9058);
or U14322 (N_14322,N_10145,N_11616);
and U14323 (N_14323,N_11771,N_10494);
or U14324 (N_14324,N_10280,N_9202);
nor U14325 (N_14325,N_10765,N_9285);
nand U14326 (N_14326,N_10581,N_11043);
or U14327 (N_14327,N_10636,N_10287);
and U14328 (N_14328,N_10548,N_11519);
nor U14329 (N_14329,N_10606,N_10290);
nor U14330 (N_14330,N_9136,N_11941);
and U14331 (N_14331,N_9922,N_10600);
and U14332 (N_14332,N_9971,N_10643);
xnor U14333 (N_14333,N_11862,N_10656);
nor U14334 (N_14334,N_10286,N_10660);
nor U14335 (N_14335,N_11235,N_10908);
and U14336 (N_14336,N_10148,N_9094);
nor U14337 (N_14337,N_9640,N_10069);
nor U14338 (N_14338,N_11576,N_11955);
or U14339 (N_14339,N_9834,N_11285);
or U14340 (N_14340,N_11702,N_11946);
nand U14341 (N_14341,N_9909,N_10743);
and U14342 (N_14342,N_10444,N_10335);
nor U14343 (N_14343,N_11214,N_11837);
nor U14344 (N_14344,N_10119,N_10634);
nor U14345 (N_14345,N_10249,N_11267);
nor U14346 (N_14346,N_9067,N_11323);
nor U14347 (N_14347,N_10993,N_11218);
or U14348 (N_14348,N_9638,N_9157);
nand U14349 (N_14349,N_10606,N_9404);
xor U14350 (N_14350,N_10614,N_10650);
and U14351 (N_14351,N_10341,N_11179);
nor U14352 (N_14352,N_9419,N_10261);
xnor U14353 (N_14353,N_9187,N_11145);
or U14354 (N_14354,N_9603,N_10287);
nor U14355 (N_14355,N_11956,N_11900);
and U14356 (N_14356,N_11370,N_11753);
nor U14357 (N_14357,N_10431,N_9435);
or U14358 (N_14358,N_9073,N_11867);
or U14359 (N_14359,N_9865,N_9558);
or U14360 (N_14360,N_10779,N_10178);
or U14361 (N_14361,N_11497,N_11626);
nor U14362 (N_14362,N_11301,N_11010);
and U14363 (N_14363,N_10955,N_9039);
nand U14364 (N_14364,N_10641,N_9040);
or U14365 (N_14365,N_11454,N_10679);
or U14366 (N_14366,N_10963,N_11174);
nor U14367 (N_14367,N_10946,N_11382);
nor U14368 (N_14368,N_11479,N_9702);
nor U14369 (N_14369,N_10411,N_10845);
or U14370 (N_14370,N_9554,N_10181);
nand U14371 (N_14371,N_10842,N_11051);
or U14372 (N_14372,N_9481,N_10040);
or U14373 (N_14373,N_10875,N_9757);
nor U14374 (N_14374,N_9048,N_10924);
nand U14375 (N_14375,N_10336,N_11404);
and U14376 (N_14376,N_9573,N_9763);
xor U14377 (N_14377,N_11612,N_9195);
or U14378 (N_14378,N_10510,N_10745);
nor U14379 (N_14379,N_9148,N_10865);
or U14380 (N_14380,N_9986,N_9900);
nor U14381 (N_14381,N_11348,N_9497);
nand U14382 (N_14382,N_10883,N_10925);
xnor U14383 (N_14383,N_11995,N_10670);
nand U14384 (N_14384,N_11466,N_10729);
or U14385 (N_14385,N_11748,N_9118);
nor U14386 (N_14386,N_11301,N_10890);
or U14387 (N_14387,N_10519,N_11355);
and U14388 (N_14388,N_10217,N_11020);
xnor U14389 (N_14389,N_10838,N_11294);
or U14390 (N_14390,N_11642,N_10064);
or U14391 (N_14391,N_10579,N_9729);
nor U14392 (N_14392,N_9992,N_9863);
xnor U14393 (N_14393,N_9161,N_9060);
xor U14394 (N_14394,N_10458,N_10796);
nor U14395 (N_14395,N_11992,N_9148);
or U14396 (N_14396,N_10440,N_10300);
and U14397 (N_14397,N_9909,N_11821);
nor U14398 (N_14398,N_11172,N_9177);
nor U14399 (N_14399,N_9658,N_11147);
nor U14400 (N_14400,N_11732,N_10295);
and U14401 (N_14401,N_9966,N_10325);
or U14402 (N_14402,N_9161,N_10328);
and U14403 (N_14403,N_9907,N_11304);
nor U14404 (N_14404,N_10307,N_9141);
or U14405 (N_14405,N_9032,N_10650);
and U14406 (N_14406,N_11986,N_10094);
nand U14407 (N_14407,N_10087,N_9006);
nor U14408 (N_14408,N_9672,N_10341);
nor U14409 (N_14409,N_10577,N_9689);
or U14410 (N_14410,N_9701,N_9041);
nor U14411 (N_14411,N_9007,N_10320);
or U14412 (N_14412,N_10253,N_10956);
and U14413 (N_14413,N_10467,N_11790);
or U14414 (N_14414,N_11174,N_9278);
nor U14415 (N_14415,N_10679,N_10180);
nor U14416 (N_14416,N_9205,N_9093);
and U14417 (N_14417,N_11511,N_10296);
xor U14418 (N_14418,N_9016,N_11827);
and U14419 (N_14419,N_11571,N_10684);
nand U14420 (N_14420,N_9965,N_9726);
or U14421 (N_14421,N_11521,N_11224);
nand U14422 (N_14422,N_11276,N_11778);
and U14423 (N_14423,N_9238,N_9256);
or U14424 (N_14424,N_9930,N_9954);
nand U14425 (N_14425,N_10953,N_10397);
xor U14426 (N_14426,N_10118,N_9904);
nor U14427 (N_14427,N_11480,N_9294);
or U14428 (N_14428,N_10487,N_11352);
or U14429 (N_14429,N_11857,N_9032);
nor U14430 (N_14430,N_9998,N_10667);
nand U14431 (N_14431,N_11037,N_10579);
or U14432 (N_14432,N_11746,N_9527);
and U14433 (N_14433,N_11883,N_11645);
nand U14434 (N_14434,N_10757,N_9151);
or U14435 (N_14435,N_11253,N_11650);
and U14436 (N_14436,N_10835,N_9114);
nor U14437 (N_14437,N_11126,N_11357);
nand U14438 (N_14438,N_11634,N_10537);
or U14439 (N_14439,N_11052,N_10171);
nand U14440 (N_14440,N_9931,N_9347);
nor U14441 (N_14441,N_9978,N_11477);
nor U14442 (N_14442,N_10778,N_11366);
nand U14443 (N_14443,N_10525,N_11667);
nand U14444 (N_14444,N_10574,N_9252);
nor U14445 (N_14445,N_9729,N_10448);
nand U14446 (N_14446,N_9296,N_9491);
xnor U14447 (N_14447,N_9825,N_10148);
nor U14448 (N_14448,N_10026,N_9680);
nor U14449 (N_14449,N_11864,N_10257);
nor U14450 (N_14450,N_9192,N_10197);
xnor U14451 (N_14451,N_10863,N_10112);
and U14452 (N_14452,N_9396,N_10928);
nor U14453 (N_14453,N_11009,N_10218);
or U14454 (N_14454,N_9904,N_11839);
xnor U14455 (N_14455,N_11656,N_11193);
or U14456 (N_14456,N_11619,N_10321);
or U14457 (N_14457,N_11322,N_11435);
xor U14458 (N_14458,N_11241,N_10226);
nand U14459 (N_14459,N_11114,N_9575);
xnor U14460 (N_14460,N_10115,N_10816);
and U14461 (N_14461,N_10276,N_9716);
nor U14462 (N_14462,N_9249,N_10662);
nor U14463 (N_14463,N_9937,N_9595);
nor U14464 (N_14464,N_10546,N_9072);
xor U14465 (N_14465,N_9747,N_9090);
nand U14466 (N_14466,N_11425,N_9505);
nor U14467 (N_14467,N_11253,N_11378);
or U14468 (N_14468,N_10515,N_10002);
nand U14469 (N_14469,N_10882,N_10004);
nor U14470 (N_14470,N_11216,N_10183);
and U14471 (N_14471,N_9363,N_9384);
xnor U14472 (N_14472,N_11741,N_11384);
nor U14473 (N_14473,N_9788,N_10548);
and U14474 (N_14474,N_9351,N_9509);
and U14475 (N_14475,N_10764,N_10096);
nor U14476 (N_14476,N_10016,N_9602);
xor U14477 (N_14477,N_10394,N_9740);
nand U14478 (N_14478,N_9864,N_10310);
xnor U14479 (N_14479,N_11393,N_10341);
nand U14480 (N_14480,N_10754,N_9211);
and U14481 (N_14481,N_10403,N_10666);
or U14482 (N_14482,N_11141,N_10550);
nor U14483 (N_14483,N_10435,N_9931);
and U14484 (N_14484,N_9501,N_11526);
nand U14485 (N_14485,N_10616,N_9804);
xnor U14486 (N_14486,N_10516,N_10986);
xor U14487 (N_14487,N_9297,N_9047);
and U14488 (N_14488,N_11294,N_10202);
xnor U14489 (N_14489,N_9499,N_10064);
nand U14490 (N_14490,N_9881,N_11237);
or U14491 (N_14491,N_9391,N_10832);
nand U14492 (N_14492,N_9875,N_9206);
nand U14493 (N_14493,N_11018,N_11767);
nor U14494 (N_14494,N_9254,N_10096);
nand U14495 (N_14495,N_11949,N_9920);
xor U14496 (N_14496,N_11812,N_9083);
and U14497 (N_14497,N_11720,N_10428);
and U14498 (N_14498,N_11190,N_9046);
and U14499 (N_14499,N_9985,N_11267);
nor U14500 (N_14500,N_9403,N_11547);
and U14501 (N_14501,N_9378,N_11185);
nor U14502 (N_14502,N_11295,N_10201);
xor U14503 (N_14503,N_9466,N_9649);
nand U14504 (N_14504,N_9278,N_10046);
xor U14505 (N_14505,N_10157,N_10756);
xnor U14506 (N_14506,N_9366,N_11257);
nand U14507 (N_14507,N_9862,N_11504);
nand U14508 (N_14508,N_11648,N_9790);
or U14509 (N_14509,N_11030,N_9990);
and U14510 (N_14510,N_11914,N_9605);
or U14511 (N_14511,N_9086,N_10515);
nor U14512 (N_14512,N_11348,N_10757);
xor U14513 (N_14513,N_11726,N_9176);
nand U14514 (N_14514,N_10661,N_10738);
nor U14515 (N_14515,N_9910,N_11562);
nand U14516 (N_14516,N_9211,N_11608);
nand U14517 (N_14517,N_10577,N_9298);
and U14518 (N_14518,N_9905,N_9199);
nor U14519 (N_14519,N_10980,N_11294);
nor U14520 (N_14520,N_9521,N_9394);
or U14521 (N_14521,N_11666,N_9726);
or U14522 (N_14522,N_11815,N_9124);
and U14523 (N_14523,N_11992,N_11258);
or U14524 (N_14524,N_10088,N_11848);
nand U14525 (N_14525,N_9222,N_11427);
nand U14526 (N_14526,N_11205,N_9481);
nor U14527 (N_14527,N_11060,N_9066);
and U14528 (N_14528,N_9182,N_11824);
or U14529 (N_14529,N_10994,N_10692);
and U14530 (N_14530,N_11712,N_9636);
or U14531 (N_14531,N_11152,N_10836);
or U14532 (N_14532,N_11381,N_9104);
xnor U14533 (N_14533,N_11658,N_10595);
nor U14534 (N_14534,N_11129,N_9586);
or U14535 (N_14535,N_11881,N_9039);
nor U14536 (N_14536,N_10689,N_11805);
and U14537 (N_14537,N_9374,N_10920);
xnor U14538 (N_14538,N_11556,N_9336);
xnor U14539 (N_14539,N_9273,N_10463);
nand U14540 (N_14540,N_9320,N_10327);
xor U14541 (N_14541,N_9112,N_10968);
or U14542 (N_14542,N_10729,N_10489);
and U14543 (N_14543,N_10776,N_10990);
or U14544 (N_14544,N_9559,N_11831);
nand U14545 (N_14545,N_11516,N_10664);
nand U14546 (N_14546,N_10661,N_10198);
nand U14547 (N_14547,N_9720,N_10558);
and U14548 (N_14548,N_9140,N_9802);
nor U14549 (N_14549,N_11304,N_9776);
nor U14550 (N_14550,N_9345,N_10659);
nor U14551 (N_14551,N_10949,N_9613);
nand U14552 (N_14552,N_9155,N_10748);
and U14553 (N_14553,N_11010,N_10073);
nand U14554 (N_14554,N_10439,N_10417);
or U14555 (N_14555,N_9912,N_11956);
nand U14556 (N_14556,N_11587,N_11546);
or U14557 (N_14557,N_9262,N_11474);
nand U14558 (N_14558,N_9270,N_10938);
and U14559 (N_14559,N_11529,N_9267);
and U14560 (N_14560,N_9172,N_11074);
or U14561 (N_14561,N_9023,N_10320);
or U14562 (N_14562,N_10403,N_10260);
or U14563 (N_14563,N_9464,N_11850);
or U14564 (N_14564,N_9257,N_11741);
nand U14565 (N_14565,N_11049,N_11707);
nand U14566 (N_14566,N_11214,N_9159);
and U14567 (N_14567,N_9672,N_11737);
nor U14568 (N_14568,N_10477,N_10823);
nor U14569 (N_14569,N_11010,N_9316);
xnor U14570 (N_14570,N_9037,N_10621);
nor U14571 (N_14571,N_11751,N_11689);
or U14572 (N_14572,N_9069,N_11048);
nand U14573 (N_14573,N_11521,N_11044);
nor U14574 (N_14574,N_9649,N_9083);
nor U14575 (N_14575,N_9791,N_10333);
and U14576 (N_14576,N_10149,N_9491);
nand U14577 (N_14577,N_10234,N_9378);
nor U14578 (N_14578,N_10013,N_10730);
nor U14579 (N_14579,N_9768,N_9598);
xnor U14580 (N_14580,N_10828,N_11932);
nand U14581 (N_14581,N_10095,N_10769);
nand U14582 (N_14582,N_9791,N_10412);
or U14583 (N_14583,N_10888,N_11306);
nand U14584 (N_14584,N_10358,N_10306);
xor U14585 (N_14585,N_11327,N_9548);
nand U14586 (N_14586,N_10332,N_10989);
nor U14587 (N_14587,N_9327,N_9145);
xor U14588 (N_14588,N_11600,N_10481);
nand U14589 (N_14589,N_9643,N_11408);
nand U14590 (N_14590,N_10975,N_11891);
and U14591 (N_14591,N_11039,N_10379);
and U14592 (N_14592,N_11374,N_10612);
and U14593 (N_14593,N_9795,N_10482);
and U14594 (N_14594,N_10532,N_9874);
or U14595 (N_14595,N_11896,N_9824);
and U14596 (N_14596,N_9245,N_10894);
nand U14597 (N_14597,N_10553,N_9829);
nand U14598 (N_14598,N_11098,N_9808);
or U14599 (N_14599,N_10706,N_9186);
xor U14600 (N_14600,N_11733,N_10090);
nand U14601 (N_14601,N_11329,N_9050);
and U14602 (N_14602,N_9758,N_10387);
and U14603 (N_14603,N_9397,N_9779);
or U14604 (N_14604,N_10233,N_10712);
and U14605 (N_14605,N_10232,N_11955);
nand U14606 (N_14606,N_9848,N_10282);
nand U14607 (N_14607,N_11678,N_10442);
or U14608 (N_14608,N_11518,N_11988);
nand U14609 (N_14609,N_9155,N_9946);
xnor U14610 (N_14610,N_9113,N_10379);
and U14611 (N_14611,N_10180,N_11226);
nand U14612 (N_14612,N_11660,N_9853);
nor U14613 (N_14613,N_10005,N_11859);
nand U14614 (N_14614,N_10753,N_9465);
xnor U14615 (N_14615,N_10393,N_9201);
or U14616 (N_14616,N_10724,N_9100);
and U14617 (N_14617,N_9366,N_9750);
or U14618 (N_14618,N_10702,N_9031);
or U14619 (N_14619,N_11348,N_9344);
nand U14620 (N_14620,N_9380,N_10163);
nor U14621 (N_14621,N_10408,N_10797);
xnor U14622 (N_14622,N_11218,N_11645);
or U14623 (N_14623,N_9093,N_10959);
nor U14624 (N_14624,N_9929,N_11470);
and U14625 (N_14625,N_11948,N_10826);
or U14626 (N_14626,N_11847,N_9084);
and U14627 (N_14627,N_10266,N_9611);
and U14628 (N_14628,N_11130,N_9756);
nand U14629 (N_14629,N_11491,N_11952);
or U14630 (N_14630,N_11064,N_9474);
xnor U14631 (N_14631,N_11753,N_11522);
and U14632 (N_14632,N_11300,N_11593);
nand U14633 (N_14633,N_10043,N_9921);
or U14634 (N_14634,N_11024,N_10347);
nor U14635 (N_14635,N_10282,N_10447);
xnor U14636 (N_14636,N_11489,N_11796);
or U14637 (N_14637,N_11498,N_10672);
nand U14638 (N_14638,N_11908,N_11184);
and U14639 (N_14639,N_10424,N_10939);
nor U14640 (N_14640,N_11952,N_11460);
and U14641 (N_14641,N_10726,N_11871);
nand U14642 (N_14642,N_9361,N_10596);
nor U14643 (N_14643,N_11649,N_11636);
nor U14644 (N_14644,N_10989,N_10643);
nor U14645 (N_14645,N_11697,N_11338);
nor U14646 (N_14646,N_10720,N_10766);
or U14647 (N_14647,N_9719,N_10330);
and U14648 (N_14648,N_10827,N_9673);
and U14649 (N_14649,N_9652,N_9691);
nand U14650 (N_14650,N_10599,N_11833);
or U14651 (N_14651,N_11711,N_10411);
nand U14652 (N_14652,N_9383,N_11473);
and U14653 (N_14653,N_11089,N_9928);
nand U14654 (N_14654,N_9569,N_10505);
nand U14655 (N_14655,N_10433,N_11744);
and U14656 (N_14656,N_10861,N_9823);
xor U14657 (N_14657,N_10567,N_11449);
and U14658 (N_14658,N_11200,N_10629);
and U14659 (N_14659,N_10578,N_10783);
and U14660 (N_14660,N_9152,N_11124);
and U14661 (N_14661,N_10945,N_11859);
and U14662 (N_14662,N_10490,N_10899);
nand U14663 (N_14663,N_9912,N_9893);
and U14664 (N_14664,N_9842,N_11372);
or U14665 (N_14665,N_11491,N_9636);
nand U14666 (N_14666,N_10699,N_10968);
nor U14667 (N_14667,N_9645,N_9962);
nor U14668 (N_14668,N_10278,N_11570);
and U14669 (N_14669,N_11847,N_11014);
and U14670 (N_14670,N_11598,N_11318);
nand U14671 (N_14671,N_11289,N_10243);
and U14672 (N_14672,N_10362,N_11154);
and U14673 (N_14673,N_9864,N_11855);
nor U14674 (N_14674,N_11343,N_11811);
or U14675 (N_14675,N_10980,N_9215);
or U14676 (N_14676,N_9628,N_10333);
or U14677 (N_14677,N_10296,N_10384);
nand U14678 (N_14678,N_10863,N_11626);
nor U14679 (N_14679,N_10809,N_11513);
or U14680 (N_14680,N_10311,N_10630);
nand U14681 (N_14681,N_9531,N_10010);
nor U14682 (N_14682,N_10378,N_9994);
and U14683 (N_14683,N_10639,N_9500);
nand U14684 (N_14684,N_10602,N_9944);
nand U14685 (N_14685,N_9630,N_11296);
nor U14686 (N_14686,N_9573,N_11687);
or U14687 (N_14687,N_9329,N_10115);
xor U14688 (N_14688,N_11636,N_9491);
and U14689 (N_14689,N_10171,N_11415);
nand U14690 (N_14690,N_9576,N_11320);
and U14691 (N_14691,N_11673,N_9656);
nand U14692 (N_14692,N_9210,N_10548);
nor U14693 (N_14693,N_11197,N_9929);
nand U14694 (N_14694,N_11591,N_11174);
xnor U14695 (N_14695,N_11505,N_10494);
and U14696 (N_14696,N_10849,N_9463);
nand U14697 (N_14697,N_11574,N_9305);
nand U14698 (N_14698,N_11457,N_9050);
and U14699 (N_14699,N_9390,N_11185);
nand U14700 (N_14700,N_11617,N_9173);
or U14701 (N_14701,N_9900,N_11474);
xor U14702 (N_14702,N_11576,N_11679);
or U14703 (N_14703,N_11021,N_10971);
nand U14704 (N_14704,N_9797,N_10316);
or U14705 (N_14705,N_11298,N_11566);
and U14706 (N_14706,N_9432,N_9033);
nand U14707 (N_14707,N_9359,N_10589);
nand U14708 (N_14708,N_10213,N_11195);
nor U14709 (N_14709,N_9403,N_9967);
nor U14710 (N_14710,N_10938,N_10866);
nor U14711 (N_14711,N_10793,N_11029);
or U14712 (N_14712,N_10293,N_9748);
nor U14713 (N_14713,N_10724,N_11742);
and U14714 (N_14714,N_11743,N_10314);
or U14715 (N_14715,N_11219,N_11419);
nor U14716 (N_14716,N_11379,N_10820);
and U14717 (N_14717,N_11971,N_9462);
and U14718 (N_14718,N_11238,N_11304);
xnor U14719 (N_14719,N_9521,N_9729);
nand U14720 (N_14720,N_9524,N_11354);
nor U14721 (N_14721,N_11268,N_9775);
or U14722 (N_14722,N_11061,N_11697);
nand U14723 (N_14723,N_10888,N_10255);
nor U14724 (N_14724,N_9218,N_11733);
or U14725 (N_14725,N_10462,N_11282);
or U14726 (N_14726,N_11764,N_10074);
or U14727 (N_14727,N_9440,N_9313);
nor U14728 (N_14728,N_9521,N_11265);
nand U14729 (N_14729,N_10710,N_11714);
nand U14730 (N_14730,N_9732,N_11411);
nand U14731 (N_14731,N_10208,N_10669);
or U14732 (N_14732,N_11958,N_10442);
or U14733 (N_14733,N_11478,N_10674);
and U14734 (N_14734,N_9862,N_10262);
xor U14735 (N_14735,N_9986,N_9066);
and U14736 (N_14736,N_9922,N_10661);
or U14737 (N_14737,N_9248,N_11586);
or U14738 (N_14738,N_11039,N_10950);
nand U14739 (N_14739,N_9900,N_10572);
or U14740 (N_14740,N_10474,N_9081);
nor U14741 (N_14741,N_11125,N_11767);
or U14742 (N_14742,N_9806,N_9476);
or U14743 (N_14743,N_9214,N_9578);
nand U14744 (N_14744,N_9602,N_9944);
xor U14745 (N_14745,N_11359,N_10171);
and U14746 (N_14746,N_10733,N_9645);
or U14747 (N_14747,N_10919,N_9872);
xnor U14748 (N_14748,N_10059,N_9560);
and U14749 (N_14749,N_9303,N_11262);
nand U14750 (N_14750,N_9956,N_9680);
or U14751 (N_14751,N_11475,N_11772);
or U14752 (N_14752,N_10571,N_10622);
or U14753 (N_14753,N_9677,N_11956);
nand U14754 (N_14754,N_10843,N_9209);
nand U14755 (N_14755,N_11055,N_11871);
and U14756 (N_14756,N_11908,N_11917);
and U14757 (N_14757,N_9068,N_11529);
xnor U14758 (N_14758,N_11887,N_9036);
and U14759 (N_14759,N_10836,N_11610);
or U14760 (N_14760,N_11094,N_10684);
and U14761 (N_14761,N_9725,N_11119);
and U14762 (N_14762,N_9427,N_10405);
nand U14763 (N_14763,N_10560,N_11352);
or U14764 (N_14764,N_9953,N_9495);
and U14765 (N_14765,N_9510,N_11554);
nor U14766 (N_14766,N_10621,N_11723);
nand U14767 (N_14767,N_10666,N_9303);
or U14768 (N_14768,N_10274,N_10128);
or U14769 (N_14769,N_9793,N_11287);
xor U14770 (N_14770,N_11257,N_9193);
and U14771 (N_14771,N_9769,N_11957);
nor U14772 (N_14772,N_11148,N_11681);
nor U14773 (N_14773,N_10421,N_11281);
nor U14774 (N_14774,N_9408,N_9002);
or U14775 (N_14775,N_10409,N_9529);
nor U14776 (N_14776,N_11093,N_9233);
nand U14777 (N_14777,N_9988,N_11551);
nand U14778 (N_14778,N_9978,N_11965);
or U14779 (N_14779,N_9650,N_10650);
nor U14780 (N_14780,N_9055,N_11930);
nand U14781 (N_14781,N_10343,N_9270);
nor U14782 (N_14782,N_9657,N_9661);
nand U14783 (N_14783,N_11639,N_10053);
or U14784 (N_14784,N_9402,N_11467);
nand U14785 (N_14785,N_9360,N_10155);
nand U14786 (N_14786,N_11234,N_10277);
or U14787 (N_14787,N_9743,N_10867);
nor U14788 (N_14788,N_10464,N_11848);
nand U14789 (N_14789,N_11542,N_11293);
nand U14790 (N_14790,N_9696,N_9229);
xnor U14791 (N_14791,N_9171,N_11128);
and U14792 (N_14792,N_11333,N_11857);
nand U14793 (N_14793,N_9216,N_11727);
or U14794 (N_14794,N_9452,N_11931);
xor U14795 (N_14795,N_11756,N_11105);
nand U14796 (N_14796,N_11011,N_9351);
and U14797 (N_14797,N_11367,N_10090);
nand U14798 (N_14798,N_10238,N_11800);
nand U14799 (N_14799,N_9418,N_10913);
nand U14800 (N_14800,N_10867,N_10580);
or U14801 (N_14801,N_10061,N_11402);
or U14802 (N_14802,N_10024,N_9444);
and U14803 (N_14803,N_11208,N_9256);
nand U14804 (N_14804,N_9745,N_11962);
nor U14805 (N_14805,N_9013,N_10697);
and U14806 (N_14806,N_11201,N_10589);
xor U14807 (N_14807,N_11233,N_10183);
nor U14808 (N_14808,N_11343,N_9484);
and U14809 (N_14809,N_9679,N_10052);
nand U14810 (N_14810,N_10642,N_9434);
nor U14811 (N_14811,N_11597,N_9249);
or U14812 (N_14812,N_9433,N_10790);
and U14813 (N_14813,N_9854,N_10410);
nand U14814 (N_14814,N_10594,N_11732);
and U14815 (N_14815,N_11629,N_10315);
xnor U14816 (N_14816,N_11426,N_9037);
nand U14817 (N_14817,N_9990,N_11730);
or U14818 (N_14818,N_11718,N_11539);
nand U14819 (N_14819,N_11557,N_11660);
or U14820 (N_14820,N_10423,N_9670);
or U14821 (N_14821,N_11136,N_11877);
and U14822 (N_14822,N_9072,N_9368);
and U14823 (N_14823,N_11603,N_9368);
nor U14824 (N_14824,N_9689,N_9013);
or U14825 (N_14825,N_11334,N_9745);
and U14826 (N_14826,N_9941,N_10873);
nand U14827 (N_14827,N_9476,N_11984);
nand U14828 (N_14828,N_9131,N_9641);
or U14829 (N_14829,N_9436,N_11950);
nand U14830 (N_14830,N_9891,N_10458);
nand U14831 (N_14831,N_9325,N_11329);
or U14832 (N_14832,N_10502,N_10862);
and U14833 (N_14833,N_10101,N_11746);
nor U14834 (N_14834,N_10133,N_11645);
nand U14835 (N_14835,N_11925,N_10698);
and U14836 (N_14836,N_9759,N_9434);
nand U14837 (N_14837,N_10499,N_11021);
and U14838 (N_14838,N_11536,N_9733);
or U14839 (N_14839,N_9059,N_11883);
or U14840 (N_14840,N_11909,N_9426);
or U14841 (N_14841,N_11697,N_9916);
or U14842 (N_14842,N_9502,N_9841);
or U14843 (N_14843,N_9195,N_10006);
or U14844 (N_14844,N_9764,N_9080);
nor U14845 (N_14845,N_10380,N_11073);
nor U14846 (N_14846,N_9041,N_9034);
or U14847 (N_14847,N_10209,N_11158);
or U14848 (N_14848,N_9615,N_11172);
nor U14849 (N_14849,N_10885,N_10694);
nand U14850 (N_14850,N_11224,N_11045);
nand U14851 (N_14851,N_11647,N_11205);
or U14852 (N_14852,N_11134,N_10123);
or U14853 (N_14853,N_10172,N_9597);
and U14854 (N_14854,N_10236,N_9394);
or U14855 (N_14855,N_9505,N_10612);
nand U14856 (N_14856,N_11201,N_9017);
and U14857 (N_14857,N_11949,N_9900);
or U14858 (N_14858,N_9998,N_9422);
nand U14859 (N_14859,N_9298,N_9136);
nand U14860 (N_14860,N_11960,N_10040);
and U14861 (N_14861,N_10873,N_10533);
xor U14862 (N_14862,N_9304,N_11532);
or U14863 (N_14863,N_10752,N_9484);
nor U14864 (N_14864,N_10501,N_10575);
xor U14865 (N_14865,N_9048,N_10963);
nand U14866 (N_14866,N_10437,N_11034);
or U14867 (N_14867,N_10224,N_10680);
nand U14868 (N_14868,N_10323,N_9947);
nor U14869 (N_14869,N_11680,N_11593);
nor U14870 (N_14870,N_11610,N_11318);
nor U14871 (N_14871,N_10601,N_9866);
nor U14872 (N_14872,N_11283,N_10618);
or U14873 (N_14873,N_10765,N_9157);
or U14874 (N_14874,N_11326,N_11063);
nor U14875 (N_14875,N_11689,N_10518);
or U14876 (N_14876,N_9397,N_9680);
nand U14877 (N_14877,N_9582,N_10317);
and U14878 (N_14878,N_10238,N_10868);
and U14879 (N_14879,N_10093,N_11337);
or U14880 (N_14880,N_9461,N_9232);
xnor U14881 (N_14881,N_9309,N_11943);
and U14882 (N_14882,N_10038,N_11591);
and U14883 (N_14883,N_10426,N_10888);
nand U14884 (N_14884,N_11066,N_9764);
and U14885 (N_14885,N_10514,N_10242);
xnor U14886 (N_14886,N_10289,N_11798);
xor U14887 (N_14887,N_9136,N_11629);
or U14888 (N_14888,N_9028,N_9984);
nand U14889 (N_14889,N_10450,N_10251);
nand U14890 (N_14890,N_10223,N_9375);
and U14891 (N_14891,N_11157,N_9025);
nor U14892 (N_14892,N_11855,N_10243);
nand U14893 (N_14893,N_11090,N_9312);
and U14894 (N_14894,N_10022,N_9915);
or U14895 (N_14895,N_10861,N_9903);
and U14896 (N_14896,N_10056,N_9793);
and U14897 (N_14897,N_9622,N_9268);
and U14898 (N_14898,N_9185,N_11426);
or U14899 (N_14899,N_10459,N_9437);
nand U14900 (N_14900,N_9809,N_11798);
nand U14901 (N_14901,N_10434,N_11084);
and U14902 (N_14902,N_9863,N_10713);
nand U14903 (N_14903,N_11505,N_11187);
xor U14904 (N_14904,N_9793,N_10494);
nor U14905 (N_14905,N_11402,N_10178);
or U14906 (N_14906,N_10221,N_10016);
and U14907 (N_14907,N_11830,N_9725);
nand U14908 (N_14908,N_11229,N_10890);
or U14909 (N_14909,N_9320,N_10411);
and U14910 (N_14910,N_11442,N_11664);
or U14911 (N_14911,N_11423,N_10848);
nand U14912 (N_14912,N_9441,N_10293);
nor U14913 (N_14913,N_10181,N_9997);
nand U14914 (N_14914,N_11165,N_11345);
nand U14915 (N_14915,N_9276,N_9210);
nand U14916 (N_14916,N_9229,N_11281);
or U14917 (N_14917,N_11498,N_9927);
or U14918 (N_14918,N_10719,N_11882);
and U14919 (N_14919,N_9012,N_9121);
xor U14920 (N_14920,N_10357,N_9771);
nand U14921 (N_14921,N_9247,N_9095);
nor U14922 (N_14922,N_10031,N_11858);
nand U14923 (N_14923,N_9164,N_10133);
nand U14924 (N_14924,N_11214,N_10911);
nand U14925 (N_14925,N_11550,N_11567);
and U14926 (N_14926,N_11062,N_11653);
or U14927 (N_14927,N_9435,N_9489);
or U14928 (N_14928,N_10132,N_9586);
or U14929 (N_14929,N_10296,N_9753);
nand U14930 (N_14930,N_9057,N_9112);
xor U14931 (N_14931,N_11747,N_9240);
nor U14932 (N_14932,N_9013,N_10110);
xnor U14933 (N_14933,N_11622,N_10597);
nor U14934 (N_14934,N_10864,N_9558);
or U14935 (N_14935,N_11674,N_10827);
nand U14936 (N_14936,N_10271,N_11022);
and U14937 (N_14937,N_11169,N_10271);
nand U14938 (N_14938,N_11308,N_10098);
nor U14939 (N_14939,N_11233,N_11309);
xor U14940 (N_14940,N_11325,N_11282);
or U14941 (N_14941,N_10799,N_11585);
nand U14942 (N_14942,N_9269,N_10150);
nor U14943 (N_14943,N_10616,N_11186);
and U14944 (N_14944,N_9112,N_9541);
nor U14945 (N_14945,N_9967,N_10751);
nor U14946 (N_14946,N_11904,N_11160);
or U14947 (N_14947,N_10719,N_10484);
nand U14948 (N_14948,N_10202,N_9251);
nor U14949 (N_14949,N_10242,N_10048);
nand U14950 (N_14950,N_11553,N_11976);
xnor U14951 (N_14951,N_11994,N_10361);
nor U14952 (N_14952,N_11438,N_11251);
or U14953 (N_14953,N_10813,N_11094);
nand U14954 (N_14954,N_9660,N_11978);
nand U14955 (N_14955,N_10262,N_9092);
xor U14956 (N_14956,N_9829,N_9395);
or U14957 (N_14957,N_10450,N_11950);
nand U14958 (N_14958,N_11470,N_11581);
nor U14959 (N_14959,N_10005,N_11381);
nor U14960 (N_14960,N_9840,N_10451);
xnor U14961 (N_14961,N_11691,N_9080);
and U14962 (N_14962,N_9575,N_9194);
nand U14963 (N_14963,N_11394,N_11680);
and U14964 (N_14964,N_9612,N_9460);
or U14965 (N_14965,N_11929,N_11297);
or U14966 (N_14966,N_11302,N_10233);
nor U14967 (N_14967,N_11178,N_11563);
and U14968 (N_14968,N_10236,N_11213);
nand U14969 (N_14969,N_10622,N_11263);
nor U14970 (N_14970,N_9101,N_11081);
or U14971 (N_14971,N_9442,N_9424);
nand U14972 (N_14972,N_9916,N_10894);
xor U14973 (N_14973,N_11586,N_10246);
and U14974 (N_14974,N_9283,N_11198);
or U14975 (N_14975,N_9907,N_9122);
nand U14976 (N_14976,N_11436,N_9400);
and U14977 (N_14977,N_10139,N_11483);
or U14978 (N_14978,N_11806,N_11229);
and U14979 (N_14979,N_11127,N_11176);
or U14980 (N_14980,N_11517,N_11833);
nand U14981 (N_14981,N_9675,N_10707);
or U14982 (N_14982,N_9489,N_10507);
and U14983 (N_14983,N_11198,N_10995);
nor U14984 (N_14984,N_9581,N_11954);
or U14985 (N_14985,N_10069,N_9738);
nor U14986 (N_14986,N_10927,N_9693);
nand U14987 (N_14987,N_10607,N_10327);
and U14988 (N_14988,N_11216,N_10730);
nor U14989 (N_14989,N_11534,N_10939);
nor U14990 (N_14990,N_10352,N_11843);
and U14991 (N_14991,N_11171,N_10601);
nor U14992 (N_14992,N_10029,N_10586);
xnor U14993 (N_14993,N_10348,N_10617);
or U14994 (N_14994,N_9515,N_11869);
or U14995 (N_14995,N_11693,N_11309);
xnor U14996 (N_14996,N_9825,N_11115);
nand U14997 (N_14997,N_10192,N_10404);
and U14998 (N_14998,N_11732,N_9655);
nand U14999 (N_14999,N_11949,N_9138);
and UO_0 (O_0,N_14218,N_12205);
xnor UO_1 (O_1,N_12252,N_12562);
nor UO_2 (O_2,N_14044,N_14008);
and UO_3 (O_3,N_12813,N_12588);
xor UO_4 (O_4,N_13447,N_13947);
nand UO_5 (O_5,N_12627,N_13411);
or UO_6 (O_6,N_12116,N_13295);
nand UO_7 (O_7,N_13938,N_13982);
nor UO_8 (O_8,N_14715,N_12210);
xnor UO_9 (O_9,N_14343,N_12648);
or UO_10 (O_10,N_12092,N_12216);
and UO_11 (O_11,N_12947,N_12482);
or UO_12 (O_12,N_12053,N_12453);
nand UO_13 (O_13,N_13766,N_12046);
or UO_14 (O_14,N_12896,N_14348);
and UO_15 (O_15,N_13016,N_14811);
nand UO_16 (O_16,N_14308,N_13155);
nand UO_17 (O_17,N_13422,N_12071);
and UO_18 (O_18,N_12891,N_12610);
nand UO_19 (O_19,N_13256,N_14472);
and UO_20 (O_20,N_13444,N_14082);
nand UO_21 (O_21,N_13736,N_13082);
and UO_22 (O_22,N_12587,N_14248);
nand UO_23 (O_23,N_13480,N_12917);
nand UO_24 (O_24,N_14532,N_12598);
xor UO_25 (O_25,N_13613,N_14279);
nand UO_26 (O_26,N_13783,N_13492);
xnor UO_27 (O_27,N_14451,N_14971);
or UO_28 (O_28,N_13590,N_14499);
and UO_29 (O_29,N_14745,N_13585);
or UO_30 (O_30,N_13934,N_13928);
nand UO_31 (O_31,N_14938,N_12282);
xnor UO_32 (O_32,N_13290,N_12854);
nand UO_33 (O_33,N_12238,N_12393);
and UO_34 (O_34,N_14447,N_13568);
or UO_35 (O_35,N_14895,N_12272);
nand UO_36 (O_36,N_13281,N_13709);
and UO_37 (O_37,N_14098,N_12439);
and UO_38 (O_38,N_12800,N_12944);
or UO_39 (O_39,N_12853,N_14739);
nor UO_40 (O_40,N_13968,N_14861);
xor UO_41 (O_41,N_14087,N_14840);
nor UO_42 (O_42,N_14870,N_13466);
xnor UO_43 (O_43,N_14776,N_12688);
nand UO_44 (O_44,N_12605,N_12007);
nand UO_45 (O_45,N_13406,N_14305);
and UO_46 (O_46,N_12994,N_13380);
and UO_47 (O_47,N_13318,N_12554);
nand UO_48 (O_48,N_14013,N_12961);
and UO_49 (O_49,N_14362,N_12114);
nand UO_50 (O_50,N_12111,N_14333);
or UO_51 (O_51,N_13743,N_14028);
and UO_52 (O_52,N_14859,N_14069);
and UO_53 (O_53,N_12228,N_14416);
and UO_54 (O_54,N_14671,N_12038);
nor UO_55 (O_55,N_12101,N_13985);
or UO_56 (O_56,N_12019,N_12715);
nand UO_57 (O_57,N_13143,N_12327);
and UO_58 (O_58,N_13080,N_13296);
nand UO_59 (O_59,N_13085,N_13469);
nand UO_60 (O_60,N_12409,N_12480);
nand UO_61 (O_61,N_13821,N_14146);
nor UO_62 (O_62,N_14823,N_13600);
nand UO_63 (O_63,N_13591,N_13701);
or UO_64 (O_64,N_14653,N_12576);
nor UO_65 (O_65,N_12886,N_13673);
and UO_66 (O_66,N_13930,N_14378);
xnor UO_67 (O_67,N_12733,N_13527);
and UO_68 (O_68,N_14595,N_12788);
and UO_69 (O_69,N_13625,N_14236);
or UO_70 (O_70,N_14303,N_14970);
or UO_71 (O_71,N_14364,N_13570);
nor UO_72 (O_72,N_13312,N_12560);
nand UO_73 (O_73,N_12615,N_14864);
nor UO_74 (O_74,N_14341,N_12000);
nor UO_75 (O_75,N_13837,N_14926);
nor UO_76 (O_76,N_13316,N_14093);
or UO_77 (O_77,N_13797,N_13587);
or UO_78 (O_78,N_13504,N_12821);
and UO_79 (O_79,N_13962,N_12028);
nor UO_80 (O_80,N_14153,N_14721);
and UO_81 (O_81,N_14126,N_13638);
nor UO_82 (O_82,N_13545,N_12481);
nand UO_83 (O_83,N_14597,N_14889);
nand UO_84 (O_84,N_13567,N_13547);
nand UO_85 (O_85,N_14462,N_14458);
nor UO_86 (O_86,N_13219,N_12218);
nor UO_87 (O_87,N_14373,N_12951);
or UO_88 (O_88,N_14273,N_12465);
or UO_89 (O_89,N_12634,N_12267);
and UO_90 (O_90,N_13394,N_14981);
nor UO_91 (O_91,N_14824,N_12100);
and UO_92 (O_92,N_14887,N_14977);
or UO_93 (O_93,N_12413,N_12270);
nand UO_94 (O_94,N_12421,N_13522);
or UO_95 (O_95,N_13734,N_12379);
nand UO_96 (O_96,N_14893,N_13706);
or UO_97 (O_97,N_13851,N_13131);
nor UO_98 (O_98,N_13999,N_12483);
nor UO_99 (O_99,N_12257,N_14152);
nand UO_100 (O_100,N_13903,N_14580);
nand UO_101 (O_101,N_12226,N_13429);
or UO_102 (O_102,N_13006,N_14581);
nand UO_103 (O_103,N_14641,N_13123);
or UO_104 (O_104,N_13328,N_12207);
nand UO_105 (O_105,N_14337,N_12713);
nor UO_106 (O_106,N_13978,N_14400);
nor UO_107 (O_107,N_12743,N_12768);
and UO_108 (O_108,N_12297,N_12645);
or UO_109 (O_109,N_14097,N_14890);
xnor UO_110 (O_110,N_14149,N_12845);
and UO_111 (O_111,N_14888,N_13848);
nand UO_112 (O_112,N_13285,N_14984);
nand UO_113 (O_113,N_13060,N_12415);
nand UO_114 (O_114,N_12241,N_14527);
xnor UO_115 (O_115,N_14592,N_12646);
nor UO_116 (O_116,N_12868,N_13307);
and UO_117 (O_117,N_14217,N_13461);
and UO_118 (O_118,N_14955,N_13643);
or UO_119 (O_119,N_13923,N_14301);
nor UO_120 (O_120,N_12495,N_13517);
and UO_121 (O_121,N_14139,N_13136);
nor UO_122 (O_122,N_14102,N_14247);
nor UO_123 (O_123,N_13824,N_12739);
nor UO_124 (O_124,N_12434,N_12949);
and UO_125 (O_125,N_14805,N_13327);
nor UO_126 (O_126,N_12815,N_13105);
nand UO_127 (O_127,N_12590,N_14531);
nand UO_128 (O_128,N_14578,N_12163);
and UO_129 (O_129,N_13456,N_12749);
nor UO_130 (O_130,N_12955,N_13214);
nand UO_131 (O_131,N_14334,N_13297);
or UO_132 (O_132,N_13449,N_14645);
nand UO_133 (O_133,N_13718,N_12844);
or UO_134 (O_134,N_12318,N_14251);
and UO_135 (O_135,N_13387,N_13166);
nor UO_136 (O_136,N_12344,N_14338);
or UO_137 (O_137,N_14120,N_13635);
nor UO_138 (O_138,N_13691,N_13656);
or UO_139 (O_139,N_14293,N_13110);
nand UO_140 (O_140,N_12303,N_13249);
xnor UO_141 (O_141,N_14090,N_14556);
nand UO_142 (O_142,N_14929,N_14414);
nand UO_143 (O_143,N_13189,N_12099);
or UO_144 (O_144,N_13306,N_13688);
nand UO_145 (O_145,N_14815,N_12472);
nor UO_146 (O_146,N_12513,N_13814);
and UO_147 (O_147,N_14567,N_12431);
and UO_148 (O_148,N_12363,N_12013);
xor UO_149 (O_149,N_12871,N_12120);
or UO_150 (O_150,N_13017,N_14468);
or UO_151 (O_151,N_13644,N_14906);
and UO_152 (O_152,N_14813,N_13030);
or UO_153 (O_153,N_12798,N_13767);
xnor UO_154 (O_154,N_14195,N_14200);
nor UO_155 (O_155,N_14322,N_12179);
or UO_156 (O_156,N_13075,N_14134);
xor UO_157 (O_157,N_12172,N_14422);
and UO_158 (O_158,N_13800,N_13258);
nand UO_159 (O_159,N_13915,N_12849);
or UO_160 (O_160,N_14335,N_14518);
xnor UO_161 (O_161,N_12682,N_13571);
nand UO_162 (O_162,N_12649,N_14446);
nor UO_163 (O_163,N_13402,N_14875);
and UO_164 (O_164,N_14467,N_13623);
nor UO_165 (O_165,N_14826,N_13437);
nand UO_166 (O_166,N_12578,N_13941);
and UO_167 (O_167,N_12325,N_13093);
nor UO_168 (O_168,N_13707,N_13605);
nand UO_169 (O_169,N_13788,N_12312);
nand UO_170 (O_170,N_12443,N_14159);
nor UO_171 (O_171,N_14219,N_13802);
nand UO_172 (O_172,N_13191,N_14212);
and UO_173 (O_173,N_13678,N_12503);
nor UO_174 (O_174,N_13112,N_13020);
nor UO_175 (O_175,N_12766,N_14729);
nor UO_176 (O_176,N_13500,N_12869);
nor UO_177 (O_177,N_13792,N_14491);
or UO_178 (O_178,N_14798,N_14554);
nand UO_179 (O_179,N_12231,N_12115);
or UO_180 (O_180,N_14872,N_13827);
and UO_181 (O_181,N_14135,N_13876);
and UO_182 (O_182,N_12076,N_12670);
nand UO_183 (O_183,N_14295,N_12102);
xnor UO_184 (O_184,N_14342,N_13597);
nor UO_185 (O_185,N_12694,N_14232);
nor UO_186 (O_186,N_14257,N_13910);
and UO_187 (O_187,N_12242,N_12804);
xnor UO_188 (O_188,N_13778,N_13637);
nor UO_189 (O_189,N_13835,N_12121);
and UO_190 (O_190,N_12736,N_13132);
and UO_191 (O_191,N_13704,N_13007);
and UO_192 (O_192,N_12109,N_12095);
and UO_193 (O_193,N_13787,N_12463);
nor UO_194 (O_194,N_14905,N_14525);
nor UO_195 (O_195,N_12012,N_14634);
or UO_196 (O_196,N_13458,N_14050);
and UO_197 (O_197,N_14281,N_14290);
nand UO_198 (O_198,N_12974,N_13419);
or UO_199 (O_199,N_14724,N_13426);
and UO_200 (O_200,N_14880,N_13231);
or UO_201 (O_201,N_12572,N_14331);
or UO_202 (O_202,N_14546,N_12760);
or UO_203 (O_203,N_13703,N_13395);
nor UO_204 (O_204,N_13984,N_13867);
or UO_205 (O_205,N_12320,N_13680);
and UO_206 (O_206,N_14151,N_12156);
nand UO_207 (O_207,N_14317,N_12208);
nor UO_208 (O_208,N_12628,N_12920);
and UO_209 (O_209,N_13323,N_13194);
and UO_210 (O_210,N_12925,N_13125);
and UO_211 (O_211,N_14372,N_12650);
and UO_212 (O_212,N_12767,N_13196);
and UO_213 (O_213,N_14019,N_12746);
nand UO_214 (O_214,N_13742,N_12685);
nor UO_215 (O_215,N_12461,N_13725);
nand UO_216 (O_216,N_14109,N_14011);
and UO_217 (O_217,N_13945,N_12151);
xnor UO_218 (O_218,N_14434,N_13081);
xor UO_219 (O_219,N_14605,N_13755);
xnor UO_220 (O_220,N_13954,N_13834);
xor UO_221 (O_221,N_12086,N_13538);
nor UO_222 (O_222,N_13119,N_12784);
nand UO_223 (O_223,N_14716,N_14586);
nand UO_224 (O_224,N_14780,N_14140);
nand UO_225 (O_225,N_13168,N_12936);
or UO_226 (O_226,N_14182,N_13385);
or UO_227 (O_227,N_13615,N_14831);
nand UO_228 (O_228,N_14616,N_14039);
or UO_229 (O_229,N_14355,N_13350);
and UO_230 (O_230,N_14316,N_14995);
nor UO_231 (O_231,N_13651,N_14101);
nand UO_232 (O_232,N_14306,N_14800);
xnor UO_233 (O_233,N_13495,N_12184);
nor UO_234 (O_234,N_14818,N_12809);
nand UO_235 (O_235,N_14145,N_12976);
and UO_236 (O_236,N_14670,N_12905);
nand UO_237 (O_237,N_12334,N_12337);
nor UO_238 (O_238,N_12211,N_12764);
and UO_239 (O_239,N_12175,N_14601);
and UO_240 (O_240,N_14261,N_12631);
nand UO_241 (O_241,N_12675,N_13404);
nand UO_242 (O_242,N_13087,N_13496);
xor UO_243 (O_243,N_13149,N_12791);
or UO_244 (O_244,N_12992,N_14137);
and UO_245 (O_245,N_14487,N_12085);
nor UO_246 (O_246,N_12504,N_14919);
and UO_247 (O_247,N_14276,N_13685);
and UO_248 (O_248,N_13282,N_12130);
and UO_249 (O_249,N_12359,N_13184);
or UO_250 (O_250,N_14899,N_12841);
or UO_251 (O_251,N_14832,N_13548);
nor UO_252 (O_252,N_12014,N_12220);
or UO_253 (O_253,N_13885,N_12331);
nor UO_254 (O_254,N_14830,N_13375);
nor UO_255 (O_255,N_14593,N_12923);
xnor UO_256 (O_256,N_14756,N_13309);
or UO_257 (O_257,N_14196,N_12607);
or UO_258 (O_258,N_12293,N_13852);
xor UO_259 (O_259,N_13510,N_13435);
and UO_260 (O_260,N_14479,N_14821);
xnor UO_261 (O_261,N_12322,N_12471);
or UO_262 (O_262,N_14561,N_12286);
and UO_263 (O_263,N_14891,N_12591);
and UO_264 (O_264,N_12098,N_14533);
xnor UO_265 (O_265,N_13407,N_13055);
nand UO_266 (O_266,N_12909,N_14631);
nor UO_267 (O_267,N_14522,N_14264);
nor UO_268 (O_268,N_14178,N_12536);
or UO_269 (O_269,N_14637,N_13433);
nand UO_270 (O_270,N_13997,N_13721);
nand UO_271 (O_271,N_14998,N_12235);
and UO_272 (O_272,N_13201,N_14792);
nor UO_273 (O_273,N_12987,N_13576);
and UO_274 (O_274,N_14509,N_14598);
nor UO_275 (O_275,N_12189,N_12150);
nor UO_276 (O_276,N_14526,N_14224);
and UO_277 (O_277,N_14231,N_13206);
or UO_278 (O_278,N_13807,N_12647);
or UO_279 (O_279,N_14494,N_13056);
nand UO_280 (O_280,N_12703,N_12149);
and UO_281 (O_281,N_13425,N_14353);
and UO_282 (O_282,N_12772,N_13209);
xor UO_283 (O_283,N_14997,N_14515);
xor UO_284 (O_284,N_13374,N_12043);
nor UO_285 (O_285,N_12903,N_12173);
and UO_286 (O_286,N_14842,N_13618);
nand UO_287 (O_287,N_13241,N_12959);
nand UO_288 (O_288,N_13135,N_14594);
and UO_289 (O_289,N_13560,N_14537);
nor UO_290 (O_290,N_13803,N_12898);
or UO_291 (O_291,N_14208,N_12787);
nand UO_292 (O_292,N_12152,N_14848);
nor UO_293 (O_293,N_12024,N_13352);
or UO_294 (O_294,N_12507,N_13544);
nor UO_295 (O_295,N_14511,N_14184);
or UO_296 (O_296,N_14636,N_13430);
or UO_297 (O_297,N_12432,N_12518);
nand UO_298 (O_298,N_14370,N_13239);
or UO_299 (O_299,N_13111,N_12187);
and UO_300 (O_300,N_13397,N_14775);
and UO_301 (O_301,N_12381,N_12351);
nand UO_302 (O_302,N_12001,N_13553);
or UO_303 (O_303,N_14603,N_13793);
nor UO_304 (O_304,N_14584,N_12661);
nand UO_305 (O_305,N_14481,N_13508);
nor UO_306 (O_306,N_13681,N_12392);
and UO_307 (O_307,N_12072,N_13959);
and UO_308 (O_308,N_13722,N_13266);
and UO_309 (O_309,N_14683,N_13744);
or UO_310 (O_310,N_12755,N_13805);
nor UO_311 (O_311,N_12428,N_13791);
xor UO_312 (O_312,N_12883,N_12902);
nor UO_313 (O_313,N_14930,N_14820);
and UO_314 (O_314,N_14829,N_14132);
and UO_315 (O_315,N_14551,N_14430);
or UO_316 (O_316,N_14454,N_12125);
nor UO_317 (O_317,N_14808,N_12213);
or UO_318 (O_318,N_13228,N_14401);
nand UO_319 (O_319,N_12146,N_14807);
and UO_320 (O_320,N_12418,N_13294);
and UO_321 (O_321,N_13593,N_14206);
nand UO_322 (O_322,N_14881,N_12888);
and UO_323 (O_323,N_13275,N_13732);
nand UO_324 (O_324,N_14769,N_12412);
nor UO_325 (O_325,N_13291,N_13035);
and UO_326 (O_326,N_13412,N_13025);
nor UO_327 (O_327,N_13153,N_13246);
nor UO_328 (O_328,N_12063,N_13097);
nor UO_329 (O_329,N_12980,N_12522);
and UO_330 (O_330,N_13631,N_13451);
nor UO_331 (O_331,N_12983,N_14863);
nand UO_332 (O_332,N_12956,N_12539);
nand UO_333 (O_333,N_13860,N_13877);
xnor UO_334 (O_334,N_14974,N_13729);
xnor UO_335 (O_335,N_13057,N_12096);
nand UO_336 (O_336,N_12273,N_12062);
or UO_337 (O_337,N_12829,N_12193);
or UO_338 (O_338,N_12679,N_14987);
or UO_339 (O_339,N_13438,N_14711);
and UO_340 (O_340,N_14398,N_13262);
xor UO_341 (O_341,N_14878,N_13471);
or UO_342 (O_342,N_13338,N_12040);
or UO_343 (O_343,N_12970,N_14412);
or UO_344 (O_344,N_12700,N_13624);
nand UO_345 (O_345,N_13520,N_12202);
or UO_346 (O_346,N_13881,N_13052);
and UO_347 (O_347,N_13401,N_14857);
nor UO_348 (O_348,N_14163,N_13315);
and UO_349 (O_349,N_12367,N_14569);
nor UO_350 (O_350,N_14274,N_13033);
nor UO_351 (O_351,N_14242,N_12438);
nor UO_352 (O_352,N_13893,N_14883);
xor UO_353 (O_353,N_12799,N_12294);
nand UO_354 (O_354,N_13353,N_13669);
nor UO_355 (O_355,N_12907,N_14731);
and UO_356 (O_356,N_14495,N_14473);
nor UO_357 (O_357,N_13666,N_12291);
nor UO_358 (O_358,N_13470,N_14988);
and UO_359 (O_359,N_13506,N_13641);
or UO_360 (O_360,N_14748,N_14148);
and UO_361 (O_361,N_12839,N_13428);
and UO_362 (O_362,N_13099,N_12306);
and UO_363 (O_363,N_13786,N_13190);
nor UO_364 (O_364,N_12553,N_14289);
nor UO_365 (O_365,N_13340,N_12158);
nand UO_366 (O_366,N_12195,N_13882);
and UO_367 (O_367,N_14426,N_13204);
nand UO_368 (O_368,N_13561,N_13695);
nand UO_369 (O_369,N_14225,N_13354);
xnor UO_370 (O_370,N_12640,N_13939);
nor UO_371 (O_371,N_12256,N_13616);
or UO_372 (O_372,N_12217,N_13858);
or UO_373 (O_373,N_12757,N_14471);
xor UO_374 (O_374,N_12748,N_14329);
or UO_375 (O_375,N_12236,N_12998);
nor UO_376 (O_376,N_13001,N_13948);
and UO_377 (O_377,N_13154,N_12874);
xnor UO_378 (O_378,N_12567,N_14629);
xnor UO_379 (O_379,N_12132,N_12851);
or UO_380 (O_380,N_13018,N_12586);
nor UO_381 (O_381,N_14119,N_14766);
or UO_382 (O_382,N_13473,N_13140);
nand UO_383 (O_383,N_14406,N_12866);
nand UO_384 (O_384,N_14523,N_14209);
nand UO_385 (O_385,N_12834,N_13465);
and UO_386 (O_386,N_14060,N_12571);
xor UO_387 (O_387,N_12953,N_12552);
or UO_388 (O_388,N_13811,N_12993);
nand UO_389 (O_389,N_13373,N_13436);
or UO_390 (O_390,N_14271,N_14049);
nand UO_391 (O_391,N_14725,N_14682);
and UO_392 (O_392,N_12289,N_12315);
xnor UO_393 (O_393,N_12614,N_14452);
and UO_394 (O_394,N_12720,N_13420);
nand UO_395 (O_395,N_14439,N_14239);
nor UO_396 (O_396,N_13672,N_13381);
nor UO_397 (O_397,N_12328,N_12881);
xor UO_398 (O_398,N_13859,N_13539);
nor UO_399 (O_399,N_14804,N_13986);
xnor UO_400 (O_400,N_14760,N_14757);
and UO_401 (O_401,N_13039,N_13053);
or UO_402 (O_402,N_14330,N_12535);
or UO_403 (O_403,N_13331,N_13841);
nor UO_404 (O_404,N_14313,N_14325);
xnor UO_405 (O_405,N_12126,N_12118);
nor UO_406 (O_406,N_14538,N_12541);
xnor UO_407 (O_407,N_14858,N_12237);
nor UO_408 (O_408,N_12088,N_14056);
nor UO_409 (O_409,N_13464,N_14345);
nand UO_410 (O_410,N_13586,N_12654);
or UO_411 (O_411,N_13043,N_13332);
and UO_412 (O_412,N_14644,N_14656);
or UO_413 (O_413,N_14954,N_14346);
nand UO_414 (O_414,N_12737,N_14583);
and UO_415 (O_415,N_13622,N_13084);
nor UO_416 (O_416,N_13998,N_12354);
xnor UO_417 (O_417,N_12164,N_14096);
nor UO_418 (O_418,N_13573,N_12050);
or UO_419 (O_419,N_14503,N_12684);
nor UO_420 (O_420,N_14038,N_14496);
nand UO_421 (O_421,N_12372,N_12835);
nand UO_422 (O_422,N_12104,N_12718);
and UO_423 (O_423,N_14612,N_13950);
and UO_424 (O_424,N_14500,N_13565);
and UO_425 (O_425,N_14186,N_13640);
or UO_426 (O_426,N_13313,N_12934);
nand UO_427 (O_427,N_14681,N_14277);
and UO_428 (O_428,N_12454,N_14570);
and UO_429 (O_429,N_13365,N_13502);
nor UO_430 (O_430,N_12765,N_12989);
xor UO_431 (O_431,N_12321,N_14141);
nand UO_432 (O_432,N_14975,N_12384);
nor UO_433 (O_433,N_12391,N_14579);
nor UO_434 (O_434,N_13243,N_13289);
or UO_435 (O_435,N_13186,N_12169);
nand UO_436 (O_436,N_13267,N_14940);
xor UO_437 (O_437,N_13247,N_14397);
or UO_438 (O_438,N_14112,N_12319);
or UO_439 (O_439,N_14202,N_12855);
and UO_440 (O_440,N_13850,N_14825);
nand UO_441 (O_441,N_14125,N_14697);
or UO_442 (O_442,N_12060,N_14391);
and UO_443 (O_443,N_14642,N_12069);
nand UO_444 (O_444,N_13490,N_12672);
nor UO_445 (O_445,N_14968,N_14782);
or UO_446 (O_446,N_13026,N_14704);
and UO_447 (O_447,N_14502,N_13162);
nor UO_448 (O_448,N_14911,N_13062);
nand UO_449 (O_449,N_13836,N_12995);
xor UO_450 (O_450,N_12681,N_13503);
or UO_451 (O_451,N_12926,N_14574);
and UO_452 (O_452,N_12514,N_14705);
and UO_453 (O_453,N_13107,N_13951);
nor UO_454 (O_454,N_12485,N_14812);
nor UO_455 (O_455,N_12622,N_14917);
or UO_456 (O_456,N_12820,N_13969);
and UO_457 (O_457,N_14118,N_13581);
and UO_458 (O_458,N_12642,N_12906);
or UO_459 (O_459,N_12112,N_13071);
and UO_460 (O_460,N_14866,N_13976);
nor UO_461 (O_461,N_14967,N_13280);
or UO_462 (O_462,N_12831,N_12999);
nand UO_463 (O_463,N_14541,N_12964);
xor UO_464 (O_464,N_14789,N_12277);
xor UO_465 (O_465,N_14969,N_13578);
or UO_466 (O_466,N_14438,N_12383);
and UO_467 (O_467,N_12143,N_14130);
nor UO_468 (O_468,N_13359,N_12254);
and UO_469 (O_469,N_13838,N_14545);
nand UO_470 (O_470,N_13603,N_13540);
nand UO_471 (O_471,N_12070,N_12908);
or UO_472 (O_472,N_14064,N_14771);
and UO_473 (O_473,N_13292,N_14684);
or UO_474 (O_474,N_13674,N_14081);
and UO_475 (O_475,N_14357,N_14104);
or UO_476 (O_476,N_12747,N_13601);
nand UO_477 (O_477,N_14175,N_12460);
or UO_478 (O_478,N_13265,N_14476);
nor UO_479 (O_479,N_14722,N_14699);
nand UO_480 (O_480,N_14730,N_13521);
and UO_481 (O_481,N_12423,N_14768);
and UO_482 (O_482,N_13453,N_14332);
and UO_483 (O_483,N_12445,N_14609);
nand UO_484 (O_484,N_13363,N_13662);
nand UO_485 (O_485,N_12105,N_13128);
nand UO_486 (O_486,N_13284,N_14896);
nand UO_487 (O_487,N_12309,N_13005);
xor UO_488 (O_488,N_14814,N_12618);
nand UO_489 (O_489,N_13205,N_12653);
nor UO_490 (O_490,N_12606,N_14059);
nor UO_491 (O_491,N_14213,N_14506);
nor UO_492 (O_492,N_13861,N_12729);
or UO_493 (O_493,N_12744,N_14220);
or UO_494 (O_494,N_13772,N_12285);
and UO_495 (O_495,N_13733,N_13455);
or UO_496 (O_496,N_14340,N_14309);
and UO_497 (O_497,N_14797,N_13106);
and UO_498 (O_498,N_13226,N_12848);
or UO_499 (O_499,N_12887,N_12353);
nor UO_500 (O_500,N_13833,N_13421);
nor UO_501 (O_501,N_13476,N_13779);
and UO_502 (O_502,N_14263,N_13314);
or UO_503 (O_503,N_12260,N_13919);
or UO_504 (O_504,N_14390,N_13856);
xor UO_505 (O_505,N_14690,N_13857);
nor UO_506 (O_506,N_13251,N_13298);
or UO_507 (O_507,N_12192,N_13546);
nand UO_508 (O_508,N_13175,N_13989);
nand UO_509 (O_509,N_13454,N_13279);
xnor UO_510 (O_510,N_14404,N_14936);
or UO_511 (O_511,N_12078,N_12074);
nor UO_512 (O_512,N_13178,N_12356);
nand UO_513 (O_513,N_13689,N_14552);
nand UO_514 (O_514,N_12933,N_12965);
nand UO_515 (O_515,N_13582,N_12693);
or UO_516 (O_516,N_13120,N_12620);
nor UO_517 (O_517,N_14686,N_13032);
or UO_518 (O_518,N_14253,N_12843);
xor UO_519 (O_519,N_12865,N_12937);
and UO_520 (O_520,N_12345,N_13609);
and UO_521 (O_521,N_12882,N_12467);
nor UO_522 (O_522,N_14727,N_14300);
or UO_523 (O_523,N_13611,N_12741);
and UO_524 (O_524,N_14924,N_14991);
nor UO_525 (O_525,N_13745,N_12442);
nand UO_526 (O_526,N_12399,N_13768);
or UO_527 (O_527,N_13238,N_12214);
and UO_528 (O_528,N_12487,N_12600);
and UO_529 (O_529,N_14121,N_12470);
and UO_530 (O_530,N_13263,N_12004);
and UO_531 (O_531,N_13617,N_14734);
nor UO_532 (O_532,N_13364,N_13574);
nand UO_533 (O_533,N_14619,N_14367);
or UO_534 (O_534,N_12911,N_12705);
or UO_535 (O_535,N_14635,N_12030);
and UO_536 (O_536,N_13965,N_13036);
and UO_537 (O_537,N_14664,N_12106);
nor UO_538 (O_538,N_14604,N_13958);
and UO_539 (O_539,N_14278,N_13723);
nand UO_540 (O_540,N_14869,N_13917);
and UO_541 (O_541,N_12641,N_14752);
and UO_542 (O_542,N_12579,N_12630);
nor UO_543 (O_543,N_12708,N_14767);
nand UO_544 (O_544,N_13368,N_13563);
nor UO_545 (O_545,N_12206,N_13160);
and UO_546 (O_546,N_13417,N_13864);
nand UO_547 (O_547,N_12284,N_14714);
or UO_548 (O_548,N_12026,N_14795);
nor UO_549 (O_549,N_14611,N_13334);
nand UO_550 (O_550,N_12701,N_14620);
and UO_551 (O_551,N_12035,N_13575);
or UO_552 (O_552,N_14444,N_14221);
xnor UO_553 (O_553,N_12611,N_13975);
nor UO_554 (O_554,N_12676,N_14607);
nand UO_555 (O_555,N_13346,N_12978);
or UO_556 (O_556,N_12407,N_12667);
or UO_557 (O_557,N_12919,N_12927);
nor UO_558 (O_558,N_13536,N_14238);
nand UO_559 (O_559,N_12346,N_13347);
nor UO_560 (O_560,N_14255,N_12696);
xor UO_561 (O_561,N_12669,N_14566);
or UO_562 (O_562,N_13188,N_14166);
or UO_563 (O_563,N_12805,N_13687);
nand UO_564 (O_564,N_12509,N_12107);
and UO_565 (O_565,N_14252,N_13993);
nor UO_566 (O_566,N_13828,N_14575);
nand UO_567 (O_567,N_13065,N_13519);
or UO_568 (O_568,N_14114,N_14855);
nand UO_569 (O_569,N_12819,N_14986);
and UO_570 (O_570,N_13233,N_12131);
nor UO_571 (O_571,N_12262,N_12316);
nor UO_572 (O_572,N_12194,N_14074);
or UO_573 (O_573,N_13255,N_13234);
and UO_574 (O_574,N_14409,N_14673);
nor UO_575 (O_575,N_14429,N_13187);
xnor UO_576 (O_576,N_13088,N_12603);
or UO_577 (O_577,N_12601,N_13596);
nor UO_578 (O_578,N_12633,N_13961);
nor UO_579 (O_579,N_14640,N_14806);
xnor UO_580 (O_580,N_14169,N_13931);
and UO_581 (O_581,N_12918,N_14173);
nand UO_582 (O_582,N_12761,N_12613);
xor UO_583 (O_583,N_13325,N_14892);
and UO_584 (O_584,N_12732,N_14078);
xor UO_585 (O_585,N_13865,N_12022);
nand UO_586 (O_586,N_13599,N_13758);
nor UO_587 (O_587,N_14587,N_12124);
xor UO_588 (O_588,N_14933,N_14973);
or UO_589 (O_589,N_12930,N_12734);
and UO_590 (O_590,N_12738,N_14469);
nor UO_591 (O_591,N_12595,N_12129);
or UO_592 (O_592,N_14661,N_14085);
and UO_593 (O_593,N_14211,N_12283);
or UO_594 (O_594,N_13826,N_13901);
nand UO_595 (O_595,N_12574,N_13063);
and UO_596 (O_596,N_12893,N_14718);
xor UO_597 (O_597,N_14267,N_12537);
and UO_598 (O_598,N_13414,N_14772);
nand UO_599 (O_599,N_13542,N_12617);
xor UO_600 (O_600,N_13432,N_14904);
and UO_601 (O_601,N_13244,N_12296);
or UO_602 (O_602,N_12540,N_12904);
nand UO_603 (O_603,N_12564,N_13874);
nor UO_604 (O_604,N_14154,N_12665);
nor UO_605 (O_605,N_12864,N_14417);
nor UO_606 (O_606,N_12361,N_14403);
nand UO_607 (O_607,N_13398,N_12735);
xor UO_608 (O_608,N_13248,N_14365);
or UO_609 (O_609,N_13463,N_12625);
nand UO_610 (O_610,N_14565,N_12643);
xnor UO_611 (O_611,N_12006,N_12015);
xor UO_612 (O_612,N_14625,N_14160);
nor UO_613 (O_613,N_14913,N_13773);
xnor UO_614 (O_614,N_14677,N_12636);
and UO_615 (O_615,N_13343,N_12982);
and UO_616 (O_616,N_12420,N_14269);
or UO_617 (O_617,N_14022,N_14199);
nor UO_618 (O_618,N_14744,N_14307);
and UO_619 (O_619,N_14053,N_14162);
or UO_620 (O_620,N_13552,N_14737);
or UO_621 (O_621,N_13627,N_14020);
and UO_622 (O_622,N_14423,N_14937);
nor UO_623 (O_623,N_13232,N_14088);
nand UO_624 (O_624,N_14327,N_12475);
nor UO_625 (O_625,N_13061,N_14946);
nor UO_626 (O_626,N_12056,N_12488);
and UO_627 (O_627,N_12374,N_13049);
or UO_628 (O_628,N_12895,N_13342);
xor UO_629 (O_629,N_14547,N_14675);
nor UO_630 (O_630,N_12244,N_12292);
nand UO_631 (O_631,N_13512,N_13580);
xor UO_632 (O_632,N_14898,N_12833);
nand UO_633 (O_633,N_13557,N_14596);
nor UO_634 (O_634,N_14606,N_12246);
or UO_635 (O_635,N_14849,N_12928);
nor UO_636 (O_636,N_12029,N_12524);
or UO_637 (O_637,N_12259,N_13224);
xnor UO_638 (O_638,N_12612,N_13174);
and UO_639 (O_639,N_14031,N_14029);
nor UO_640 (O_640,N_13528,N_12263);
or UO_641 (O_641,N_13221,N_13900);
nand UO_642 (O_642,N_12341,N_12135);
nor UO_643 (O_643,N_14702,N_13059);
xnor UO_644 (O_644,N_13497,N_13308);
nor UO_645 (O_645,N_13818,N_13358);
or UO_646 (O_646,N_14351,N_12496);
or UO_647 (O_647,N_14665,N_12814);
nand UO_648 (O_648,N_13029,N_13367);
nor UO_649 (O_649,N_13907,N_12812);
or UO_650 (O_650,N_12714,N_13844);
and UO_651 (O_651,N_14781,N_12890);
xnor UO_652 (O_652,N_14408,N_14553);
nor UO_653 (O_653,N_12066,N_12330);
nor UO_654 (O_654,N_13477,N_13849);
nand UO_655 (O_655,N_14799,N_13064);
or UO_656 (O_656,N_12561,N_13785);
nor UO_657 (O_657,N_14810,N_12021);
nand UO_658 (O_658,N_13400,N_13970);
nand UO_659 (O_659,N_12530,N_12240);
and UO_660 (O_660,N_14250,N_12033);
nor UO_661 (O_661,N_14867,N_12358);
or UO_662 (O_662,N_13102,N_13932);
or UO_663 (O_663,N_12527,N_14318);
and UO_664 (O_664,N_13474,N_13764);
and UO_665 (O_665,N_14215,N_12677);
or UO_666 (O_666,N_14407,N_13416);
and UO_667 (O_667,N_14167,N_12599);
and UO_668 (O_668,N_12338,N_13090);
nor UO_669 (O_669,N_13878,N_14608);
and UO_670 (O_670,N_13604,N_13069);
xnor UO_671 (O_671,N_14431,N_14876);
xor UO_672 (O_672,N_13264,N_13485);
and UO_673 (O_673,N_12087,N_12229);
and UO_674 (O_674,N_12860,N_13914);
nand UO_675 (O_675,N_12079,N_12656);
nor UO_676 (O_676,N_13753,N_14498);
nand UO_677 (O_677,N_12077,N_13550);
and UO_678 (O_678,N_13794,N_14485);
and UO_679 (O_679,N_13278,N_14827);
nor UO_680 (O_680,N_14262,N_12502);
nand UO_681 (O_681,N_12516,N_14902);
and UO_682 (O_682,N_12427,N_13379);
nand UO_683 (O_683,N_13781,N_12089);
and UO_684 (O_684,N_13482,N_14755);
and UO_685 (O_685,N_13330,N_13964);
nor UO_686 (O_686,N_12377,N_12783);
nor UO_687 (O_687,N_12177,N_14868);
and UO_688 (O_688,N_13151,N_13801);
nor UO_689 (O_689,N_14280,N_12879);
xor UO_690 (O_690,N_12133,N_13823);
and UO_691 (O_691,N_13620,N_13457);
nor UO_692 (O_692,N_14953,N_13460);
xor UO_693 (O_693,N_14360,N_13276);
nor UO_694 (O_694,N_13782,N_14504);
xnor UO_695 (O_695,N_13252,N_14433);
nor UO_696 (O_696,N_14676,N_12559);
or UO_697 (O_697,N_12652,N_12662);
nand UO_698 (O_698,N_14270,N_13804);
and UO_699 (O_699,N_12093,N_14990);
nor UO_700 (O_700,N_13362,N_14529);
or UO_701 (O_701,N_13037,N_14623);
or UO_702 (O_702,N_14413,N_14461);
and UO_703 (O_703,N_14695,N_14490);
nor UO_704 (O_704,N_12668,N_13013);
nand UO_705 (O_705,N_12268,N_14122);
and UO_706 (O_706,N_14363,N_14386);
xnor UO_707 (O_707,N_12635,N_14111);
or UO_708 (O_708,N_13543,N_14512);
or UO_709 (O_709,N_13183,N_13237);
or UO_710 (O_710,N_13126,N_12597);
nor UO_711 (O_711,N_13665,N_13329);
xor UO_712 (O_712,N_14294,N_14012);
and UO_713 (O_713,N_13431,N_12857);
or UO_714 (O_714,N_14836,N_13769);
xnor UO_715 (O_715,N_13443,N_12247);
or UO_716 (O_716,N_14582,N_12778);
and UO_717 (O_717,N_14067,N_14918);
nand UO_718 (O_718,N_13840,N_12140);
xnor UO_719 (O_719,N_14657,N_12117);
and UO_720 (O_720,N_13632,N_12144);
nand UO_721 (O_721,N_14728,N_12565);
and UO_722 (O_722,N_14435,N_12782);
and UO_723 (O_723,N_13370,N_13717);
and UO_724 (O_724,N_12711,N_14713);
or UO_725 (O_725,N_12153,N_13446);
or UO_726 (O_726,N_14205,N_14685);
nand UO_727 (O_727,N_14483,N_12436);
or UO_728 (O_728,N_14689,N_13336);
and UO_729 (O_729,N_13891,N_13288);
and UO_730 (O_730,N_13777,N_12996);
nand UO_731 (O_731,N_14801,N_12873);
nand UO_732 (O_732,N_14484,N_14359);
or UO_733 (O_733,N_13647,N_13198);
and UO_734 (O_734,N_14909,N_14951);
nor UO_735 (O_735,N_14501,N_14129);
xor UO_736 (O_736,N_13809,N_14079);
or UO_737 (O_737,N_13091,N_14505);
or UO_738 (O_738,N_12786,N_12913);
and UO_739 (O_739,N_12458,N_12139);
or UO_740 (O_740,N_13389,N_12108);
nor UO_741 (O_741,N_12792,N_14751);
or UO_742 (O_742,N_14568,N_14632);
nor UO_743 (O_743,N_13634,N_12638);
nand UO_744 (O_744,N_12119,N_14004);
and UO_745 (O_745,N_14174,N_12929);
nor UO_746 (O_746,N_14043,N_12825);
and UO_747 (O_747,N_12299,N_14287);
and UO_748 (O_748,N_14198,N_13906);
nor UO_749 (O_749,N_14630,N_12390);
and UO_750 (O_750,N_14017,N_12424);
nand UO_751 (O_751,N_14187,N_13629);
nand UO_752 (O_752,N_14016,N_13748);
nand UO_753 (O_753,N_14249,N_13671);
or UO_754 (O_754,N_14048,N_13731);
nand UO_755 (O_755,N_12975,N_12914);
or UO_756 (O_756,N_14610,N_12529);
or UO_757 (O_757,N_14941,N_13977);
nor UO_758 (O_758,N_12660,N_13583);
nor UO_759 (O_759,N_14035,N_13988);
nor UO_760 (O_760,N_14063,N_14962);
xnor UO_761 (O_761,N_14897,N_14315);
and UO_762 (O_762,N_14072,N_12416);
nand UO_763 (O_763,N_14550,N_14055);
or UO_764 (O_764,N_12203,N_14131);
nand UO_765 (O_765,N_13747,N_12141);
nor UO_766 (O_766,N_12261,N_12136);
xnor UO_767 (O_767,N_14717,N_14358);
nand UO_768 (O_768,N_14158,N_13418);
and UO_769 (O_769,N_13784,N_12555);
or UO_770 (O_770,N_13268,N_14190);
nor UO_771 (O_771,N_12160,N_14051);
or UO_772 (O_772,N_13776,N_14319);
and UO_773 (O_773,N_14648,N_13619);
and UO_774 (O_774,N_13890,N_14384);
and UO_775 (O_775,N_12828,N_13905);
and UO_776 (O_776,N_14292,N_12773);
nor UO_777 (O_777,N_14948,N_13771);
nand UO_778 (O_778,N_12632,N_12250);
or UO_779 (O_779,N_14666,N_12478);
xnor UO_780 (O_780,N_13646,N_14624);
nor UO_781 (O_781,N_13366,N_13253);
nand UO_782 (O_782,N_12279,N_13514);
nor UO_783 (O_783,N_13475,N_14176);
and UO_784 (O_784,N_13949,N_12499);
or UO_785 (O_785,N_13213,N_14788);
nor UO_786 (O_786,N_12371,N_13390);
nor UO_787 (O_787,N_13486,N_14256);
nand UO_788 (O_788,N_12249,N_13283);
nand UO_789 (O_789,N_12064,N_13716);
nand UO_790 (O_790,N_14299,N_12304);
nor UO_791 (O_791,N_12543,N_13642);
and UO_792 (O_792,N_12186,N_14517);
nand UO_793 (O_793,N_13301,N_12759);
or UO_794 (O_794,N_14845,N_14521);
nor UO_795 (O_795,N_14680,N_13556);
or UO_796 (O_796,N_14254,N_14709);
xnor UO_797 (O_797,N_13240,N_12771);
nand UO_798 (O_798,N_12355,N_13774);
or UO_799 (O_799,N_13300,N_13670);
nor UO_800 (O_800,N_13274,N_14742);
nand UO_801 (O_801,N_14985,N_13108);
nor UO_802 (O_802,N_14674,N_13038);
nor UO_803 (O_803,N_13022,N_12215);
and UO_804 (O_804,N_13212,N_12538);
or UO_805 (O_805,N_12433,N_14115);
or UO_806 (O_806,N_14188,N_13708);
nor UO_807 (O_807,N_12958,N_13339);
nor UO_808 (O_808,N_14191,N_13741);
nand UO_809 (O_809,N_14787,N_13208);
nor UO_810 (O_810,N_13478,N_12544);
and UO_811 (O_811,N_14534,N_12168);
nor UO_812 (O_812,N_14046,N_12592);
nand UO_813 (O_813,N_12626,N_12616);
nand UO_814 (O_814,N_12161,N_13819);
or UO_815 (O_815,N_12426,N_14966);
and UO_816 (O_816,N_13488,N_12253);
nand UO_817 (O_817,N_12589,N_12084);
and UO_818 (O_818,N_13319,N_13750);
nor UO_819 (O_819,N_13902,N_13158);
or UO_820 (O_820,N_13661,N_13740);
and UO_821 (O_821,N_13127,N_12255);
or UO_822 (O_822,N_13511,N_12510);
nand UO_823 (O_823,N_12476,N_12912);
and UO_824 (O_824,N_13050,N_13074);
and UO_825 (O_825,N_12666,N_12200);
xnor UO_826 (O_826,N_14847,N_13994);
nor UO_827 (O_827,N_13655,N_12957);
xnor UO_828 (O_828,N_14207,N_12332);
nand UO_829 (O_829,N_14480,N_14229);
nand UO_830 (O_830,N_14785,N_12429);
nor UO_831 (O_831,N_14536,N_12474);
and UO_832 (O_832,N_14475,N_13572);
nand UO_833 (O_833,N_12802,N_14576);
nor UO_834 (O_834,N_12823,N_12290);
nor UO_835 (O_835,N_12447,N_14142);
nand UO_836 (O_836,N_14877,N_14907);
xor UO_837 (O_837,N_14759,N_12410);
or UO_838 (O_838,N_14696,N_14233);
nor UO_839 (O_839,N_12266,N_14732);
nor UO_840 (O_840,N_14062,N_13806);
or UO_841 (O_841,N_13499,N_12569);
nor UO_842 (O_842,N_14113,N_12425);
nand UO_843 (O_843,N_13382,N_13242);
nor UO_844 (O_844,N_14934,N_12534);
or UO_845 (O_845,N_14244,N_14275);
or UO_846 (O_846,N_14996,N_12659);
nor UO_847 (O_847,N_12979,N_14449);
or UO_848 (O_848,N_14260,N_14381);
nand UO_849 (O_849,N_13927,N_12988);
and UO_850 (O_850,N_13531,N_13664);
xor UO_851 (O_851,N_12068,N_14703);
nand UO_852 (O_852,N_14389,N_14375);
and UO_853 (O_853,N_14694,N_12440);
nor UO_854 (O_854,N_12878,N_12837);
or UO_855 (O_855,N_12818,N_13752);
and UO_856 (O_856,N_14915,N_12859);
nor UO_857 (O_857,N_12897,N_14054);
xor UO_858 (O_858,N_14976,N_12756);
nor UO_859 (O_859,N_12437,N_12501);
xor UO_860 (O_860,N_12180,N_12446);
or UO_861 (O_861,N_12585,N_12699);
xor UO_862 (O_862,N_13524,N_12932);
or UO_863 (O_863,N_13657,N_12310);
nand UO_864 (O_864,N_12832,N_13825);
nor UO_865 (O_865,N_14856,N_12142);
or UO_866 (O_866,N_13981,N_12686);
nor UO_867 (O_867,N_14980,N_12885);
nor UO_868 (O_868,N_12167,N_12145);
nor UO_869 (O_869,N_12404,N_14099);
or UO_870 (O_870,N_12324,N_13855);
and UO_871 (O_871,N_12558,N_14040);
and UO_872 (O_872,N_12486,N_12090);
nand UO_873 (O_873,N_12811,N_14573);
or UO_874 (O_874,N_14572,N_13163);
and UO_875 (O_875,N_12269,N_14235);
or UO_876 (O_876,N_12985,N_14424);
xor UO_877 (O_877,N_12342,N_12080);
nor UO_878 (O_878,N_14773,N_13875);
or UO_879 (O_879,N_13286,N_14528);
nand UO_880 (O_880,N_13372,N_12774);
nor UO_881 (O_881,N_13217,N_14488);
nor UO_882 (O_882,N_14443,N_14463);
and UO_883 (O_883,N_12128,N_12637);
xnor UO_884 (O_884,N_14177,N_12872);
or UO_885 (O_885,N_12032,N_13498);
and UO_886 (O_886,N_12380,N_12449);
or UO_887 (O_887,N_12045,N_13173);
nor UO_888 (O_888,N_13146,N_14455);
xor UO_889 (O_889,N_14961,N_14803);
or UO_890 (O_890,N_12960,N_14802);
and UO_891 (O_891,N_14147,N_14465);
or UO_892 (O_892,N_12387,N_12967);
or UO_893 (O_893,N_14761,N_13648);
xnor UO_894 (O_894,N_13739,N_13710);
nand UO_895 (O_895,N_12824,N_13351);
nand UO_896 (O_896,N_12274,N_14720);
or UO_897 (O_897,N_13697,N_14809);
nor UO_898 (O_898,N_13889,N_14548);
nor UO_899 (O_899,N_13886,N_14850);
xor UO_900 (O_900,N_12459,N_12251);
nor UO_901 (O_901,N_12199,N_12624);
and UO_902 (O_902,N_14687,N_14577);
or UO_903 (O_903,N_13410,N_14080);
nand UO_904 (O_904,N_14647,N_14246);
nor UO_905 (O_905,N_14086,N_14908);
nor UO_906 (O_906,N_14590,N_13424);
and UO_907 (O_907,N_13820,N_14972);
nor UO_908 (O_908,N_12395,N_14710);
nand UO_909 (O_909,N_13667,N_14379);
or UO_910 (O_910,N_12357,N_12822);
or UO_911 (O_911,N_12333,N_13089);
nand UO_912 (O_912,N_14817,N_12233);
xor UO_913 (O_913,N_12191,N_13348);
nand UO_914 (O_914,N_14032,N_14589);
and UO_915 (O_915,N_12924,N_12110);
or UO_916 (O_916,N_13448,N_13098);
nor UO_917 (O_917,N_14100,N_12212);
or UO_918 (O_918,N_13079,N_14005);
nor UO_919 (O_919,N_13558,N_13780);
xor UO_920 (O_920,N_13139,N_14777);
nand UO_921 (O_921,N_13015,N_12058);
and UO_922 (O_922,N_12969,N_12227);
nand UO_923 (O_923,N_13694,N_13645);
nor UO_924 (O_924,N_13713,N_13101);
nand UO_925 (O_925,N_14507,N_14754);
nand UO_926 (O_926,N_12862,N_12695);
nand UO_927 (O_927,N_12889,N_12629);
xnor UO_928 (O_928,N_12663,N_14786);
nor UO_929 (O_929,N_14486,N_13829);
nor UO_930 (O_930,N_13369,N_13103);
or UO_931 (O_931,N_12706,N_14819);
nor UO_932 (O_932,N_12008,N_13654);
nand UO_933 (O_933,N_14094,N_12219);
and UO_934 (O_934,N_12789,N_14952);
or UO_935 (O_935,N_12323,N_13356);
and UO_936 (O_936,N_13895,N_13357);
and UO_937 (O_937,N_14436,N_12769);
or UO_938 (O_938,N_14083,N_14712);
or UO_939 (O_939,N_13027,N_14288);
nand UO_940 (O_940,N_12847,N_14396);
or UO_941 (O_941,N_13355,N_14950);
nand UO_942 (O_942,N_13159,N_13405);
nor UO_943 (O_943,N_13533,N_14298);
nor UO_944 (O_944,N_12243,N_14457);
and UO_945 (O_945,N_13215,N_14382);
nor UO_946 (O_946,N_13501,N_13912);
nor UO_947 (O_947,N_14497,N_12948);
and UO_948 (O_948,N_12305,N_13361);
nand UO_949 (O_949,N_14352,N_12609);
nor UO_950 (O_950,N_13759,N_12462);
and UO_951 (O_951,N_12517,N_12054);
nor UO_952 (O_952,N_12657,N_14838);
nand UO_953 (O_953,N_13936,N_14165);
or UO_954 (O_954,N_12968,N_12602);
nor UO_955 (O_955,N_14774,N_14571);
nand UO_956 (O_956,N_14743,N_12170);
and UO_957 (O_957,N_13138,N_12584);
and UO_958 (O_958,N_14784,N_13754);
nor UO_959 (O_959,N_13967,N_13869);
and UO_960 (O_960,N_13095,N_14258);
and UO_961 (O_961,N_12492,N_14380);
nor UO_962 (O_962,N_13633,N_14314);
or UO_963 (O_963,N_14659,N_13211);
nand UO_964 (O_964,N_14873,N_14992);
and UO_965 (O_965,N_14108,N_14230);
and UO_966 (O_966,N_13795,N_14110);
nor UO_967 (O_967,N_12477,N_13076);
or UO_968 (O_968,N_13677,N_12508);
nor UO_969 (O_969,N_13048,N_13909);
or UO_970 (O_970,N_14442,N_13916);
and UO_971 (O_971,N_12302,N_12596);
or UO_972 (O_972,N_14172,N_14448);
or UO_973 (O_973,N_12511,N_12348);
nand UO_974 (O_974,N_13439,N_12023);
and UO_975 (O_975,N_14344,N_13702);
or UO_976 (O_976,N_14749,N_13579);
nand UO_977 (O_977,N_12621,N_12057);
nor UO_978 (O_978,N_14979,N_14633);
nand UO_979 (O_979,N_12515,N_14927);
nor UO_980 (O_980,N_12880,N_14222);
or UO_981 (O_981,N_12059,N_14791);
nand UO_982 (O_982,N_12300,N_13880);
and UO_983 (O_983,N_12687,N_13360);
nor UO_984 (O_984,N_13728,N_12910);
nand UO_985 (O_985,N_13911,N_13167);
nand UO_986 (O_986,N_14700,N_12148);
or UO_987 (O_987,N_13549,N_13047);
or UO_988 (O_988,N_14092,N_12547);
nand UO_989 (O_989,N_13888,N_12858);
and UO_990 (O_990,N_12287,N_13972);
nand UO_991 (O_991,N_14006,N_13973);
nand UO_992 (O_992,N_14535,N_12990);
xor UO_993 (O_993,N_14369,N_14920);
nor UO_994 (O_994,N_14021,N_14066);
or UO_995 (O_995,N_12347,N_13044);
xnor UO_996 (O_996,N_14516,N_12224);
nor UO_997 (O_997,N_12984,N_13971);
nand UO_998 (O_998,N_13845,N_14900);
nor UO_999 (O_999,N_13200,N_12573);
or UO_1000 (O_1000,N_12159,N_14420);
nand UO_1001 (O_1001,N_14425,N_12570);
nor UO_1002 (O_1002,N_14658,N_14018);
nand UO_1003 (O_1003,N_13679,N_12939);
and UO_1004 (O_1004,N_13333,N_14394);
nor UO_1005 (O_1005,N_12803,N_12417);
and UO_1006 (O_1006,N_14914,N_14628);
nor UO_1007 (O_1007,N_13068,N_13185);
and UO_1008 (O_1008,N_12278,N_13933);
or UO_1009 (O_1009,N_12551,N_12493);
and UO_1010 (O_1010,N_13137,N_13897);
nor UO_1011 (O_1011,N_12394,N_12375);
or UO_1012 (O_1012,N_14026,N_12122);
nor UO_1013 (O_1013,N_13172,N_13562);
nor UO_1014 (O_1014,N_14068,N_13853);
nand UO_1015 (O_1015,N_12034,N_14192);
nor UO_1016 (O_1016,N_13386,N_13147);
nor UO_1017 (O_1017,N_12047,N_12365);
and UO_1018 (O_1018,N_14445,N_13727);
nor UO_1019 (O_1019,N_14377,N_12712);
or UO_1020 (O_1020,N_13415,N_14852);
xnor UO_1021 (O_1021,N_13134,N_14155);
nand UO_1022 (O_1022,N_13003,N_12288);
or UO_1023 (O_1023,N_14245,N_13399);
or UO_1024 (O_1024,N_13960,N_12582);
nand UO_1025 (O_1025,N_13693,N_13207);
and UO_1026 (O_1026,N_13245,N_13010);
nor UO_1027 (O_1027,N_12742,N_12940);
nand UO_1028 (O_1028,N_13344,N_12892);
or UO_1029 (O_1029,N_13918,N_12875);
nand UO_1030 (O_1030,N_14667,N_12945);
nand UO_1031 (O_1031,N_14223,N_12311);
or UO_1032 (O_1032,N_14639,N_14540);
nor UO_1033 (O_1033,N_13293,N_12339);
nor UO_1034 (O_1034,N_14779,N_12166);
nand UO_1035 (O_1035,N_13045,N_13577);
xnor UO_1036 (O_1036,N_14958,N_13031);
nor UO_1037 (O_1037,N_14834,N_14324);
or UO_1038 (O_1038,N_13526,N_13197);
nor UO_1039 (O_1039,N_14701,N_13317);
nor UO_1040 (O_1040,N_14106,N_12397);
and UO_1041 (O_1041,N_13956,N_13427);
and UO_1042 (O_1042,N_12840,N_12877);
nand UO_1043 (O_1043,N_14034,N_12797);
or UO_1044 (O_1044,N_12223,N_13873);
nand UO_1045 (O_1045,N_12209,N_13652);
xnor UO_1046 (O_1046,N_14259,N_12489);
nand UO_1047 (O_1047,N_14923,N_12916);
nor UO_1048 (O_1048,N_13479,N_12127);
and UO_1049 (O_1049,N_14161,N_13979);
or UO_1050 (O_1050,N_13121,N_13770);
xor UO_1051 (O_1051,N_13724,N_12557);
or UO_1052 (O_1052,N_12265,N_13684);
or UO_1053 (O_1053,N_12484,N_13413);
and UO_1054 (O_1054,N_12876,N_13595);
nor UO_1055 (O_1055,N_13396,N_13649);
nand UO_1056 (O_1056,N_13584,N_13320);
or UO_1057 (O_1057,N_12020,N_13847);
and UO_1058 (O_1058,N_14865,N_13165);
or UO_1059 (O_1059,N_12336,N_12264);
xnor UO_1060 (O_1060,N_14672,N_14268);
or UO_1061 (O_1061,N_13002,N_13483);
nor UO_1062 (O_1062,N_13434,N_13810);
nor UO_1063 (O_1063,N_13614,N_13113);
nor UO_1064 (O_1064,N_12991,N_12232);
and UO_1065 (O_1065,N_14128,N_13324);
and UO_1066 (O_1066,N_13943,N_14841);
or UO_1067 (O_1067,N_12061,N_12276);
nor UO_1068 (O_1068,N_12781,N_12491);
nor UO_1069 (O_1069,N_12846,N_14945);
and UO_1070 (O_1070,N_12870,N_14025);
and UO_1071 (O_1071,N_14204,N_13925);
and UO_1072 (O_1072,N_14957,N_12113);
and UO_1073 (O_1073,N_12722,N_12450);
and UO_1074 (O_1074,N_14643,N_12899);
and UO_1075 (O_1075,N_13676,N_14939);
nand UO_1076 (O_1076,N_13765,N_14181);
nor UO_1077 (O_1077,N_14790,N_12370);
and UO_1078 (O_1078,N_13974,N_13491);
nand UO_1079 (O_1079,N_13349,N_14691);
nor UO_1080 (O_1080,N_12707,N_12313);
and UO_1081 (O_1081,N_14978,N_12673);
nor UO_1082 (O_1082,N_13518,N_13534);
nor UO_1083 (O_1083,N_12103,N_14555);
and UO_1084 (O_1084,N_14226,N_13124);
or UO_1085 (O_1085,N_14626,N_13726);
nand UO_1086 (O_1086,N_12753,N_13484);
nand UO_1087 (O_1087,N_13639,N_12009);
nor UO_1088 (O_1088,N_13335,N_13756);
nor UO_1089 (O_1089,N_14539,N_14669);
and UO_1090 (O_1090,N_14921,N_14460);
or UO_1091 (O_1091,N_13831,N_14197);
nand UO_1092 (O_1092,N_14084,N_14544);
nand UO_1093 (O_1093,N_13564,N_14514);
and UO_1094 (O_1094,N_13513,N_14563);
or UO_1095 (O_1095,N_12731,N_12176);
nor UO_1096 (O_1096,N_14103,N_12350);
and UO_1097 (O_1097,N_12776,N_12566);
nor UO_1098 (O_1098,N_13863,N_12580);
and UO_1099 (O_1099,N_14943,N_12435);
xor UO_1100 (O_1100,N_14000,N_13230);
and UO_1101 (O_1101,N_13675,N_12709);
nor UO_1102 (O_1102,N_13176,N_13735);
or UO_1103 (O_1103,N_14839,N_12542);
or UO_1104 (O_1104,N_12915,N_14912);
or UO_1105 (O_1105,N_14470,N_13225);
xnor UO_1106 (O_1106,N_12763,N_14105);
nand UO_1107 (O_1107,N_14349,N_14618);
or UO_1108 (O_1108,N_13592,N_13653);
or UO_1109 (O_1109,N_13898,N_14740);
xor UO_1110 (O_1110,N_13116,N_13554);
nor UO_1111 (O_1111,N_13493,N_13218);
nand UO_1112 (O_1112,N_13607,N_13843);
nand UO_1113 (O_1113,N_14284,N_13272);
and UO_1114 (O_1114,N_12082,N_14002);
xor UO_1115 (O_1115,N_12473,N_14822);
or UO_1116 (O_1116,N_13509,N_13612);
nand UO_1117 (O_1117,N_13602,N_12577);
and UO_1118 (O_1118,N_12275,N_13170);
or UO_1119 (O_1119,N_13870,N_13630);
nor UO_1120 (O_1120,N_13450,N_14057);
nand UO_1121 (O_1121,N_12075,N_13302);
nand UO_1122 (O_1122,N_14478,N_14543);
or UO_1123 (O_1123,N_13305,N_12065);
nand UO_1124 (O_1124,N_12779,N_13846);
and UO_1125 (O_1125,N_12697,N_14965);
and UO_1126 (O_1126,N_13223,N_12147);
nand UO_1127 (O_1127,N_13341,N_13009);
nand UO_1128 (O_1128,N_14376,N_12581);
xor UO_1129 (O_1129,N_14123,N_12385);
or UO_1130 (O_1130,N_14023,N_14668);
nand UO_1131 (O_1131,N_12523,N_14796);
nand UO_1132 (O_1132,N_13273,N_12005);
nor UO_1133 (O_1133,N_12730,N_12777);
xor UO_1134 (O_1134,N_12188,N_12444);
nor UO_1135 (O_1135,N_13594,N_12422);
and UO_1136 (O_1136,N_13887,N_13516);
or UO_1137 (O_1137,N_12850,N_14214);
or UO_1138 (O_1138,N_13610,N_13193);
and UO_1139 (O_1139,N_14266,N_13070);
nor UO_1140 (O_1140,N_14464,N_12619);
nand UO_1141 (O_1141,N_13751,N_13705);
nand UO_1142 (O_1142,N_13660,N_14427);
nor UO_1143 (O_1143,N_14562,N_12329);
or UO_1144 (O_1144,N_14441,N_13487);
or UO_1145 (O_1145,N_13148,N_13812);
nor UO_1146 (O_1146,N_12921,N_12655);
nor UO_1147 (O_1147,N_12011,N_13711);
and UO_1148 (O_1148,N_13532,N_12190);
xnor UO_1149 (O_1149,N_14095,N_13686);
nor UO_1150 (O_1150,N_12094,N_13408);
nor UO_1151 (O_1151,N_12352,N_14520);
and UO_1152 (O_1152,N_14310,N_13203);
nor UO_1153 (O_1153,N_13606,N_14033);
or UO_1154 (O_1154,N_14726,N_14846);
nand UO_1155 (O_1155,N_13195,N_12052);
and UO_1156 (O_1156,N_12307,N_12137);
or UO_1157 (O_1157,N_13157,N_13129);
or UO_1158 (O_1158,N_14558,N_13494);
nor UO_1159 (O_1159,N_14688,N_14052);
and UO_1160 (O_1160,N_12512,N_13164);
nor UO_1161 (O_1161,N_14758,N_13179);
nand UO_1162 (O_1162,N_13481,N_12479);
and UO_1163 (O_1163,N_14828,N_12856);
nand UO_1164 (O_1164,N_13371,N_12083);
or UO_1165 (O_1165,N_14853,N_12806);
nor UO_1166 (O_1166,N_14402,N_12154);
or UO_1167 (O_1167,N_12222,N_14627);
or UO_1168 (O_1168,N_13384,N_14493);
or UO_1169 (O_1169,N_13141,N_14193);
nor UO_1170 (O_1170,N_12780,N_12027);
xor UO_1171 (O_1171,N_13391,N_13525);
and UO_1172 (O_1172,N_14071,N_14770);
or UO_1173 (O_1173,N_12225,N_12181);
nand UO_1174 (O_1174,N_12922,N_14837);
nor UO_1175 (O_1175,N_14835,N_13796);
nor UO_1176 (O_1176,N_12376,N_14871);
and UO_1177 (O_1177,N_14652,N_13277);
nor UO_1178 (O_1178,N_13118,N_14692);
nand UO_1179 (O_1179,N_12466,N_13260);
nand UO_1180 (O_1180,N_13690,N_12674);
nand UO_1181 (O_1181,N_14894,N_12931);
nand UO_1182 (O_1182,N_13842,N_14719);
or UO_1183 (O_1183,N_13808,N_13523);
or UO_1184 (O_1184,N_14180,N_14477);
nand UO_1185 (O_1185,N_13042,N_12532);
nor UO_1186 (O_1186,N_13096,N_14366);
or UO_1187 (O_1187,N_12031,N_14164);
nand UO_1188 (O_1188,N_12456,N_14061);
nand UO_1189 (O_1189,N_13393,N_12972);
nand UO_1190 (O_1190,N_13626,N_14194);
or UO_1191 (O_1191,N_14650,N_12952);
and UO_1192 (O_1192,N_12455,N_12308);
nand UO_1193 (O_1193,N_14210,N_14884);
or UO_1194 (O_1194,N_13004,N_14089);
xor UO_1195 (O_1195,N_14041,N_14617);
nor UO_1196 (O_1196,N_12097,N_13872);
and UO_1197 (O_1197,N_14989,N_14437);
nor UO_1198 (O_1198,N_12962,N_12664);
nand UO_1199 (O_1199,N_12548,N_14009);
and UO_1200 (O_1200,N_14285,N_12295);
nand UO_1201 (O_1201,N_12704,N_14459);
nor UO_1202 (O_1202,N_14419,N_13083);
or UO_1203 (O_1203,N_12977,N_12816);
or UO_1204 (O_1204,N_14272,N_14456);
or UO_1205 (O_1205,N_13066,N_12795);
xor UO_1206 (O_1206,N_13117,N_12651);
or UO_1207 (O_1207,N_12702,N_13467);
nand UO_1208 (O_1208,N_14851,N_13862);
or UO_1209 (O_1209,N_12451,N_13034);
nor UO_1210 (O_1210,N_14024,N_14833);
or UO_1211 (O_1211,N_12942,N_12568);
or UO_1212 (O_1212,N_14762,N_14649);
or UO_1213 (O_1213,N_14282,N_12725);
and UO_1214 (O_1214,N_14885,N_13892);
and UO_1215 (O_1215,N_14286,N_12545);
and UO_1216 (O_1216,N_14723,N_13924);
nor UO_1217 (O_1217,N_14171,N_12003);
nand UO_1218 (O_1218,N_12067,N_12689);
or UO_1219 (O_1219,N_13257,N_12963);
and UO_1220 (O_1220,N_12464,N_12867);
nand UO_1221 (O_1221,N_12494,N_12138);
nor UO_1222 (O_1222,N_13730,N_13311);
or UO_1223 (O_1223,N_14127,N_12521);
nor UO_1224 (O_1224,N_12754,N_13555);
or UO_1225 (O_1225,N_13051,N_12165);
nand UO_1226 (O_1226,N_13761,N_12049);
xnor UO_1227 (O_1227,N_12055,N_12025);
xnor UO_1228 (O_1228,N_13866,N_12531);
nor UO_1229 (O_1229,N_12680,N_12441);
nor UO_1230 (O_1230,N_14410,N_13799);
and UO_1231 (O_1231,N_13608,N_12943);
and UO_1232 (O_1232,N_13299,N_12301);
and UO_1233 (O_1233,N_12842,N_14138);
and UO_1234 (O_1234,N_12018,N_14302);
and UO_1235 (O_1235,N_12997,N_14075);
nand UO_1236 (O_1236,N_12042,N_14432);
nand UO_1237 (O_1237,N_13322,N_13636);
xnor UO_1238 (O_1238,N_13749,N_12037);
nand UO_1239 (O_1239,N_12234,N_12448);
nor UO_1240 (O_1240,N_13345,N_14843);
or UO_1241 (O_1241,N_14564,N_14764);
nand UO_1242 (O_1242,N_13021,N_13529);
xor UO_1243 (O_1243,N_14615,N_12623);
nor UO_1244 (O_1244,N_13023,N_13682);
nand UO_1245 (O_1245,N_13459,N_13058);
and UO_1246 (O_1246,N_14983,N_12349);
nor UO_1247 (O_1247,N_12556,N_14117);
xnor UO_1248 (O_1248,N_13922,N_14693);
and UO_1249 (O_1249,N_14003,N_12593);
or UO_1250 (O_1250,N_14530,N_14599);
nor UO_1251 (O_1251,N_13310,N_13182);
xor UO_1252 (O_1252,N_14237,N_13326);
and UO_1253 (O_1253,N_12364,N_14030);
nor UO_1254 (O_1254,N_14045,N_13569);
nor UO_1255 (O_1255,N_13259,N_14297);
xnor UO_1256 (O_1256,N_12728,N_14228);
nand UO_1257 (O_1257,N_12183,N_12726);
xnor UO_1258 (O_1258,N_12519,N_13894);
nand UO_1259 (O_1259,N_14091,N_13388);
nand UO_1260 (O_1260,N_14949,N_13952);
nor UO_1261 (O_1261,N_14492,N_13321);
nand UO_1262 (O_1262,N_12398,N_12469);
xor UO_1263 (O_1263,N_14513,N_13658);
xor UO_1264 (O_1264,N_14706,N_12002);
nand UO_1265 (O_1265,N_14201,N_12317);
or UO_1266 (O_1266,N_14654,N_13192);
nor UO_1267 (O_1267,N_14794,N_12378);
and UO_1268 (O_1268,N_13790,N_13775);
and UO_1269 (O_1269,N_12826,N_12196);
nand UO_1270 (O_1270,N_12044,N_13181);
or UO_1271 (O_1271,N_13012,N_13746);
and UO_1272 (O_1272,N_14879,N_13442);
nand UO_1273 (O_1273,N_14698,N_13987);
or UO_1274 (O_1274,N_13980,N_12658);
and UO_1275 (O_1275,N_13122,N_13937);
nand UO_1276 (O_1276,N_12691,N_14392);
and UO_1277 (O_1277,N_12386,N_13692);
and UO_1278 (O_1278,N_13996,N_12836);
or UO_1279 (O_1279,N_13041,N_12248);
nor UO_1280 (O_1280,N_12505,N_12134);
xor UO_1281 (O_1281,N_13991,N_13403);
nor UO_1282 (O_1282,N_13896,N_14133);
and UO_1283 (O_1283,N_12389,N_12894);
nor UO_1284 (O_1284,N_14549,N_12155);
or UO_1285 (O_1285,N_13489,N_13452);
or UO_1286 (O_1286,N_14646,N_14638);
and UO_1287 (O_1287,N_12698,N_12750);
nor UO_1288 (O_1288,N_14116,N_14999);
and UO_1289 (O_1289,N_14124,N_13054);
and UO_1290 (O_1290,N_12162,N_12280);
nand UO_1291 (O_1291,N_12745,N_13832);
or UO_1292 (O_1292,N_12526,N_13668);
nand UO_1293 (O_1293,N_14076,N_14746);
xnor UO_1294 (O_1294,N_12986,N_14415);
nor UO_1295 (O_1295,N_13229,N_13078);
nand UO_1296 (O_1296,N_14942,N_13798);
or UO_1297 (O_1297,N_13929,N_12827);
nor UO_1298 (O_1298,N_12401,N_12810);
or UO_1299 (O_1299,N_13202,N_13817);
or UO_1300 (O_1300,N_14489,N_13024);
nor UO_1301 (O_1301,N_12817,N_13966);
xnor UO_1302 (O_1302,N_14007,N_14156);
nor UO_1303 (O_1303,N_13014,N_13377);
or UO_1304 (O_1304,N_13220,N_13720);
and UO_1305 (O_1305,N_14678,N_12801);
and UO_1306 (O_1306,N_13535,N_12724);
nand UO_1307 (O_1307,N_12639,N_12498);
nand UO_1308 (O_1308,N_14010,N_13983);
nor UO_1309 (O_1309,N_14042,N_14816);
or UO_1310 (O_1310,N_12884,N_12048);
xor UO_1311 (O_1311,N_12298,N_13505);
or UO_1312 (O_1312,N_14077,N_14960);
nand UO_1313 (O_1313,N_12950,N_12719);
nor UO_1314 (O_1314,N_14679,N_12388);
and UO_1315 (O_1315,N_12490,N_13100);
and UO_1316 (O_1316,N_12710,N_12406);
xor UO_1317 (O_1317,N_13589,N_12073);
nand UO_1318 (O_1318,N_12644,N_13008);
nor UO_1319 (O_1319,N_14707,N_12550);
nand UO_1320 (O_1320,N_14750,N_14935);
or UO_1321 (O_1321,N_13236,N_14738);
nor UO_1322 (O_1322,N_14860,N_14393);
nand UO_1323 (O_1323,N_13177,N_13663);
nor UO_1324 (O_1324,N_13541,N_14203);
and UO_1325 (O_1325,N_12971,N_14265);
or UO_1326 (O_1326,N_14559,N_12717);
or UO_1327 (O_1327,N_14170,N_13133);
and UO_1328 (O_1328,N_12281,N_13019);
nand UO_1329 (O_1329,N_12690,N_12221);
nand UO_1330 (O_1330,N_13995,N_13822);
nand UO_1331 (O_1331,N_14107,N_14240);
and UO_1332 (O_1332,N_13169,N_14557);
nor UO_1333 (O_1333,N_13094,N_14482);
and UO_1334 (O_1334,N_12201,N_14959);
or UO_1335 (O_1335,N_13712,N_13261);
or UO_1336 (O_1336,N_12457,N_13235);
and UO_1337 (O_1337,N_14931,N_13698);
xor UO_1338 (O_1338,N_13150,N_14336);
xnor UO_1339 (O_1339,N_14736,N_13719);
or UO_1340 (O_1340,N_14886,N_14234);
nand UO_1341 (O_1341,N_12683,N_14733);
or UO_1342 (O_1342,N_12400,N_12520);
nor UO_1343 (O_1343,N_13559,N_14662);
nand UO_1344 (O_1344,N_12594,N_14862);
nand UO_1345 (O_1345,N_14901,N_12830);
or UO_1346 (O_1346,N_12966,N_14922);
nor UO_1347 (O_1347,N_12770,N_13462);
nor UO_1348 (O_1348,N_12583,N_13472);
nor UO_1349 (O_1349,N_13884,N_14708);
nor UO_1350 (O_1350,N_14371,N_14291);
nor UO_1351 (O_1351,N_14296,N_14374);
and UO_1352 (O_1352,N_14944,N_13287);
and UO_1353 (O_1353,N_13304,N_13946);
or UO_1354 (O_1354,N_13696,N_12405);
nor UO_1355 (O_1355,N_12185,N_14560);
nand UO_1356 (O_1356,N_14150,N_12230);
nand UO_1357 (O_1357,N_12403,N_12174);
nand UO_1358 (O_1358,N_14741,N_13067);
and UO_1359 (O_1359,N_12762,N_14428);
and UO_1360 (O_1360,N_13383,N_12402);
and UO_1361 (O_1361,N_14735,N_14510);
nor UO_1362 (O_1362,N_14015,N_14321);
nand UO_1363 (O_1363,N_13423,N_14356);
nor UO_1364 (O_1364,N_12245,N_14168);
and UO_1365 (O_1365,N_13659,N_13171);
or UO_1366 (O_1366,N_12157,N_14421);
and UO_1367 (O_1367,N_14753,N_13789);
or UO_1368 (O_1368,N_13920,N_13963);
or UO_1369 (O_1369,N_14903,N_14304);
and UO_1370 (O_1370,N_13378,N_14387);
or UO_1371 (O_1371,N_14183,N_13303);
and UO_1372 (O_1372,N_14585,N_14747);
nor UO_1373 (O_1373,N_13145,N_13935);
nor UO_1374 (O_1374,N_12366,N_12271);
nand UO_1375 (O_1375,N_13737,N_13942);
or UO_1376 (O_1376,N_13854,N_14144);
and UO_1377 (O_1377,N_14136,N_12419);
and UO_1378 (O_1378,N_14037,N_14602);
nor UO_1379 (O_1379,N_14323,N_13270);
nor UO_1380 (O_1380,N_12807,N_14227);
nand UO_1381 (O_1381,N_14185,N_13871);
or UO_1382 (O_1382,N_12678,N_14783);
or UO_1383 (O_1383,N_12946,N_14411);
nand UO_1384 (O_1384,N_14368,N_13813);
nand UO_1385 (O_1385,N_12340,N_12941);
nand UO_1386 (O_1386,N_12343,N_13957);
nand UO_1387 (O_1387,N_14910,N_12981);
nand UO_1388 (O_1388,N_14065,N_13000);
xor UO_1389 (O_1389,N_14765,N_13714);
or UO_1390 (O_1390,N_13515,N_13040);
nor UO_1391 (O_1391,N_14519,N_14854);
nand UO_1392 (O_1392,N_12036,N_14189);
nor UO_1393 (O_1393,N_12808,N_13104);
nor UO_1394 (O_1394,N_13990,N_14328);
xnor UO_1395 (O_1395,N_14014,N_12671);
xnor UO_1396 (O_1396,N_14614,N_12468);
xnor UO_1397 (O_1397,N_12382,N_12051);
nand UO_1398 (O_1398,N_12017,N_13683);
and UO_1399 (O_1399,N_13114,N_14964);
xor UO_1400 (O_1400,N_13926,N_12794);
or UO_1401 (O_1401,N_14073,N_13254);
and UO_1402 (O_1402,N_14243,N_14047);
or UO_1403 (O_1403,N_12861,N_13440);
or UO_1404 (O_1404,N_13757,N_12528);
xor UO_1405 (O_1405,N_14157,N_14036);
nand UO_1406 (O_1406,N_12608,N_12852);
xnor UO_1407 (O_1407,N_12081,N_12692);
nand UO_1408 (O_1408,N_14405,N_13468);
nand UO_1409 (O_1409,N_12533,N_13760);
nor UO_1410 (O_1410,N_14216,N_14311);
xnor UO_1411 (O_1411,N_14179,N_14241);
nor UO_1412 (O_1412,N_12368,N_14916);
and UO_1413 (O_1413,N_14588,N_12838);
xnor UO_1414 (O_1414,N_13072,N_13953);
nor UO_1415 (O_1415,N_14143,N_12204);
or UO_1416 (O_1416,N_14383,N_14070);
and UO_1417 (O_1417,N_12740,N_13028);
or UO_1418 (O_1418,N_14844,N_12016);
nor UO_1419 (O_1419,N_12369,N_12408);
nor UO_1420 (O_1420,N_12396,N_14993);
or UO_1421 (O_1421,N_12039,N_12010);
nor UO_1422 (O_1422,N_12411,N_13738);
nand UO_1423 (O_1423,N_12751,N_14418);
or UO_1424 (O_1424,N_14474,N_12935);
nor UO_1425 (O_1425,N_13011,N_13921);
nor UO_1426 (O_1426,N_13161,N_13762);
xnor UO_1427 (O_1427,N_12938,N_13222);
nor UO_1428 (O_1428,N_12239,N_14450);
xnor UO_1429 (O_1429,N_14963,N_14283);
nand UO_1430 (O_1430,N_12326,N_14354);
or UO_1431 (O_1431,N_12863,N_12182);
xor UO_1432 (O_1432,N_12796,N_13507);
and UO_1433 (O_1433,N_13566,N_12563);
or UO_1434 (O_1434,N_14600,N_12430);
and UO_1435 (O_1435,N_14651,N_12546);
and UO_1436 (O_1436,N_12758,N_12500);
nand UO_1437 (O_1437,N_12362,N_14001);
nor UO_1438 (O_1438,N_13092,N_13913);
nor UO_1439 (O_1439,N_13598,N_13940);
or UO_1440 (O_1440,N_12901,N_12373);
or UO_1441 (O_1441,N_13816,N_13955);
or UO_1442 (O_1442,N_14928,N_13700);
nor UO_1443 (O_1443,N_14778,N_14339);
and UO_1444 (O_1444,N_13879,N_13839);
xor UO_1445 (O_1445,N_14347,N_13763);
and UO_1446 (O_1446,N_14874,N_13883);
nand UO_1447 (O_1447,N_14385,N_12197);
nand UO_1448 (O_1448,N_14361,N_14622);
and UO_1449 (O_1449,N_14655,N_13868);
and UO_1450 (O_1450,N_13073,N_12198);
nand UO_1451 (O_1451,N_12314,N_14453);
nor UO_1452 (O_1452,N_12793,N_14440);
xor UO_1453 (O_1453,N_12258,N_14660);
xor UO_1454 (O_1454,N_13944,N_13699);
nand UO_1455 (O_1455,N_13815,N_13109);
nor UO_1456 (O_1456,N_13392,N_13077);
and UO_1457 (O_1457,N_12785,N_12091);
and UO_1458 (O_1458,N_12171,N_14882);
nand UO_1459 (O_1459,N_14994,N_13908);
nor UO_1460 (O_1460,N_14312,N_14591);
or UO_1461 (O_1461,N_13621,N_14388);
or UO_1462 (O_1462,N_13271,N_14947);
and UO_1463 (O_1463,N_12954,N_13250);
nor UO_1464 (O_1464,N_14466,N_12335);
xor UO_1465 (O_1465,N_12752,N_12727);
or UO_1466 (O_1466,N_14663,N_14982);
or UO_1467 (O_1467,N_13715,N_13227);
and UO_1468 (O_1468,N_13441,N_14399);
xor UO_1469 (O_1469,N_13899,N_13144);
xnor UO_1470 (O_1470,N_14320,N_12716);
nor UO_1471 (O_1471,N_12506,N_13086);
nor UO_1472 (O_1472,N_14058,N_14763);
nor UO_1473 (O_1473,N_12525,N_13337);
or UO_1474 (O_1474,N_14027,N_13409);
nand UO_1475 (O_1475,N_14956,N_12123);
nand UO_1476 (O_1476,N_14350,N_14326);
xor UO_1477 (O_1477,N_13445,N_13130);
or UO_1478 (O_1478,N_14613,N_14508);
and UO_1479 (O_1479,N_12575,N_12360);
nor UO_1480 (O_1480,N_12973,N_13152);
or UO_1481 (O_1481,N_13269,N_13588);
and UO_1482 (O_1482,N_12414,N_12721);
or UO_1483 (O_1483,N_12790,N_14542);
and UO_1484 (O_1484,N_12900,N_13199);
nor UO_1485 (O_1485,N_13142,N_13650);
nand UO_1486 (O_1486,N_14395,N_13046);
nand UO_1487 (O_1487,N_12178,N_12452);
nor UO_1488 (O_1488,N_12775,N_13156);
and UO_1489 (O_1489,N_13551,N_14621);
and UO_1490 (O_1490,N_12549,N_13537);
nor UO_1491 (O_1491,N_13115,N_13376);
nand UO_1492 (O_1492,N_14925,N_14524);
or UO_1493 (O_1493,N_13830,N_13530);
and UO_1494 (O_1494,N_12041,N_13628);
or UO_1495 (O_1495,N_12497,N_12604);
and UO_1496 (O_1496,N_14793,N_13216);
xor UO_1497 (O_1497,N_13180,N_13904);
and UO_1498 (O_1498,N_12723,N_13992);
and UO_1499 (O_1499,N_14932,N_13210);
and UO_1500 (O_1500,N_12968,N_12283);
nand UO_1501 (O_1501,N_13912,N_12833);
or UO_1502 (O_1502,N_12727,N_13299);
and UO_1503 (O_1503,N_14967,N_13757);
nor UO_1504 (O_1504,N_13950,N_12033);
xnor UO_1505 (O_1505,N_14970,N_13127);
and UO_1506 (O_1506,N_13894,N_13377);
and UO_1507 (O_1507,N_14790,N_13899);
nand UO_1508 (O_1508,N_12163,N_13728);
and UO_1509 (O_1509,N_13890,N_12763);
nand UO_1510 (O_1510,N_14858,N_12037);
nor UO_1511 (O_1511,N_13532,N_14715);
and UO_1512 (O_1512,N_13788,N_14931);
or UO_1513 (O_1513,N_12318,N_12770);
nand UO_1514 (O_1514,N_14024,N_13946);
nand UO_1515 (O_1515,N_13786,N_13271);
and UO_1516 (O_1516,N_14287,N_14256);
nand UO_1517 (O_1517,N_14859,N_13936);
or UO_1518 (O_1518,N_14725,N_12566);
xnor UO_1519 (O_1519,N_12910,N_13933);
xnor UO_1520 (O_1520,N_13089,N_14652);
nand UO_1521 (O_1521,N_12528,N_14513);
nand UO_1522 (O_1522,N_12660,N_13513);
xor UO_1523 (O_1523,N_12823,N_14131);
nor UO_1524 (O_1524,N_12745,N_14239);
xnor UO_1525 (O_1525,N_14797,N_12420);
or UO_1526 (O_1526,N_12425,N_12173);
and UO_1527 (O_1527,N_14939,N_13328);
and UO_1528 (O_1528,N_14809,N_14049);
nor UO_1529 (O_1529,N_12460,N_13866);
xor UO_1530 (O_1530,N_12557,N_13002);
nand UO_1531 (O_1531,N_14386,N_14512);
or UO_1532 (O_1532,N_13874,N_14080);
nor UO_1533 (O_1533,N_14825,N_14260);
nor UO_1534 (O_1534,N_14238,N_14618);
or UO_1535 (O_1535,N_13839,N_13561);
nor UO_1536 (O_1536,N_14859,N_14923);
and UO_1537 (O_1537,N_14866,N_13086);
nand UO_1538 (O_1538,N_12462,N_13487);
nand UO_1539 (O_1539,N_14159,N_13966);
nor UO_1540 (O_1540,N_13817,N_12804);
and UO_1541 (O_1541,N_14370,N_13376);
or UO_1542 (O_1542,N_13796,N_13536);
nor UO_1543 (O_1543,N_12353,N_13885);
xnor UO_1544 (O_1544,N_13932,N_14657);
xnor UO_1545 (O_1545,N_13218,N_14592);
or UO_1546 (O_1546,N_14342,N_12849);
nand UO_1547 (O_1547,N_14310,N_12518);
nand UO_1548 (O_1548,N_12481,N_14805);
nand UO_1549 (O_1549,N_14959,N_12178);
or UO_1550 (O_1550,N_14358,N_12646);
nor UO_1551 (O_1551,N_14317,N_12204);
or UO_1552 (O_1552,N_14959,N_12284);
or UO_1553 (O_1553,N_12461,N_12322);
nand UO_1554 (O_1554,N_14620,N_12502);
nor UO_1555 (O_1555,N_14628,N_13980);
nand UO_1556 (O_1556,N_14798,N_14710);
nand UO_1557 (O_1557,N_14283,N_14850);
nor UO_1558 (O_1558,N_13655,N_14020);
and UO_1559 (O_1559,N_14808,N_12300);
xor UO_1560 (O_1560,N_14250,N_13115);
and UO_1561 (O_1561,N_14826,N_14199);
xor UO_1562 (O_1562,N_14699,N_12053);
xor UO_1563 (O_1563,N_14668,N_12357);
nor UO_1564 (O_1564,N_12156,N_13549);
or UO_1565 (O_1565,N_12685,N_13120);
nor UO_1566 (O_1566,N_14740,N_13894);
nor UO_1567 (O_1567,N_14003,N_14531);
xor UO_1568 (O_1568,N_13103,N_12594);
or UO_1569 (O_1569,N_12338,N_13182);
and UO_1570 (O_1570,N_13953,N_13981);
xor UO_1571 (O_1571,N_14836,N_12541);
nand UO_1572 (O_1572,N_14974,N_12235);
nand UO_1573 (O_1573,N_12842,N_12836);
or UO_1574 (O_1574,N_13863,N_12598);
nand UO_1575 (O_1575,N_12393,N_13471);
xnor UO_1576 (O_1576,N_13533,N_14809);
nand UO_1577 (O_1577,N_12241,N_13812);
or UO_1578 (O_1578,N_14401,N_14137);
and UO_1579 (O_1579,N_12078,N_14309);
or UO_1580 (O_1580,N_12064,N_14595);
nor UO_1581 (O_1581,N_14290,N_14210);
nand UO_1582 (O_1582,N_13236,N_13005);
or UO_1583 (O_1583,N_13602,N_12002);
or UO_1584 (O_1584,N_13396,N_13042);
nor UO_1585 (O_1585,N_13408,N_13236);
nor UO_1586 (O_1586,N_14828,N_13740);
and UO_1587 (O_1587,N_12405,N_14272);
nand UO_1588 (O_1588,N_14464,N_12534);
xnor UO_1589 (O_1589,N_12428,N_12522);
nor UO_1590 (O_1590,N_14265,N_14027);
or UO_1591 (O_1591,N_14234,N_14020);
nor UO_1592 (O_1592,N_14576,N_13151);
nand UO_1593 (O_1593,N_13286,N_14041);
nand UO_1594 (O_1594,N_12457,N_14721);
or UO_1595 (O_1595,N_13889,N_13278);
and UO_1596 (O_1596,N_12314,N_13591);
nor UO_1597 (O_1597,N_12864,N_13857);
nand UO_1598 (O_1598,N_14792,N_13520);
nand UO_1599 (O_1599,N_12803,N_14738);
nand UO_1600 (O_1600,N_13994,N_14144);
nand UO_1601 (O_1601,N_13829,N_12530);
or UO_1602 (O_1602,N_12268,N_13113);
and UO_1603 (O_1603,N_14034,N_13290);
or UO_1604 (O_1604,N_12863,N_12106);
nor UO_1605 (O_1605,N_12667,N_12891);
nor UO_1606 (O_1606,N_12534,N_13407);
or UO_1607 (O_1607,N_12819,N_13706);
nand UO_1608 (O_1608,N_12278,N_14449);
and UO_1609 (O_1609,N_14897,N_12647);
xor UO_1610 (O_1610,N_13671,N_12471);
nand UO_1611 (O_1611,N_13113,N_13119);
and UO_1612 (O_1612,N_13458,N_14140);
and UO_1613 (O_1613,N_13516,N_12366);
and UO_1614 (O_1614,N_14676,N_13809);
or UO_1615 (O_1615,N_14148,N_12786);
nor UO_1616 (O_1616,N_13748,N_14000);
or UO_1617 (O_1617,N_13047,N_13397);
nand UO_1618 (O_1618,N_12964,N_14826);
nand UO_1619 (O_1619,N_14921,N_12976);
nor UO_1620 (O_1620,N_12396,N_13385);
xnor UO_1621 (O_1621,N_14186,N_12270);
and UO_1622 (O_1622,N_14851,N_14461);
nor UO_1623 (O_1623,N_14109,N_12563);
nor UO_1624 (O_1624,N_13096,N_13355);
nand UO_1625 (O_1625,N_12336,N_12900);
or UO_1626 (O_1626,N_13659,N_14005);
xnor UO_1627 (O_1627,N_13273,N_12568);
nor UO_1628 (O_1628,N_13200,N_13093);
nor UO_1629 (O_1629,N_13147,N_12592);
or UO_1630 (O_1630,N_13707,N_14060);
and UO_1631 (O_1631,N_14032,N_13946);
nor UO_1632 (O_1632,N_14170,N_14493);
nand UO_1633 (O_1633,N_12342,N_13407);
nand UO_1634 (O_1634,N_13526,N_12672);
nand UO_1635 (O_1635,N_12981,N_14096);
nand UO_1636 (O_1636,N_13651,N_14982);
or UO_1637 (O_1637,N_13825,N_13627);
xnor UO_1638 (O_1638,N_12214,N_12818);
xnor UO_1639 (O_1639,N_12265,N_14336);
xor UO_1640 (O_1640,N_13917,N_14449);
nor UO_1641 (O_1641,N_13809,N_13390);
nor UO_1642 (O_1642,N_14474,N_13950);
nor UO_1643 (O_1643,N_14401,N_12124);
nand UO_1644 (O_1644,N_13228,N_14426);
or UO_1645 (O_1645,N_14883,N_14394);
nand UO_1646 (O_1646,N_12858,N_12501);
xor UO_1647 (O_1647,N_12491,N_13464);
nand UO_1648 (O_1648,N_13389,N_14859);
xor UO_1649 (O_1649,N_14236,N_14243);
xnor UO_1650 (O_1650,N_13352,N_13536);
or UO_1651 (O_1651,N_12614,N_12792);
nand UO_1652 (O_1652,N_12120,N_14816);
or UO_1653 (O_1653,N_12264,N_14282);
and UO_1654 (O_1654,N_12235,N_12782);
and UO_1655 (O_1655,N_13363,N_12707);
xor UO_1656 (O_1656,N_12616,N_12515);
or UO_1657 (O_1657,N_14481,N_13821);
xor UO_1658 (O_1658,N_12580,N_13238);
and UO_1659 (O_1659,N_13745,N_13020);
and UO_1660 (O_1660,N_14757,N_13712);
nor UO_1661 (O_1661,N_14352,N_14583);
and UO_1662 (O_1662,N_13678,N_12128);
or UO_1663 (O_1663,N_14131,N_12017);
nor UO_1664 (O_1664,N_12983,N_14326);
nor UO_1665 (O_1665,N_13157,N_13552);
nor UO_1666 (O_1666,N_14057,N_12527);
nand UO_1667 (O_1667,N_14296,N_12459);
and UO_1668 (O_1668,N_14234,N_14752);
and UO_1669 (O_1669,N_14887,N_14589);
or UO_1670 (O_1670,N_14473,N_14963);
nand UO_1671 (O_1671,N_12528,N_12175);
or UO_1672 (O_1672,N_13089,N_14617);
nand UO_1673 (O_1673,N_12946,N_12242);
and UO_1674 (O_1674,N_14897,N_12494);
and UO_1675 (O_1675,N_14327,N_14693);
or UO_1676 (O_1676,N_12167,N_12842);
or UO_1677 (O_1677,N_14870,N_12533);
and UO_1678 (O_1678,N_13453,N_14887);
or UO_1679 (O_1679,N_14256,N_13838);
or UO_1680 (O_1680,N_12198,N_12373);
nor UO_1681 (O_1681,N_12510,N_14084);
nand UO_1682 (O_1682,N_12357,N_13083);
and UO_1683 (O_1683,N_12807,N_13013);
xor UO_1684 (O_1684,N_12185,N_13849);
nand UO_1685 (O_1685,N_13230,N_14508);
and UO_1686 (O_1686,N_14571,N_14677);
or UO_1687 (O_1687,N_14156,N_12900);
or UO_1688 (O_1688,N_12529,N_12501);
nor UO_1689 (O_1689,N_14646,N_12457);
nor UO_1690 (O_1690,N_12001,N_14637);
nand UO_1691 (O_1691,N_12613,N_14572);
nand UO_1692 (O_1692,N_14451,N_13118);
xnor UO_1693 (O_1693,N_14096,N_13186);
or UO_1694 (O_1694,N_13640,N_14035);
xnor UO_1695 (O_1695,N_12184,N_13214);
nand UO_1696 (O_1696,N_12540,N_13924);
and UO_1697 (O_1697,N_13296,N_14003);
nor UO_1698 (O_1698,N_13634,N_13438);
nor UO_1699 (O_1699,N_13918,N_13312);
nor UO_1700 (O_1700,N_14829,N_12041);
xnor UO_1701 (O_1701,N_14566,N_12038);
nand UO_1702 (O_1702,N_12514,N_14785);
and UO_1703 (O_1703,N_12245,N_13985);
or UO_1704 (O_1704,N_12390,N_14056);
or UO_1705 (O_1705,N_12538,N_12922);
nor UO_1706 (O_1706,N_13140,N_14311);
and UO_1707 (O_1707,N_14119,N_13271);
xor UO_1708 (O_1708,N_14164,N_13459);
and UO_1709 (O_1709,N_12638,N_12034);
or UO_1710 (O_1710,N_13625,N_12097);
or UO_1711 (O_1711,N_12230,N_13325);
nand UO_1712 (O_1712,N_14120,N_13626);
nand UO_1713 (O_1713,N_13248,N_13544);
and UO_1714 (O_1714,N_13445,N_13515);
nor UO_1715 (O_1715,N_14199,N_12750);
or UO_1716 (O_1716,N_14034,N_13552);
nand UO_1717 (O_1717,N_12333,N_13241);
nor UO_1718 (O_1718,N_14951,N_13587);
xor UO_1719 (O_1719,N_13113,N_14970);
and UO_1720 (O_1720,N_13346,N_13768);
nor UO_1721 (O_1721,N_13609,N_13668);
xnor UO_1722 (O_1722,N_14381,N_14148);
nor UO_1723 (O_1723,N_12179,N_13340);
or UO_1724 (O_1724,N_12053,N_12267);
or UO_1725 (O_1725,N_14414,N_12109);
and UO_1726 (O_1726,N_12379,N_12724);
or UO_1727 (O_1727,N_13377,N_14145);
or UO_1728 (O_1728,N_14176,N_14813);
xnor UO_1729 (O_1729,N_14232,N_12599);
nand UO_1730 (O_1730,N_12015,N_12150);
or UO_1731 (O_1731,N_13391,N_14998);
nand UO_1732 (O_1732,N_13128,N_12862);
or UO_1733 (O_1733,N_13514,N_14133);
or UO_1734 (O_1734,N_12308,N_13841);
xor UO_1735 (O_1735,N_12810,N_13164);
and UO_1736 (O_1736,N_12584,N_12219);
or UO_1737 (O_1737,N_13794,N_13697);
nand UO_1738 (O_1738,N_12449,N_13543);
or UO_1739 (O_1739,N_13060,N_12598);
xnor UO_1740 (O_1740,N_12266,N_14739);
and UO_1741 (O_1741,N_12838,N_14485);
and UO_1742 (O_1742,N_14993,N_14132);
nand UO_1743 (O_1743,N_13579,N_13493);
xor UO_1744 (O_1744,N_14114,N_13414);
nand UO_1745 (O_1745,N_13160,N_14754);
or UO_1746 (O_1746,N_14665,N_13396);
and UO_1747 (O_1747,N_13042,N_14165);
xnor UO_1748 (O_1748,N_12123,N_14126);
nor UO_1749 (O_1749,N_14407,N_14223);
or UO_1750 (O_1750,N_14979,N_14706);
nor UO_1751 (O_1751,N_12335,N_12450);
or UO_1752 (O_1752,N_13863,N_12590);
xor UO_1753 (O_1753,N_14451,N_12496);
nand UO_1754 (O_1754,N_12056,N_13474);
nand UO_1755 (O_1755,N_14700,N_13972);
nand UO_1756 (O_1756,N_12328,N_12260);
or UO_1757 (O_1757,N_13556,N_13559);
or UO_1758 (O_1758,N_13850,N_12332);
and UO_1759 (O_1759,N_12682,N_12797);
xor UO_1760 (O_1760,N_14485,N_12387);
nor UO_1761 (O_1761,N_13531,N_13755);
or UO_1762 (O_1762,N_13159,N_12581);
or UO_1763 (O_1763,N_12990,N_14078);
nand UO_1764 (O_1764,N_12831,N_14287);
nor UO_1765 (O_1765,N_12041,N_13924);
or UO_1766 (O_1766,N_13915,N_14172);
nand UO_1767 (O_1767,N_13172,N_14101);
nand UO_1768 (O_1768,N_13946,N_14205);
nand UO_1769 (O_1769,N_13063,N_14708);
nand UO_1770 (O_1770,N_12000,N_13127);
nor UO_1771 (O_1771,N_13821,N_13003);
or UO_1772 (O_1772,N_14961,N_14185);
nand UO_1773 (O_1773,N_13453,N_12080);
and UO_1774 (O_1774,N_12471,N_12126);
xnor UO_1775 (O_1775,N_14604,N_14291);
nand UO_1776 (O_1776,N_12101,N_12457);
nand UO_1777 (O_1777,N_13803,N_12800);
and UO_1778 (O_1778,N_12094,N_14284);
and UO_1779 (O_1779,N_13239,N_14085);
nor UO_1780 (O_1780,N_12633,N_13613);
and UO_1781 (O_1781,N_14326,N_14384);
nor UO_1782 (O_1782,N_13377,N_13654);
nor UO_1783 (O_1783,N_12993,N_14351);
nor UO_1784 (O_1784,N_12518,N_13190);
or UO_1785 (O_1785,N_13540,N_12459);
or UO_1786 (O_1786,N_14121,N_12147);
and UO_1787 (O_1787,N_14059,N_12904);
nor UO_1788 (O_1788,N_12207,N_12445);
and UO_1789 (O_1789,N_13841,N_12402);
and UO_1790 (O_1790,N_13571,N_13985);
and UO_1791 (O_1791,N_14256,N_14414);
nand UO_1792 (O_1792,N_12347,N_12449);
and UO_1793 (O_1793,N_14618,N_12612);
or UO_1794 (O_1794,N_12398,N_14664);
and UO_1795 (O_1795,N_14075,N_13272);
nor UO_1796 (O_1796,N_12986,N_14729);
or UO_1797 (O_1797,N_14309,N_12180);
nand UO_1798 (O_1798,N_12690,N_13671);
or UO_1799 (O_1799,N_12964,N_12276);
nor UO_1800 (O_1800,N_12738,N_12059);
nand UO_1801 (O_1801,N_14339,N_14666);
or UO_1802 (O_1802,N_12663,N_13791);
xnor UO_1803 (O_1803,N_14943,N_13309);
and UO_1804 (O_1804,N_13741,N_12424);
xnor UO_1805 (O_1805,N_14121,N_14025);
and UO_1806 (O_1806,N_13828,N_14777);
nand UO_1807 (O_1807,N_14404,N_14644);
and UO_1808 (O_1808,N_12852,N_13102);
nor UO_1809 (O_1809,N_13752,N_13259);
nand UO_1810 (O_1810,N_13973,N_13394);
or UO_1811 (O_1811,N_13262,N_13633);
and UO_1812 (O_1812,N_14106,N_13171);
nor UO_1813 (O_1813,N_13502,N_14465);
and UO_1814 (O_1814,N_13850,N_13235);
nor UO_1815 (O_1815,N_12227,N_13619);
and UO_1816 (O_1816,N_13515,N_13275);
and UO_1817 (O_1817,N_14117,N_13422);
nand UO_1818 (O_1818,N_14112,N_13654);
or UO_1819 (O_1819,N_13293,N_12883);
and UO_1820 (O_1820,N_12844,N_14258);
xnor UO_1821 (O_1821,N_13037,N_13033);
nor UO_1822 (O_1822,N_12139,N_14091);
or UO_1823 (O_1823,N_13478,N_12174);
and UO_1824 (O_1824,N_13489,N_14136);
or UO_1825 (O_1825,N_13545,N_13378);
and UO_1826 (O_1826,N_12909,N_12901);
or UO_1827 (O_1827,N_14228,N_12062);
nor UO_1828 (O_1828,N_14795,N_13953);
nor UO_1829 (O_1829,N_13197,N_12394);
nand UO_1830 (O_1830,N_12369,N_14536);
nor UO_1831 (O_1831,N_13350,N_13256);
and UO_1832 (O_1832,N_14602,N_13485);
or UO_1833 (O_1833,N_13971,N_13667);
nand UO_1834 (O_1834,N_12553,N_12837);
nand UO_1835 (O_1835,N_14891,N_13496);
xnor UO_1836 (O_1836,N_13951,N_14496);
or UO_1837 (O_1837,N_14982,N_13312);
xor UO_1838 (O_1838,N_13014,N_12123);
or UO_1839 (O_1839,N_12662,N_13752);
and UO_1840 (O_1840,N_14642,N_12692);
nand UO_1841 (O_1841,N_12209,N_14051);
or UO_1842 (O_1842,N_14396,N_13363);
and UO_1843 (O_1843,N_12545,N_12898);
or UO_1844 (O_1844,N_12882,N_13103);
nand UO_1845 (O_1845,N_12811,N_14257);
nor UO_1846 (O_1846,N_12382,N_14804);
and UO_1847 (O_1847,N_12411,N_12399);
nor UO_1848 (O_1848,N_12481,N_14056);
xor UO_1849 (O_1849,N_12403,N_13153);
nand UO_1850 (O_1850,N_12559,N_14454);
xor UO_1851 (O_1851,N_12842,N_14452);
xnor UO_1852 (O_1852,N_14653,N_14697);
nand UO_1853 (O_1853,N_12381,N_12956);
nor UO_1854 (O_1854,N_14254,N_14225);
and UO_1855 (O_1855,N_14816,N_13596);
and UO_1856 (O_1856,N_12607,N_14747);
xnor UO_1857 (O_1857,N_14368,N_13469);
or UO_1858 (O_1858,N_12711,N_14134);
nand UO_1859 (O_1859,N_14983,N_14735);
nor UO_1860 (O_1860,N_14830,N_12564);
nor UO_1861 (O_1861,N_14850,N_13350);
and UO_1862 (O_1862,N_13708,N_12354);
xnor UO_1863 (O_1863,N_12144,N_14371);
nand UO_1864 (O_1864,N_14307,N_14817);
or UO_1865 (O_1865,N_12598,N_13976);
nand UO_1866 (O_1866,N_14118,N_13996);
and UO_1867 (O_1867,N_13125,N_12476);
and UO_1868 (O_1868,N_14818,N_13803);
nor UO_1869 (O_1869,N_13909,N_13583);
nand UO_1870 (O_1870,N_14147,N_14854);
nor UO_1871 (O_1871,N_13344,N_13192);
and UO_1872 (O_1872,N_14422,N_13640);
xor UO_1873 (O_1873,N_14741,N_12234);
and UO_1874 (O_1874,N_12309,N_14826);
or UO_1875 (O_1875,N_12887,N_12378);
nor UO_1876 (O_1876,N_13240,N_12997);
nor UO_1877 (O_1877,N_14800,N_14350);
nor UO_1878 (O_1878,N_12191,N_12773);
or UO_1879 (O_1879,N_14263,N_13234);
and UO_1880 (O_1880,N_12637,N_12275);
xor UO_1881 (O_1881,N_12751,N_13052);
or UO_1882 (O_1882,N_14320,N_13944);
or UO_1883 (O_1883,N_14461,N_14909);
or UO_1884 (O_1884,N_13089,N_14146);
nor UO_1885 (O_1885,N_14957,N_12084);
nor UO_1886 (O_1886,N_12912,N_14217);
and UO_1887 (O_1887,N_14576,N_12018);
nor UO_1888 (O_1888,N_12686,N_12775);
and UO_1889 (O_1889,N_14962,N_13399);
nor UO_1890 (O_1890,N_13636,N_12465);
nand UO_1891 (O_1891,N_12269,N_13104);
and UO_1892 (O_1892,N_14373,N_12358);
nor UO_1893 (O_1893,N_12115,N_13426);
nand UO_1894 (O_1894,N_12164,N_12892);
or UO_1895 (O_1895,N_14872,N_14003);
nand UO_1896 (O_1896,N_12347,N_12128);
or UO_1897 (O_1897,N_14485,N_12793);
nand UO_1898 (O_1898,N_13869,N_12616);
or UO_1899 (O_1899,N_12427,N_12882);
or UO_1900 (O_1900,N_14190,N_13112);
and UO_1901 (O_1901,N_12983,N_14035);
nand UO_1902 (O_1902,N_12232,N_12506);
or UO_1903 (O_1903,N_14174,N_13075);
xor UO_1904 (O_1904,N_12906,N_13406);
and UO_1905 (O_1905,N_13960,N_12895);
nor UO_1906 (O_1906,N_12397,N_12751);
nor UO_1907 (O_1907,N_12353,N_14343);
and UO_1908 (O_1908,N_14345,N_12744);
nor UO_1909 (O_1909,N_13950,N_14549);
xnor UO_1910 (O_1910,N_13852,N_13577);
xor UO_1911 (O_1911,N_13121,N_13158);
nor UO_1912 (O_1912,N_12228,N_13698);
or UO_1913 (O_1913,N_13170,N_14989);
or UO_1914 (O_1914,N_14458,N_14493);
xnor UO_1915 (O_1915,N_14446,N_12677);
and UO_1916 (O_1916,N_14621,N_14401);
nor UO_1917 (O_1917,N_12973,N_13082);
and UO_1918 (O_1918,N_12176,N_14814);
or UO_1919 (O_1919,N_13621,N_12433);
nor UO_1920 (O_1920,N_14358,N_12413);
nand UO_1921 (O_1921,N_12458,N_12812);
nand UO_1922 (O_1922,N_12142,N_14128);
nand UO_1923 (O_1923,N_13408,N_13982);
or UO_1924 (O_1924,N_13288,N_14172);
nor UO_1925 (O_1925,N_12401,N_14144);
and UO_1926 (O_1926,N_13801,N_14989);
and UO_1927 (O_1927,N_13118,N_14417);
nor UO_1928 (O_1928,N_14272,N_12848);
nand UO_1929 (O_1929,N_12860,N_12158);
nand UO_1930 (O_1930,N_13124,N_12608);
and UO_1931 (O_1931,N_14598,N_12625);
nor UO_1932 (O_1932,N_13318,N_14944);
nand UO_1933 (O_1933,N_13411,N_13503);
or UO_1934 (O_1934,N_14272,N_13731);
or UO_1935 (O_1935,N_13409,N_13985);
and UO_1936 (O_1936,N_13598,N_12564);
or UO_1937 (O_1937,N_13891,N_13531);
or UO_1938 (O_1938,N_14256,N_12432);
and UO_1939 (O_1939,N_14569,N_13811);
nand UO_1940 (O_1940,N_12753,N_13400);
or UO_1941 (O_1941,N_12369,N_13510);
xnor UO_1942 (O_1942,N_12647,N_14814);
nand UO_1943 (O_1943,N_13934,N_12789);
and UO_1944 (O_1944,N_13575,N_13693);
or UO_1945 (O_1945,N_14619,N_12536);
nor UO_1946 (O_1946,N_13626,N_14094);
nand UO_1947 (O_1947,N_14951,N_12739);
or UO_1948 (O_1948,N_12658,N_12661);
nand UO_1949 (O_1949,N_12477,N_14100);
or UO_1950 (O_1950,N_12724,N_14147);
nand UO_1951 (O_1951,N_12036,N_12903);
xor UO_1952 (O_1952,N_14738,N_12453);
nand UO_1953 (O_1953,N_13903,N_12574);
xor UO_1954 (O_1954,N_12296,N_14617);
or UO_1955 (O_1955,N_14082,N_14688);
or UO_1956 (O_1956,N_12768,N_13823);
or UO_1957 (O_1957,N_13759,N_14484);
or UO_1958 (O_1958,N_12126,N_12070);
or UO_1959 (O_1959,N_12299,N_13354);
xnor UO_1960 (O_1960,N_13701,N_12670);
nor UO_1961 (O_1961,N_14543,N_12263);
nor UO_1962 (O_1962,N_14943,N_14408);
nand UO_1963 (O_1963,N_14767,N_13938);
nand UO_1964 (O_1964,N_13687,N_12956);
or UO_1965 (O_1965,N_13686,N_13838);
xor UO_1966 (O_1966,N_13103,N_13044);
nor UO_1967 (O_1967,N_12751,N_12715);
nor UO_1968 (O_1968,N_13025,N_13399);
nor UO_1969 (O_1969,N_13720,N_14951);
nand UO_1970 (O_1970,N_12393,N_12137);
nor UO_1971 (O_1971,N_12184,N_13177);
xnor UO_1972 (O_1972,N_12507,N_12431);
or UO_1973 (O_1973,N_14053,N_12259);
or UO_1974 (O_1974,N_13119,N_12191);
nor UO_1975 (O_1975,N_12811,N_13063);
nand UO_1976 (O_1976,N_13377,N_12482);
xor UO_1977 (O_1977,N_13964,N_12823);
or UO_1978 (O_1978,N_14073,N_14929);
or UO_1979 (O_1979,N_12758,N_13816);
or UO_1980 (O_1980,N_12237,N_14071);
nor UO_1981 (O_1981,N_12918,N_14591);
xnor UO_1982 (O_1982,N_13687,N_13010);
nand UO_1983 (O_1983,N_14317,N_12944);
nor UO_1984 (O_1984,N_13363,N_13876);
nor UO_1985 (O_1985,N_14273,N_13305);
or UO_1986 (O_1986,N_13104,N_14430);
and UO_1987 (O_1987,N_13664,N_13918);
and UO_1988 (O_1988,N_14383,N_14483);
nand UO_1989 (O_1989,N_13792,N_13366);
or UO_1990 (O_1990,N_13305,N_14868);
or UO_1991 (O_1991,N_14362,N_12087);
nand UO_1992 (O_1992,N_14183,N_13787);
or UO_1993 (O_1993,N_12498,N_12331);
or UO_1994 (O_1994,N_12768,N_13977);
or UO_1995 (O_1995,N_12708,N_13258);
and UO_1996 (O_1996,N_12387,N_12012);
xnor UO_1997 (O_1997,N_13599,N_12944);
and UO_1998 (O_1998,N_13717,N_14679);
nor UO_1999 (O_1999,N_14498,N_12376);
endmodule