module basic_2000_20000_2500_4_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1721,In_1146);
nor U1 (N_1,In_462,In_1950);
and U2 (N_2,In_269,In_235);
nor U3 (N_3,In_110,In_897);
and U4 (N_4,In_711,In_1022);
nor U5 (N_5,In_150,In_1301);
xnor U6 (N_6,In_1198,In_1317);
xnor U7 (N_7,In_877,In_427);
nand U8 (N_8,In_1722,In_1527);
nand U9 (N_9,In_445,In_1152);
nand U10 (N_10,In_1759,In_1487);
nor U11 (N_11,In_899,In_68);
or U12 (N_12,In_1193,In_1444);
nand U13 (N_13,In_1741,In_1299);
nand U14 (N_14,In_1265,In_739);
or U15 (N_15,In_1206,In_277);
or U16 (N_16,In_1506,In_1900);
nor U17 (N_17,In_1421,In_831);
or U18 (N_18,In_122,In_886);
nor U19 (N_19,In_1336,In_746);
or U20 (N_20,In_271,In_1368);
or U21 (N_21,In_1024,In_102);
nand U22 (N_22,In_284,In_450);
nor U23 (N_23,In_1188,In_1312);
and U24 (N_24,In_1320,In_1877);
and U25 (N_25,In_1075,In_151);
nor U26 (N_26,In_1219,In_1748);
and U27 (N_27,In_755,In_49);
and U28 (N_28,In_708,In_722);
and U29 (N_29,In_1752,In_1513);
nand U30 (N_30,In_806,In_1957);
and U31 (N_31,In_1625,In_1925);
and U32 (N_32,In_1038,In_570);
and U33 (N_33,In_1686,In_1184);
or U34 (N_34,In_536,In_338);
nand U35 (N_35,In_407,In_157);
and U36 (N_36,In_1137,In_1550);
xor U37 (N_37,In_1366,In_1943);
and U38 (N_38,In_1581,In_890);
xor U39 (N_39,In_399,In_1584);
nor U40 (N_40,In_1253,In_1933);
nand U41 (N_41,In_291,In_695);
and U42 (N_42,In_1263,In_1996);
nand U43 (N_43,In_280,In_416);
nand U44 (N_44,In_1113,In_676);
or U45 (N_45,In_825,In_987);
nor U46 (N_46,In_1826,In_753);
and U47 (N_47,In_42,In_1836);
nor U48 (N_48,In_718,In_1539);
and U49 (N_49,In_1754,In_1335);
or U50 (N_50,In_678,In_1955);
xnor U51 (N_51,In_1059,In_17);
or U52 (N_52,In_507,In_1777);
nor U53 (N_53,In_696,In_537);
or U54 (N_54,In_1494,In_1960);
or U55 (N_55,In_489,In_1132);
xor U56 (N_56,In_369,In_1678);
nand U57 (N_57,In_752,In_1736);
nand U58 (N_58,In_193,In_1389);
or U59 (N_59,In_655,In_1094);
nand U60 (N_60,In_1273,In_1369);
nor U61 (N_61,In_1287,In_1018);
nand U62 (N_62,In_1390,In_220);
and U63 (N_63,In_1426,In_805);
or U64 (N_64,In_1873,In_1847);
nand U65 (N_65,In_10,In_440);
and U66 (N_66,In_74,In_207);
xor U67 (N_67,In_479,In_750);
or U68 (N_68,In_146,In_1638);
and U69 (N_69,In_347,In_776);
nor U70 (N_70,In_1191,In_632);
or U71 (N_71,In_448,In_1055);
xnor U72 (N_72,In_749,In_1670);
nor U73 (N_73,In_541,In_1982);
nand U74 (N_74,In_1577,In_251);
nand U75 (N_75,In_1056,In_1082);
nor U76 (N_76,In_578,In_590);
xor U77 (N_77,In_63,In_759);
or U78 (N_78,In_513,In_1802);
xnor U79 (N_79,In_1610,In_30);
nor U80 (N_80,In_14,In_998);
or U81 (N_81,In_691,In_470);
and U82 (N_82,In_893,In_1234);
nor U83 (N_83,In_309,In_661);
nor U84 (N_84,In_41,In_1237);
xnor U85 (N_85,In_60,In_1461);
or U86 (N_86,In_249,In_248);
or U87 (N_87,In_438,In_1293);
and U88 (N_88,In_1092,In_234);
nor U89 (N_89,In_861,In_159);
and U90 (N_90,In_907,In_1425);
nor U91 (N_91,In_3,In_422);
or U92 (N_92,In_414,In_1154);
or U93 (N_93,In_892,In_835);
nand U94 (N_94,In_233,In_1372);
nor U95 (N_95,In_1655,In_257);
nor U96 (N_96,In_1185,In_1109);
and U97 (N_97,In_1037,In_1538);
or U98 (N_98,In_1182,In_1928);
nand U99 (N_99,In_183,In_1159);
and U100 (N_100,In_245,In_1541);
nor U101 (N_101,In_804,In_16);
or U102 (N_102,In_1986,In_1868);
or U103 (N_103,In_32,In_1961);
and U104 (N_104,In_1131,In_1609);
nor U105 (N_105,In_1411,In_794);
nand U106 (N_106,In_1888,In_962);
nand U107 (N_107,In_1825,In_1385);
nand U108 (N_108,In_1173,In_679);
nor U109 (N_109,In_630,In_1787);
nor U110 (N_110,In_1498,In_765);
or U111 (N_111,In_1735,In_1731);
nand U112 (N_112,In_261,In_884);
and U113 (N_113,In_1079,In_993);
and U114 (N_114,In_1375,In_1861);
or U115 (N_115,In_845,In_611);
nand U116 (N_116,In_1290,In_1837);
xor U117 (N_117,In_540,In_1081);
nand U118 (N_118,In_1813,In_686);
or U119 (N_119,In_1102,In_1598);
nor U120 (N_120,In_289,In_1358);
nor U121 (N_121,In_705,In_1653);
nor U122 (N_122,In_848,In_1009);
nor U123 (N_123,In_71,In_1623);
and U124 (N_124,In_36,In_641);
nand U125 (N_125,In_816,In_964);
or U126 (N_126,In_1542,In_626);
xor U127 (N_127,In_1612,In_721);
or U128 (N_128,In_428,In_1050);
or U129 (N_129,In_1879,In_1382);
and U130 (N_130,In_1809,In_734);
nor U131 (N_131,In_1637,In_1895);
and U132 (N_132,In_290,In_1397);
and U133 (N_133,In_996,In_179);
and U134 (N_134,In_894,In_1099);
and U135 (N_135,In_137,In_662);
nand U136 (N_136,In_916,In_480);
and U137 (N_137,In_598,In_891);
nor U138 (N_138,In_1403,In_498);
xor U139 (N_139,In_1854,In_84);
and U140 (N_140,In_500,In_1746);
or U141 (N_141,In_1669,In_70);
nand U142 (N_142,In_593,In_688);
nand U143 (N_143,In_777,In_1098);
and U144 (N_144,In_45,In_1891);
nor U145 (N_145,In_976,In_1027);
or U146 (N_146,In_1449,In_176);
or U147 (N_147,In_46,In_1571);
xnor U148 (N_148,In_94,In_128);
and U149 (N_149,In_954,In_18);
and U150 (N_150,In_454,In_1651);
nor U151 (N_151,In_37,In_173);
and U152 (N_152,In_1819,In_1371);
nor U153 (N_153,In_79,In_1747);
nand U154 (N_154,In_358,In_1294);
and U155 (N_155,In_505,In_1945);
nand U156 (N_156,In_1919,In_1572);
nand U157 (N_157,In_1395,In_949);
nand U158 (N_158,In_1916,In_785);
or U159 (N_159,In_382,In_673);
nor U160 (N_160,In_852,In_1189);
or U161 (N_161,In_1217,In_548);
and U162 (N_162,In_198,In_1215);
and U163 (N_163,In_1829,In_463);
nor U164 (N_164,In_799,In_1093);
nand U165 (N_165,In_573,In_1695);
nand U166 (N_166,In_1857,In_1799);
xnor U167 (N_167,In_324,In_1681);
nand U168 (N_168,In_608,In_228);
and U169 (N_169,In_394,In_1316);
nor U170 (N_170,In_250,In_1624);
nand U171 (N_171,In_1357,In_1241);
or U172 (N_172,In_1295,In_177);
nor U173 (N_173,In_105,In_1463);
nand U174 (N_174,In_1349,In_1871);
nand U175 (N_175,In_951,In_1186);
nor U176 (N_176,In_1264,In_1980);
nor U177 (N_177,In_1008,In_621);
nand U178 (N_178,In_111,In_239);
or U179 (N_179,In_1650,In_11);
xnor U180 (N_180,In_1238,In_1717);
nand U181 (N_181,In_216,In_39);
nand U182 (N_182,In_1780,In_983);
nand U183 (N_183,In_1604,In_531);
or U184 (N_184,In_778,In_491);
nor U185 (N_185,In_1012,In_1483);
or U186 (N_186,In_944,In_1204);
and U187 (N_187,In_1633,In_227);
nand U188 (N_188,In_1148,In_1907);
and U189 (N_189,In_1972,In_1797);
nor U190 (N_190,In_388,In_1201);
nor U191 (N_191,In_1046,In_850);
xor U192 (N_192,In_923,In_1177);
nand U193 (N_193,In_1279,In_123);
and U194 (N_194,In_499,In_380);
nor U195 (N_195,In_485,In_1926);
and U196 (N_196,In_1790,In_1235);
or U197 (N_197,In_254,In_1356);
nand U198 (N_198,In_55,In_1798);
or U199 (N_199,In_1063,In_374);
and U200 (N_200,In_483,In_542);
nand U201 (N_201,In_1326,In_116);
nand U202 (N_202,In_560,In_999);
or U203 (N_203,In_1940,In_855);
xnor U204 (N_204,In_634,In_1884);
xnor U205 (N_205,In_1405,In_172);
or U206 (N_206,In_1812,In_372);
and U207 (N_207,In_1901,In_1416);
nand U208 (N_208,In_62,In_288);
or U209 (N_209,In_1307,In_1782);
xnor U210 (N_210,In_455,In_1123);
and U211 (N_211,In_265,In_675);
nand U212 (N_212,In_909,In_1902);
xnor U213 (N_213,In_109,In_404);
and U214 (N_214,In_534,In_965);
nand U215 (N_215,In_348,In_694);
nor U216 (N_216,In_905,In_1851);
nand U217 (N_217,In_1938,In_1761);
nor U218 (N_218,In_1242,In_947);
or U219 (N_219,In_314,In_167);
nand U220 (N_220,In_1288,In_795);
xnor U221 (N_221,In_1553,In_278);
nand U222 (N_222,In_551,In_1864);
nand U223 (N_223,In_218,In_1057);
and U224 (N_224,In_417,In_466);
nor U225 (N_225,In_262,In_1726);
and U226 (N_226,In_1115,In_15);
or U227 (N_227,In_140,In_136);
xor U228 (N_228,In_1514,In_1480);
and U229 (N_229,In_1255,In_1387);
nor U230 (N_230,In_600,In_1540);
and U231 (N_231,In_1116,In_1406);
or U232 (N_232,In_436,In_1134);
nor U233 (N_233,In_1558,In_614);
nor U234 (N_234,In_1164,In_1985);
or U235 (N_235,In_1345,In_760);
nor U236 (N_236,In_800,In_625);
nand U237 (N_237,In_430,In_325);
and U238 (N_238,In_1816,In_1086);
nand U239 (N_239,In_1200,In_1500);
nand U240 (N_240,In_135,In_1872);
nor U241 (N_241,In_281,In_639);
nor U242 (N_242,In_1744,In_687);
and U243 (N_243,In_212,In_860);
nand U244 (N_244,In_148,In_824);
and U245 (N_245,In_664,In_1646);
and U246 (N_246,In_1642,In_165);
and U247 (N_247,In_1605,In_1552);
and U248 (N_248,In_1060,In_644);
nand U249 (N_249,In_840,In_240);
nand U250 (N_250,In_581,In_230);
nand U251 (N_251,In_846,In_465);
and U252 (N_252,In_1254,In_612);
nand U253 (N_253,In_636,In_1419);
or U254 (N_254,In_1862,In_972);
nor U255 (N_255,In_336,In_563);
or U256 (N_256,In_384,In_1276);
or U257 (N_257,In_1310,In_1935);
nor U258 (N_258,In_67,In_981);
or U259 (N_259,In_833,In_510);
nor U260 (N_260,In_960,In_810);
nor U261 (N_261,In_156,In_152);
or U262 (N_262,In_616,In_955);
nand U263 (N_263,In_1247,In_1652);
nand U264 (N_264,In_35,In_1268);
nand U265 (N_265,In_171,In_1608);
nor U266 (N_266,In_525,In_665);
or U267 (N_267,In_1640,In_270);
and U268 (N_268,In_1260,In_379);
nor U269 (N_269,In_1522,In_1001);
xnor U270 (N_270,In_1465,In_595);
nand U271 (N_271,In_287,In_8);
xnor U272 (N_272,In_1026,In_754);
nor U273 (N_273,In_320,In_1054);
nor U274 (N_274,In_1554,In_1543);
or U275 (N_275,In_124,In_969);
nand U276 (N_276,In_723,In_975);
nor U277 (N_277,In_1233,In_1436);
nand U278 (N_278,In_1750,In_556);
xnor U279 (N_279,In_1679,In_607);
nand U280 (N_280,In_1053,In_1029);
nor U281 (N_281,In_1105,In_1114);
or U282 (N_282,In_874,In_720);
and U283 (N_283,In_126,In_1784);
and U284 (N_284,In_559,In_82);
and U285 (N_285,In_1757,In_1166);
or U286 (N_286,In_995,In_252);
and U287 (N_287,In_1091,In_756);
or U288 (N_288,In_1775,In_1947);
or U289 (N_289,In_1367,In_1163);
and U290 (N_290,In_343,In_1485);
or U291 (N_291,In_1899,In_415);
or U292 (N_292,In_1756,In_1414);
xnor U293 (N_293,In_1319,In_1302);
xnor U294 (N_294,In_895,In_974);
or U295 (N_295,In_400,In_312);
xnor U296 (N_296,In_1030,In_1337);
and U297 (N_297,In_628,In_1126);
nand U298 (N_298,In_20,In_1509);
xnor U299 (N_299,In_1831,In_564);
and U300 (N_300,In_1941,In_1992);
or U301 (N_301,In_202,In_1903);
and U302 (N_302,In_1077,In_937);
or U303 (N_303,In_1573,In_1064);
or U304 (N_304,In_610,In_1250);
nor U305 (N_305,In_575,In_12);
or U306 (N_306,In_475,In_1594);
or U307 (N_307,In_194,In_1631);
and U308 (N_308,In_701,In_175);
or U309 (N_309,In_1392,In_170);
nor U310 (N_310,In_1709,In_1800);
nand U311 (N_311,In_856,In_361);
nand U312 (N_312,In_1607,In_1013);
nand U313 (N_313,In_1621,In_1869);
nor U314 (N_314,In_1489,In_1089);
or U315 (N_315,In_1967,In_129);
nand U316 (N_316,In_624,In_1236);
nand U317 (N_317,In_263,In_579);
and U318 (N_318,In_622,In_1674);
nor U319 (N_319,In_562,In_1684);
nor U320 (N_320,In_1453,In_266);
nand U321 (N_321,In_1025,In_1391);
nor U322 (N_322,In_1785,In_1303);
and U323 (N_323,In_1227,In_1632);
and U324 (N_324,In_1835,In_786);
and U325 (N_325,In_939,In_1781);
or U326 (N_326,In_762,In_323);
xor U327 (N_327,In_149,In_487);
nand U328 (N_328,In_1020,In_1424);
and U329 (N_329,In_571,In_927);
and U330 (N_330,In_189,In_389);
nor U331 (N_331,In_490,In_550);
xnor U332 (N_332,In_1939,In_1010);
or U333 (N_333,In_121,In_792);
nand U334 (N_334,In_1229,In_61);
or U335 (N_335,In_851,In_1853);
xor U336 (N_336,In_1776,In_629);
nor U337 (N_337,In_594,In_980);
nand U338 (N_338,In_1561,In_1508);
xnor U339 (N_339,In_1745,In_1922);
nor U340 (N_340,In_707,In_832);
xnor U341 (N_341,In_1432,In_1065);
and U342 (N_342,In_638,In_908);
or U343 (N_343,In_160,In_1628);
and U344 (N_344,In_1913,In_1378);
nand U345 (N_345,In_353,In_434);
nor U346 (N_346,In_566,In_1773);
and U347 (N_347,In_1138,In_633);
xor U348 (N_348,In_643,In_1833);
or U349 (N_349,In_1015,In_1129);
or U350 (N_350,In_375,In_1074);
nand U351 (N_351,In_657,In_28);
or U352 (N_352,In_1194,In_1306);
nand U353 (N_353,In_1979,In_85);
xor U354 (N_354,In_1546,In_512);
nor U355 (N_355,In_504,In_1145);
or U356 (N_356,In_424,In_1427);
nand U357 (N_357,In_1753,In_431);
nor U358 (N_358,In_132,In_605);
and U359 (N_359,In_118,In_1420);
nor U360 (N_360,In_1417,In_315);
and U361 (N_361,In_1495,In_553);
nand U362 (N_362,In_1751,In_1231);
nand U363 (N_363,In_1051,In_1874);
nand U364 (N_364,In_1520,In_818);
nor U365 (N_365,In_1445,In_1121);
xor U366 (N_366,In_1530,In_6);
or U367 (N_367,In_1153,In_476);
or U368 (N_368,In_1275,In_1647);
nor U369 (N_369,In_1687,In_264);
nor U370 (N_370,In_1591,In_93);
nand U371 (N_371,In_1708,In_1300);
nand U372 (N_372,In_1999,In_58);
or U373 (N_373,In_812,In_519);
xor U374 (N_374,In_714,In_1497);
and U375 (N_375,In_528,In_328);
nor U376 (N_376,In_255,In_1354);
or U377 (N_377,In_1883,In_997);
nor U378 (N_378,In_143,In_1820);
nand U379 (N_379,In_526,In_113);
nor U380 (N_380,In_1711,In_724);
nor U381 (N_381,In_853,In_1556);
and U382 (N_382,In_337,In_758);
xor U383 (N_383,In_1314,In_1507);
and U384 (N_384,In_301,In_572);
or U385 (N_385,In_467,In_1203);
nor U386 (N_386,In_19,In_1796);
or U387 (N_387,In_1965,In_1398);
or U388 (N_388,In_1412,In_1593);
nor U389 (N_389,In_728,In_789);
or U390 (N_390,In_656,In_1150);
and U391 (N_391,In_1724,In_730);
and U392 (N_392,In_1764,In_1692);
and U393 (N_393,In_1220,In_1228);
nor U394 (N_394,In_209,In_1704);
nand U395 (N_395,In_1127,In_161);
and U396 (N_396,In_1702,In_1739);
nor U397 (N_397,In_1071,In_933);
or U398 (N_398,In_557,In_1328);
nor U399 (N_399,In_1524,In_322);
nand U400 (N_400,In_1682,In_232);
and U401 (N_401,In_1376,In_1286);
nor U402 (N_402,In_992,In_341);
nand U403 (N_403,In_1794,In_1824);
nor U404 (N_404,In_936,In_1858);
nor U405 (N_405,In_1330,In_1266);
or U406 (N_406,In_1434,In_1023);
or U407 (N_407,In_1322,In_1443);
nor U408 (N_408,In_390,In_1795);
nor U409 (N_409,In_1517,In_521);
nor U410 (N_410,In_1600,In_1430);
and U411 (N_411,In_213,In_373);
xor U412 (N_412,In_1968,In_1732);
and U413 (N_413,In_1208,In_1755);
or U414 (N_414,In_1963,In_530);
and U415 (N_415,In_418,In_86);
and U416 (N_416,In_1450,In_565);
and U417 (N_417,In_319,In_583);
nand U418 (N_418,In_1881,In_1088);
or U419 (N_419,In_1855,In_1654);
or U420 (N_420,In_1713,In_815);
nand U421 (N_421,In_1918,In_114);
nand U422 (N_422,In_1476,In_1779);
or U423 (N_423,In_967,In_188);
xor U424 (N_424,In_9,In_1688);
nor U425 (N_425,In_1243,In_1849);
nand U426 (N_426,In_774,In_351);
nor U427 (N_427,In_1087,In_1122);
or U428 (N_428,In_841,In_1923);
xnor U429 (N_429,In_843,In_915);
nand U430 (N_430,In_1696,In_1338);
and U431 (N_431,In_1135,In_326);
nor U432 (N_432,In_1418,In_441);
nand U433 (N_433,In_1484,In_669);
nor U434 (N_434,In_1379,In_1165);
nor U435 (N_435,In_862,In_1048);
nand U436 (N_436,In_1665,In_241);
and U437 (N_437,In_1568,In_588);
or U438 (N_438,In_1937,In_313);
or U439 (N_439,In_1212,In_1578);
or U440 (N_440,In_1162,In_1155);
nor U441 (N_441,In_1723,In_5);
nand U442 (N_442,In_1441,In_1887);
or U443 (N_443,In_357,In_1246);
xor U444 (N_444,In_520,In_1249);
nand U445 (N_445,In_1124,In_1564);
nor U446 (N_446,In_1758,In_1422);
xor U447 (N_447,In_1596,In_830);
and U448 (N_448,In_811,In_1587);
nor U449 (N_449,In_561,In_737);
and U450 (N_450,In_757,In_511);
nor U451 (N_451,In_1616,In_1334);
and U452 (N_452,In_1467,In_1141);
or U453 (N_453,In_236,In_1742);
nand U454 (N_454,In_403,In_1214);
and U455 (N_455,In_1906,In_104);
nor U456 (N_456,In_1180,In_1728);
nand U457 (N_457,In_1474,In_1705);
nand U458 (N_458,In_371,In_1977);
nand U459 (N_459,In_921,In_1987);
nor U460 (N_460,In_1332,In_1984);
and U461 (N_461,In_206,In_1559);
nand U462 (N_462,In_69,In_1997);
nor U463 (N_463,In_1142,In_208);
and U464 (N_464,In_1396,In_1639);
and U465 (N_465,In_751,In_959);
or U466 (N_466,In_1280,In_743);
nor U467 (N_467,In_552,In_163);
nand U468 (N_468,In_331,In_168);
or U469 (N_469,In_780,In_934);
nand U470 (N_470,In_574,In_1481);
nor U471 (N_471,In_429,In_1643);
nand U472 (N_472,In_1927,In_1394);
or U473 (N_473,In_1144,In_247);
nand U474 (N_474,In_292,In_1285);
nand U475 (N_475,In_1662,In_606);
and U476 (N_476,In_1663,In_514);
nor U477 (N_477,In_748,In_710);
and U478 (N_478,In_931,In_237);
xor U479 (N_479,In_1716,In_1492);
and U480 (N_480,In_1363,In_596);
nor U481 (N_481,In_1856,In_659);
nand U482 (N_482,In_702,In_200);
or U483 (N_483,In_1457,In_1582);
and U484 (N_484,In_1325,In_637);
and U485 (N_485,In_615,In_139);
nand U486 (N_486,In_1232,In_1488);
or U487 (N_487,In_847,In_620);
or U488 (N_488,In_1034,In_517);
xnor U489 (N_489,In_1599,In_142);
and U490 (N_490,In_1072,In_318);
xor U491 (N_491,In_1904,In_1315);
nor U492 (N_492,In_1039,In_1525);
nand U493 (N_493,In_1763,In_107);
or U494 (N_494,In_735,In_1331);
nand U495 (N_495,In_1021,In_27);
or U496 (N_496,In_619,In_464);
xor U497 (N_497,In_1181,In_77);
nand U498 (N_498,In_138,In_327);
or U499 (N_499,In_1618,In_1240);
or U500 (N_500,In_1017,In_1499);
or U501 (N_501,In_670,In_942);
and U502 (N_502,In_1112,In_221);
nand U503 (N_503,In_370,In_186);
nor U504 (N_504,In_885,In_1442);
and U505 (N_505,In_1437,In_875);
or U506 (N_506,In_225,In_1719);
and U507 (N_507,In_43,In_346);
nand U508 (N_508,In_732,In_97);
or U509 (N_509,In_1090,In_599);
nand U510 (N_510,In_642,In_1042);
nor U511 (N_511,In_1282,In_1932);
and U512 (N_512,In_803,In_854);
or U513 (N_513,In_535,In_1976);
nand U514 (N_514,In_1893,In_547);
and U515 (N_515,In_446,In_305);
and U516 (N_516,In_1769,In_1804);
nor U517 (N_517,In_1626,In_793);
and U518 (N_518,In_1580,In_1211);
xnor U519 (N_519,In_1289,In_769);
nand U520 (N_520,In_1516,In_1834);
or U521 (N_521,In_872,In_1533);
nand U522 (N_522,In_81,In_568);
and U523 (N_523,In_335,In_449);
nand U524 (N_524,In_1168,In_647);
or U525 (N_525,In_1413,In_1333);
and U526 (N_526,In_1676,In_99);
nor U527 (N_527,In_496,In_809);
or U528 (N_528,In_73,In_1158);
nand U529 (N_529,In_1019,In_1668);
nand U530 (N_530,In_989,In_1830);
nor U531 (N_531,In_681,In_672);
nand U532 (N_532,In_90,In_408);
xnor U533 (N_533,In_367,In_344);
and U534 (N_534,In_1710,In_1601);
nand U535 (N_535,In_1401,In_259);
or U536 (N_536,In_376,In_796);
xor U537 (N_537,In_1084,In_219);
nand U538 (N_538,In_13,In_1622);
nand U539 (N_539,In_1700,In_377);
nand U540 (N_540,In_1917,In_1399);
and U541 (N_541,In_1210,In_1706);
nor U542 (N_542,In_692,In_587);
nand U543 (N_543,In_683,In_1482);
or U544 (N_544,In_580,In_1521);
nand U545 (N_545,In_340,In_1197);
nand U546 (N_546,In_395,In_719);
or U547 (N_547,In_47,In_362);
and U548 (N_548,In_1466,In_1171);
nand U549 (N_549,In_1503,In_658);
and U550 (N_550,In_383,In_419);
nand U551 (N_551,In_1880,In_1067);
or U552 (N_552,In_1630,In_1562);
or U553 (N_553,In_1036,In_503);
or U554 (N_554,In_386,In_460);
or U555 (N_555,In_1823,In_920);
and U556 (N_556,In_1791,In_1801);
xnor U557 (N_557,In_1821,In_1360);
and U558 (N_558,In_1551,In_546);
xnor U559 (N_559,In_210,In_260);
or U560 (N_560,In_911,In_204);
nor U561 (N_561,In_1318,In_1951);
nor U562 (N_562,In_350,In_823);
nor U563 (N_563,In_141,In_779);
nor U564 (N_564,In_772,In_807);
nand U565 (N_565,In_761,In_693);
or U566 (N_566,In_1496,In_1740);
nand U567 (N_567,In_1693,In_1657);
nand U568 (N_568,In_985,In_1680);
xnor U569 (N_569,In_516,In_1028);
or U570 (N_570,In_1890,In_297);
nor U571 (N_571,In_447,In_1699);
or U572 (N_572,In_1321,In_898);
nand U573 (N_573,In_192,In_442);
nand U574 (N_574,In_1518,In_387);
nor U575 (N_575,In_162,In_1230);
and U576 (N_576,In_56,In_914);
nand U577 (N_577,In_1061,In_474);
nor U578 (N_578,In_334,In_943);
nor U579 (N_579,In_164,In_524);
and U580 (N_580,In_889,In_787);
or U581 (N_581,In_21,In_984);
nand U582 (N_582,In_274,In_1415);
xnor U583 (N_583,In_838,In_345);
or U584 (N_584,In_1505,In_1946);
nor U585 (N_585,In_1712,In_866);
and U586 (N_586,In_1440,In_34);
and U587 (N_587,In_501,In_273);
and U588 (N_588,In_59,In_709);
and U589 (N_589,In_1267,In_1729);
and U590 (N_590,In_1586,In_1169);
or U591 (N_591,In_704,In_865);
xnor U592 (N_592,In_1218,In_1340);
and U593 (N_593,In_901,In_1878);
nand U594 (N_594,In_900,In_968);
or U595 (N_595,In_130,In_842);
and U596 (N_596,In_929,In_767);
or U597 (N_597,In_1435,In_613);
and U598 (N_598,In_576,In_654);
and U599 (N_599,In_1566,In_1101);
nor U600 (N_600,In_508,In_1078);
nor U601 (N_601,In_869,In_932);
and U602 (N_602,In_922,In_978);
or U603 (N_603,In_770,In_342);
nor U604 (N_604,In_1743,In_1803);
nor U605 (N_605,In_131,In_1187);
xor U606 (N_606,In_829,In_1531);
and U607 (N_607,In_333,In_100);
or U608 (N_608,In_51,In_1000);
or U609 (N_609,In_1774,In_1393);
or U610 (N_610,In_1404,In_396);
nor U611 (N_611,In_1004,In_529);
nand U612 (N_612,In_1661,In_990);
nand U613 (N_613,In_1603,In_203);
nor U614 (N_614,In_982,In_1793);
nor U615 (N_615,In_1355,In_896);
nor U616 (N_616,In_458,In_849);
and U617 (N_617,In_1130,In_586);
and U618 (N_618,In_1298,In_482);
and U619 (N_619,In_1119,In_1136);
nor U620 (N_620,In_1147,In_591);
nor U621 (N_621,In_1590,In_421);
or U622 (N_622,In_256,In_356);
and U623 (N_623,In_1718,In_1140);
and U624 (N_624,In_1560,In_763);
nand U625 (N_625,In_1644,In_1448);
nand U626 (N_626,In_1106,In_23);
nor U627 (N_627,In_392,In_321);
nor U628 (N_628,In_1433,In_1156);
xnor U629 (N_629,In_1974,In_979);
nand U630 (N_630,In_700,In_1068);
nand U631 (N_631,In_1178,In_1822);
nor U632 (N_632,In_668,In_1634);
nand U633 (N_633,In_857,In_1843);
and U634 (N_634,In_1846,In_1157);
nand U635 (N_635,In_1613,In_222);
nand U636 (N_636,In_1576,In_1534);
nand U637 (N_637,In_1083,In_1167);
nor U638 (N_638,In_1730,In_1244);
and U639 (N_639,In_1707,In_788);
xor U640 (N_640,In_185,In_1677);
and U641 (N_641,In_316,In_1765);
nor U642 (N_642,In_745,In_1914);
nand U643 (N_643,In_545,In_492);
or U644 (N_644,In_1971,In_1579);
nor U645 (N_645,In_1685,In_477);
or U646 (N_646,In_1006,In_729);
xor U647 (N_647,In_115,In_1995);
nor U648 (N_648,In_1511,In_1076);
nor U649 (N_649,In_349,In_881);
and U650 (N_650,In_108,In_432);
or U651 (N_651,In_1339,In_1451);
xor U652 (N_652,In_1139,In_1381);
and U653 (N_653,In_1898,In_1959);
or U654 (N_654,In_1555,In_1860);
or U655 (N_655,In_868,In_1786);
or U656 (N_656,In_258,In_1563);
or U657 (N_657,In_1380,In_1973);
or U658 (N_658,In_469,In_1278);
and U659 (N_659,In_826,In_1737);
xnor U660 (N_660,In_1683,In_481);
nand U661 (N_661,In_1792,In_584);
nand U662 (N_662,In_515,In_1248);
and U663 (N_663,In_1305,In_635);
xor U664 (N_664,In_1574,In_468);
nand U665 (N_665,In_790,In_1341);
nor U666 (N_666,In_1170,In_1766);
nand U667 (N_667,In_569,In_935);
nor U668 (N_668,In_1544,In_912);
or U669 (N_669,In_155,In_802);
nor U670 (N_670,In_827,In_178);
or U671 (N_671,In_1954,In_1047);
nand U672 (N_672,In_1714,In_727);
nor U673 (N_673,In_650,In_294);
nor U674 (N_674,In_782,In_1245);
nand U675 (N_675,In_385,In_48);
xor U676 (N_676,In_1103,In_1350);
xnor U677 (N_677,In_406,In_437);
or U678 (N_678,In_381,In_870);
xnor U679 (N_679,In_1892,In_1327);
or U680 (N_680,In_443,In_439);
nand U681 (N_681,In_180,In_1636);
nor U682 (N_682,In_538,In_1125);
nand U683 (N_683,In_1364,In_522);
xor U684 (N_684,In_783,In_275);
and U685 (N_685,In_1671,In_1477);
nor U686 (N_686,In_1512,In_1216);
or U687 (N_687,In_201,In_1840);
nand U688 (N_688,In_1003,In_1172);
or U689 (N_689,In_1468,In_651);
nand U690 (N_690,In_518,In_1535);
or U691 (N_691,In_558,In_801);
nor U692 (N_692,In_1062,In_938);
nand U693 (N_693,In_423,In_740);
nand U694 (N_694,In_1383,In_352);
or U695 (N_695,In_299,In_1911);
or U696 (N_696,In_1176,In_953);
nand U697 (N_697,In_1859,In_1174);
nand U698 (N_698,In_1510,In_913);
and U699 (N_699,In_1896,In_1479);
nand U700 (N_700,In_267,In_928);
nand U701 (N_701,In_409,In_87);
nor U702 (N_702,In_433,In_1400);
and U703 (N_703,In_653,In_253);
or U704 (N_704,In_741,In_359);
or U705 (N_705,In_1183,In_1844);
or U706 (N_706,In_1532,In_1842);
nand U707 (N_707,In_38,In_1767);
xnor U708 (N_708,In_1715,In_1456);
and U709 (N_709,In_92,In_187);
and U710 (N_710,In_543,In_1066);
or U711 (N_711,In_1557,In_478);
nor U712 (N_712,In_1269,In_1770);
nand U713 (N_713,In_226,In_773);
or U714 (N_714,In_360,In_717);
or U715 (N_715,In_1221,In_1205);
nand U716 (N_716,In_91,In_1455);
nand U717 (N_717,In_1274,In_1226);
nand U718 (N_718,In_195,In_863);
xor U719 (N_719,In_604,In_420);
or U720 (N_720,In_1548,In_1277);
nor U721 (N_721,In_1005,In_952);
nand U722 (N_722,In_1251,In_1402);
or U723 (N_723,In_882,In_645);
nand U724 (N_724,In_1297,In_601);
and U725 (N_725,In_1930,In_52);
or U726 (N_726,In_1490,In_354);
or U727 (N_727,In_1885,In_332);
and U728 (N_728,In_1195,In_95);
nor U729 (N_729,In_1850,In_286);
or U730 (N_730,In_768,In_112);
nand U731 (N_731,In_495,In_497);
nand U732 (N_732,In_1944,In_1151);
and U733 (N_733,In_1948,In_205);
nor U734 (N_734,In_1291,In_1464);
nand U735 (N_735,In_1270,In_1032);
nand U736 (N_736,In_133,In_725);
nand U737 (N_737,In_1909,In_1691);
and U738 (N_738,In_65,In_677);
or U739 (N_739,In_1080,In_1239);
xor U740 (N_740,In_925,In_828);
and U741 (N_741,In_733,In_1031);
nor U742 (N_742,In_555,In_1828);
xnor U743 (N_743,In_134,In_1377);
xnor U744 (N_744,In_1936,In_1202);
nand U745 (N_745,In_1648,In_617);
xnor U746 (N_746,In_731,In_1952);
and U747 (N_747,In_1438,In_211);
or U748 (N_748,In_1673,In_308);
nand U749 (N_749,In_1588,In_926);
nand U750 (N_750,In_1359,In_1656);
xnor U751 (N_751,In_244,In_726);
and U752 (N_752,In_1473,In_1570);
or U753 (N_753,In_1611,In_1475);
nand U754 (N_754,In_425,In_961);
nand U755 (N_755,In_1118,In_1108);
nand U756 (N_756,In_1875,In_1589);
nand U757 (N_757,In_1128,In_72);
and U758 (N_758,In_1296,In_680);
nand U759 (N_759,In_1347,In_640);
or U760 (N_760,In_991,In_506);
nand U761 (N_761,In_75,In_597);
nand U762 (N_762,In_1629,In_1133);
nand U763 (N_763,In_29,In_53);
and U764 (N_764,In_402,In_1614);
and U765 (N_765,In_1460,In_988);
or U766 (N_766,In_1664,In_268);
and U767 (N_767,In_1096,In_1929);
and U768 (N_768,In_391,In_1052);
and U769 (N_769,In_703,In_1990);
or U770 (N_770,In_243,In_296);
xnor U771 (N_771,In_603,In_1196);
nor U772 (N_772,In_1595,In_1447);
nand U773 (N_773,In_1889,In_887);
nand U774 (N_774,In_242,In_1033);
or U775 (N_775,In_471,In_963);
or U776 (N_776,In_451,In_1814);
nor U777 (N_777,In_89,In_456);
or U778 (N_778,In_930,In_1361);
nor U779 (N_779,In_1768,In_1343);
xnor U780 (N_780,In_410,In_401);
xor U781 (N_781,In_652,In_715);
xor U782 (N_782,In_1733,In_1592);
nand U783 (N_783,In_1470,In_1324);
and U784 (N_784,In_145,In_1374);
and U785 (N_785,In_813,In_646);
nand U786 (N_786,In_950,In_1725);
and U787 (N_787,In_1547,In_303);
nand U788 (N_788,In_1069,In_1585);
nand U789 (N_789,In_876,In_1529);
or U790 (N_790,In_365,In_649);
nor U791 (N_791,In_1942,In_1675);
or U792 (N_792,In_706,In_1259);
and U793 (N_793,In_317,In_1910);
nand U794 (N_794,In_1257,In_1620);
nand U795 (N_795,In_836,In_1222);
and U796 (N_796,In_363,In_1658);
nand U797 (N_797,In_1994,In_532);
nor U798 (N_798,In_329,In_7);
nor U799 (N_799,In_1817,In_689);
or U800 (N_800,In_582,In_1815);
or U801 (N_801,In_903,In_158);
and U802 (N_802,In_1549,In_1649);
or U803 (N_803,In_627,In_1058);
or U804 (N_804,In_1905,In_1117);
and U805 (N_805,In_791,In_592);
and U806 (N_806,In_1924,In_1931);
and U807 (N_807,In_31,In_1697);
or U808 (N_808,In_994,In_1810);
and U809 (N_809,In_1388,In_368);
or U810 (N_810,In_966,In_986);
nor U811 (N_811,In_1897,In_1283);
xor U812 (N_812,In_4,In_839);
and U813 (N_813,In_879,In_1110);
and U814 (N_814,In_411,In_1070);
nand U815 (N_815,In_1738,In_1698);
nand U816 (N_816,In_66,In_1575);
or U817 (N_817,In_1313,In_486);
nand U818 (N_818,In_33,In_567);
xor U819 (N_819,In_1915,In_648);
and U820 (N_820,In_1838,In_1848);
nor U821 (N_821,In_117,In_1807);
and U822 (N_822,In_1870,In_1694);
nor U823 (N_823,In_1469,In_1045);
and U824 (N_824,In_1720,In_924);
or U825 (N_825,In_1597,In_0);
and U826 (N_826,In_1160,In_1690);
and U827 (N_827,In_302,In_1865);
and U828 (N_828,In_902,In_147);
or U829 (N_829,In_945,In_919);
nor U830 (N_830,In_1284,In_1983);
or U831 (N_831,In_191,In_1373);
nor U832 (N_832,In_223,In_742);
xnor U833 (N_833,In_1252,In_917);
or U834 (N_834,In_1839,In_667);
or U835 (N_835,In_1143,In_837);
or U836 (N_836,In_144,In_1428);
nor U837 (N_837,In_1523,In_197);
or U838 (N_838,In_817,In_1149);
or U839 (N_839,In_154,In_24);
and U840 (N_840,In_26,In_906);
and U841 (N_841,In_304,In_660);
and U842 (N_842,In_609,In_1308);
xor U843 (N_843,In_1966,In_215);
nand U844 (N_844,In_22,In_106);
nor U845 (N_845,In_1111,In_457);
nand U846 (N_846,In_1501,In_880);
and U847 (N_847,In_946,In_1998);
nand U848 (N_848,In_523,In_1365);
and U849 (N_849,In_858,In_1701);
or U850 (N_850,In_819,In_1471);
nand U851 (N_851,In_83,In_918);
nand U852 (N_852,In_405,In_285);
xnor U853 (N_853,In_1262,In_1258);
nor U854 (N_854,In_1446,In_1014);
and U855 (N_855,In_1958,In_1353);
and U856 (N_856,In_311,In_1863);
xor U857 (N_857,In_366,In_663);
nor U858 (N_858,In_293,In_1439);
nor U859 (N_859,In_1016,In_279);
or U860 (N_860,In_1602,In_1789);
nor U861 (N_861,In_549,In_618);
and U862 (N_862,In_867,In_814);
or U863 (N_863,In_956,In_398);
or U864 (N_864,In_585,In_1049);
nor U865 (N_865,In_1431,In_1519);
and U866 (N_866,In_747,In_1841);
and U867 (N_867,In_217,In_527);
nor U868 (N_868,In_1459,In_904);
and U869 (N_869,In_1627,In_1876);
nand U870 (N_870,In_859,In_1727);
nand U871 (N_871,In_781,In_494);
xor U872 (N_872,In_821,In_1040);
nand U873 (N_873,In_1348,In_1407);
nand U874 (N_874,In_1043,In_282);
and U875 (N_875,In_1225,In_1866);
nor U876 (N_876,In_1256,In_54);
or U877 (N_877,In_844,In_1956);
xnor U878 (N_878,In_378,In_1097);
nor U879 (N_879,In_1962,In_539);
nor U880 (N_880,In_1429,In_1526);
xor U881 (N_881,In_1179,In_1949);
nor U882 (N_882,In_1569,In_1981);
and U883 (N_883,In_698,In_276);
xnor U884 (N_884,In_973,In_1894);
nand U885 (N_885,In_1528,In_224);
nor U886 (N_886,In_1689,In_306);
xor U887 (N_887,In_797,In_25);
nand U888 (N_888,In_1209,In_1329);
xor U889 (N_889,In_1085,In_671);
or U890 (N_890,In_958,In_426);
nand U891 (N_891,In_1778,In_1734);
nand U892 (N_892,In_1504,In_957);
or U893 (N_893,In_238,In_229);
or U894 (N_894,In_1472,In_1199);
or U895 (N_895,In_1771,In_246);
nor U896 (N_896,In_1213,In_971);
and U897 (N_897,In_602,In_169);
and U898 (N_898,In_120,In_1565);
and U899 (N_899,In_1617,In_1120);
and U900 (N_900,In_1515,In_822);
or U901 (N_901,In_940,In_1934);
and U902 (N_902,In_330,In_941);
and U903 (N_903,In_1311,In_1458);
and U904 (N_904,In_1352,In_544);
or U905 (N_905,In_50,In_910);
or U906 (N_906,In_1619,In_1281);
nor U907 (N_907,In_716,In_1762);
nand U908 (N_908,In_690,In_307);
nand U909 (N_909,In_1410,In_1615);
or U910 (N_910,In_461,In_1409);
xor U911 (N_911,In_166,In_808);
nand U912 (N_912,In_1703,In_1953);
nand U913 (N_913,In_1351,In_1104);
or U914 (N_914,In_1292,In_452);
nor U915 (N_915,In_1912,In_1666);
nand U916 (N_916,In_125,In_295);
xnor U917 (N_917,In_674,In_1095);
nand U918 (N_918,In_1811,In_1107);
or U919 (N_919,In_1583,In_1175);
nand U920 (N_920,In_1667,In_784);
and U921 (N_921,In_80,In_2);
xnor U922 (N_922,In_1882,In_1408);
and U923 (N_923,In_1190,In_682);
or U924 (N_924,In_413,In_1486);
nand U925 (N_925,In_1537,In_127);
and U926 (N_926,In_444,In_1660);
nand U927 (N_927,In_1384,In_339);
nand U928 (N_928,In_196,In_744);
nor U929 (N_929,In_96,In_502);
or U930 (N_930,In_1641,In_1645);
or U931 (N_931,In_623,In_1772);
nor U932 (N_932,In_1969,In_412);
and U933 (N_933,In_1635,In_272);
nor U934 (N_934,In_1309,In_948);
nor U935 (N_935,In_184,In_214);
nand U936 (N_936,In_631,In_1002);
or U937 (N_937,In_355,In_834);
nor U938 (N_938,In_1867,In_103);
and U939 (N_939,In_775,In_1749);
nor U940 (N_940,In_181,In_1964);
and U941 (N_941,In_699,In_589);
and U942 (N_942,In_713,In_1808);
or U943 (N_943,In_883,In_577);
nand U944 (N_944,In_1011,In_1100);
and U945 (N_945,In_1224,In_697);
or U946 (N_946,In_44,In_878);
xor U947 (N_947,In_484,In_1041);
nor U948 (N_948,In_1993,In_453);
and U949 (N_949,In_685,In_57);
nor U950 (N_950,In_864,In_666);
nand U951 (N_951,In_970,In_771);
and U952 (N_952,In_712,In_153);
and U953 (N_953,In_764,In_473);
nor U954 (N_954,In_1044,In_1073);
or U955 (N_955,In_1192,In_1344);
or U956 (N_956,In_76,In_1271);
nand U957 (N_957,In_1272,In_1536);
or U958 (N_958,In_1978,In_1659);
and U959 (N_959,In_977,In_1672);
nor U960 (N_960,In_1304,In_1261);
nor U961 (N_961,In_64,In_873);
or U962 (N_962,In_1207,In_1852);
nor U963 (N_963,In_1970,In_1502);
or U964 (N_964,In_1370,In_459);
nor U965 (N_965,In_1827,In_393);
or U966 (N_966,In_78,In_736);
nor U967 (N_967,In_1362,In_1920);
and U968 (N_968,In_1478,In_766);
nand U969 (N_969,In_300,In_1462);
and U970 (N_970,In_488,In_1606);
and U971 (N_971,In_1423,In_820);
nand U972 (N_972,In_199,In_1035);
nor U973 (N_973,In_1908,In_888);
and U974 (N_974,In_1386,In_1452);
and U975 (N_975,In_283,In_684);
nand U976 (N_976,In_1818,In_472);
and U977 (N_977,In_98,In_871);
and U978 (N_978,In_298,In_1991);
nand U979 (N_979,In_190,In_88);
nor U980 (N_980,In_231,In_1491);
and U981 (N_981,In_174,In_554);
or U982 (N_982,In_1760,In_1845);
or U983 (N_983,In_435,In_1988);
or U984 (N_984,In_364,In_1975);
nand U985 (N_985,In_509,In_1454);
nor U986 (N_986,In_1886,In_738);
nor U987 (N_987,In_1921,In_1806);
or U988 (N_988,In_493,In_182);
and U989 (N_989,In_1342,In_1832);
and U990 (N_990,In_1346,In_1161);
nor U991 (N_991,In_1493,In_1788);
nor U992 (N_992,In_1989,In_1805);
nor U993 (N_993,In_40,In_119);
nor U994 (N_994,In_1567,In_397);
or U995 (N_995,In_1545,In_1);
and U996 (N_996,In_101,In_1007);
nor U997 (N_997,In_1323,In_533);
and U998 (N_998,In_1223,In_798);
or U999 (N_999,In_310,In_1783);
nor U1000 (N_1000,In_410,In_172);
xnor U1001 (N_1001,In_300,In_603);
or U1002 (N_1002,In_1141,In_1572);
nor U1003 (N_1003,In_1614,In_1760);
nor U1004 (N_1004,In_1566,In_461);
nor U1005 (N_1005,In_1475,In_533);
nor U1006 (N_1006,In_331,In_888);
xnor U1007 (N_1007,In_71,In_79);
or U1008 (N_1008,In_1838,In_195);
nand U1009 (N_1009,In_1618,In_799);
xnor U1010 (N_1010,In_1733,In_1850);
nand U1011 (N_1011,In_1682,In_821);
or U1012 (N_1012,In_1065,In_1455);
or U1013 (N_1013,In_152,In_1240);
nand U1014 (N_1014,In_41,In_265);
and U1015 (N_1015,In_795,In_699);
nor U1016 (N_1016,In_419,In_151);
nand U1017 (N_1017,In_1086,In_974);
nand U1018 (N_1018,In_416,In_1550);
or U1019 (N_1019,In_1031,In_82);
or U1020 (N_1020,In_89,In_126);
or U1021 (N_1021,In_1582,In_700);
nor U1022 (N_1022,In_127,In_1084);
nand U1023 (N_1023,In_1831,In_1268);
nor U1024 (N_1024,In_677,In_1403);
and U1025 (N_1025,In_1233,In_20);
and U1026 (N_1026,In_226,In_1212);
nand U1027 (N_1027,In_821,In_1853);
or U1028 (N_1028,In_1322,In_1750);
nor U1029 (N_1029,In_418,In_975);
and U1030 (N_1030,In_190,In_1609);
xnor U1031 (N_1031,In_371,In_38);
nor U1032 (N_1032,In_65,In_405);
or U1033 (N_1033,In_1718,In_725);
nor U1034 (N_1034,In_779,In_1288);
xnor U1035 (N_1035,In_1719,In_1162);
nor U1036 (N_1036,In_1453,In_1782);
or U1037 (N_1037,In_27,In_1051);
nand U1038 (N_1038,In_1956,In_24);
nor U1039 (N_1039,In_359,In_651);
nand U1040 (N_1040,In_1214,In_1405);
or U1041 (N_1041,In_57,In_1145);
xor U1042 (N_1042,In_834,In_975);
xor U1043 (N_1043,In_1021,In_760);
or U1044 (N_1044,In_87,In_700);
and U1045 (N_1045,In_867,In_454);
nand U1046 (N_1046,In_739,In_558);
or U1047 (N_1047,In_873,In_192);
and U1048 (N_1048,In_1678,In_1609);
and U1049 (N_1049,In_278,In_328);
or U1050 (N_1050,In_1225,In_1322);
and U1051 (N_1051,In_1288,In_1583);
or U1052 (N_1052,In_1301,In_31);
nand U1053 (N_1053,In_238,In_577);
and U1054 (N_1054,In_1185,In_1677);
nand U1055 (N_1055,In_1140,In_453);
nand U1056 (N_1056,In_1797,In_1503);
and U1057 (N_1057,In_1658,In_950);
and U1058 (N_1058,In_235,In_245);
xnor U1059 (N_1059,In_1395,In_915);
nor U1060 (N_1060,In_1918,In_1098);
nand U1061 (N_1061,In_1194,In_36);
and U1062 (N_1062,In_1378,In_434);
and U1063 (N_1063,In_1825,In_842);
nand U1064 (N_1064,In_758,In_244);
or U1065 (N_1065,In_1491,In_1426);
and U1066 (N_1066,In_384,In_585);
or U1067 (N_1067,In_435,In_1311);
xnor U1068 (N_1068,In_1150,In_1303);
or U1069 (N_1069,In_1650,In_571);
or U1070 (N_1070,In_1407,In_973);
nor U1071 (N_1071,In_1935,In_534);
nor U1072 (N_1072,In_206,In_1466);
nand U1073 (N_1073,In_1675,In_450);
and U1074 (N_1074,In_689,In_728);
xor U1075 (N_1075,In_1089,In_989);
nand U1076 (N_1076,In_1254,In_1774);
nand U1077 (N_1077,In_806,In_1559);
and U1078 (N_1078,In_1511,In_168);
or U1079 (N_1079,In_1799,In_183);
xnor U1080 (N_1080,In_1138,In_919);
nor U1081 (N_1081,In_1783,In_2);
nor U1082 (N_1082,In_1480,In_1537);
xnor U1083 (N_1083,In_11,In_250);
nand U1084 (N_1084,In_1407,In_1318);
nand U1085 (N_1085,In_252,In_1538);
nor U1086 (N_1086,In_394,In_1252);
and U1087 (N_1087,In_873,In_681);
nand U1088 (N_1088,In_336,In_1699);
and U1089 (N_1089,In_869,In_894);
and U1090 (N_1090,In_908,In_1874);
nor U1091 (N_1091,In_1982,In_464);
nand U1092 (N_1092,In_183,In_1760);
and U1093 (N_1093,In_1634,In_1620);
xor U1094 (N_1094,In_1743,In_33);
nor U1095 (N_1095,In_1375,In_1478);
or U1096 (N_1096,In_693,In_179);
and U1097 (N_1097,In_471,In_731);
nand U1098 (N_1098,In_1965,In_1442);
or U1099 (N_1099,In_1096,In_1607);
or U1100 (N_1100,In_915,In_138);
and U1101 (N_1101,In_1796,In_319);
and U1102 (N_1102,In_409,In_544);
nor U1103 (N_1103,In_1169,In_762);
and U1104 (N_1104,In_986,In_983);
nand U1105 (N_1105,In_1833,In_690);
nor U1106 (N_1106,In_475,In_1557);
nor U1107 (N_1107,In_1474,In_1378);
or U1108 (N_1108,In_1423,In_937);
or U1109 (N_1109,In_1458,In_1371);
xor U1110 (N_1110,In_1042,In_707);
xor U1111 (N_1111,In_878,In_905);
xor U1112 (N_1112,In_201,In_1495);
xnor U1113 (N_1113,In_1424,In_1365);
nand U1114 (N_1114,In_910,In_46);
or U1115 (N_1115,In_1469,In_1618);
nor U1116 (N_1116,In_244,In_836);
or U1117 (N_1117,In_849,In_1533);
or U1118 (N_1118,In_159,In_322);
and U1119 (N_1119,In_1823,In_721);
nor U1120 (N_1120,In_1633,In_246);
and U1121 (N_1121,In_1059,In_404);
nor U1122 (N_1122,In_702,In_1771);
and U1123 (N_1123,In_1453,In_1705);
or U1124 (N_1124,In_1657,In_347);
or U1125 (N_1125,In_1440,In_1572);
or U1126 (N_1126,In_412,In_1960);
and U1127 (N_1127,In_683,In_1235);
xnor U1128 (N_1128,In_161,In_1800);
or U1129 (N_1129,In_673,In_999);
and U1130 (N_1130,In_1095,In_235);
and U1131 (N_1131,In_454,In_1538);
nor U1132 (N_1132,In_1660,In_1084);
or U1133 (N_1133,In_634,In_1010);
nor U1134 (N_1134,In_519,In_631);
nand U1135 (N_1135,In_4,In_435);
nand U1136 (N_1136,In_1515,In_1805);
and U1137 (N_1137,In_0,In_1044);
and U1138 (N_1138,In_1327,In_1808);
and U1139 (N_1139,In_1203,In_369);
or U1140 (N_1140,In_1628,In_819);
and U1141 (N_1141,In_50,In_825);
or U1142 (N_1142,In_545,In_384);
nand U1143 (N_1143,In_1144,In_691);
or U1144 (N_1144,In_1393,In_1136);
and U1145 (N_1145,In_1668,In_330);
nand U1146 (N_1146,In_1472,In_1754);
nand U1147 (N_1147,In_1613,In_890);
or U1148 (N_1148,In_1799,In_1297);
xnor U1149 (N_1149,In_1958,In_674);
or U1150 (N_1150,In_1209,In_1534);
xor U1151 (N_1151,In_812,In_1901);
xnor U1152 (N_1152,In_1252,In_135);
and U1153 (N_1153,In_276,In_397);
nand U1154 (N_1154,In_949,In_1161);
nand U1155 (N_1155,In_289,In_1415);
or U1156 (N_1156,In_218,In_1405);
or U1157 (N_1157,In_912,In_93);
or U1158 (N_1158,In_359,In_1104);
and U1159 (N_1159,In_168,In_806);
or U1160 (N_1160,In_181,In_544);
nand U1161 (N_1161,In_1357,In_1654);
and U1162 (N_1162,In_1162,In_1026);
xnor U1163 (N_1163,In_1003,In_1097);
and U1164 (N_1164,In_1211,In_1378);
nor U1165 (N_1165,In_1868,In_1171);
xnor U1166 (N_1166,In_766,In_862);
nand U1167 (N_1167,In_119,In_103);
nand U1168 (N_1168,In_1775,In_767);
nand U1169 (N_1169,In_489,In_1942);
or U1170 (N_1170,In_146,In_1575);
or U1171 (N_1171,In_0,In_643);
nand U1172 (N_1172,In_525,In_609);
nor U1173 (N_1173,In_573,In_1086);
or U1174 (N_1174,In_1220,In_476);
and U1175 (N_1175,In_1606,In_502);
nand U1176 (N_1176,In_1368,In_1256);
or U1177 (N_1177,In_1955,In_1398);
nor U1178 (N_1178,In_1979,In_1864);
and U1179 (N_1179,In_158,In_496);
xor U1180 (N_1180,In_1413,In_1838);
or U1181 (N_1181,In_325,In_1337);
nor U1182 (N_1182,In_15,In_1008);
nor U1183 (N_1183,In_579,In_1255);
xor U1184 (N_1184,In_1854,In_1401);
or U1185 (N_1185,In_787,In_908);
and U1186 (N_1186,In_637,In_773);
or U1187 (N_1187,In_1695,In_527);
nand U1188 (N_1188,In_1282,In_382);
and U1189 (N_1189,In_846,In_1717);
and U1190 (N_1190,In_1559,In_486);
nand U1191 (N_1191,In_1940,In_479);
nand U1192 (N_1192,In_46,In_245);
nor U1193 (N_1193,In_60,In_65);
or U1194 (N_1194,In_538,In_1225);
nand U1195 (N_1195,In_1929,In_1742);
nand U1196 (N_1196,In_1321,In_1162);
or U1197 (N_1197,In_1838,In_1323);
xnor U1198 (N_1198,In_1366,In_485);
or U1199 (N_1199,In_1263,In_1113);
nor U1200 (N_1200,In_1802,In_178);
xor U1201 (N_1201,In_1158,In_1400);
or U1202 (N_1202,In_168,In_407);
and U1203 (N_1203,In_1260,In_993);
nand U1204 (N_1204,In_1835,In_1696);
nand U1205 (N_1205,In_1752,In_695);
nand U1206 (N_1206,In_1946,In_1738);
and U1207 (N_1207,In_1549,In_284);
or U1208 (N_1208,In_1574,In_1549);
nor U1209 (N_1209,In_1157,In_1310);
xor U1210 (N_1210,In_1398,In_420);
or U1211 (N_1211,In_1799,In_455);
and U1212 (N_1212,In_490,In_1734);
and U1213 (N_1213,In_1104,In_1987);
and U1214 (N_1214,In_1199,In_1825);
nand U1215 (N_1215,In_1313,In_18);
or U1216 (N_1216,In_728,In_790);
nor U1217 (N_1217,In_504,In_1062);
and U1218 (N_1218,In_27,In_1119);
nor U1219 (N_1219,In_1486,In_546);
nor U1220 (N_1220,In_605,In_216);
and U1221 (N_1221,In_1458,In_241);
nor U1222 (N_1222,In_1687,In_1063);
xor U1223 (N_1223,In_1799,In_1278);
and U1224 (N_1224,In_1276,In_49);
nor U1225 (N_1225,In_628,In_1891);
nor U1226 (N_1226,In_1130,In_733);
and U1227 (N_1227,In_1112,In_1270);
nor U1228 (N_1228,In_1999,In_1114);
nor U1229 (N_1229,In_392,In_1941);
nor U1230 (N_1230,In_1163,In_1544);
nand U1231 (N_1231,In_853,In_1922);
nor U1232 (N_1232,In_985,In_1032);
nand U1233 (N_1233,In_276,In_1564);
xor U1234 (N_1234,In_618,In_1103);
or U1235 (N_1235,In_50,In_1134);
nor U1236 (N_1236,In_767,In_1418);
nand U1237 (N_1237,In_1579,In_534);
or U1238 (N_1238,In_814,In_1819);
xnor U1239 (N_1239,In_1445,In_376);
nor U1240 (N_1240,In_1263,In_1859);
nor U1241 (N_1241,In_1423,In_1265);
nor U1242 (N_1242,In_331,In_1525);
and U1243 (N_1243,In_473,In_384);
nand U1244 (N_1244,In_688,In_1146);
and U1245 (N_1245,In_50,In_790);
nor U1246 (N_1246,In_498,In_595);
or U1247 (N_1247,In_1677,In_9);
nor U1248 (N_1248,In_1639,In_307);
nand U1249 (N_1249,In_58,In_1285);
and U1250 (N_1250,In_1492,In_629);
and U1251 (N_1251,In_1936,In_71);
or U1252 (N_1252,In_487,In_514);
nand U1253 (N_1253,In_1474,In_814);
and U1254 (N_1254,In_741,In_1330);
nand U1255 (N_1255,In_345,In_861);
nor U1256 (N_1256,In_1439,In_88);
and U1257 (N_1257,In_541,In_545);
or U1258 (N_1258,In_947,In_814);
nand U1259 (N_1259,In_343,In_1375);
nand U1260 (N_1260,In_1104,In_928);
nand U1261 (N_1261,In_1827,In_1436);
xor U1262 (N_1262,In_272,In_137);
or U1263 (N_1263,In_1847,In_1970);
and U1264 (N_1264,In_1221,In_12);
and U1265 (N_1265,In_1704,In_1306);
and U1266 (N_1266,In_1897,In_1886);
nand U1267 (N_1267,In_1546,In_610);
xnor U1268 (N_1268,In_152,In_1476);
nor U1269 (N_1269,In_1699,In_1179);
and U1270 (N_1270,In_927,In_1473);
or U1271 (N_1271,In_535,In_974);
nand U1272 (N_1272,In_1996,In_42);
nor U1273 (N_1273,In_961,In_1325);
nand U1274 (N_1274,In_130,In_1891);
or U1275 (N_1275,In_600,In_1736);
nor U1276 (N_1276,In_1631,In_196);
nand U1277 (N_1277,In_329,In_826);
xnor U1278 (N_1278,In_1818,In_416);
and U1279 (N_1279,In_1094,In_1382);
and U1280 (N_1280,In_1796,In_757);
or U1281 (N_1281,In_1562,In_982);
nor U1282 (N_1282,In_1548,In_1686);
nand U1283 (N_1283,In_1780,In_371);
nand U1284 (N_1284,In_1415,In_1817);
nand U1285 (N_1285,In_1987,In_1070);
or U1286 (N_1286,In_1913,In_889);
nand U1287 (N_1287,In_280,In_1594);
or U1288 (N_1288,In_943,In_46);
nor U1289 (N_1289,In_1956,In_789);
or U1290 (N_1290,In_1626,In_1220);
and U1291 (N_1291,In_1993,In_677);
nand U1292 (N_1292,In_748,In_480);
nand U1293 (N_1293,In_1800,In_588);
nand U1294 (N_1294,In_1810,In_1625);
nand U1295 (N_1295,In_1341,In_1512);
and U1296 (N_1296,In_900,In_378);
xnor U1297 (N_1297,In_1026,In_850);
xnor U1298 (N_1298,In_1279,In_129);
xnor U1299 (N_1299,In_1354,In_966);
nor U1300 (N_1300,In_1783,In_33);
nand U1301 (N_1301,In_1280,In_1762);
and U1302 (N_1302,In_1080,In_1060);
nand U1303 (N_1303,In_429,In_739);
and U1304 (N_1304,In_444,In_1141);
nand U1305 (N_1305,In_1730,In_334);
xnor U1306 (N_1306,In_1375,In_259);
or U1307 (N_1307,In_570,In_1691);
nor U1308 (N_1308,In_198,In_58);
nor U1309 (N_1309,In_1109,In_1324);
nor U1310 (N_1310,In_1470,In_132);
or U1311 (N_1311,In_1442,In_863);
nand U1312 (N_1312,In_1662,In_1520);
xnor U1313 (N_1313,In_1647,In_1995);
and U1314 (N_1314,In_439,In_1073);
nand U1315 (N_1315,In_444,In_654);
and U1316 (N_1316,In_1563,In_1101);
nand U1317 (N_1317,In_1941,In_237);
nor U1318 (N_1318,In_456,In_606);
nand U1319 (N_1319,In_460,In_1437);
xor U1320 (N_1320,In_1387,In_1335);
nor U1321 (N_1321,In_376,In_543);
or U1322 (N_1322,In_694,In_283);
or U1323 (N_1323,In_32,In_296);
or U1324 (N_1324,In_1747,In_1839);
nor U1325 (N_1325,In_154,In_1521);
nor U1326 (N_1326,In_667,In_703);
and U1327 (N_1327,In_610,In_77);
nor U1328 (N_1328,In_165,In_789);
xnor U1329 (N_1329,In_1308,In_872);
nor U1330 (N_1330,In_1794,In_1088);
nor U1331 (N_1331,In_537,In_83);
nand U1332 (N_1332,In_456,In_179);
and U1333 (N_1333,In_1937,In_1958);
and U1334 (N_1334,In_932,In_1981);
or U1335 (N_1335,In_1388,In_229);
and U1336 (N_1336,In_737,In_1142);
and U1337 (N_1337,In_1559,In_249);
and U1338 (N_1338,In_1226,In_671);
nor U1339 (N_1339,In_672,In_974);
xor U1340 (N_1340,In_976,In_359);
nor U1341 (N_1341,In_562,In_1437);
and U1342 (N_1342,In_677,In_1446);
and U1343 (N_1343,In_1550,In_89);
and U1344 (N_1344,In_112,In_32);
nor U1345 (N_1345,In_1713,In_128);
nand U1346 (N_1346,In_1369,In_1915);
or U1347 (N_1347,In_724,In_1987);
and U1348 (N_1348,In_1538,In_755);
or U1349 (N_1349,In_1595,In_975);
nand U1350 (N_1350,In_1054,In_1588);
xnor U1351 (N_1351,In_707,In_236);
nand U1352 (N_1352,In_532,In_364);
and U1353 (N_1353,In_1603,In_60);
nor U1354 (N_1354,In_343,In_1203);
or U1355 (N_1355,In_598,In_233);
or U1356 (N_1356,In_794,In_611);
nor U1357 (N_1357,In_236,In_515);
and U1358 (N_1358,In_316,In_1796);
or U1359 (N_1359,In_929,In_1349);
nor U1360 (N_1360,In_1654,In_422);
nand U1361 (N_1361,In_1519,In_945);
nor U1362 (N_1362,In_1531,In_904);
nand U1363 (N_1363,In_690,In_303);
nand U1364 (N_1364,In_1181,In_264);
nor U1365 (N_1365,In_448,In_1121);
and U1366 (N_1366,In_33,In_546);
nand U1367 (N_1367,In_1625,In_947);
and U1368 (N_1368,In_204,In_578);
and U1369 (N_1369,In_314,In_1510);
xnor U1370 (N_1370,In_1963,In_1501);
nor U1371 (N_1371,In_1508,In_539);
or U1372 (N_1372,In_135,In_468);
or U1373 (N_1373,In_1479,In_71);
nand U1374 (N_1374,In_1379,In_1431);
or U1375 (N_1375,In_723,In_73);
or U1376 (N_1376,In_876,In_993);
or U1377 (N_1377,In_995,In_244);
or U1378 (N_1378,In_1412,In_245);
nand U1379 (N_1379,In_1982,In_284);
or U1380 (N_1380,In_352,In_501);
or U1381 (N_1381,In_1625,In_435);
or U1382 (N_1382,In_751,In_118);
nand U1383 (N_1383,In_1050,In_1792);
nor U1384 (N_1384,In_1268,In_1104);
or U1385 (N_1385,In_72,In_1146);
or U1386 (N_1386,In_1931,In_1852);
or U1387 (N_1387,In_381,In_1122);
nand U1388 (N_1388,In_720,In_668);
nand U1389 (N_1389,In_1456,In_478);
and U1390 (N_1390,In_1657,In_842);
nand U1391 (N_1391,In_524,In_1597);
nand U1392 (N_1392,In_400,In_1822);
or U1393 (N_1393,In_909,In_257);
nor U1394 (N_1394,In_864,In_809);
or U1395 (N_1395,In_1288,In_1174);
xnor U1396 (N_1396,In_1387,In_1116);
and U1397 (N_1397,In_456,In_700);
nor U1398 (N_1398,In_1546,In_258);
nand U1399 (N_1399,In_665,In_300);
nand U1400 (N_1400,In_1347,In_1281);
nor U1401 (N_1401,In_767,In_1127);
nand U1402 (N_1402,In_834,In_843);
nor U1403 (N_1403,In_1479,In_846);
and U1404 (N_1404,In_437,In_651);
xnor U1405 (N_1405,In_77,In_797);
nor U1406 (N_1406,In_999,In_1260);
and U1407 (N_1407,In_993,In_1948);
and U1408 (N_1408,In_921,In_945);
nor U1409 (N_1409,In_398,In_2);
nor U1410 (N_1410,In_1158,In_465);
nand U1411 (N_1411,In_1297,In_1316);
and U1412 (N_1412,In_773,In_202);
xnor U1413 (N_1413,In_685,In_1256);
nand U1414 (N_1414,In_218,In_661);
nor U1415 (N_1415,In_24,In_1292);
and U1416 (N_1416,In_1442,In_892);
or U1417 (N_1417,In_1764,In_926);
nand U1418 (N_1418,In_1023,In_236);
nand U1419 (N_1419,In_1227,In_1847);
or U1420 (N_1420,In_1584,In_1764);
or U1421 (N_1421,In_844,In_1602);
nor U1422 (N_1422,In_1438,In_1529);
xnor U1423 (N_1423,In_1651,In_336);
or U1424 (N_1424,In_1648,In_986);
nor U1425 (N_1425,In_349,In_780);
nor U1426 (N_1426,In_143,In_784);
or U1427 (N_1427,In_1559,In_1641);
or U1428 (N_1428,In_89,In_179);
or U1429 (N_1429,In_478,In_582);
nand U1430 (N_1430,In_1866,In_472);
nor U1431 (N_1431,In_344,In_391);
nand U1432 (N_1432,In_663,In_1136);
nor U1433 (N_1433,In_1119,In_1168);
nor U1434 (N_1434,In_594,In_673);
nand U1435 (N_1435,In_509,In_1039);
or U1436 (N_1436,In_1676,In_104);
nand U1437 (N_1437,In_925,In_1480);
nor U1438 (N_1438,In_1567,In_714);
nand U1439 (N_1439,In_1187,In_1043);
or U1440 (N_1440,In_819,In_539);
or U1441 (N_1441,In_1567,In_1409);
and U1442 (N_1442,In_143,In_186);
xnor U1443 (N_1443,In_1606,In_148);
nor U1444 (N_1444,In_542,In_1982);
or U1445 (N_1445,In_1540,In_659);
nor U1446 (N_1446,In_269,In_307);
nand U1447 (N_1447,In_721,In_1283);
or U1448 (N_1448,In_1537,In_822);
or U1449 (N_1449,In_759,In_397);
nor U1450 (N_1450,In_1986,In_650);
nor U1451 (N_1451,In_1990,In_1746);
nand U1452 (N_1452,In_290,In_1587);
and U1453 (N_1453,In_515,In_1288);
nand U1454 (N_1454,In_1306,In_444);
nor U1455 (N_1455,In_232,In_1335);
or U1456 (N_1456,In_1548,In_408);
and U1457 (N_1457,In_996,In_1906);
or U1458 (N_1458,In_796,In_329);
nor U1459 (N_1459,In_1602,In_469);
nand U1460 (N_1460,In_916,In_1917);
or U1461 (N_1461,In_1752,In_1152);
and U1462 (N_1462,In_1254,In_1599);
or U1463 (N_1463,In_525,In_218);
xor U1464 (N_1464,In_691,In_26);
nor U1465 (N_1465,In_492,In_1710);
nor U1466 (N_1466,In_1543,In_1140);
and U1467 (N_1467,In_982,In_14);
and U1468 (N_1468,In_1340,In_851);
and U1469 (N_1469,In_87,In_1462);
or U1470 (N_1470,In_74,In_1384);
and U1471 (N_1471,In_1683,In_552);
or U1472 (N_1472,In_574,In_675);
xor U1473 (N_1473,In_1585,In_681);
and U1474 (N_1474,In_904,In_73);
nor U1475 (N_1475,In_1021,In_582);
nand U1476 (N_1476,In_1555,In_154);
xor U1477 (N_1477,In_705,In_29);
nor U1478 (N_1478,In_877,In_1412);
or U1479 (N_1479,In_1125,In_1711);
nand U1480 (N_1480,In_1030,In_508);
and U1481 (N_1481,In_1675,In_1562);
and U1482 (N_1482,In_547,In_1428);
xor U1483 (N_1483,In_1656,In_1329);
nand U1484 (N_1484,In_983,In_521);
and U1485 (N_1485,In_404,In_1215);
or U1486 (N_1486,In_1922,In_713);
and U1487 (N_1487,In_825,In_40);
and U1488 (N_1488,In_60,In_1846);
and U1489 (N_1489,In_1016,In_1208);
nor U1490 (N_1490,In_1865,In_626);
or U1491 (N_1491,In_287,In_132);
and U1492 (N_1492,In_995,In_27);
nand U1493 (N_1493,In_1140,In_52);
or U1494 (N_1494,In_302,In_1307);
nand U1495 (N_1495,In_1510,In_966);
nor U1496 (N_1496,In_1888,In_1328);
nor U1497 (N_1497,In_1774,In_986);
and U1498 (N_1498,In_307,In_988);
and U1499 (N_1499,In_1778,In_1652);
nor U1500 (N_1500,In_653,In_883);
nand U1501 (N_1501,In_908,In_962);
nand U1502 (N_1502,In_431,In_1258);
nor U1503 (N_1503,In_579,In_1561);
or U1504 (N_1504,In_1948,In_317);
and U1505 (N_1505,In_1888,In_244);
nand U1506 (N_1506,In_1820,In_731);
xnor U1507 (N_1507,In_214,In_1500);
nor U1508 (N_1508,In_800,In_873);
or U1509 (N_1509,In_647,In_1378);
nand U1510 (N_1510,In_1682,In_1470);
and U1511 (N_1511,In_1262,In_1122);
or U1512 (N_1512,In_752,In_1272);
or U1513 (N_1513,In_1057,In_113);
nor U1514 (N_1514,In_623,In_1924);
nor U1515 (N_1515,In_1866,In_291);
xor U1516 (N_1516,In_729,In_1036);
or U1517 (N_1517,In_1299,In_235);
or U1518 (N_1518,In_262,In_238);
or U1519 (N_1519,In_1345,In_660);
and U1520 (N_1520,In_1125,In_464);
or U1521 (N_1521,In_856,In_1208);
or U1522 (N_1522,In_1147,In_449);
and U1523 (N_1523,In_582,In_670);
xor U1524 (N_1524,In_245,In_1889);
nor U1525 (N_1525,In_121,In_694);
nor U1526 (N_1526,In_937,In_33);
nand U1527 (N_1527,In_1942,In_926);
or U1528 (N_1528,In_1935,In_959);
or U1529 (N_1529,In_599,In_208);
nor U1530 (N_1530,In_739,In_249);
xnor U1531 (N_1531,In_2,In_499);
and U1532 (N_1532,In_1717,In_1854);
xor U1533 (N_1533,In_1877,In_460);
nand U1534 (N_1534,In_688,In_718);
nor U1535 (N_1535,In_1737,In_1433);
and U1536 (N_1536,In_604,In_1440);
nor U1537 (N_1537,In_857,In_1464);
and U1538 (N_1538,In_1875,In_227);
xor U1539 (N_1539,In_1642,In_1924);
or U1540 (N_1540,In_138,In_1726);
and U1541 (N_1541,In_970,In_1076);
nand U1542 (N_1542,In_1542,In_695);
nand U1543 (N_1543,In_1833,In_133);
xnor U1544 (N_1544,In_763,In_352);
xnor U1545 (N_1545,In_324,In_1754);
nand U1546 (N_1546,In_1547,In_1557);
nor U1547 (N_1547,In_239,In_1257);
nand U1548 (N_1548,In_439,In_197);
or U1549 (N_1549,In_232,In_1252);
nor U1550 (N_1550,In_1762,In_1412);
nor U1551 (N_1551,In_1205,In_1858);
or U1552 (N_1552,In_1568,In_240);
nand U1553 (N_1553,In_271,In_1284);
nand U1554 (N_1554,In_1181,In_916);
nor U1555 (N_1555,In_627,In_1288);
or U1556 (N_1556,In_919,In_549);
nand U1557 (N_1557,In_1137,In_1197);
and U1558 (N_1558,In_1622,In_1852);
nor U1559 (N_1559,In_838,In_479);
xor U1560 (N_1560,In_1431,In_1020);
nand U1561 (N_1561,In_40,In_1108);
or U1562 (N_1562,In_1808,In_819);
and U1563 (N_1563,In_1728,In_1802);
nand U1564 (N_1564,In_472,In_922);
and U1565 (N_1565,In_694,In_1766);
nand U1566 (N_1566,In_1444,In_1959);
or U1567 (N_1567,In_914,In_1545);
nand U1568 (N_1568,In_861,In_1527);
nand U1569 (N_1569,In_875,In_1637);
or U1570 (N_1570,In_1947,In_1426);
and U1571 (N_1571,In_390,In_1343);
or U1572 (N_1572,In_1352,In_856);
or U1573 (N_1573,In_843,In_1024);
nand U1574 (N_1574,In_1611,In_1508);
and U1575 (N_1575,In_1849,In_375);
and U1576 (N_1576,In_711,In_953);
nor U1577 (N_1577,In_1754,In_1179);
and U1578 (N_1578,In_1624,In_154);
or U1579 (N_1579,In_1264,In_714);
nor U1580 (N_1580,In_287,In_828);
nor U1581 (N_1581,In_1099,In_1319);
nand U1582 (N_1582,In_425,In_1072);
nand U1583 (N_1583,In_1749,In_1500);
or U1584 (N_1584,In_1492,In_1225);
xor U1585 (N_1585,In_63,In_41);
and U1586 (N_1586,In_1431,In_232);
and U1587 (N_1587,In_305,In_917);
nand U1588 (N_1588,In_864,In_1328);
or U1589 (N_1589,In_63,In_1876);
or U1590 (N_1590,In_34,In_1539);
xor U1591 (N_1591,In_1013,In_283);
nand U1592 (N_1592,In_1915,In_1729);
and U1593 (N_1593,In_104,In_253);
nand U1594 (N_1594,In_267,In_1222);
and U1595 (N_1595,In_527,In_1607);
xor U1596 (N_1596,In_1989,In_526);
and U1597 (N_1597,In_1893,In_428);
xnor U1598 (N_1598,In_1071,In_1509);
nor U1599 (N_1599,In_1760,In_1606);
or U1600 (N_1600,In_412,In_656);
xnor U1601 (N_1601,In_698,In_1779);
nor U1602 (N_1602,In_1113,In_1407);
nor U1603 (N_1603,In_439,In_231);
nor U1604 (N_1604,In_159,In_300);
nand U1605 (N_1605,In_1453,In_30);
or U1606 (N_1606,In_1337,In_1634);
nor U1607 (N_1607,In_885,In_251);
and U1608 (N_1608,In_1181,In_80);
nand U1609 (N_1609,In_1052,In_1334);
nor U1610 (N_1610,In_1318,In_1482);
or U1611 (N_1611,In_1456,In_661);
and U1612 (N_1612,In_613,In_69);
and U1613 (N_1613,In_762,In_1447);
nor U1614 (N_1614,In_571,In_1895);
and U1615 (N_1615,In_366,In_1172);
nor U1616 (N_1616,In_1228,In_482);
and U1617 (N_1617,In_1117,In_1941);
and U1618 (N_1618,In_439,In_1775);
or U1619 (N_1619,In_1441,In_191);
and U1620 (N_1620,In_208,In_1982);
nor U1621 (N_1621,In_1749,In_1852);
or U1622 (N_1622,In_1751,In_1355);
and U1623 (N_1623,In_1763,In_57);
or U1624 (N_1624,In_184,In_1043);
nand U1625 (N_1625,In_1177,In_1639);
nor U1626 (N_1626,In_125,In_211);
or U1627 (N_1627,In_1727,In_97);
nor U1628 (N_1628,In_28,In_643);
nand U1629 (N_1629,In_891,In_1861);
nor U1630 (N_1630,In_1744,In_56);
or U1631 (N_1631,In_1170,In_1096);
nor U1632 (N_1632,In_74,In_1989);
or U1633 (N_1633,In_1442,In_453);
or U1634 (N_1634,In_1406,In_364);
and U1635 (N_1635,In_1892,In_1898);
and U1636 (N_1636,In_743,In_137);
nor U1637 (N_1637,In_1835,In_629);
xor U1638 (N_1638,In_897,In_354);
nand U1639 (N_1639,In_1243,In_325);
and U1640 (N_1640,In_126,In_1466);
nand U1641 (N_1641,In_1139,In_379);
nand U1642 (N_1642,In_1071,In_1800);
and U1643 (N_1643,In_525,In_980);
nor U1644 (N_1644,In_623,In_1257);
nand U1645 (N_1645,In_406,In_1813);
xnor U1646 (N_1646,In_122,In_1959);
or U1647 (N_1647,In_1136,In_937);
nor U1648 (N_1648,In_172,In_1454);
and U1649 (N_1649,In_428,In_1614);
nor U1650 (N_1650,In_1854,In_988);
and U1651 (N_1651,In_1666,In_285);
nor U1652 (N_1652,In_1217,In_1732);
nand U1653 (N_1653,In_1177,In_320);
nand U1654 (N_1654,In_908,In_1968);
and U1655 (N_1655,In_1814,In_1834);
and U1656 (N_1656,In_868,In_1905);
nor U1657 (N_1657,In_597,In_727);
nand U1658 (N_1658,In_1684,In_1827);
or U1659 (N_1659,In_1908,In_1808);
xor U1660 (N_1660,In_976,In_594);
or U1661 (N_1661,In_1488,In_915);
and U1662 (N_1662,In_1650,In_1420);
nor U1663 (N_1663,In_1705,In_863);
or U1664 (N_1664,In_1376,In_1514);
and U1665 (N_1665,In_696,In_52);
or U1666 (N_1666,In_434,In_206);
xnor U1667 (N_1667,In_241,In_562);
or U1668 (N_1668,In_496,In_977);
nor U1669 (N_1669,In_1703,In_1699);
and U1670 (N_1670,In_528,In_1090);
or U1671 (N_1671,In_751,In_1904);
or U1672 (N_1672,In_205,In_891);
or U1673 (N_1673,In_1423,In_573);
and U1674 (N_1674,In_768,In_1721);
and U1675 (N_1675,In_1358,In_1243);
and U1676 (N_1676,In_629,In_867);
nor U1677 (N_1677,In_300,In_1240);
xnor U1678 (N_1678,In_290,In_881);
nand U1679 (N_1679,In_764,In_1641);
nor U1680 (N_1680,In_562,In_391);
or U1681 (N_1681,In_937,In_1171);
and U1682 (N_1682,In_104,In_519);
and U1683 (N_1683,In_522,In_263);
nand U1684 (N_1684,In_49,In_422);
or U1685 (N_1685,In_1229,In_761);
nor U1686 (N_1686,In_695,In_146);
nor U1687 (N_1687,In_1626,In_842);
xnor U1688 (N_1688,In_1725,In_838);
nor U1689 (N_1689,In_1935,In_1134);
nor U1690 (N_1690,In_856,In_1244);
nand U1691 (N_1691,In_388,In_1861);
and U1692 (N_1692,In_306,In_1969);
and U1693 (N_1693,In_289,In_1739);
or U1694 (N_1694,In_1601,In_80);
or U1695 (N_1695,In_956,In_1000);
and U1696 (N_1696,In_1413,In_1647);
nor U1697 (N_1697,In_349,In_454);
xnor U1698 (N_1698,In_620,In_1056);
or U1699 (N_1699,In_486,In_1670);
nor U1700 (N_1700,In_357,In_1005);
or U1701 (N_1701,In_1358,In_834);
nand U1702 (N_1702,In_1478,In_1563);
nand U1703 (N_1703,In_1057,In_1169);
or U1704 (N_1704,In_1114,In_1705);
xor U1705 (N_1705,In_1752,In_508);
nand U1706 (N_1706,In_849,In_984);
nand U1707 (N_1707,In_1129,In_437);
nand U1708 (N_1708,In_1933,In_171);
and U1709 (N_1709,In_420,In_639);
and U1710 (N_1710,In_158,In_1128);
xnor U1711 (N_1711,In_1748,In_938);
and U1712 (N_1712,In_1659,In_1178);
nor U1713 (N_1713,In_663,In_122);
nand U1714 (N_1714,In_1647,In_1148);
nor U1715 (N_1715,In_286,In_1124);
and U1716 (N_1716,In_173,In_1706);
xnor U1717 (N_1717,In_1877,In_1054);
and U1718 (N_1718,In_200,In_1074);
and U1719 (N_1719,In_235,In_467);
nand U1720 (N_1720,In_1010,In_425);
or U1721 (N_1721,In_1045,In_755);
nand U1722 (N_1722,In_1243,In_1413);
or U1723 (N_1723,In_111,In_964);
or U1724 (N_1724,In_863,In_871);
nand U1725 (N_1725,In_1534,In_1449);
nor U1726 (N_1726,In_1759,In_468);
xor U1727 (N_1727,In_1007,In_482);
xnor U1728 (N_1728,In_612,In_944);
nand U1729 (N_1729,In_283,In_240);
or U1730 (N_1730,In_655,In_1829);
nor U1731 (N_1731,In_62,In_1329);
nand U1732 (N_1732,In_584,In_1823);
nor U1733 (N_1733,In_1164,In_1454);
or U1734 (N_1734,In_1586,In_1364);
or U1735 (N_1735,In_648,In_1766);
or U1736 (N_1736,In_1912,In_181);
or U1737 (N_1737,In_98,In_802);
nand U1738 (N_1738,In_1451,In_631);
or U1739 (N_1739,In_996,In_1605);
nand U1740 (N_1740,In_636,In_73);
nor U1741 (N_1741,In_1801,In_380);
or U1742 (N_1742,In_865,In_22);
nand U1743 (N_1743,In_1639,In_189);
nand U1744 (N_1744,In_1595,In_619);
nand U1745 (N_1745,In_509,In_750);
or U1746 (N_1746,In_1051,In_233);
and U1747 (N_1747,In_1117,In_1152);
xor U1748 (N_1748,In_1422,In_1833);
xnor U1749 (N_1749,In_562,In_117);
and U1750 (N_1750,In_316,In_1943);
and U1751 (N_1751,In_774,In_1974);
and U1752 (N_1752,In_1918,In_1538);
nand U1753 (N_1753,In_1711,In_1762);
nand U1754 (N_1754,In_989,In_368);
xnor U1755 (N_1755,In_821,In_1235);
xnor U1756 (N_1756,In_209,In_1039);
and U1757 (N_1757,In_461,In_471);
and U1758 (N_1758,In_534,In_1653);
nor U1759 (N_1759,In_1471,In_928);
or U1760 (N_1760,In_1087,In_1572);
nor U1761 (N_1761,In_1063,In_1548);
nand U1762 (N_1762,In_1559,In_510);
and U1763 (N_1763,In_1291,In_338);
nor U1764 (N_1764,In_1849,In_1612);
nand U1765 (N_1765,In_310,In_178);
or U1766 (N_1766,In_81,In_1313);
and U1767 (N_1767,In_388,In_415);
nor U1768 (N_1768,In_461,In_1180);
and U1769 (N_1769,In_327,In_1159);
nor U1770 (N_1770,In_1813,In_714);
and U1771 (N_1771,In_649,In_223);
or U1772 (N_1772,In_1667,In_546);
nor U1773 (N_1773,In_880,In_660);
nor U1774 (N_1774,In_1769,In_1454);
nor U1775 (N_1775,In_1310,In_83);
nand U1776 (N_1776,In_1758,In_1537);
nor U1777 (N_1777,In_1692,In_803);
nand U1778 (N_1778,In_1163,In_1627);
nand U1779 (N_1779,In_800,In_1819);
xor U1780 (N_1780,In_834,In_885);
or U1781 (N_1781,In_1760,In_648);
or U1782 (N_1782,In_773,In_90);
nand U1783 (N_1783,In_542,In_1997);
nor U1784 (N_1784,In_335,In_864);
or U1785 (N_1785,In_199,In_1114);
nor U1786 (N_1786,In_503,In_1235);
nand U1787 (N_1787,In_1622,In_99);
xnor U1788 (N_1788,In_1292,In_1099);
nor U1789 (N_1789,In_1142,In_738);
nand U1790 (N_1790,In_983,In_1996);
nor U1791 (N_1791,In_372,In_442);
or U1792 (N_1792,In_1401,In_1549);
nor U1793 (N_1793,In_678,In_957);
xor U1794 (N_1794,In_1233,In_787);
and U1795 (N_1795,In_1155,In_8);
xnor U1796 (N_1796,In_1477,In_239);
xnor U1797 (N_1797,In_91,In_815);
nor U1798 (N_1798,In_1524,In_1140);
nor U1799 (N_1799,In_939,In_300);
nand U1800 (N_1800,In_1933,In_78);
and U1801 (N_1801,In_1276,In_1366);
nand U1802 (N_1802,In_1552,In_727);
or U1803 (N_1803,In_1396,In_362);
nor U1804 (N_1804,In_269,In_286);
nand U1805 (N_1805,In_1289,In_76);
nand U1806 (N_1806,In_299,In_340);
and U1807 (N_1807,In_454,In_578);
and U1808 (N_1808,In_579,In_1550);
nor U1809 (N_1809,In_1245,In_1263);
nand U1810 (N_1810,In_1625,In_360);
or U1811 (N_1811,In_142,In_803);
or U1812 (N_1812,In_510,In_1691);
and U1813 (N_1813,In_1776,In_928);
xnor U1814 (N_1814,In_1460,In_144);
nand U1815 (N_1815,In_1031,In_491);
xnor U1816 (N_1816,In_312,In_1652);
or U1817 (N_1817,In_448,In_702);
nor U1818 (N_1818,In_1738,In_1915);
and U1819 (N_1819,In_993,In_541);
or U1820 (N_1820,In_1396,In_1048);
and U1821 (N_1821,In_1223,In_234);
or U1822 (N_1822,In_595,In_928);
xor U1823 (N_1823,In_245,In_1501);
or U1824 (N_1824,In_575,In_555);
nor U1825 (N_1825,In_711,In_1985);
nand U1826 (N_1826,In_975,In_1928);
nor U1827 (N_1827,In_771,In_1954);
or U1828 (N_1828,In_1721,In_1761);
and U1829 (N_1829,In_72,In_1701);
xor U1830 (N_1830,In_1751,In_878);
or U1831 (N_1831,In_924,In_235);
xor U1832 (N_1832,In_935,In_354);
or U1833 (N_1833,In_899,In_822);
nand U1834 (N_1834,In_1051,In_1865);
nand U1835 (N_1835,In_1697,In_625);
nor U1836 (N_1836,In_1302,In_328);
or U1837 (N_1837,In_1012,In_697);
nand U1838 (N_1838,In_389,In_1735);
xnor U1839 (N_1839,In_1752,In_1910);
or U1840 (N_1840,In_590,In_832);
and U1841 (N_1841,In_653,In_823);
nand U1842 (N_1842,In_1883,In_114);
nor U1843 (N_1843,In_625,In_188);
nor U1844 (N_1844,In_1399,In_1462);
and U1845 (N_1845,In_511,In_278);
nand U1846 (N_1846,In_892,In_366);
nand U1847 (N_1847,In_868,In_858);
xnor U1848 (N_1848,In_1226,In_1154);
nor U1849 (N_1849,In_1038,In_277);
and U1850 (N_1850,In_1328,In_12);
or U1851 (N_1851,In_1791,In_1093);
and U1852 (N_1852,In_1733,In_1334);
and U1853 (N_1853,In_910,In_1775);
nor U1854 (N_1854,In_997,In_81);
nor U1855 (N_1855,In_1130,In_1940);
nand U1856 (N_1856,In_1262,In_705);
or U1857 (N_1857,In_140,In_723);
or U1858 (N_1858,In_710,In_1587);
and U1859 (N_1859,In_1882,In_1089);
xnor U1860 (N_1860,In_1921,In_1947);
and U1861 (N_1861,In_1446,In_916);
nor U1862 (N_1862,In_141,In_418);
and U1863 (N_1863,In_1001,In_1140);
nand U1864 (N_1864,In_1827,In_1699);
or U1865 (N_1865,In_1753,In_1799);
or U1866 (N_1866,In_273,In_1379);
or U1867 (N_1867,In_1263,In_1908);
nand U1868 (N_1868,In_677,In_1449);
or U1869 (N_1869,In_530,In_1239);
nand U1870 (N_1870,In_1978,In_1299);
or U1871 (N_1871,In_127,In_651);
nand U1872 (N_1872,In_1331,In_1205);
nand U1873 (N_1873,In_1113,In_1991);
nand U1874 (N_1874,In_284,In_1770);
nand U1875 (N_1875,In_343,In_851);
nor U1876 (N_1876,In_775,In_1937);
nand U1877 (N_1877,In_317,In_1419);
and U1878 (N_1878,In_212,In_1458);
nor U1879 (N_1879,In_1133,In_1286);
or U1880 (N_1880,In_1531,In_705);
xor U1881 (N_1881,In_896,In_1861);
and U1882 (N_1882,In_408,In_1155);
and U1883 (N_1883,In_1910,In_1894);
nor U1884 (N_1884,In_501,In_243);
and U1885 (N_1885,In_1969,In_276);
nand U1886 (N_1886,In_1136,In_1302);
or U1887 (N_1887,In_647,In_1852);
or U1888 (N_1888,In_1648,In_1308);
or U1889 (N_1889,In_64,In_233);
nand U1890 (N_1890,In_1605,In_1239);
and U1891 (N_1891,In_608,In_578);
and U1892 (N_1892,In_1815,In_201);
xnor U1893 (N_1893,In_1984,In_1548);
nand U1894 (N_1894,In_302,In_496);
nor U1895 (N_1895,In_393,In_267);
nor U1896 (N_1896,In_1693,In_382);
nand U1897 (N_1897,In_1817,In_1743);
and U1898 (N_1898,In_766,In_754);
nor U1899 (N_1899,In_1698,In_527);
nor U1900 (N_1900,In_1529,In_53);
nor U1901 (N_1901,In_1383,In_464);
xor U1902 (N_1902,In_994,In_1635);
or U1903 (N_1903,In_1681,In_691);
or U1904 (N_1904,In_844,In_1123);
and U1905 (N_1905,In_224,In_1341);
xnor U1906 (N_1906,In_552,In_1269);
or U1907 (N_1907,In_466,In_1195);
or U1908 (N_1908,In_1742,In_1479);
nand U1909 (N_1909,In_1345,In_1711);
xor U1910 (N_1910,In_837,In_182);
and U1911 (N_1911,In_312,In_1663);
or U1912 (N_1912,In_710,In_634);
nor U1913 (N_1913,In_1048,In_1785);
or U1914 (N_1914,In_1784,In_1363);
xnor U1915 (N_1915,In_154,In_127);
nand U1916 (N_1916,In_934,In_1997);
nand U1917 (N_1917,In_1546,In_733);
nor U1918 (N_1918,In_1727,In_298);
nor U1919 (N_1919,In_1696,In_108);
xor U1920 (N_1920,In_1372,In_759);
xor U1921 (N_1921,In_13,In_1303);
nand U1922 (N_1922,In_894,In_1175);
nor U1923 (N_1923,In_180,In_937);
nor U1924 (N_1924,In_1647,In_1292);
and U1925 (N_1925,In_1616,In_236);
and U1926 (N_1926,In_1988,In_1908);
nand U1927 (N_1927,In_886,In_1810);
nand U1928 (N_1928,In_1259,In_987);
and U1929 (N_1929,In_120,In_735);
xor U1930 (N_1930,In_395,In_1495);
nor U1931 (N_1931,In_206,In_1188);
xnor U1932 (N_1932,In_1224,In_1588);
nand U1933 (N_1933,In_690,In_657);
xnor U1934 (N_1934,In_1971,In_275);
nand U1935 (N_1935,In_1324,In_523);
nand U1936 (N_1936,In_224,In_1555);
and U1937 (N_1937,In_1315,In_980);
nand U1938 (N_1938,In_1048,In_524);
or U1939 (N_1939,In_398,In_1037);
nand U1940 (N_1940,In_1976,In_110);
nor U1941 (N_1941,In_1539,In_900);
nor U1942 (N_1942,In_1872,In_1807);
nand U1943 (N_1943,In_276,In_1451);
nor U1944 (N_1944,In_1307,In_1229);
nand U1945 (N_1945,In_1965,In_1488);
xor U1946 (N_1946,In_1040,In_1418);
or U1947 (N_1947,In_1452,In_1846);
and U1948 (N_1948,In_917,In_31);
and U1949 (N_1949,In_1125,In_1520);
nand U1950 (N_1950,In_1614,In_89);
xnor U1951 (N_1951,In_893,In_1412);
or U1952 (N_1952,In_1117,In_184);
and U1953 (N_1953,In_994,In_1582);
and U1954 (N_1954,In_1129,In_243);
and U1955 (N_1955,In_1403,In_1913);
nor U1956 (N_1956,In_209,In_1557);
and U1957 (N_1957,In_83,In_284);
nor U1958 (N_1958,In_1623,In_531);
nor U1959 (N_1959,In_1134,In_333);
nand U1960 (N_1960,In_1975,In_1685);
or U1961 (N_1961,In_1986,In_512);
nor U1962 (N_1962,In_534,In_797);
nor U1963 (N_1963,In_968,In_1121);
and U1964 (N_1964,In_1065,In_777);
and U1965 (N_1965,In_1108,In_340);
and U1966 (N_1966,In_217,In_1114);
nand U1967 (N_1967,In_1593,In_775);
nor U1968 (N_1968,In_406,In_1812);
nor U1969 (N_1969,In_1073,In_582);
nor U1970 (N_1970,In_1531,In_118);
nor U1971 (N_1971,In_973,In_822);
nand U1972 (N_1972,In_715,In_705);
or U1973 (N_1973,In_1530,In_39);
nor U1974 (N_1974,In_1494,In_1533);
or U1975 (N_1975,In_12,In_1816);
xor U1976 (N_1976,In_530,In_1037);
nor U1977 (N_1977,In_1076,In_985);
and U1978 (N_1978,In_704,In_1856);
nor U1979 (N_1979,In_1230,In_823);
nor U1980 (N_1980,In_40,In_786);
nor U1981 (N_1981,In_154,In_497);
nor U1982 (N_1982,In_924,In_1077);
and U1983 (N_1983,In_272,In_1708);
nand U1984 (N_1984,In_349,In_1702);
xnor U1985 (N_1985,In_21,In_1019);
or U1986 (N_1986,In_577,In_940);
nor U1987 (N_1987,In_797,In_1468);
xor U1988 (N_1988,In_1421,In_1692);
nand U1989 (N_1989,In_358,In_1259);
nor U1990 (N_1990,In_586,In_1715);
and U1991 (N_1991,In_974,In_1551);
nor U1992 (N_1992,In_946,In_265);
or U1993 (N_1993,In_1676,In_1613);
nor U1994 (N_1994,In_836,In_453);
nand U1995 (N_1995,In_373,In_393);
and U1996 (N_1996,In_1050,In_1107);
or U1997 (N_1997,In_1707,In_1920);
or U1998 (N_1998,In_252,In_985);
nor U1999 (N_1999,In_1028,In_1904);
and U2000 (N_2000,In_252,In_1562);
nand U2001 (N_2001,In_283,In_915);
or U2002 (N_2002,In_1064,In_1501);
nand U2003 (N_2003,In_1452,In_655);
or U2004 (N_2004,In_1458,In_223);
nor U2005 (N_2005,In_1552,In_902);
nand U2006 (N_2006,In_1740,In_1399);
and U2007 (N_2007,In_1924,In_1805);
and U2008 (N_2008,In_1851,In_1094);
xor U2009 (N_2009,In_1897,In_60);
nand U2010 (N_2010,In_1007,In_1550);
and U2011 (N_2011,In_1853,In_1100);
nor U2012 (N_2012,In_1140,In_893);
or U2013 (N_2013,In_129,In_1571);
nand U2014 (N_2014,In_919,In_215);
or U2015 (N_2015,In_837,In_1163);
nor U2016 (N_2016,In_1983,In_1058);
nor U2017 (N_2017,In_1861,In_1039);
nor U2018 (N_2018,In_1273,In_1214);
and U2019 (N_2019,In_98,In_1703);
nor U2020 (N_2020,In_1981,In_229);
or U2021 (N_2021,In_1740,In_759);
or U2022 (N_2022,In_688,In_1241);
nor U2023 (N_2023,In_1681,In_596);
nand U2024 (N_2024,In_1885,In_356);
or U2025 (N_2025,In_1971,In_907);
and U2026 (N_2026,In_506,In_1479);
nor U2027 (N_2027,In_382,In_212);
nand U2028 (N_2028,In_479,In_954);
nand U2029 (N_2029,In_1428,In_740);
nand U2030 (N_2030,In_837,In_1302);
and U2031 (N_2031,In_477,In_849);
nor U2032 (N_2032,In_404,In_988);
nor U2033 (N_2033,In_921,In_1916);
nand U2034 (N_2034,In_453,In_697);
and U2035 (N_2035,In_1631,In_1027);
and U2036 (N_2036,In_941,In_219);
xor U2037 (N_2037,In_392,In_1709);
or U2038 (N_2038,In_1017,In_524);
nor U2039 (N_2039,In_887,In_1914);
or U2040 (N_2040,In_1849,In_303);
or U2041 (N_2041,In_25,In_1018);
or U2042 (N_2042,In_34,In_1454);
xnor U2043 (N_2043,In_1169,In_348);
and U2044 (N_2044,In_346,In_214);
nand U2045 (N_2045,In_1885,In_66);
and U2046 (N_2046,In_1167,In_888);
and U2047 (N_2047,In_863,In_1336);
nand U2048 (N_2048,In_780,In_1105);
or U2049 (N_2049,In_102,In_535);
and U2050 (N_2050,In_1728,In_299);
nand U2051 (N_2051,In_545,In_1540);
nand U2052 (N_2052,In_887,In_641);
nand U2053 (N_2053,In_40,In_1925);
nand U2054 (N_2054,In_1001,In_248);
nand U2055 (N_2055,In_1058,In_437);
nand U2056 (N_2056,In_1259,In_1819);
or U2057 (N_2057,In_843,In_619);
and U2058 (N_2058,In_1901,In_339);
and U2059 (N_2059,In_1515,In_1355);
or U2060 (N_2060,In_1309,In_380);
and U2061 (N_2061,In_1713,In_1902);
nor U2062 (N_2062,In_1274,In_1584);
and U2063 (N_2063,In_1994,In_1450);
and U2064 (N_2064,In_945,In_1621);
and U2065 (N_2065,In_189,In_1268);
nor U2066 (N_2066,In_833,In_354);
nor U2067 (N_2067,In_605,In_1893);
nand U2068 (N_2068,In_742,In_193);
nand U2069 (N_2069,In_1516,In_100);
nand U2070 (N_2070,In_1987,In_1865);
or U2071 (N_2071,In_1433,In_32);
or U2072 (N_2072,In_740,In_659);
nor U2073 (N_2073,In_1793,In_915);
xnor U2074 (N_2074,In_126,In_1474);
and U2075 (N_2075,In_640,In_1317);
and U2076 (N_2076,In_228,In_1966);
nor U2077 (N_2077,In_158,In_1831);
xnor U2078 (N_2078,In_1195,In_722);
and U2079 (N_2079,In_388,In_313);
and U2080 (N_2080,In_619,In_866);
xnor U2081 (N_2081,In_890,In_1839);
nor U2082 (N_2082,In_1900,In_935);
xnor U2083 (N_2083,In_55,In_1552);
nor U2084 (N_2084,In_1384,In_1060);
and U2085 (N_2085,In_594,In_557);
nand U2086 (N_2086,In_1592,In_326);
or U2087 (N_2087,In_97,In_919);
xor U2088 (N_2088,In_701,In_927);
and U2089 (N_2089,In_748,In_364);
or U2090 (N_2090,In_1600,In_1764);
or U2091 (N_2091,In_458,In_230);
or U2092 (N_2092,In_844,In_306);
and U2093 (N_2093,In_808,In_1176);
and U2094 (N_2094,In_1381,In_857);
nand U2095 (N_2095,In_1926,In_1019);
nor U2096 (N_2096,In_1295,In_1167);
nand U2097 (N_2097,In_101,In_408);
and U2098 (N_2098,In_1321,In_1649);
nor U2099 (N_2099,In_1469,In_1442);
and U2100 (N_2100,In_522,In_225);
nand U2101 (N_2101,In_1443,In_1915);
and U2102 (N_2102,In_842,In_42);
nor U2103 (N_2103,In_847,In_918);
or U2104 (N_2104,In_1506,In_1261);
and U2105 (N_2105,In_658,In_1971);
and U2106 (N_2106,In_1625,In_1529);
and U2107 (N_2107,In_1130,In_41);
or U2108 (N_2108,In_713,In_1395);
nand U2109 (N_2109,In_1501,In_1338);
and U2110 (N_2110,In_608,In_773);
and U2111 (N_2111,In_747,In_187);
or U2112 (N_2112,In_1190,In_1086);
or U2113 (N_2113,In_987,In_19);
xor U2114 (N_2114,In_202,In_530);
nand U2115 (N_2115,In_217,In_219);
and U2116 (N_2116,In_590,In_192);
nand U2117 (N_2117,In_360,In_25);
or U2118 (N_2118,In_771,In_131);
nand U2119 (N_2119,In_1715,In_1290);
and U2120 (N_2120,In_1420,In_1641);
or U2121 (N_2121,In_296,In_758);
or U2122 (N_2122,In_987,In_272);
nand U2123 (N_2123,In_876,In_1060);
nor U2124 (N_2124,In_4,In_1230);
nand U2125 (N_2125,In_843,In_669);
or U2126 (N_2126,In_1737,In_1708);
nand U2127 (N_2127,In_666,In_109);
nand U2128 (N_2128,In_1016,In_344);
and U2129 (N_2129,In_519,In_1943);
or U2130 (N_2130,In_1786,In_1667);
xnor U2131 (N_2131,In_460,In_1784);
or U2132 (N_2132,In_1125,In_892);
nand U2133 (N_2133,In_277,In_1561);
or U2134 (N_2134,In_1058,In_555);
or U2135 (N_2135,In_442,In_1219);
nand U2136 (N_2136,In_278,In_1029);
nand U2137 (N_2137,In_1600,In_204);
nor U2138 (N_2138,In_454,In_372);
nor U2139 (N_2139,In_632,In_1400);
and U2140 (N_2140,In_1065,In_1738);
nand U2141 (N_2141,In_452,In_1553);
xnor U2142 (N_2142,In_542,In_1522);
nor U2143 (N_2143,In_1632,In_918);
nor U2144 (N_2144,In_1780,In_1737);
and U2145 (N_2145,In_844,In_545);
and U2146 (N_2146,In_430,In_591);
nand U2147 (N_2147,In_655,In_1380);
nor U2148 (N_2148,In_1937,In_750);
nand U2149 (N_2149,In_1141,In_1502);
nand U2150 (N_2150,In_1381,In_1957);
or U2151 (N_2151,In_1961,In_293);
xnor U2152 (N_2152,In_1829,In_495);
nor U2153 (N_2153,In_1124,In_1127);
nand U2154 (N_2154,In_496,In_1912);
xnor U2155 (N_2155,In_1628,In_1875);
or U2156 (N_2156,In_755,In_189);
and U2157 (N_2157,In_559,In_657);
nor U2158 (N_2158,In_1545,In_942);
or U2159 (N_2159,In_755,In_1665);
or U2160 (N_2160,In_1939,In_1512);
nand U2161 (N_2161,In_150,In_386);
nand U2162 (N_2162,In_363,In_72);
nand U2163 (N_2163,In_1232,In_1024);
and U2164 (N_2164,In_1794,In_287);
and U2165 (N_2165,In_539,In_1476);
nand U2166 (N_2166,In_1568,In_1779);
nor U2167 (N_2167,In_1554,In_207);
or U2168 (N_2168,In_1572,In_1937);
or U2169 (N_2169,In_540,In_1150);
nand U2170 (N_2170,In_1796,In_1236);
nand U2171 (N_2171,In_1881,In_756);
nand U2172 (N_2172,In_1206,In_600);
or U2173 (N_2173,In_1493,In_1687);
or U2174 (N_2174,In_233,In_667);
nor U2175 (N_2175,In_493,In_462);
and U2176 (N_2176,In_341,In_543);
xor U2177 (N_2177,In_26,In_1342);
nor U2178 (N_2178,In_617,In_328);
or U2179 (N_2179,In_1324,In_149);
nand U2180 (N_2180,In_1152,In_1351);
nand U2181 (N_2181,In_1798,In_477);
or U2182 (N_2182,In_433,In_1712);
and U2183 (N_2183,In_879,In_58);
nor U2184 (N_2184,In_735,In_926);
and U2185 (N_2185,In_854,In_701);
and U2186 (N_2186,In_749,In_61);
and U2187 (N_2187,In_756,In_1821);
or U2188 (N_2188,In_1611,In_237);
xnor U2189 (N_2189,In_1338,In_511);
and U2190 (N_2190,In_1657,In_993);
nor U2191 (N_2191,In_1520,In_242);
or U2192 (N_2192,In_563,In_1938);
or U2193 (N_2193,In_1340,In_1409);
nand U2194 (N_2194,In_1799,In_1835);
and U2195 (N_2195,In_1547,In_1197);
nand U2196 (N_2196,In_1567,In_862);
nor U2197 (N_2197,In_1241,In_942);
xor U2198 (N_2198,In_1270,In_989);
nand U2199 (N_2199,In_1913,In_1329);
and U2200 (N_2200,In_1429,In_386);
xor U2201 (N_2201,In_969,In_1541);
nand U2202 (N_2202,In_1867,In_873);
nand U2203 (N_2203,In_498,In_432);
xor U2204 (N_2204,In_105,In_447);
nand U2205 (N_2205,In_1127,In_1398);
xnor U2206 (N_2206,In_1821,In_1909);
nor U2207 (N_2207,In_532,In_1269);
nand U2208 (N_2208,In_1620,In_843);
and U2209 (N_2209,In_1624,In_1772);
nor U2210 (N_2210,In_329,In_187);
and U2211 (N_2211,In_998,In_1190);
nor U2212 (N_2212,In_1219,In_436);
nand U2213 (N_2213,In_1344,In_1043);
or U2214 (N_2214,In_391,In_1858);
xor U2215 (N_2215,In_557,In_1507);
nand U2216 (N_2216,In_1093,In_634);
nand U2217 (N_2217,In_597,In_1085);
nor U2218 (N_2218,In_1571,In_1436);
or U2219 (N_2219,In_1996,In_1044);
and U2220 (N_2220,In_631,In_550);
nor U2221 (N_2221,In_1089,In_315);
or U2222 (N_2222,In_1303,In_592);
xnor U2223 (N_2223,In_1957,In_1816);
or U2224 (N_2224,In_1861,In_1121);
nor U2225 (N_2225,In_584,In_986);
nor U2226 (N_2226,In_630,In_494);
and U2227 (N_2227,In_13,In_63);
or U2228 (N_2228,In_1500,In_125);
nand U2229 (N_2229,In_1220,In_1304);
nor U2230 (N_2230,In_1792,In_1825);
nand U2231 (N_2231,In_466,In_13);
nand U2232 (N_2232,In_1435,In_874);
and U2233 (N_2233,In_1228,In_1957);
and U2234 (N_2234,In_1351,In_1218);
and U2235 (N_2235,In_135,In_1736);
nand U2236 (N_2236,In_1020,In_1704);
nand U2237 (N_2237,In_620,In_1619);
and U2238 (N_2238,In_1049,In_81);
nand U2239 (N_2239,In_167,In_292);
and U2240 (N_2240,In_991,In_1029);
and U2241 (N_2241,In_249,In_1206);
or U2242 (N_2242,In_1751,In_56);
nor U2243 (N_2243,In_802,In_888);
or U2244 (N_2244,In_765,In_1075);
and U2245 (N_2245,In_1761,In_757);
nor U2246 (N_2246,In_826,In_908);
or U2247 (N_2247,In_1157,In_481);
or U2248 (N_2248,In_157,In_1007);
nand U2249 (N_2249,In_1709,In_817);
or U2250 (N_2250,In_1312,In_115);
nand U2251 (N_2251,In_1202,In_1405);
xor U2252 (N_2252,In_1016,In_1105);
nor U2253 (N_2253,In_113,In_507);
nand U2254 (N_2254,In_1387,In_897);
nand U2255 (N_2255,In_1571,In_383);
and U2256 (N_2256,In_6,In_1976);
or U2257 (N_2257,In_842,In_1991);
and U2258 (N_2258,In_1949,In_1705);
nor U2259 (N_2259,In_758,In_1702);
nor U2260 (N_2260,In_402,In_612);
nand U2261 (N_2261,In_1245,In_68);
or U2262 (N_2262,In_253,In_1847);
or U2263 (N_2263,In_235,In_670);
or U2264 (N_2264,In_530,In_1602);
and U2265 (N_2265,In_158,In_371);
and U2266 (N_2266,In_921,In_1356);
nor U2267 (N_2267,In_1974,In_1419);
nand U2268 (N_2268,In_1607,In_1120);
or U2269 (N_2269,In_495,In_869);
nor U2270 (N_2270,In_944,In_815);
nand U2271 (N_2271,In_257,In_1406);
and U2272 (N_2272,In_1238,In_124);
nor U2273 (N_2273,In_1049,In_1874);
and U2274 (N_2274,In_728,In_752);
xnor U2275 (N_2275,In_1337,In_586);
xnor U2276 (N_2276,In_519,In_1852);
or U2277 (N_2277,In_1444,In_1575);
nor U2278 (N_2278,In_1420,In_1700);
nor U2279 (N_2279,In_1472,In_1435);
or U2280 (N_2280,In_1127,In_764);
or U2281 (N_2281,In_1758,In_1426);
nand U2282 (N_2282,In_195,In_1439);
nand U2283 (N_2283,In_1978,In_1603);
nor U2284 (N_2284,In_695,In_1240);
nand U2285 (N_2285,In_1250,In_889);
or U2286 (N_2286,In_1087,In_787);
or U2287 (N_2287,In_708,In_1380);
nor U2288 (N_2288,In_1626,In_818);
nand U2289 (N_2289,In_1122,In_1295);
nor U2290 (N_2290,In_1875,In_1043);
nand U2291 (N_2291,In_1028,In_68);
or U2292 (N_2292,In_1120,In_1305);
or U2293 (N_2293,In_428,In_766);
nand U2294 (N_2294,In_530,In_806);
and U2295 (N_2295,In_888,In_1517);
and U2296 (N_2296,In_1371,In_1213);
nor U2297 (N_2297,In_192,In_965);
nand U2298 (N_2298,In_1682,In_1746);
or U2299 (N_2299,In_1397,In_35);
or U2300 (N_2300,In_1778,In_200);
or U2301 (N_2301,In_1781,In_1724);
or U2302 (N_2302,In_1597,In_1840);
or U2303 (N_2303,In_639,In_955);
and U2304 (N_2304,In_357,In_1380);
and U2305 (N_2305,In_1490,In_1730);
nand U2306 (N_2306,In_563,In_1141);
and U2307 (N_2307,In_443,In_214);
nand U2308 (N_2308,In_289,In_1724);
nor U2309 (N_2309,In_1367,In_1801);
nor U2310 (N_2310,In_500,In_1988);
nor U2311 (N_2311,In_435,In_1733);
nand U2312 (N_2312,In_487,In_1121);
or U2313 (N_2313,In_1868,In_1524);
xor U2314 (N_2314,In_132,In_736);
or U2315 (N_2315,In_1091,In_1370);
nor U2316 (N_2316,In_577,In_827);
or U2317 (N_2317,In_1132,In_543);
xor U2318 (N_2318,In_1413,In_1480);
nor U2319 (N_2319,In_1332,In_402);
or U2320 (N_2320,In_1514,In_110);
or U2321 (N_2321,In_1458,In_1744);
nor U2322 (N_2322,In_890,In_1524);
nand U2323 (N_2323,In_1805,In_1834);
xor U2324 (N_2324,In_1818,In_947);
nand U2325 (N_2325,In_708,In_386);
nor U2326 (N_2326,In_31,In_1015);
or U2327 (N_2327,In_1349,In_658);
and U2328 (N_2328,In_1201,In_771);
or U2329 (N_2329,In_1284,In_1399);
nor U2330 (N_2330,In_1097,In_940);
nor U2331 (N_2331,In_1388,In_372);
nor U2332 (N_2332,In_1948,In_874);
and U2333 (N_2333,In_18,In_800);
or U2334 (N_2334,In_851,In_1000);
and U2335 (N_2335,In_304,In_681);
nand U2336 (N_2336,In_766,In_179);
nor U2337 (N_2337,In_1488,In_547);
nor U2338 (N_2338,In_1876,In_381);
and U2339 (N_2339,In_1832,In_1391);
nor U2340 (N_2340,In_457,In_1314);
nand U2341 (N_2341,In_1195,In_1155);
nor U2342 (N_2342,In_1273,In_1792);
nand U2343 (N_2343,In_1140,In_792);
nand U2344 (N_2344,In_1201,In_761);
nor U2345 (N_2345,In_1230,In_511);
xnor U2346 (N_2346,In_613,In_457);
nor U2347 (N_2347,In_439,In_1310);
and U2348 (N_2348,In_1608,In_681);
and U2349 (N_2349,In_39,In_1008);
and U2350 (N_2350,In_1833,In_1125);
nand U2351 (N_2351,In_25,In_38);
nor U2352 (N_2352,In_1744,In_1264);
or U2353 (N_2353,In_1857,In_111);
nor U2354 (N_2354,In_376,In_351);
nor U2355 (N_2355,In_1224,In_1088);
nor U2356 (N_2356,In_403,In_467);
and U2357 (N_2357,In_954,In_486);
nor U2358 (N_2358,In_348,In_1384);
nor U2359 (N_2359,In_1477,In_1308);
or U2360 (N_2360,In_1506,In_801);
and U2361 (N_2361,In_973,In_595);
xor U2362 (N_2362,In_1069,In_1756);
nand U2363 (N_2363,In_1032,In_460);
or U2364 (N_2364,In_26,In_583);
nand U2365 (N_2365,In_1765,In_223);
and U2366 (N_2366,In_787,In_1453);
or U2367 (N_2367,In_715,In_1918);
and U2368 (N_2368,In_1687,In_982);
and U2369 (N_2369,In_1019,In_257);
or U2370 (N_2370,In_754,In_8);
nor U2371 (N_2371,In_345,In_364);
or U2372 (N_2372,In_432,In_1448);
or U2373 (N_2373,In_527,In_1078);
nand U2374 (N_2374,In_1723,In_1889);
or U2375 (N_2375,In_182,In_1156);
and U2376 (N_2376,In_1531,In_1912);
nand U2377 (N_2377,In_1649,In_575);
or U2378 (N_2378,In_1844,In_1791);
or U2379 (N_2379,In_418,In_1449);
or U2380 (N_2380,In_86,In_1218);
nor U2381 (N_2381,In_629,In_968);
and U2382 (N_2382,In_317,In_958);
or U2383 (N_2383,In_238,In_1045);
and U2384 (N_2384,In_1025,In_859);
xnor U2385 (N_2385,In_1813,In_995);
and U2386 (N_2386,In_1153,In_1882);
or U2387 (N_2387,In_1608,In_220);
xor U2388 (N_2388,In_1711,In_1000);
nor U2389 (N_2389,In_1613,In_1825);
nor U2390 (N_2390,In_884,In_1679);
and U2391 (N_2391,In_1915,In_479);
or U2392 (N_2392,In_1242,In_569);
and U2393 (N_2393,In_109,In_125);
nand U2394 (N_2394,In_216,In_261);
xnor U2395 (N_2395,In_419,In_179);
nand U2396 (N_2396,In_831,In_1460);
nand U2397 (N_2397,In_1715,In_856);
nand U2398 (N_2398,In_1867,In_1075);
or U2399 (N_2399,In_875,In_1682);
nor U2400 (N_2400,In_1691,In_1774);
or U2401 (N_2401,In_177,In_1606);
nand U2402 (N_2402,In_1812,In_1710);
and U2403 (N_2403,In_1033,In_776);
or U2404 (N_2404,In_500,In_945);
and U2405 (N_2405,In_1619,In_1007);
xnor U2406 (N_2406,In_1991,In_226);
nand U2407 (N_2407,In_1791,In_1414);
nor U2408 (N_2408,In_983,In_1208);
xor U2409 (N_2409,In_1623,In_1871);
xnor U2410 (N_2410,In_953,In_1014);
xor U2411 (N_2411,In_562,In_773);
nor U2412 (N_2412,In_1871,In_527);
or U2413 (N_2413,In_430,In_1660);
and U2414 (N_2414,In_1453,In_1344);
nor U2415 (N_2415,In_1307,In_534);
nor U2416 (N_2416,In_616,In_933);
xor U2417 (N_2417,In_119,In_560);
nor U2418 (N_2418,In_1353,In_544);
nand U2419 (N_2419,In_183,In_312);
nor U2420 (N_2420,In_261,In_279);
and U2421 (N_2421,In_1884,In_1109);
nand U2422 (N_2422,In_215,In_855);
nor U2423 (N_2423,In_413,In_1293);
nand U2424 (N_2424,In_26,In_516);
nand U2425 (N_2425,In_348,In_1672);
nor U2426 (N_2426,In_1201,In_969);
nand U2427 (N_2427,In_960,In_1837);
and U2428 (N_2428,In_180,In_1131);
nor U2429 (N_2429,In_137,In_1081);
nand U2430 (N_2430,In_1345,In_625);
and U2431 (N_2431,In_1691,In_472);
nor U2432 (N_2432,In_611,In_38);
and U2433 (N_2433,In_817,In_1285);
and U2434 (N_2434,In_889,In_1849);
nor U2435 (N_2435,In_1187,In_318);
nand U2436 (N_2436,In_1422,In_1554);
nor U2437 (N_2437,In_1279,In_1514);
xor U2438 (N_2438,In_1626,In_1209);
nand U2439 (N_2439,In_528,In_1430);
nor U2440 (N_2440,In_111,In_1415);
nand U2441 (N_2441,In_369,In_39);
or U2442 (N_2442,In_177,In_1075);
nor U2443 (N_2443,In_1221,In_787);
or U2444 (N_2444,In_791,In_1130);
or U2445 (N_2445,In_1517,In_1775);
xor U2446 (N_2446,In_90,In_1848);
and U2447 (N_2447,In_1142,In_1792);
and U2448 (N_2448,In_1256,In_1716);
nand U2449 (N_2449,In_1123,In_199);
xor U2450 (N_2450,In_798,In_325);
or U2451 (N_2451,In_865,In_969);
and U2452 (N_2452,In_1407,In_1219);
and U2453 (N_2453,In_801,In_1287);
nor U2454 (N_2454,In_1955,In_478);
nor U2455 (N_2455,In_1012,In_1187);
or U2456 (N_2456,In_1497,In_815);
xnor U2457 (N_2457,In_14,In_158);
or U2458 (N_2458,In_8,In_486);
or U2459 (N_2459,In_1882,In_1754);
and U2460 (N_2460,In_1389,In_1728);
nor U2461 (N_2461,In_1997,In_195);
or U2462 (N_2462,In_1960,In_82);
xnor U2463 (N_2463,In_1086,In_346);
nor U2464 (N_2464,In_1559,In_645);
nand U2465 (N_2465,In_707,In_1742);
and U2466 (N_2466,In_1318,In_1581);
and U2467 (N_2467,In_1840,In_1780);
nand U2468 (N_2468,In_1455,In_1819);
nor U2469 (N_2469,In_1864,In_654);
nand U2470 (N_2470,In_1593,In_219);
nor U2471 (N_2471,In_1407,In_167);
xor U2472 (N_2472,In_1212,In_1873);
or U2473 (N_2473,In_1518,In_1370);
or U2474 (N_2474,In_28,In_796);
nand U2475 (N_2475,In_1369,In_1131);
or U2476 (N_2476,In_188,In_1912);
or U2477 (N_2477,In_1420,In_1246);
nand U2478 (N_2478,In_1339,In_807);
nor U2479 (N_2479,In_1119,In_1839);
nor U2480 (N_2480,In_1109,In_220);
and U2481 (N_2481,In_126,In_538);
nor U2482 (N_2482,In_1759,In_832);
and U2483 (N_2483,In_848,In_10);
nand U2484 (N_2484,In_1053,In_636);
or U2485 (N_2485,In_262,In_226);
and U2486 (N_2486,In_26,In_340);
nor U2487 (N_2487,In_818,In_1394);
nor U2488 (N_2488,In_417,In_1876);
nor U2489 (N_2489,In_882,In_1654);
and U2490 (N_2490,In_244,In_1204);
or U2491 (N_2491,In_930,In_466);
nor U2492 (N_2492,In_427,In_1669);
or U2493 (N_2493,In_868,In_1515);
xor U2494 (N_2494,In_987,In_1078);
nor U2495 (N_2495,In_997,In_1175);
or U2496 (N_2496,In_187,In_1389);
nand U2497 (N_2497,In_1265,In_1276);
or U2498 (N_2498,In_214,In_646);
nand U2499 (N_2499,In_689,In_851);
xor U2500 (N_2500,In_604,In_750);
nand U2501 (N_2501,In_1053,In_1133);
nand U2502 (N_2502,In_1394,In_444);
nor U2503 (N_2503,In_1115,In_776);
and U2504 (N_2504,In_1149,In_719);
and U2505 (N_2505,In_218,In_768);
nor U2506 (N_2506,In_1670,In_981);
nor U2507 (N_2507,In_739,In_1327);
and U2508 (N_2508,In_496,In_1560);
xor U2509 (N_2509,In_1416,In_1799);
and U2510 (N_2510,In_1502,In_27);
or U2511 (N_2511,In_1198,In_1091);
or U2512 (N_2512,In_1057,In_510);
nor U2513 (N_2513,In_1452,In_987);
nand U2514 (N_2514,In_604,In_617);
xor U2515 (N_2515,In_838,In_1957);
or U2516 (N_2516,In_308,In_472);
nand U2517 (N_2517,In_1859,In_1448);
nor U2518 (N_2518,In_125,In_1901);
and U2519 (N_2519,In_328,In_18);
or U2520 (N_2520,In_1172,In_1765);
and U2521 (N_2521,In_1336,In_690);
and U2522 (N_2522,In_1408,In_1263);
nor U2523 (N_2523,In_969,In_1146);
nand U2524 (N_2524,In_389,In_245);
nand U2525 (N_2525,In_1423,In_317);
or U2526 (N_2526,In_958,In_540);
nor U2527 (N_2527,In_1289,In_1808);
nand U2528 (N_2528,In_673,In_1205);
nor U2529 (N_2529,In_0,In_949);
nor U2530 (N_2530,In_934,In_1242);
or U2531 (N_2531,In_1384,In_1205);
nor U2532 (N_2532,In_1527,In_1568);
and U2533 (N_2533,In_727,In_1638);
and U2534 (N_2534,In_1433,In_1638);
nand U2535 (N_2535,In_1634,In_552);
xnor U2536 (N_2536,In_737,In_105);
nor U2537 (N_2537,In_804,In_1083);
nor U2538 (N_2538,In_76,In_632);
xnor U2539 (N_2539,In_997,In_1325);
or U2540 (N_2540,In_1572,In_475);
or U2541 (N_2541,In_654,In_411);
nor U2542 (N_2542,In_1780,In_1182);
or U2543 (N_2543,In_1704,In_1933);
nor U2544 (N_2544,In_1367,In_1634);
nor U2545 (N_2545,In_763,In_445);
nand U2546 (N_2546,In_565,In_1051);
nor U2547 (N_2547,In_927,In_1239);
or U2548 (N_2548,In_111,In_999);
and U2549 (N_2549,In_1991,In_228);
and U2550 (N_2550,In_1252,In_781);
nor U2551 (N_2551,In_1663,In_541);
or U2552 (N_2552,In_35,In_1731);
nand U2553 (N_2553,In_290,In_961);
nor U2554 (N_2554,In_807,In_55);
nor U2555 (N_2555,In_1550,In_1895);
or U2556 (N_2556,In_1778,In_1942);
xnor U2557 (N_2557,In_456,In_1271);
xnor U2558 (N_2558,In_1438,In_1460);
nor U2559 (N_2559,In_1402,In_462);
or U2560 (N_2560,In_1728,In_1492);
or U2561 (N_2561,In_653,In_1210);
or U2562 (N_2562,In_1378,In_1730);
or U2563 (N_2563,In_613,In_1649);
nor U2564 (N_2564,In_899,In_1674);
or U2565 (N_2565,In_315,In_116);
nor U2566 (N_2566,In_365,In_1528);
and U2567 (N_2567,In_641,In_715);
nand U2568 (N_2568,In_1591,In_1605);
and U2569 (N_2569,In_1157,In_330);
nor U2570 (N_2570,In_1388,In_774);
nor U2571 (N_2571,In_857,In_1287);
nor U2572 (N_2572,In_919,In_441);
or U2573 (N_2573,In_1651,In_1925);
and U2574 (N_2574,In_1328,In_1158);
nor U2575 (N_2575,In_1833,In_1755);
or U2576 (N_2576,In_1199,In_540);
xor U2577 (N_2577,In_781,In_1065);
xor U2578 (N_2578,In_1363,In_1757);
or U2579 (N_2579,In_116,In_347);
nand U2580 (N_2580,In_1240,In_855);
nand U2581 (N_2581,In_1995,In_1684);
nor U2582 (N_2582,In_559,In_1518);
or U2583 (N_2583,In_437,In_1095);
nand U2584 (N_2584,In_1799,In_1527);
and U2585 (N_2585,In_621,In_622);
or U2586 (N_2586,In_1437,In_1345);
xnor U2587 (N_2587,In_62,In_336);
nand U2588 (N_2588,In_1833,In_1807);
nor U2589 (N_2589,In_1318,In_170);
nor U2590 (N_2590,In_165,In_337);
and U2591 (N_2591,In_24,In_1232);
and U2592 (N_2592,In_1488,In_404);
and U2593 (N_2593,In_1242,In_1453);
nor U2594 (N_2594,In_808,In_611);
or U2595 (N_2595,In_1757,In_445);
and U2596 (N_2596,In_175,In_938);
nand U2597 (N_2597,In_432,In_1683);
nor U2598 (N_2598,In_96,In_26);
xor U2599 (N_2599,In_33,In_803);
nand U2600 (N_2600,In_615,In_78);
and U2601 (N_2601,In_1033,In_1834);
nand U2602 (N_2602,In_1207,In_1061);
xor U2603 (N_2603,In_955,In_171);
nor U2604 (N_2604,In_853,In_1653);
nor U2605 (N_2605,In_47,In_233);
and U2606 (N_2606,In_1726,In_851);
or U2607 (N_2607,In_1531,In_1476);
nor U2608 (N_2608,In_1218,In_728);
and U2609 (N_2609,In_1107,In_79);
nand U2610 (N_2610,In_929,In_1292);
and U2611 (N_2611,In_182,In_720);
nor U2612 (N_2612,In_49,In_1424);
nand U2613 (N_2613,In_944,In_949);
nand U2614 (N_2614,In_1322,In_691);
nand U2615 (N_2615,In_113,In_756);
xnor U2616 (N_2616,In_143,In_937);
or U2617 (N_2617,In_1444,In_606);
and U2618 (N_2618,In_1129,In_1702);
or U2619 (N_2619,In_761,In_664);
nand U2620 (N_2620,In_687,In_532);
nor U2621 (N_2621,In_1175,In_1004);
or U2622 (N_2622,In_907,In_1763);
or U2623 (N_2623,In_1771,In_970);
and U2624 (N_2624,In_203,In_788);
xor U2625 (N_2625,In_1268,In_1160);
nor U2626 (N_2626,In_311,In_1742);
or U2627 (N_2627,In_708,In_728);
nor U2628 (N_2628,In_1377,In_916);
nand U2629 (N_2629,In_1888,In_323);
or U2630 (N_2630,In_1287,In_818);
nand U2631 (N_2631,In_1344,In_736);
and U2632 (N_2632,In_695,In_300);
xor U2633 (N_2633,In_226,In_1828);
nand U2634 (N_2634,In_551,In_1090);
nor U2635 (N_2635,In_1754,In_1909);
nand U2636 (N_2636,In_1411,In_1824);
nor U2637 (N_2637,In_1111,In_434);
nor U2638 (N_2638,In_1409,In_1100);
and U2639 (N_2639,In_1115,In_613);
nand U2640 (N_2640,In_1554,In_1829);
nor U2641 (N_2641,In_521,In_139);
nor U2642 (N_2642,In_1683,In_1467);
nor U2643 (N_2643,In_1398,In_62);
nand U2644 (N_2644,In_1232,In_295);
nor U2645 (N_2645,In_38,In_1757);
nand U2646 (N_2646,In_1885,In_1388);
xor U2647 (N_2647,In_692,In_1651);
nand U2648 (N_2648,In_1243,In_47);
and U2649 (N_2649,In_1089,In_1004);
and U2650 (N_2650,In_1843,In_1878);
nand U2651 (N_2651,In_1791,In_1246);
nor U2652 (N_2652,In_525,In_747);
and U2653 (N_2653,In_119,In_1247);
xnor U2654 (N_2654,In_1964,In_590);
and U2655 (N_2655,In_699,In_880);
xnor U2656 (N_2656,In_1910,In_732);
nand U2657 (N_2657,In_994,In_451);
nor U2658 (N_2658,In_1257,In_126);
or U2659 (N_2659,In_507,In_1794);
nor U2660 (N_2660,In_454,In_1372);
xnor U2661 (N_2661,In_413,In_1700);
xor U2662 (N_2662,In_437,In_950);
xor U2663 (N_2663,In_942,In_1281);
and U2664 (N_2664,In_2,In_82);
and U2665 (N_2665,In_1351,In_1144);
nor U2666 (N_2666,In_1953,In_682);
and U2667 (N_2667,In_573,In_1819);
and U2668 (N_2668,In_20,In_912);
nor U2669 (N_2669,In_130,In_159);
nand U2670 (N_2670,In_752,In_1846);
nor U2671 (N_2671,In_1735,In_224);
nand U2672 (N_2672,In_1514,In_1895);
nand U2673 (N_2673,In_1819,In_31);
xor U2674 (N_2674,In_1909,In_1054);
nor U2675 (N_2675,In_478,In_279);
nor U2676 (N_2676,In_1645,In_887);
nand U2677 (N_2677,In_1855,In_1642);
and U2678 (N_2678,In_1607,In_572);
xor U2679 (N_2679,In_553,In_361);
nand U2680 (N_2680,In_380,In_387);
or U2681 (N_2681,In_1701,In_1961);
or U2682 (N_2682,In_1055,In_768);
nand U2683 (N_2683,In_1406,In_1103);
nand U2684 (N_2684,In_456,In_600);
nand U2685 (N_2685,In_1473,In_458);
and U2686 (N_2686,In_732,In_1777);
xor U2687 (N_2687,In_1108,In_396);
and U2688 (N_2688,In_678,In_1382);
nand U2689 (N_2689,In_1981,In_900);
xor U2690 (N_2690,In_1575,In_1387);
or U2691 (N_2691,In_278,In_804);
xnor U2692 (N_2692,In_1856,In_557);
or U2693 (N_2693,In_1395,In_1473);
nor U2694 (N_2694,In_1693,In_1069);
and U2695 (N_2695,In_685,In_305);
and U2696 (N_2696,In_24,In_1032);
or U2697 (N_2697,In_630,In_1455);
xor U2698 (N_2698,In_1962,In_485);
nand U2699 (N_2699,In_1739,In_1697);
nor U2700 (N_2700,In_830,In_601);
nand U2701 (N_2701,In_462,In_195);
nand U2702 (N_2702,In_1845,In_1755);
or U2703 (N_2703,In_1699,In_1866);
nor U2704 (N_2704,In_634,In_1859);
nand U2705 (N_2705,In_1246,In_1963);
or U2706 (N_2706,In_826,In_1862);
nand U2707 (N_2707,In_579,In_188);
or U2708 (N_2708,In_83,In_298);
and U2709 (N_2709,In_1687,In_1517);
and U2710 (N_2710,In_61,In_1991);
or U2711 (N_2711,In_1786,In_1699);
nor U2712 (N_2712,In_251,In_1654);
and U2713 (N_2713,In_341,In_1061);
and U2714 (N_2714,In_121,In_1519);
nand U2715 (N_2715,In_541,In_1081);
nand U2716 (N_2716,In_1170,In_1059);
or U2717 (N_2717,In_1119,In_723);
or U2718 (N_2718,In_1206,In_286);
or U2719 (N_2719,In_1594,In_1292);
xor U2720 (N_2720,In_971,In_517);
nor U2721 (N_2721,In_1283,In_391);
nor U2722 (N_2722,In_1147,In_470);
and U2723 (N_2723,In_1864,In_922);
or U2724 (N_2724,In_1523,In_1355);
and U2725 (N_2725,In_104,In_748);
nand U2726 (N_2726,In_1595,In_821);
nor U2727 (N_2727,In_896,In_1218);
nand U2728 (N_2728,In_633,In_455);
and U2729 (N_2729,In_1051,In_136);
nor U2730 (N_2730,In_358,In_1467);
and U2731 (N_2731,In_1903,In_266);
and U2732 (N_2732,In_1836,In_1386);
nor U2733 (N_2733,In_1432,In_1473);
nand U2734 (N_2734,In_396,In_1816);
nand U2735 (N_2735,In_1636,In_717);
nand U2736 (N_2736,In_1831,In_1053);
and U2737 (N_2737,In_1648,In_242);
nand U2738 (N_2738,In_1826,In_231);
or U2739 (N_2739,In_739,In_1767);
nor U2740 (N_2740,In_1890,In_1917);
or U2741 (N_2741,In_1224,In_852);
and U2742 (N_2742,In_687,In_744);
or U2743 (N_2743,In_1382,In_1743);
nor U2744 (N_2744,In_478,In_561);
or U2745 (N_2745,In_1047,In_1505);
or U2746 (N_2746,In_16,In_1890);
nand U2747 (N_2747,In_444,In_781);
and U2748 (N_2748,In_1236,In_1955);
and U2749 (N_2749,In_2,In_1169);
and U2750 (N_2750,In_190,In_1573);
nand U2751 (N_2751,In_382,In_1479);
nor U2752 (N_2752,In_1503,In_1866);
and U2753 (N_2753,In_833,In_16);
nor U2754 (N_2754,In_606,In_1679);
or U2755 (N_2755,In_851,In_710);
or U2756 (N_2756,In_558,In_369);
nor U2757 (N_2757,In_1141,In_1955);
nor U2758 (N_2758,In_1844,In_663);
or U2759 (N_2759,In_792,In_1322);
nor U2760 (N_2760,In_621,In_1039);
or U2761 (N_2761,In_1230,In_1210);
xnor U2762 (N_2762,In_1949,In_1170);
nand U2763 (N_2763,In_1425,In_1430);
nor U2764 (N_2764,In_401,In_1822);
nor U2765 (N_2765,In_1538,In_685);
and U2766 (N_2766,In_547,In_1279);
and U2767 (N_2767,In_1570,In_1619);
xor U2768 (N_2768,In_722,In_548);
or U2769 (N_2769,In_1321,In_1423);
nor U2770 (N_2770,In_1036,In_1159);
or U2771 (N_2771,In_1131,In_77);
or U2772 (N_2772,In_1560,In_187);
and U2773 (N_2773,In_356,In_1746);
and U2774 (N_2774,In_886,In_463);
nor U2775 (N_2775,In_1836,In_1879);
nor U2776 (N_2776,In_1315,In_1045);
nand U2777 (N_2777,In_1995,In_906);
nand U2778 (N_2778,In_1418,In_469);
nand U2779 (N_2779,In_754,In_1369);
and U2780 (N_2780,In_1808,In_423);
nand U2781 (N_2781,In_1518,In_510);
and U2782 (N_2782,In_609,In_1675);
nor U2783 (N_2783,In_1782,In_958);
nand U2784 (N_2784,In_911,In_1478);
or U2785 (N_2785,In_1760,In_175);
or U2786 (N_2786,In_1212,In_1449);
or U2787 (N_2787,In_1111,In_375);
or U2788 (N_2788,In_1030,In_1252);
xnor U2789 (N_2789,In_1173,In_1638);
xor U2790 (N_2790,In_149,In_1158);
and U2791 (N_2791,In_471,In_1698);
and U2792 (N_2792,In_362,In_983);
or U2793 (N_2793,In_931,In_1179);
and U2794 (N_2794,In_259,In_634);
nor U2795 (N_2795,In_769,In_553);
nor U2796 (N_2796,In_890,In_528);
nand U2797 (N_2797,In_493,In_805);
nand U2798 (N_2798,In_1071,In_640);
nand U2799 (N_2799,In_1388,In_1917);
nor U2800 (N_2800,In_1744,In_1429);
nand U2801 (N_2801,In_263,In_998);
or U2802 (N_2802,In_1267,In_483);
nand U2803 (N_2803,In_317,In_266);
nor U2804 (N_2804,In_1074,In_1076);
xnor U2805 (N_2805,In_309,In_1412);
or U2806 (N_2806,In_170,In_458);
nor U2807 (N_2807,In_20,In_1215);
or U2808 (N_2808,In_1399,In_819);
nand U2809 (N_2809,In_667,In_1694);
nor U2810 (N_2810,In_738,In_512);
nor U2811 (N_2811,In_476,In_60);
nor U2812 (N_2812,In_268,In_1533);
xor U2813 (N_2813,In_1228,In_53);
nand U2814 (N_2814,In_1238,In_1170);
nor U2815 (N_2815,In_405,In_1857);
or U2816 (N_2816,In_1257,In_639);
nor U2817 (N_2817,In_1786,In_151);
nand U2818 (N_2818,In_1752,In_14);
and U2819 (N_2819,In_1509,In_211);
nor U2820 (N_2820,In_1293,In_804);
or U2821 (N_2821,In_1974,In_1810);
nand U2822 (N_2822,In_1923,In_1670);
nor U2823 (N_2823,In_1484,In_53);
nor U2824 (N_2824,In_1810,In_700);
nor U2825 (N_2825,In_726,In_176);
nand U2826 (N_2826,In_1659,In_715);
nor U2827 (N_2827,In_356,In_1279);
or U2828 (N_2828,In_1591,In_1760);
nor U2829 (N_2829,In_740,In_753);
nor U2830 (N_2830,In_1563,In_265);
and U2831 (N_2831,In_1610,In_1569);
nor U2832 (N_2832,In_498,In_553);
nand U2833 (N_2833,In_825,In_1090);
nand U2834 (N_2834,In_1097,In_110);
or U2835 (N_2835,In_1488,In_935);
nor U2836 (N_2836,In_1376,In_1056);
nand U2837 (N_2837,In_1599,In_1542);
xnor U2838 (N_2838,In_158,In_852);
nor U2839 (N_2839,In_1688,In_1081);
nand U2840 (N_2840,In_989,In_1475);
and U2841 (N_2841,In_116,In_845);
or U2842 (N_2842,In_1400,In_98);
nand U2843 (N_2843,In_1199,In_1802);
or U2844 (N_2844,In_276,In_614);
or U2845 (N_2845,In_330,In_71);
and U2846 (N_2846,In_1084,In_1042);
or U2847 (N_2847,In_386,In_1980);
nor U2848 (N_2848,In_1010,In_21);
or U2849 (N_2849,In_1125,In_98);
nand U2850 (N_2850,In_1058,In_949);
nor U2851 (N_2851,In_1848,In_1487);
or U2852 (N_2852,In_1933,In_1013);
nand U2853 (N_2853,In_1939,In_1501);
xor U2854 (N_2854,In_541,In_589);
and U2855 (N_2855,In_1809,In_351);
and U2856 (N_2856,In_1521,In_884);
or U2857 (N_2857,In_1077,In_716);
and U2858 (N_2858,In_1708,In_1736);
nor U2859 (N_2859,In_1024,In_1499);
nor U2860 (N_2860,In_1985,In_1780);
nor U2861 (N_2861,In_1412,In_1091);
or U2862 (N_2862,In_1411,In_1438);
nor U2863 (N_2863,In_815,In_1370);
nand U2864 (N_2864,In_217,In_342);
nand U2865 (N_2865,In_216,In_404);
nor U2866 (N_2866,In_995,In_751);
nor U2867 (N_2867,In_8,In_715);
nor U2868 (N_2868,In_1758,In_25);
and U2869 (N_2869,In_959,In_130);
nand U2870 (N_2870,In_958,In_1255);
or U2871 (N_2871,In_1526,In_227);
nand U2872 (N_2872,In_1335,In_263);
nand U2873 (N_2873,In_1373,In_1285);
nor U2874 (N_2874,In_322,In_218);
nor U2875 (N_2875,In_1358,In_939);
nor U2876 (N_2876,In_585,In_1299);
or U2877 (N_2877,In_1589,In_1068);
or U2878 (N_2878,In_1304,In_1129);
nand U2879 (N_2879,In_903,In_74);
nand U2880 (N_2880,In_1040,In_882);
or U2881 (N_2881,In_288,In_1125);
nand U2882 (N_2882,In_1934,In_1035);
xor U2883 (N_2883,In_1042,In_1432);
nand U2884 (N_2884,In_656,In_4);
nor U2885 (N_2885,In_170,In_1547);
nand U2886 (N_2886,In_500,In_250);
or U2887 (N_2887,In_721,In_1652);
nand U2888 (N_2888,In_784,In_650);
or U2889 (N_2889,In_842,In_191);
nand U2890 (N_2890,In_37,In_1355);
nor U2891 (N_2891,In_290,In_1227);
nand U2892 (N_2892,In_1096,In_1727);
nor U2893 (N_2893,In_899,In_132);
or U2894 (N_2894,In_799,In_772);
and U2895 (N_2895,In_1296,In_531);
or U2896 (N_2896,In_374,In_243);
nor U2897 (N_2897,In_1416,In_32);
xnor U2898 (N_2898,In_1227,In_953);
xnor U2899 (N_2899,In_162,In_1101);
and U2900 (N_2900,In_991,In_400);
or U2901 (N_2901,In_1875,In_1800);
xor U2902 (N_2902,In_1752,In_1334);
nand U2903 (N_2903,In_7,In_56);
or U2904 (N_2904,In_727,In_525);
nor U2905 (N_2905,In_891,In_1703);
and U2906 (N_2906,In_270,In_762);
nor U2907 (N_2907,In_560,In_1046);
or U2908 (N_2908,In_410,In_1903);
nand U2909 (N_2909,In_1322,In_415);
or U2910 (N_2910,In_1158,In_226);
and U2911 (N_2911,In_186,In_610);
nor U2912 (N_2912,In_1369,In_1502);
xor U2913 (N_2913,In_1012,In_686);
nand U2914 (N_2914,In_974,In_395);
or U2915 (N_2915,In_650,In_126);
and U2916 (N_2916,In_381,In_289);
or U2917 (N_2917,In_728,In_956);
nand U2918 (N_2918,In_1375,In_1249);
nor U2919 (N_2919,In_448,In_92);
nor U2920 (N_2920,In_1094,In_57);
or U2921 (N_2921,In_732,In_1988);
or U2922 (N_2922,In_842,In_1037);
nand U2923 (N_2923,In_575,In_796);
or U2924 (N_2924,In_553,In_1726);
xor U2925 (N_2925,In_1379,In_260);
nand U2926 (N_2926,In_1884,In_604);
or U2927 (N_2927,In_90,In_436);
nand U2928 (N_2928,In_415,In_1871);
nand U2929 (N_2929,In_1412,In_1284);
nor U2930 (N_2930,In_949,In_508);
and U2931 (N_2931,In_1697,In_368);
nand U2932 (N_2932,In_196,In_408);
nor U2933 (N_2933,In_1657,In_1430);
or U2934 (N_2934,In_811,In_1555);
xnor U2935 (N_2935,In_873,In_1904);
or U2936 (N_2936,In_683,In_816);
nand U2937 (N_2937,In_270,In_1257);
nand U2938 (N_2938,In_1921,In_234);
or U2939 (N_2939,In_1602,In_336);
or U2940 (N_2940,In_184,In_863);
nor U2941 (N_2941,In_1522,In_97);
nor U2942 (N_2942,In_1331,In_982);
nand U2943 (N_2943,In_622,In_1575);
and U2944 (N_2944,In_620,In_943);
nor U2945 (N_2945,In_1476,In_495);
and U2946 (N_2946,In_675,In_936);
nand U2947 (N_2947,In_1650,In_529);
nor U2948 (N_2948,In_670,In_1012);
xor U2949 (N_2949,In_50,In_609);
and U2950 (N_2950,In_1279,In_550);
and U2951 (N_2951,In_286,In_1513);
xnor U2952 (N_2952,In_1482,In_1453);
or U2953 (N_2953,In_1832,In_1063);
and U2954 (N_2954,In_866,In_239);
and U2955 (N_2955,In_1106,In_1827);
and U2956 (N_2956,In_1286,In_1142);
nand U2957 (N_2957,In_1060,In_1432);
and U2958 (N_2958,In_573,In_1102);
or U2959 (N_2959,In_1450,In_406);
nand U2960 (N_2960,In_854,In_619);
and U2961 (N_2961,In_988,In_1502);
or U2962 (N_2962,In_510,In_692);
and U2963 (N_2963,In_780,In_1900);
or U2964 (N_2964,In_1219,In_985);
or U2965 (N_2965,In_1197,In_1439);
xor U2966 (N_2966,In_314,In_1292);
nor U2967 (N_2967,In_1202,In_957);
nor U2968 (N_2968,In_1901,In_921);
nand U2969 (N_2969,In_1859,In_545);
xnor U2970 (N_2970,In_1214,In_1649);
nor U2971 (N_2971,In_8,In_721);
or U2972 (N_2972,In_116,In_1106);
nand U2973 (N_2973,In_38,In_444);
or U2974 (N_2974,In_991,In_817);
and U2975 (N_2975,In_1820,In_1841);
nor U2976 (N_2976,In_1757,In_1679);
and U2977 (N_2977,In_1203,In_10);
or U2978 (N_2978,In_875,In_1578);
nor U2979 (N_2979,In_662,In_1991);
nand U2980 (N_2980,In_207,In_450);
nand U2981 (N_2981,In_426,In_931);
or U2982 (N_2982,In_1615,In_245);
nor U2983 (N_2983,In_1667,In_180);
and U2984 (N_2984,In_611,In_927);
xnor U2985 (N_2985,In_815,In_632);
nand U2986 (N_2986,In_1721,In_1768);
nand U2987 (N_2987,In_93,In_46);
nand U2988 (N_2988,In_176,In_1480);
nand U2989 (N_2989,In_1432,In_1315);
and U2990 (N_2990,In_1685,In_1531);
xnor U2991 (N_2991,In_1422,In_1993);
nor U2992 (N_2992,In_1047,In_752);
or U2993 (N_2993,In_64,In_1525);
nor U2994 (N_2994,In_561,In_332);
and U2995 (N_2995,In_150,In_22);
xor U2996 (N_2996,In_403,In_214);
nand U2997 (N_2997,In_137,In_18);
nand U2998 (N_2998,In_1119,In_1813);
or U2999 (N_2999,In_626,In_1235);
or U3000 (N_3000,In_8,In_1881);
nand U3001 (N_3001,In_948,In_1464);
nand U3002 (N_3002,In_1881,In_1485);
or U3003 (N_3003,In_1058,In_443);
and U3004 (N_3004,In_1754,In_849);
xor U3005 (N_3005,In_432,In_1076);
nor U3006 (N_3006,In_1391,In_899);
nand U3007 (N_3007,In_347,In_1830);
and U3008 (N_3008,In_1302,In_194);
or U3009 (N_3009,In_1212,In_14);
and U3010 (N_3010,In_1797,In_344);
nor U3011 (N_3011,In_393,In_183);
and U3012 (N_3012,In_1899,In_1050);
or U3013 (N_3013,In_1597,In_1092);
or U3014 (N_3014,In_687,In_1423);
and U3015 (N_3015,In_644,In_722);
or U3016 (N_3016,In_342,In_481);
nand U3017 (N_3017,In_603,In_1075);
and U3018 (N_3018,In_1104,In_1111);
nor U3019 (N_3019,In_121,In_115);
and U3020 (N_3020,In_260,In_1864);
nor U3021 (N_3021,In_594,In_1029);
nor U3022 (N_3022,In_461,In_1705);
nand U3023 (N_3023,In_1576,In_233);
or U3024 (N_3024,In_1017,In_1785);
nor U3025 (N_3025,In_614,In_6);
nor U3026 (N_3026,In_1719,In_56);
or U3027 (N_3027,In_1658,In_469);
nor U3028 (N_3028,In_111,In_429);
and U3029 (N_3029,In_1117,In_1356);
nor U3030 (N_3030,In_906,In_431);
and U3031 (N_3031,In_1922,In_1769);
and U3032 (N_3032,In_212,In_1203);
and U3033 (N_3033,In_732,In_1799);
and U3034 (N_3034,In_1642,In_960);
xor U3035 (N_3035,In_1003,In_1851);
nor U3036 (N_3036,In_646,In_701);
nor U3037 (N_3037,In_293,In_1871);
or U3038 (N_3038,In_1978,In_938);
nor U3039 (N_3039,In_680,In_260);
nand U3040 (N_3040,In_1483,In_1521);
and U3041 (N_3041,In_1567,In_361);
or U3042 (N_3042,In_1535,In_231);
or U3043 (N_3043,In_1444,In_483);
or U3044 (N_3044,In_732,In_559);
nor U3045 (N_3045,In_330,In_1494);
xnor U3046 (N_3046,In_1739,In_1520);
or U3047 (N_3047,In_734,In_1230);
and U3048 (N_3048,In_794,In_1638);
or U3049 (N_3049,In_320,In_717);
nor U3050 (N_3050,In_746,In_838);
nand U3051 (N_3051,In_1756,In_415);
xor U3052 (N_3052,In_614,In_909);
or U3053 (N_3053,In_116,In_20);
and U3054 (N_3054,In_185,In_1342);
and U3055 (N_3055,In_1601,In_1979);
and U3056 (N_3056,In_730,In_748);
xor U3057 (N_3057,In_749,In_1882);
nor U3058 (N_3058,In_1141,In_1634);
or U3059 (N_3059,In_1865,In_523);
and U3060 (N_3060,In_1219,In_1379);
nand U3061 (N_3061,In_274,In_1876);
or U3062 (N_3062,In_329,In_1313);
and U3063 (N_3063,In_1491,In_651);
nor U3064 (N_3064,In_805,In_293);
nand U3065 (N_3065,In_1795,In_1550);
nand U3066 (N_3066,In_1474,In_330);
nor U3067 (N_3067,In_919,In_1419);
nor U3068 (N_3068,In_1528,In_33);
nand U3069 (N_3069,In_1175,In_1848);
nand U3070 (N_3070,In_973,In_1290);
and U3071 (N_3071,In_1828,In_147);
nor U3072 (N_3072,In_577,In_1501);
or U3073 (N_3073,In_954,In_1889);
nand U3074 (N_3074,In_1154,In_1632);
nor U3075 (N_3075,In_228,In_759);
xor U3076 (N_3076,In_1052,In_1721);
nand U3077 (N_3077,In_1609,In_586);
nor U3078 (N_3078,In_75,In_1812);
nor U3079 (N_3079,In_633,In_442);
nor U3080 (N_3080,In_1317,In_348);
nand U3081 (N_3081,In_883,In_645);
nor U3082 (N_3082,In_469,In_748);
nand U3083 (N_3083,In_657,In_360);
nor U3084 (N_3084,In_135,In_1788);
and U3085 (N_3085,In_206,In_190);
nand U3086 (N_3086,In_1492,In_1700);
or U3087 (N_3087,In_149,In_1064);
nor U3088 (N_3088,In_285,In_1641);
or U3089 (N_3089,In_1881,In_659);
nand U3090 (N_3090,In_1458,In_1113);
nor U3091 (N_3091,In_1485,In_1098);
xnor U3092 (N_3092,In_1046,In_1458);
or U3093 (N_3093,In_1517,In_1578);
and U3094 (N_3094,In_1293,In_769);
and U3095 (N_3095,In_1666,In_218);
or U3096 (N_3096,In_917,In_610);
or U3097 (N_3097,In_433,In_1255);
nand U3098 (N_3098,In_141,In_1174);
and U3099 (N_3099,In_1497,In_1291);
nor U3100 (N_3100,In_137,In_875);
or U3101 (N_3101,In_1941,In_1249);
nand U3102 (N_3102,In_1236,In_199);
xor U3103 (N_3103,In_1601,In_1704);
or U3104 (N_3104,In_639,In_1922);
or U3105 (N_3105,In_606,In_193);
nand U3106 (N_3106,In_601,In_1291);
or U3107 (N_3107,In_509,In_1932);
and U3108 (N_3108,In_70,In_1927);
nand U3109 (N_3109,In_450,In_1504);
or U3110 (N_3110,In_267,In_574);
and U3111 (N_3111,In_1566,In_571);
and U3112 (N_3112,In_1295,In_1567);
nand U3113 (N_3113,In_548,In_1658);
or U3114 (N_3114,In_971,In_1680);
nor U3115 (N_3115,In_94,In_1539);
and U3116 (N_3116,In_1118,In_951);
or U3117 (N_3117,In_1142,In_23);
nand U3118 (N_3118,In_1962,In_1646);
nand U3119 (N_3119,In_1590,In_1671);
nand U3120 (N_3120,In_1135,In_483);
and U3121 (N_3121,In_323,In_1026);
nand U3122 (N_3122,In_1236,In_422);
and U3123 (N_3123,In_1229,In_1208);
and U3124 (N_3124,In_175,In_1138);
nor U3125 (N_3125,In_1054,In_488);
xnor U3126 (N_3126,In_1785,In_1140);
nand U3127 (N_3127,In_994,In_1998);
nor U3128 (N_3128,In_1451,In_363);
nor U3129 (N_3129,In_1330,In_1585);
or U3130 (N_3130,In_917,In_664);
nand U3131 (N_3131,In_1334,In_1171);
xnor U3132 (N_3132,In_1323,In_1024);
nand U3133 (N_3133,In_1363,In_661);
xnor U3134 (N_3134,In_59,In_717);
nor U3135 (N_3135,In_990,In_1868);
or U3136 (N_3136,In_358,In_1540);
and U3137 (N_3137,In_742,In_190);
or U3138 (N_3138,In_1811,In_684);
nor U3139 (N_3139,In_868,In_1061);
or U3140 (N_3140,In_1475,In_1642);
nor U3141 (N_3141,In_1104,In_883);
or U3142 (N_3142,In_351,In_1780);
and U3143 (N_3143,In_1702,In_1884);
and U3144 (N_3144,In_1666,In_1781);
xor U3145 (N_3145,In_846,In_1086);
or U3146 (N_3146,In_515,In_667);
and U3147 (N_3147,In_1160,In_873);
nand U3148 (N_3148,In_1350,In_22);
xnor U3149 (N_3149,In_203,In_1649);
or U3150 (N_3150,In_1699,In_1963);
and U3151 (N_3151,In_344,In_1812);
nand U3152 (N_3152,In_1066,In_909);
nor U3153 (N_3153,In_634,In_1738);
nor U3154 (N_3154,In_744,In_1580);
or U3155 (N_3155,In_151,In_777);
nor U3156 (N_3156,In_28,In_739);
nor U3157 (N_3157,In_1943,In_1052);
and U3158 (N_3158,In_990,In_913);
nand U3159 (N_3159,In_156,In_1999);
nor U3160 (N_3160,In_1643,In_1760);
or U3161 (N_3161,In_1770,In_315);
nor U3162 (N_3162,In_778,In_505);
nor U3163 (N_3163,In_1443,In_1176);
or U3164 (N_3164,In_1414,In_1777);
or U3165 (N_3165,In_1314,In_1756);
nand U3166 (N_3166,In_1611,In_1422);
xnor U3167 (N_3167,In_1185,In_1407);
and U3168 (N_3168,In_1478,In_1815);
and U3169 (N_3169,In_539,In_1333);
nand U3170 (N_3170,In_1593,In_1240);
or U3171 (N_3171,In_987,In_805);
or U3172 (N_3172,In_914,In_1936);
nand U3173 (N_3173,In_1681,In_1269);
and U3174 (N_3174,In_154,In_1883);
or U3175 (N_3175,In_920,In_162);
xor U3176 (N_3176,In_1745,In_670);
or U3177 (N_3177,In_189,In_1269);
and U3178 (N_3178,In_384,In_1416);
nor U3179 (N_3179,In_290,In_1600);
nor U3180 (N_3180,In_598,In_1750);
or U3181 (N_3181,In_1166,In_72);
nor U3182 (N_3182,In_471,In_1231);
or U3183 (N_3183,In_1928,In_1060);
and U3184 (N_3184,In_929,In_1999);
nor U3185 (N_3185,In_367,In_638);
nand U3186 (N_3186,In_633,In_1121);
and U3187 (N_3187,In_837,In_732);
or U3188 (N_3188,In_1180,In_1770);
nand U3189 (N_3189,In_1309,In_420);
or U3190 (N_3190,In_1335,In_1188);
or U3191 (N_3191,In_542,In_101);
nand U3192 (N_3192,In_734,In_101);
or U3193 (N_3193,In_28,In_167);
or U3194 (N_3194,In_1126,In_1434);
nand U3195 (N_3195,In_59,In_434);
nand U3196 (N_3196,In_1459,In_988);
and U3197 (N_3197,In_1614,In_127);
xor U3198 (N_3198,In_202,In_540);
nor U3199 (N_3199,In_1879,In_735);
nand U3200 (N_3200,In_980,In_502);
and U3201 (N_3201,In_1684,In_1197);
or U3202 (N_3202,In_1418,In_1054);
or U3203 (N_3203,In_1529,In_1583);
nand U3204 (N_3204,In_131,In_604);
nor U3205 (N_3205,In_1371,In_1268);
nor U3206 (N_3206,In_353,In_1980);
or U3207 (N_3207,In_376,In_1786);
nand U3208 (N_3208,In_1947,In_1011);
nor U3209 (N_3209,In_1219,In_303);
nand U3210 (N_3210,In_1880,In_1590);
nor U3211 (N_3211,In_1663,In_1896);
or U3212 (N_3212,In_68,In_98);
nand U3213 (N_3213,In_1277,In_270);
and U3214 (N_3214,In_476,In_1121);
or U3215 (N_3215,In_1145,In_984);
nand U3216 (N_3216,In_660,In_557);
nor U3217 (N_3217,In_753,In_62);
nand U3218 (N_3218,In_513,In_1624);
xor U3219 (N_3219,In_270,In_1232);
or U3220 (N_3220,In_686,In_1041);
nor U3221 (N_3221,In_1879,In_292);
nand U3222 (N_3222,In_99,In_746);
nand U3223 (N_3223,In_1633,In_1959);
xnor U3224 (N_3224,In_1209,In_1494);
and U3225 (N_3225,In_1373,In_1969);
and U3226 (N_3226,In_1477,In_784);
nor U3227 (N_3227,In_490,In_1497);
nor U3228 (N_3228,In_1606,In_1309);
nor U3229 (N_3229,In_33,In_1740);
or U3230 (N_3230,In_1831,In_128);
or U3231 (N_3231,In_42,In_932);
or U3232 (N_3232,In_31,In_1545);
or U3233 (N_3233,In_1723,In_630);
nor U3234 (N_3234,In_648,In_86);
or U3235 (N_3235,In_1422,In_1792);
nor U3236 (N_3236,In_1055,In_1107);
nor U3237 (N_3237,In_589,In_1421);
or U3238 (N_3238,In_1922,In_746);
nand U3239 (N_3239,In_920,In_504);
and U3240 (N_3240,In_1635,In_211);
nor U3241 (N_3241,In_1271,In_882);
nand U3242 (N_3242,In_753,In_1308);
and U3243 (N_3243,In_1023,In_721);
or U3244 (N_3244,In_1184,In_635);
nor U3245 (N_3245,In_981,In_141);
xor U3246 (N_3246,In_1592,In_1702);
and U3247 (N_3247,In_838,In_39);
or U3248 (N_3248,In_1387,In_1699);
nand U3249 (N_3249,In_1235,In_489);
nand U3250 (N_3250,In_266,In_1805);
and U3251 (N_3251,In_256,In_1801);
or U3252 (N_3252,In_465,In_1045);
nand U3253 (N_3253,In_142,In_1037);
and U3254 (N_3254,In_787,In_984);
nor U3255 (N_3255,In_1254,In_204);
and U3256 (N_3256,In_1020,In_507);
nor U3257 (N_3257,In_1696,In_1873);
nand U3258 (N_3258,In_918,In_1215);
and U3259 (N_3259,In_1323,In_441);
or U3260 (N_3260,In_540,In_1826);
or U3261 (N_3261,In_11,In_1807);
or U3262 (N_3262,In_271,In_587);
or U3263 (N_3263,In_47,In_1035);
or U3264 (N_3264,In_512,In_1819);
and U3265 (N_3265,In_865,In_1288);
and U3266 (N_3266,In_1827,In_779);
nand U3267 (N_3267,In_827,In_225);
nand U3268 (N_3268,In_1396,In_1060);
nor U3269 (N_3269,In_128,In_814);
xnor U3270 (N_3270,In_67,In_616);
or U3271 (N_3271,In_665,In_1656);
nor U3272 (N_3272,In_709,In_1615);
or U3273 (N_3273,In_1867,In_1615);
nand U3274 (N_3274,In_619,In_596);
nand U3275 (N_3275,In_124,In_1829);
xnor U3276 (N_3276,In_1897,In_1801);
nand U3277 (N_3277,In_1873,In_1101);
xor U3278 (N_3278,In_867,In_951);
nor U3279 (N_3279,In_1268,In_874);
nor U3280 (N_3280,In_638,In_836);
or U3281 (N_3281,In_1930,In_1397);
nand U3282 (N_3282,In_20,In_509);
and U3283 (N_3283,In_1677,In_751);
and U3284 (N_3284,In_616,In_1253);
xor U3285 (N_3285,In_745,In_1723);
and U3286 (N_3286,In_126,In_1203);
nand U3287 (N_3287,In_1071,In_1317);
or U3288 (N_3288,In_406,In_1369);
nor U3289 (N_3289,In_1060,In_1883);
or U3290 (N_3290,In_82,In_1193);
or U3291 (N_3291,In_508,In_1087);
nor U3292 (N_3292,In_1727,In_1823);
nand U3293 (N_3293,In_1989,In_1749);
or U3294 (N_3294,In_744,In_663);
and U3295 (N_3295,In_670,In_860);
nand U3296 (N_3296,In_1610,In_132);
and U3297 (N_3297,In_1429,In_1341);
nand U3298 (N_3298,In_531,In_673);
xor U3299 (N_3299,In_1302,In_1499);
nor U3300 (N_3300,In_520,In_1418);
and U3301 (N_3301,In_1089,In_1352);
nand U3302 (N_3302,In_144,In_552);
and U3303 (N_3303,In_1649,In_409);
nor U3304 (N_3304,In_149,In_1964);
nand U3305 (N_3305,In_1538,In_234);
or U3306 (N_3306,In_1832,In_547);
xor U3307 (N_3307,In_1701,In_216);
and U3308 (N_3308,In_977,In_1330);
nor U3309 (N_3309,In_758,In_662);
nand U3310 (N_3310,In_354,In_574);
or U3311 (N_3311,In_1034,In_664);
nand U3312 (N_3312,In_1763,In_1776);
nor U3313 (N_3313,In_1666,In_104);
nor U3314 (N_3314,In_785,In_466);
nor U3315 (N_3315,In_81,In_115);
and U3316 (N_3316,In_1205,In_91);
nor U3317 (N_3317,In_1957,In_84);
nand U3318 (N_3318,In_1610,In_185);
or U3319 (N_3319,In_643,In_914);
and U3320 (N_3320,In_1769,In_574);
and U3321 (N_3321,In_936,In_1106);
and U3322 (N_3322,In_1588,In_934);
xor U3323 (N_3323,In_1605,In_1370);
or U3324 (N_3324,In_1120,In_516);
or U3325 (N_3325,In_1603,In_1438);
nor U3326 (N_3326,In_688,In_813);
and U3327 (N_3327,In_999,In_668);
and U3328 (N_3328,In_186,In_1403);
and U3329 (N_3329,In_1681,In_1031);
or U3330 (N_3330,In_671,In_120);
xor U3331 (N_3331,In_933,In_1513);
nand U3332 (N_3332,In_1709,In_748);
nor U3333 (N_3333,In_1243,In_132);
nand U3334 (N_3334,In_75,In_1059);
nor U3335 (N_3335,In_777,In_1155);
or U3336 (N_3336,In_567,In_930);
and U3337 (N_3337,In_1811,In_1848);
nand U3338 (N_3338,In_1064,In_974);
or U3339 (N_3339,In_1665,In_1487);
nand U3340 (N_3340,In_1505,In_880);
nand U3341 (N_3341,In_727,In_1284);
or U3342 (N_3342,In_618,In_646);
nand U3343 (N_3343,In_1640,In_1499);
and U3344 (N_3344,In_1154,In_706);
nor U3345 (N_3345,In_1842,In_1699);
nand U3346 (N_3346,In_1260,In_752);
and U3347 (N_3347,In_990,In_377);
or U3348 (N_3348,In_891,In_402);
nand U3349 (N_3349,In_709,In_1916);
nand U3350 (N_3350,In_231,In_544);
and U3351 (N_3351,In_1253,In_1755);
nand U3352 (N_3352,In_32,In_315);
nand U3353 (N_3353,In_765,In_405);
nand U3354 (N_3354,In_10,In_1713);
nor U3355 (N_3355,In_1129,In_497);
nor U3356 (N_3356,In_1280,In_1678);
nor U3357 (N_3357,In_853,In_1206);
and U3358 (N_3358,In_432,In_48);
nor U3359 (N_3359,In_654,In_868);
and U3360 (N_3360,In_95,In_1595);
or U3361 (N_3361,In_399,In_1015);
or U3362 (N_3362,In_93,In_1348);
or U3363 (N_3363,In_993,In_516);
nand U3364 (N_3364,In_1483,In_1533);
and U3365 (N_3365,In_1338,In_1432);
nor U3366 (N_3366,In_989,In_1170);
nor U3367 (N_3367,In_153,In_1444);
and U3368 (N_3368,In_113,In_470);
nand U3369 (N_3369,In_428,In_1793);
nand U3370 (N_3370,In_1646,In_1723);
or U3371 (N_3371,In_1726,In_18);
nand U3372 (N_3372,In_470,In_1804);
nand U3373 (N_3373,In_603,In_595);
xor U3374 (N_3374,In_1221,In_1780);
and U3375 (N_3375,In_558,In_1266);
nand U3376 (N_3376,In_1714,In_1302);
nor U3377 (N_3377,In_95,In_1137);
or U3378 (N_3378,In_387,In_695);
or U3379 (N_3379,In_617,In_1300);
nor U3380 (N_3380,In_1487,In_948);
nand U3381 (N_3381,In_1353,In_1000);
xor U3382 (N_3382,In_105,In_1156);
and U3383 (N_3383,In_589,In_1040);
xnor U3384 (N_3384,In_478,In_976);
and U3385 (N_3385,In_937,In_1974);
or U3386 (N_3386,In_921,In_1675);
and U3387 (N_3387,In_1365,In_1843);
nor U3388 (N_3388,In_160,In_1176);
and U3389 (N_3389,In_1934,In_1675);
and U3390 (N_3390,In_1983,In_1132);
nor U3391 (N_3391,In_387,In_108);
and U3392 (N_3392,In_1820,In_910);
or U3393 (N_3393,In_936,In_486);
and U3394 (N_3394,In_1886,In_1215);
and U3395 (N_3395,In_3,In_247);
xor U3396 (N_3396,In_1622,In_862);
and U3397 (N_3397,In_1351,In_532);
and U3398 (N_3398,In_616,In_1152);
or U3399 (N_3399,In_276,In_1769);
nand U3400 (N_3400,In_146,In_1879);
xor U3401 (N_3401,In_306,In_1166);
or U3402 (N_3402,In_946,In_1108);
xnor U3403 (N_3403,In_714,In_504);
nand U3404 (N_3404,In_1046,In_991);
and U3405 (N_3405,In_1750,In_317);
and U3406 (N_3406,In_391,In_1035);
nor U3407 (N_3407,In_1039,In_1181);
xor U3408 (N_3408,In_1342,In_207);
and U3409 (N_3409,In_1563,In_761);
nand U3410 (N_3410,In_87,In_1684);
nor U3411 (N_3411,In_74,In_580);
and U3412 (N_3412,In_778,In_1093);
and U3413 (N_3413,In_1764,In_1904);
nand U3414 (N_3414,In_1464,In_1973);
or U3415 (N_3415,In_46,In_1370);
nor U3416 (N_3416,In_55,In_1333);
nor U3417 (N_3417,In_1735,In_534);
nor U3418 (N_3418,In_1017,In_1583);
or U3419 (N_3419,In_493,In_347);
nand U3420 (N_3420,In_881,In_1453);
nand U3421 (N_3421,In_591,In_1299);
or U3422 (N_3422,In_234,In_740);
xor U3423 (N_3423,In_329,In_974);
or U3424 (N_3424,In_1716,In_932);
or U3425 (N_3425,In_1443,In_25);
or U3426 (N_3426,In_1452,In_131);
or U3427 (N_3427,In_383,In_5);
nand U3428 (N_3428,In_1710,In_767);
nor U3429 (N_3429,In_279,In_492);
nor U3430 (N_3430,In_1241,In_364);
and U3431 (N_3431,In_420,In_714);
or U3432 (N_3432,In_94,In_1019);
and U3433 (N_3433,In_255,In_1813);
and U3434 (N_3434,In_709,In_508);
nor U3435 (N_3435,In_474,In_929);
and U3436 (N_3436,In_1398,In_1793);
and U3437 (N_3437,In_1264,In_810);
or U3438 (N_3438,In_712,In_1386);
or U3439 (N_3439,In_663,In_1854);
nor U3440 (N_3440,In_1506,In_1240);
xor U3441 (N_3441,In_332,In_1020);
nand U3442 (N_3442,In_833,In_819);
xnor U3443 (N_3443,In_1032,In_771);
nor U3444 (N_3444,In_1757,In_1580);
nand U3445 (N_3445,In_1501,In_1992);
nor U3446 (N_3446,In_1495,In_373);
or U3447 (N_3447,In_1166,In_1678);
or U3448 (N_3448,In_788,In_442);
nor U3449 (N_3449,In_1435,In_1162);
or U3450 (N_3450,In_133,In_426);
and U3451 (N_3451,In_1757,In_391);
and U3452 (N_3452,In_487,In_1826);
nand U3453 (N_3453,In_238,In_790);
and U3454 (N_3454,In_376,In_336);
nand U3455 (N_3455,In_1050,In_1157);
and U3456 (N_3456,In_1597,In_1991);
or U3457 (N_3457,In_371,In_676);
or U3458 (N_3458,In_1126,In_488);
or U3459 (N_3459,In_1530,In_667);
and U3460 (N_3460,In_231,In_1287);
nor U3461 (N_3461,In_1629,In_667);
nand U3462 (N_3462,In_340,In_339);
nor U3463 (N_3463,In_1276,In_231);
nand U3464 (N_3464,In_619,In_1760);
xnor U3465 (N_3465,In_1576,In_114);
nand U3466 (N_3466,In_197,In_1557);
and U3467 (N_3467,In_1787,In_580);
xor U3468 (N_3468,In_18,In_1575);
or U3469 (N_3469,In_1882,In_1817);
nor U3470 (N_3470,In_1450,In_705);
nor U3471 (N_3471,In_878,In_248);
nand U3472 (N_3472,In_545,In_49);
nor U3473 (N_3473,In_1070,In_1451);
nand U3474 (N_3474,In_381,In_1124);
nor U3475 (N_3475,In_303,In_402);
xor U3476 (N_3476,In_1476,In_729);
and U3477 (N_3477,In_383,In_460);
and U3478 (N_3478,In_1887,In_459);
nand U3479 (N_3479,In_405,In_1310);
or U3480 (N_3480,In_159,In_683);
xnor U3481 (N_3481,In_1169,In_1291);
xnor U3482 (N_3482,In_528,In_1031);
or U3483 (N_3483,In_1097,In_910);
or U3484 (N_3484,In_992,In_1755);
nand U3485 (N_3485,In_362,In_1712);
or U3486 (N_3486,In_1908,In_785);
nand U3487 (N_3487,In_489,In_1607);
and U3488 (N_3488,In_1188,In_340);
nand U3489 (N_3489,In_646,In_1685);
and U3490 (N_3490,In_1609,In_1017);
xnor U3491 (N_3491,In_487,In_751);
nor U3492 (N_3492,In_1559,In_784);
nand U3493 (N_3493,In_1522,In_871);
nand U3494 (N_3494,In_1670,In_418);
nand U3495 (N_3495,In_53,In_527);
or U3496 (N_3496,In_1771,In_202);
nor U3497 (N_3497,In_48,In_504);
nor U3498 (N_3498,In_686,In_1063);
or U3499 (N_3499,In_1104,In_229);
xnor U3500 (N_3500,In_353,In_1639);
and U3501 (N_3501,In_1950,In_604);
or U3502 (N_3502,In_229,In_592);
nand U3503 (N_3503,In_92,In_1998);
or U3504 (N_3504,In_954,In_1360);
or U3505 (N_3505,In_1500,In_656);
nand U3506 (N_3506,In_1506,In_815);
nor U3507 (N_3507,In_1086,In_1112);
or U3508 (N_3508,In_493,In_1588);
or U3509 (N_3509,In_665,In_910);
and U3510 (N_3510,In_137,In_644);
nand U3511 (N_3511,In_1502,In_1894);
nor U3512 (N_3512,In_1522,In_936);
xor U3513 (N_3513,In_1783,In_1116);
xor U3514 (N_3514,In_1015,In_382);
nor U3515 (N_3515,In_265,In_387);
and U3516 (N_3516,In_179,In_1858);
nor U3517 (N_3517,In_563,In_1928);
or U3518 (N_3518,In_1794,In_1354);
xnor U3519 (N_3519,In_1604,In_639);
nand U3520 (N_3520,In_1306,In_916);
xor U3521 (N_3521,In_1968,In_765);
and U3522 (N_3522,In_1515,In_1359);
and U3523 (N_3523,In_1837,In_1400);
nor U3524 (N_3524,In_275,In_1907);
or U3525 (N_3525,In_500,In_754);
nand U3526 (N_3526,In_282,In_287);
and U3527 (N_3527,In_664,In_353);
or U3528 (N_3528,In_356,In_316);
and U3529 (N_3529,In_1305,In_447);
nor U3530 (N_3530,In_449,In_1994);
or U3531 (N_3531,In_1345,In_1329);
or U3532 (N_3532,In_1436,In_111);
or U3533 (N_3533,In_889,In_82);
or U3534 (N_3534,In_789,In_502);
nor U3535 (N_3535,In_276,In_391);
xor U3536 (N_3536,In_369,In_765);
nor U3537 (N_3537,In_700,In_589);
and U3538 (N_3538,In_1303,In_948);
and U3539 (N_3539,In_1076,In_907);
xor U3540 (N_3540,In_324,In_1868);
and U3541 (N_3541,In_1456,In_259);
nor U3542 (N_3542,In_398,In_1049);
and U3543 (N_3543,In_229,In_1888);
or U3544 (N_3544,In_1520,In_1126);
nand U3545 (N_3545,In_1654,In_151);
and U3546 (N_3546,In_608,In_450);
and U3547 (N_3547,In_162,In_142);
or U3548 (N_3548,In_800,In_294);
and U3549 (N_3549,In_258,In_767);
xor U3550 (N_3550,In_930,In_759);
and U3551 (N_3551,In_140,In_110);
and U3552 (N_3552,In_529,In_941);
nand U3553 (N_3553,In_1211,In_1014);
or U3554 (N_3554,In_684,In_889);
or U3555 (N_3555,In_314,In_1074);
nand U3556 (N_3556,In_1879,In_1761);
and U3557 (N_3557,In_253,In_1452);
xor U3558 (N_3558,In_1341,In_856);
nor U3559 (N_3559,In_658,In_1516);
and U3560 (N_3560,In_1138,In_947);
nor U3561 (N_3561,In_1114,In_0);
xnor U3562 (N_3562,In_31,In_1749);
and U3563 (N_3563,In_926,In_728);
and U3564 (N_3564,In_1992,In_899);
nand U3565 (N_3565,In_378,In_878);
nor U3566 (N_3566,In_274,In_1914);
xor U3567 (N_3567,In_367,In_1535);
and U3568 (N_3568,In_1260,In_1932);
nand U3569 (N_3569,In_945,In_592);
nand U3570 (N_3570,In_1993,In_1080);
and U3571 (N_3571,In_829,In_1242);
nand U3572 (N_3572,In_1756,In_411);
or U3573 (N_3573,In_465,In_1435);
or U3574 (N_3574,In_25,In_39);
nor U3575 (N_3575,In_1007,In_1962);
xor U3576 (N_3576,In_85,In_1795);
and U3577 (N_3577,In_751,In_1063);
nand U3578 (N_3578,In_1432,In_1760);
nor U3579 (N_3579,In_436,In_1442);
nor U3580 (N_3580,In_1907,In_115);
or U3581 (N_3581,In_1633,In_1814);
nand U3582 (N_3582,In_214,In_213);
nor U3583 (N_3583,In_1577,In_1643);
nand U3584 (N_3584,In_584,In_1686);
or U3585 (N_3585,In_1758,In_1565);
and U3586 (N_3586,In_421,In_444);
nand U3587 (N_3587,In_1065,In_1473);
nand U3588 (N_3588,In_632,In_1251);
nand U3589 (N_3589,In_1777,In_53);
nand U3590 (N_3590,In_1907,In_1536);
and U3591 (N_3591,In_1528,In_1735);
and U3592 (N_3592,In_1565,In_748);
nand U3593 (N_3593,In_1634,In_986);
or U3594 (N_3594,In_481,In_720);
xnor U3595 (N_3595,In_1781,In_747);
or U3596 (N_3596,In_774,In_1514);
xor U3597 (N_3597,In_914,In_1528);
or U3598 (N_3598,In_1649,In_429);
or U3599 (N_3599,In_1794,In_182);
or U3600 (N_3600,In_741,In_5);
or U3601 (N_3601,In_1940,In_1268);
and U3602 (N_3602,In_1205,In_309);
xor U3603 (N_3603,In_30,In_1323);
nand U3604 (N_3604,In_1442,In_1508);
and U3605 (N_3605,In_107,In_527);
nor U3606 (N_3606,In_1645,In_54);
xor U3607 (N_3607,In_1770,In_1905);
nor U3608 (N_3608,In_721,In_260);
xnor U3609 (N_3609,In_231,In_1717);
nand U3610 (N_3610,In_107,In_359);
xnor U3611 (N_3611,In_1547,In_409);
or U3612 (N_3612,In_294,In_1695);
and U3613 (N_3613,In_1514,In_1568);
nand U3614 (N_3614,In_1871,In_794);
or U3615 (N_3615,In_86,In_304);
nand U3616 (N_3616,In_602,In_1054);
or U3617 (N_3617,In_166,In_268);
or U3618 (N_3618,In_495,In_633);
and U3619 (N_3619,In_1092,In_1003);
nand U3620 (N_3620,In_358,In_1);
nor U3621 (N_3621,In_95,In_1590);
or U3622 (N_3622,In_161,In_1237);
or U3623 (N_3623,In_155,In_1065);
nand U3624 (N_3624,In_1340,In_65);
or U3625 (N_3625,In_75,In_538);
or U3626 (N_3626,In_871,In_670);
and U3627 (N_3627,In_1777,In_555);
xor U3628 (N_3628,In_1602,In_309);
and U3629 (N_3629,In_817,In_399);
and U3630 (N_3630,In_144,In_1275);
and U3631 (N_3631,In_1317,In_1643);
or U3632 (N_3632,In_641,In_173);
and U3633 (N_3633,In_1372,In_1911);
and U3634 (N_3634,In_853,In_302);
nor U3635 (N_3635,In_462,In_1322);
or U3636 (N_3636,In_1573,In_833);
nor U3637 (N_3637,In_1690,In_1223);
nand U3638 (N_3638,In_486,In_451);
or U3639 (N_3639,In_225,In_1989);
or U3640 (N_3640,In_950,In_1318);
and U3641 (N_3641,In_264,In_1572);
nand U3642 (N_3642,In_311,In_1484);
or U3643 (N_3643,In_1923,In_996);
or U3644 (N_3644,In_1176,In_590);
and U3645 (N_3645,In_1883,In_988);
and U3646 (N_3646,In_1220,In_288);
nor U3647 (N_3647,In_543,In_924);
nand U3648 (N_3648,In_1417,In_965);
and U3649 (N_3649,In_672,In_1765);
or U3650 (N_3650,In_892,In_958);
and U3651 (N_3651,In_262,In_488);
and U3652 (N_3652,In_1503,In_1403);
xor U3653 (N_3653,In_1930,In_80);
or U3654 (N_3654,In_110,In_1835);
and U3655 (N_3655,In_61,In_1344);
and U3656 (N_3656,In_1613,In_1648);
xor U3657 (N_3657,In_496,In_1214);
or U3658 (N_3658,In_1355,In_1983);
and U3659 (N_3659,In_1193,In_1867);
nand U3660 (N_3660,In_434,In_1097);
nand U3661 (N_3661,In_1292,In_417);
and U3662 (N_3662,In_1997,In_549);
or U3663 (N_3663,In_1319,In_629);
or U3664 (N_3664,In_1663,In_802);
nand U3665 (N_3665,In_1655,In_963);
nand U3666 (N_3666,In_149,In_871);
or U3667 (N_3667,In_1581,In_623);
nor U3668 (N_3668,In_442,In_699);
nand U3669 (N_3669,In_59,In_1990);
or U3670 (N_3670,In_1475,In_368);
and U3671 (N_3671,In_515,In_946);
xor U3672 (N_3672,In_792,In_740);
xnor U3673 (N_3673,In_1271,In_99);
and U3674 (N_3674,In_1633,In_1154);
nor U3675 (N_3675,In_983,In_1707);
and U3676 (N_3676,In_886,In_1086);
and U3677 (N_3677,In_260,In_280);
and U3678 (N_3678,In_305,In_135);
nand U3679 (N_3679,In_411,In_690);
or U3680 (N_3680,In_374,In_1552);
and U3681 (N_3681,In_1926,In_1215);
nand U3682 (N_3682,In_1219,In_70);
xor U3683 (N_3683,In_569,In_321);
and U3684 (N_3684,In_602,In_1801);
or U3685 (N_3685,In_1411,In_480);
nand U3686 (N_3686,In_1823,In_1378);
or U3687 (N_3687,In_1161,In_951);
and U3688 (N_3688,In_250,In_643);
nor U3689 (N_3689,In_1862,In_1537);
or U3690 (N_3690,In_821,In_1473);
nand U3691 (N_3691,In_1139,In_1142);
nand U3692 (N_3692,In_1345,In_1217);
or U3693 (N_3693,In_1024,In_437);
or U3694 (N_3694,In_201,In_146);
nand U3695 (N_3695,In_1918,In_748);
or U3696 (N_3696,In_607,In_843);
and U3697 (N_3697,In_438,In_450);
nor U3698 (N_3698,In_524,In_1439);
nor U3699 (N_3699,In_47,In_1669);
nor U3700 (N_3700,In_566,In_235);
and U3701 (N_3701,In_1160,In_795);
nand U3702 (N_3702,In_662,In_254);
nor U3703 (N_3703,In_76,In_178);
and U3704 (N_3704,In_332,In_811);
nor U3705 (N_3705,In_1519,In_1121);
or U3706 (N_3706,In_1371,In_1521);
nor U3707 (N_3707,In_1044,In_1818);
and U3708 (N_3708,In_990,In_539);
and U3709 (N_3709,In_95,In_284);
xor U3710 (N_3710,In_568,In_1045);
and U3711 (N_3711,In_1447,In_451);
xnor U3712 (N_3712,In_1523,In_891);
nand U3713 (N_3713,In_1915,In_406);
nor U3714 (N_3714,In_831,In_1380);
or U3715 (N_3715,In_732,In_28);
and U3716 (N_3716,In_278,In_458);
nor U3717 (N_3717,In_31,In_1932);
nor U3718 (N_3718,In_1109,In_1500);
and U3719 (N_3719,In_1342,In_1585);
nor U3720 (N_3720,In_516,In_816);
or U3721 (N_3721,In_1034,In_754);
nand U3722 (N_3722,In_1449,In_1485);
xnor U3723 (N_3723,In_921,In_1871);
nor U3724 (N_3724,In_1402,In_1408);
nand U3725 (N_3725,In_901,In_314);
or U3726 (N_3726,In_100,In_767);
nor U3727 (N_3727,In_1468,In_860);
or U3728 (N_3728,In_990,In_20);
nand U3729 (N_3729,In_656,In_1230);
nor U3730 (N_3730,In_717,In_1292);
or U3731 (N_3731,In_547,In_104);
nand U3732 (N_3732,In_873,In_1156);
and U3733 (N_3733,In_1677,In_671);
and U3734 (N_3734,In_1704,In_1544);
or U3735 (N_3735,In_128,In_970);
nand U3736 (N_3736,In_1157,In_630);
nor U3737 (N_3737,In_1546,In_898);
and U3738 (N_3738,In_666,In_1341);
or U3739 (N_3739,In_1344,In_1670);
nand U3740 (N_3740,In_1346,In_1115);
and U3741 (N_3741,In_1832,In_860);
or U3742 (N_3742,In_1570,In_1448);
nand U3743 (N_3743,In_41,In_1933);
nor U3744 (N_3744,In_1638,In_1824);
and U3745 (N_3745,In_797,In_557);
nor U3746 (N_3746,In_982,In_496);
nand U3747 (N_3747,In_1340,In_1139);
and U3748 (N_3748,In_1723,In_1205);
or U3749 (N_3749,In_1606,In_135);
nor U3750 (N_3750,In_1871,In_1420);
nor U3751 (N_3751,In_1180,In_1226);
and U3752 (N_3752,In_1853,In_343);
and U3753 (N_3753,In_1103,In_1169);
and U3754 (N_3754,In_1646,In_863);
and U3755 (N_3755,In_697,In_1995);
or U3756 (N_3756,In_1788,In_1618);
and U3757 (N_3757,In_1298,In_484);
xnor U3758 (N_3758,In_1796,In_1890);
nand U3759 (N_3759,In_1122,In_1938);
or U3760 (N_3760,In_1415,In_748);
nor U3761 (N_3761,In_1306,In_543);
and U3762 (N_3762,In_1760,In_148);
xor U3763 (N_3763,In_668,In_521);
and U3764 (N_3764,In_1717,In_1064);
nand U3765 (N_3765,In_1187,In_1980);
and U3766 (N_3766,In_220,In_403);
nor U3767 (N_3767,In_1690,In_573);
xor U3768 (N_3768,In_1215,In_387);
and U3769 (N_3769,In_330,In_1240);
or U3770 (N_3770,In_70,In_354);
nand U3771 (N_3771,In_1288,In_1792);
nand U3772 (N_3772,In_1003,In_609);
nand U3773 (N_3773,In_1447,In_528);
or U3774 (N_3774,In_1125,In_1345);
or U3775 (N_3775,In_1300,In_36);
nor U3776 (N_3776,In_1549,In_1928);
and U3777 (N_3777,In_719,In_881);
nand U3778 (N_3778,In_234,In_885);
nand U3779 (N_3779,In_769,In_1437);
and U3780 (N_3780,In_1308,In_1961);
and U3781 (N_3781,In_565,In_795);
nand U3782 (N_3782,In_1860,In_1846);
nor U3783 (N_3783,In_1312,In_1564);
nor U3784 (N_3784,In_1420,In_881);
xnor U3785 (N_3785,In_1957,In_1201);
and U3786 (N_3786,In_786,In_1887);
and U3787 (N_3787,In_950,In_1981);
nand U3788 (N_3788,In_305,In_698);
or U3789 (N_3789,In_1089,In_1314);
xnor U3790 (N_3790,In_774,In_720);
nor U3791 (N_3791,In_1049,In_1414);
or U3792 (N_3792,In_34,In_149);
and U3793 (N_3793,In_1611,In_1108);
nor U3794 (N_3794,In_189,In_194);
nand U3795 (N_3795,In_1486,In_1795);
or U3796 (N_3796,In_809,In_196);
or U3797 (N_3797,In_1544,In_1079);
nor U3798 (N_3798,In_275,In_606);
nand U3799 (N_3799,In_1764,In_1335);
nor U3800 (N_3800,In_113,In_988);
nor U3801 (N_3801,In_1837,In_1301);
nor U3802 (N_3802,In_1306,In_662);
and U3803 (N_3803,In_507,In_217);
xnor U3804 (N_3804,In_171,In_1371);
nand U3805 (N_3805,In_1355,In_1409);
nor U3806 (N_3806,In_865,In_1861);
or U3807 (N_3807,In_471,In_1677);
or U3808 (N_3808,In_4,In_1330);
nor U3809 (N_3809,In_1869,In_110);
and U3810 (N_3810,In_1129,In_662);
nand U3811 (N_3811,In_1318,In_1645);
nor U3812 (N_3812,In_509,In_588);
nand U3813 (N_3813,In_1469,In_116);
and U3814 (N_3814,In_1743,In_1153);
or U3815 (N_3815,In_1303,In_1312);
or U3816 (N_3816,In_1318,In_217);
nand U3817 (N_3817,In_1017,In_1561);
and U3818 (N_3818,In_233,In_695);
xnor U3819 (N_3819,In_1157,In_1252);
xor U3820 (N_3820,In_595,In_735);
and U3821 (N_3821,In_1319,In_198);
or U3822 (N_3822,In_1586,In_1527);
nor U3823 (N_3823,In_616,In_1135);
and U3824 (N_3824,In_1317,In_673);
xnor U3825 (N_3825,In_1459,In_1499);
nand U3826 (N_3826,In_231,In_367);
nand U3827 (N_3827,In_1542,In_912);
and U3828 (N_3828,In_406,In_73);
nand U3829 (N_3829,In_1110,In_1576);
or U3830 (N_3830,In_1924,In_1857);
nand U3831 (N_3831,In_1366,In_1668);
xnor U3832 (N_3832,In_1599,In_808);
nor U3833 (N_3833,In_1005,In_1732);
nor U3834 (N_3834,In_1036,In_543);
or U3835 (N_3835,In_25,In_367);
nor U3836 (N_3836,In_1290,In_312);
and U3837 (N_3837,In_1177,In_1123);
xor U3838 (N_3838,In_1021,In_63);
and U3839 (N_3839,In_1384,In_1458);
nor U3840 (N_3840,In_1588,In_1690);
or U3841 (N_3841,In_716,In_1092);
or U3842 (N_3842,In_695,In_1070);
nand U3843 (N_3843,In_741,In_1349);
nand U3844 (N_3844,In_302,In_339);
nand U3845 (N_3845,In_969,In_334);
and U3846 (N_3846,In_1032,In_647);
nor U3847 (N_3847,In_1244,In_1949);
nand U3848 (N_3848,In_1484,In_1390);
or U3849 (N_3849,In_1928,In_900);
nor U3850 (N_3850,In_465,In_566);
nor U3851 (N_3851,In_1542,In_142);
and U3852 (N_3852,In_410,In_1472);
and U3853 (N_3853,In_1842,In_1225);
nor U3854 (N_3854,In_1623,In_1549);
or U3855 (N_3855,In_533,In_546);
or U3856 (N_3856,In_1013,In_1779);
nor U3857 (N_3857,In_1015,In_1699);
nor U3858 (N_3858,In_566,In_1374);
nand U3859 (N_3859,In_1862,In_1474);
nor U3860 (N_3860,In_779,In_1168);
and U3861 (N_3861,In_1725,In_1648);
and U3862 (N_3862,In_193,In_566);
and U3863 (N_3863,In_480,In_1928);
nor U3864 (N_3864,In_1409,In_1328);
or U3865 (N_3865,In_576,In_1948);
nand U3866 (N_3866,In_875,In_1102);
or U3867 (N_3867,In_1301,In_1387);
nor U3868 (N_3868,In_1911,In_364);
or U3869 (N_3869,In_337,In_1797);
and U3870 (N_3870,In_1319,In_1605);
or U3871 (N_3871,In_887,In_1852);
nand U3872 (N_3872,In_1093,In_415);
or U3873 (N_3873,In_453,In_1661);
and U3874 (N_3874,In_1325,In_1331);
or U3875 (N_3875,In_144,In_1188);
or U3876 (N_3876,In_1943,In_1689);
or U3877 (N_3877,In_1789,In_1542);
or U3878 (N_3878,In_1321,In_1622);
or U3879 (N_3879,In_904,In_1647);
and U3880 (N_3880,In_718,In_1910);
nor U3881 (N_3881,In_1797,In_1933);
nor U3882 (N_3882,In_1117,In_1689);
and U3883 (N_3883,In_1883,In_856);
nor U3884 (N_3884,In_518,In_110);
xor U3885 (N_3885,In_1105,In_1456);
nand U3886 (N_3886,In_1221,In_241);
and U3887 (N_3887,In_574,In_1352);
nand U3888 (N_3888,In_1284,In_685);
nor U3889 (N_3889,In_888,In_1209);
nor U3890 (N_3890,In_947,In_1674);
nor U3891 (N_3891,In_540,In_1009);
or U3892 (N_3892,In_189,In_575);
and U3893 (N_3893,In_487,In_858);
or U3894 (N_3894,In_278,In_143);
and U3895 (N_3895,In_618,In_438);
and U3896 (N_3896,In_1197,In_1000);
and U3897 (N_3897,In_259,In_1115);
and U3898 (N_3898,In_1301,In_1142);
and U3899 (N_3899,In_1507,In_1597);
nand U3900 (N_3900,In_1739,In_202);
nand U3901 (N_3901,In_1057,In_1705);
nor U3902 (N_3902,In_785,In_1561);
nor U3903 (N_3903,In_1052,In_174);
and U3904 (N_3904,In_348,In_630);
and U3905 (N_3905,In_1037,In_1446);
and U3906 (N_3906,In_1218,In_892);
or U3907 (N_3907,In_1998,In_179);
nand U3908 (N_3908,In_103,In_1798);
and U3909 (N_3909,In_1744,In_311);
or U3910 (N_3910,In_42,In_1297);
xnor U3911 (N_3911,In_783,In_1102);
nand U3912 (N_3912,In_1727,In_337);
and U3913 (N_3913,In_919,In_792);
or U3914 (N_3914,In_1269,In_795);
nor U3915 (N_3915,In_151,In_1204);
and U3916 (N_3916,In_101,In_572);
nor U3917 (N_3917,In_1758,In_1115);
nand U3918 (N_3918,In_49,In_1162);
nand U3919 (N_3919,In_37,In_1346);
and U3920 (N_3920,In_1071,In_134);
xnor U3921 (N_3921,In_1614,In_975);
nor U3922 (N_3922,In_741,In_1611);
nor U3923 (N_3923,In_1269,In_69);
or U3924 (N_3924,In_1700,In_492);
or U3925 (N_3925,In_371,In_110);
and U3926 (N_3926,In_1425,In_1897);
and U3927 (N_3927,In_878,In_1587);
and U3928 (N_3928,In_1054,In_481);
nand U3929 (N_3929,In_483,In_1067);
nand U3930 (N_3930,In_1402,In_1927);
xor U3931 (N_3931,In_760,In_1180);
or U3932 (N_3932,In_597,In_818);
and U3933 (N_3933,In_498,In_1369);
or U3934 (N_3934,In_1201,In_1718);
nor U3935 (N_3935,In_253,In_355);
xnor U3936 (N_3936,In_567,In_346);
or U3937 (N_3937,In_743,In_1777);
xnor U3938 (N_3938,In_1501,In_1485);
nand U3939 (N_3939,In_1223,In_1797);
nor U3940 (N_3940,In_1422,In_37);
nor U3941 (N_3941,In_963,In_972);
nand U3942 (N_3942,In_1783,In_1950);
nor U3943 (N_3943,In_397,In_576);
or U3944 (N_3944,In_1654,In_381);
and U3945 (N_3945,In_278,In_1348);
nor U3946 (N_3946,In_934,In_824);
or U3947 (N_3947,In_537,In_444);
and U3948 (N_3948,In_821,In_1189);
nand U3949 (N_3949,In_1183,In_1158);
and U3950 (N_3950,In_310,In_479);
and U3951 (N_3951,In_1508,In_141);
nor U3952 (N_3952,In_9,In_904);
or U3953 (N_3953,In_1729,In_1584);
nand U3954 (N_3954,In_896,In_1808);
nor U3955 (N_3955,In_176,In_1134);
and U3956 (N_3956,In_274,In_1751);
and U3957 (N_3957,In_1462,In_1802);
xor U3958 (N_3958,In_317,In_1316);
nor U3959 (N_3959,In_1210,In_1340);
or U3960 (N_3960,In_1211,In_1779);
and U3961 (N_3961,In_181,In_724);
nor U3962 (N_3962,In_701,In_1508);
and U3963 (N_3963,In_979,In_1910);
nand U3964 (N_3964,In_1696,In_644);
or U3965 (N_3965,In_428,In_1006);
and U3966 (N_3966,In_1038,In_41);
xnor U3967 (N_3967,In_760,In_6);
or U3968 (N_3968,In_634,In_1983);
nor U3969 (N_3969,In_1784,In_1258);
xnor U3970 (N_3970,In_1311,In_1900);
nand U3971 (N_3971,In_1683,In_1862);
and U3972 (N_3972,In_715,In_1608);
nor U3973 (N_3973,In_1184,In_1162);
and U3974 (N_3974,In_1679,In_1230);
or U3975 (N_3975,In_1884,In_174);
and U3976 (N_3976,In_1985,In_301);
and U3977 (N_3977,In_869,In_1328);
or U3978 (N_3978,In_751,In_1944);
or U3979 (N_3979,In_573,In_1492);
nand U3980 (N_3980,In_1055,In_1003);
nand U3981 (N_3981,In_447,In_1200);
and U3982 (N_3982,In_10,In_1786);
xnor U3983 (N_3983,In_474,In_1136);
or U3984 (N_3984,In_598,In_405);
nand U3985 (N_3985,In_180,In_1603);
nand U3986 (N_3986,In_1005,In_128);
or U3987 (N_3987,In_150,In_983);
or U3988 (N_3988,In_861,In_261);
xor U3989 (N_3989,In_586,In_913);
and U3990 (N_3990,In_805,In_201);
nor U3991 (N_3991,In_246,In_1748);
and U3992 (N_3992,In_1849,In_32);
nand U3993 (N_3993,In_1095,In_958);
or U3994 (N_3994,In_139,In_1218);
and U3995 (N_3995,In_235,In_246);
xor U3996 (N_3996,In_1066,In_329);
and U3997 (N_3997,In_920,In_596);
and U3998 (N_3998,In_1237,In_971);
nand U3999 (N_3999,In_1157,In_714);
xor U4000 (N_4000,In_1633,In_1229);
and U4001 (N_4001,In_1945,In_391);
nor U4002 (N_4002,In_286,In_311);
nand U4003 (N_4003,In_1356,In_37);
or U4004 (N_4004,In_439,In_1182);
or U4005 (N_4005,In_1072,In_1691);
nor U4006 (N_4006,In_28,In_111);
nor U4007 (N_4007,In_694,In_982);
or U4008 (N_4008,In_1710,In_502);
nand U4009 (N_4009,In_698,In_1492);
or U4010 (N_4010,In_133,In_540);
nand U4011 (N_4011,In_220,In_1605);
nand U4012 (N_4012,In_211,In_1581);
or U4013 (N_4013,In_1643,In_235);
nor U4014 (N_4014,In_675,In_1646);
or U4015 (N_4015,In_533,In_731);
nand U4016 (N_4016,In_530,In_1919);
xor U4017 (N_4017,In_1682,In_1154);
or U4018 (N_4018,In_193,In_1268);
nand U4019 (N_4019,In_415,In_468);
and U4020 (N_4020,In_675,In_251);
and U4021 (N_4021,In_167,In_1802);
nand U4022 (N_4022,In_513,In_895);
nor U4023 (N_4023,In_1798,In_1444);
and U4024 (N_4024,In_1346,In_301);
and U4025 (N_4025,In_401,In_1545);
or U4026 (N_4026,In_476,In_138);
nor U4027 (N_4027,In_1301,In_346);
nand U4028 (N_4028,In_953,In_244);
nand U4029 (N_4029,In_225,In_870);
nand U4030 (N_4030,In_1981,In_1632);
or U4031 (N_4031,In_1810,In_1455);
xor U4032 (N_4032,In_1696,In_1576);
xnor U4033 (N_4033,In_352,In_931);
xnor U4034 (N_4034,In_581,In_323);
or U4035 (N_4035,In_997,In_1863);
nor U4036 (N_4036,In_803,In_1416);
nand U4037 (N_4037,In_334,In_953);
nor U4038 (N_4038,In_114,In_883);
nor U4039 (N_4039,In_276,In_114);
or U4040 (N_4040,In_1062,In_1917);
or U4041 (N_4041,In_374,In_1450);
nor U4042 (N_4042,In_715,In_854);
and U4043 (N_4043,In_231,In_575);
or U4044 (N_4044,In_1229,In_174);
and U4045 (N_4045,In_222,In_305);
and U4046 (N_4046,In_1007,In_1110);
nor U4047 (N_4047,In_190,In_1660);
or U4048 (N_4048,In_1058,In_489);
or U4049 (N_4049,In_186,In_1034);
and U4050 (N_4050,In_142,In_1104);
nand U4051 (N_4051,In_363,In_555);
xor U4052 (N_4052,In_530,In_130);
or U4053 (N_4053,In_660,In_638);
nor U4054 (N_4054,In_822,In_850);
nor U4055 (N_4055,In_1481,In_1422);
nand U4056 (N_4056,In_994,In_1369);
nor U4057 (N_4057,In_571,In_97);
nand U4058 (N_4058,In_790,In_1182);
and U4059 (N_4059,In_134,In_156);
or U4060 (N_4060,In_82,In_1277);
and U4061 (N_4061,In_661,In_733);
nand U4062 (N_4062,In_1895,In_559);
nand U4063 (N_4063,In_962,In_1215);
nand U4064 (N_4064,In_1827,In_1119);
or U4065 (N_4065,In_855,In_431);
nand U4066 (N_4066,In_1264,In_651);
or U4067 (N_4067,In_18,In_1609);
nor U4068 (N_4068,In_933,In_556);
and U4069 (N_4069,In_624,In_636);
nor U4070 (N_4070,In_1019,In_1631);
or U4071 (N_4071,In_1934,In_382);
nor U4072 (N_4072,In_349,In_1164);
nand U4073 (N_4073,In_1005,In_1434);
and U4074 (N_4074,In_1107,In_30);
or U4075 (N_4075,In_1759,In_1525);
nand U4076 (N_4076,In_269,In_1103);
or U4077 (N_4077,In_1437,In_157);
nor U4078 (N_4078,In_32,In_720);
nand U4079 (N_4079,In_997,In_1211);
nor U4080 (N_4080,In_370,In_1223);
xor U4081 (N_4081,In_1581,In_1849);
nor U4082 (N_4082,In_423,In_564);
or U4083 (N_4083,In_1043,In_1228);
and U4084 (N_4084,In_631,In_991);
and U4085 (N_4085,In_1160,In_1822);
nor U4086 (N_4086,In_691,In_1268);
or U4087 (N_4087,In_1328,In_721);
nand U4088 (N_4088,In_770,In_887);
and U4089 (N_4089,In_719,In_1502);
and U4090 (N_4090,In_313,In_1207);
nor U4091 (N_4091,In_661,In_400);
xor U4092 (N_4092,In_1002,In_663);
and U4093 (N_4093,In_1351,In_1868);
nor U4094 (N_4094,In_664,In_694);
and U4095 (N_4095,In_1712,In_1564);
nor U4096 (N_4096,In_1260,In_1335);
or U4097 (N_4097,In_1308,In_686);
nor U4098 (N_4098,In_756,In_961);
or U4099 (N_4099,In_1160,In_737);
or U4100 (N_4100,In_988,In_1671);
nor U4101 (N_4101,In_1142,In_1929);
and U4102 (N_4102,In_1645,In_560);
and U4103 (N_4103,In_1259,In_886);
and U4104 (N_4104,In_1116,In_1452);
nand U4105 (N_4105,In_1542,In_130);
and U4106 (N_4106,In_784,In_496);
nand U4107 (N_4107,In_263,In_941);
or U4108 (N_4108,In_33,In_613);
or U4109 (N_4109,In_114,In_1645);
nand U4110 (N_4110,In_865,In_1273);
and U4111 (N_4111,In_1186,In_1867);
or U4112 (N_4112,In_259,In_1452);
nor U4113 (N_4113,In_132,In_534);
and U4114 (N_4114,In_1419,In_73);
or U4115 (N_4115,In_918,In_1508);
or U4116 (N_4116,In_593,In_1031);
or U4117 (N_4117,In_1266,In_1429);
nor U4118 (N_4118,In_1682,In_1343);
xor U4119 (N_4119,In_1318,In_1451);
or U4120 (N_4120,In_1753,In_182);
and U4121 (N_4121,In_1448,In_414);
or U4122 (N_4122,In_773,In_1924);
and U4123 (N_4123,In_358,In_867);
and U4124 (N_4124,In_145,In_622);
nor U4125 (N_4125,In_131,In_1347);
nor U4126 (N_4126,In_742,In_71);
and U4127 (N_4127,In_492,In_1916);
or U4128 (N_4128,In_636,In_802);
nor U4129 (N_4129,In_703,In_494);
xor U4130 (N_4130,In_216,In_1798);
nand U4131 (N_4131,In_921,In_457);
and U4132 (N_4132,In_213,In_1664);
nand U4133 (N_4133,In_1860,In_402);
or U4134 (N_4134,In_1356,In_783);
and U4135 (N_4135,In_393,In_1808);
nand U4136 (N_4136,In_1468,In_667);
and U4137 (N_4137,In_182,In_1493);
nand U4138 (N_4138,In_158,In_1741);
and U4139 (N_4139,In_527,In_216);
xor U4140 (N_4140,In_854,In_683);
xor U4141 (N_4141,In_1974,In_193);
xnor U4142 (N_4142,In_1776,In_1356);
and U4143 (N_4143,In_1697,In_1835);
nor U4144 (N_4144,In_1926,In_1300);
xor U4145 (N_4145,In_1946,In_304);
xnor U4146 (N_4146,In_1044,In_1546);
nor U4147 (N_4147,In_1013,In_1403);
and U4148 (N_4148,In_1551,In_342);
or U4149 (N_4149,In_1619,In_1518);
and U4150 (N_4150,In_514,In_1471);
and U4151 (N_4151,In_1431,In_139);
or U4152 (N_4152,In_8,In_756);
nand U4153 (N_4153,In_542,In_478);
nand U4154 (N_4154,In_1181,In_1124);
and U4155 (N_4155,In_198,In_829);
xnor U4156 (N_4156,In_1341,In_1681);
nor U4157 (N_4157,In_455,In_812);
nor U4158 (N_4158,In_644,In_495);
or U4159 (N_4159,In_900,In_556);
nand U4160 (N_4160,In_420,In_1414);
nand U4161 (N_4161,In_800,In_576);
and U4162 (N_4162,In_527,In_499);
or U4163 (N_4163,In_1763,In_656);
nand U4164 (N_4164,In_1395,In_623);
xnor U4165 (N_4165,In_1857,In_1534);
or U4166 (N_4166,In_1878,In_1545);
and U4167 (N_4167,In_638,In_1983);
or U4168 (N_4168,In_1245,In_1760);
or U4169 (N_4169,In_0,In_1237);
and U4170 (N_4170,In_1270,In_266);
nor U4171 (N_4171,In_1989,In_1020);
or U4172 (N_4172,In_87,In_359);
nand U4173 (N_4173,In_909,In_172);
nor U4174 (N_4174,In_780,In_1649);
and U4175 (N_4175,In_424,In_1570);
and U4176 (N_4176,In_1172,In_929);
or U4177 (N_4177,In_1429,In_573);
and U4178 (N_4178,In_1827,In_1310);
nand U4179 (N_4179,In_112,In_1874);
and U4180 (N_4180,In_876,In_720);
nand U4181 (N_4181,In_1222,In_144);
and U4182 (N_4182,In_1242,In_1265);
nand U4183 (N_4183,In_1977,In_1111);
nand U4184 (N_4184,In_616,In_1188);
or U4185 (N_4185,In_929,In_282);
nor U4186 (N_4186,In_1475,In_1762);
nand U4187 (N_4187,In_1814,In_1025);
or U4188 (N_4188,In_285,In_608);
nor U4189 (N_4189,In_967,In_1508);
and U4190 (N_4190,In_70,In_796);
nand U4191 (N_4191,In_578,In_828);
nand U4192 (N_4192,In_798,In_346);
nand U4193 (N_4193,In_1817,In_1913);
or U4194 (N_4194,In_1470,In_299);
nor U4195 (N_4195,In_198,In_1277);
nor U4196 (N_4196,In_1459,In_405);
nand U4197 (N_4197,In_471,In_1494);
nor U4198 (N_4198,In_1072,In_1168);
nand U4199 (N_4199,In_672,In_1311);
or U4200 (N_4200,In_994,In_366);
or U4201 (N_4201,In_965,In_31);
nor U4202 (N_4202,In_1407,In_411);
nand U4203 (N_4203,In_102,In_901);
and U4204 (N_4204,In_1142,In_107);
nor U4205 (N_4205,In_1512,In_982);
nand U4206 (N_4206,In_1604,In_1506);
or U4207 (N_4207,In_1095,In_123);
nor U4208 (N_4208,In_1372,In_791);
or U4209 (N_4209,In_1790,In_1830);
and U4210 (N_4210,In_455,In_817);
and U4211 (N_4211,In_62,In_995);
and U4212 (N_4212,In_1501,In_132);
nor U4213 (N_4213,In_893,In_1221);
and U4214 (N_4214,In_1206,In_157);
nand U4215 (N_4215,In_1444,In_256);
or U4216 (N_4216,In_1793,In_1918);
xnor U4217 (N_4217,In_321,In_1658);
and U4218 (N_4218,In_210,In_1452);
nand U4219 (N_4219,In_1875,In_1490);
or U4220 (N_4220,In_772,In_629);
xnor U4221 (N_4221,In_123,In_1872);
and U4222 (N_4222,In_1601,In_1625);
or U4223 (N_4223,In_434,In_339);
or U4224 (N_4224,In_598,In_30);
xnor U4225 (N_4225,In_1623,In_757);
or U4226 (N_4226,In_919,In_1040);
and U4227 (N_4227,In_501,In_1382);
nand U4228 (N_4228,In_1771,In_551);
nand U4229 (N_4229,In_412,In_1962);
nor U4230 (N_4230,In_1203,In_1841);
nand U4231 (N_4231,In_1007,In_1598);
nor U4232 (N_4232,In_1051,In_683);
or U4233 (N_4233,In_1949,In_1002);
and U4234 (N_4234,In_608,In_1881);
and U4235 (N_4235,In_1596,In_115);
nand U4236 (N_4236,In_1325,In_747);
nand U4237 (N_4237,In_1989,In_1431);
or U4238 (N_4238,In_1631,In_1911);
or U4239 (N_4239,In_839,In_1828);
nand U4240 (N_4240,In_1753,In_1969);
nand U4241 (N_4241,In_1627,In_541);
and U4242 (N_4242,In_1069,In_140);
xnor U4243 (N_4243,In_1122,In_1415);
or U4244 (N_4244,In_1619,In_463);
nand U4245 (N_4245,In_1335,In_841);
and U4246 (N_4246,In_434,In_1654);
and U4247 (N_4247,In_823,In_1004);
nand U4248 (N_4248,In_1985,In_496);
nor U4249 (N_4249,In_145,In_424);
xnor U4250 (N_4250,In_1990,In_856);
nand U4251 (N_4251,In_954,In_733);
and U4252 (N_4252,In_1696,In_99);
nor U4253 (N_4253,In_149,In_1284);
or U4254 (N_4254,In_726,In_471);
and U4255 (N_4255,In_1752,In_1994);
or U4256 (N_4256,In_447,In_1558);
nor U4257 (N_4257,In_443,In_986);
and U4258 (N_4258,In_1200,In_1914);
or U4259 (N_4259,In_1042,In_1916);
nor U4260 (N_4260,In_848,In_194);
and U4261 (N_4261,In_645,In_319);
nor U4262 (N_4262,In_76,In_715);
nand U4263 (N_4263,In_1433,In_426);
nor U4264 (N_4264,In_90,In_235);
xnor U4265 (N_4265,In_987,In_1538);
and U4266 (N_4266,In_822,In_1806);
nand U4267 (N_4267,In_266,In_1103);
and U4268 (N_4268,In_1612,In_1467);
and U4269 (N_4269,In_829,In_1530);
or U4270 (N_4270,In_1672,In_608);
or U4271 (N_4271,In_1013,In_1021);
nor U4272 (N_4272,In_1033,In_1076);
nor U4273 (N_4273,In_215,In_1838);
and U4274 (N_4274,In_799,In_1740);
nor U4275 (N_4275,In_1930,In_1914);
nor U4276 (N_4276,In_934,In_472);
xor U4277 (N_4277,In_708,In_363);
nor U4278 (N_4278,In_1524,In_1720);
and U4279 (N_4279,In_893,In_1633);
xor U4280 (N_4280,In_813,In_1580);
xor U4281 (N_4281,In_1495,In_101);
xnor U4282 (N_4282,In_369,In_1938);
or U4283 (N_4283,In_1158,In_1745);
and U4284 (N_4284,In_514,In_1516);
and U4285 (N_4285,In_221,In_1853);
or U4286 (N_4286,In_457,In_1195);
or U4287 (N_4287,In_1368,In_1567);
nor U4288 (N_4288,In_1769,In_335);
nand U4289 (N_4289,In_1630,In_357);
nand U4290 (N_4290,In_1056,In_752);
nor U4291 (N_4291,In_1019,In_597);
xnor U4292 (N_4292,In_1534,In_1030);
xor U4293 (N_4293,In_1568,In_1608);
or U4294 (N_4294,In_1439,In_1624);
and U4295 (N_4295,In_819,In_1966);
or U4296 (N_4296,In_1190,In_339);
nor U4297 (N_4297,In_330,In_1626);
and U4298 (N_4298,In_1599,In_566);
or U4299 (N_4299,In_1674,In_881);
nand U4300 (N_4300,In_1281,In_1024);
and U4301 (N_4301,In_1549,In_955);
nand U4302 (N_4302,In_434,In_1513);
or U4303 (N_4303,In_1127,In_1578);
nand U4304 (N_4304,In_1590,In_410);
and U4305 (N_4305,In_298,In_1164);
or U4306 (N_4306,In_1168,In_347);
and U4307 (N_4307,In_1176,In_1851);
nand U4308 (N_4308,In_1088,In_1330);
or U4309 (N_4309,In_1680,In_204);
nand U4310 (N_4310,In_407,In_1762);
nor U4311 (N_4311,In_1223,In_1115);
nor U4312 (N_4312,In_216,In_1215);
nand U4313 (N_4313,In_1111,In_230);
nor U4314 (N_4314,In_940,In_1891);
or U4315 (N_4315,In_729,In_1924);
xor U4316 (N_4316,In_202,In_1309);
and U4317 (N_4317,In_1141,In_1927);
nand U4318 (N_4318,In_62,In_1609);
nand U4319 (N_4319,In_585,In_1519);
nand U4320 (N_4320,In_1048,In_834);
and U4321 (N_4321,In_827,In_864);
and U4322 (N_4322,In_1895,In_382);
and U4323 (N_4323,In_1769,In_1593);
nor U4324 (N_4324,In_750,In_212);
and U4325 (N_4325,In_49,In_1613);
or U4326 (N_4326,In_1880,In_411);
nor U4327 (N_4327,In_1366,In_779);
or U4328 (N_4328,In_168,In_839);
and U4329 (N_4329,In_377,In_1135);
nor U4330 (N_4330,In_1343,In_1980);
xnor U4331 (N_4331,In_1606,In_1421);
nand U4332 (N_4332,In_994,In_234);
or U4333 (N_4333,In_840,In_1973);
or U4334 (N_4334,In_1747,In_1966);
or U4335 (N_4335,In_390,In_291);
nand U4336 (N_4336,In_1374,In_1305);
nor U4337 (N_4337,In_393,In_1653);
or U4338 (N_4338,In_1947,In_1650);
or U4339 (N_4339,In_776,In_1796);
xor U4340 (N_4340,In_252,In_1626);
and U4341 (N_4341,In_658,In_1353);
nor U4342 (N_4342,In_1619,In_142);
nand U4343 (N_4343,In_1290,In_103);
nand U4344 (N_4344,In_780,In_242);
and U4345 (N_4345,In_1002,In_1921);
nor U4346 (N_4346,In_1523,In_1966);
or U4347 (N_4347,In_1883,In_1700);
or U4348 (N_4348,In_1030,In_1706);
xor U4349 (N_4349,In_1770,In_1267);
nand U4350 (N_4350,In_956,In_1308);
nand U4351 (N_4351,In_1988,In_216);
and U4352 (N_4352,In_1954,In_1712);
nand U4353 (N_4353,In_1089,In_21);
nand U4354 (N_4354,In_853,In_261);
nand U4355 (N_4355,In_1119,In_207);
nor U4356 (N_4356,In_754,In_635);
and U4357 (N_4357,In_805,In_1995);
or U4358 (N_4358,In_431,In_698);
xnor U4359 (N_4359,In_1427,In_333);
nand U4360 (N_4360,In_307,In_1656);
nor U4361 (N_4361,In_124,In_1097);
nor U4362 (N_4362,In_1053,In_369);
or U4363 (N_4363,In_1839,In_1189);
nand U4364 (N_4364,In_60,In_1247);
nor U4365 (N_4365,In_486,In_973);
or U4366 (N_4366,In_1071,In_1583);
nand U4367 (N_4367,In_1162,In_639);
nand U4368 (N_4368,In_1069,In_557);
nor U4369 (N_4369,In_75,In_1138);
and U4370 (N_4370,In_1636,In_1019);
nand U4371 (N_4371,In_1497,In_723);
or U4372 (N_4372,In_1560,In_1258);
nand U4373 (N_4373,In_332,In_87);
nor U4374 (N_4374,In_223,In_1498);
or U4375 (N_4375,In_259,In_1238);
xor U4376 (N_4376,In_828,In_872);
nor U4377 (N_4377,In_1237,In_140);
or U4378 (N_4378,In_1595,In_1239);
and U4379 (N_4379,In_1254,In_718);
or U4380 (N_4380,In_81,In_1245);
nand U4381 (N_4381,In_1152,In_1972);
nand U4382 (N_4382,In_1364,In_116);
nand U4383 (N_4383,In_1846,In_1140);
or U4384 (N_4384,In_977,In_1405);
or U4385 (N_4385,In_1719,In_1489);
nor U4386 (N_4386,In_1815,In_1011);
xnor U4387 (N_4387,In_1012,In_1030);
nor U4388 (N_4388,In_437,In_595);
and U4389 (N_4389,In_1337,In_430);
and U4390 (N_4390,In_1284,In_774);
or U4391 (N_4391,In_1516,In_989);
nand U4392 (N_4392,In_692,In_1472);
nand U4393 (N_4393,In_673,In_1101);
and U4394 (N_4394,In_372,In_1250);
and U4395 (N_4395,In_220,In_122);
or U4396 (N_4396,In_417,In_1950);
nand U4397 (N_4397,In_404,In_337);
and U4398 (N_4398,In_222,In_1396);
nand U4399 (N_4399,In_1711,In_1484);
or U4400 (N_4400,In_404,In_1420);
nand U4401 (N_4401,In_1309,In_734);
or U4402 (N_4402,In_1222,In_479);
and U4403 (N_4403,In_1129,In_600);
xnor U4404 (N_4404,In_712,In_694);
nand U4405 (N_4405,In_1093,In_488);
xnor U4406 (N_4406,In_809,In_714);
and U4407 (N_4407,In_1473,In_1068);
and U4408 (N_4408,In_83,In_1213);
and U4409 (N_4409,In_699,In_1578);
and U4410 (N_4410,In_1672,In_1035);
nor U4411 (N_4411,In_1608,In_94);
and U4412 (N_4412,In_85,In_1711);
nand U4413 (N_4413,In_1448,In_306);
xnor U4414 (N_4414,In_407,In_392);
and U4415 (N_4415,In_124,In_1975);
and U4416 (N_4416,In_353,In_1781);
or U4417 (N_4417,In_641,In_1908);
nor U4418 (N_4418,In_1302,In_282);
and U4419 (N_4419,In_680,In_1316);
and U4420 (N_4420,In_1057,In_1233);
or U4421 (N_4421,In_695,In_787);
nor U4422 (N_4422,In_318,In_403);
nor U4423 (N_4423,In_1002,In_360);
nor U4424 (N_4424,In_1722,In_1137);
xor U4425 (N_4425,In_1729,In_1884);
and U4426 (N_4426,In_1428,In_1908);
nor U4427 (N_4427,In_213,In_538);
nor U4428 (N_4428,In_1739,In_1914);
nand U4429 (N_4429,In_629,In_1619);
and U4430 (N_4430,In_1541,In_1251);
and U4431 (N_4431,In_823,In_534);
and U4432 (N_4432,In_1298,In_1016);
nand U4433 (N_4433,In_200,In_1888);
nor U4434 (N_4434,In_970,In_1460);
and U4435 (N_4435,In_1424,In_1607);
and U4436 (N_4436,In_313,In_1706);
nand U4437 (N_4437,In_1261,In_1488);
or U4438 (N_4438,In_1331,In_795);
xnor U4439 (N_4439,In_1288,In_1240);
xor U4440 (N_4440,In_1935,In_1379);
and U4441 (N_4441,In_1611,In_997);
xor U4442 (N_4442,In_1092,In_190);
or U4443 (N_4443,In_1395,In_596);
nand U4444 (N_4444,In_950,In_193);
nand U4445 (N_4445,In_1197,In_423);
or U4446 (N_4446,In_992,In_1521);
nor U4447 (N_4447,In_700,In_1655);
nor U4448 (N_4448,In_607,In_1635);
nor U4449 (N_4449,In_1588,In_1004);
xnor U4450 (N_4450,In_1439,In_909);
nand U4451 (N_4451,In_706,In_1903);
and U4452 (N_4452,In_1669,In_1086);
nor U4453 (N_4453,In_583,In_1583);
or U4454 (N_4454,In_1129,In_290);
nor U4455 (N_4455,In_1429,In_1691);
and U4456 (N_4456,In_964,In_1733);
nand U4457 (N_4457,In_1587,In_1896);
nand U4458 (N_4458,In_102,In_1619);
nand U4459 (N_4459,In_1051,In_1180);
nor U4460 (N_4460,In_1452,In_1362);
and U4461 (N_4461,In_1797,In_748);
nand U4462 (N_4462,In_789,In_66);
nor U4463 (N_4463,In_389,In_91);
xor U4464 (N_4464,In_135,In_1320);
nor U4465 (N_4465,In_1970,In_1742);
and U4466 (N_4466,In_856,In_321);
nor U4467 (N_4467,In_419,In_893);
or U4468 (N_4468,In_1836,In_688);
nand U4469 (N_4469,In_1987,In_335);
nand U4470 (N_4470,In_1180,In_881);
nand U4471 (N_4471,In_1499,In_1823);
xnor U4472 (N_4472,In_1278,In_445);
or U4473 (N_4473,In_327,In_163);
nor U4474 (N_4474,In_1681,In_1421);
and U4475 (N_4475,In_1996,In_621);
nand U4476 (N_4476,In_1176,In_1790);
and U4477 (N_4477,In_1206,In_616);
nand U4478 (N_4478,In_1040,In_978);
or U4479 (N_4479,In_1537,In_720);
nand U4480 (N_4480,In_428,In_1209);
nand U4481 (N_4481,In_770,In_814);
nand U4482 (N_4482,In_1575,In_1857);
or U4483 (N_4483,In_327,In_301);
or U4484 (N_4484,In_517,In_87);
nor U4485 (N_4485,In_1070,In_789);
and U4486 (N_4486,In_393,In_2);
and U4487 (N_4487,In_923,In_371);
nand U4488 (N_4488,In_1255,In_965);
or U4489 (N_4489,In_432,In_759);
nand U4490 (N_4490,In_1301,In_1342);
or U4491 (N_4491,In_1098,In_1976);
nand U4492 (N_4492,In_10,In_1912);
and U4493 (N_4493,In_82,In_1600);
nand U4494 (N_4494,In_1944,In_1211);
nand U4495 (N_4495,In_440,In_351);
xnor U4496 (N_4496,In_544,In_840);
nand U4497 (N_4497,In_1128,In_469);
nor U4498 (N_4498,In_1691,In_1832);
or U4499 (N_4499,In_828,In_294);
nor U4500 (N_4500,In_900,In_1870);
or U4501 (N_4501,In_398,In_301);
xnor U4502 (N_4502,In_1868,In_116);
and U4503 (N_4503,In_302,In_1032);
xor U4504 (N_4504,In_1931,In_1252);
nor U4505 (N_4505,In_1015,In_1994);
nor U4506 (N_4506,In_685,In_1064);
nand U4507 (N_4507,In_168,In_587);
nor U4508 (N_4508,In_909,In_539);
nor U4509 (N_4509,In_1095,In_1926);
and U4510 (N_4510,In_1381,In_693);
or U4511 (N_4511,In_1800,In_838);
nand U4512 (N_4512,In_676,In_61);
nand U4513 (N_4513,In_410,In_1267);
nor U4514 (N_4514,In_1676,In_1586);
nor U4515 (N_4515,In_645,In_445);
nand U4516 (N_4516,In_48,In_199);
nor U4517 (N_4517,In_1552,In_1828);
nor U4518 (N_4518,In_110,In_689);
and U4519 (N_4519,In_264,In_1590);
xor U4520 (N_4520,In_1915,In_1409);
nor U4521 (N_4521,In_474,In_791);
nand U4522 (N_4522,In_1508,In_1221);
nand U4523 (N_4523,In_1520,In_142);
nand U4524 (N_4524,In_428,In_557);
or U4525 (N_4525,In_1990,In_1777);
and U4526 (N_4526,In_1533,In_1366);
or U4527 (N_4527,In_677,In_1998);
nor U4528 (N_4528,In_804,In_115);
nor U4529 (N_4529,In_483,In_230);
nor U4530 (N_4530,In_1069,In_1258);
or U4531 (N_4531,In_1954,In_331);
and U4532 (N_4532,In_1571,In_1433);
xor U4533 (N_4533,In_1548,In_1532);
or U4534 (N_4534,In_1471,In_79);
and U4535 (N_4535,In_1929,In_761);
nand U4536 (N_4536,In_157,In_90);
and U4537 (N_4537,In_190,In_932);
xor U4538 (N_4538,In_173,In_910);
or U4539 (N_4539,In_1925,In_737);
and U4540 (N_4540,In_11,In_58);
nor U4541 (N_4541,In_1816,In_1459);
or U4542 (N_4542,In_689,In_1397);
nand U4543 (N_4543,In_1123,In_1279);
xor U4544 (N_4544,In_1704,In_377);
nor U4545 (N_4545,In_138,In_1210);
nand U4546 (N_4546,In_1943,In_118);
nor U4547 (N_4547,In_884,In_1153);
and U4548 (N_4548,In_1093,In_1849);
or U4549 (N_4549,In_172,In_1684);
and U4550 (N_4550,In_1552,In_1170);
nand U4551 (N_4551,In_701,In_762);
nand U4552 (N_4552,In_908,In_277);
nand U4553 (N_4553,In_466,In_52);
nor U4554 (N_4554,In_626,In_15);
xnor U4555 (N_4555,In_144,In_729);
nand U4556 (N_4556,In_393,In_1933);
xnor U4557 (N_4557,In_1898,In_521);
nor U4558 (N_4558,In_62,In_94);
and U4559 (N_4559,In_343,In_380);
nand U4560 (N_4560,In_1530,In_914);
nand U4561 (N_4561,In_282,In_1892);
or U4562 (N_4562,In_1928,In_518);
nor U4563 (N_4563,In_715,In_1356);
nor U4564 (N_4564,In_1810,In_1861);
nor U4565 (N_4565,In_727,In_1745);
or U4566 (N_4566,In_1278,In_1717);
nand U4567 (N_4567,In_1155,In_664);
nand U4568 (N_4568,In_954,In_768);
or U4569 (N_4569,In_1525,In_816);
nor U4570 (N_4570,In_969,In_9);
xor U4571 (N_4571,In_1435,In_154);
nor U4572 (N_4572,In_1765,In_27);
nor U4573 (N_4573,In_450,In_1552);
nor U4574 (N_4574,In_1109,In_180);
xnor U4575 (N_4575,In_1291,In_1279);
or U4576 (N_4576,In_862,In_342);
nor U4577 (N_4577,In_1487,In_1656);
nand U4578 (N_4578,In_597,In_1679);
nor U4579 (N_4579,In_1953,In_1227);
xnor U4580 (N_4580,In_1512,In_68);
nand U4581 (N_4581,In_497,In_1665);
nand U4582 (N_4582,In_945,In_321);
xnor U4583 (N_4583,In_613,In_1579);
and U4584 (N_4584,In_1205,In_1135);
nor U4585 (N_4585,In_1415,In_282);
or U4586 (N_4586,In_1280,In_190);
or U4587 (N_4587,In_1701,In_673);
or U4588 (N_4588,In_376,In_1854);
nand U4589 (N_4589,In_722,In_534);
and U4590 (N_4590,In_1688,In_207);
xor U4591 (N_4591,In_220,In_306);
nor U4592 (N_4592,In_1078,In_938);
nor U4593 (N_4593,In_950,In_1215);
nand U4594 (N_4594,In_1524,In_1547);
xnor U4595 (N_4595,In_1572,In_1252);
xor U4596 (N_4596,In_1849,In_1416);
nor U4597 (N_4597,In_224,In_919);
nor U4598 (N_4598,In_771,In_48);
or U4599 (N_4599,In_1846,In_802);
nor U4600 (N_4600,In_672,In_197);
or U4601 (N_4601,In_169,In_1579);
or U4602 (N_4602,In_1858,In_1576);
and U4603 (N_4603,In_1095,In_1920);
nor U4604 (N_4604,In_337,In_329);
and U4605 (N_4605,In_306,In_72);
nand U4606 (N_4606,In_189,In_513);
and U4607 (N_4607,In_1081,In_1099);
or U4608 (N_4608,In_69,In_1702);
nand U4609 (N_4609,In_1417,In_1205);
nor U4610 (N_4610,In_1821,In_380);
nor U4611 (N_4611,In_809,In_1716);
or U4612 (N_4612,In_194,In_666);
nor U4613 (N_4613,In_1649,In_1793);
or U4614 (N_4614,In_1422,In_1142);
and U4615 (N_4615,In_606,In_1208);
xor U4616 (N_4616,In_1240,In_1554);
and U4617 (N_4617,In_1029,In_1121);
xnor U4618 (N_4618,In_312,In_465);
and U4619 (N_4619,In_167,In_1895);
or U4620 (N_4620,In_1050,In_1288);
and U4621 (N_4621,In_452,In_223);
or U4622 (N_4622,In_774,In_1882);
or U4623 (N_4623,In_803,In_128);
nor U4624 (N_4624,In_1891,In_346);
nand U4625 (N_4625,In_1071,In_1298);
or U4626 (N_4626,In_1537,In_1170);
and U4627 (N_4627,In_1541,In_427);
and U4628 (N_4628,In_1561,In_342);
nand U4629 (N_4629,In_837,In_6);
nor U4630 (N_4630,In_439,In_965);
nand U4631 (N_4631,In_133,In_1469);
nor U4632 (N_4632,In_302,In_664);
and U4633 (N_4633,In_638,In_721);
or U4634 (N_4634,In_1840,In_1156);
nand U4635 (N_4635,In_406,In_1676);
nor U4636 (N_4636,In_336,In_704);
and U4637 (N_4637,In_776,In_1962);
or U4638 (N_4638,In_660,In_1019);
and U4639 (N_4639,In_649,In_1736);
nor U4640 (N_4640,In_1456,In_1039);
nor U4641 (N_4641,In_1757,In_188);
nand U4642 (N_4642,In_1362,In_214);
or U4643 (N_4643,In_1987,In_1539);
and U4644 (N_4644,In_1988,In_1896);
xor U4645 (N_4645,In_214,In_769);
nand U4646 (N_4646,In_696,In_372);
nand U4647 (N_4647,In_1589,In_1746);
nor U4648 (N_4648,In_702,In_1908);
or U4649 (N_4649,In_1255,In_1269);
and U4650 (N_4650,In_1105,In_1092);
nor U4651 (N_4651,In_1367,In_399);
or U4652 (N_4652,In_728,In_360);
nand U4653 (N_4653,In_631,In_1838);
xor U4654 (N_4654,In_1313,In_1474);
or U4655 (N_4655,In_1387,In_1033);
nand U4656 (N_4656,In_1822,In_1238);
nand U4657 (N_4657,In_236,In_961);
and U4658 (N_4658,In_374,In_900);
or U4659 (N_4659,In_1475,In_237);
xor U4660 (N_4660,In_395,In_1003);
and U4661 (N_4661,In_832,In_320);
xnor U4662 (N_4662,In_839,In_3);
or U4663 (N_4663,In_1012,In_1815);
and U4664 (N_4664,In_200,In_1894);
nand U4665 (N_4665,In_3,In_297);
and U4666 (N_4666,In_1840,In_395);
and U4667 (N_4667,In_1989,In_282);
nand U4668 (N_4668,In_1976,In_154);
or U4669 (N_4669,In_508,In_1757);
or U4670 (N_4670,In_1398,In_39);
nor U4671 (N_4671,In_79,In_253);
and U4672 (N_4672,In_1938,In_1066);
nor U4673 (N_4673,In_1551,In_186);
nor U4674 (N_4674,In_1837,In_59);
nand U4675 (N_4675,In_763,In_1305);
nor U4676 (N_4676,In_1248,In_976);
nand U4677 (N_4677,In_338,In_1017);
nor U4678 (N_4678,In_1960,In_624);
or U4679 (N_4679,In_1584,In_921);
and U4680 (N_4680,In_843,In_1885);
nor U4681 (N_4681,In_195,In_146);
nor U4682 (N_4682,In_1656,In_483);
or U4683 (N_4683,In_1029,In_1158);
or U4684 (N_4684,In_1254,In_650);
xor U4685 (N_4685,In_115,In_1484);
nand U4686 (N_4686,In_207,In_757);
or U4687 (N_4687,In_1118,In_1901);
or U4688 (N_4688,In_1303,In_1952);
xnor U4689 (N_4689,In_1749,In_986);
or U4690 (N_4690,In_1075,In_400);
xor U4691 (N_4691,In_1726,In_1385);
or U4692 (N_4692,In_326,In_1132);
and U4693 (N_4693,In_649,In_1008);
nor U4694 (N_4694,In_1580,In_750);
nor U4695 (N_4695,In_1338,In_1592);
nand U4696 (N_4696,In_695,In_116);
and U4697 (N_4697,In_446,In_1678);
and U4698 (N_4698,In_1668,In_33);
and U4699 (N_4699,In_419,In_735);
nor U4700 (N_4700,In_86,In_1783);
nor U4701 (N_4701,In_21,In_756);
nand U4702 (N_4702,In_609,In_95);
xor U4703 (N_4703,In_282,In_870);
nor U4704 (N_4704,In_339,In_842);
or U4705 (N_4705,In_1846,In_1170);
and U4706 (N_4706,In_240,In_1270);
or U4707 (N_4707,In_1922,In_413);
nand U4708 (N_4708,In_448,In_729);
xnor U4709 (N_4709,In_674,In_679);
nand U4710 (N_4710,In_1179,In_1285);
nor U4711 (N_4711,In_715,In_1839);
and U4712 (N_4712,In_997,In_1504);
nand U4713 (N_4713,In_670,In_1221);
and U4714 (N_4714,In_98,In_22);
nand U4715 (N_4715,In_1188,In_1212);
nand U4716 (N_4716,In_481,In_1050);
or U4717 (N_4717,In_1088,In_1724);
nand U4718 (N_4718,In_1319,In_126);
and U4719 (N_4719,In_1230,In_1328);
nor U4720 (N_4720,In_1857,In_1880);
or U4721 (N_4721,In_1397,In_713);
nor U4722 (N_4722,In_734,In_781);
or U4723 (N_4723,In_256,In_375);
and U4724 (N_4724,In_519,In_1763);
nor U4725 (N_4725,In_1908,In_220);
nor U4726 (N_4726,In_773,In_624);
nor U4727 (N_4727,In_489,In_47);
nor U4728 (N_4728,In_1339,In_1319);
or U4729 (N_4729,In_1398,In_937);
and U4730 (N_4730,In_554,In_140);
xnor U4731 (N_4731,In_110,In_1043);
nor U4732 (N_4732,In_1936,In_1406);
and U4733 (N_4733,In_1803,In_1160);
xnor U4734 (N_4734,In_312,In_1288);
or U4735 (N_4735,In_63,In_405);
or U4736 (N_4736,In_1023,In_1747);
nand U4737 (N_4737,In_329,In_805);
nand U4738 (N_4738,In_665,In_1092);
xor U4739 (N_4739,In_735,In_1389);
or U4740 (N_4740,In_1750,In_1736);
and U4741 (N_4741,In_1507,In_478);
and U4742 (N_4742,In_495,In_827);
nand U4743 (N_4743,In_777,In_183);
nand U4744 (N_4744,In_939,In_1958);
or U4745 (N_4745,In_960,In_498);
and U4746 (N_4746,In_470,In_1775);
or U4747 (N_4747,In_743,In_355);
and U4748 (N_4748,In_830,In_1889);
nand U4749 (N_4749,In_1539,In_358);
nand U4750 (N_4750,In_1861,In_795);
nand U4751 (N_4751,In_359,In_1707);
and U4752 (N_4752,In_61,In_1604);
or U4753 (N_4753,In_473,In_281);
nor U4754 (N_4754,In_763,In_850);
nand U4755 (N_4755,In_485,In_1930);
xnor U4756 (N_4756,In_905,In_939);
or U4757 (N_4757,In_1877,In_1729);
or U4758 (N_4758,In_1337,In_926);
nor U4759 (N_4759,In_892,In_1836);
or U4760 (N_4760,In_499,In_355);
nand U4761 (N_4761,In_959,In_1120);
and U4762 (N_4762,In_1672,In_1281);
or U4763 (N_4763,In_1012,In_827);
nand U4764 (N_4764,In_1336,In_1542);
nor U4765 (N_4765,In_346,In_461);
nor U4766 (N_4766,In_1793,In_1550);
nand U4767 (N_4767,In_747,In_1817);
nor U4768 (N_4768,In_1003,In_167);
and U4769 (N_4769,In_1299,In_218);
nor U4770 (N_4770,In_116,In_73);
and U4771 (N_4771,In_1422,In_333);
nand U4772 (N_4772,In_1456,In_358);
nor U4773 (N_4773,In_84,In_218);
or U4774 (N_4774,In_483,In_1224);
xor U4775 (N_4775,In_732,In_573);
and U4776 (N_4776,In_1324,In_436);
nor U4777 (N_4777,In_695,In_1098);
or U4778 (N_4778,In_1650,In_663);
and U4779 (N_4779,In_441,In_1090);
and U4780 (N_4780,In_1214,In_694);
or U4781 (N_4781,In_1776,In_656);
nand U4782 (N_4782,In_48,In_117);
nand U4783 (N_4783,In_1750,In_553);
and U4784 (N_4784,In_1869,In_982);
and U4785 (N_4785,In_1922,In_1525);
and U4786 (N_4786,In_892,In_1823);
nor U4787 (N_4787,In_1692,In_1713);
nor U4788 (N_4788,In_1263,In_1432);
xnor U4789 (N_4789,In_587,In_719);
nand U4790 (N_4790,In_255,In_232);
or U4791 (N_4791,In_909,In_1921);
nor U4792 (N_4792,In_1307,In_433);
nand U4793 (N_4793,In_787,In_26);
or U4794 (N_4794,In_1737,In_693);
or U4795 (N_4795,In_1325,In_576);
or U4796 (N_4796,In_1254,In_686);
or U4797 (N_4797,In_151,In_310);
nand U4798 (N_4798,In_182,In_853);
nor U4799 (N_4799,In_1749,In_660);
xor U4800 (N_4800,In_103,In_985);
or U4801 (N_4801,In_1193,In_1742);
nor U4802 (N_4802,In_1188,In_1014);
nand U4803 (N_4803,In_1430,In_1161);
nor U4804 (N_4804,In_353,In_1529);
nor U4805 (N_4805,In_400,In_842);
or U4806 (N_4806,In_1207,In_150);
or U4807 (N_4807,In_386,In_376);
or U4808 (N_4808,In_510,In_874);
nand U4809 (N_4809,In_1114,In_1322);
nand U4810 (N_4810,In_101,In_394);
or U4811 (N_4811,In_1837,In_781);
nor U4812 (N_4812,In_227,In_523);
nor U4813 (N_4813,In_1100,In_141);
nor U4814 (N_4814,In_1859,In_1224);
and U4815 (N_4815,In_1310,In_273);
or U4816 (N_4816,In_358,In_1184);
or U4817 (N_4817,In_1608,In_1511);
and U4818 (N_4818,In_210,In_1725);
nor U4819 (N_4819,In_106,In_21);
nand U4820 (N_4820,In_1939,In_1144);
nor U4821 (N_4821,In_1602,In_402);
or U4822 (N_4822,In_1881,In_1314);
or U4823 (N_4823,In_175,In_1643);
and U4824 (N_4824,In_469,In_1871);
nand U4825 (N_4825,In_1957,In_1025);
xor U4826 (N_4826,In_1591,In_1219);
and U4827 (N_4827,In_1345,In_1923);
and U4828 (N_4828,In_381,In_1043);
and U4829 (N_4829,In_1655,In_763);
nor U4830 (N_4830,In_983,In_1788);
xnor U4831 (N_4831,In_1412,In_974);
nand U4832 (N_4832,In_1190,In_1575);
nand U4833 (N_4833,In_1367,In_1673);
and U4834 (N_4834,In_1949,In_1430);
and U4835 (N_4835,In_823,In_437);
nand U4836 (N_4836,In_205,In_617);
nor U4837 (N_4837,In_1827,In_973);
or U4838 (N_4838,In_1354,In_1011);
nor U4839 (N_4839,In_1523,In_1487);
nand U4840 (N_4840,In_491,In_1064);
and U4841 (N_4841,In_1762,In_1956);
and U4842 (N_4842,In_725,In_606);
and U4843 (N_4843,In_1359,In_1613);
xnor U4844 (N_4844,In_710,In_904);
or U4845 (N_4845,In_241,In_638);
or U4846 (N_4846,In_1251,In_1041);
and U4847 (N_4847,In_258,In_265);
xor U4848 (N_4848,In_878,In_762);
nand U4849 (N_4849,In_390,In_1896);
nor U4850 (N_4850,In_1090,In_1244);
nand U4851 (N_4851,In_1530,In_656);
nor U4852 (N_4852,In_1427,In_512);
nor U4853 (N_4853,In_1984,In_250);
xnor U4854 (N_4854,In_1292,In_1148);
or U4855 (N_4855,In_1599,In_1364);
or U4856 (N_4856,In_1172,In_343);
and U4857 (N_4857,In_242,In_1208);
nand U4858 (N_4858,In_482,In_1778);
and U4859 (N_4859,In_1685,In_1482);
xnor U4860 (N_4860,In_1054,In_1060);
nand U4861 (N_4861,In_731,In_717);
or U4862 (N_4862,In_1242,In_225);
and U4863 (N_4863,In_1109,In_1754);
nand U4864 (N_4864,In_1033,In_1514);
nand U4865 (N_4865,In_1824,In_1235);
nand U4866 (N_4866,In_863,In_1984);
nand U4867 (N_4867,In_39,In_476);
and U4868 (N_4868,In_812,In_1110);
nand U4869 (N_4869,In_1381,In_1187);
nand U4870 (N_4870,In_1594,In_871);
and U4871 (N_4871,In_1348,In_104);
and U4872 (N_4872,In_323,In_1071);
or U4873 (N_4873,In_1391,In_918);
nor U4874 (N_4874,In_1659,In_461);
and U4875 (N_4875,In_696,In_1061);
nand U4876 (N_4876,In_1850,In_1228);
and U4877 (N_4877,In_544,In_283);
and U4878 (N_4878,In_851,In_1425);
and U4879 (N_4879,In_1672,In_255);
or U4880 (N_4880,In_825,In_541);
xnor U4881 (N_4881,In_296,In_731);
or U4882 (N_4882,In_748,In_1195);
and U4883 (N_4883,In_1340,In_1901);
and U4884 (N_4884,In_640,In_794);
xnor U4885 (N_4885,In_735,In_563);
nand U4886 (N_4886,In_1933,In_1819);
xor U4887 (N_4887,In_1864,In_240);
and U4888 (N_4888,In_215,In_654);
or U4889 (N_4889,In_149,In_1825);
or U4890 (N_4890,In_772,In_1899);
or U4891 (N_4891,In_1476,In_605);
or U4892 (N_4892,In_1773,In_1002);
nand U4893 (N_4893,In_1174,In_1366);
and U4894 (N_4894,In_299,In_1316);
or U4895 (N_4895,In_1418,In_831);
xnor U4896 (N_4896,In_538,In_137);
nor U4897 (N_4897,In_1385,In_379);
or U4898 (N_4898,In_147,In_743);
nor U4899 (N_4899,In_1761,In_1382);
nor U4900 (N_4900,In_475,In_1822);
xor U4901 (N_4901,In_270,In_1685);
or U4902 (N_4902,In_442,In_1945);
xnor U4903 (N_4903,In_1230,In_1567);
or U4904 (N_4904,In_173,In_1452);
nand U4905 (N_4905,In_1993,In_1386);
nor U4906 (N_4906,In_1197,In_1248);
nand U4907 (N_4907,In_756,In_740);
or U4908 (N_4908,In_762,In_155);
nor U4909 (N_4909,In_1879,In_725);
or U4910 (N_4910,In_1222,In_1947);
nor U4911 (N_4911,In_103,In_695);
nor U4912 (N_4912,In_1145,In_1158);
or U4913 (N_4913,In_963,In_771);
and U4914 (N_4914,In_56,In_642);
nand U4915 (N_4915,In_1714,In_1853);
or U4916 (N_4916,In_1699,In_346);
or U4917 (N_4917,In_1267,In_324);
and U4918 (N_4918,In_598,In_1619);
nand U4919 (N_4919,In_525,In_1495);
xnor U4920 (N_4920,In_1379,In_860);
xor U4921 (N_4921,In_1178,In_1441);
and U4922 (N_4922,In_1333,In_532);
nand U4923 (N_4923,In_136,In_1633);
nand U4924 (N_4924,In_1741,In_1084);
and U4925 (N_4925,In_1666,In_1404);
or U4926 (N_4926,In_1175,In_736);
and U4927 (N_4927,In_874,In_930);
or U4928 (N_4928,In_504,In_1998);
xor U4929 (N_4929,In_1245,In_1828);
and U4930 (N_4930,In_1806,In_395);
nor U4931 (N_4931,In_747,In_1668);
and U4932 (N_4932,In_1135,In_1816);
or U4933 (N_4933,In_685,In_1955);
nand U4934 (N_4934,In_567,In_1599);
or U4935 (N_4935,In_1007,In_93);
xnor U4936 (N_4936,In_806,In_375);
and U4937 (N_4937,In_723,In_980);
nor U4938 (N_4938,In_1805,In_1455);
and U4939 (N_4939,In_1972,In_521);
nor U4940 (N_4940,In_1208,In_1158);
and U4941 (N_4941,In_1797,In_128);
or U4942 (N_4942,In_1411,In_1796);
or U4943 (N_4943,In_1197,In_1889);
nand U4944 (N_4944,In_1793,In_1351);
and U4945 (N_4945,In_137,In_226);
xnor U4946 (N_4946,In_1469,In_1235);
nand U4947 (N_4947,In_1557,In_1072);
nor U4948 (N_4948,In_174,In_1050);
or U4949 (N_4949,In_359,In_367);
nor U4950 (N_4950,In_1982,In_1802);
or U4951 (N_4951,In_1115,In_1495);
and U4952 (N_4952,In_1491,In_892);
or U4953 (N_4953,In_307,In_1509);
nor U4954 (N_4954,In_49,In_1934);
nor U4955 (N_4955,In_548,In_678);
nand U4956 (N_4956,In_1696,In_1540);
nand U4957 (N_4957,In_1312,In_1305);
xnor U4958 (N_4958,In_1123,In_1076);
nand U4959 (N_4959,In_285,In_1997);
or U4960 (N_4960,In_1715,In_1801);
and U4961 (N_4961,In_1848,In_1100);
xor U4962 (N_4962,In_1131,In_216);
nand U4963 (N_4963,In_489,In_611);
xnor U4964 (N_4964,In_1882,In_1504);
and U4965 (N_4965,In_1738,In_531);
nor U4966 (N_4966,In_1378,In_965);
and U4967 (N_4967,In_455,In_1818);
xor U4968 (N_4968,In_11,In_1023);
or U4969 (N_4969,In_99,In_1078);
xor U4970 (N_4970,In_788,In_1295);
and U4971 (N_4971,In_428,In_205);
or U4972 (N_4972,In_1533,In_143);
nand U4973 (N_4973,In_478,In_596);
and U4974 (N_4974,In_1970,In_1245);
xnor U4975 (N_4975,In_1586,In_1273);
nand U4976 (N_4976,In_1850,In_384);
or U4977 (N_4977,In_1511,In_1908);
nand U4978 (N_4978,In_924,In_404);
nand U4979 (N_4979,In_607,In_530);
and U4980 (N_4980,In_919,In_1639);
or U4981 (N_4981,In_261,In_522);
nor U4982 (N_4982,In_368,In_621);
xor U4983 (N_4983,In_450,In_1962);
and U4984 (N_4984,In_179,In_1775);
or U4985 (N_4985,In_1148,In_1416);
xor U4986 (N_4986,In_979,In_290);
nor U4987 (N_4987,In_1962,In_1103);
nand U4988 (N_4988,In_1301,In_1386);
nor U4989 (N_4989,In_440,In_826);
or U4990 (N_4990,In_446,In_439);
and U4991 (N_4991,In_1743,In_358);
xor U4992 (N_4992,In_670,In_1028);
nor U4993 (N_4993,In_1842,In_1718);
xor U4994 (N_4994,In_1452,In_27);
or U4995 (N_4995,In_346,In_401);
nand U4996 (N_4996,In_602,In_114);
and U4997 (N_4997,In_1474,In_1352);
nor U4998 (N_4998,In_771,In_1342);
or U4999 (N_4999,In_1139,In_436);
or U5000 (N_5000,N_2065,N_1128);
nand U5001 (N_5001,N_372,N_212);
and U5002 (N_5002,N_4833,N_1281);
or U5003 (N_5003,N_4357,N_3672);
nand U5004 (N_5004,N_836,N_4474);
nor U5005 (N_5005,N_1982,N_646);
or U5006 (N_5006,N_1344,N_2122);
nor U5007 (N_5007,N_2584,N_2177);
or U5008 (N_5008,N_2201,N_2355);
nand U5009 (N_5009,N_2029,N_4301);
and U5010 (N_5010,N_4804,N_1846);
and U5011 (N_5011,N_1820,N_2986);
nor U5012 (N_5012,N_3922,N_3183);
and U5013 (N_5013,N_3342,N_2024);
nor U5014 (N_5014,N_1648,N_3288);
nor U5015 (N_5015,N_1000,N_1441);
nand U5016 (N_5016,N_1288,N_2540);
nor U5017 (N_5017,N_3262,N_2157);
or U5018 (N_5018,N_1657,N_2794);
nor U5019 (N_5019,N_4038,N_3446);
and U5020 (N_5020,N_3792,N_2600);
nand U5021 (N_5021,N_50,N_4839);
nor U5022 (N_5022,N_1445,N_2840);
nand U5023 (N_5023,N_2740,N_2070);
nor U5024 (N_5024,N_713,N_3799);
nor U5025 (N_5025,N_1094,N_4448);
or U5026 (N_5026,N_4813,N_1237);
nand U5027 (N_5027,N_363,N_3217);
nand U5028 (N_5028,N_2638,N_4486);
and U5029 (N_5029,N_835,N_1766);
xor U5030 (N_5030,N_1834,N_4120);
and U5031 (N_5031,N_91,N_2333);
or U5032 (N_5032,N_3177,N_4792);
and U5033 (N_5033,N_3381,N_2532);
or U5034 (N_5034,N_1419,N_3335);
or U5035 (N_5035,N_3461,N_2906);
and U5036 (N_5036,N_4197,N_782);
xor U5037 (N_5037,N_2612,N_1059);
nand U5038 (N_5038,N_3762,N_3598);
or U5039 (N_5039,N_52,N_4519);
nor U5040 (N_5040,N_3736,N_1244);
or U5041 (N_5041,N_3425,N_3948);
nand U5042 (N_5042,N_678,N_522);
xnor U5043 (N_5043,N_657,N_2008);
nor U5044 (N_5044,N_2851,N_2508);
nor U5045 (N_5045,N_3710,N_2243);
or U5046 (N_5046,N_720,N_2132);
or U5047 (N_5047,N_2002,N_970);
or U5048 (N_5048,N_2888,N_1105);
and U5049 (N_5049,N_2464,N_350);
or U5050 (N_5050,N_1721,N_2629);
xor U5051 (N_5051,N_4642,N_1394);
or U5052 (N_5052,N_4171,N_4596);
and U5053 (N_5053,N_4941,N_127);
xnor U5054 (N_5054,N_3773,N_4442);
nand U5055 (N_5055,N_532,N_3173);
nand U5056 (N_5056,N_3210,N_1850);
and U5057 (N_5057,N_2302,N_1051);
xnor U5058 (N_5058,N_3485,N_1476);
or U5059 (N_5059,N_1465,N_2968);
or U5060 (N_5060,N_4317,N_445);
nor U5061 (N_5061,N_4506,N_3546);
and U5062 (N_5062,N_130,N_4084);
and U5063 (N_5063,N_563,N_821);
xor U5064 (N_5064,N_510,N_1907);
and U5065 (N_5065,N_2783,N_811);
xor U5066 (N_5066,N_3236,N_3976);
nand U5067 (N_5067,N_1985,N_3194);
nor U5068 (N_5068,N_2007,N_635);
or U5069 (N_5069,N_2488,N_496);
nor U5070 (N_5070,N_1359,N_1936);
nand U5071 (N_5071,N_2556,N_2330);
and U5072 (N_5072,N_2490,N_4022);
or U5073 (N_5073,N_3121,N_136);
nand U5074 (N_5074,N_3149,N_3369);
xor U5075 (N_5075,N_723,N_4940);
nand U5076 (N_5076,N_1809,N_1799);
nor U5077 (N_5077,N_3140,N_83);
or U5078 (N_5078,N_3768,N_2087);
and U5079 (N_5079,N_96,N_2475);
nor U5080 (N_5080,N_2032,N_1172);
or U5081 (N_5081,N_2604,N_2648);
or U5082 (N_5082,N_3919,N_4966);
and U5083 (N_5083,N_1602,N_253);
or U5084 (N_5084,N_1792,N_2745);
nor U5085 (N_5085,N_3480,N_3650);
nand U5086 (N_5086,N_829,N_775);
and U5087 (N_5087,N_1502,N_4153);
nor U5088 (N_5088,N_2420,N_3915);
nand U5089 (N_5089,N_1005,N_3017);
and U5090 (N_5090,N_3315,N_693);
nand U5091 (N_5091,N_1246,N_4330);
and U5092 (N_5092,N_1925,N_4849);
xnor U5093 (N_5093,N_3793,N_4081);
nor U5094 (N_5094,N_4321,N_3327);
and U5095 (N_5095,N_3898,N_4706);
or U5096 (N_5096,N_77,N_1510);
and U5097 (N_5097,N_2790,N_3040);
nand U5098 (N_5098,N_2390,N_3797);
nand U5099 (N_5099,N_4622,N_2014);
and U5100 (N_5100,N_4551,N_4463);
and U5101 (N_5101,N_567,N_1975);
or U5102 (N_5102,N_4384,N_3463);
or U5103 (N_5103,N_3239,N_1178);
xor U5104 (N_5104,N_1739,N_3902);
or U5105 (N_5105,N_1628,N_3503);
nand U5106 (N_5106,N_1368,N_3712);
and U5107 (N_5107,N_2690,N_1836);
and U5108 (N_5108,N_1221,N_3864);
nand U5109 (N_5109,N_4736,N_1670);
and U5110 (N_5110,N_2356,N_383);
and U5111 (N_5111,N_1578,N_3355);
or U5112 (N_5112,N_4238,N_4006);
or U5113 (N_5113,N_3493,N_118);
xor U5114 (N_5114,N_2166,N_2130);
and U5115 (N_5115,N_2416,N_147);
nand U5116 (N_5116,N_1370,N_2715);
nand U5117 (N_5117,N_3548,N_3527);
or U5118 (N_5118,N_979,N_4897);
or U5119 (N_5119,N_3855,N_568);
and U5120 (N_5120,N_1631,N_4196);
and U5121 (N_5121,N_4776,N_349);
xnor U5122 (N_5122,N_1129,N_852);
xnor U5123 (N_5123,N_733,N_2077);
nand U5124 (N_5124,N_2587,N_2304);
nand U5125 (N_5125,N_1560,N_272);
or U5126 (N_5126,N_1802,N_1414);
and U5127 (N_5127,N_1483,N_4845);
or U5128 (N_5128,N_1046,N_287);
nor U5129 (N_5129,N_1467,N_4447);
or U5130 (N_5130,N_184,N_3406);
nor U5131 (N_5131,N_3636,N_1352);
and U5132 (N_5132,N_3639,N_2607);
and U5133 (N_5133,N_3723,N_3640);
nand U5134 (N_5134,N_433,N_4546);
and U5135 (N_5135,N_3229,N_4691);
nor U5136 (N_5136,N_1089,N_1515);
nand U5137 (N_5137,N_4669,N_999);
or U5138 (N_5138,N_3404,N_3714);
nand U5139 (N_5139,N_4404,N_2322);
and U5140 (N_5140,N_3721,N_3862);
nor U5141 (N_5141,N_2621,N_4053);
or U5142 (N_5142,N_3302,N_931);
nor U5143 (N_5143,N_3811,N_3757);
nand U5144 (N_5144,N_1615,N_4619);
nand U5145 (N_5145,N_3600,N_3705);
or U5146 (N_5146,N_3963,N_834);
or U5147 (N_5147,N_2897,N_4856);
and U5148 (N_5148,N_2868,N_1138);
xnor U5149 (N_5149,N_4117,N_3336);
nand U5150 (N_5150,N_4959,N_1685);
and U5151 (N_5151,N_355,N_735);
nand U5152 (N_5152,N_3087,N_2610);
and U5153 (N_5153,N_842,N_235);
nand U5154 (N_5154,N_3682,N_4139);
or U5155 (N_5155,N_3502,N_1176);
or U5156 (N_5156,N_3621,N_4620);
xor U5157 (N_5157,N_4590,N_4103);
or U5158 (N_5158,N_181,N_2431);
xnor U5159 (N_5159,N_1098,N_3585);
nand U5160 (N_5160,N_345,N_4871);
xor U5161 (N_5161,N_3088,N_2775);
or U5162 (N_5162,N_61,N_1842);
nand U5163 (N_5163,N_1960,N_3899);
nor U5164 (N_5164,N_5,N_3993);
or U5165 (N_5165,N_647,N_4394);
nor U5166 (N_5166,N_110,N_525);
and U5167 (N_5167,N_407,N_66);
nor U5168 (N_5168,N_4921,N_1177);
nand U5169 (N_5169,N_3876,N_4502);
xor U5170 (N_5170,N_692,N_3592);
nor U5171 (N_5171,N_3286,N_92);
nor U5172 (N_5172,N_2440,N_387);
nor U5173 (N_5173,N_2729,N_1010);
or U5174 (N_5174,N_2593,N_1054);
nand U5175 (N_5175,N_4529,N_295);
nand U5176 (N_5176,N_4070,N_4294);
or U5177 (N_5177,N_4743,N_280);
and U5178 (N_5178,N_4418,N_3354);
nor U5179 (N_5179,N_4499,N_892);
xnor U5180 (N_5180,N_1438,N_2493);
nand U5181 (N_5181,N_1191,N_1035);
nand U5182 (N_5182,N_3588,N_4949);
and U5183 (N_5183,N_544,N_1447);
or U5184 (N_5184,N_204,N_3159);
and U5185 (N_5185,N_4641,N_710);
or U5186 (N_5186,N_2052,N_3371);
xor U5187 (N_5187,N_164,N_312);
nor U5188 (N_5188,N_1422,N_4326);
or U5189 (N_5189,N_2927,N_1524);
or U5190 (N_5190,N_4489,N_2108);
and U5191 (N_5191,N_401,N_2206);
and U5192 (N_5192,N_113,N_1143);
and U5193 (N_5193,N_4808,N_3624);
nand U5194 (N_5194,N_3142,N_1120);
or U5195 (N_5195,N_2997,N_1998);
xor U5196 (N_5196,N_4775,N_2458);
and U5197 (N_5197,N_3104,N_3412);
and U5198 (N_5198,N_1558,N_565);
and U5199 (N_5199,N_1999,N_4824);
and U5200 (N_5200,N_785,N_2387);
nor U5201 (N_5201,N_2164,N_4251);
or U5202 (N_5202,N_648,N_4112);
nand U5203 (N_5203,N_4748,N_4476);
nor U5204 (N_5204,N_236,N_4780);
nand U5205 (N_5205,N_1231,N_3826);
nor U5206 (N_5206,N_4073,N_1581);
and U5207 (N_5207,N_2375,N_3587);
nand U5208 (N_5208,N_1145,N_3802);
nand U5209 (N_5209,N_3998,N_644);
and U5210 (N_5210,N_3837,N_4246);
nor U5211 (N_5211,N_4388,N_1884);
and U5212 (N_5212,N_1482,N_3781);
and U5213 (N_5213,N_4977,N_1630);
nor U5214 (N_5214,N_4284,N_4511);
and U5215 (N_5215,N_40,N_2925);
xnor U5216 (N_5216,N_537,N_3035);
or U5217 (N_5217,N_2882,N_3528);
and U5218 (N_5218,N_2218,N_1015);
nand U5219 (N_5219,N_3994,N_2209);
or U5220 (N_5220,N_4342,N_1421);
or U5221 (N_5221,N_4708,N_2161);
nor U5222 (N_5222,N_2739,N_2011);
nand U5223 (N_5223,N_279,N_2564);
and U5224 (N_5224,N_405,N_3324);
and U5225 (N_5225,N_768,N_882);
or U5226 (N_5226,N_1317,N_4344);
nor U5227 (N_5227,N_584,N_4233);
nand U5228 (N_5228,N_143,N_3407);
and U5229 (N_5229,N_4170,N_2038);
or U5230 (N_5230,N_3408,N_3658);
nor U5231 (N_5231,N_4850,N_4677);
nand U5232 (N_5232,N_1210,N_4547);
or U5233 (N_5233,N_1179,N_1541);
nand U5234 (N_5234,N_1978,N_4297);
nand U5235 (N_5235,N_14,N_192);
nor U5236 (N_5236,N_4907,N_3863);
or U5237 (N_5237,N_2449,N_4525);
nand U5238 (N_5238,N_2513,N_3129);
nor U5239 (N_5239,N_2833,N_1305);
nor U5240 (N_5240,N_2034,N_3794);
and U5241 (N_5241,N_1588,N_663);
or U5242 (N_5242,N_968,N_1226);
nor U5243 (N_5243,N_2760,N_331);
or U5244 (N_5244,N_3379,N_511);
nor U5245 (N_5245,N_4761,N_2784);
or U5246 (N_5246,N_912,N_4762);
nand U5247 (N_5247,N_4879,N_2048);
nand U5248 (N_5248,N_159,N_1045);
nor U5249 (N_5249,N_1082,N_131);
or U5250 (N_5250,N_2677,N_2598);
or U5251 (N_5251,N_4024,N_333);
and U5252 (N_5252,N_2365,N_1997);
nand U5253 (N_5253,N_2393,N_426);
xor U5254 (N_5254,N_1393,N_4711);
nand U5255 (N_5255,N_2175,N_4558);
nand U5256 (N_5256,N_357,N_4578);
or U5257 (N_5257,N_1885,N_2377);
nand U5258 (N_5258,N_1298,N_124);
nand U5259 (N_5259,N_1521,N_533);
nand U5260 (N_5260,N_3554,N_1617);
or U5261 (N_5261,N_20,N_1901);
nand U5262 (N_5262,N_3516,N_4473);
xnor U5263 (N_5263,N_1390,N_2310);
and U5264 (N_5264,N_753,N_589);
nand U5265 (N_5265,N_3929,N_2084);
and U5266 (N_5266,N_2191,N_3941);
and U5267 (N_5267,N_3137,N_1835);
nor U5268 (N_5268,N_701,N_960);
and U5269 (N_5269,N_930,N_4713);
nor U5270 (N_5270,N_4407,N_4655);
nand U5271 (N_5271,N_2703,N_4000);
or U5272 (N_5272,N_4605,N_1609);
nand U5273 (N_5273,N_1455,N_1944);
nand U5274 (N_5274,N_624,N_3534);
xnor U5275 (N_5275,N_2911,N_4247);
nor U5276 (N_5276,N_3633,N_4020);
and U5277 (N_5277,N_2866,N_3618);
and U5278 (N_5278,N_1469,N_2278);
and U5279 (N_5279,N_1994,N_4864);
nand U5280 (N_5280,N_2141,N_2114);
nor U5281 (N_5281,N_1036,N_865);
xnor U5282 (N_5282,N_1785,N_304);
nand U5283 (N_5283,N_2296,N_1109);
or U5284 (N_5284,N_2533,N_795);
xnor U5285 (N_5285,N_37,N_1219);
xnor U5286 (N_5286,N_4142,N_2263);
or U5287 (N_5287,N_2549,N_1879);
and U5288 (N_5288,N_2518,N_2428);
or U5289 (N_5289,N_3872,N_4441);
or U5290 (N_5290,N_1241,N_4143);
or U5291 (N_5291,N_4359,N_711);
or U5292 (N_5292,N_3367,N_1891);
nand U5293 (N_5293,N_1733,N_3535);
nor U5294 (N_5294,N_3244,N_1475);
or U5295 (N_5295,N_4696,N_2510);
xor U5296 (N_5296,N_237,N_3240);
and U5297 (N_5297,N_109,N_4612);
nor U5298 (N_5298,N_1584,N_247);
xnor U5299 (N_5299,N_4787,N_1488);
nor U5300 (N_5300,N_368,N_3257);
and U5301 (N_5301,N_4906,N_4099);
nor U5302 (N_5302,N_4094,N_1289);
nand U5303 (N_5303,N_4191,N_1740);
nand U5304 (N_5304,N_1201,N_318);
nand U5305 (N_5305,N_3195,N_794);
or U5306 (N_5306,N_4160,N_4505);
or U5307 (N_5307,N_3179,N_1550);
and U5308 (N_5308,N_807,N_594);
and U5309 (N_5309,N_2127,N_1913);
nor U5310 (N_5310,N_1424,N_7);
or U5311 (N_5311,N_798,N_1619);
nor U5312 (N_5312,N_1187,N_2687);
xnor U5313 (N_5313,N_144,N_1092);
or U5314 (N_5314,N_620,N_1800);
xnor U5315 (N_5315,N_2948,N_1859);
nor U5316 (N_5316,N_1634,N_1302);
nand U5317 (N_5317,N_1374,N_2168);
nand U5318 (N_5318,N_3048,N_3519);
nor U5319 (N_5319,N_277,N_1784);
and U5320 (N_5320,N_4935,N_1658);
and U5321 (N_5321,N_2244,N_1490);
and U5322 (N_5322,N_2592,N_4346);
nand U5323 (N_5323,N_3575,N_3847);
nor U5324 (N_5324,N_161,N_1681);
nand U5325 (N_5325,N_745,N_2696);
xor U5326 (N_5326,N_2438,N_728);
xnor U5327 (N_5327,N_1304,N_3831);
or U5328 (N_5328,N_3114,N_4415);
nor U5329 (N_5329,N_689,N_121);
nor U5330 (N_5330,N_634,N_1813);
and U5331 (N_5331,N_895,N_4784);
and U5332 (N_5332,N_1434,N_4789);
xor U5333 (N_5333,N_998,N_2324);
and U5334 (N_5334,N_2219,N_1941);
and U5335 (N_5335,N_2022,N_797);
nand U5336 (N_5336,N_410,N_4203);
nor U5337 (N_5337,N_2369,N_705);
and U5338 (N_5338,N_4456,N_2266);
and U5339 (N_5339,N_3850,N_397);
nand U5340 (N_5340,N_4887,N_4996);
nand U5341 (N_5341,N_4176,N_2234);
nor U5342 (N_5342,N_3440,N_1906);
and U5343 (N_5343,N_2863,N_4127);
xnor U5344 (N_5344,N_4704,N_3126);
nor U5345 (N_5345,N_412,N_1690);
xor U5346 (N_5346,N_427,N_1535);
nor U5347 (N_5347,N_721,N_4295);
or U5348 (N_5348,N_3134,N_2381);
nor U5349 (N_5349,N_1217,N_2554);
nor U5350 (N_5350,N_3127,N_3427);
or U5351 (N_5351,N_3190,N_1659);
nor U5352 (N_5352,N_1860,N_2712);
nor U5353 (N_5353,N_2994,N_1576);
nand U5354 (N_5354,N_1607,N_78);
nand U5355 (N_5355,N_2750,N_4583);
nor U5356 (N_5356,N_3096,N_849);
nand U5357 (N_5357,N_1212,N_4177);
or U5358 (N_5358,N_2290,N_3981);
and U5359 (N_5359,N_3489,N_1736);
and U5360 (N_5360,N_1349,N_3038);
and U5361 (N_5361,N_651,N_4594);
nor U5362 (N_5362,N_3321,N_18);
and U5363 (N_5363,N_1542,N_3323);
nand U5364 (N_5364,N_1009,N_12);
nor U5365 (N_5365,N_1471,N_2574);
and U5366 (N_5366,N_501,N_2853);
nor U5367 (N_5367,N_1182,N_4230);
or U5368 (N_5368,N_3816,N_3778);
xnor U5369 (N_5369,N_4403,N_3944);
or U5370 (N_5370,N_3277,N_676);
nand U5371 (N_5371,N_3809,N_2060);
xor U5372 (N_5372,N_4627,N_2432);
or U5373 (N_5373,N_289,N_826);
nor U5374 (N_5374,N_2547,N_2155);
nand U5375 (N_5375,N_1893,N_2625);
or U5376 (N_5376,N_53,N_838);
xnor U5377 (N_5377,N_2481,N_1153);
nand U5378 (N_5378,N_4178,N_3775);
and U5379 (N_5379,N_3281,N_2842);
nand U5380 (N_5380,N_2881,N_2992);
or U5381 (N_5381,N_2885,N_4148);
nor U5382 (N_5382,N_379,N_3662);
and U5383 (N_5383,N_1321,N_3078);
and U5384 (N_5384,N_1767,N_2681);
or U5385 (N_5385,N_3077,N_4210);
nand U5386 (N_5386,N_564,N_685);
or U5387 (N_5387,N_2269,N_4937);
xnor U5388 (N_5388,N_2981,N_3276);
or U5389 (N_5389,N_4125,N_1166);
and U5390 (N_5390,N_2688,N_2072);
nand U5391 (N_5391,N_2555,N_4309);
nor U5392 (N_5392,N_2661,N_2836);
or U5393 (N_5393,N_708,N_2928);
nor U5394 (N_5394,N_4207,N_3352);
and U5395 (N_5395,N_2673,N_2553);
and U5396 (N_5396,N_3258,N_4149);
nand U5397 (N_5397,N_2286,N_1222);
nor U5398 (N_5398,N_3569,N_3436);
nor U5399 (N_5399,N_530,N_3093);
xnor U5400 (N_5400,N_2485,N_1961);
or U5401 (N_5401,N_4324,N_4461);
nand U5402 (N_5402,N_44,N_3983);
or U5403 (N_5403,N_854,N_4009);
xnor U5404 (N_5404,N_1130,N_609);
nand U5405 (N_5405,N_3973,N_3168);
nor U5406 (N_5406,N_839,N_2829);
nor U5407 (N_5407,N_2765,N_3526);
nand U5408 (N_5408,N_937,N_702);
nor U5409 (N_5409,N_4698,N_758);
nand U5410 (N_5410,N_2354,N_1018);
nor U5411 (N_5411,N_54,N_3764);
or U5412 (N_5412,N_3691,N_2374);
nor U5413 (N_5413,N_416,N_1306);
or U5414 (N_5414,N_643,N_117);
nand U5415 (N_5415,N_2626,N_951);
nor U5416 (N_5416,N_1318,N_4422);
nand U5417 (N_5417,N_2147,N_2620);
and U5418 (N_5418,N_4678,N_2826);
nand U5419 (N_5419,N_2467,N_4090);
and U5420 (N_5420,N_4063,N_2382);
nand U5421 (N_5421,N_1077,N_3437);
nand U5422 (N_5422,N_2543,N_4536);
nand U5423 (N_5423,N_1671,N_536);
nor U5424 (N_5424,N_814,N_2216);
xor U5425 (N_5425,N_1559,N_3492);
xor U5426 (N_5426,N_3504,N_3115);
xor U5427 (N_5427,N_1292,N_1613);
or U5428 (N_5428,N_2635,N_1199);
and U5429 (N_5429,N_669,N_3709);
and U5430 (N_5430,N_1741,N_3499);
nand U5431 (N_5431,N_4161,N_1979);
or U5432 (N_5432,N_3590,N_2248);
or U5433 (N_5433,N_3197,N_3905);
or U5434 (N_5434,N_220,N_2531);
xnor U5435 (N_5435,N_3695,N_3843);
nand U5436 (N_5436,N_3267,N_2309);
nor U5437 (N_5437,N_995,N_3387);
or U5438 (N_5438,N_502,N_3042);
nand U5439 (N_5439,N_2086,N_4773);
and U5440 (N_5440,N_2984,N_894);
xnor U5441 (N_5441,N_4296,N_3685);
or U5442 (N_5442,N_3219,N_1543);
and U5443 (N_5443,N_4769,N_4255);
nor U5444 (N_5444,N_2349,N_600);
or U5445 (N_5445,N_2887,N_4540);
or U5446 (N_5446,N_4397,N_4962);
and U5447 (N_5447,N_3316,N_3012);
nor U5448 (N_5448,N_516,N_4515);
or U5449 (N_5449,N_439,N_1282);
xnor U5450 (N_5450,N_4348,N_4076);
nor U5451 (N_5451,N_945,N_3671);
nor U5452 (N_5452,N_3651,N_3942);
and U5453 (N_5453,N_2197,N_4895);
and U5454 (N_5454,N_314,N_3906);
xor U5455 (N_5455,N_4724,N_395);
nor U5456 (N_5456,N_2606,N_1732);
nor U5457 (N_5457,N_3334,N_281);
nand U5458 (N_5458,N_3604,N_3023);
and U5459 (N_5459,N_4570,N_4521);
nor U5460 (N_5460,N_3791,N_695);
and U5461 (N_5461,N_2207,N_60);
nor U5462 (N_5462,N_1726,N_1395);
nand U5463 (N_5463,N_1930,N_837);
and U5464 (N_5464,N_2639,N_4554);
or U5465 (N_5465,N_98,N_1874);
nand U5466 (N_5466,N_2644,N_805);
or U5467 (N_5467,N_2346,N_3946);
nor U5468 (N_5468,N_4756,N_4088);
nand U5469 (N_5469,N_2165,N_2757);
and U5470 (N_5470,N_4624,N_4308);
xor U5471 (N_5471,N_3909,N_1605);
and U5472 (N_5472,N_2489,N_467);
nand U5473 (N_5473,N_2242,N_1431);
nand U5474 (N_5474,N_4058,N_4152);
nor U5475 (N_5475,N_2423,N_541);
and U5476 (N_5476,N_1157,N_3388);
nand U5477 (N_5477,N_1058,N_1564);
or U5478 (N_5478,N_3046,N_2769);
xor U5479 (N_5479,N_3083,N_4078);
and U5480 (N_5480,N_2873,N_1752);
nor U5481 (N_5481,N_339,N_990);
nor U5482 (N_5482,N_2529,N_2507);
or U5483 (N_5483,N_2366,N_2869);
xnor U5484 (N_5484,N_340,N_2803);
or U5485 (N_5485,N_1066,N_2822);
and U5486 (N_5486,N_1808,N_812);
nor U5487 (N_5487,N_3573,N_732);
or U5488 (N_5488,N_3089,N_4817);
nor U5489 (N_5489,N_4145,N_347);
nand U5490 (N_5490,N_4368,N_4905);
or U5491 (N_5491,N_2223,N_598);
and U5492 (N_5492,N_4918,N_3410);
xnor U5493 (N_5493,N_4557,N_1383);
or U5494 (N_5494,N_4390,N_2395);
and U5495 (N_5495,N_950,N_3581);
xor U5496 (N_5496,N_2353,N_3674);
or U5497 (N_5497,N_3347,N_1517);
or U5498 (N_5498,N_1108,N_3664);
nand U5499 (N_5499,N_1055,N_1427);
nor U5500 (N_5500,N_2137,N_3506);
or U5501 (N_5501,N_375,N_4810);
and U5502 (N_5502,N_1562,N_4331);
or U5503 (N_5503,N_2515,N_3584);
nand U5504 (N_5504,N_3022,N_1173);
nor U5505 (N_5505,N_1450,N_3343);
nor U5506 (N_5506,N_4467,N_303);
nand U5507 (N_5507,N_1470,N_264);
nand U5508 (N_5508,N_2858,N_1996);
and U5509 (N_5509,N_762,N_1125);
and U5510 (N_5510,N_1698,N_4944);
and U5511 (N_5511,N_3079,N_4370);
nor U5512 (N_5512,N_3949,N_99);
and U5513 (N_5513,N_2443,N_4659);
xor U5514 (N_5514,N_4956,N_1420);
nand U5515 (N_5515,N_683,N_4183);
or U5516 (N_5516,N_4276,N_820);
or U5517 (N_5517,N_3214,N_2987);
nor U5518 (N_5518,N_1200,N_2267);
or U5519 (N_5519,N_788,N_454);
nor U5520 (N_5520,N_3629,N_35);
and U5521 (N_5521,N_1478,N_1870);
nor U5522 (N_5522,N_2561,N_1014);
nor U5523 (N_5523,N_2396,N_1667);
and U5524 (N_5524,N_2979,N_4179);
nand U5525 (N_5525,N_4782,N_2503);
and U5526 (N_5526,N_1225,N_2581);
xor U5527 (N_5527,N_2590,N_4236);
nand U5528 (N_5528,N_2328,N_4938);
or U5529 (N_5529,N_1132,N_474);
or U5530 (N_5530,N_2415,N_1594);
or U5531 (N_5531,N_2040,N_2728);
nand U5532 (N_5532,N_2941,N_167);
and U5533 (N_5533,N_760,N_3325);
and U5534 (N_5534,N_483,N_2670);
nand U5535 (N_5535,N_741,N_1086);
or U5536 (N_5536,N_883,N_3058);
nand U5537 (N_5537,N_3804,N_3027);
or U5538 (N_5538,N_887,N_953);
nand U5539 (N_5539,N_2138,N_963);
nor U5540 (N_5540,N_1012,N_1273);
nand U5541 (N_5541,N_4932,N_3734);
or U5542 (N_5542,N_4185,N_450);
nor U5543 (N_5543,N_480,N_2524);
or U5544 (N_5544,N_3481,N_444);
or U5545 (N_5545,N_463,N_49);
xnor U5546 (N_5546,N_1795,N_4548);
nand U5547 (N_5547,N_4232,N_1504);
and U5548 (N_5548,N_2398,N_1358);
nor U5549 (N_5549,N_3943,N_4593);
nor U5550 (N_5550,N_4023,N_1235);
or U5551 (N_5551,N_3419,N_1593);
and U5552 (N_5552,N_1480,N_4881);
nand U5553 (N_5553,N_1762,N_2158);
and U5554 (N_5554,N_3830,N_4873);
nor U5555 (N_5555,N_3402,N_3591);
xor U5556 (N_5556,N_4587,N_4705);
nand U5557 (N_5557,N_3808,N_4340);
or U5558 (N_5558,N_1165,N_4549);
nor U5559 (N_5559,N_462,N_1067);
and U5560 (N_5560,N_3543,N_94);
nand U5561 (N_5561,N_2808,N_4640);
or U5562 (N_5562,N_4616,N_4721);
and U5563 (N_5563,N_4507,N_2841);
nand U5564 (N_5564,N_3256,N_3004);
and U5565 (N_5565,N_2249,N_1328);
nor U5566 (N_5566,N_2496,N_818);
and U5567 (N_5567,N_1029,N_876);
nor U5568 (N_5568,N_222,N_307);
nor U5569 (N_5569,N_1319,N_266);
or U5570 (N_5570,N_911,N_1914);
and U5571 (N_5571,N_3181,N_1921);
nand U5572 (N_5572,N_4980,N_4971);
or U5573 (N_5573,N_3759,N_2289);
and U5574 (N_5574,N_627,N_4638);
nand U5575 (N_5575,N_1033,N_404);
and U5576 (N_5576,N_3202,N_3227);
xnor U5577 (N_5577,N_2856,N_4011);
and U5578 (N_5578,N_3927,N_4175);
and U5579 (N_5579,N_2058,N_3163);
nor U5580 (N_5580,N_476,N_55);
or U5581 (N_5581,N_3076,N_2832);
or U5582 (N_5582,N_1429,N_3536);
nand U5583 (N_5583,N_548,N_4685);
nand U5584 (N_5584,N_2228,N_4960);
or U5585 (N_5585,N_275,N_4983);
and U5586 (N_5586,N_1002,N_3098);
and U5587 (N_5587,N_2407,N_2131);
and U5588 (N_5588,N_1063,N_4768);
nand U5589 (N_5589,N_4173,N_3132);
nor U5590 (N_5590,N_3686,N_4989);
xor U5591 (N_5591,N_4652,N_19);
nor U5592 (N_5592,N_42,N_268);
nor U5593 (N_5593,N_3541,N_3072);
and U5594 (N_5594,N_2344,N_1674);
nand U5595 (N_5595,N_2215,N_4381);
nand U5596 (N_5596,N_4131,N_2892);
nand U5597 (N_5597,N_4633,N_3445);
and U5598 (N_5598,N_3241,N_4113);
and U5599 (N_5599,N_1582,N_3418);
nor U5600 (N_5600,N_4121,N_1342);
or U5601 (N_5601,N_2337,N_258);
or U5602 (N_5602,N_2419,N_4032);
nand U5603 (N_5603,N_400,N_1662);
or U5604 (N_5604,N_1436,N_1805);
or U5605 (N_5605,N_1192,N_1849);
or U5606 (N_5606,N_3468,N_3423);
or U5607 (N_5607,N_2492,N_3531);
nand U5608 (N_5608,N_2666,N_514);
or U5609 (N_5609,N_3208,N_1410);
nand U5610 (N_5610,N_3198,N_1144);
and U5611 (N_5611,N_2001,N_869);
nand U5612 (N_5612,N_4867,N_4455);
nor U5613 (N_5613,N_1057,N_3928);
or U5614 (N_5614,N_2772,N_4796);
and U5615 (N_5615,N_2950,N_4007);
nand U5616 (N_5616,N_2149,N_4414);
nor U5617 (N_5617,N_3124,N_1247);
nand U5618 (N_5618,N_4757,N_3297);
nor U5619 (N_5619,N_3363,N_2179);
nand U5620 (N_5620,N_868,N_3259);
nand U5621 (N_5621,N_4383,N_804);
or U5622 (N_5622,N_3391,N_59);
nor U5623 (N_5623,N_2701,N_1248);
and U5624 (N_5624,N_595,N_4292);
or U5625 (N_5625,N_3740,N_1791);
or U5626 (N_5626,N_3971,N_2726);
and U5627 (N_5627,N_1655,N_2886);
nor U5628 (N_5628,N_493,N_681);
nand U5629 (N_5629,N_4432,N_813);
and U5630 (N_5630,N_1730,N_3);
and U5631 (N_5631,N_1404,N_1768);
nor U5632 (N_5632,N_4831,N_1325);
and U5633 (N_5633,N_4195,N_4739);
and U5634 (N_5634,N_4577,N_904);
and U5635 (N_5635,N_193,N_601);
nand U5636 (N_5636,N_2283,N_2350);
and U5637 (N_5637,N_3986,N_1656);
or U5638 (N_5638,N_3366,N_4213);
or U5639 (N_5639,N_3075,N_2689);
or U5640 (N_5640,N_2568,N_2734);
xnor U5641 (N_5641,N_2285,N_3754);
xor U5642 (N_5642,N_155,N_1976);
nor U5643 (N_5643,N_2500,N_2408);
or U5644 (N_5644,N_4319,N_1380);
nand U5645 (N_5645,N_2499,N_2314);
or U5646 (N_5646,N_586,N_2232);
or U5647 (N_5647,N_4936,N_377);
nand U5648 (N_5648,N_2342,N_4199);
xnor U5649 (N_5649,N_4500,N_4673);
nand U5650 (N_5650,N_2009,N_142);
nand U5651 (N_5651,N_4778,N_4068);
or U5652 (N_5652,N_4910,N_2089);
and U5653 (N_5653,N_1696,N_2862);
or U5654 (N_5654,N_273,N_4483);
or U5655 (N_5655,N_342,N_152);
nor U5656 (N_5656,N_3825,N_4150);
nor U5657 (N_5657,N_3559,N_1214);
nand U5658 (N_5658,N_3693,N_2742);
xor U5659 (N_5659,N_513,N_3215);
nand U5660 (N_5660,N_428,N_2860);
nand U5661 (N_5661,N_3890,N_1196);
or U5662 (N_5662,N_3450,N_3356);
xnor U5663 (N_5663,N_4835,N_4315);
and U5664 (N_5664,N_4657,N_3774);
nor U5665 (N_5665,N_3951,N_3034);
nand U5666 (N_5666,N_1995,N_2471);
or U5667 (N_5667,N_4731,N_862);
xnor U5668 (N_5668,N_884,N_2692);
nand U5669 (N_5669,N_2572,N_1381);
nor U5670 (N_5670,N_621,N_2204);
and U5671 (N_5671,N_500,N_3143);
or U5672 (N_5672,N_2329,N_4764);
and U5673 (N_5673,N_1495,N_441);
xnor U5674 (N_5674,N_2251,N_2063);
nand U5675 (N_5675,N_3218,N_3698);
xor U5676 (N_5676,N_2291,N_2537);
or U5677 (N_5677,N_1206,N_1796);
or U5678 (N_5678,N_1308,N_4903);
or U5679 (N_5679,N_901,N_22);
or U5680 (N_5680,N_494,N_3991);
and U5681 (N_5681,N_1080,N_498);
or U5682 (N_5682,N_4338,N_3669);
nand U5683 (N_5683,N_1371,N_4137);
xnor U5684 (N_5684,N_2261,N_3966);
and U5685 (N_5685,N_1484,N_100);
and U5686 (N_5686,N_3886,N_3910);
and U5687 (N_5687,N_486,N_2482);
nor U5688 (N_5688,N_1453,N_2360);
nor U5689 (N_5689,N_1186,N_1324);
and U5690 (N_5690,N_1185,N_497);
nor U5691 (N_5691,N_3273,N_2447);
or U5692 (N_5692,N_3939,N_1496);
nand U5693 (N_5693,N_1664,N_4563);
nand U5694 (N_5694,N_373,N_1536);
nand U5695 (N_5695,N_3510,N_358);
xor U5696 (N_5696,N_3160,N_2270);
and U5697 (N_5697,N_1728,N_398);
nand U5698 (N_5698,N_1056,N_2934);
nand U5699 (N_5699,N_709,N_3787);
nor U5700 (N_5700,N_2939,N_528);
nor U5701 (N_5701,N_424,N_3311);
nor U5702 (N_5702,N_51,N_257);
and U5703 (N_5703,N_15,N_4235);
and U5704 (N_5704,N_393,N_1332);
nor U5705 (N_5705,N_1897,N_2047);
or U5706 (N_5706,N_2255,N_93);
xnor U5707 (N_5707,N_3401,N_2099);
nand U5708 (N_5708,N_3249,N_1399);
xnor U5709 (N_5709,N_3678,N_82);
or U5710 (N_5710,N_2352,N_4016);
and U5711 (N_5711,N_981,N_3434);
nand U5712 (N_5712,N_1303,N_227);
or U5713 (N_5713,N_301,N_382);
nand U5714 (N_5714,N_2918,N_543);
nor U5715 (N_5715,N_1649,N_4259);
and U5716 (N_5716,N_4880,N_1296);
and U5717 (N_5717,N_359,N_1113);
nor U5718 (N_5718,N_1873,N_3199);
nor U5719 (N_5719,N_4033,N_2233);
nor U5720 (N_5720,N_3421,N_4510);
and U5721 (N_5721,N_1398,N_3766);
and U5722 (N_5722,N_2849,N_4608);
and U5723 (N_5723,N_2383,N_1771);
nor U5724 (N_5724,N_1597,N_4401);
nor U5725 (N_5725,N_1744,N_3790);
nand U5726 (N_5726,N_1202,N_3652);
nor U5727 (N_5727,N_947,N_2682);
xnor U5728 (N_5728,N_3064,N_4818);
and U5729 (N_5729,N_2617,N_4846);
nor U5730 (N_5730,N_4805,N_194);
and U5731 (N_5731,N_3871,N_4082);
xnor U5732 (N_5732,N_4564,N_1259);
and U5733 (N_5733,N_45,N_2154);
xor U5734 (N_5734,N_4375,N_827);
or U5735 (N_5735,N_3550,N_2284);
nor U5736 (N_5736,N_1793,N_3289);
or U5737 (N_5737,N_4891,N_2630);
nand U5738 (N_5738,N_1853,N_2172);
xor U5739 (N_5739,N_2295,N_2954);
xnor U5740 (N_5740,N_1623,N_2010);
nand U5741 (N_5741,N_1865,N_2117);
or U5742 (N_5742,N_3661,N_112);
nor U5743 (N_5743,N_982,N_1391);
nor U5744 (N_5744,N_1280,N_3280);
nand U5745 (N_5745,N_4968,N_596);
nand U5746 (N_5746,N_2414,N_4478);
xor U5747 (N_5747,N_4987,N_4475);
nor U5748 (N_5748,N_3833,N_1703);
xor U5749 (N_5749,N_2916,N_2469);
and U5750 (N_5750,N_1085,N_3688);
nor U5751 (N_5751,N_330,N_505);
nand U5752 (N_5752,N_1804,N_897);
or U5753 (N_5753,N_1746,N_4227);
and U5754 (N_5754,N_1966,N_4809);
nand U5755 (N_5755,N_4172,N_2491);
and U5756 (N_5756,N_4779,N_2614);
xor U5757 (N_5757,N_2318,N_334);
nand U5758 (N_5758,N_390,N_4783);
nor U5759 (N_5759,N_3989,N_1121);
or U5760 (N_5760,N_3341,N_1030);
nand U5761 (N_5761,N_4050,N_3429);
nor U5762 (N_5762,N_3978,N_1497);
or U5763 (N_5763,N_4343,N_1251);
xor U5764 (N_5764,N_2406,N_2317);
or U5765 (N_5765,N_3119,N_4039);
nand U5766 (N_5766,N_2605,N_3647);
nor U5767 (N_5767,N_1435,N_3996);
or U5768 (N_5768,N_3812,N_3310);
nor U5769 (N_5769,N_3300,N_3888);
nor U5770 (N_5770,N_2112,N_4814);
nand U5771 (N_5771,N_1331,N_2030);
xor U5772 (N_5772,N_1673,N_1076);
nand U5773 (N_5773,N_846,N_605);
and U5774 (N_5774,N_3500,N_3977);
nor U5775 (N_5775,N_4325,N_3488);
nand U5776 (N_5776,N_3081,N_2960);
nand U5777 (N_5777,N_321,N_2453);
and U5778 (N_5778,N_3853,N_3107);
xnor U5779 (N_5779,N_2770,N_952);
xor U5780 (N_5780,N_389,N_1596);
and U5781 (N_5781,N_4603,N_3224);
nor U5782 (N_5782,N_3508,N_3200);
nand U5783 (N_5783,N_717,N_3765);
or U5784 (N_5784,N_4169,N_4806);
nor U5785 (N_5785,N_1461,N_520);
nand U5786 (N_5786,N_242,N_1106);
and U5787 (N_5787,N_1375,N_2964);
or U5788 (N_5788,N_2327,N_771);
and U5789 (N_5789,N_2111,N_2474);
nor U5790 (N_5790,N_2830,N_87);
and U5791 (N_5791,N_3789,N_4306);
xor U5792 (N_5792,N_694,N_3490);
nand U5793 (N_5793,N_1048,N_2798);
nand U5794 (N_5794,N_3921,N_3033);
nand U5795 (N_5795,N_940,N_352);
nand U5796 (N_5796,N_3561,N_579);
nor U5797 (N_5797,N_954,N_929);
nand U5798 (N_5798,N_4201,N_4927);
nor U5799 (N_5799,N_809,N_1787);
and U5800 (N_5800,N_2972,N_4044);
or U5801 (N_5801,N_2430,N_3438);
and U5802 (N_5802,N_1672,N_1064);
nor U5803 (N_5803,N_38,N_4367);
nor U5804 (N_5804,N_3801,N_2404);
and U5805 (N_5805,N_1487,N_3841);
or U5806 (N_5806,N_4275,N_2025);
and U5807 (N_5807,N_4209,N_249);
or U5808 (N_5808,N_1474,N_4794);
nand U5809 (N_5809,N_4561,N_2502);
nor U5810 (N_5810,N_4360,N_33);
nand U5811 (N_5811,N_2551,N_187);
nor U5812 (N_5812,N_3211,N_2075);
nand U5813 (N_5813,N_364,N_3512);
or U5814 (N_5814,N_1022,N_1180);
nor U5815 (N_5815,N_2615,N_3563);
nand U5816 (N_5816,N_4763,N_1844);
or U5817 (N_5817,N_216,N_2991);
nor U5818 (N_5818,N_729,N_1079);
nand U5819 (N_5819,N_857,N_4328);
nand U5820 (N_5820,N_2871,N_8);
nand U5821 (N_5821,N_4840,N_2573);
nor U5822 (N_5822,N_119,N_4553);
and U5823 (N_5823,N_1931,N_1050);
nor U5824 (N_5824,N_1892,N_311);
xnor U5825 (N_5825,N_773,N_2744);
nor U5826 (N_5826,N_4189,N_335);
nand U5827 (N_5827,N_4140,N_4501);
xnor U5828 (N_5828,N_1156,N_975);
and U5829 (N_5829,N_4573,N_2711);
xnor U5830 (N_5830,N_3415,N_3479);
nor U5831 (N_5831,N_1112,N_2998);
xor U5832 (N_5832,N_3061,N_2667);
nor U5833 (N_5833,N_3221,N_2512);
and U5834 (N_5834,N_4872,N_2668);
or U5835 (N_5835,N_1616,N_3861);
or U5836 (N_5836,N_2409,N_3469);
nor U5837 (N_5837,N_1939,N_3278);
nand U5838 (N_5838,N_3819,N_1001);
and U5839 (N_5839,N_3907,N_2427);
nor U5840 (N_5840,N_531,N_919);
nand U5841 (N_5841,N_3255,N_36);
xnor U5842 (N_5842,N_4575,N_971);
nor U5843 (N_5843,N_3884,N_1345);
nor U5844 (N_5844,N_2758,N_965);
and U5845 (N_5845,N_4254,N_4843);
and U5846 (N_5846,N_1230,N_316);
nand U5847 (N_5847,N_2982,N_392);
nor U5848 (N_5848,N_1339,N_158);
and U5849 (N_5849,N_2281,N_1340);
nor U5850 (N_5850,N_3011,N_4602);
and U5851 (N_5851,N_2616,N_765);
nor U5852 (N_5852,N_4043,N_2128);
nand U5853 (N_5853,N_4645,N_2118);
or U5854 (N_5854,N_3663,N_552);
or U5855 (N_5855,N_4061,N_4035);
or U5856 (N_5856,N_30,N_65);
or U5857 (N_5857,N_2526,N_2875);
nand U5858 (N_5858,N_3068,N_3213);
and U5859 (N_5859,N_2088,N_2624);
nor U5860 (N_5860,N_2791,N_2716);
nand U5861 (N_5861,N_3008,N_1981);
nand U5862 (N_5862,N_4821,N_4569);
nand U5863 (N_5863,N_3956,N_4466);
nand U5864 (N_5864,N_4372,N_2766);
xor U5865 (N_5865,N_3448,N_2120);
nor U5866 (N_5866,N_4807,N_900);
or U5867 (N_5867,N_2288,N_3753);
and U5868 (N_5868,N_138,N_2664);
and U5869 (N_5869,N_2240,N_1032);
or U5870 (N_5870,N_3845,N_3242);
xor U5871 (N_5871,N_934,N_3216);
and U5872 (N_5872,N_3416,N_2193);
or U5873 (N_5873,N_1544,N_3649);
and U5874 (N_5874,N_3066,N_299);
nor U5875 (N_5875,N_2521,N_4538);
and U5876 (N_5876,N_4664,N_4305);
and U5877 (N_5877,N_374,N_1258);
xnor U5878 (N_5878,N_4093,N_1532);
and U5879 (N_5879,N_4277,N_3285);
nand U5880 (N_5880,N_1405,N_3641);
xnor U5881 (N_5881,N_2971,N_610);
nand U5882 (N_5882,N_399,N_677);
nor U5883 (N_5883,N_1141,N_3494);
nor U5884 (N_5884,N_2720,N_2326);
and U5885 (N_5885,N_936,N_3795);
or U5886 (N_5886,N_402,N_1356);
nor U5887 (N_5887,N_3666,N_1934);
and U5888 (N_5888,N_4613,N_302);
nor U5889 (N_5889,N_636,N_1862);
nand U5890 (N_5890,N_4857,N_2339);
and U5891 (N_5891,N_3611,N_3453);
and U5892 (N_5892,N_1848,N_4709);
nand U5893 (N_5893,N_3230,N_160);
nor U5894 (N_5894,N_2698,N_4454);
nor U5895 (N_5895,N_2913,N_980);
nand U5896 (N_5896,N_4589,N_4298);
or U5897 (N_5897,N_1253,N_4477);
or U5898 (N_5898,N_2347,N_2776);
nand U5899 (N_5899,N_1464,N_3063);
and U5900 (N_5900,N_3495,N_1611);
and U5901 (N_5901,N_2123,N_802);
nor U5902 (N_5902,N_3839,N_4314);
nand U5903 (N_5903,N_3465,N_873);
nor U5904 (N_5904,N_556,N_137);
nand U5905 (N_5905,N_738,N_4075);
nor U5906 (N_5906,N_2403,N_1406);
or U5907 (N_5907,N_1152,N_1114);
nor U5908 (N_5908,N_3138,N_3635);
or U5909 (N_5909,N_1189,N_1701);
and U5910 (N_5910,N_1887,N_1351);
nand U5911 (N_5911,N_1603,N_1555);
nor U5912 (N_5912,N_421,N_58);
xor U5913 (N_5913,N_3062,N_3542);
or U5914 (N_5914,N_4079,N_1494);
nor U5915 (N_5915,N_2455,N_4599);
and U5916 (N_5916,N_938,N_3630);
nand U5917 (N_5917,N_3191,N_4811);
nand U5918 (N_5918,N_3294,N_1101);
nand U5919 (N_5919,N_1183,N_1871);
nor U5920 (N_5920,N_415,N_1004);
nor U5921 (N_5921,N_4464,N_380);
nor U5922 (N_5922,N_4335,N_4064);
or U5923 (N_5923,N_4676,N_4733);
xor U5924 (N_5924,N_4098,N_3196);
and U5925 (N_5925,N_4545,N_269);
nor U5926 (N_5926,N_4222,N_2990);
or U5927 (N_5927,N_4815,N_2199);
nand U5928 (N_5928,N_4504,N_1661);
nand U5929 (N_5929,N_542,N_4036);
nand U5930 (N_5930,N_4648,N_1147);
xnor U5931 (N_5931,N_1621,N_3185);
and U5932 (N_5932,N_4883,N_1330);
nor U5933 (N_5933,N_1660,N_1942);
and U5934 (N_5934,N_1606,N_2876);
or U5935 (N_5935,N_4830,N_4376);
nand U5936 (N_5936,N_470,N_200);
nand U5937 (N_5937,N_1341,N_1139);
xor U5938 (N_5938,N_2436,N_3703);
nand U5939 (N_5939,N_3858,N_2680);
xnor U5940 (N_5940,N_4495,N_2710);
or U5941 (N_5941,N_2239,N_417);
nor U5942 (N_5942,N_163,N_2079);
and U5943 (N_5943,N_1133,N_1350);
or U5944 (N_5944,N_1964,N_864);
nor U5945 (N_5945,N_3665,N_3209);
and U5946 (N_5946,N_3822,N_4686);
or U5947 (N_5947,N_4097,N_4958);
xnor U5948 (N_5948,N_4924,N_4387);
or U5949 (N_5949,N_1573,N_2671);
nand U5950 (N_5950,N_2341,N_4482);
xor U5951 (N_5951,N_3657,N_4337);
and U5952 (N_5952,N_4188,N_1007);
nor U5953 (N_5953,N_1400,N_4994);
or U5954 (N_5954,N_2878,N_2434);
nand U5955 (N_5955,N_4202,N_4832);
or U5956 (N_5956,N_1908,N_1254);
and U5957 (N_5957,N_4133,N_2678);
nand U5958 (N_5958,N_2908,N_3487);
or U5959 (N_5959,N_4834,N_675);
nand U5960 (N_5960,N_653,N_2202);
or U5961 (N_5961,N_3462,N_3454);
and U5962 (N_5962,N_1423,N_4056);
nor U5963 (N_5963,N_3518,N_209);
and U5964 (N_5964,N_3614,N_148);
nor U5965 (N_5965,N_1572,N_1204);
or U5966 (N_5966,N_1437,N_1919);
nor U5967 (N_5967,N_3474,N_2665);
or U5968 (N_5968,N_1823,N_3084);
and U5969 (N_5969,N_21,N_2292);
nand U5970 (N_5970,N_4862,N_2411);
nand U5971 (N_5971,N_1411,N_1801);
nor U5972 (N_5972,N_4797,N_4984);
and U5973 (N_5973,N_391,N_448);
or U5974 (N_5974,N_1181,N_1146);
and U5975 (N_5975,N_1546,N_3032);
or U5976 (N_5976,N_4894,N_2357);
and U5977 (N_5977,N_414,N_973);
nor U5978 (N_5978,N_4302,N_4861);
nor U5979 (N_5979,N_591,N_3491);
or U5980 (N_5980,N_2189,N_3866);
nor U5981 (N_5981,N_265,N_25);
or U5982 (N_5982,N_2272,N_1917);
and U5983 (N_5983,N_376,N_515);
and U5984 (N_5984,N_1236,N_2893);
nand U5985 (N_5985,N_3339,N_527);
or U5986 (N_5986,N_3136,N_1197);
nand U5987 (N_5987,N_1753,N_1093);
or U5988 (N_5988,N_3439,N_899);
or U5989 (N_5989,N_3254,N_3400);
and U5990 (N_5990,N_1622,N_4758);
or U5991 (N_5991,N_2245,N_108);
or U5992 (N_5992,N_3477,N_3623);
nand U5993 (N_5993,N_1717,N_111);
nand U5994 (N_5994,N_4490,N_381);
and U5995 (N_5995,N_3283,N_2902);
and U5996 (N_5996,N_215,N_2545);
xnor U5997 (N_5997,N_3889,N_2134);
and U5998 (N_5998,N_2727,N_3364);
and U5999 (N_5999,N_4369,N_4610);
xnor U6000 (N_6000,N_3950,N_1268);
or U6001 (N_6001,N_2083,N_422);
nor U6002 (N_6002,N_4838,N_46);
nor U6003 (N_6003,N_4219,N_759);
and U6004 (N_6004,N_1402,N_2280);
and U6005 (N_6005,N_2180,N_2591);
nand U6006 (N_6006,N_1610,N_2788);
nor U6007 (N_6007,N_1019,N_535);
xnor U6008 (N_6008,N_593,N_4374);
and U6009 (N_6009,N_3471,N_4484);
or U6010 (N_6010,N_458,N_2684);
nor U6011 (N_6011,N_4406,N_1316);
or U6012 (N_6012,N_2373,N_3622);
nand U6013 (N_6013,N_1354,N_3376);
or U6014 (N_6014,N_3849,N_3578);
or U6015 (N_6015,N_3940,N_1126);
or U6016 (N_6016,N_1700,N_916);
nand U6017 (N_6017,N_4262,N_4517);
or U6018 (N_6018,N_4067,N_1096);
or U6019 (N_6019,N_2931,N_487);
or U6020 (N_6020,N_1971,N_570);
nand U6021 (N_6021,N_987,N_3028);
or U6022 (N_6022,N_3836,N_1687);
nand U6023 (N_6023,N_1131,N_2575);
or U6024 (N_6024,N_73,N_3859);
or U6025 (N_6025,N_2944,N_958);
and U6026 (N_6026,N_4261,N_3458);
nor U6027 (N_6027,N_1773,N_2566);
nor U6028 (N_6028,N_972,N_1169);
nand U6029 (N_6029,N_612,N_89);
xor U6030 (N_6030,N_815,N_171);
nand U6031 (N_6031,N_3739,N_4115);
and U6032 (N_6032,N_1090,N_1935);
and U6033 (N_6033,N_2477,N_2904);
and U6034 (N_6034,N_2848,N_910);
xnor U6035 (N_6035,N_1905,N_4574);
and U6036 (N_6036,N_1881,N_1110);
nor U6037 (N_6037,N_1909,N_3627);
nand U6038 (N_6038,N_2777,N_1122);
nor U6039 (N_6039,N_4625,N_2321);
or U6040 (N_6040,N_4136,N_4240);
xor U6041 (N_6041,N_850,N_244);
xnor U6042 (N_6042,N_1520,N_3857);
and U6043 (N_6043,N_3838,N_2429);
and U6044 (N_6044,N_2852,N_313);
nand U6045 (N_6045,N_4072,N_2708);
xnor U6046 (N_6046,N_260,N_2596);
and U6047 (N_6047,N_3997,N_4423);
xnor U6048 (N_6048,N_3694,N_2926);
or U6049 (N_6049,N_4742,N_2816);
and U6050 (N_6050,N_69,N_908);
nor U6051 (N_6051,N_4703,N_56);
nand U6052 (N_6052,N_1587,N_2618);
nor U6053 (N_6053,N_1583,N_4530);
nor U6054 (N_6054,N_1620,N_4005);
nor U6055 (N_6055,N_2585,N_4774);
or U6056 (N_6056,N_726,N_4243);
and U6057 (N_6057,N_2313,N_1044);
and U6058 (N_6058,N_1608,N_2525);
and U6059 (N_6059,N_2637,N_1833);
xor U6060 (N_6060,N_3346,N_889);
and U6061 (N_6061,N_891,N_1712);
nand U6062 (N_6062,N_671,N_3988);
or U6063 (N_6063,N_4637,N_2985);
and U6064 (N_6064,N_2586,N_1407);
nor U6065 (N_6065,N_2764,N_4556);
or U6066 (N_6066,N_655,N_3676);
xor U6067 (N_6067,N_384,N_4679);
nor U6068 (N_6068,N_4771,N_1175);
nand U6069 (N_6069,N_288,N_3945);
or U6070 (N_6070,N_4018,N_3470);
nor U6071 (N_6071,N_4135,N_907);
nand U6072 (N_6072,N_1293,N_1194);
and U6073 (N_6073,N_3186,N_1772);
nand U6074 (N_6074,N_4291,N_985);
nand U6075 (N_6075,N_4457,N_4666);
nor U6076 (N_6076,N_4753,N_3891);
nor U6077 (N_6077,N_4860,N_1988);
or U6078 (N_6078,N_3247,N_888);
nand U6079 (N_6079,N_4639,N_1285);
nand U6080 (N_6080,N_2457,N_2505);
and U6081 (N_6081,N_4722,N_545);
and U6082 (N_6082,N_3603,N_344);
nand U6083 (N_6083,N_1845,N_1972);
or U6084 (N_6084,N_2534,N_323);
nand U6085 (N_6085,N_1683,N_823);
xnor U6086 (N_6086,N_4623,N_667);
xnor U6087 (N_6087,N_1384,N_4916);
and U6088 (N_6088,N_1439,N_3505);
or U6089 (N_6089,N_4781,N_1249);
xor U6090 (N_6090,N_4287,N_2957);
nor U6091 (N_6091,N_310,N_4013);
nand U6092 (N_6092,N_696,N_4665);
xor U6093 (N_6093,N_246,N_3842);
nor U6094 (N_6094,N_1827,N_4433);
or U6095 (N_6095,N_4738,N_3913);
nand U6096 (N_6096,N_3507,N_1570);
or U6097 (N_6097,N_3105,N_2162);
nand U6098 (N_6098,N_3756,N_4408);
or U6099 (N_6099,N_3301,N_1551);
xnor U6100 (N_6100,N_3037,N_1203);
or U6101 (N_6101,N_1774,N_4318);
or U6102 (N_6102,N_4208,N_3074);
nand U6103 (N_6103,N_451,N_1947);
and U6104 (N_6104,N_4727,N_3441);
nor U6105 (N_6105,N_3135,N_4270);
and U6106 (N_6106,N_2709,N_90);
nand U6107 (N_6107,N_1568,N_174);
nand U6108 (N_6108,N_2143,N_1689);
and U6109 (N_6109,N_1922,N_1759);
or U6110 (N_6110,N_491,N_4948);
nand U6111 (N_6111,N_1557,N_1575);
nor U6112 (N_6112,N_4225,N_3044);
or U6113 (N_6113,N_2116,N_2730);
nor U6114 (N_6114,N_4431,N_3720);
nor U6115 (N_6115,N_3287,N_2802);
and U6116 (N_6116,N_115,N_3608);
and U6117 (N_6117,N_432,N_1269);
nor U6118 (N_6118,N_1069,N_3699);
and U6119 (N_6119,N_4559,N_3337);
xnor U6120 (N_6120,N_4239,N_2704);
nor U6121 (N_6121,N_489,N_4154);
xnor U6122 (N_6122,N_4726,N_2844);
and U6123 (N_6123,N_4029,N_1068);
nand U6124 (N_6124,N_3226,N_1160);
nor U6125 (N_6125,N_425,N_2444);
and U6126 (N_6126,N_2051,N_177);
and U6127 (N_6127,N_369,N_3368);
nand U6128 (N_6128,N_2965,N_1088);
nor U6129 (N_6129,N_459,N_1127);
or U6130 (N_6130,N_955,N_662);
nand U6131 (N_6131,N_4520,N_2190);
nor U6132 (N_6132,N_2801,N_2276);
and U6133 (N_6133,N_4045,N_224);
nor U6134 (N_6134,N_3047,N_4576);
and U6135 (N_6135,N_3045,N_727);
or U6136 (N_6136,N_1207,N_1433);
or U6137 (N_6137,N_2343,N_3532);
xor U6138 (N_6138,N_2601,N_172);
xnor U6139 (N_6139,N_3304,N_3687);
nand U6140 (N_6140,N_534,N_2250);
and U6141 (N_6141,N_1738,N_2187);
and U6142 (N_6142,N_966,N_3732);
nor U6143 (N_6143,N_211,N_2792);
and U6144 (N_6144,N_4799,N_2388);
or U6145 (N_6145,N_4054,N_3746);
xor U6146 (N_6146,N_1492,N_4410);
or U6147 (N_6147,N_3296,N_3722);
nor U6148 (N_6148,N_2656,N_3307);
or U6149 (N_6149,N_1637,N_3755);
nor U6150 (N_6150,N_1075,N_1243);
or U6151 (N_6151,N_3667,N_1750);
xor U6152 (N_6152,N_1643,N_4107);
or U6153 (N_6153,N_3150,N_1162);
or U6154 (N_6154,N_1116,N_1336);
nor U6155 (N_6155,N_4405,N_2675);
or U6156 (N_6156,N_1749,N_2460);
xor U6157 (N_6157,N_2061,N_2311);
or U6158 (N_6158,N_3203,N_1757);
or U6159 (N_6159,N_640,N_4765);
or U6160 (N_6160,N_4629,N_921);
nor U6161 (N_6161,N_2023,N_2150);
xnor U6162 (N_6162,N_3577,N_3644);
nand U6163 (N_6163,N_3798,N_4231);
nand U6164 (N_6164,N_4224,N_254);
or U6165 (N_6165,N_4290,N_4822);
and U6166 (N_6166,N_4132,N_57);
or U6167 (N_6167,N_2003,N_2700);
or U6168 (N_6168,N_4524,N_4151);
and U6169 (N_6169,N_3261,N_1250);
and U6170 (N_6170,N_2186,N_2368);
or U6171 (N_6171,N_1916,N_1355);
nor U6172 (N_6172,N_1362,N_2956);
nor U6173 (N_6173,N_687,N_3960);
xnor U6174 (N_6174,N_699,N_1238);
xor U6175 (N_6175,N_915,N_4320);
and U6176 (N_6176,N_2103,N_1417);
and U6177 (N_6177,N_3646,N_2043);
nand U6178 (N_6178,N_2294,N_126);
or U6179 (N_6179,N_4885,N_1119);
and U6180 (N_6180,N_3874,N_3738);
nor U6181 (N_6181,N_4280,N_4158);
xnor U6182 (N_6182,N_3852,N_2473);
nand U6183 (N_6183,N_2535,N_4693);
nor U6184 (N_6184,N_784,N_3628);
nand U6185 (N_6185,N_4249,N_3979);
or U6186 (N_6186,N_2093,N_1828);
nand U6187 (N_6187,N_932,N_341);
nor U6188 (N_6188,N_3593,N_4714);
and U6189 (N_6189,N_4533,N_3353);
and U6190 (N_6190,N_2940,N_1632);
nand U6191 (N_6191,N_3271,N_4402);
nor U6192 (N_6192,N_509,N_388);
and U6193 (N_6193,N_1886,N_4901);
or U6194 (N_6194,N_285,N_1595);
or U6195 (N_6195,N_3511,N_150);
nand U6196 (N_6196,N_4492,N_637);
and U6197 (N_6197,N_3716,N_2697);
or U6198 (N_6198,N_4730,N_2041);
nor U6199 (N_6199,N_1071,N_2795);
or U6200 (N_6200,N_3779,N_4606);
nand U6201 (N_6201,N_2109,N_608);
and U6202 (N_6202,N_239,N_704);
and U6203 (N_6203,N_1794,N_122);
xnor U6204 (N_6204,N_1781,N_1713);
and U6205 (N_6205,N_4531,N_4584);
nor U6206 (N_6206,N_3883,N_2773);
or U6207 (N_6207,N_4988,N_27);
and U6208 (N_6208,N_4963,N_4786);
and U6209 (N_6209,N_3974,N_3018);
or U6210 (N_6210,N_4904,N_3409);
nor U6211 (N_6211,N_3467,N_4411);
or U6212 (N_6212,N_2933,N_3270);
xor U6213 (N_6213,N_2050,N_4972);
nor U6214 (N_6214,N_29,N_2225);
nand U6215 (N_6215,N_2105,N_4702);
nand U6216 (N_6216,N_4970,N_3700);
nand U6217 (N_6217,N_603,N_1896);
nor U6218 (N_6218,N_103,N_4630);
nand U6219 (N_6219,N_2046,N_1446);
nand U6220 (N_6220,N_4718,N_4379);
or U6221 (N_6221,N_4552,N_39);
or U6222 (N_6222,N_4282,N_1161);
and U6223 (N_6223,N_1691,N_866);
and U6224 (N_6224,N_3615,N_1822);
nand U6225 (N_6225,N_4386,N_2980);
or U6226 (N_6226,N_1501,N_3953);
and U6227 (N_6227,N_1224,N_583);
xnor U6228 (N_6228,N_508,N_3599);
or U6229 (N_6229,N_845,N_786);
nand U6230 (N_6230,N_3602,N_4820);
or U6231 (N_6231,N_3509,N_1266);
nand U6232 (N_6232,N_1547,N_597);
xnor U6233 (N_6233,N_157,N_4995);
and U6234 (N_6234,N_4200,N_1984);
or U6235 (N_6235,N_751,N_2796);
and U6236 (N_6236,N_670,N_3620);
xor U6237 (N_6237,N_507,N_3172);
xor U6238 (N_6238,N_2236,N_431);
and U6239 (N_6239,N_2989,N_917);
nand U6240 (N_6240,N_4186,N_1676);
nand U6241 (N_6241,N_2966,N_145);
and U6242 (N_6242,N_661,N_3424);
nor U6243 (N_6243,N_4770,N_1872);
xor U6244 (N_6244,N_2247,N_4741);
nand U6245 (N_6245,N_4017,N_4479);
nor U6246 (N_6246,N_2160,N_4981);
and U6247 (N_6247,N_994,N_3055);
nand U6248 (N_6248,N_394,N_3073);
and U6249 (N_6249,N_1279,N_3013);
or U6250 (N_6250,N_2501,N_4697);
and U6251 (N_6251,N_1508,N_3151);
nand U6252 (N_6252,N_2140,N_752);
nand U6253 (N_6253,N_2217,N_4926);
nand U6254 (N_6254,N_4435,N_4893);
nor U6255 (N_6255,N_3631,N_2380);
nand U6256 (N_6256,N_2522,N_3112);
xor U6257 (N_6257,N_468,N_3394);
and U6258 (N_6258,N_2552,N_4226);
and U6259 (N_6259,N_898,N_1283);
or U6260 (N_6260,N_4668,N_4122);
nor U6261 (N_6261,N_3308,N_3206);
nand U6262 (N_6262,N_2706,N_2622);
nand U6263 (N_6263,N_3783,N_2005);
and U6264 (N_6264,N_2576,N_189);
nand U6265 (N_6265,N_3332,N_3187);
nand U6266 (N_6266,N_3459,N_4532);
xnor U6267 (N_6267,N_2597,N_2905);
nand U6268 (N_6268,N_1505,N_948);
or U6269 (N_6269,N_614,N_2121);
nor U6270 (N_6270,N_3770,N_208);
nor U6271 (N_6271,N_2435,N_512);
nor U6272 (N_6272,N_2662,N_602);
and U6273 (N_6273,N_1878,N_4567);
nor U6274 (N_6274,N_1814,N_3313);
xor U6275 (N_6275,N_4256,N_4055);
nand U6276 (N_6276,N_4487,N_3020);
xnor U6277 (N_6277,N_2071,N_2577);
or U6278 (N_6278,N_935,N_2642);
nor U6279 (N_6279,N_855,N_4954);
or U6280 (N_6280,N_2016,N_4965);
nor U6281 (N_6281,N_2136,N_4710);
nand U6282 (N_6282,N_743,N_3564);
or U6283 (N_6283,N_3677,N_518);
nor U6284 (N_6284,N_1500,N_4992);
or U6285 (N_6285,N_2019,N_628);
nor U6286 (N_6286,N_430,N_1668);
or U6287 (N_6287,N_1016,N_4130);
nand U6288 (N_6288,N_3748,N_3231);
xnor U6289 (N_6289,N_141,N_2085);
or U6290 (N_6290,N_434,N_4544);
and U6291 (N_6291,N_3146,N_2176);
nor U6292 (N_6292,N_2098,N_2312);
nand U6293 (N_6293,N_2793,N_4156);
nand U6294 (N_6294,N_2951,N_3634);
xor U6295 (N_6295,N_4420,N_1401);
xor U6296 (N_6296,N_1275,N_154);
nor U6297 (N_6297,N_2306,N_4723);
and U6298 (N_6298,N_566,N_2679);
and U6299 (N_6299,N_2896,N_1911);
nor U6300 (N_6300,N_2487,N_1950);
or U6301 (N_6301,N_4683,N_3656);
nor U6302 (N_6302,N_2771,N_1300);
nor U6303 (N_6303,N_2080,N_3574);
xor U6304 (N_6304,N_1554,N_1242);
nand U6305 (N_6305,N_4692,N_1776);
or U6306 (N_6306,N_3553,N_631);
nand U6307 (N_6307,N_1387,N_3298);
or U6308 (N_6308,N_2520,N_996);
xor U6309 (N_6309,N_1457,N_2362);
nand U6310 (N_6310,N_1509,N_4307);
or U6311 (N_6311,N_1856,N_700);
and U6312 (N_6312,N_4795,N_251);
nor U6313 (N_6313,N_686,N_471);
xnor U6314 (N_6314,N_4790,N_3475);
nor U6315 (N_6315,N_4440,N_4353);
nand U6316 (N_6316,N_1216,N_3309);
xor U6317 (N_6317,N_828,N_4993);
or U6318 (N_6318,N_1763,N_2264);
nor U6319 (N_6319,N_1412,N_4398);
nand U6320 (N_6320,N_553,N_1747);
and U6321 (N_6321,N_300,N_3551);
and U6322 (N_6322,N_4539,N_1499);
nand U6323 (N_6323,N_63,N_306);
nand U6324 (N_6324,N_3384,N_2609);
and U6325 (N_6325,N_2231,N_1049);
or U6326 (N_6326,N_296,N_3846);
xnor U6327 (N_6327,N_824,N_24);
and U6328 (N_6328,N_1851,N_4164);
nor U6329 (N_6329,N_1556,N_3730);
or U6330 (N_6330,N_747,N_3052);
or U6331 (N_6331,N_2736,N_4027);
or U6332 (N_6332,N_3413,N_2753);
nand U6333 (N_6333,N_3616,N_3097);
and U6334 (N_6334,N_1516,N_4896);
and U6335 (N_6335,N_477,N_4681);
or U6336 (N_6336,N_2104,N_3274);
nor U6337 (N_6337,N_4211,N_2752);
nand U6338 (N_6338,N_3498,N_332);
nor U6339 (N_6339,N_197,N_4204);
nor U6340 (N_6340,N_619,N_4311);
nand U6341 (N_6341,N_3805,N_2999);
and U6342 (N_6342,N_4198,N_517);
nor U6343 (N_6343,N_4890,N_746);
and U6344 (N_6344,N_867,N_796);
and U6345 (N_6345,N_225,N_62);
xor U6346 (N_6346,N_969,N_1898);
nor U6347 (N_6347,N_465,N_4105);
nor U6348 (N_6348,N_2867,N_4400);
or U6349 (N_6349,N_1023,N_880);
nor U6350 (N_6350,N_185,N_626);
or U6351 (N_6351,N_2580,N_734);
or U6352 (N_6352,N_803,N_2735);
or U6353 (N_6353,N_3452,N_4220);
and U6354 (N_6354,N_1706,N_1924);
nor U6355 (N_6355,N_1257,N_1920);
xor U6356 (N_6356,N_4632,N_3617);
xnor U6357 (N_6357,N_1024,N_4946);
nor U6358 (N_6358,N_4051,N_4373);
or U6359 (N_6359,N_408,N_1348);
or U6360 (N_6360,N_4363,N_2756);
nor U6361 (N_6361,N_764,N_2751);
xnor U6362 (N_6362,N_3555,N_4793);
nor U6363 (N_6363,N_1065,N_1963);
and U6364 (N_6364,N_4333,N_1218);
or U6365 (N_6365,N_2583,N_4116);
and U6366 (N_6366,N_2340,N_2741);
nand U6367 (N_6367,N_722,N_2208);
and U6368 (N_6368,N_403,N_2737);
or U6369 (N_6369,N_3390,N_34);
xnor U6370 (N_6370,N_3840,N_198);
and U6371 (N_6371,N_941,N_939);
nand U6372 (N_6372,N_3930,N_1653);
nand U6373 (N_6373,N_830,N_3005);
and U6374 (N_6374,N_2663,N_1137);
or U6375 (N_6375,N_3238,N_67);
or U6376 (N_6376,N_3545,N_1215);
nor U6377 (N_6377,N_4089,N_4241);
or U6378 (N_6378,N_1449,N_2303);
nor U6379 (N_6379,N_1826,N_1159);
and U6380 (N_6380,N_4752,N_1091);
nand U6381 (N_6381,N_4855,N_1864);
and U6382 (N_6382,N_4124,N_1854);
nor U6383 (N_6383,N_3655,N_4091);
nor U6384 (N_6384,N_4159,N_3051);
nor U6385 (N_6385,N_2054,N_1751);
nand U6386 (N_6386,N_1952,N_2588);
nand U6387 (N_6387,N_1227,N_4555);
nand U6388 (N_6388,N_2567,N_361);
nor U6389 (N_6389,N_4065,N_3675);
nor U6390 (N_6390,N_3525,N_4615);
nand U6391 (N_6391,N_1148,N_2845);
and U6392 (N_6392,N_1392,N_3006);
xnor U6393 (N_6393,N_2749,N_449);
xor U6394 (N_6394,N_4425,N_3625);
nand U6395 (N_6395,N_210,N_3193);
or U6396 (N_6396,N_977,N_590);
or U6397 (N_6397,N_3266,N_1585);
nor U6398 (N_6398,N_4041,N_2691);
nand U6399 (N_6399,N_1840,N_1503);
nor U6400 (N_6400,N_3482,N_1103);
or U6401 (N_6401,N_4345,N_2814);
and U6402 (N_6402,N_4527,N_71);
nand U6403 (N_6403,N_4452,N_1600);
nand U6404 (N_6404,N_3153,N_1413);
nor U6405 (N_6405,N_3455,N_2889);
xnor U6406 (N_6406,N_3225,N_4618);
xnor U6407 (N_6407,N_2402,N_1107);
nand U6408 (N_6408,N_2156,N_825);
nand U6409 (N_6409,N_4443,N_2053);
and U6410 (N_6410,N_4206,N_4380);
or U6411 (N_6411,N_2799,N_2640);
nor U6412 (N_6412,N_4066,N_1454);
nand U6413 (N_6413,N_1378,N_4286);
or U6414 (N_6414,N_1364,N_2301);
xor U6415 (N_6415,N_615,N_893);
nor U6416 (N_6416,N_4293,N_2943);
xnor U6417 (N_6417,N_1473,N_943);
nand U6418 (N_6418,N_2613,N_3567);
and U6419 (N_6419,N_2917,N_1315);
xor U6420 (N_6420,N_3595,N_3750);
or U6421 (N_6421,N_2693,N_292);
or U6422 (N_6422,N_4092,N_3349);
and U6423 (N_6423,N_2110,N_1);
nand U6424 (N_6424,N_156,N_2623);
or U6425 (N_6425,N_4436,N_2571);
nand U6426 (N_6426,N_3815,N_70);
nand U6427 (N_6427,N_3060,N_3832);
nand U6428 (N_6428,N_4163,N_1081);
and U6429 (N_6429,N_3810,N_1040);
or U6430 (N_6430,N_2073,N_2367);
or U6431 (N_6431,N_2082,N_365);
nor U6432 (N_6432,N_914,N_2441);
nor U6433 (N_6433,N_2909,N_440);
or U6434 (N_6434,N_2185,N_3021);
xor U6435 (N_6435,N_2589,N_578);
nand U6436 (N_6436,N_3513,N_2222);
nor U6437 (N_6437,N_1333,N_3771);
xnor U6438 (N_6438,N_688,N_896);
and U6439 (N_6439,N_286,N_2426);
and U6440 (N_6440,N_853,N_1363);
nor U6441 (N_6441,N_3540,N_324);
or U6442 (N_6442,N_271,N_679);
and U6443 (N_6443,N_625,N_2817);
xor U6444 (N_6444,N_4942,N_1904);
nand U6445 (N_6445,N_2299,N_737);
nand U6446 (N_6446,N_3442,N_3727);
or U6447 (N_6447,N_3704,N_592);
and U6448 (N_6448,N_3660,N_3501);
nand U6449 (N_6449,N_419,N_4228);
or U6450 (N_6450,N_2631,N_178);
nand U6451 (N_6451,N_1624,N_2372);
nand U6452 (N_6452,N_9,N_962);
nand U6453 (N_6453,N_2548,N_2824);
nand U6454 (N_6454,N_571,N_4788);
or U6455 (N_6455,N_1343,N_878);
and U6456 (N_6456,N_282,N_4754);
or U6457 (N_6457,N_4427,N_2394);
or U6458 (N_6458,N_495,N_3800);
or U6459 (N_6459,N_547,N_2963);
xor U6460 (N_6460,N_1638,N_2466);
or U6461 (N_6461,N_2536,N_3161);
nor U6462 (N_6462,N_3016,N_3917);
and U6463 (N_6463,N_327,N_4653);
and U6464 (N_6464,N_666,N_2476);
or U6465 (N_6465,N_1875,N_263);
nand U6466 (N_6466,N_4382,N_2178);
or U6467 (N_6467,N_3580,N_1038);
nand U6468 (N_6468,N_1902,N_2707);
xor U6469 (N_6469,N_4412,N_2850);
and U6470 (N_6470,N_2056,N_3360);
or U6471 (N_6471,N_3123,N_2308);
and U6472 (N_6472,N_3958,N_4767);
xor U6473 (N_6473,N_607,N_1561);
nor U6474 (N_6474,N_4611,N_3312);
xnor U6475 (N_6475,N_4434,N_351);
and U6476 (N_6476,N_4281,N_353);
and U6477 (N_6477,N_1636,N_4334);
nand U6478 (N_6478,N_3697,N_322);
or U6479 (N_6479,N_2929,N_2883);
and U6480 (N_6480,N_2782,N_3782);
or U6481 (N_6481,N_1727,N_2184);
or U6482 (N_6482,N_4801,N_4347);
and U6483 (N_6483,N_3935,N_4395);
or U6484 (N_6484,N_276,N_274);
nand U6485 (N_6485,N_4385,N_3019);
nor U6486 (N_6486,N_2498,N_4060);
nor U6487 (N_6487,N_4080,N_1365);
or U6488 (N_6488,N_4749,N_2932);
nor U6489 (N_6489,N_2358,N_325);
nor U6490 (N_6490,N_2686,N_703);
or U6491 (N_6491,N_2039,N_2017);
or U6492 (N_6492,N_3856,N_1456);
and U6493 (N_6493,N_793,N_2962);
xor U6494 (N_6494,N_3282,N_4823);
and U6495 (N_6495,N_783,N_85);
nor U6496 (N_6496,N_68,N_724);
nand U6497 (N_6497,N_698,N_2076);
nand U6498 (N_6498,N_4923,N_4493);
nor U6499 (N_6499,N_2818,N_3147);
or U6500 (N_6500,N_1807,N_2797);
xor U6501 (N_6501,N_4174,N_4134);
nand U6502 (N_6502,N_4194,N_455);
nor U6503 (N_6503,N_2599,N_2733);
nor U6504 (N_6504,N_3887,N_3362);
xnor U6505 (N_6505,N_1171,N_2838);
xnor U6506 (N_6506,N_1168,N_2870);
nor U6507 (N_6507,N_1312,N_1646);
xnor U6508 (N_6508,N_217,N_1601);
nor U6509 (N_6509,N_2611,N_4647);
or U6510 (N_6510,N_3521,N_443);
nand U6511 (N_6511,N_2319,N_2930);
nand U6512 (N_6512,N_3728,N_1912);
and U6513 (N_6513,N_3692,N_769);
xnor U6514 (N_6514,N_2452,N_1326);
or U6515 (N_6515,N_206,N_2252);
or U6516 (N_6516,N_3331,N_4470);
xnor U6517 (N_6517,N_4190,N_1579);
nor U6518 (N_6518,N_748,N_2152);
nand U6519 (N_6519,N_2021,N_4902);
and U6520 (N_6520,N_1635,N_104);
and U6521 (N_6521,N_4366,N_4046);
nand U6522 (N_6522,N_928,N_3414);
nand U6523 (N_6523,N_3175,N_1719);
nand U6524 (N_6524,N_4720,N_3937);
nand U6525 (N_6525,N_3870,N_4453);
nor U6526 (N_6526,N_4882,N_1880);
nor U6527 (N_6527,N_3464,N_4217);
and U6528 (N_6528,N_1386,N_2907);
nor U6529 (N_6529,N_1973,N_3189);
xor U6530 (N_6530,N_1385,N_203);
or U6531 (N_6531,N_1566,N_3517);
and U6532 (N_6532,N_3102,N_4323);
or U6533 (N_6533,N_1338,N_2901);
and U6534 (N_6534,N_4866,N_1782);
nor U6535 (N_6535,N_526,N_461);
nor U6536 (N_6536,N_3737,N_1778);
xor U6537 (N_6537,N_4327,N_918);
nand U6538 (N_6538,N_2594,N_4560);
or U6539 (N_6539,N_1633,N_4265);
nand U6540 (N_6540,N_169,N_1663);
or U6541 (N_6541,N_3120,N_320);
nand U6542 (N_6542,N_3306,N_3835);
nor U6543 (N_6543,N_4,N_3824);
or U6544 (N_6544,N_1514,N_166);
or U6545 (N_6545,N_944,N_877);
or U6546 (N_6546,N_348,N_4049);
nand U6547 (N_6547,N_847,N_2230);
or U6548 (N_6548,N_179,N_756);
nand U6549 (N_6549,N_2254,N_1290);
or U6550 (N_6550,N_618,N_4667);
or U6551 (N_6551,N_559,N_309);
xnor U6552 (N_6552,N_3719,N_4920);
nand U6553 (N_6553,N_1831,N_1008);
and U6554 (N_6554,N_2371,N_3947);
and U6555 (N_6555,N_1397,N_442);
nor U6556 (N_6556,N_3911,N_191);
and U6557 (N_6557,N_1229,N_2557);
xor U6558 (N_6558,N_2425,N_1078);
nor U6559 (N_6559,N_2174,N_3726);
xnor U6560 (N_6560,N_4362,N_3430);
and U6561 (N_6561,N_3460,N_3818);
nand U6562 (N_6562,N_2439,N_294);
nand U6563 (N_6563,N_2401,N_3432);
nand U6564 (N_6564,N_3378,N_1533);
nand U6565 (N_6565,N_3031,N_4349);
or U6566 (N_6566,N_4446,N_3619);
and U6567 (N_6567,N_4234,N_4074);
nand U6568 (N_6568,N_1918,N_1095);
and U6569 (N_6569,N_1678,N_2293);
or U6570 (N_6570,N_367,N_4166);
nor U6571 (N_6571,N_3314,N_766);
nor U6572 (N_6572,N_642,N_1769);
and U6573 (N_6573,N_4316,N_3579);
or U6574 (N_6574,N_3711,N_582);
nor U6575 (N_6575,N_613,N_2504);
and U6576 (N_6576,N_2258,N_2676);
or U6577 (N_6577,N_245,N_202);
xnor U6578 (N_6578,N_3562,N_924);
nand U6579 (N_6579,N_3154,N_2097);
and U6580 (N_6580,N_4180,N_886);
nand U6581 (N_6581,N_2163,N_4271);
and U6582 (N_6582,N_1735,N_3155);
and U6583 (N_6583,N_1260,N_1193);
nor U6584 (N_6584,N_3220,N_2655);
or U6585 (N_6585,N_4444,N_787);
nand U6586 (N_6586,N_2124,N_3069);
nor U6587 (N_6587,N_2006,N_4263);
xnor U6588 (N_6588,N_790,N_4313);
nand U6589 (N_6589,N_4214,N_1722);
xor U6590 (N_6590,N_1970,N_290);
and U6591 (N_6591,N_3558,N_902);
nor U6592 (N_6592,N_4892,N_3007);
nand U6593 (N_6593,N_3041,N_2778);
nand U6594 (N_6594,N_2643,N_4437);
and U6595 (N_6595,N_871,N_3092);
or U6596 (N_6596,N_1540,N_740);
xnor U6597 (N_6597,N_4244,N_1764);
and U6598 (N_6598,N_909,N_4591);
xor U6599 (N_6599,N_4104,N_4184);
xor U6600 (N_6600,N_4223,N_456);
nand U6601 (N_6601,N_1135,N_967);
nand U6602 (N_6602,N_1327,N_870);
xnor U6603 (N_6603,N_2282,N_1209);
or U6604 (N_6604,N_767,N_757);
xnor U6605 (N_6605,N_3834,N_2976);
nor U6606 (N_6606,N_3176,N_1428);
nand U6607 (N_6607,N_2153,N_2702);
or U6608 (N_6608,N_1967,N_3556);
xor U6609 (N_6609,N_125,N_4635);
or U6610 (N_6610,N_3036,N_2854);
or U6611 (N_6611,N_1272,N_2952);
nor U6612 (N_6612,N_3689,N_2903);
nor U6613 (N_6613,N_4979,N_175);
or U6614 (N_6614,N_2210,N_4147);
or U6615 (N_6615,N_2970,N_80);
xor U6616 (N_6616,N_1839,N_2045);
nor U6617 (N_6617,N_4523,N_3696);
and U6618 (N_6618,N_2806,N_1640);
nand U6619 (N_6619,N_1396,N_1910);
xnor U6620 (N_6620,N_4982,N_4508);
and U6621 (N_6621,N_4976,N_3613);
xnor U6622 (N_6622,N_4568,N_1530);
and U6623 (N_6623,N_3851,N_2345);
nand U6624 (N_6624,N_3895,N_1198);
nor U6625 (N_6625,N_3473,N_76);
and U6626 (N_6626,N_1825,N_1817);
nor U6627 (N_6627,N_2800,N_2837);
and U6628 (N_6628,N_1565,N_3108);
or U6629 (N_6629,N_1346,N_2542);
or U6630 (N_6630,N_162,N_2634);
nand U6631 (N_6631,N_2780,N_1779);
nor U6632 (N_6632,N_1188,N_1789);
nor U6633 (N_6633,N_1760,N_2718);
xnor U6634 (N_6634,N_3484,N_1025);
or U6635 (N_6635,N_2714,N_1682);
nand U6636 (N_6636,N_3632,N_2653);
nand U6637 (N_6637,N_956,N_4329);
or U6638 (N_6638,N_4586,N_1329);
or U6639 (N_6639,N_2456,N_2511);
and U6640 (N_6640,N_4650,N_885);
xnor U6641 (N_6641,N_3533,N_3875);
or U6642 (N_6642,N_1211,N_1639);
and U6643 (N_6643,N_1761,N_4592);
nand U6644 (N_6644,N_1299,N_2969);
and U6645 (N_6645,N_3317,N_4644);
nor U6646 (N_6646,N_1832,N_2721);
and U6647 (N_6647,N_2363,N_4798);
nor U6648 (N_6648,N_4859,N_1379);
nand U6649 (N_6649,N_816,N_3529);
or U6650 (N_6650,N_4365,N_4028);
or U6651 (N_6651,N_2378,N_781);
and U6652 (N_6652,N_4732,N_4019);
nor U6653 (N_6653,N_2483,N_238);
nor U6654 (N_6654,N_1489,N_1295);
and U6655 (N_6655,N_43,N_1745);
and U6656 (N_6656,N_305,N_3925);
nor U6657 (N_6657,N_1313,N_4847);
nor U6658 (N_6658,N_229,N_4389);
or U6659 (N_6659,N_2171,N_2959);
and U6660 (N_6660,N_3319,N_4791);
and U6661 (N_6661,N_4101,N_3706);
nor U6662 (N_6662,N_3417,N_874);
nand U6663 (N_6663,N_1665,N_1213);
nor U6664 (N_6664,N_270,N_3233);
nand U6665 (N_6665,N_1651,N_2213);
xor U6666 (N_6666,N_3610,N_3827);
xnor U6667 (N_6667,N_859,N_1692);
nor U6668 (N_6668,N_3001,N_2351);
nand U6669 (N_6669,N_3570,N_3934);
and U6670 (N_6670,N_2405,N_241);
and U6671 (N_6671,N_4572,N_1945);
or U6672 (N_6672,N_1277,N_4212);
xor U6673 (N_6673,N_770,N_4735);
and U6674 (N_6674,N_4167,N_716);
or U6675 (N_6675,N_1527,N_2523);
nor U6676 (N_6676,N_844,N_3250);
or U6677 (N_6677,N_366,N_3054);
nand U6678 (N_6678,N_660,N_2012);
nor U6679 (N_6679,N_4628,N_3292);
or U6680 (N_6680,N_974,N_1377);
and U6681 (N_6681,N_297,N_1440);
and U6682 (N_6682,N_429,N_1590);
xnor U6683 (N_6683,N_1261,N_243);
or U6684 (N_6684,N_1847,N_3544);
and U6685 (N_6685,N_3515,N_4245);
or U6686 (N_6686,N_2462,N_95);
nor U6687 (N_6687,N_4836,N_555);
nor U6688 (N_6688,N_4242,N_503);
nor U6689 (N_6689,N_3848,N_105);
nand U6690 (N_6690,N_2884,N_4672);
and U6691 (N_6691,N_3969,N_3752);
nand U6692 (N_6692,N_1810,N_4579);
or U6693 (N_6693,N_1418,N_2694);
nand U6694 (N_6694,N_1158,N_1134);
or U6695 (N_6695,N_1857,N_1815);
and U6696 (N_6696,N_2386,N_3679);
nand U6697 (N_6697,N_4631,N_4974);
and U6698 (N_6698,N_2095,N_1552);
or U6699 (N_6699,N_1255,N_1534);
or U6700 (N_6700,N_3708,N_2660);
xnor U6701 (N_6701,N_4488,N_4967);
or U6702 (N_6702,N_3626,N_3653);
nand U6703 (N_6703,N_1959,N_3601);
nand U6704 (N_6704,N_1938,N_2214);
nand U6705 (N_6705,N_3029,N_3328);
nand U6706 (N_6706,N_3496,N_4929);
nor U6707 (N_6707,N_1991,N_2748);
nand U6708 (N_6708,N_4565,N_725);
nor U6709 (N_6709,N_3248,N_1256);
nand U6710 (N_6710,N_3744,N_2835);
nand U6711 (N_6711,N_1403,N_1233);
nand U6712 (N_6712,N_4562,N_2993);
or U6713 (N_6713,N_2937,N_3923);
nor U6714 (N_6714,N_2000,N_4848);
and U6715 (N_6715,N_3358,N_1956);
or U6716 (N_6716,N_3279,N_3952);
xor U6717 (N_6717,N_3392,N_4429);
nand U6718 (N_6718,N_3099,N_3449);
and U6719 (N_6719,N_1903,N_2094);
nand U6720 (N_6720,N_1861,N_186);
or U6721 (N_6721,N_4868,N_2092);
and U6722 (N_6722,N_4825,N_4025);
nand U6723 (N_6723,N_1704,N_1149);
nand U6724 (N_6724,N_2967,N_3428);
nand U6725 (N_6725,N_1479,N_1711);
and U6726 (N_6726,N_114,N_3169);
nand U6727 (N_6727,N_2685,N_262);
and U6728 (N_6728,N_546,N_4014);
and U6729 (N_6729,N_2101,N_3965);
or U6730 (N_6730,N_4085,N_3351);
nand U6731 (N_6731,N_3386,N_4945);
and U6732 (N_6732,N_48,N_641);
or U6733 (N_6733,N_654,N_4898);
or U6734 (N_6734,N_3049,N_2958);
or U6735 (N_6735,N_1710,N_2899);
and U6736 (N_6736,N_4914,N_4975);
and U6737 (N_6737,N_1932,N_4278);
and U6738 (N_6738,N_3263,N_1923);
and U6739 (N_6739,N_4930,N_473);
or U6740 (N_6740,N_2338,N_1589);
nand U6741 (N_6741,N_3938,N_691);
and U6742 (N_6742,N_2807,N_984);
or U6743 (N_6743,N_3389,N_4001);
or U6744 (N_6744,N_1838,N_2746);
nand U6745 (N_6745,N_4604,N_1866);
nand U6746 (N_6746,N_2067,N_2450);
and U6747 (N_6747,N_3067,N_1491);
nand U6748 (N_6748,N_2298,N_4462);
nor U6749 (N_6749,N_2731,N_4267);
or U6750 (N_6750,N_3659,N_1699);
nand U6751 (N_6751,N_2603,N_4973);
nand U6752 (N_6752,N_3476,N_2983);
xnor U6753 (N_6753,N_2081,N_1026);
and U6754 (N_6754,N_2713,N_4909);
and U6755 (N_6755,N_1697,N_165);
nand U6756 (N_6756,N_949,N_1150);
or U6757 (N_6757,N_550,N_690);
and U6758 (N_6758,N_3128,N_539);
nand U6759 (N_6759,N_3245,N_2376);
nand U6760 (N_6760,N_988,N_2221);
nor U6761 (N_6761,N_4512,N_4816);
xor U6762 (N_6762,N_4042,N_577);
nor U6763 (N_6763,N_2872,N_504);
and U6764 (N_6764,N_3162,N_3605);
or U6765 (N_6765,N_817,N_1937);
nor U6766 (N_6766,N_3130,N_2271);
and U6767 (N_6767,N_4842,N_3320);
nand U6768 (N_6768,N_2323,N_3968);
nor U6769 (N_6769,N_4052,N_4108);
or U6770 (N_6770,N_3295,N_420);
or U6771 (N_6771,N_3583,N_13);
and U6772 (N_6772,N_102,N_1577);
nand U6773 (N_6773,N_2785,N_3926);
and U6774 (N_6774,N_2,N_3232);
and U6775 (N_6775,N_3868,N_1271);
or U6776 (N_6776,N_2145,N_3340);
nor U6777 (N_6777,N_3702,N_4118);
xnor U6778 (N_6778,N_153,N_199);
nor U6779 (N_6779,N_3122,N_207);
nor U6780 (N_6780,N_4129,N_4496);
or U6781 (N_6781,N_3901,N_833);
or U6782 (N_6782,N_4759,N_2755);
nor U6783 (N_6783,N_1052,N_1020);
xnor U6784 (N_6784,N_1286,N_4875);
xnor U6785 (N_6785,N_4417,N_3080);
nand U6786 (N_6786,N_1099,N_2253);
or U6787 (N_6787,N_2335,N_4465);
or U6788 (N_6788,N_1369,N_1357);
nor U6789 (N_6789,N_1522,N_2015);
nand U6790 (N_6790,N_2042,N_2096);
or U6791 (N_6791,N_3291,N_4356);
or U6792 (N_6792,N_2277,N_925);
or U6793 (N_6793,N_214,N_1837);
nand U6794 (N_6794,N_1136,N_317);
and U6795 (N_6795,N_4917,N_4680);
nand U6796 (N_6796,N_4258,N_2133);
or U6797 (N_6797,N_2843,N_47);
nand U6798 (N_6798,N_4737,N_173);
nand U6799 (N_6799,N_2169,N_3293);
nand U6800 (N_6800,N_706,N_284);
nor U6801 (N_6801,N_1863,N_2119);
and U6802 (N_6802,N_2562,N_2224);
and U6803 (N_6803,N_2463,N_2651);
or U6804 (N_6804,N_2879,N_606);
nand U6805 (N_6805,N_1006,N_1311);
or U6806 (N_6806,N_4237,N_1511);
or U6807 (N_6807,N_1477,N_2385);
or U6808 (N_6808,N_3398,N_4953);
nand U6809 (N_6809,N_1830,N_707);
or U6810 (N_6810,N_1729,N_3201);
or U6811 (N_6811,N_4155,N_3141);
nor U6812 (N_6812,N_3222,N_1062);
or U6813 (N_6813,N_4413,N_413);
and U6814 (N_6814,N_1087,N_4250);
or U6815 (N_6815,N_1310,N_1841);
nor U6816 (N_6816,N_772,N_4391);
nand U6817 (N_6817,N_903,N_2113);
nand U6818 (N_6818,N_4671,N_4955);
nor U6819 (N_6819,N_4912,N_3435);
nor U6820 (N_6820,N_1462,N_4528);
or U6821 (N_6821,N_4716,N_3043);
and U6822 (N_6822,N_2495,N_2334);
nand U6823 (N_6823,N_79,N_1694);
or U6824 (N_6824,N_819,N_3443);
and U6825 (N_6825,N_2107,N_1708);
nor U6826 (N_6826,N_3820,N_2996);
and U6827 (N_6827,N_3002,N_2151);
or U6828 (N_6828,N_638,N_4858);
or U6829 (N_6829,N_1083,N_3761);
nor U6830 (N_6830,N_3009,N_1987);
nand U6831 (N_6831,N_2220,N_1580);
nor U6832 (N_6832,N_1526,N_3399);
xor U6833 (N_6833,N_4598,N_2738);
or U6834 (N_6834,N_2148,N_3985);
and U6835 (N_6835,N_4925,N_469);
nand U6836 (N_6836,N_4952,N_3565);
nor U6837 (N_6837,N_3444,N_4837);
nor U6838 (N_6838,N_3025,N_2645);
nand U6839 (N_6839,N_588,N_4978);
or U6840 (N_6840,N_1513,N_1195);
nor U6841 (N_6841,N_4509,N_3920);
and U6842 (N_6842,N_3813,N_665);
nand U6843 (N_6843,N_1990,N_622);
or U6844 (N_6844,N_4802,N_1969);
nor U6845 (N_6845,N_1858,N_3865);
and U6846 (N_6846,N_554,N_1965);
nand U6847 (N_6847,N_1883,N_3786);
or U6848 (N_6848,N_4257,N_231);
nor U6849 (N_6849,N_1876,N_2237);
or U6850 (N_6850,N_4396,N_848);
and U6851 (N_6851,N_1074,N_4997);
nand U6852 (N_6852,N_4853,N_1684);
nand U6853 (N_6853,N_4119,N_385);
nor U6854 (N_6854,N_3880,N_2859);
nand U6855 (N_6855,N_2212,N_3014);
nor U6856 (N_6856,N_478,N_4273);
or U6857 (N_6857,N_3961,N_4285);
nand U6858 (N_6858,N_4260,N_4580);
or U6859 (N_6859,N_3918,N_4071);
and U6860 (N_6860,N_2717,N_4869);
or U6861 (N_6861,N_4656,N_346);
or U6862 (N_6862,N_1974,N_1073);
and U6863 (N_6863,N_652,N_2320);
xor U6864 (N_6864,N_3365,N_1376);
xnor U6865 (N_6865,N_3070,N_3829);
nand U6866 (N_6866,N_1867,N_2068);
nor U6867 (N_6867,N_2506,N_2364);
and U6868 (N_6868,N_4111,N_993);
or U6869 (N_6869,N_3745,N_2139);
or U6870 (N_6870,N_4421,N_714);
nand U6871 (N_6871,N_1100,N_674);
or U6872 (N_6872,N_4908,N_697);
and U6873 (N_6873,N_4595,N_2484);
xnor U6874 (N_6874,N_4800,N_337);
and U6875 (N_6875,N_4699,N_549);
nor U6876 (N_6876,N_1549,N_3668);
and U6877 (N_6877,N_506,N_1432);
nand U6878 (N_6878,N_4888,N_2135);
and U6879 (N_6879,N_2955,N_1949);
or U6880 (N_6880,N_2563,N_4636);
nor U6881 (N_6881,N_3735,N_1816);
nor U6882 (N_6882,N_1895,N_2762);
and U6883 (N_6883,N_3954,N_4350);
nand U6884 (N_6884,N_3987,N_256);
nand U6885 (N_6885,N_2839,N_1571);
xnor U6886 (N_6886,N_2945,N_2921);
and U6887 (N_6887,N_1486,N_3763);
or U6888 (N_6888,N_1946,N_4491);
and U6889 (N_6889,N_1915,N_2725);
and U6890 (N_6890,N_386,N_3305);
or U6891 (N_6891,N_1373,N_650);
nand U6892 (N_6892,N_4745,N_343);
and U6893 (N_6893,N_4168,N_789);
nor U6894 (N_6894,N_1140,N_4690);
xnor U6895 (N_6895,N_872,N_792);
or U6896 (N_6896,N_3654,N_3713);
xor U6897 (N_6897,N_3207,N_3094);
nand U6898 (N_6898,N_3572,N_2539);
or U6899 (N_6899,N_218,N_64);
or U6900 (N_6900,N_780,N_4248);
and U6901 (N_6901,N_540,N_3100);
and U6902 (N_6902,N_3860,N_2834);
xnor U6903 (N_6903,N_4874,N_1115);
or U6904 (N_6904,N_2953,N_3568);
nor U6905 (N_6905,N_196,N_1821);
and U6906 (N_6906,N_4747,N_1986);
nand U6907 (N_6907,N_1803,N_658);
xor U6908 (N_6908,N_2936,N_629);
nand U6909 (N_6909,N_1263,N_1780);
or U6910 (N_6910,N_2608,N_2857);
nand U6911 (N_6911,N_2546,N_107);
nand U6912 (N_6912,N_3984,N_2786);
nor U6913 (N_6913,N_4469,N_2057);
xor U6914 (N_6914,N_149,N_664);
xor U6915 (N_6915,N_3751,N_1693);
and U6916 (N_6916,N_1039,N_4886);
nand U6917 (N_6917,N_3522,N_1042);
nor U6918 (N_6918,N_4253,N_1812);
and U6919 (N_6919,N_139,N_2211);
nor U6920 (N_6920,N_1335,N_4717);
and U6921 (N_6921,N_1239,N_3010);
and U6922 (N_6922,N_4494,N_3056);
and U6923 (N_6923,N_396,N_3144);
and U6924 (N_6924,N_3760,N_4428);
xnor U6925 (N_6925,N_4034,N_731);
and U6926 (N_6926,N_2004,N_1425);
and U6927 (N_6927,N_1043,N_3707);
xor U6928 (N_6928,N_581,N_1929);
xnor U6929 (N_6929,N_1614,N_3867);
nand U6930 (N_6930,N_3606,N_519);
and U6931 (N_6931,N_3894,N_4026);
or U6932 (N_6932,N_2020,N_3403);
and U6933 (N_6933,N_3039,N_3090);
or U6934 (N_6934,N_2924,N_4695);
and U6935 (N_6935,N_2259,N_482);
and U6936 (N_6936,N_1855,N_4393);
or U6937 (N_6937,N_2442,N_2433);
or U6938 (N_6938,N_2789,N_1797);
and U6939 (N_6939,N_633,N_81);
nor U6940 (N_6940,N_3085,N_1220);
or U6941 (N_6941,N_336,N_3192);
and U6942 (N_6942,N_2632,N_806);
xnor U6943 (N_6943,N_2754,N_2569);
nand U6944 (N_6944,N_2238,N_3936);
xor U6945 (N_6945,N_1888,N_3205);
nand U6946 (N_6946,N_1829,N_1783);
nor U6947 (N_6947,N_1347,N_4728);
or U6948 (N_6948,N_2325,N_2914);
nand U6949 (N_6949,N_1868,N_1506);
nor U6950 (N_6950,N_2768,N_1705);
or U6951 (N_6951,N_484,N_1754);
or U6952 (N_6952,N_4037,N_453);
nor U6953 (N_6953,N_2129,N_151);
and U6954 (N_6954,N_2761,N_4682);
xor U6955 (N_6955,N_255,N_3053);
or U6956 (N_6956,N_1240,N_1123);
nand U6957 (N_6957,N_4649,N_3050);
nor U6958 (N_6958,N_1737,N_569);
or U6959 (N_6959,N_1742,N_2874);
nor U6960 (N_6960,N_1824,N_4513);
and U6961 (N_6961,N_3359,N_2628);
or U6962 (N_6962,N_261,N_3725);
xor U6963 (N_6963,N_2100,N_3265);
xnor U6964 (N_6964,N_1642,N_2370);
and U6965 (N_6965,N_3900,N_2479);
and U6966 (N_6966,N_4947,N_4059);
nand U6967 (N_6967,N_2412,N_3821);
nor U6968 (N_6968,N_4535,N_4643);
nand U6969 (N_6969,N_4310,N_3571);
nor U6970 (N_6970,N_3817,N_1430);
or U6971 (N_6971,N_2809,N_4047);
xnor U6972 (N_6972,N_3729,N_1167);
and U6973 (N_6973,N_3877,N_1786);
nor U6974 (N_6974,N_1337,N_3684);
or U6975 (N_6975,N_315,N_2126);
or U6976 (N_6976,N_574,N_2763);
and U6977 (N_6977,N_810,N_3788);
nor U6978 (N_6978,N_2275,N_4110);
nand U6979 (N_6979,N_755,N_3372);
nand U6980 (N_6980,N_3523,N_1452);
nand U6981 (N_6981,N_3243,N_604);
nor U6982 (N_6982,N_2451,N_1629);
nand U6983 (N_6983,N_832,N_4424);
and U6984 (N_6984,N_3931,N_4889);
or U6985 (N_6985,N_1748,N_4922);
or U6986 (N_6986,N_41,N_3896);
and U6987 (N_6987,N_976,N_1591);
and U6988 (N_6988,N_3701,N_3749);
and U6989 (N_6989,N_3767,N_2106);
or U6990 (N_6990,N_356,N_1451);
nor U6991 (N_6991,N_28,N_3681);
or U6992 (N_6992,N_4468,N_4581);
and U6993 (N_6993,N_371,N_749);
nand U6994 (N_6994,N_3329,N_2975);
and U6995 (N_6995,N_3758,N_1900);
and U6996 (N_6996,N_283,N_4715);
and U6997 (N_6997,N_3370,N_2805);
nand U6998 (N_6998,N_3486,N_4162);
nand U6999 (N_6999,N_3433,N_2091);
xnor U7000 (N_7000,N_2167,N_2399);
nand U7001 (N_7001,N_1448,N_2602);
xor U7002 (N_7002,N_4481,N_2988);
xor U7003 (N_7003,N_1408,N_4986);
or U7004 (N_7004,N_2595,N_170);
nand U7005 (N_7005,N_4304,N_4734);
nand U7006 (N_7006,N_4812,N_84);
xnor U7007 (N_7007,N_1652,N_3380);
nand U7008 (N_7008,N_4919,N_1695);
and U7009 (N_7009,N_992,N_2257);
and U7010 (N_7010,N_2182,N_1518);
nor U7011 (N_7011,N_1426,N_2961);
or U7012 (N_7012,N_1627,N_3422);
xor U7013 (N_7013,N_2336,N_1598);
and U7014 (N_7014,N_4100,N_233);
nor U7015 (N_7015,N_1415,N_2558);
and U7016 (N_7016,N_190,N_712);
nand U7017 (N_7017,N_1037,N_3330);
or U7018 (N_7018,N_2470,N_3071);
or U7019 (N_7019,N_4751,N_2946);
and U7020 (N_7020,N_4884,N_2035);
or U7021 (N_7021,N_1993,N_4409);
xnor U7022 (N_7022,N_1320,N_1714);
nor U7023 (N_7023,N_4192,N_3125);
or U7024 (N_7024,N_2650,N_4663);
or U7025 (N_7025,N_3776,N_3269);
nand U7026 (N_7026,N_4030,N_2192);
nand U7027 (N_7027,N_881,N_1677);
and U7028 (N_7028,N_3589,N_3457);
and U7029 (N_7029,N_3420,N_4057);
or U7030 (N_7030,N_3264,N_1072);
nand U7031 (N_7031,N_736,N_3893);
or U7032 (N_7032,N_3164,N_2949);
nor U7033 (N_7033,N_4141,N_1528);
nand U7034 (N_7034,N_1569,N_3607);
xor U7035 (N_7035,N_4863,N_906);
nand U7036 (N_7036,N_4299,N_2847);
nand U7037 (N_7037,N_2695,N_2229);
nand U7038 (N_7038,N_485,N_562);
or U7039 (N_7039,N_0,N_2669);
and U7040 (N_7040,N_3892,N_1102);
and U7041 (N_7041,N_3171,N_2538);
and U7042 (N_7042,N_1563,N_1625);
and U7043 (N_7043,N_1151,N_1190);
and U7044 (N_7044,N_101,N_4961);
xnor U7045 (N_7045,N_3967,N_2361);
nor U7046 (N_7046,N_2033,N_2066);
or U7047 (N_7047,N_4205,N_3101);
and U7048 (N_7048,N_4430,N_2815);
and U7049 (N_7049,N_1843,N_2384);
nand U7050 (N_7050,N_1070,N_492);
and U7051 (N_7051,N_1034,N_1707);
xnor U7052 (N_7052,N_3796,N_3743);
nand U7053 (N_7053,N_3003,N_3530);
or U7054 (N_7054,N_3345,N_132);
and U7055 (N_7055,N_4746,N_799);
nand U7056 (N_7056,N_3253,N_3466);
nand U7057 (N_7057,N_3348,N_4852);
or U7058 (N_7058,N_978,N_2480);
or U7059 (N_7059,N_2173,N_3643);
nor U7060 (N_7060,N_2864,N_3234);
nor U7061 (N_7061,N_1723,N_4634);
and U7062 (N_7062,N_3514,N_1334);
nor U7063 (N_7063,N_2494,N_4123);
and U7064 (N_7064,N_464,N_120);
and U7065 (N_7065,N_2421,N_4566);
nor U7066 (N_7066,N_10,N_2379);
nor U7067 (N_7067,N_2307,N_2300);
or U7068 (N_7068,N_3990,N_146);
or U7069 (N_7069,N_3897,N_1267);
nor U7070 (N_7070,N_2144,N_4913);
nand U7071 (N_7071,N_3139,N_2256);
and U7072 (N_7072,N_4614,N_3299);
and U7073 (N_7073,N_128,N_1252);
or U7074 (N_7074,N_16,N_2747);
nand U7075 (N_7075,N_3718,N_4215);
or U7076 (N_7076,N_1537,N_4660);
nor U7077 (N_7077,N_1743,N_1567);
or U7078 (N_7078,N_3784,N_3086);
nand U7079 (N_7079,N_1124,N_362);
nor U7080 (N_7080,N_2855,N_3246);
or U7081 (N_7081,N_4361,N_3690);
nor U7082 (N_7082,N_4355,N_3456);
or U7083 (N_7083,N_4828,N_232);
nor U7084 (N_7084,N_116,N_1758);
or U7085 (N_7085,N_1382,N_183);
nor U7086 (N_7086,N_2090,N_2641);
nand U7087 (N_7087,N_3237,N_3539);
nand U7088 (N_7088,N_1291,N_1287);
nor U7089 (N_7089,N_3777,N_2331);
nand U7090 (N_7090,N_423,N_2541);
nand U7091 (N_7091,N_761,N_2478);
nor U7092 (N_7092,N_2759,N_4048);
or U7093 (N_7093,N_1265,N_4459);
or U7094 (N_7094,N_4012,N_1031);
and U7095 (N_7095,N_2181,N_234);
nor U7096 (N_7096,N_180,N_1529);
nand U7097 (N_7097,N_599,N_4670);
or U7098 (N_7098,N_1047,N_2514);
or U7099 (N_7099,N_1955,N_4844);
and U7100 (N_7100,N_3377,N_2468);
and U7101 (N_7101,N_4658,N_3165);
nand U7102 (N_7102,N_3326,N_1675);
or U7103 (N_7103,N_1977,N_2724);
or U7104 (N_7104,N_2279,N_778);
nand U7105 (N_7105,N_4438,N_3594);
and U7106 (N_7106,N_2241,N_3166);
or U7107 (N_7107,N_2821,N_452);
and U7108 (N_7108,N_1507,N_3065);
and U7109 (N_7109,N_4102,N_411);
nand U7110 (N_7110,N_2647,N_4841);
and U7111 (N_7111,N_3823,N_1388);
nor U7112 (N_7112,N_4700,N_2274);
or U7113 (N_7113,N_3560,N_3431);
or U7114 (N_7114,N_680,N_4336);
nand U7115 (N_7115,N_2781,N_2235);
nand U7116 (N_7116,N_3957,N_2827);
or U7117 (N_7117,N_1953,N_3117);
or U7118 (N_7118,N_97,N_3103);
nor U7119 (N_7119,N_3167,N_135);
or U7120 (N_7120,N_3180,N_4687);
xor U7121 (N_7121,N_4878,N_3383);
nor U7122 (N_7122,N_2227,N_1531);
and U7123 (N_7123,N_457,N_460);
and U7124 (N_7124,N_1519,N_3497);
and U7125 (N_7125,N_3878,N_1389);
or U7126 (N_7126,N_3638,N_1104);
nor U7127 (N_7127,N_2920,N_370);
and U7128 (N_7128,N_3290,N_3188);
or U7129 (N_7129,N_248,N_2812);
nand U7130 (N_7130,N_3596,N_2418);
nor U7131 (N_7131,N_31,N_2305);
and U7132 (N_7132,N_2880,N_3537);
or U7133 (N_7133,N_319,N_438);
and U7134 (N_7134,N_879,N_1084);
nand U7135 (N_7135,N_4095,N_4264);
or U7136 (N_7136,N_2722,N_1372);
and U7137 (N_7137,N_529,N_4157);
xor U7138 (N_7138,N_659,N_587);
nand U7139 (N_7139,N_3015,N_3785);
nand U7140 (N_7140,N_4729,N_2059);
nor U7141 (N_7141,N_1458,N_672);
nor U7142 (N_7142,N_4015,N_338);
or U7143 (N_7143,N_3717,N_4601);
xnor U7144 (N_7144,N_2049,N_2912);
or U7145 (N_7145,N_742,N_4609);
nand U7146 (N_7146,N_2519,N_2516);
and U7147 (N_7147,N_2919,N_2978);
nand U7148 (N_7148,N_2018,N_3057);
nand U7149 (N_7149,N_3145,N_3566);
nand U7150 (N_7150,N_2454,N_4621);
nor U7151 (N_7151,N_1361,N_2811);
nand U7152 (N_7152,N_1463,N_4187);
xor U7153 (N_7153,N_3609,N_3814);
and U7154 (N_7154,N_2497,N_1940);
xnor U7155 (N_7155,N_1765,N_326);
nand U7156 (N_7156,N_2183,N_856);
nand U7157 (N_7157,N_2198,N_1962);
nor U7158 (N_7158,N_4010,N_1539);
xor U7159 (N_7159,N_133,N_851);
or U7160 (N_7160,N_4969,N_3182);
xor U7161 (N_7161,N_4654,N_1142);
and U7162 (N_7162,N_250,N_2705);
nand U7163 (N_7163,N_4689,N_1163);
nand U7164 (N_7164,N_3447,N_1485);
or U7165 (N_7165,N_1017,N_2417);
nor U7166 (N_7166,N_2037,N_4933);
nand U7167 (N_7167,N_4626,N_4498);
nor U7168 (N_7168,N_354,N_1818);
nand U7169 (N_7169,N_1882,N_2527);
and U7170 (N_7170,N_2935,N_4077);
or U7171 (N_7171,N_3109,N_3252);
and U7172 (N_7172,N_4701,N_4449);
and U7173 (N_7173,N_1644,N_3648);
nand U7174 (N_7174,N_1574,N_2026);
and U7175 (N_7175,N_2062,N_1223);
xnor U7176 (N_7176,N_913,N_946);
xnor U7177 (N_7177,N_3030,N_1278);
and U7178 (N_7178,N_4439,N_1270);
nand U7179 (N_7179,N_4364,N_4694);
nand U7180 (N_7180,N_2315,N_1899);
nand U7181 (N_7181,N_875,N_1060);
and U7182 (N_7182,N_3549,N_1679);
and U7183 (N_7183,N_3426,N_2915);
or U7184 (N_7184,N_4785,N_3576);
or U7185 (N_7185,N_3133,N_4939);
or U7186 (N_7186,N_3026,N_205);
and U7187 (N_7187,N_2195,N_106);
and U7188 (N_7188,N_1184,N_195);
nand U7189 (N_7189,N_3260,N_4928);
or U7190 (N_7190,N_2947,N_4083);
nor U7191 (N_7191,N_1208,N_1309);
and U7192 (N_7192,N_4915,N_4911);
nand U7193 (N_7193,N_1709,N_3357);
nand U7194 (N_7194,N_3106,N_1322);
nor U7195 (N_7195,N_1927,N_1869);
nand U7196 (N_7196,N_538,N_3904);
or U7197 (N_7197,N_843,N_2923);
nand U7198 (N_7198,N_3552,N_4322);
or U7199 (N_7199,N_4069,N_2410);
xor U7200 (N_7200,N_3806,N_4266);
or U7201 (N_7201,N_2013,N_630);
nand U7202 (N_7202,N_3747,N_1775);
nor U7203 (N_7203,N_2579,N_4600);
and U7204 (N_7204,N_3170,N_1459);
nand U7205 (N_7205,N_3780,N_3586);
xor U7206 (N_7206,N_4541,N_3110);
and U7207 (N_7207,N_472,N_4312);
or U7208 (N_7208,N_572,N_1545);
nand U7209 (N_7209,N_718,N_4371);
nor U7210 (N_7210,N_226,N_3478);
nand U7211 (N_7211,N_436,N_561);
and U7212 (N_7212,N_259,N_4617);
xor U7213 (N_7213,N_4819,N_986);
or U7214 (N_7214,N_1061,N_2649);
nor U7215 (N_7215,N_1718,N_4218);
or U7216 (N_7216,N_744,N_1626);
nor U7217 (N_7217,N_3212,N_4537);
or U7218 (N_7218,N_2877,N_4725);
or U7219 (N_7219,N_267,N_4419);
xnor U7220 (N_7220,N_3375,N_585);
nor U7221 (N_7221,N_575,N_1852);
xnor U7222 (N_7222,N_4445,N_3344);
or U7223 (N_7223,N_2732,N_4031);
or U7224 (N_7224,N_4900,N_4661);
and U7225 (N_7225,N_2657,N_3982);
nor U7226 (N_7226,N_4008,N_3157);
nor U7227 (N_7227,N_4354,N_4518);
xor U7228 (N_7228,N_1980,N_890);
and U7229 (N_7229,N_4087,N_3932);
nand U7230 (N_7230,N_4542,N_2036);
nor U7231 (N_7231,N_4114,N_1724);
nand U7232 (N_7232,N_2898,N_4339);
and U7233 (N_7233,N_2767,N_801);
and U7234 (N_7234,N_1957,N_3000);
or U7235 (N_7235,N_409,N_2633);
xnor U7236 (N_7236,N_3803,N_3873);
and U7237 (N_7237,N_2743,N_4279);
nand U7238 (N_7238,N_2188,N_4352);
nand U7239 (N_7239,N_293,N_623);
and U7240 (N_7240,N_4109,N_580);
and U7241 (N_7241,N_715,N_2683);
and U7242 (N_7242,N_252,N_168);
nand U7243 (N_7243,N_4934,N_730);
and U7244 (N_7244,N_4719,N_3148);
nand U7245 (N_7245,N_1155,N_3869);
xor U7246 (N_7246,N_1205,N_831);
nand U7247 (N_7247,N_2142,N_3116);
or U7248 (N_7248,N_4096,N_3272);
nor U7249 (N_7249,N_2069,N_1468);
nor U7250 (N_7250,N_2831,N_2205);
nor U7251 (N_7251,N_4268,N_3396);
or U7252 (N_7252,N_763,N_3095);
nand U7253 (N_7253,N_2159,N_4128);
nor U7254 (N_7254,N_2565,N_2894);
nand U7255 (N_7255,N_2530,N_6);
or U7256 (N_7256,N_4750,N_4181);
xor U7257 (N_7257,N_942,N_1877);
nand U7258 (N_7258,N_1234,N_479);
and U7259 (N_7259,N_499,N_3903);
or U7260 (N_7260,N_964,N_201);
or U7261 (N_7261,N_4588,N_2246);
and U7262 (N_7262,N_2268,N_4651);
and U7263 (N_7263,N_4216,N_2448);
xor U7264 (N_7264,N_2461,N_4712);
nand U7265 (N_7265,N_1811,N_3999);
and U7266 (N_7266,N_1669,N_684);
nand U7267 (N_7267,N_437,N_3451);
nor U7268 (N_7268,N_4480,N_2820);
nand U7269 (N_7269,N_1890,N_4138);
nand U7270 (N_7270,N_3385,N_2846);
nand U7271 (N_7271,N_4526,N_2659);
and U7272 (N_7272,N_3223,N_1798);
or U7273 (N_7273,N_4272,N_2654);
or U7274 (N_7274,N_858,N_4851);
nand U7275 (N_7275,N_3741,N_521);
nor U7276 (N_7276,N_2865,N_2422);
nand U7277 (N_7277,N_17,N_4485);
or U7278 (N_7278,N_475,N_3174);
xnor U7279 (N_7279,N_3972,N_611);
and U7280 (N_7280,N_3557,N_3397);
or U7281 (N_7281,N_1013,N_3333);
xnor U7282 (N_7282,N_2397,N_4943);
or U7283 (N_7283,N_4303,N_1111);
nand U7284 (N_7284,N_4503,N_2196);
nor U7285 (N_7285,N_4146,N_1164);
nand U7286 (N_7286,N_3962,N_3322);
and U7287 (N_7287,N_1992,N_1443);
nand U7288 (N_7288,N_4144,N_1027);
nor U7289 (N_7289,N_1790,N_1770);
or U7290 (N_7290,N_774,N_308);
nand U7291 (N_7291,N_1734,N_2359);
xnor U7292 (N_7292,N_3828,N_176);
nand U7293 (N_7293,N_4870,N_140);
nor U7294 (N_7294,N_88,N_3373);
and U7295 (N_7295,N_4165,N_2813);
or U7296 (N_7296,N_3924,N_3268);
or U7297 (N_7297,N_406,N_4003);
xor U7298 (N_7298,N_1525,N_649);
nand U7299 (N_7299,N_719,N_4899);
and U7300 (N_7300,N_2636,N_4471);
nand U7301 (N_7301,N_523,N_3964);
nor U7302 (N_7302,N_4571,N_2890);
and U7303 (N_7303,N_4341,N_4534);
nor U7304 (N_7304,N_2895,N_645);
nor U7305 (N_7305,N_4269,N_2544);
xnor U7306 (N_7306,N_4766,N_3582);
nor U7307 (N_7307,N_4582,N_3854);
or U7308 (N_7308,N_1592,N_2078);
nor U7309 (N_7309,N_221,N_2891);
nand U7310 (N_7310,N_2973,N_1367);
nand U7311 (N_7311,N_3683,N_4991);
or U7312 (N_7312,N_1731,N_1688);
nor U7313 (N_7313,N_2646,N_2027);
nand U7314 (N_7314,N_1232,N_466);
or U7315 (N_7315,N_2942,N_3178);
nor U7316 (N_7316,N_4998,N_2074);
and U7317 (N_7317,N_1512,N_1444);
or U7318 (N_7318,N_2582,N_86);
nor U7319 (N_7319,N_4597,N_134);
nor U7320 (N_7320,N_524,N_2203);
xnor U7321 (N_7321,N_750,N_573);
nor U7322 (N_7322,N_4458,N_481);
xor U7323 (N_7323,N_4288,N_3520);
nor U7324 (N_7324,N_1416,N_3955);
xnor U7325 (N_7325,N_278,N_298);
xor U7326 (N_7326,N_4760,N_4675);
and U7327 (N_7327,N_4550,N_551);
nor U7328 (N_7328,N_435,N_1466);
and U7329 (N_7329,N_1604,N_1314);
or U7330 (N_7330,N_3645,N_2200);
and U7331 (N_7331,N_3382,N_3538);
and U7332 (N_7332,N_4451,N_1819);
or U7333 (N_7333,N_4854,N_3670);
and U7334 (N_7334,N_4740,N_488);
and U7335 (N_7335,N_1889,N_490);
and U7336 (N_7336,N_1442,N_2779);
nand U7337 (N_7337,N_800,N_328);
nand U7338 (N_7338,N_4472,N_3156);
or U7339 (N_7339,N_4829,N_1715);
xor U7340 (N_7340,N_3912,N_2297);
nand U7341 (N_7341,N_182,N_4289);
or U7342 (N_7342,N_1641,N_4450);
xnor U7343 (N_7343,N_4607,N_4877);
or U7344 (N_7344,N_3881,N_4957);
nor U7345 (N_7345,N_777,N_3091);
nor U7346 (N_7346,N_1612,N_4040);
nor U7347 (N_7347,N_4876,N_1284);
and U7348 (N_7348,N_3995,N_1460);
nor U7349 (N_7349,N_668,N_822);
nor U7350 (N_7350,N_3980,N_4999);
and U7351 (N_7351,N_4182,N_2559);
and U7352 (N_7352,N_3350,N_1021);
nor U7353 (N_7353,N_213,N_3251);
or U7354 (N_7354,N_446,N_4392);
xor U7355 (N_7355,N_3733,N_3374);
and U7356 (N_7356,N_639,N_4021);
or U7357 (N_7357,N_3338,N_3082);
or U7358 (N_7358,N_3742,N_1943);
or U7359 (N_7359,N_1788,N_4283);
and U7360 (N_7360,N_3807,N_4193);
and U7361 (N_7361,N_2031,N_3882);
nand U7362 (N_7362,N_2974,N_617);
nor U7363 (N_7363,N_557,N_2064);
nand U7364 (N_7364,N_576,N_3235);
or U7365 (N_7365,N_922,N_2804);
nor U7366 (N_7366,N_3393,N_4460);
nor U7367 (N_7367,N_2391,N_1297);
xnor U7368 (N_7368,N_927,N_3111);
nor U7369 (N_7369,N_3637,N_1548);
nand U7370 (N_7370,N_223,N_2472);
nand U7371 (N_7371,N_4274,N_2570);
and U7372 (N_7372,N_1498,N_2627);
and U7373 (N_7373,N_3992,N_2446);
nand U7374 (N_7374,N_2578,N_1958);
nand U7375 (N_7375,N_4674,N_3113);
or U7376 (N_7376,N_4827,N_2389);
nor U7377 (N_7377,N_4826,N_1725);
nand U7378 (N_7378,N_2674,N_2146);
nand U7379 (N_7379,N_2774,N_2995);
nor U7380 (N_7380,N_2723,N_3184);
or U7381 (N_7381,N_4646,N_3204);
and U7382 (N_7382,N_2287,N_3933);
nor U7383 (N_7383,N_2332,N_920);
nor U7384 (N_7384,N_2509,N_616);
or U7385 (N_7385,N_2044,N_3975);
xor U7386 (N_7386,N_4399,N_2528);
nand U7387 (N_7387,N_3885,N_4300);
nand U7388 (N_7388,N_905,N_1716);
and U7389 (N_7389,N_2424,N_3844);
nor U7390 (N_7390,N_1118,N_3724);
nor U7391 (N_7391,N_4004,N_2102);
nand U7392 (N_7392,N_1954,N_2861);
or U7393 (N_7393,N_4497,N_1041);
or U7394 (N_7394,N_1933,N_188);
or U7395 (N_7395,N_2170,N_1989);
and U7396 (N_7396,N_1680,N_791);
nand U7397 (N_7397,N_3959,N_3284);
nand U7398 (N_7398,N_1262,N_2719);
and U7399 (N_7399,N_1523,N_3914);
xor U7400 (N_7400,N_1686,N_2550);
nand U7401 (N_7401,N_923,N_1264);
and U7402 (N_7402,N_1894,N_1011);
xor U7403 (N_7403,N_1720,N_1228);
nand U7404 (N_7404,N_230,N_4002);
or U7405 (N_7405,N_2194,N_926);
and U7406 (N_7406,N_632,N_2486);
nor U7407 (N_7407,N_860,N_4351);
or U7408 (N_7408,N_4865,N_841);
or U7409 (N_7409,N_240,N_4951);
nand U7410 (N_7410,N_1028,N_2922);
or U7411 (N_7411,N_219,N_1654);
nand U7412 (N_7412,N_4377,N_72);
and U7413 (N_7413,N_4416,N_1053);
nor U7414 (N_7414,N_2699,N_997);
nand U7415 (N_7415,N_3118,N_779);
nand U7416 (N_7416,N_1170,N_4755);
nor U7417 (N_7417,N_1481,N_4252);
nand U7418 (N_7418,N_4585,N_1274);
or U7419 (N_7419,N_1174,N_4985);
nand U7420 (N_7420,N_2055,N_23);
and U7421 (N_7421,N_1755,N_961);
xor U7422 (N_7422,N_4662,N_1599);
nor U7423 (N_7423,N_291,N_3411);
xnor U7424 (N_7424,N_1553,N_75);
and U7425 (N_7425,N_2560,N_4426);
and U7426 (N_7426,N_378,N_4688);
or U7427 (N_7427,N_1983,N_1117);
nor U7428 (N_7428,N_4522,N_558);
nor U7429 (N_7429,N_1777,N_3275);
and U7430 (N_7430,N_1928,N_2262);
and U7431 (N_7431,N_3158,N_863);
nor U7432 (N_7432,N_1276,N_1951);
nand U7433 (N_7433,N_3916,N_4772);
nand U7434 (N_7434,N_4803,N_1948);
xor U7435 (N_7435,N_991,N_2348);
and U7436 (N_7436,N_2226,N_2619);
and U7437 (N_7437,N_2672,N_3597);
nor U7438 (N_7438,N_4931,N_2392);
nor U7439 (N_7439,N_1154,N_1645);
nor U7440 (N_7440,N_1618,N_933);
xnor U7441 (N_7441,N_2517,N_1366);
or U7442 (N_7442,N_2273,N_4990);
nand U7443 (N_7443,N_3680,N_754);
or U7444 (N_7444,N_4126,N_3642);
or U7445 (N_7445,N_3547,N_1301);
nand U7446 (N_7446,N_560,N_1323);
and U7447 (N_7447,N_3879,N_3228);
and U7448 (N_7448,N_957,N_4684);
and U7449 (N_7449,N_808,N_2938);
nand U7450 (N_7450,N_2658,N_2465);
and U7451 (N_7451,N_2265,N_4514);
nand U7452 (N_7452,N_3131,N_129);
or U7453 (N_7453,N_989,N_74);
xnor U7454 (N_7454,N_1360,N_2437);
nor U7455 (N_7455,N_360,N_1472);
nand U7456 (N_7456,N_4543,N_1245);
xor U7457 (N_7457,N_1806,N_2125);
or U7458 (N_7458,N_4950,N_2828);
xnor U7459 (N_7459,N_1307,N_2900);
and U7460 (N_7460,N_1294,N_3731);
nand U7461 (N_7461,N_1650,N_2028);
and U7462 (N_7462,N_4106,N_3361);
and U7463 (N_7463,N_739,N_3024);
or U7464 (N_7464,N_2910,N_2652);
or U7465 (N_7465,N_4516,N_329);
nand U7466 (N_7466,N_1926,N_3318);
nor U7467 (N_7467,N_123,N_861);
xor U7468 (N_7468,N_2823,N_2459);
nor U7469 (N_7469,N_3769,N_2977);
and U7470 (N_7470,N_4707,N_1756);
and U7471 (N_7471,N_1586,N_2819);
xor U7472 (N_7472,N_3772,N_3059);
or U7473 (N_7473,N_1647,N_2316);
nand U7474 (N_7474,N_4744,N_2787);
and U7475 (N_7475,N_673,N_3673);
nor U7476 (N_7476,N_4221,N_1702);
nor U7477 (N_7477,N_2115,N_4086);
or U7478 (N_7478,N_682,N_840);
nor U7479 (N_7479,N_983,N_2260);
nor U7480 (N_7480,N_3472,N_776);
nor U7481 (N_7481,N_2445,N_228);
or U7482 (N_7482,N_3524,N_32);
nand U7483 (N_7483,N_26,N_3612);
or U7484 (N_7484,N_4332,N_1493);
nor U7485 (N_7485,N_1003,N_2413);
and U7486 (N_7486,N_4378,N_2810);
nor U7487 (N_7487,N_2825,N_418);
nand U7488 (N_7488,N_4358,N_959);
nor U7489 (N_7489,N_4777,N_4229);
or U7490 (N_7490,N_1409,N_4964);
and U7491 (N_7491,N_3908,N_1353);
nand U7492 (N_7492,N_2400,N_656);
xor U7493 (N_7493,N_11,N_3715);
and U7494 (N_7494,N_3395,N_3970);
or U7495 (N_7495,N_4062,N_1666);
or U7496 (N_7496,N_3483,N_1968);
nor U7497 (N_7497,N_3303,N_3405);
nor U7498 (N_7498,N_1538,N_1097);
nand U7499 (N_7499,N_3152,N_447);
nand U7500 (N_7500,N_915,N_416);
and U7501 (N_7501,N_3365,N_1223);
xnor U7502 (N_7502,N_3758,N_687);
or U7503 (N_7503,N_352,N_2140);
xor U7504 (N_7504,N_656,N_2707);
or U7505 (N_7505,N_959,N_4547);
nor U7506 (N_7506,N_2094,N_1351);
and U7507 (N_7507,N_1694,N_3504);
or U7508 (N_7508,N_1303,N_3168);
and U7509 (N_7509,N_4161,N_1626);
and U7510 (N_7510,N_1887,N_1330);
and U7511 (N_7511,N_4245,N_4436);
or U7512 (N_7512,N_1074,N_62);
or U7513 (N_7513,N_1201,N_4752);
nor U7514 (N_7514,N_928,N_4930);
nor U7515 (N_7515,N_180,N_4042);
or U7516 (N_7516,N_2907,N_3447);
and U7517 (N_7517,N_929,N_2350);
nand U7518 (N_7518,N_4837,N_2554);
and U7519 (N_7519,N_3039,N_2222);
and U7520 (N_7520,N_502,N_773);
nor U7521 (N_7521,N_3024,N_1952);
or U7522 (N_7522,N_1300,N_2744);
nand U7523 (N_7523,N_1440,N_4168);
or U7524 (N_7524,N_699,N_4581);
nand U7525 (N_7525,N_4891,N_748);
and U7526 (N_7526,N_3281,N_1348);
nor U7527 (N_7527,N_3312,N_3476);
nand U7528 (N_7528,N_4885,N_235);
nor U7529 (N_7529,N_2815,N_2768);
nand U7530 (N_7530,N_3372,N_2387);
and U7531 (N_7531,N_2569,N_814);
nand U7532 (N_7532,N_1810,N_1610);
and U7533 (N_7533,N_3459,N_1539);
or U7534 (N_7534,N_3961,N_4822);
and U7535 (N_7535,N_4307,N_4309);
nor U7536 (N_7536,N_4283,N_121);
nand U7537 (N_7537,N_18,N_3452);
or U7538 (N_7538,N_4945,N_1270);
and U7539 (N_7539,N_2199,N_4546);
and U7540 (N_7540,N_1361,N_645);
nor U7541 (N_7541,N_2025,N_954);
nand U7542 (N_7542,N_1897,N_2412);
nand U7543 (N_7543,N_3544,N_4788);
xnor U7544 (N_7544,N_4781,N_2630);
nand U7545 (N_7545,N_1593,N_344);
nand U7546 (N_7546,N_2940,N_1911);
nor U7547 (N_7547,N_2909,N_4542);
or U7548 (N_7548,N_1179,N_4012);
and U7549 (N_7549,N_2317,N_222);
or U7550 (N_7550,N_4022,N_2413);
and U7551 (N_7551,N_2611,N_3858);
nand U7552 (N_7552,N_4644,N_4304);
nand U7553 (N_7553,N_2833,N_1681);
nor U7554 (N_7554,N_1348,N_2009);
or U7555 (N_7555,N_4430,N_630);
and U7556 (N_7556,N_1114,N_1907);
nor U7557 (N_7557,N_4293,N_3907);
nor U7558 (N_7558,N_1766,N_1119);
nor U7559 (N_7559,N_2269,N_713);
or U7560 (N_7560,N_3627,N_2459);
nand U7561 (N_7561,N_2691,N_4300);
nand U7562 (N_7562,N_4134,N_1247);
xor U7563 (N_7563,N_4414,N_726);
and U7564 (N_7564,N_3449,N_2977);
or U7565 (N_7565,N_80,N_1496);
or U7566 (N_7566,N_1038,N_2535);
nor U7567 (N_7567,N_317,N_1888);
nor U7568 (N_7568,N_986,N_1225);
nand U7569 (N_7569,N_204,N_3884);
or U7570 (N_7570,N_1038,N_1568);
or U7571 (N_7571,N_3533,N_324);
xnor U7572 (N_7572,N_1111,N_1144);
or U7573 (N_7573,N_3084,N_4610);
or U7574 (N_7574,N_2654,N_4298);
or U7575 (N_7575,N_4661,N_4557);
and U7576 (N_7576,N_1887,N_1082);
and U7577 (N_7577,N_2075,N_2751);
or U7578 (N_7578,N_1842,N_404);
nor U7579 (N_7579,N_3664,N_2078);
xor U7580 (N_7580,N_3017,N_3225);
nor U7581 (N_7581,N_1403,N_656);
and U7582 (N_7582,N_1656,N_4989);
and U7583 (N_7583,N_712,N_2886);
and U7584 (N_7584,N_2391,N_3356);
nor U7585 (N_7585,N_350,N_401);
nand U7586 (N_7586,N_3813,N_1855);
and U7587 (N_7587,N_2408,N_1125);
nor U7588 (N_7588,N_4341,N_2181);
nand U7589 (N_7589,N_3598,N_3190);
or U7590 (N_7590,N_65,N_2482);
or U7591 (N_7591,N_4726,N_622);
and U7592 (N_7592,N_4962,N_4854);
nand U7593 (N_7593,N_1408,N_4677);
and U7594 (N_7594,N_2372,N_2561);
or U7595 (N_7595,N_134,N_658);
or U7596 (N_7596,N_3305,N_3300);
xor U7597 (N_7597,N_4709,N_846);
nand U7598 (N_7598,N_1739,N_3319);
xnor U7599 (N_7599,N_4911,N_4553);
nor U7600 (N_7600,N_3295,N_4726);
or U7601 (N_7601,N_3215,N_466);
and U7602 (N_7602,N_1288,N_4870);
xor U7603 (N_7603,N_1738,N_4771);
nand U7604 (N_7604,N_592,N_4926);
and U7605 (N_7605,N_1057,N_2335);
nor U7606 (N_7606,N_11,N_3200);
xnor U7607 (N_7607,N_1003,N_2960);
and U7608 (N_7608,N_3377,N_1296);
nor U7609 (N_7609,N_4683,N_2452);
nand U7610 (N_7610,N_4125,N_585);
or U7611 (N_7611,N_3694,N_1414);
or U7612 (N_7612,N_2663,N_600);
xnor U7613 (N_7613,N_1915,N_3297);
nand U7614 (N_7614,N_1177,N_833);
or U7615 (N_7615,N_4073,N_675);
or U7616 (N_7616,N_2575,N_1707);
or U7617 (N_7617,N_1451,N_859);
nand U7618 (N_7618,N_2714,N_4380);
nand U7619 (N_7619,N_4432,N_3130);
and U7620 (N_7620,N_503,N_1963);
nand U7621 (N_7621,N_3070,N_2435);
nand U7622 (N_7622,N_664,N_3146);
nor U7623 (N_7623,N_2281,N_2225);
xor U7624 (N_7624,N_2700,N_3283);
and U7625 (N_7625,N_399,N_694);
or U7626 (N_7626,N_532,N_4302);
and U7627 (N_7627,N_2410,N_4721);
or U7628 (N_7628,N_2298,N_4238);
nand U7629 (N_7629,N_3589,N_3942);
or U7630 (N_7630,N_4214,N_1732);
or U7631 (N_7631,N_3998,N_2365);
or U7632 (N_7632,N_265,N_3338);
and U7633 (N_7633,N_1427,N_2125);
and U7634 (N_7634,N_2155,N_1667);
and U7635 (N_7635,N_1388,N_3740);
and U7636 (N_7636,N_1755,N_2742);
and U7637 (N_7637,N_4767,N_1693);
nor U7638 (N_7638,N_344,N_3274);
or U7639 (N_7639,N_4944,N_984);
and U7640 (N_7640,N_1292,N_1678);
nor U7641 (N_7641,N_4717,N_3104);
and U7642 (N_7642,N_1253,N_3338);
nor U7643 (N_7643,N_2214,N_998);
nor U7644 (N_7644,N_3062,N_16);
nand U7645 (N_7645,N_2794,N_1239);
and U7646 (N_7646,N_2105,N_2877);
nor U7647 (N_7647,N_220,N_1921);
and U7648 (N_7648,N_4470,N_667);
nand U7649 (N_7649,N_3143,N_132);
nor U7650 (N_7650,N_2415,N_1416);
nor U7651 (N_7651,N_4493,N_2871);
nor U7652 (N_7652,N_4207,N_1825);
nand U7653 (N_7653,N_4987,N_2);
and U7654 (N_7654,N_2808,N_928);
nand U7655 (N_7655,N_270,N_861);
or U7656 (N_7656,N_4823,N_292);
nand U7657 (N_7657,N_4911,N_791);
and U7658 (N_7658,N_4727,N_4658);
and U7659 (N_7659,N_3454,N_4549);
and U7660 (N_7660,N_97,N_1712);
and U7661 (N_7661,N_2064,N_19);
nand U7662 (N_7662,N_1572,N_3064);
and U7663 (N_7663,N_533,N_440);
xor U7664 (N_7664,N_1218,N_156);
or U7665 (N_7665,N_4842,N_17);
and U7666 (N_7666,N_976,N_556);
nor U7667 (N_7667,N_3642,N_633);
nand U7668 (N_7668,N_1966,N_3111);
nand U7669 (N_7669,N_3625,N_1407);
or U7670 (N_7670,N_2704,N_3976);
or U7671 (N_7671,N_4290,N_3208);
or U7672 (N_7672,N_591,N_2508);
nor U7673 (N_7673,N_3051,N_2897);
or U7674 (N_7674,N_1767,N_4706);
and U7675 (N_7675,N_1231,N_4644);
nand U7676 (N_7676,N_3049,N_2602);
nand U7677 (N_7677,N_291,N_4771);
and U7678 (N_7678,N_2576,N_459);
or U7679 (N_7679,N_4974,N_24);
or U7680 (N_7680,N_127,N_1389);
xnor U7681 (N_7681,N_1423,N_1607);
and U7682 (N_7682,N_4687,N_2331);
or U7683 (N_7683,N_513,N_4066);
nor U7684 (N_7684,N_2634,N_1869);
nor U7685 (N_7685,N_736,N_3772);
xor U7686 (N_7686,N_1850,N_4262);
and U7687 (N_7687,N_4927,N_845);
xor U7688 (N_7688,N_737,N_2893);
nand U7689 (N_7689,N_2001,N_1851);
and U7690 (N_7690,N_3420,N_1884);
xnor U7691 (N_7691,N_1030,N_251);
nor U7692 (N_7692,N_823,N_2039);
and U7693 (N_7693,N_603,N_4669);
or U7694 (N_7694,N_1363,N_2210);
and U7695 (N_7695,N_3476,N_916);
nand U7696 (N_7696,N_567,N_623);
nand U7697 (N_7697,N_3621,N_2218);
and U7698 (N_7698,N_4163,N_4778);
nor U7699 (N_7699,N_1643,N_794);
and U7700 (N_7700,N_1057,N_890);
nor U7701 (N_7701,N_3268,N_3823);
or U7702 (N_7702,N_541,N_3958);
nand U7703 (N_7703,N_105,N_1225);
or U7704 (N_7704,N_886,N_3521);
or U7705 (N_7705,N_3042,N_1178);
nor U7706 (N_7706,N_4767,N_3478);
xnor U7707 (N_7707,N_3099,N_4877);
nand U7708 (N_7708,N_886,N_33);
or U7709 (N_7709,N_3323,N_3770);
nand U7710 (N_7710,N_4505,N_485);
or U7711 (N_7711,N_3389,N_1568);
or U7712 (N_7712,N_1547,N_93);
nor U7713 (N_7713,N_3130,N_779);
nand U7714 (N_7714,N_3603,N_4383);
nand U7715 (N_7715,N_1607,N_1593);
or U7716 (N_7716,N_1414,N_4066);
and U7717 (N_7717,N_1729,N_2991);
nor U7718 (N_7718,N_4161,N_143);
and U7719 (N_7719,N_947,N_2752);
xnor U7720 (N_7720,N_445,N_3311);
and U7721 (N_7721,N_3472,N_3780);
or U7722 (N_7722,N_4381,N_2803);
or U7723 (N_7723,N_1844,N_3775);
nand U7724 (N_7724,N_2187,N_719);
xnor U7725 (N_7725,N_4264,N_1055);
nor U7726 (N_7726,N_3438,N_1114);
nand U7727 (N_7727,N_4018,N_2820);
and U7728 (N_7728,N_1484,N_3096);
or U7729 (N_7729,N_2380,N_3674);
nor U7730 (N_7730,N_4306,N_2483);
and U7731 (N_7731,N_213,N_3709);
or U7732 (N_7732,N_2926,N_1036);
and U7733 (N_7733,N_449,N_3551);
nand U7734 (N_7734,N_2296,N_175);
and U7735 (N_7735,N_1017,N_859);
xor U7736 (N_7736,N_2779,N_2715);
or U7737 (N_7737,N_822,N_682);
or U7738 (N_7738,N_4668,N_2837);
or U7739 (N_7739,N_2998,N_1773);
or U7740 (N_7740,N_2459,N_2265);
nand U7741 (N_7741,N_1383,N_3180);
or U7742 (N_7742,N_4493,N_1750);
nor U7743 (N_7743,N_4916,N_3905);
nor U7744 (N_7744,N_2998,N_881);
and U7745 (N_7745,N_2271,N_1597);
nor U7746 (N_7746,N_674,N_4232);
nor U7747 (N_7747,N_1134,N_3333);
xnor U7748 (N_7748,N_1294,N_1375);
nor U7749 (N_7749,N_1405,N_1052);
or U7750 (N_7750,N_4831,N_2968);
nor U7751 (N_7751,N_2150,N_4913);
nand U7752 (N_7752,N_4692,N_3989);
and U7753 (N_7753,N_4223,N_4082);
nor U7754 (N_7754,N_1545,N_2204);
xnor U7755 (N_7755,N_1644,N_1280);
nand U7756 (N_7756,N_4772,N_2718);
and U7757 (N_7757,N_2071,N_3900);
nand U7758 (N_7758,N_3075,N_358);
and U7759 (N_7759,N_2869,N_4817);
and U7760 (N_7760,N_4647,N_73);
nand U7761 (N_7761,N_4196,N_4883);
or U7762 (N_7762,N_3192,N_1053);
nand U7763 (N_7763,N_4684,N_3021);
nor U7764 (N_7764,N_3179,N_2117);
nor U7765 (N_7765,N_554,N_4455);
and U7766 (N_7766,N_3876,N_3737);
and U7767 (N_7767,N_898,N_2413);
and U7768 (N_7768,N_905,N_3253);
nor U7769 (N_7769,N_3220,N_4558);
and U7770 (N_7770,N_1165,N_1173);
nor U7771 (N_7771,N_4259,N_3405);
and U7772 (N_7772,N_465,N_2963);
and U7773 (N_7773,N_3982,N_4100);
nand U7774 (N_7774,N_198,N_4993);
nor U7775 (N_7775,N_519,N_2226);
nand U7776 (N_7776,N_777,N_3283);
and U7777 (N_7777,N_4224,N_781);
and U7778 (N_7778,N_3678,N_4739);
or U7779 (N_7779,N_431,N_3018);
and U7780 (N_7780,N_2554,N_407);
nand U7781 (N_7781,N_3807,N_2866);
or U7782 (N_7782,N_3932,N_3367);
or U7783 (N_7783,N_2979,N_3073);
nand U7784 (N_7784,N_1436,N_99);
and U7785 (N_7785,N_4573,N_2394);
xnor U7786 (N_7786,N_708,N_3230);
and U7787 (N_7787,N_1209,N_3094);
nor U7788 (N_7788,N_3236,N_1754);
and U7789 (N_7789,N_3140,N_1832);
nand U7790 (N_7790,N_4600,N_230);
nor U7791 (N_7791,N_3637,N_1337);
xnor U7792 (N_7792,N_667,N_324);
nand U7793 (N_7793,N_1662,N_1087);
nor U7794 (N_7794,N_4610,N_1926);
or U7795 (N_7795,N_3561,N_2446);
xnor U7796 (N_7796,N_1686,N_2642);
nor U7797 (N_7797,N_1238,N_175);
nand U7798 (N_7798,N_3533,N_4594);
or U7799 (N_7799,N_2215,N_167);
nor U7800 (N_7800,N_3449,N_2807);
and U7801 (N_7801,N_3848,N_4442);
and U7802 (N_7802,N_1,N_3208);
xnor U7803 (N_7803,N_1372,N_4962);
nor U7804 (N_7804,N_2837,N_1134);
or U7805 (N_7805,N_3754,N_4637);
nor U7806 (N_7806,N_2354,N_1025);
nor U7807 (N_7807,N_4693,N_460);
or U7808 (N_7808,N_4232,N_2878);
nor U7809 (N_7809,N_201,N_1926);
or U7810 (N_7810,N_164,N_4553);
nor U7811 (N_7811,N_2884,N_2043);
or U7812 (N_7812,N_246,N_2928);
nand U7813 (N_7813,N_2923,N_4887);
nor U7814 (N_7814,N_3294,N_3001);
and U7815 (N_7815,N_4142,N_2759);
nand U7816 (N_7816,N_1128,N_1179);
and U7817 (N_7817,N_446,N_713);
nor U7818 (N_7818,N_4676,N_360);
nand U7819 (N_7819,N_886,N_3784);
nor U7820 (N_7820,N_4863,N_3798);
or U7821 (N_7821,N_160,N_4572);
and U7822 (N_7822,N_3859,N_978);
or U7823 (N_7823,N_1571,N_2547);
and U7824 (N_7824,N_587,N_619);
nand U7825 (N_7825,N_3593,N_3534);
nor U7826 (N_7826,N_2468,N_3076);
or U7827 (N_7827,N_1294,N_2906);
nand U7828 (N_7828,N_1667,N_52);
and U7829 (N_7829,N_3021,N_3599);
nor U7830 (N_7830,N_671,N_4675);
or U7831 (N_7831,N_3739,N_807);
and U7832 (N_7832,N_3848,N_1054);
and U7833 (N_7833,N_1256,N_2679);
nand U7834 (N_7834,N_2361,N_3294);
and U7835 (N_7835,N_1910,N_4177);
or U7836 (N_7836,N_3532,N_3117);
nor U7837 (N_7837,N_3552,N_2907);
or U7838 (N_7838,N_1942,N_4435);
xnor U7839 (N_7839,N_4088,N_4541);
or U7840 (N_7840,N_3606,N_112);
or U7841 (N_7841,N_1875,N_3054);
nand U7842 (N_7842,N_3230,N_716);
and U7843 (N_7843,N_2714,N_3382);
and U7844 (N_7844,N_1736,N_1413);
or U7845 (N_7845,N_2623,N_264);
nor U7846 (N_7846,N_3684,N_1822);
nand U7847 (N_7847,N_1727,N_203);
and U7848 (N_7848,N_465,N_2080);
nand U7849 (N_7849,N_1581,N_3064);
and U7850 (N_7850,N_3941,N_4946);
nand U7851 (N_7851,N_1124,N_418);
xnor U7852 (N_7852,N_2981,N_4976);
nand U7853 (N_7853,N_3390,N_224);
nand U7854 (N_7854,N_1120,N_3989);
xor U7855 (N_7855,N_149,N_4315);
or U7856 (N_7856,N_4165,N_4937);
nor U7857 (N_7857,N_936,N_3096);
and U7858 (N_7858,N_2822,N_973);
or U7859 (N_7859,N_1121,N_2565);
xor U7860 (N_7860,N_2246,N_4748);
or U7861 (N_7861,N_1026,N_1687);
or U7862 (N_7862,N_2480,N_3507);
nand U7863 (N_7863,N_420,N_1695);
and U7864 (N_7864,N_622,N_1702);
nand U7865 (N_7865,N_4561,N_686);
or U7866 (N_7866,N_419,N_3296);
or U7867 (N_7867,N_562,N_4473);
or U7868 (N_7868,N_392,N_2165);
nand U7869 (N_7869,N_2479,N_1385);
nand U7870 (N_7870,N_4281,N_2414);
or U7871 (N_7871,N_152,N_2109);
nor U7872 (N_7872,N_4109,N_2177);
nor U7873 (N_7873,N_2192,N_4684);
or U7874 (N_7874,N_808,N_1037);
nand U7875 (N_7875,N_1309,N_1218);
and U7876 (N_7876,N_729,N_2967);
or U7877 (N_7877,N_2622,N_3553);
or U7878 (N_7878,N_2390,N_4849);
nand U7879 (N_7879,N_2024,N_2002);
nand U7880 (N_7880,N_3532,N_919);
or U7881 (N_7881,N_2887,N_513);
and U7882 (N_7882,N_3500,N_1943);
and U7883 (N_7883,N_520,N_2449);
or U7884 (N_7884,N_4078,N_2700);
nand U7885 (N_7885,N_4202,N_603);
or U7886 (N_7886,N_1952,N_1864);
and U7887 (N_7887,N_3096,N_2401);
and U7888 (N_7888,N_4980,N_591);
xor U7889 (N_7889,N_2266,N_2306);
nand U7890 (N_7890,N_2367,N_1188);
xor U7891 (N_7891,N_127,N_2123);
nand U7892 (N_7892,N_4345,N_3575);
or U7893 (N_7893,N_2658,N_4500);
and U7894 (N_7894,N_3326,N_3259);
nand U7895 (N_7895,N_2025,N_1750);
or U7896 (N_7896,N_4876,N_2547);
or U7897 (N_7897,N_689,N_1332);
nor U7898 (N_7898,N_965,N_3669);
or U7899 (N_7899,N_1145,N_3610);
or U7900 (N_7900,N_2585,N_1871);
nand U7901 (N_7901,N_4112,N_941);
and U7902 (N_7902,N_1135,N_3670);
and U7903 (N_7903,N_3970,N_1534);
nand U7904 (N_7904,N_3011,N_3186);
nor U7905 (N_7905,N_1299,N_2852);
nor U7906 (N_7906,N_2637,N_3235);
or U7907 (N_7907,N_764,N_316);
or U7908 (N_7908,N_3465,N_1727);
nand U7909 (N_7909,N_4171,N_1788);
and U7910 (N_7910,N_2065,N_2120);
and U7911 (N_7911,N_3847,N_4297);
nand U7912 (N_7912,N_651,N_2038);
or U7913 (N_7913,N_1074,N_1020);
or U7914 (N_7914,N_3966,N_3019);
xor U7915 (N_7915,N_4039,N_4861);
nor U7916 (N_7916,N_2550,N_296);
or U7917 (N_7917,N_4545,N_865);
nor U7918 (N_7918,N_2681,N_596);
or U7919 (N_7919,N_4532,N_4345);
or U7920 (N_7920,N_2956,N_4103);
or U7921 (N_7921,N_3661,N_402);
or U7922 (N_7922,N_2896,N_3883);
xnor U7923 (N_7923,N_359,N_3069);
and U7924 (N_7924,N_3957,N_4195);
nor U7925 (N_7925,N_1631,N_3618);
nand U7926 (N_7926,N_868,N_398);
or U7927 (N_7927,N_1773,N_1739);
and U7928 (N_7928,N_2231,N_143);
nand U7929 (N_7929,N_3283,N_3242);
or U7930 (N_7930,N_3237,N_780);
and U7931 (N_7931,N_4663,N_4338);
nand U7932 (N_7932,N_2017,N_1695);
and U7933 (N_7933,N_4068,N_1091);
or U7934 (N_7934,N_506,N_4898);
or U7935 (N_7935,N_2889,N_4218);
and U7936 (N_7936,N_3584,N_2894);
xnor U7937 (N_7937,N_4895,N_3458);
nand U7938 (N_7938,N_1752,N_230);
nand U7939 (N_7939,N_391,N_3179);
nand U7940 (N_7940,N_4700,N_368);
nor U7941 (N_7941,N_4706,N_4508);
and U7942 (N_7942,N_575,N_2059);
xnor U7943 (N_7943,N_2259,N_1963);
and U7944 (N_7944,N_1991,N_3385);
and U7945 (N_7945,N_4149,N_322);
xor U7946 (N_7946,N_2742,N_1076);
nor U7947 (N_7947,N_2477,N_4179);
nand U7948 (N_7948,N_4817,N_3339);
nand U7949 (N_7949,N_4994,N_3634);
or U7950 (N_7950,N_3877,N_2825);
nor U7951 (N_7951,N_1890,N_4396);
nor U7952 (N_7952,N_545,N_2233);
or U7953 (N_7953,N_2340,N_4292);
nor U7954 (N_7954,N_217,N_3643);
or U7955 (N_7955,N_3666,N_1778);
nand U7956 (N_7956,N_594,N_1577);
nor U7957 (N_7957,N_831,N_686);
and U7958 (N_7958,N_1494,N_4398);
nor U7959 (N_7959,N_4240,N_3649);
or U7960 (N_7960,N_3121,N_938);
nor U7961 (N_7961,N_2752,N_3154);
and U7962 (N_7962,N_3134,N_659);
nand U7963 (N_7963,N_4556,N_1484);
nand U7964 (N_7964,N_832,N_2926);
and U7965 (N_7965,N_3741,N_3377);
and U7966 (N_7966,N_4740,N_2317);
nor U7967 (N_7967,N_4066,N_421);
nand U7968 (N_7968,N_2662,N_896);
nand U7969 (N_7969,N_540,N_2488);
or U7970 (N_7970,N_2558,N_2307);
nand U7971 (N_7971,N_3519,N_4492);
or U7972 (N_7972,N_1581,N_851);
or U7973 (N_7973,N_2640,N_3874);
and U7974 (N_7974,N_1541,N_3366);
or U7975 (N_7975,N_4619,N_1811);
and U7976 (N_7976,N_1323,N_2768);
or U7977 (N_7977,N_1553,N_1573);
or U7978 (N_7978,N_3235,N_900);
and U7979 (N_7979,N_588,N_2575);
nand U7980 (N_7980,N_2523,N_1303);
or U7981 (N_7981,N_1590,N_450);
nand U7982 (N_7982,N_802,N_684);
nor U7983 (N_7983,N_1030,N_1777);
and U7984 (N_7984,N_2271,N_1825);
nor U7985 (N_7985,N_4796,N_649);
nor U7986 (N_7986,N_4850,N_3566);
nand U7987 (N_7987,N_4811,N_3950);
nor U7988 (N_7988,N_2790,N_2087);
xnor U7989 (N_7989,N_982,N_913);
xnor U7990 (N_7990,N_2906,N_3647);
or U7991 (N_7991,N_3820,N_55);
nand U7992 (N_7992,N_4055,N_2210);
and U7993 (N_7993,N_1562,N_1009);
or U7994 (N_7994,N_4157,N_4786);
nor U7995 (N_7995,N_3473,N_252);
and U7996 (N_7996,N_3534,N_4037);
nand U7997 (N_7997,N_1251,N_1642);
or U7998 (N_7998,N_1357,N_3435);
xnor U7999 (N_7999,N_2369,N_1197);
nor U8000 (N_8000,N_1997,N_1573);
and U8001 (N_8001,N_1117,N_4242);
or U8002 (N_8002,N_2925,N_2744);
nand U8003 (N_8003,N_4668,N_2521);
nand U8004 (N_8004,N_1223,N_597);
or U8005 (N_8005,N_1071,N_3483);
or U8006 (N_8006,N_396,N_4353);
nand U8007 (N_8007,N_2158,N_4535);
and U8008 (N_8008,N_1412,N_3932);
xnor U8009 (N_8009,N_3193,N_2018);
xor U8010 (N_8010,N_104,N_2802);
xnor U8011 (N_8011,N_3083,N_3109);
nand U8012 (N_8012,N_2274,N_1985);
nor U8013 (N_8013,N_1692,N_4323);
nor U8014 (N_8014,N_1238,N_2738);
or U8015 (N_8015,N_4175,N_1808);
and U8016 (N_8016,N_4165,N_175);
and U8017 (N_8017,N_1477,N_1445);
xnor U8018 (N_8018,N_4408,N_2554);
or U8019 (N_8019,N_4775,N_4546);
and U8020 (N_8020,N_2901,N_4530);
or U8021 (N_8021,N_2774,N_1169);
nor U8022 (N_8022,N_1404,N_2680);
nand U8023 (N_8023,N_4486,N_4235);
and U8024 (N_8024,N_4273,N_849);
or U8025 (N_8025,N_1057,N_2774);
or U8026 (N_8026,N_119,N_2816);
nor U8027 (N_8027,N_112,N_2369);
or U8028 (N_8028,N_1203,N_1559);
or U8029 (N_8029,N_3069,N_2628);
nor U8030 (N_8030,N_2492,N_3974);
nor U8031 (N_8031,N_3083,N_3891);
and U8032 (N_8032,N_4466,N_1006);
nor U8033 (N_8033,N_3048,N_2522);
nand U8034 (N_8034,N_2626,N_1082);
nor U8035 (N_8035,N_4125,N_2078);
nor U8036 (N_8036,N_440,N_4640);
or U8037 (N_8037,N_1446,N_321);
nand U8038 (N_8038,N_2819,N_2222);
nand U8039 (N_8039,N_1935,N_3110);
and U8040 (N_8040,N_1640,N_98);
nor U8041 (N_8041,N_1849,N_3787);
nor U8042 (N_8042,N_2640,N_3882);
and U8043 (N_8043,N_4383,N_2789);
nor U8044 (N_8044,N_3361,N_1393);
xnor U8045 (N_8045,N_3360,N_2869);
and U8046 (N_8046,N_1354,N_590);
or U8047 (N_8047,N_581,N_1596);
or U8048 (N_8048,N_511,N_2956);
and U8049 (N_8049,N_308,N_1838);
and U8050 (N_8050,N_2943,N_3788);
xnor U8051 (N_8051,N_2548,N_3311);
nand U8052 (N_8052,N_4563,N_85);
xnor U8053 (N_8053,N_3647,N_3364);
nor U8054 (N_8054,N_1760,N_3247);
and U8055 (N_8055,N_3204,N_3673);
nand U8056 (N_8056,N_1142,N_4893);
nor U8057 (N_8057,N_482,N_637);
nor U8058 (N_8058,N_3786,N_3749);
xor U8059 (N_8059,N_3014,N_4578);
or U8060 (N_8060,N_333,N_2748);
xor U8061 (N_8061,N_4626,N_3216);
nand U8062 (N_8062,N_3600,N_3741);
nor U8063 (N_8063,N_1182,N_1385);
nand U8064 (N_8064,N_3177,N_4702);
and U8065 (N_8065,N_1270,N_1368);
and U8066 (N_8066,N_1273,N_2008);
and U8067 (N_8067,N_4053,N_3317);
and U8068 (N_8068,N_1661,N_4838);
xor U8069 (N_8069,N_108,N_2151);
or U8070 (N_8070,N_1437,N_4691);
or U8071 (N_8071,N_723,N_3848);
nor U8072 (N_8072,N_2405,N_3767);
and U8073 (N_8073,N_2247,N_3400);
nor U8074 (N_8074,N_278,N_3576);
nand U8075 (N_8075,N_2419,N_3304);
nor U8076 (N_8076,N_2752,N_429);
nand U8077 (N_8077,N_749,N_3993);
nor U8078 (N_8078,N_2338,N_1717);
nand U8079 (N_8079,N_4397,N_3080);
nor U8080 (N_8080,N_4859,N_4020);
nor U8081 (N_8081,N_2057,N_863);
nand U8082 (N_8082,N_3744,N_1291);
nand U8083 (N_8083,N_2021,N_1595);
and U8084 (N_8084,N_1387,N_4286);
or U8085 (N_8085,N_4776,N_2981);
xnor U8086 (N_8086,N_4908,N_1133);
nor U8087 (N_8087,N_1728,N_3312);
and U8088 (N_8088,N_565,N_1132);
and U8089 (N_8089,N_1968,N_2541);
or U8090 (N_8090,N_1665,N_2506);
xor U8091 (N_8091,N_3925,N_736);
nor U8092 (N_8092,N_3736,N_1778);
and U8093 (N_8093,N_2874,N_2582);
or U8094 (N_8094,N_427,N_4505);
and U8095 (N_8095,N_1214,N_485);
nor U8096 (N_8096,N_4300,N_3561);
nor U8097 (N_8097,N_1838,N_2232);
and U8098 (N_8098,N_4942,N_66);
nand U8099 (N_8099,N_3440,N_3720);
nand U8100 (N_8100,N_4694,N_1575);
xnor U8101 (N_8101,N_2264,N_904);
nand U8102 (N_8102,N_611,N_4753);
nand U8103 (N_8103,N_4491,N_1632);
or U8104 (N_8104,N_3898,N_1699);
nor U8105 (N_8105,N_3736,N_1725);
nor U8106 (N_8106,N_62,N_2931);
xnor U8107 (N_8107,N_3113,N_3800);
or U8108 (N_8108,N_791,N_2406);
nand U8109 (N_8109,N_973,N_3755);
nor U8110 (N_8110,N_4651,N_1712);
nand U8111 (N_8111,N_1500,N_2766);
and U8112 (N_8112,N_2274,N_24);
and U8113 (N_8113,N_1090,N_1143);
nor U8114 (N_8114,N_4249,N_224);
or U8115 (N_8115,N_1206,N_1897);
nor U8116 (N_8116,N_2295,N_13);
or U8117 (N_8117,N_1008,N_4480);
xor U8118 (N_8118,N_806,N_4777);
nand U8119 (N_8119,N_466,N_2563);
or U8120 (N_8120,N_4536,N_954);
nor U8121 (N_8121,N_3018,N_403);
nor U8122 (N_8122,N_4912,N_2365);
or U8123 (N_8123,N_3780,N_2064);
nand U8124 (N_8124,N_2022,N_165);
and U8125 (N_8125,N_3531,N_743);
and U8126 (N_8126,N_584,N_4519);
nor U8127 (N_8127,N_3280,N_2838);
nand U8128 (N_8128,N_46,N_592);
nand U8129 (N_8129,N_2870,N_2924);
nor U8130 (N_8130,N_522,N_1026);
and U8131 (N_8131,N_4856,N_4504);
or U8132 (N_8132,N_2929,N_3700);
and U8133 (N_8133,N_4308,N_17);
nand U8134 (N_8134,N_2591,N_2461);
or U8135 (N_8135,N_1801,N_3659);
nand U8136 (N_8136,N_3467,N_3816);
nand U8137 (N_8137,N_2480,N_1860);
nor U8138 (N_8138,N_467,N_2022);
nor U8139 (N_8139,N_3614,N_1894);
and U8140 (N_8140,N_3637,N_4744);
and U8141 (N_8141,N_3190,N_4948);
nor U8142 (N_8142,N_4942,N_3545);
and U8143 (N_8143,N_3271,N_4932);
and U8144 (N_8144,N_1701,N_1279);
nand U8145 (N_8145,N_2461,N_4743);
xnor U8146 (N_8146,N_1125,N_1760);
nor U8147 (N_8147,N_3491,N_1488);
nor U8148 (N_8148,N_4254,N_144);
or U8149 (N_8149,N_3413,N_4890);
or U8150 (N_8150,N_1396,N_1639);
and U8151 (N_8151,N_3169,N_4259);
and U8152 (N_8152,N_2580,N_3907);
nand U8153 (N_8153,N_1880,N_2397);
nor U8154 (N_8154,N_3231,N_290);
nand U8155 (N_8155,N_2270,N_2307);
and U8156 (N_8156,N_4601,N_2559);
or U8157 (N_8157,N_492,N_4826);
or U8158 (N_8158,N_276,N_2362);
nand U8159 (N_8159,N_2435,N_4236);
or U8160 (N_8160,N_3387,N_2002);
or U8161 (N_8161,N_3939,N_3273);
nand U8162 (N_8162,N_1608,N_4750);
nor U8163 (N_8163,N_2776,N_4565);
nand U8164 (N_8164,N_320,N_2620);
or U8165 (N_8165,N_1335,N_4946);
nor U8166 (N_8166,N_4233,N_4283);
nor U8167 (N_8167,N_1218,N_11);
and U8168 (N_8168,N_1925,N_2430);
nand U8169 (N_8169,N_169,N_1455);
or U8170 (N_8170,N_3452,N_1167);
nand U8171 (N_8171,N_2822,N_3858);
or U8172 (N_8172,N_1066,N_25);
and U8173 (N_8173,N_4315,N_3542);
and U8174 (N_8174,N_638,N_2972);
nand U8175 (N_8175,N_4820,N_1064);
nor U8176 (N_8176,N_4706,N_332);
nand U8177 (N_8177,N_1488,N_2501);
or U8178 (N_8178,N_1257,N_443);
or U8179 (N_8179,N_1156,N_2232);
nor U8180 (N_8180,N_1442,N_4697);
or U8181 (N_8181,N_10,N_4207);
xnor U8182 (N_8182,N_2273,N_1113);
xnor U8183 (N_8183,N_4623,N_1822);
nand U8184 (N_8184,N_3100,N_3292);
nor U8185 (N_8185,N_3304,N_2135);
and U8186 (N_8186,N_1593,N_1064);
nand U8187 (N_8187,N_2669,N_4507);
or U8188 (N_8188,N_2955,N_2337);
and U8189 (N_8189,N_4096,N_3639);
or U8190 (N_8190,N_2475,N_2471);
or U8191 (N_8191,N_2341,N_2114);
or U8192 (N_8192,N_671,N_4225);
nand U8193 (N_8193,N_832,N_2027);
nand U8194 (N_8194,N_3458,N_1897);
nand U8195 (N_8195,N_1571,N_2556);
or U8196 (N_8196,N_3752,N_358);
nor U8197 (N_8197,N_1061,N_827);
nand U8198 (N_8198,N_3360,N_4371);
and U8199 (N_8199,N_2573,N_4480);
nor U8200 (N_8200,N_1363,N_2970);
xor U8201 (N_8201,N_3103,N_1659);
nand U8202 (N_8202,N_4353,N_1176);
and U8203 (N_8203,N_3863,N_936);
xnor U8204 (N_8204,N_3024,N_4251);
and U8205 (N_8205,N_4241,N_43);
or U8206 (N_8206,N_2942,N_1414);
nor U8207 (N_8207,N_1664,N_88);
nand U8208 (N_8208,N_4197,N_2583);
xor U8209 (N_8209,N_659,N_1251);
and U8210 (N_8210,N_1778,N_3569);
or U8211 (N_8211,N_3684,N_4757);
and U8212 (N_8212,N_4139,N_3063);
nor U8213 (N_8213,N_2183,N_1285);
and U8214 (N_8214,N_4666,N_4762);
and U8215 (N_8215,N_2603,N_740);
or U8216 (N_8216,N_1266,N_4314);
nor U8217 (N_8217,N_3199,N_1731);
or U8218 (N_8218,N_4414,N_522);
or U8219 (N_8219,N_4805,N_2758);
or U8220 (N_8220,N_4287,N_2798);
nor U8221 (N_8221,N_901,N_4223);
and U8222 (N_8222,N_503,N_778);
nand U8223 (N_8223,N_340,N_2319);
or U8224 (N_8224,N_4013,N_2603);
and U8225 (N_8225,N_460,N_4807);
or U8226 (N_8226,N_1726,N_1760);
and U8227 (N_8227,N_2638,N_975);
or U8228 (N_8228,N_604,N_4681);
and U8229 (N_8229,N_2304,N_4107);
nand U8230 (N_8230,N_4,N_1266);
xnor U8231 (N_8231,N_2699,N_3893);
or U8232 (N_8232,N_3786,N_1643);
nand U8233 (N_8233,N_3361,N_2967);
and U8234 (N_8234,N_1595,N_1216);
or U8235 (N_8235,N_871,N_1863);
nand U8236 (N_8236,N_1874,N_4863);
nand U8237 (N_8237,N_3975,N_2034);
nand U8238 (N_8238,N_895,N_87);
nand U8239 (N_8239,N_2847,N_780);
nor U8240 (N_8240,N_3240,N_730);
or U8241 (N_8241,N_4476,N_762);
nor U8242 (N_8242,N_4305,N_2047);
or U8243 (N_8243,N_1354,N_1077);
and U8244 (N_8244,N_4296,N_1901);
and U8245 (N_8245,N_2894,N_3285);
nor U8246 (N_8246,N_2995,N_3624);
and U8247 (N_8247,N_2970,N_3711);
nor U8248 (N_8248,N_3456,N_2371);
xor U8249 (N_8249,N_2441,N_3674);
and U8250 (N_8250,N_1609,N_4547);
nor U8251 (N_8251,N_4371,N_1991);
xor U8252 (N_8252,N_3918,N_1378);
nor U8253 (N_8253,N_2398,N_1441);
and U8254 (N_8254,N_1243,N_1694);
or U8255 (N_8255,N_364,N_4737);
nand U8256 (N_8256,N_2148,N_3285);
nand U8257 (N_8257,N_3815,N_1305);
nand U8258 (N_8258,N_3685,N_2200);
or U8259 (N_8259,N_3960,N_3801);
and U8260 (N_8260,N_299,N_1611);
xor U8261 (N_8261,N_2589,N_3160);
and U8262 (N_8262,N_2684,N_2391);
nand U8263 (N_8263,N_4049,N_3867);
or U8264 (N_8264,N_4050,N_3123);
nor U8265 (N_8265,N_1439,N_1461);
nand U8266 (N_8266,N_2798,N_1374);
nor U8267 (N_8267,N_2688,N_3847);
nor U8268 (N_8268,N_89,N_1080);
nor U8269 (N_8269,N_1777,N_742);
and U8270 (N_8270,N_4240,N_182);
nand U8271 (N_8271,N_2895,N_1573);
nor U8272 (N_8272,N_1268,N_4314);
nand U8273 (N_8273,N_2644,N_2405);
and U8274 (N_8274,N_2619,N_1889);
xor U8275 (N_8275,N_4263,N_4599);
and U8276 (N_8276,N_4531,N_2303);
xnor U8277 (N_8277,N_3503,N_4914);
or U8278 (N_8278,N_3573,N_2041);
and U8279 (N_8279,N_2815,N_81);
nand U8280 (N_8280,N_1748,N_3590);
nor U8281 (N_8281,N_1113,N_4904);
or U8282 (N_8282,N_604,N_1088);
nor U8283 (N_8283,N_1992,N_2741);
and U8284 (N_8284,N_4918,N_1294);
nand U8285 (N_8285,N_2383,N_481);
nor U8286 (N_8286,N_1066,N_3483);
nor U8287 (N_8287,N_3896,N_591);
nor U8288 (N_8288,N_3085,N_3521);
and U8289 (N_8289,N_3812,N_3647);
xor U8290 (N_8290,N_649,N_1480);
and U8291 (N_8291,N_4745,N_3485);
nand U8292 (N_8292,N_4162,N_2652);
nor U8293 (N_8293,N_2063,N_3277);
or U8294 (N_8294,N_2110,N_2080);
or U8295 (N_8295,N_2747,N_113);
nand U8296 (N_8296,N_1329,N_2853);
nand U8297 (N_8297,N_3129,N_1508);
nor U8298 (N_8298,N_3946,N_1491);
and U8299 (N_8299,N_2226,N_2375);
nand U8300 (N_8300,N_2005,N_669);
and U8301 (N_8301,N_3926,N_391);
nand U8302 (N_8302,N_2328,N_2952);
or U8303 (N_8303,N_4080,N_1774);
and U8304 (N_8304,N_681,N_2070);
or U8305 (N_8305,N_522,N_894);
nor U8306 (N_8306,N_336,N_682);
and U8307 (N_8307,N_939,N_666);
nor U8308 (N_8308,N_1828,N_2813);
and U8309 (N_8309,N_2455,N_211);
nand U8310 (N_8310,N_1116,N_3012);
nand U8311 (N_8311,N_3625,N_3446);
or U8312 (N_8312,N_4809,N_444);
xnor U8313 (N_8313,N_1506,N_3360);
nand U8314 (N_8314,N_492,N_1025);
and U8315 (N_8315,N_2361,N_694);
nor U8316 (N_8316,N_4162,N_4827);
xor U8317 (N_8317,N_181,N_3582);
nor U8318 (N_8318,N_3309,N_3796);
or U8319 (N_8319,N_1304,N_592);
xor U8320 (N_8320,N_3394,N_2433);
and U8321 (N_8321,N_3150,N_3147);
nand U8322 (N_8322,N_3676,N_1500);
nor U8323 (N_8323,N_1092,N_2183);
and U8324 (N_8324,N_1393,N_3355);
and U8325 (N_8325,N_3359,N_1741);
or U8326 (N_8326,N_2928,N_4640);
nor U8327 (N_8327,N_3383,N_724);
nor U8328 (N_8328,N_3263,N_496);
and U8329 (N_8329,N_236,N_2644);
and U8330 (N_8330,N_1507,N_3899);
nand U8331 (N_8331,N_4852,N_1114);
and U8332 (N_8332,N_4488,N_1016);
or U8333 (N_8333,N_3129,N_4544);
and U8334 (N_8334,N_4399,N_114);
and U8335 (N_8335,N_4366,N_416);
nor U8336 (N_8336,N_2765,N_111);
nand U8337 (N_8337,N_1820,N_3239);
and U8338 (N_8338,N_4821,N_493);
nor U8339 (N_8339,N_1734,N_2473);
nand U8340 (N_8340,N_3641,N_1235);
xnor U8341 (N_8341,N_1390,N_4828);
or U8342 (N_8342,N_4732,N_2134);
nor U8343 (N_8343,N_3720,N_1192);
nand U8344 (N_8344,N_1709,N_3017);
nor U8345 (N_8345,N_4035,N_2546);
xnor U8346 (N_8346,N_4243,N_3205);
and U8347 (N_8347,N_4221,N_3670);
and U8348 (N_8348,N_824,N_1975);
xor U8349 (N_8349,N_4514,N_1205);
or U8350 (N_8350,N_2247,N_4478);
nor U8351 (N_8351,N_1699,N_739);
nand U8352 (N_8352,N_3733,N_4877);
nand U8353 (N_8353,N_3570,N_3992);
or U8354 (N_8354,N_3198,N_287);
nand U8355 (N_8355,N_4729,N_2937);
and U8356 (N_8356,N_4152,N_1244);
and U8357 (N_8357,N_1875,N_3135);
and U8358 (N_8358,N_2412,N_1036);
nor U8359 (N_8359,N_3179,N_189);
and U8360 (N_8360,N_3194,N_499);
nand U8361 (N_8361,N_4518,N_3951);
and U8362 (N_8362,N_450,N_2018);
nand U8363 (N_8363,N_2650,N_828);
nand U8364 (N_8364,N_4190,N_2557);
nand U8365 (N_8365,N_2942,N_1239);
and U8366 (N_8366,N_1812,N_1250);
nor U8367 (N_8367,N_343,N_4611);
or U8368 (N_8368,N_2156,N_3031);
nor U8369 (N_8369,N_2366,N_4285);
or U8370 (N_8370,N_4127,N_969);
xnor U8371 (N_8371,N_3287,N_261);
nand U8372 (N_8372,N_4887,N_2197);
and U8373 (N_8373,N_121,N_2134);
nand U8374 (N_8374,N_712,N_270);
and U8375 (N_8375,N_2627,N_1021);
xnor U8376 (N_8376,N_1068,N_2517);
and U8377 (N_8377,N_3603,N_3089);
xor U8378 (N_8378,N_1188,N_4027);
or U8379 (N_8379,N_3128,N_1284);
xnor U8380 (N_8380,N_2187,N_786);
xnor U8381 (N_8381,N_3223,N_3744);
or U8382 (N_8382,N_3850,N_866);
or U8383 (N_8383,N_3238,N_2850);
or U8384 (N_8384,N_4955,N_692);
and U8385 (N_8385,N_4436,N_3406);
or U8386 (N_8386,N_757,N_3094);
nand U8387 (N_8387,N_2702,N_1775);
nor U8388 (N_8388,N_320,N_4511);
or U8389 (N_8389,N_4099,N_607);
and U8390 (N_8390,N_614,N_4344);
nor U8391 (N_8391,N_2897,N_170);
or U8392 (N_8392,N_968,N_118);
and U8393 (N_8393,N_827,N_4404);
nand U8394 (N_8394,N_1366,N_1188);
and U8395 (N_8395,N_2491,N_2250);
nand U8396 (N_8396,N_4125,N_2524);
nor U8397 (N_8397,N_2229,N_1014);
xnor U8398 (N_8398,N_1915,N_719);
nor U8399 (N_8399,N_1217,N_743);
or U8400 (N_8400,N_3223,N_1147);
nor U8401 (N_8401,N_768,N_661);
nand U8402 (N_8402,N_859,N_1939);
nand U8403 (N_8403,N_699,N_1452);
and U8404 (N_8404,N_1907,N_1719);
or U8405 (N_8405,N_3076,N_3323);
nor U8406 (N_8406,N_901,N_4548);
or U8407 (N_8407,N_4986,N_3173);
nand U8408 (N_8408,N_4062,N_2316);
xnor U8409 (N_8409,N_4192,N_3325);
xnor U8410 (N_8410,N_4573,N_4890);
nand U8411 (N_8411,N_4781,N_226);
and U8412 (N_8412,N_1697,N_2902);
nand U8413 (N_8413,N_782,N_3007);
and U8414 (N_8414,N_3996,N_1124);
nand U8415 (N_8415,N_4560,N_2523);
xnor U8416 (N_8416,N_1223,N_3381);
nor U8417 (N_8417,N_1665,N_3629);
nor U8418 (N_8418,N_375,N_272);
nand U8419 (N_8419,N_458,N_4030);
and U8420 (N_8420,N_2964,N_414);
or U8421 (N_8421,N_2794,N_1002);
and U8422 (N_8422,N_1017,N_3681);
nand U8423 (N_8423,N_1340,N_4361);
or U8424 (N_8424,N_2869,N_2058);
and U8425 (N_8425,N_4820,N_3612);
xor U8426 (N_8426,N_2025,N_3276);
nand U8427 (N_8427,N_2522,N_207);
nand U8428 (N_8428,N_3937,N_2514);
nor U8429 (N_8429,N_168,N_2697);
and U8430 (N_8430,N_4061,N_3118);
xor U8431 (N_8431,N_1410,N_1285);
nor U8432 (N_8432,N_4496,N_2302);
or U8433 (N_8433,N_4999,N_4165);
nand U8434 (N_8434,N_1977,N_2664);
xnor U8435 (N_8435,N_1453,N_4235);
nor U8436 (N_8436,N_783,N_3777);
or U8437 (N_8437,N_705,N_3878);
and U8438 (N_8438,N_2147,N_2164);
or U8439 (N_8439,N_1683,N_2256);
nor U8440 (N_8440,N_2049,N_4446);
nor U8441 (N_8441,N_3859,N_3735);
nor U8442 (N_8442,N_4303,N_1627);
and U8443 (N_8443,N_2277,N_4017);
or U8444 (N_8444,N_1431,N_3116);
and U8445 (N_8445,N_1100,N_2411);
or U8446 (N_8446,N_213,N_1414);
nor U8447 (N_8447,N_4453,N_3758);
xor U8448 (N_8448,N_3095,N_4302);
nor U8449 (N_8449,N_1304,N_3353);
and U8450 (N_8450,N_325,N_4252);
and U8451 (N_8451,N_2219,N_1262);
nand U8452 (N_8452,N_4976,N_1671);
xnor U8453 (N_8453,N_2132,N_3099);
nand U8454 (N_8454,N_2891,N_3027);
and U8455 (N_8455,N_3104,N_1166);
and U8456 (N_8456,N_886,N_808);
and U8457 (N_8457,N_4905,N_419);
nor U8458 (N_8458,N_1469,N_2711);
xnor U8459 (N_8459,N_2162,N_2246);
nand U8460 (N_8460,N_3186,N_4993);
or U8461 (N_8461,N_2477,N_58);
nand U8462 (N_8462,N_2380,N_3124);
nor U8463 (N_8463,N_3607,N_3463);
nand U8464 (N_8464,N_1785,N_4372);
nand U8465 (N_8465,N_2875,N_4778);
or U8466 (N_8466,N_2287,N_3336);
and U8467 (N_8467,N_99,N_183);
nor U8468 (N_8468,N_2035,N_3200);
xor U8469 (N_8469,N_2119,N_3114);
and U8470 (N_8470,N_3478,N_886);
nor U8471 (N_8471,N_344,N_1053);
or U8472 (N_8472,N_311,N_1968);
nand U8473 (N_8473,N_1984,N_1281);
nor U8474 (N_8474,N_2471,N_1111);
nor U8475 (N_8475,N_3332,N_1448);
xor U8476 (N_8476,N_2185,N_2215);
and U8477 (N_8477,N_4062,N_936);
or U8478 (N_8478,N_1664,N_997);
or U8479 (N_8479,N_584,N_4725);
nand U8480 (N_8480,N_4696,N_4265);
and U8481 (N_8481,N_1062,N_2755);
nor U8482 (N_8482,N_3797,N_1681);
nor U8483 (N_8483,N_1371,N_4736);
and U8484 (N_8484,N_872,N_1176);
nor U8485 (N_8485,N_4156,N_2791);
nand U8486 (N_8486,N_472,N_1188);
or U8487 (N_8487,N_1993,N_843);
nor U8488 (N_8488,N_3302,N_485);
or U8489 (N_8489,N_4554,N_3602);
or U8490 (N_8490,N_726,N_1791);
nor U8491 (N_8491,N_438,N_4953);
nand U8492 (N_8492,N_3764,N_2368);
or U8493 (N_8493,N_1691,N_4868);
and U8494 (N_8494,N_4500,N_3909);
xnor U8495 (N_8495,N_2537,N_2236);
nand U8496 (N_8496,N_1292,N_778);
nor U8497 (N_8497,N_2488,N_669);
xor U8498 (N_8498,N_1725,N_218);
nand U8499 (N_8499,N_149,N_4722);
nand U8500 (N_8500,N_4249,N_1941);
nand U8501 (N_8501,N_1277,N_2547);
nand U8502 (N_8502,N_491,N_3025);
or U8503 (N_8503,N_850,N_269);
and U8504 (N_8504,N_3062,N_1389);
nand U8505 (N_8505,N_848,N_3009);
and U8506 (N_8506,N_1269,N_634);
nand U8507 (N_8507,N_1245,N_2495);
nand U8508 (N_8508,N_4558,N_4918);
and U8509 (N_8509,N_2464,N_3394);
or U8510 (N_8510,N_1106,N_2526);
nor U8511 (N_8511,N_3882,N_4263);
or U8512 (N_8512,N_1216,N_3819);
nand U8513 (N_8513,N_2401,N_3146);
and U8514 (N_8514,N_849,N_710);
nor U8515 (N_8515,N_2727,N_4644);
nor U8516 (N_8516,N_4095,N_2781);
and U8517 (N_8517,N_1985,N_4015);
nor U8518 (N_8518,N_1879,N_4943);
or U8519 (N_8519,N_506,N_4034);
nor U8520 (N_8520,N_3744,N_2813);
nand U8521 (N_8521,N_1146,N_3140);
nand U8522 (N_8522,N_4848,N_1957);
nand U8523 (N_8523,N_4535,N_53);
nor U8524 (N_8524,N_4097,N_1068);
and U8525 (N_8525,N_4808,N_3149);
xor U8526 (N_8526,N_1247,N_4982);
xor U8527 (N_8527,N_1521,N_532);
and U8528 (N_8528,N_4141,N_2758);
nand U8529 (N_8529,N_60,N_578);
nand U8530 (N_8530,N_2403,N_469);
nor U8531 (N_8531,N_320,N_3745);
nor U8532 (N_8532,N_2347,N_154);
nand U8533 (N_8533,N_3388,N_2484);
nor U8534 (N_8534,N_3031,N_3833);
and U8535 (N_8535,N_2942,N_3371);
nand U8536 (N_8536,N_2505,N_1534);
nor U8537 (N_8537,N_2509,N_3442);
nor U8538 (N_8538,N_1974,N_546);
nor U8539 (N_8539,N_2493,N_1550);
nand U8540 (N_8540,N_4407,N_3399);
nor U8541 (N_8541,N_2589,N_3191);
and U8542 (N_8542,N_2535,N_3443);
nor U8543 (N_8543,N_4748,N_3972);
nand U8544 (N_8544,N_3878,N_2901);
nor U8545 (N_8545,N_3483,N_150);
nor U8546 (N_8546,N_4071,N_1566);
and U8547 (N_8547,N_3789,N_4149);
nand U8548 (N_8548,N_3737,N_4509);
nor U8549 (N_8549,N_3469,N_4159);
nor U8550 (N_8550,N_3152,N_1862);
and U8551 (N_8551,N_4793,N_124);
xnor U8552 (N_8552,N_2328,N_4463);
or U8553 (N_8553,N_262,N_3443);
or U8554 (N_8554,N_1263,N_2206);
or U8555 (N_8555,N_2699,N_1420);
nand U8556 (N_8556,N_4906,N_3753);
nand U8557 (N_8557,N_3216,N_2905);
nor U8558 (N_8558,N_1615,N_2477);
and U8559 (N_8559,N_4198,N_2581);
and U8560 (N_8560,N_439,N_4961);
nand U8561 (N_8561,N_2356,N_3198);
and U8562 (N_8562,N_4146,N_748);
or U8563 (N_8563,N_1775,N_1856);
and U8564 (N_8564,N_2006,N_498);
nor U8565 (N_8565,N_2286,N_2394);
or U8566 (N_8566,N_4767,N_3932);
nor U8567 (N_8567,N_862,N_1809);
nor U8568 (N_8568,N_709,N_3232);
and U8569 (N_8569,N_117,N_3676);
and U8570 (N_8570,N_3371,N_1332);
or U8571 (N_8571,N_2521,N_4955);
and U8572 (N_8572,N_412,N_4700);
and U8573 (N_8573,N_132,N_4955);
nand U8574 (N_8574,N_4097,N_3644);
or U8575 (N_8575,N_2578,N_3469);
nand U8576 (N_8576,N_1474,N_2622);
and U8577 (N_8577,N_2449,N_2978);
or U8578 (N_8578,N_1532,N_1334);
nand U8579 (N_8579,N_2365,N_2539);
nor U8580 (N_8580,N_117,N_4706);
xor U8581 (N_8581,N_4866,N_4254);
nand U8582 (N_8582,N_2549,N_1063);
nor U8583 (N_8583,N_139,N_2798);
nand U8584 (N_8584,N_2405,N_4613);
nor U8585 (N_8585,N_3867,N_4529);
or U8586 (N_8586,N_4189,N_420);
and U8587 (N_8587,N_3718,N_3130);
and U8588 (N_8588,N_1750,N_4740);
nor U8589 (N_8589,N_3375,N_4121);
nor U8590 (N_8590,N_2385,N_4775);
xor U8591 (N_8591,N_3257,N_3778);
and U8592 (N_8592,N_2889,N_4629);
xor U8593 (N_8593,N_25,N_3933);
or U8594 (N_8594,N_2832,N_1533);
nand U8595 (N_8595,N_464,N_4734);
nor U8596 (N_8596,N_2141,N_2442);
and U8597 (N_8597,N_434,N_3770);
xnor U8598 (N_8598,N_655,N_2155);
xor U8599 (N_8599,N_4130,N_3302);
nand U8600 (N_8600,N_2592,N_3949);
or U8601 (N_8601,N_4662,N_1839);
nor U8602 (N_8602,N_4591,N_1534);
xor U8603 (N_8603,N_3434,N_1559);
nand U8604 (N_8604,N_4259,N_2831);
and U8605 (N_8605,N_3458,N_2570);
and U8606 (N_8606,N_4330,N_3328);
xor U8607 (N_8607,N_1580,N_4697);
or U8608 (N_8608,N_3585,N_2419);
or U8609 (N_8609,N_3889,N_1660);
nand U8610 (N_8610,N_2609,N_1747);
and U8611 (N_8611,N_2102,N_1622);
nand U8612 (N_8612,N_1814,N_814);
xor U8613 (N_8613,N_2215,N_2961);
or U8614 (N_8614,N_4300,N_1422);
xor U8615 (N_8615,N_3926,N_4644);
or U8616 (N_8616,N_2669,N_4086);
nand U8617 (N_8617,N_3405,N_4161);
xnor U8618 (N_8618,N_1655,N_4092);
nand U8619 (N_8619,N_2085,N_4623);
nor U8620 (N_8620,N_2626,N_3395);
nor U8621 (N_8621,N_825,N_1975);
nand U8622 (N_8622,N_4867,N_4268);
or U8623 (N_8623,N_1593,N_470);
xnor U8624 (N_8624,N_592,N_2379);
nand U8625 (N_8625,N_2084,N_1356);
nor U8626 (N_8626,N_908,N_3844);
nor U8627 (N_8627,N_720,N_4654);
nand U8628 (N_8628,N_3760,N_382);
nor U8629 (N_8629,N_1441,N_2911);
nor U8630 (N_8630,N_1216,N_3990);
nand U8631 (N_8631,N_1016,N_3956);
and U8632 (N_8632,N_1547,N_2757);
and U8633 (N_8633,N_1906,N_3284);
or U8634 (N_8634,N_1052,N_1326);
nand U8635 (N_8635,N_3874,N_546);
nand U8636 (N_8636,N_3464,N_2960);
nand U8637 (N_8637,N_3657,N_4407);
or U8638 (N_8638,N_2837,N_987);
or U8639 (N_8639,N_4606,N_660);
xor U8640 (N_8640,N_1168,N_4321);
and U8641 (N_8641,N_1366,N_4652);
and U8642 (N_8642,N_4506,N_4640);
nor U8643 (N_8643,N_3878,N_2184);
or U8644 (N_8644,N_3140,N_416);
or U8645 (N_8645,N_3075,N_511);
or U8646 (N_8646,N_1883,N_2202);
or U8647 (N_8647,N_4101,N_274);
and U8648 (N_8648,N_1299,N_2566);
xor U8649 (N_8649,N_1055,N_2688);
or U8650 (N_8650,N_751,N_2530);
nand U8651 (N_8651,N_4057,N_587);
or U8652 (N_8652,N_2611,N_205);
and U8653 (N_8653,N_2365,N_3734);
nand U8654 (N_8654,N_4432,N_856);
nand U8655 (N_8655,N_959,N_3460);
nand U8656 (N_8656,N_1558,N_3810);
nor U8657 (N_8657,N_4460,N_2817);
nor U8658 (N_8658,N_4005,N_520);
or U8659 (N_8659,N_4466,N_1839);
nand U8660 (N_8660,N_2026,N_1271);
and U8661 (N_8661,N_2509,N_2826);
nor U8662 (N_8662,N_4460,N_4117);
nand U8663 (N_8663,N_1058,N_4917);
and U8664 (N_8664,N_276,N_2344);
nand U8665 (N_8665,N_3448,N_2862);
nor U8666 (N_8666,N_2103,N_1968);
and U8667 (N_8667,N_3737,N_2243);
nand U8668 (N_8668,N_4921,N_3333);
xor U8669 (N_8669,N_4636,N_1971);
nor U8670 (N_8670,N_2863,N_2342);
or U8671 (N_8671,N_331,N_379);
or U8672 (N_8672,N_772,N_4132);
xor U8673 (N_8673,N_3746,N_895);
or U8674 (N_8674,N_4584,N_2577);
or U8675 (N_8675,N_4952,N_304);
and U8676 (N_8676,N_1436,N_3677);
nor U8677 (N_8677,N_4610,N_2182);
nor U8678 (N_8678,N_262,N_2968);
nand U8679 (N_8679,N_3675,N_4714);
nand U8680 (N_8680,N_1823,N_1919);
nor U8681 (N_8681,N_3023,N_692);
and U8682 (N_8682,N_4403,N_2907);
nand U8683 (N_8683,N_1643,N_884);
nor U8684 (N_8684,N_4665,N_4297);
xnor U8685 (N_8685,N_1640,N_1770);
nand U8686 (N_8686,N_2822,N_4638);
xnor U8687 (N_8687,N_33,N_1662);
xnor U8688 (N_8688,N_2382,N_2697);
nand U8689 (N_8689,N_700,N_210);
nand U8690 (N_8690,N_4097,N_1486);
and U8691 (N_8691,N_4322,N_2066);
nor U8692 (N_8692,N_3235,N_3499);
and U8693 (N_8693,N_985,N_2284);
xor U8694 (N_8694,N_1837,N_1209);
and U8695 (N_8695,N_1611,N_1009);
or U8696 (N_8696,N_1016,N_4205);
or U8697 (N_8697,N_4008,N_1188);
and U8698 (N_8698,N_4633,N_2679);
or U8699 (N_8699,N_2193,N_4629);
nor U8700 (N_8700,N_4983,N_1547);
and U8701 (N_8701,N_347,N_3528);
and U8702 (N_8702,N_4457,N_46);
or U8703 (N_8703,N_2835,N_4842);
nor U8704 (N_8704,N_2280,N_2744);
xnor U8705 (N_8705,N_4087,N_12);
and U8706 (N_8706,N_3326,N_552);
nand U8707 (N_8707,N_4485,N_925);
or U8708 (N_8708,N_1760,N_2643);
nor U8709 (N_8709,N_4786,N_2015);
nand U8710 (N_8710,N_3834,N_825);
nor U8711 (N_8711,N_210,N_3558);
nor U8712 (N_8712,N_709,N_4247);
nor U8713 (N_8713,N_4912,N_851);
or U8714 (N_8714,N_2614,N_422);
and U8715 (N_8715,N_4129,N_3967);
or U8716 (N_8716,N_1399,N_4950);
nand U8717 (N_8717,N_1705,N_491);
xnor U8718 (N_8718,N_4649,N_4911);
and U8719 (N_8719,N_3810,N_4213);
or U8720 (N_8720,N_3829,N_1543);
nand U8721 (N_8721,N_4723,N_1107);
or U8722 (N_8722,N_3116,N_3947);
nand U8723 (N_8723,N_1225,N_3936);
nand U8724 (N_8724,N_456,N_1249);
or U8725 (N_8725,N_6,N_2491);
nand U8726 (N_8726,N_4833,N_3033);
or U8727 (N_8727,N_3071,N_1598);
and U8728 (N_8728,N_4503,N_648);
nand U8729 (N_8729,N_1918,N_330);
and U8730 (N_8730,N_3485,N_4790);
nand U8731 (N_8731,N_2592,N_469);
xnor U8732 (N_8732,N_2487,N_4363);
nand U8733 (N_8733,N_923,N_749);
nand U8734 (N_8734,N_2653,N_3453);
nor U8735 (N_8735,N_3196,N_1754);
nor U8736 (N_8736,N_2770,N_4894);
nor U8737 (N_8737,N_4637,N_2380);
xnor U8738 (N_8738,N_632,N_218);
xnor U8739 (N_8739,N_1954,N_4885);
and U8740 (N_8740,N_4078,N_4507);
xor U8741 (N_8741,N_3750,N_3882);
nand U8742 (N_8742,N_4706,N_3254);
or U8743 (N_8743,N_4902,N_307);
nor U8744 (N_8744,N_3796,N_3863);
or U8745 (N_8745,N_3093,N_1137);
nand U8746 (N_8746,N_3494,N_381);
or U8747 (N_8747,N_4096,N_3854);
nor U8748 (N_8748,N_875,N_3387);
and U8749 (N_8749,N_325,N_1960);
and U8750 (N_8750,N_823,N_2768);
and U8751 (N_8751,N_1003,N_3876);
or U8752 (N_8752,N_3756,N_1476);
nand U8753 (N_8753,N_661,N_152);
nor U8754 (N_8754,N_4518,N_1793);
nor U8755 (N_8755,N_107,N_3935);
or U8756 (N_8756,N_924,N_3523);
nor U8757 (N_8757,N_3886,N_3746);
nand U8758 (N_8758,N_2342,N_2090);
nand U8759 (N_8759,N_330,N_452);
xnor U8760 (N_8760,N_4105,N_4141);
nor U8761 (N_8761,N_4823,N_1725);
and U8762 (N_8762,N_4946,N_928);
and U8763 (N_8763,N_4011,N_4349);
nand U8764 (N_8764,N_4076,N_572);
nor U8765 (N_8765,N_2789,N_3490);
and U8766 (N_8766,N_1214,N_2182);
nor U8767 (N_8767,N_4355,N_709);
nor U8768 (N_8768,N_382,N_2627);
nand U8769 (N_8769,N_3412,N_3084);
nand U8770 (N_8770,N_1681,N_2188);
nor U8771 (N_8771,N_1473,N_4965);
and U8772 (N_8772,N_3543,N_98);
and U8773 (N_8773,N_3252,N_3110);
and U8774 (N_8774,N_1509,N_2895);
nand U8775 (N_8775,N_3293,N_2391);
nor U8776 (N_8776,N_4528,N_760);
or U8777 (N_8777,N_1325,N_1485);
or U8778 (N_8778,N_3509,N_638);
and U8779 (N_8779,N_1730,N_460);
nand U8780 (N_8780,N_623,N_3195);
and U8781 (N_8781,N_1867,N_2642);
nand U8782 (N_8782,N_2170,N_4216);
nor U8783 (N_8783,N_1822,N_3511);
nand U8784 (N_8784,N_3179,N_214);
or U8785 (N_8785,N_4747,N_4491);
nor U8786 (N_8786,N_1627,N_3963);
or U8787 (N_8787,N_2672,N_4193);
nand U8788 (N_8788,N_3412,N_981);
nor U8789 (N_8789,N_31,N_4339);
and U8790 (N_8790,N_4410,N_1867);
nand U8791 (N_8791,N_2812,N_4267);
or U8792 (N_8792,N_1411,N_3698);
or U8793 (N_8793,N_3897,N_989);
nor U8794 (N_8794,N_1857,N_4638);
nor U8795 (N_8795,N_1412,N_1069);
nand U8796 (N_8796,N_1852,N_2121);
and U8797 (N_8797,N_2536,N_1469);
and U8798 (N_8798,N_2389,N_4556);
nor U8799 (N_8799,N_4834,N_269);
and U8800 (N_8800,N_1229,N_2320);
nand U8801 (N_8801,N_4553,N_3275);
and U8802 (N_8802,N_4179,N_1953);
nor U8803 (N_8803,N_1432,N_29);
nand U8804 (N_8804,N_2862,N_3842);
nor U8805 (N_8805,N_2844,N_38);
or U8806 (N_8806,N_4123,N_4804);
and U8807 (N_8807,N_4652,N_3383);
nor U8808 (N_8808,N_3924,N_4110);
nor U8809 (N_8809,N_3951,N_400);
or U8810 (N_8810,N_4074,N_2248);
nand U8811 (N_8811,N_584,N_4935);
and U8812 (N_8812,N_3450,N_4450);
nand U8813 (N_8813,N_953,N_4868);
and U8814 (N_8814,N_4343,N_682);
or U8815 (N_8815,N_118,N_4038);
or U8816 (N_8816,N_2342,N_4946);
xnor U8817 (N_8817,N_1642,N_2391);
nand U8818 (N_8818,N_4775,N_2139);
nand U8819 (N_8819,N_3796,N_4600);
or U8820 (N_8820,N_1507,N_845);
nor U8821 (N_8821,N_215,N_202);
or U8822 (N_8822,N_591,N_1251);
and U8823 (N_8823,N_3407,N_3939);
and U8824 (N_8824,N_2764,N_907);
nor U8825 (N_8825,N_1386,N_3947);
and U8826 (N_8826,N_1989,N_4990);
and U8827 (N_8827,N_1795,N_1787);
and U8828 (N_8828,N_3594,N_1510);
nor U8829 (N_8829,N_1499,N_3426);
nand U8830 (N_8830,N_3295,N_1827);
or U8831 (N_8831,N_4828,N_2488);
nand U8832 (N_8832,N_2878,N_4800);
or U8833 (N_8833,N_4550,N_3211);
or U8834 (N_8834,N_4242,N_4047);
or U8835 (N_8835,N_3233,N_4802);
or U8836 (N_8836,N_4766,N_2212);
and U8837 (N_8837,N_4124,N_2226);
and U8838 (N_8838,N_3005,N_1324);
or U8839 (N_8839,N_1998,N_960);
nand U8840 (N_8840,N_3286,N_4646);
or U8841 (N_8841,N_4282,N_2039);
nand U8842 (N_8842,N_946,N_4292);
or U8843 (N_8843,N_2656,N_4140);
or U8844 (N_8844,N_3363,N_1747);
nand U8845 (N_8845,N_1154,N_418);
and U8846 (N_8846,N_3788,N_880);
nand U8847 (N_8847,N_3840,N_2240);
nor U8848 (N_8848,N_3021,N_2348);
and U8849 (N_8849,N_908,N_4501);
nand U8850 (N_8850,N_2558,N_2317);
xnor U8851 (N_8851,N_1780,N_1410);
or U8852 (N_8852,N_4100,N_2230);
or U8853 (N_8853,N_355,N_864);
nor U8854 (N_8854,N_4570,N_384);
or U8855 (N_8855,N_2920,N_1572);
nor U8856 (N_8856,N_766,N_61);
nand U8857 (N_8857,N_4100,N_2774);
and U8858 (N_8858,N_3940,N_3240);
nand U8859 (N_8859,N_4757,N_314);
and U8860 (N_8860,N_1738,N_106);
or U8861 (N_8861,N_1664,N_2129);
and U8862 (N_8862,N_1260,N_4531);
and U8863 (N_8863,N_3881,N_3502);
nor U8864 (N_8864,N_381,N_4737);
and U8865 (N_8865,N_2881,N_3097);
xnor U8866 (N_8866,N_4873,N_4930);
nand U8867 (N_8867,N_3269,N_4712);
xnor U8868 (N_8868,N_647,N_1695);
nand U8869 (N_8869,N_3655,N_3890);
xor U8870 (N_8870,N_4582,N_4614);
xnor U8871 (N_8871,N_1655,N_2115);
and U8872 (N_8872,N_1217,N_3419);
nor U8873 (N_8873,N_539,N_1927);
nor U8874 (N_8874,N_1770,N_641);
or U8875 (N_8875,N_422,N_4345);
and U8876 (N_8876,N_4425,N_3680);
or U8877 (N_8877,N_825,N_1168);
nand U8878 (N_8878,N_776,N_2829);
nor U8879 (N_8879,N_1039,N_3922);
nand U8880 (N_8880,N_4014,N_4483);
nand U8881 (N_8881,N_713,N_3813);
and U8882 (N_8882,N_4389,N_3167);
xnor U8883 (N_8883,N_62,N_3183);
nor U8884 (N_8884,N_3866,N_1820);
nor U8885 (N_8885,N_3239,N_4795);
xor U8886 (N_8886,N_810,N_1641);
or U8887 (N_8887,N_1289,N_4135);
nor U8888 (N_8888,N_3389,N_4327);
nand U8889 (N_8889,N_4527,N_4744);
xnor U8890 (N_8890,N_4613,N_3613);
xor U8891 (N_8891,N_3707,N_4007);
xor U8892 (N_8892,N_1181,N_898);
and U8893 (N_8893,N_434,N_195);
nand U8894 (N_8894,N_4010,N_60);
and U8895 (N_8895,N_370,N_528);
nand U8896 (N_8896,N_4719,N_3383);
nand U8897 (N_8897,N_3699,N_2104);
nand U8898 (N_8898,N_521,N_4794);
and U8899 (N_8899,N_2658,N_3989);
or U8900 (N_8900,N_1619,N_643);
nand U8901 (N_8901,N_3670,N_3885);
or U8902 (N_8902,N_3996,N_2243);
and U8903 (N_8903,N_1455,N_4592);
or U8904 (N_8904,N_538,N_3890);
or U8905 (N_8905,N_371,N_274);
nor U8906 (N_8906,N_1255,N_2322);
and U8907 (N_8907,N_983,N_2836);
or U8908 (N_8908,N_1254,N_4392);
nand U8909 (N_8909,N_2959,N_1800);
or U8910 (N_8910,N_2977,N_1150);
and U8911 (N_8911,N_1877,N_1241);
nand U8912 (N_8912,N_1789,N_4738);
nand U8913 (N_8913,N_827,N_2126);
nand U8914 (N_8914,N_745,N_1756);
nand U8915 (N_8915,N_3822,N_3221);
and U8916 (N_8916,N_3485,N_1361);
or U8917 (N_8917,N_2399,N_3435);
or U8918 (N_8918,N_3858,N_875);
and U8919 (N_8919,N_4245,N_2690);
and U8920 (N_8920,N_42,N_660);
nor U8921 (N_8921,N_3880,N_4230);
and U8922 (N_8922,N_2112,N_434);
nand U8923 (N_8923,N_876,N_455);
xnor U8924 (N_8924,N_2860,N_856);
or U8925 (N_8925,N_3880,N_734);
or U8926 (N_8926,N_1107,N_700);
nor U8927 (N_8927,N_699,N_4263);
and U8928 (N_8928,N_2444,N_3945);
or U8929 (N_8929,N_1932,N_4999);
and U8930 (N_8930,N_4331,N_1181);
xor U8931 (N_8931,N_744,N_4158);
xor U8932 (N_8932,N_3097,N_429);
or U8933 (N_8933,N_189,N_3045);
nand U8934 (N_8934,N_1728,N_3401);
xor U8935 (N_8935,N_805,N_4142);
nand U8936 (N_8936,N_1151,N_2817);
nand U8937 (N_8937,N_3398,N_3358);
and U8938 (N_8938,N_2972,N_36);
and U8939 (N_8939,N_548,N_3902);
or U8940 (N_8940,N_2698,N_308);
xor U8941 (N_8941,N_181,N_2349);
nand U8942 (N_8942,N_4381,N_1662);
and U8943 (N_8943,N_4494,N_1031);
and U8944 (N_8944,N_4910,N_1922);
xor U8945 (N_8945,N_969,N_4755);
nor U8946 (N_8946,N_4606,N_881);
xnor U8947 (N_8947,N_2191,N_1581);
or U8948 (N_8948,N_1839,N_3776);
nand U8949 (N_8949,N_4910,N_3894);
nand U8950 (N_8950,N_4868,N_1308);
nand U8951 (N_8951,N_1224,N_170);
and U8952 (N_8952,N_4442,N_1268);
and U8953 (N_8953,N_888,N_262);
nand U8954 (N_8954,N_3553,N_3478);
and U8955 (N_8955,N_4541,N_1506);
and U8956 (N_8956,N_4304,N_4268);
and U8957 (N_8957,N_1014,N_2971);
xor U8958 (N_8958,N_4649,N_204);
or U8959 (N_8959,N_1684,N_2044);
nor U8960 (N_8960,N_1259,N_4204);
or U8961 (N_8961,N_3241,N_1474);
nor U8962 (N_8962,N_2704,N_3958);
and U8963 (N_8963,N_4960,N_4197);
xor U8964 (N_8964,N_1572,N_137);
or U8965 (N_8965,N_3667,N_2084);
nor U8966 (N_8966,N_3383,N_682);
and U8967 (N_8967,N_1277,N_2267);
nor U8968 (N_8968,N_1344,N_3583);
or U8969 (N_8969,N_3016,N_2096);
and U8970 (N_8970,N_2101,N_414);
nor U8971 (N_8971,N_4009,N_922);
or U8972 (N_8972,N_4138,N_4137);
nand U8973 (N_8973,N_4139,N_380);
nand U8974 (N_8974,N_3194,N_2844);
nand U8975 (N_8975,N_3157,N_4146);
nand U8976 (N_8976,N_4010,N_3976);
nor U8977 (N_8977,N_3563,N_3849);
nand U8978 (N_8978,N_983,N_1583);
nand U8979 (N_8979,N_1967,N_507);
nor U8980 (N_8980,N_3180,N_4028);
or U8981 (N_8981,N_4077,N_3983);
and U8982 (N_8982,N_610,N_3444);
or U8983 (N_8983,N_490,N_4538);
or U8984 (N_8984,N_4268,N_720);
or U8985 (N_8985,N_1222,N_2587);
and U8986 (N_8986,N_1799,N_4283);
and U8987 (N_8987,N_1341,N_2360);
or U8988 (N_8988,N_1094,N_4120);
nor U8989 (N_8989,N_1316,N_2922);
and U8990 (N_8990,N_2436,N_1253);
nand U8991 (N_8991,N_4248,N_4640);
nand U8992 (N_8992,N_3794,N_874);
or U8993 (N_8993,N_1093,N_376);
or U8994 (N_8994,N_4552,N_1052);
nor U8995 (N_8995,N_224,N_2774);
and U8996 (N_8996,N_26,N_4664);
or U8997 (N_8997,N_956,N_2296);
nand U8998 (N_8998,N_3069,N_3487);
xor U8999 (N_8999,N_359,N_1640);
nand U9000 (N_9000,N_1415,N_1571);
xor U9001 (N_9001,N_1741,N_2158);
xor U9002 (N_9002,N_4966,N_1284);
or U9003 (N_9003,N_2833,N_1238);
and U9004 (N_9004,N_534,N_2817);
and U9005 (N_9005,N_2831,N_2593);
nor U9006 (N_9006,N_2992,N_229);
nor U9007 (N_9007,N_3762,N_4048);
or U9008 (N_9008,N_4544,N_2648);
nand U9009 (N_9009,N_2970,N_3180);
or U9010 (N_9010,N_4621,N_2128);
nor U9011 (N_9011,N_2778,N_4052);
or U9012 (N_9012,N_1598,N_2757);
nand U9013 (N_9013,N_4693,N_191);
and U9014 (N_9014,N_129,N_1571);
nor U9015 (N_9015,N_2799,N_3985);
nand U9016 (N_9016,N_2512,N_1366);
nand U9017 (N_9017,N_873,N_3723);
nor U9018 (N_9018,N_2251,N_2016);
nand U9019 (N_9019,N_4797,N_160);
nand U9020 (N_9020,N_792,N_3260);
nand U9021 (N_9021,N_4579,N_4126);
and U9022 (N_9022,N_2838,N_4792);
or U9023 (N_9023,N_2854,N_2054);
and U9024 (N_9024,N_2698,N_2290);
or U9025 (N_9025,N_2199,N_3361);
or U9026 (N_9026,N_1896,N_3568);
nand U9027 (N_9027,N_573,N_4717);
nand U9028 (N_9028,N_2746,N_3842);
nand U9029 (N_9029,N_343,N_515);
and U9030 (N_9030,N_3610,N_37);
nor U9031 (N_9031,N_4081,N_1516);
and U9032 (N_9032,N_7,N_510);
and U9033 (N_9033,N_2041,N_619);
xor U9034 (N_9034,N_1043,N_1518);
nor U9035 (N_9035,N_3797,N_3593);
nand U9036 (N_9036,N_3664,N_144);
nand U9037 (N_9037,N_4492,N_1353);
or U9038 (N_9038,N_4804,N_1004);
nor U9039 (N_9039,N_4375,N_2070);
or U9040 (N_9040,N_19,N_768);
nor U9041 (N_9041,N_4517,N_1931);
and U9042 (N_9042,N_2352,N_789);
and U9043 (N_9043,N_3470,N_4133);
or U9044 (N_9044,N_1357,N_1730);
xor U9045 (N_9045,N_1014,N_4077);
nor U9046 (N_9046,N_4319,N_2497);
nor U9047 (N_9047,N_164,N_828);
nor U9048 (N_9048,N_2896,N_4949);
and U9049 (N_9049,N_1828,N_4701);
nand U9050 (N_9050,N_1438,N_2117);
or U9051 (N_9051,N_722,N_2108);
and U9052 (N_9052,N_2811,N_2739);
xor U9053 (N_9053,N_4875,N_1572);
nor U9054 (N_9054,N_4502,N_3355);
nor U9055 (N_9055,N_125,N_2729);
nand U9056 (N_9056,N_1535,N_1595);
xnor U9057 (N_9057,N_684,N_2894);
nor U9058 (N_9058,N_2763,N_2404);
and U9059 (N_9059,N_1470,N_2468);
nand U9060 (N_9060,N_2549,N_3529);
and U9061 (N_9061,N_3920,N_3367);
nor U9062 (N_9062,N_1041,N_3290);
nand U9063 (N_9063,N_1285,N_3266);
and U9064 (N_9064,N_3861,N_2161);
and U9065 (N_9065,N_2861,N_3985);
and U9066 (N_9066,N_1492,N_4167);
nor U9067 (N_9067,N_1961,N_1991);
and U9068 (N_9068,N_1317,N_409);
nand U9069 (N_9069,N_4688,N_3840);
nand U9070 (N_9070,N_4613,N_3596);
or U9071 (N_9071,N_3003,N_4021);
nand U9072 (N_9072,N_3600,N_4510);
and U9073 (N_9073,N_1590,N_58);
xnor U9074 (N_9074,N_2513,N_3268);
nand U9075 (N_9075,N_4982,N_1570);
and U9076 (N_9076,N_4639,N_1851);
xnor U9077 (N_9077,N_498,N_3857);
or U9078 (N_9078,N_3185,N_3062);
or U9079 (N_9079,N_2616,N_3184);
or U9080 (N_9080,N_3601,N_431);
nor U9081 (N_9081,N_414,N_353);
nor U9082 (N_9082,N_1791,N_4607);
and U9083 (N_9083,N_3669,N_1055);
or U9084 (N_9084,N_4239,N_2837);
and U9085 (N_9085,N_3130,N_3532);
and U9086 (N_9086,N_3000,N_475);
nor U9087 (N_9087,N_3546,N_2442);
and U9088 (N_9088,N_3515,N_2891);
and U9089 (N_9089,N_1341,N_2762);
nand U9090 (N_9090,N_4019,N_4004);
nand U9091 (N_9091,N_21,N_1127);
nand U9092 (N_9092,N_3592,N_1398);
nand U9093 (N_9093,N_1575,N_3877);
or U9094 (N_9094,N_1556,N_3243);
nor U9095 (N_9095,N_2262,N_385);
xnor U9096 (N_9096,N_3546,N_2114);
nand U9097 (N_9097,N_2563,N_4826);
and U9098 (N_9098,N_373,N_1941);
nor U9099 (N_9099,N_1563,N_4142);
nand U9100 (N_9100,N_3441,N_2459);
nor U9101 (N_9101,N_114,N_3810);
nand U9102 (N_9102,N_2237,N_2056);
xnor U9103 (N_9103,N_4198,N_4102);
nand U9104 (N_9104,N_501,N_303);
nor U9105 (N_9105,N_2963,N_1330);
nand U9106 (N_9106,N_4962,N_4614);
or U9107 (N_9107,N_1585,N_2367);
and U9108 (N_9108,N_4842,N_4135);
and U9109 (N_9109,N_2923,N_4840);
and U9110 (N_9110,N_2725,N_4318);
and U9111 (N_9111,N_2533,N_4586);
and U9112 (N_9112,N_4016,N_3917);
and U9113 (N_9113,N_563,N_3326);
or U9114 (N_9114,N_1500,N_2880);
and U9115 (N_9115,N_4151,N_910);
nand U9116 (N_9116,N_1183,N_1054);
nand U9117 (N_9117,N_3591,N_1665);
or U9118 (N_9118,N_4677,N_2447);
nor U9119 (N_9119,N_3940,N_1119);
and U9120 (N_9120,N_628,N_903);
nand U9121 (N_9121,N_4680,N_3282);
or U9122 (N_9122,N_2964,N_3260);
nand U9123 (N_9123,N_2258,N_409);
nor U9124 (N_9124,N_3217,N_4545);
or U9125 (N_9125,N_1242,N_889);
or U9126 (N_9126,N_1076,N_2190);
nand U9127 (N_9127,N_4646,N_4691);
nand U9128 (N_9128,N_4080,N_713);
nor U9129 (N_9129,N_1370,N_1059);
nor U9130 (N_9130,N_4812,N_1690);
or U9131 (N_9131,N_3809,N_2232);
nand U9132 (N_9132,N_1501,N_3324);
nand U9133 (N_9133,N_2889,N_3732);
and U9134 (N_9134,N_1825,N_2958);
nand U9135 (N_9135,N_1178,N_836);
and U9136 (N_9136,N_3999,N_2748);
nand U9137 (N_9137,N_4005,N_4138);
nor U9138 (N_9138,N_3276,N_1998);
and U9139 (N_9139,N_1084,N_1687);
xor U9140 (N_9140,N_4501,N_629);
and U9141 (N_9141,N_4528,N_263);
and U9142 (N_9142,N_1887,N_335);
and U9143 (N_9143,N_543,N_312);
nor U9144 (N_9144,N_2196,N_1825);
nor U9145 (N_9145,N_2054,N_2967);
nand U9146 (N_9146,N_3151,N_4834);
and U9147 (N_9147,N_1047,N_675);
or U9148 (N_9148,N_260,N_1301);
nor U9149 (N_9149,N_1556,N_3936);
and U9150 (N_9150,N_1394,N_1056);
and U9151 (N_9151,N_819,N_917);
nor U9152 (N_9152,N_4365,N_3386);
nand U9153 (N_9153,N_4239,N_4544);
nor U9154 (N_9154,N_4675,N_2337);
nor U9155 (N_9155,N_357,N_4976);
or U9156 (N_9156,N_643,N_3055);
nand U9157 (N_9157,N_3826,N_207);
xnor U9158 (N_9158,N_1733,N_3219);
nand U9159 (N_9159,N_1325,N_3745);
xor U9160 (N_9160,N_1144,N_1602);
or U9161 (N_9161,N_1117,N_4768);
and U9162 (N_9162,N_3747,N_1798);
or U9163 (N_9163,N_4561,N_4632);
nor U9164 (N_9164,N_2200,N_4836);
nand U9165 (N_9165,N_775,N_860);
nor U9166 (N_9166,N_4078,N_3377);
and U9167 (N_9167,N_783,N_2708);
xnor U9168 (N_9168,N_2365,N_1645);
or U9169 (N_9169,N_3709,N_2536);
nor U9170 (N_9170,N_4493,N_3643);
nand U9171 (N_9171,N_2512,N_3634);
or U9172 (N_9172,N_2082,N_223);
and U9173 (N_9173,N_366,N_2942);
xor U9174 (N_9174,N_747,N_4349);
xor U9175 (N_9175,N_102,N_3603);
or U9176 (N_9176,N_330,N_876);
or U9177 (N_9177,N_3188,N_110);
nor U9178 (N_9178,N_213,N_3313);
and U9179 (N_9179,N_3693,N_129);
nor U9180 (N_9180,N_4695,N_141);
or U9181 (N_9181,N_1373,N_2274);
or U9182 (N_9182,N_3547,N_2511);
nor U9183 (N_9183,N_4634,N_3621);
and U9184 (N_9184,N_4622,N_1765);
or U9185 (N_9185,N_4431,N_3462);
xnor U9186 (N_9186,N_4574,N_800);
nor U9187 (N_9187,N_1412,N_4490);
nor U9188 (N_9188,N_2298,N_644);
and U9189 (N_9189,N_663,N_4987);
or U9190 (N_9190,N_4460,N_1401);
xor U9191 (N_9191,N_663,N_2732);
nor U9192 (N_9192,N_2277,N_2457);
nor U9193 (N_9193,N_1563,N_2808);
nor U9194 (N_9194,N_302,N_4404);
nand U9195 (N_9195,N_4684,N_4500);
nand U9196 (N_9196,N_1458,N_46);
and U9197 (N_9197,N_275,N_1946);
or U9198 (N_9198,N_3806,N_209);
nor U9199 (N_9199,N_3243,N_235);
nand U9200 (N_9200,N_3217,N_1427);
nor U9201 (N_9201,N_2064,N_3858);
and U9202 (N_9202,N_2014,N_3047);
nor U9203 (N_9203,N_3134,N_2830);
nor U9204 (N_9204,N_3632,N_1688);
nand U9205 (N_9205,N_4834,N_1956);
or U9206 (N_9206,N_3453,N_3988);
nand U9207 (N_9207,N_494,N_2859);
nand U9208 (N_9208,N_4316,N_1701);
nand U9209 (N_9209,N_1341,N_808);
nand U9210 (N_9210,N_3935,N_3536);
or U9211 (N_9211,N_107,N_1376);
nor U9212 (N_9212,N_3549,N_3191);
or U9213 (N_9213,N_2051,N_1589);
nor U9214 (N_9214,N_14,N_4546);
nand U9215 (N_9215,N_2692,N_889);
nand U9216 (N_9216,N_324,N_350);
or U9217 (N_9217,N_590,N_4678);
nor U9218 (N_9218,N_4827,N_3894);
and U9219 (N_9219,N_315,N_1699);
or U9220 (N_9220,N_1461,N_4258);
and U9221 (N_9221,N_2096,N_1379);
and U9222 (N_9222,N_4785,N_3371);
nor U9223 (N_9223,N_4535,N_695);
nor U9224 (N_9224,N_2916,N_294);
nor U9225 (N_9225,N_2806,N_2566);
and U9226 (N_9226,N_4516,N_3559);
or U9227 (N_9227,N_1494,N_390);
and U9228 (N_9228,N_2957,N_4870);
and U9229 (N_9229,N_1933,N_4323);
or U9230 (N_9230,N_2837,N_474);
xnor U9231 (N_9231,N_2774,N_3147);
nand U9232 (N_9232,N_1836,N_3165);
or U9233 (N_9233,N_2797,N_1692);
or U9234 (N_9234,N_4704,N_163);
and U9235 (N_9235,N_4915,N_3223);
and U9236 (N_9236,N_1207,N_2052);
and U9237 (N_9237,N_2006,N_2079);
nor U9238 (N_9238,N_2617,N_3556);
nor U9239 (N_9239,N_4864,N_2281);
or U9240 (N_9240,N_1505,N_139);
or U9241 (N_9241,N_4267,N_4262);
or U9242 (N_9242,N_1775,N_2243);
or U9243 (N_9243,N_3129,N_1554);
nor U9244 (N_9244,N_3687,N_2419);
nor U9245 (N_9245,N_3661,N_878);
and U9246 (N_9246,N_4430,N_3288);
or U9247 (N_9247,N_2244,N_1530);
xnor U9248 (N_9248,N_2597,N_2986);
and U9249 (N_9249,N_3329,N_2645);
nor U9250 (N_9250,N_2044,N_324);
and U9251 (N_9251,N_1146,N_3059);
or U9252 (N_9252,N_3111,N_1275);
xor U9253 (N_9253,N_4243,N_4901);
or U9254 (N_9254,N_355,N_1151);
and U9255 (N_9255,N_4225,N_4831);
or U9256 (N_9256,N_2003,N_2936);
and U9257 (N_9257,N_4108,N_1217);
nand U9258 (N_9258,N_515,N_1246);
nor U9259 (N_9259,N_3385,N_3280);
and U9260 (N_9260,N_1166,N_2014);
nor U9261 (N_9261,N_4166,N_3180);
or U9262 (N_9262,N_3683,N_3922);
xnor U9263 (N_9263,N_4174,N_4942);
nand U9264 (N_9264,N_431,N_4062);
and U9265 (N_9265,N_4319,N_434);
or U9266 (N_9266,N_4853,N_133);
nand U9267 (N_9267,N_4177,N_2956);
nand U9268 (N_9268,N_92,N_2497);
nand U9269 (N_9269,N_2961,N_3297);
nor U9270 (N_9270,N_4101,N_253);
xnor U9271 (N_9271,N_2685,N_3752);
and U9272 (N_9272,N_3192,N_4276);
nand U9273 (N_9273,N_1538,N_3863);
and U9274 (N_9274,N_224,N_959);
nand U9275 (N_9275,N_2663,N_1404);
nand U9276 (N_9276,N_4533,N_3954);
xor U9277 (N_9277,N_4654,N_493);
and U9278 (N_9278,N_4468,N_392);
and U9279 (N_9279,N_4769,N_3177);
nand U9280 (N_9280,N_2052,N_3663);
nor U9281 (N_9281,N_3510,N_795);
or U9282 (N_9282,N_1520,N_2094);
or U9283 (N_9283,N_990,N_1121);
or U9284 (N_9284,N_2891,N_2362);
nand U9285 (N_9285,N_2302,N_3815);
nand U9286 (N_9286,N_2831,N_721);
or U9287 (N_9287,N_594,N_4296);
nand U9288 (N_9288,N_3688,N_4265);
and U9289 (N_9289,N_3142,N_3584);
or U9290 (N_9290,N_4412,N_1446);
or U9291 (N_9291,N_3690,N_4063);
or U9292 (N_9292,N_63,N_3078);
nand U9293 (N_9293,N_1303,N_4005);
and U9294 (N_9294,N_1319,N_3514);
nor U9295 (N_9295,N_3436,N_4475);
and U9296 (N_9296,N_3279,N_4802);
nand U9297 (N_9297,N_4937,N_835);
and U9298 (N_9298,N_4004,N_3774);
nor U9299 (N_9299,N_3323,N_1662);
nor U9300 (N_9300,N_522,N_4624);
or U9301 (N_9301,N_2305,N_4944);
or U9302 (N_9302,N_2403,N_2114);
nand U9303 (N_9303,N_4275,N_2049);
nand U9304 (N_9304,N_254,N_708);
nor U9305 (N_9305,N_4319,N_2977);
and U9306 (N_9306,N_87,N_1692);
nor U9307 (N_9307,N_531,N_2714);
or U9308 (N_9308,N_4480,N_2031);
and U9309 (N_9309,N_478,N_4818);
nor U9310 (N_9310,N_4561,N_2058);
or U9311 (N_9311,N_2593,N_4422);
and U9312 (N_9312,N_2980,N_3870);
or U9313 (N_9313,N_3032,N_3655);
and U9314 (N_9314,N_2332,N_2032);
and U9315 (N_9315,N_955,N_3340);
nand U9316 (N_9316,N_2093,N_1180);
and U9317 (N_9317,N_3016,N_312);
and U9318 (N_9318,N_2895,N_4350);
nand U9319 (N_9319,N_1420,N_4249);
and U9320 (N_9320,N_3548,N_502);
nand U9321 (N_9321,N_1719,N_3366);
nand U9322 (N_9322,N_2206,N_3504);
nand U9323 (N_9323,N_3878,N_3467);
nand U9324 (N_9324,N_1912,N_870);
nand U9325 (N_9325,N_2095,N_1176);
nand U9326 (N_9326,N_1047,N_1937);
or U9327 (N_9327,N_3256,N_4206);
or U9328 (N_9328,N_3195,N_3847);
nor U9329 (N_9329,N_2549,N_4580);
nor U9330 (N_9330,N_2815,N_2965);
nor U9331 (N_9331,N_1521,N_1538);
nor U9332 (N_9332,N_1376,N_289);
or U9333 (N_9333,N_3658,N_3097);
and U9334 (N_9334,N_3637,N_1130);
and U9335 (N_9335,N_2380,N_76);
and U9336 (N_9336,N_3994,N_3873);
and U9337 (N_9337,N_1513,N_4562);
or U9338 (N_9338,N_1007,N_3384);
and U9339 (N_9339,N_3965,N_241);
nor U9340 (N_9340,N_2362,N_3473);
and U9341 (N_9341,N_1593,N_4540);
or U9342 (N_9342,N_4819,N_550);
nand U9343 (N_9343,N_3112,N_1917);
nand U9344 (N_9344,N_1612,N_1851);
nor U9345 (N_9345,N_1390,N_3777);
or U9346 (N_9346,N_2075,N_3164);
and U9347 (N_9347,N_3912,N_2093);
and U9348 (N_9348,N_2610,N_2935);
and U9349 (N_9349,N_2800,N_2310);
or U9350 (N_9350,N_1269,N_3052);
nand U9351 (N_9351,N_3834,N_3238);
nand U9352 (N_9352,N_4994,N_328);
nand U9353 (N_9353,N_3900,N_1667);
or U9354 (N_9354,N_3398,N_804);
and U9355 (N_9355,N_1045,N_3969);
or U9356 (N_9356,N_4088,N_337);
nand U9357 (N_9357,N_432,N_1469);
and U9358 (N_9358,N_1347,N_2019);
nor U9359 (N_9359,N_4224,N_1886);
nor U9360 (N_9360,N_4279,N_1978);
and U9361 (N_9361,N_659,N_1485);
nor U9362 (N_9362,N_3954,N_3495);
or U9363 (N_9363,N_650,N_3255);
and U9364 (N_9364,N_2561,N_4644);
nor U9365 (N_9365,N_3735,N_312);
or U9366 (N_9366,N_1440,N_3672);
nor U9367 (N_9367,N_3187,N_242);
nand U9368 (N_9368,N_4135,N_1199);
nand U9369 (N_9369,N_3826,N_4008);
nor U9370 (N_9370,N_515,N_1063);
or U9371 (N_9371,N_3596,N_21);
nand U9372 (N_9372,N_463,N_4577);
nor U9373 (N_9373,N_3324,N_1784);
nand U9374 (N_9374,N_918,N_3898);
and U9375 (N_9375,N_4659,N_2772);
nand U9376 (N_9376,N_4502,N_4305);
and U9377 (N_9377,N_3161,N_665);
and U9378 (N_9378,N_2484,N_2751);
nand U9379 (N_9379,N_3332,N_2868);
nor U9380 (N_9380,N_2897,N_2966);
and U9381 (N_9381,N_3864,N_1960);
nand U9382 (N_9382,N_154,N_1054);
nor U9383 (N_9383,N_3482,N_1562);
nor U9384 (N_9384,N_111,N_1860);
nor U9385 (N_9385,N_3551,N_3514);
or U9386 (N_9386,N_2252,N_4017);
and U9387 (N_9387,N_3922,N_751);
nor U9388 (N_9388,N_4444,N_1225);
nand U9389 (N_9389,N_209,N_1741);
xnor U9390 (N_9390,N_504,N_3479);
xnor U9391 (N_9391,N_482,N_4034);
or U9392 (N_9392,N_4767,N_2892);
or U9393 (N_9393,N_1492,N_1694);
nor U9394 (N_9394,N_823,N_4241);
and U9395 (N_9395,N_1272,N_4722);
and U9396 (N_9396,N_2264,N_733);
nand U9397 (N_9397,N_1497,N_1669);
or U9398 (N_9398,N_1749,N_2570);
nor U9399 (N_9399,N_4199,N_4700);
and U9400 (N_9400,N_2939,N_4977);
nand U9401 (N_9401,N_146,N_4693);
nor U9402 (N_9402,N_3139,N_117);
nand U9403 (N_9403,N_3064,N_1136);
nand U9404 (N_9404,N_1963,N_46);
nand U9405 (N_9405,N_4721,N_951);
nor U9406 (N_9406,N_1429,N_3105);
nor U9407 (N_9407,N_3736,N_1959);
xnor U9408 (N_9408,N_1975,N_861);
and U9409 (N_9409,N_1613,N_4805);
nand U9410 (N_9410,N_1247,N_2463);
or U9411 (N_9411,N_2523,N_2049);
and U9412 (N_9412,N_4239,N_1088);
nand U9413 (N_9413,N_556,N_1669);
xnor U9414 (N_9414,N_106,N_1670);
and U9415 (N_9415,N_4788,N_2911);
and U9416 (N_9416,N_1534,N_1214);
nor U9417 (N_9417,N_3514,N_3147);
nor U9418 (N_9418,N_806,N_2422);
or U9419 (N_9419,N_2745,N_4177);
xnor U9420 (N_9420,N_536,N_2934);
xor U9421 (N_9421,N_4452,N_790);
nor U9422 (N_9422,N_3507,N_4713);
nor U9423 (N_9423,N_2854,N_1870);
and U9424 (N_9424,N_393,N_3526);
or U9425 (N_9425,N_835,N_452);
or U9426 (N_9426,N_1813,N_2656);
xnor U9427 (N_9427,N_4679,N_1668);
or U9428 (N_9428,N_4235,N_411);
or U9429 (N_9429,N_4568,N_2524);
or U9430 (N_9430,N_1390,N_2837);
xnor U9431 (N_9431,N_3144,N_4455);
nand U9432 (N_9432,N_3802,N_1698);
nand U9433 (N_9433,N_3643,N_4658);
nor U9434 (N_9434,N_3396,N_2995);
nand U9435 (N_9435,N_930,N_4880);
nor U9436 (N_9436,N_1713,N_2940);
xor U9437 (N_9437,N_2466,N_1137);
and U9438 (N_9438,N_8,N_4025);
nor U9439 (N_9439,N_4999,N_4684);
and U9440 (N_9440,N_3156,N_847);
and U9441 (N_9441,N_4686,N_2005);
nand U9442 (N_9442,N_898,N_4476);
or U9443 (N_9443,N_3297,N_709);
and U9444 (N_9444,N_371,N_1624);
nor U9445 (N_9445,N_3066,N_3953);
nor U9446 (N_9446,N_712,N_530);
xnor U9447 (N_9447,N_77,N_553);
nor U9448 (N_9448,N_664,N_4182);
and U9449 (N_9449,N_152,N_389);
nand U9450 (N_9450,N_747,N_1827);
and U9451 (N_9451,N_2362,N_4414);
and U9452 (N_9452,N_1995,N_277);
nand U9453 (N_9453,N_466,N_1623);
or U9454 (N_9454,N_3997,N_2417);
and U9455 (N_9455,N_2312,N_1846);
nor U9456 (N_9456,N_3829,N_1475);
or U9457 (N_9457,N_4367,N_450);
nand U9458 (N_9458,N_3722,N_4869);
nor U9459 (N_9459,N_3283,N_3900);
xnor U9460 (N_9460,N_467,N_671);
and U9461 (N_9461,N_4484,N_4702);
or U9462 (N_9462,N_4946,N_306);
and U9463 (N_9463,N_4703,N_406);
and U9464 (N_9464,N_1677,N_576);
and U9465 (N_9465,N_4340,N_1393);
nor U9466 (N_9466,N_2783,N_1739);
nor U9467 (N_9467,N_3801,N_863);
nor U9468 (N_9468,N_2840,N_3538);
nand U9469 (N_9469,N_2478,N_615);
or U9470 (N_9470,N_593,N_2006);
and U9471 (N_9471,N_4248,N_1023);
nand U9472 (N_9472,N_3271,N_4810);
or U9473 (N_9473,N_1336,N_1891);
or U9474 (N_9474,N_187,N_1918);
nor U9475 (N_9475,N_4335,N_4956);
and U9476 (N_9476,N_745,N_2156);
and U9477 (N_9477,N_4295,N_4736);
nand U9478 (N_9478,N_1226,N_4269);
nor U9479 (N_9479,N_2728,N_1971);
and U9480 (N_9480,N_1288,N_2619);
nor U9481 (N_9481,N_3842,N_2330);
xnor U9482 (N_9482,N_3809,N_4845);
and U9483 (N_9483,N_4926,N_1809);
xor U9484 (N_9484,N_1438,N_1900);
or U9485 (N_9485,N_2626,N_802);
nor U9486 (N_9486,N_1532,N_3951);
xnor U9487 (N_9487,N_811,N_2645);
xor U9488 (N_9488,N_2357,N_2638);
nor U9489 (N_9489,N_1272,N_1430);
nand U9490 (N_9490,N_4201,N_2397);
or U9491 (N_9491,N_2344,N_3911);
nor U9492 (N_9492,N_2692,N_4317);
nand U9493 (N_9493,N_3334,N_1100);
or U9494 (N_9494,N_4743,N_4230);
and U9495 (N_9495,N_3946,N_350);
nor U9496 (N_9496,N_726,N_689);
nand U9497 (N_9497,N_4936,N_4180);
or U9498 (N_9498,N_757,N_1099);
or U9499 (N_9499,N_3048,N_1656);
nor U9500 (N_9500,N_4563,N_1029);
nor U9501 (N_9501,N_614,N_228);
nor U9502 (N_9502,N_1340,N_2969);
or U9503 (N_9503,N_2724,N_2744);
nor U9504 (N_9504,N_242,N_1392);
and U9505 (N_9505,N_2921,N_3449);
nor U9506 (N_9506,N_880,N_20);
nor U9507 (N_9507,N_4561,N_4995);
or U9508 (N_9508,N_2609,N_309);
nor U9509 (N_9509,N_4604,N_571);
and U9510 (N_9510,N_1914,N_313);
nor U9511 (N_9511,N_839,N_4978);
or U9512 (N_9512,N_1698,N_2746);
or U9513 (N_9513,N_78,N_2305);
or U9514 (N_9514,N_4674,N_1872);
and U9515 (N_9515,N_2295,N_2026);
nor U9516 (N_9516,N_2420,N_1903);
nor U9517 (N_9517,N_2450,N_371);
and U9518 (N_9518,N_492,N_4949);
nand U9519 (N_9519,N_2941,N_3499);
or U9520 (N_9520,N_2860,N_2845);
nor U9521 (N_9521,N_4928,N_4734);
and U9522 (N_9522,N_1264,N_4818);
or U9523 (N_9523,N_3319,N_2428);
nand U9524 (N_9524,N_3493,N_565);
nor U9525 (N_9525,N_275,N_1981);
or U9526 (N_9526,N_4278,N_3946);
or U9527 (N_9527,N_1270,N_2417);
and U9528 (N_9528,N_134,N_4885);
nand U9529 (N_9529,N_139,N_2123);
or U9530 (N_9530,N_2806,N_1034);
or U9531 (N_9531,N_4448,N_1005);
nand U9532 (N_9532,N_116,N_3111);
and U9533 (N_9533,N_1025,N_2988);
nor U9534 (N_9534,N_2410,N_4879);
nor U9535 (N_9535,N_493,N_183);
nand U9536 (N_9536,N_990,N_4357);
xnor U9537 (N_9537,N_4828,N_3898);
nand U9538 (N_9538,N_2085,N_4073);
nor U9539 (N_9539,N_962,N_2579);
nand U9540 (N_9540,N_317,N_3120);
nand U9541 (N_9541,N_615,N_207);
nand U9542 (N_9542,N_2091,N_1843);
and U9543 (N_9543,N_3192,N_1424);
nor U9544 (N_9544,N_3505,N_3561);
nand U9545 (N_9545,N_3133,N_451);
xor U9546 (N_9546,N_466,N_3526);
nor U9547 (N_9547,N_4420,N_1006);
nor U9548 (N_9548,N_3013,N_4350);
and U9549 (N_9549,N_365,N_453);
or U9550 (N_9550,N_1627,N_4424);
or U9551 (N_9551,N_606,N_1187);
nand U9552 (N_9552,N_1958,N_3605);
nor U9553 (N_9553,N_2815,N_364);
nand U9554 (N_9554,N_134,N_3415);
nor U9555 (N_9555,N_2918,N_1082);
and U9556 (N_9556,N_3074,N_4614);
nor U9557 (N_9557,N_1770,N_3621);
and U9558 (N_9558,N_3899,N_4619);
and U9559 (N_9559,N_1160,N_1858);
xnor U9560 (N_9560,N_503,N_1582);
nand U9561 (N_9561,N_3243,N_3316);
and U9562 (N_9562,N_952,N_4544);
nand U9563 (N_9563,N_1250,N_844);
nand U9564 (N_9564,N_3209,N_4046);
nand U9565 (N_9565,N_4236,N_1549);
or U9566 (N_9566,N_1490,N_1956);
nand U9567 (N_9567,N_1127,N_1493);
or U9568 (N_9568,N_3255,N_3615);
and U9569 (N_9569,N_546,N_4710);
xnor U9570 (N_9570,N_2903,N_441);
nor U9571 (N_9571,N_1357,N_1441);
nand U9572 (N_9572,N_2394,N_181);
and U9573 (N_9573,N_170,N_2493);
or U9574 (N_9574,N_1019,N_3657);
nor U9575 (N_9575,N_1804,N_3433);
xor U9576 (N_9576,N_3144,N_2275);
or U9577 (N_9577,N_1273,N_3173);
or U9578 (N_9578,N_4098,N_4795);
nor U9579 (N_9579,N_3756,N_2969);
nand U9580 (N_9580,N_3822,N_3568);
or U9581 (N_9581,N_3801,N_2733);
nor U9582 (N_9582,N_263,N_1133);
or U9583 (N_9583,N_1423,N_4547);
and U9584 (N_9584,N_696,N_249);
nand U9585 (N_9585,N_3334,N_371);
nor U9586 (N_9586,N_4367,N_4613);
or U9587 (N_9587,N_965,N_978);
or U9588 (N_9588,N_3940,N_2023);
and U9589 (N_9589,N_3100,N_3533);
nand U9590 (N_9590,N_4074,N_2747);
xor U9591 (N_9591,N_1384,N_2690);
nand U9592 (N_9592,N_4913,N_4969);
or U9593 (N_9593,N_2429,N_848);
and U9594 (N_9594,N_3673,N_1399);
nand U9595 (N_9595,N_2290,N_3019);
and U9596 (N_9596,N_699,N_3042);
nor U9597 (N_9597,N_3564,N_1888);
nand U9598 (N_9598,N_3048,N_1846);
nand U9599 (N_9599,N_3952,N_2953);
and U9600 (N_9600,N_931,N_472);
or U9601 (N_9601,N_677,N_4053);
and U9602 (N_9602,N_3095,N_1652);
nand U9603 (N_9603,N_2990,N_4565);
nand U9604 (N_9604,N_844,N_770);
nor U9605 (N_9605,N_4643,N_130);
nor U9606 (N_9606,N_4529,N_1230);
or U9607 (N_9607,N_3468,N_2926);
or U9608 (N_9608,N_2516,N_2975);
nand U9609 (N_9609,N_4744,N_97);
nand U9610 (N_9610,N_1293,N_3833);
or U9611 (N_9611,N_2029,N_3613);
nor U9612 (N_9612,N_1580,N_2996);
nor U9613 (N_9613,N_2458,N_2167);
or U9614 (N_9614,N_243,N_3127);
and U9615 (N_9615,N_3905,N_1813);
nand U9616 (N_9616,N_4325,N_1201);
nand U9617 (N_9617,N_2934,N_1718);
and U9618 (N_9618,N_642,N_1531);
nor U9619 (N_9619,N_4528,N_4243);
nand U9620 (N_9620,N_799,N_2231);
nor U9621 (N_9621,N_253,N_3886);
or U9622 (N_9622,N_4401,N_3578);
or U9623 (N_9623,N_4538,N_3848);
xor U9624 (N_9624,N_3877,N_4973);
nand U9625 (N_9625,N_4205,N_3373);
or U9626 (N_9626,N_3004,N_3483);
xor U9627 (N_9627,N_3442,N_121);
nor U9628 (N_9628,N_4409,N_323);
nor U9629 (N_9629,N_710,N_2715);
nor U9630 (N_9630,N_1876,N_2012);
and U9631 (N_9631,N_4338,N_2653);
nand U9632 (N_9632,N_1460,N_2023);
nand U9633 (N_9633,N_1278,N_991);
and U9634 (N_9634,N_773,N_1877);
or U9635 (N_9635,N_38,N_1345);
nand U9636 (N_9636,N_2665,N_4954);
nand U9637 (N_9637,N_4536,N_2393);
nor U9638 (N_9638,N_2064,N_4620);
xor U9639 (N_9639,N_19,N_4371);
or U9640 (N_9640,N_4951,N_1831);
and U9641 (N_9641,N_421,N_2376);
nand U9642 (N_9642,N_426,N_1072);
nand U9643 (N_9643,N_2603,N_11);
nor U9644 (N_9644,N_3551,N_1702);
or U9645 (N_9645,N_687,N_253);
or U9646 (N_9646,N_2157,N_4607);
and U9647 (N_9647,N_3000,N_3675);
and U9648 (N_9648,N_3910,N_4752);
or U9649 (N_9649,N_3249,N_132);
nand U9650 (N_9650,N_3723,N_4506);
or U9651 (N_9651,N_4334,N_3075);
nand U9652 (N_9652,N_3254,N_4692);
or U9653 (N_9653,N_2492,N_3485);
and U9654 (N_9654,N_3132,N_4069);
and U9655 (N_9655,N_3937,N_4212);
nor U9656 (N_9656,N_2418,N_4072);
nor U9657 (N_9657,N_4611,N_516);
and U9658 (N_9658,N_4555,N_4819);
nand U9659 (N_9659,N_4588,N_4056);
nand U9660 (N_9660,N_1597,N_3590);
nor U9661 (N_9661,N_155,N_761);
nor U9662 (N_9662,N_2322,N_552);
nand U9663 (N_9663,N_2072,N_2945);
nand U9664 (N_9664,N_2142,N_424);
nand U9665 (N_9665,N_3510,N_2653);
nand U9666 (N_9666,N_3386,N_646);
and U9667 (N_9667,N_2384,N_2135);
and U9668 (N_9668,N_2587,N_2728);
nor U9669 (N_9669,N_2570,N_2916);
or U9670 (N_9670,N_560,N_1223);
xor U9671 (N_9671,N_3162,N_3189);
xnor U9672 (N_9672,N_866,N_2726);
nand U9673 (N_9673,N_2535,N_4568);
and U9674 (N_9674,N_3924,N_3042);
or U9675 (N_9675,N_4344,N_3324);
nor U9676 (N_9676,N_182,N_3173);
and U9677 (N_9677,N_807,N_2621);
nand U9678 (N_9678,N_3611,N_3373);
and U9679 (N_9679,N_3663,N_661);
nand U9680 (N_9680,N_499,N_59);
and U9681 (N_9681,N_4304,N_2296);
nor U9682 (N_9682,N_1649,N_72);
xor U9683 (N_9683,N_2988,N_3872);
nand U9684 (N_9684,N_2906,N_3931);
nand U9685 (N_9685,N_4486,N_2692);
xnor U9686 (N_9686,N_116,N_3820);
and U9687 (N_9687,N_4336,N_792);
and U9688 (N_9688,N_628,N_1951);
nand U9689 (N_9689,N_3262,N_4807);
and U9690 (N_9690,N_2073,N_4994);
nand U9691 (N_9691,N_3206,N_421);
and U9692 (N_9692,N_100,N_1096);
or U9693 (N_9693,N_1122,N_4072);
nand U9694 (N_9694,N_3719,N_3417);
and U9695 (N_9695,N_2738,N_1232);
or U9696 (N_9696,N_574,N_1958);
nand U9697 (N_9697,N_775,N_4403);
and U9698 (N_9698,N_2138,N_2679);
and U9699 (N_9699,N_920,N_117);
nor U9700 (N_9700,N_1492,N_3950);
or U9701 (N_9701,N_3409,N_3139);
nand U9702 (N_9702,N_3708,N_508);
or U9703 (N_9703,N_4159,N_7);
and U9704 (N_9704,N_461,N_1442);
and U9705 (N_9705,N_4423,N_1102);
nand U9706 (N_9706,N_2514,N_1268);
and U9707 (N_9707,N_2283,N_1308);
or U9708 (N_9708,N_2473,N_4344);
or U9709 (N_9709,N_4979,N_476);
and U9710 (N_9710,N_2323,N_1012);
and U9711 (N_9711,N_2686,N_4702);
nor U9712 (N_9712,N_1523,N_194);
nand U9713 (N_9713,N_3400,N_2899);
or U9714 (N_9714,N_33,N_2377);
nor U9715 (N_9715,N_4209,N_4350);
nor U9716 (N_9716,N_3751,N_4469);
nor U9717 (N_9717,N_3729,N_2157);
nand U9718 (N_9718,N_3423,N_3572);
and U9719 (N_9719,N_288,N_3433);
nor U9720 (N_9720,N_3703,N_1317);
or U9721 (N_9721,N_4923,N_4112);
nor U9722 (N_9722,N_3377,N_1702);
nor U9723 (N_9723,N_2704,N_741);
nor U9724 (N_9724,N_1504,N_3300);
xnor U9725 (N_9725,N_32,N_3299);
or U9726 (N_9726,N_1259,N_4044);
or U9727 (N_9727,N_2736,N_521);
nor U9728 (N_9728,N_2013,N_420);
and U9729 (N_9729,N_1381,N_4504);
and U9730 (N_9730,N_1454,N_695);
nor U9731 (N_9731,N_2075,N_2374);
nand U9732 (N_9732,N_3258,N_1480);
nand U9733 (N_9733,N_2270,N_1730);
and U9734 (N_9734,N_2794,N_3625);
nand U9735 (N_9735,N_3620,N_2819);
nor U9736 (N_9736,N_676,N_4808);
xor U9737 (N_9737,N_381,N_4817);
or U9738 (N_9738,N_2784,N_2872);
xor U9739 (N_9739,N_3782,N_1796);
nor U9740 (N_9740,N_1775,N_2910);
nor U9741 (N_9741,N_985,N_4507);
xnor U9742 (N_9742,N_189,N_840);
nor U9743 (N_9743,N_315,N_1306);
nor U9744 (N_9744,N_4842,N_3550);
and U9745 (N_9745,N_221,N_919);
nand U9746 (N_9746,N_1979,N_4640);
or U9747 (N_9747,N_3297,N_1362);
xnor U9748 (N_9748,N_2617,N_639);
nor U9749 (N_9749,N_2206,N_3739);
or U9750 (N_9750,N_3871,N_4698);
or U9751 (N_9751,N_3176,N_3029);
or U9752 (N_9752,N_214,N_3198);
nor U9753 (N_9753,N_4320,N_2977);
nor U9754 (N_9754,N_3570,N_4757);
or U9755 (N_9755,N_2557,N_3660);
nand U9756 (N_9756,N_3014,N_1720);
nor U9757 (N_9757,N_3991,N_3533);
nand U9758 (N_9758,N_2778,N_884);
and U9759 (N_9759,N_4097,N_79);
xnor U9760 (N_9760,N_3142,N_3916);
nor U9761 (N_9761,N_3325,N_862);
or U9762 (N_9762,N_1881,N_3925);
or U9763 (N_9763,N_4287,N_1629);
nor U9764 (N_9764,N_4190,N_886);
and U9765 (N_9765,N_4919,N_1281);
or U9766 (N_9766,N_4925,N_3514);
nor U9767 (N_9767,N_4282,N_2236);
or U9768 (N_9768,N_4164,N_1729);
nor U9769 (N_9769,N_3826,N_1589);
nand U9770 (N_9770,N_1064,N_3369);
nor U9771 (N_9771,N_1749,N_3130);
nand U9772 (N_9772,N_2095,N_4884);
and U9773 (N_9773,N_1304,N_4559);
nand U9774 (N_9774,N_1740,N_4007);
nand U9775 (N_9775,N_1026,N_2332);
and U9776 (N_9776,N_4978,N_3077);
or U9777 (N_9777,N_827,N_919);
and U9778 (N_9778,N_3740,N_1233);
or U9779 (N_9779,N_800,N_501);
nor U9780 (N_9780,N_4703,N_1362);
or U9781 (N_9781,N_4724,N_3366);
xnor U9782 (N_9782,N_1243,N_4177);
nor U9783 (N_9783,N_937,N_2343);
nand U9784 (N_9784,N_4328,N_3784);
and U9785 (N_9785,N_888,N_1368);
nor U9786 (N_9786,N_643,N_3475);
nand U9787 (N_9787,N_3988,N_4744);
nand U9788 (N_9788,N_558,N_1582);
and U9789 (N_9789,N_3823,N_3680);
or U9790 (N_9790,N_2255,N_2490);
nor U9791 (N_9791,N_4397,N_3136);
and U9792 (N_9792,N_3082,N_3375);
or U9793 (N_9793,N_4160,N_4193);
or U9794 (N_9794,N_4840,N_3965);
nor U9795 (N_9795,N_4816,N_1433);
nor U9796 (N_9796,N_391,N_201);
nand U9797 (N_9797,N_3161,N_3072);
and U9798 (N_9798,N_752,N_2241);
nor U9799 (N_9799,N_1224,N_3203);
and U9800 (N_9800,N_2216,N_1421);
and U9801 (N_9801,N_2261,N_1438);
and U9802 (N_9802,N_3317,N_703);
nand U9803 (N_9803,N_531,N_3289);
nor U9804 (N_9804,N_3840,N_4965);
nor U9805 (N_9805,N_1355,N_748);
and U9806 (N_9806,N_2823,N_2977);
xor U9807 (N_9807,N_2689,N_844);
nor U9808 (N_9808,N_1579,N_3099);
nor U9809 (N_9809,N_1873,N_4183);
nor U9810 (N_9810,N_481,N_302);
and U9811 (N_9811,N_3909,N_4553);
and U9812 (N_9812,N_1596,N_346);
or U9813 (N_9813,N_3181,N_4578);
and U9814 (N_9814,N_1812,N_2219);
and U9815 (N_9815,N_1029,N_2137);
or U9816 (N_9816,N_355,N_441);
xor U9817 (N_9817,N_1580,N_540);
nand U9818 (N_9818,N_77,N_3365);
xor U9819 (N_9819,N_773,N_836);
nor U9820 (N_9820,N_761,N_239);
and U9821 (N_9821,N_2523,N_3373);
and U9822 (N_9822,N_3405,N_1361);
and U9823 (N_9823,N_2164,N_2969);
nor U9824 (N_9824,N_1753,N_2649);
xnor U9825 (N_9825,N_3044,N_2236);
nand U9826 (N_9826,N_4889,N_168);
and U9827 (N_9827,N_2733,N_4867);
xor U9828 (N_9828,N_1423,N_3486);
nor U9829 (N_9829,N_2849,N_3507);
xor U9830 (N_9830,N_3179,N_2482);
and U9831 (N_9831,N_2291,N_3473);
or U9832 (N_9832,N_32,N_3671);
xnor U9833 (N_9833,N_3228,N_3816);
and U9834 (N_9834,N_3302,N_1194);
and U9835 (N_9835,N_3305,N_2783);
xor U9836 (N_9836,N_4063,N_415);
or U9837 (N_9837,N_1562,N_4324);
xnor U9838 (N_9838,N_4509,N_544);
nor U9839 (N_9839,N_1083,N_2943);
nand U9840 (N_9840,N_4597,N_2257);
and U9841 (N_9841,N_1191,N_1533);
nor U9842 (N_9842,N_4169,N_882);
and U9843 (N_9843,N_3194,N_3022);
or U9844 (N_9844,N_1370,N_3608);
and U9845 (N_9845,N_1902,N_3337);
and U9846 (N_9846,N_2750,N_1079);
nand U9847 (N_9847,N_3971,N_2590);
nor U9848 (N_9848,N_1942,N_860);
nor U9849 (N_9849,N_2328,N_978);
nand U9850 (N_9850,N_2035,N_857);
nor U9851 (N_9851,N_3415,N_4969);
nor U9852 (N_9852,N_1942,N_1604);
nand U9853 (N_9853,N_2423,N_3828);
and U9854 (N_9854,N_2251,N_4065);
nand U9855 (N_9855,N_834,N_3641);
nor U9856 (N_9856,N_2198,N_680);
or U9857 (N_9857,N_4867,N_4649);
nor U9858 (N_9858,N_3161,N_4016);
nand U9859 (N_9859,N_1672,N_4095);
or U9860 (N_9860,N_1038,N_4304);
or U9861 (N_9861,N_488,N_1774);
nor U9862 (N_9862,N_109,N_826);
nand U9863 (N_9863,N_2447,N_3169);
or U9864 (N_9864,N_1553,N_3885);
nand U9865 (N_9865,N_2404,N_4473);
and U9866 (N_9866,N_3103,N_4451);
nand U9867 (N_9867,N_2645,N_927);
or U9868 (N_9868,N_2327,N_2320);
or U9869 (N_9869,N_499,N_2021);
or U9870 (N_9870,N_1046,N_1011);
nand U9871 (N_9871,N_2585,N_4205);
nand U9872 (N_9872,N_3181,N_2013);
and U9873 (N_9873,N_3351,N_2699);
and U9874 (N_9874,N_1467,N_136);
or U9875 (N_9875,N_3169,N_3634);
or U9876 (N_9876,N_815,N_3987);
nor U9877 (N_9877,N_4325,N_611);
or U9878 (N_9878,N_88,N_2914);
and U9879 (N_9879,N_621,N_728);
or U9880 (N_9880,N_2553,N_4833);
and U9881 (N_9881,N_2007,N_702);
nand U9882 (N_9882,N_742,N_373);
and U9883 (N_9883,N_3620,N_80);
or U9884 (N_9884,N_1362,N_1072);
nor U9885 (N_9885,N_852,N_1872);
nand U9886 (N_9886,N_712,N_4143);
and U9887 (N_9887,N_1537,N_61);
nor U9888 (N_9888,N_4224,N_99);
or U9889 (N_9889,N_1344,N_3553);
nor U9890 (N_9890,N_969,N_1992);
or U9891 (N_9891,N_841,N_4072);
or U9892 (N_9892,N_2741,N_1762);
and U9893 (N_9893,N_581,N_895);
nand U9894 (N_9894,N_3514,N_328);
nor U9895 (N_9895,N_2120,N_3600);
nand U9896 (N_9896,N_3842,N_3449);
nand U9897 (N_9897,N_4828,N_2150);
xnor U9898 (N_9898,N_440,N_3505);
nand U9899 (N_9899,N_4406,N_3349);
nor U9900 (N_9900,N_661,N_2130);
or U9901 (N_9901,N_1903,N_1466);
or U9902 (N_9902,N_2813,N_3796);
nor U9903 (N_9903,N_3919,N_3498);
nand U9904 (N_9904,N_1674,N_178);
xor U9905 (N_9905,N_4855,N_2671);
and U9906 (N_9906,N_2534,N_3043);
nor U9907 (N_9907,N_1547,N_315);
xor U9908 (N_9908,N_1602,N_1476);
or U9909 (N_9909,N_904,N_2842);
nor U9910 (N_9910,N_4428,N_481);
nor U9911 (N_9911,N_4540,N_2114);
or U9912 (N_9912,N_3397,N_2152);
nor U9913 (N_9913,N_4055,N_4398);
nand U9914 (N_9914,N_813,N_1255);
and U9915 (N_9915,N_12,N_4887);
and U9916 (N_9916,N_1139,N_1216);
nor U9917 (N_9917,N_62,N_838);
or U9918 (N_9918,N_2286,N_2705);
nand U9919 (N_9919,N_4245,N_3253);
or U9920 (N_9920,N_4918,N_1818);
xnor U9921 (N_9921,N_1236,N_3098);
and U9922 (N_9922,N_1647,N_1586);
nor U9923 (N_9923,N_373,N_1957);
nor U9924 (N_9924,N_446,N_2817);
or U9925 (N_9925,N_3972,N_882);
or U9926 (N_9926,N_1360,N_4438);
xor U9927 (N_9927,N_1933,N_99);
or U9928 (N_9928,N_2480,N_1256);
or U9929 (N_9929,N_2510,N_4945);
or U9930 (N_9930,N_1526,N_201);
nand U9931 (N_9931,N_4863,N_3586);
nor U9932 (N_9932,N_3701,N_4064);
nand U9933 (N_9933,N_4996,N_1174);
xnor U9934 (N_9934,N_1249,N_3630);
or U9935 (N_9935,N_1559,N_1258);
and U9936 (N_9936,N_2028,N_1286);
nand U9937 (N_9937,N_199,N_2661);
nand U9938 (N_9938,N_4821,N_3412);
nor U9939 (N_9939,N_1329,N_241);
or U9940 (N_9940,N_3141,N_249);
and U9941 (N_9941,N_2116,N_868);
nand U9942 (N_9942,N_1500,N_1559);
nor U9943 (N_9943,N_2998,N_838);
or U9944 (N_9944,N_4324,N_3129);
nand U9945 (N_9945,N_1124,N_4448);
or U9946 (N_9946,N_1736,N_996);
nor U9947 (N_9947,N_3114,N_3889);
and U9948 (N_9948,N_425,N_920);
nor U9949 (N_9949,N_2771,N_112);
xnor U9950 (N_9950,N_2967,N_2716);
xor U9951 (N_9951,N_1215,N_1424);
or U9952 (N_9952,N_2038,N_87);
nor U9953 (N_9953,N_1459,N_48);
nand U9954 (N_9954,N_2316,N_2880);
or U9955 (N_9955,N_2331,N_3060);
or U9956 (N_9956,N_1561,N_4171);
and U9957 (N_9957,N_1439,N_2482);
or U9958 (N_9958,N_3059,N_2930);
xor U9959 (N_9959,N_3835,N_140);
nand U9960 (N_9960,N_2031,N_3444);
nor U9961 (N_9961,N_3986,N_3488);
nand U9962 (N_9962,N_4579,N_3349);
or U9963 (N_9963,N_3128,N_2326);
nor U9964 (N_9964,N_4790,N_4910);
nor U9965 (N_9965,N_1740,N_3278);
xor U9966 (N_9966,N_2813,N_3872);
xor U9967 (N_9967,N_1060,N_1298);
or U9968 (N_9968,N_4166,N_4518);
and U9969 (N_9969,N_4125,N_4538);
xnor U9970 (N_9970,N_447,N_4821);
and U9971 (N_9971,N_3959,N_3319);
or U9972 (N_9972,N_3267,N_2989);
nor U9973 (N_9973,N_3147,N_3911);
nor U9974 (N_9974,N_1691,N_812);
or U9975 (N_9975,N_3407,N_30);
or U9976 (N_9976,N_1438,N_1149);
or U9977 (N_9977,N_4829,N_161);
xnor U9978 (N_9978,N_2279,N_4343);
or U9979 (N_9979,N_3229,N_2666);
xnor U9980 (N_9980,N_2122,N_4503);
nand U9981 (N_9981,N_2384,N_4419);
and U9982 (N_9982,N_423,N_1967);
nand U9983 (N_9983,N_3541,N_46);
nand U9984 (N_9984,N_3358,N_511);
xor U9985 (N_9985,N_1081,N_1840);
and U9986 (N_9986,N_3640,N_2022);
nor U9987 (N_9987,N_687,N_4025);
or U9988 (N_9988,N_3085,N_2814);
or U9989 (N_9989,N_1843,N_4686);
or U9990 (N_9990,N_4810,N_3775);
xnor U9991 (N_9991,N_3319,N_1013);
or U9992 (N_9992,N_3842,N_2811);
and U9993 (N_9993,N_2028,N_1293);
nand U9994 (N_9994,N_1121,N_3631);
or U9995 (N_9995,N_761,N_3026);
and U9996 (N_9996,N_772,N_1114);
nand U9997 (N_9997,N_2414,N_1862);
and U9998 (N_9998,N_536,N_3126);
nand U9999 (N_9999,N_2832,N_472);
nand U10000 (N_10000,N_7029,N_5491);
and U10001 (N_10001,N_5381,N_5673);
and U10002 (N_10002,N_7150,N_6077);
and U10003 (N_10003,N_5337,N_5256);
or U10004 (N_10004,N_7425,N_5984);
nand U10005 (N_10005,N_6862,N_6307);
nor U10006 (N_10006,N_7534,N_6145);
and U10007 (N_10007,N_9589,N_9816);
or U10008 (N_10008,N_6331,N_8367);
xor U10009 (N_10009,N_6128,N_9558);
nor U10010 (N_10010,N_9683,N_8541);
nand U10011 (N_10011,N_8113,N_8967);
nand U10012 (N_10012,N_9295,N_7268);
and U10013 (N_10013,N_8843,N_8819);
nand U10014 (N_10014,N_9093,N_5027);
xor U10015 (N_10015,N_9294,N_6433);
xor U10016 (N_10016,N_7048,N_7627);
and U10017 (N_10017,N_9389,N_6515);
or U10018 (N_10018,N_9702,N_5891);
nor U10019 (N_10019,N_8701,N_5841);
xnor U10020 (N_10020,N_7372,N_8879);
nor U10021 (N_10021,N_9238,N_6166);
xnor U10022 (N_10022,N_8384,N_7892);
or U10023 (N_10023,N_9820,N_5534);
nor U10024 (N_10024,N_5261,N_8213);
nand U10025 (N_10025,N_5908,N_6774);
nand U10026 (N_10026,N_9957,N_6035);
and U10027 (N_10027,N_9296,N_6189);
or U10028 (N_10028,N_6414,N_6398);
or U10029 (N_10029,N_8586,N_8506);
xnor U10030 (N_10030,N_9579,N_8450);
and U10031 (N_10031,N_6306,N_9189);
nand U10032 (N_10032,N_7617,N_9614);
xnor U10033 (N_10033,N_6704,N_9607);
and U10034 (N_10034,N_5959,N_7232);
nor U10035 (N_10035,N_8426,N_5203);
xnor U10036 (N_10036,N_7273,N_9317);
nand U10037 (N_10037,N_5761,N_9139);
nand U10038 (N_10038,N_6878,N_7985);
nor U10039 (N_10039,N_9541,N_9948);
nor U10040 (N_10040,N_5039,N_7996);
xor U10041 (N_10041,N_7964,N_9976);
or U10042 (N_10042,N_5016,N_9038);
nor U10043 (N_10043,N_9393,N_9584);
nor U10044 (N_10044,N_8465,N_8300);
or U10045 (N_10045,N_9627,N_6354);
nor U10046 (N_10046,N_5901,N_6164);
xor U10047 (N_10047,N_8456,N_8996);
xnor U10048 (N_10048,N_6048,N_7791);
or U10049 (N_10049,N_6987,N_6881);
nand U10050 (N_10050,N_8614,N_5421);
nand U10051 (N_10051,N_7552,N_7278);
and U10052 (N_10052,N_7885,N_5651);
nor U10053 (N_10053,N_8666,N_6640);
nand U10054 (N_10054,N_8890,N_6495);
and U10055 (N_10055,N_5024,N_7112);
and U10056 (N_10056,N_8258,N_9117);
and U10057 (N_10057,N_9237,N_9719);
and U10058 (N_10058,N_5946,N_9866);
nor U10059 (N_10059,N_9555,N_6126);
xnor U10060 (N_10060,N_5063,N_9568);
and U10061 (N_10061,N_6663,N_7899);
and U10062 (N_10062,N_9698,N_5793);
nor U10063 (N_10063,N_8236,N_5558);
xnor U10064 (N_10064,N_7438,N_5813);
nor U10065 (N_10065,N_9126,N_9367);
nor U10066 (N_10066,N_8404,N_5759);
nand U10067 (N_10067,N_6115,N_9397);
nand U10068 (N_10068,N_7124,N_9751);
or U10069 (N_10069,N_9373,N_5607);
nand U10070 (N_10070,N_6489,N_9082);
nand U10071 (N_10071,N_8853,N_5242);
and U10072 (N_10072,N_7190,N_5300);
or U10073 (N_10073,N_8266,N_7975);
nand U10074 (N_10074,N_5153,N_9372);
or U10075 (N_10075,N_8664,N_7873);
or U10076 (N_10076,N_5232,N_9500);
or U10077 (N_10077,N_6814,N_8772);
nand U10078 (N_10078,N_9713,N_7420);
nor U10079 (N_10079,N_8679,N_5279);
or U10080 (N_10080,N_8974,N_7111);
and U10081 (N_10081,N_5964,N_8119);
nor U10082 (N_10082,N_6131,N_8876);
and U10083 (N_10083,N_9011,N_5129);
and U10084 (N_10084,N_7369,N_8662);
or U10085 (N_10085,N_8729,N_5087);
nand U10086 (N_10086,N_5177,N_5393);
and U10087 (N_10087,N_9973,N_9123);
and U10088 (N_10088,N_5081,N_6948);
nand U10089 (N_10089,N_9546,N_5022);
or U10090 (N_10090,N_5495,N_8167);
or U10091 (N_10091,N_6876,N_7948);
nand U10092 (N_10092,N_9186,N_6154);
nand U10093 (N_10093,N_7168,N_8648);
or U10094 (N_10094,N_5319,N_9076);
nor U10095 (N_10095,N_7570,N_8108);
nor U10096 (N_10096,N_7160,N_7832);
or U10097 (N_10097,N_7915,N_8842);
xnor U10098 (N_10098,N_6159,N_7239);
nor U10099 (N_10099,N_9983,N_8143);
nand U10100 (N_10100,N_5522,N_6431);
nor U10101 (N_10101,N_7847,N_5795);
nor U10102 (N_10102,N_7909,N_5453);
nor U10103 (N_10103,N_7246,N_6929);
nand U10104 (N_10104,N_8329,N_9756);
and U10105 (N_10105,N_9759,N_7220);
nor U10106 (N_10106,N_5896,N_7392);
nor U10107 (N_10107,N_6375,N_8757);
and U10108 (N_10108,N_7411,N_7184);
nor U10109 (N_10109,N_6963,N_6247);
xor U10110 (N_10110,N_7585,N_9239);
and U10111 (N_10111,N_5322,N_8289);
or U10112 (N_10112,N_7368,N_7859);
or U10113 (N_10113,N_8406,N_9599);
nand U10114 (N_10114,N_5125,N_9581);
or U10115 (N_10115,N_7102,N_9963);
and U10116 (N_10116,N_7837,N_9663);
nand U10117 (N_10117,N_8838,N_9498);
and U10118 (N_10118,N_6429,N_9769);
and U10119 (N_10119,N_8668,N_9302);
and U10120 (N_10120,N_5862,N_8282);
or U10121 (N_10121,N_9644,N_9489);
or U10122 (N_10122,N_8179,N_5995);
and U10123 (N_10123,N_7141,N_6295);
and U10124 (N_10124,N_5549,N_6356);
and U10125 (N_10125,N_9703,N_7713);
or U10126 (N_10126,N_5267,N_7366);
or U10127 (N_10127,N_6540,N_5137);
and U10128 (N_10128,N_5556,N_7077);
nor U10129 (N_10129,N_8631,N_8771);
and U10130 (N_10130,N_6969,N_5363);
or U10131 (N_10131,N_5678,N_9320);
xor U10132 (N_10132,N_8116,N_5349);
nand U10133 (N_10133,N_8643,N_8240);
nand U10134 (N_10134,N_7108,N_5914);
nor U10135 (N_10135,N_5683,N_7040);
or U10136 (N_10136,N_7231,N_7787);
xnor U10137 (N_10137,N_8029,N_5796);
nor U10138 (N_10138,N_5680,N_9593);
and U10139 (N_10139,N_5462,N_8122);
nand U10140 (N_10140,N_6090,N_5711);
and U10141 (N_10141,N_5542,N_8502);
nand U10142 (N_10142,N_5539,N_6709);
nor U10143 (N_10143,N_5445,N_8935);
nand U10144 (N_10144,N_9492,N_7092);
nand U10145 (N_10145,N_7076,N_5827);
and U10146 (N_10146,N_5624,N_7854);
nand U10147 (N_10147,N_8459,N_6989);
nand U10148 (N_10148,N_9553,N_6759);
or U10149 (N_10149,N_7062,N_6682);
nand U10150 (N_10150,N_7318,N_9945);
or U10151 (N_10151,N_7148,N_6454);
and U10152 (N_10152,N_9336,N_7628);
nand U10153 (N_10153,N_9376,N_7543);
or U10154 (N_10154,N_7325,N_9423);
or U10155 (N_10155,N_5266,N_8877);
xnor U10156 (N_10156,N_7591,N_6190);
nor U10157 (N_10157,N_8553,N_6024);
or U10158 (N_10158,N_6754,N_8903);
nand U10159 (N_10159,N_8521,N_8626);
or U10160 (N_10160,N_9814,N_7460);
nand U10161 (N_10161,N_5655,N_7050);
xor U10162 (N_10162,N_5224,N_8373);
or U10163 (N_10163,N_6137,N_9802);
nand U10164 (N_10164,N_8339,N_5511);
or U10165 (N_10165,N_8046,N_8234);
xnor U10166 (N_10166,N_8222,N_6171);
or U10167 (N_10167,N_8202,N_8565);
nor U10168 (N_10168,N_7700,N_8888);
or U10169 (N_10169,N_7026,N_6797);
nor U10170 (N_10170,N_9244,N_8128);
nor U10171 (N_10171,N_8627,N_6636);
and U10172 (N_10172,N_6148,N_9267);
nor U10173 (N_10173,N_5978,N_8944);
nand U10174 (N_10174,N_9308,N_5150);
xnor U10175 (N_10175,N_8607,N_5287);
nor U10176 (N_10176,N_6563,N_6986);
and U10177 (N_10177,N_6106,N_9152);
nand U10178 (N_10178,N_9356,N_9691);
and U10179 (N_10179,N_5693,N_8558);
nor U10180 (N_10180,N_8059,N_7690);
nand U10181 (N_10181,N_7991,N_7673);
or U10182 (N_10182,N_8170,N_7021);
nand U10183 (N_10183,N_6758,N_8809);
xor U10184 (N_10184,N_7352,N_8462);
nor U10185 (N_10185,N_9622,N_8957);
nand U10186 (N_10186,N_5653,N_8672);
nor U10187 (N_10187,N_7131,N_9594);
or U10188 (N_10188,N_9853,N_8791);
and U10189 (N_10189,N_7512,N_7398);
nand U10190 (N_10190,N_7637,N_5882);
nand U10191 (N_10191,N_7444,N_7665);
nand U10192 (N_10192,N_8697,N_7868);
xnor U10193 (N_10193,N_8617,N_8682);
or U10194 (N_10194,N_9467,N_6235);
nand U10195 (N_10195,N_6458,N_5632);
or U10196 (N_10196,N_8325,N_7401);
or U10197 (N_10197,N_9327,N_5851);
nand U10198 (N_10198,N_5292,N_7773);
or U10199 (N_10199,N_7751,N_9155);
nor U10200 (N_10200,N_8706,N_7195);
xnor U10201 (N_10201,N_7233,N_7117);
or U10202 (N_10202,N_9758,N_8358);
nor U10203 (N_10203,N_9045,N_5874);
nor U10204 (N_10204,N_5091,N_5760);
or U10205 (N_10205,N_8345,N_6026);
nand U10206 (N_10206,N_6303,N_5702);
and U10207 (N_10207,N_6947,N_8986);
nor U10208 (N_10208,N_8650,N_7661);
xnor U10209 (N_10209,N_8420,N_9564);
or U10210 (N_10210,N_7463,N_7987);
nand U10211 (N_10211,N_6453,N_7770);
or U10212 (N_10212,N_8220,N_9289);
or U10213 (N_10213,N_8782,N_5784);
or U10214 (N_10214,N_9226,N_9242);
nor U10215 (N_10215,N_7450,N_7950);
nand U10216 (N_10216,N_8239,N_5822);
nand U10217 (N_10217,N_9146,N_7484);
xor U10218 (N_10218,N_7490,N_7138);
nand U10219 (N_10219,N_5193,N_8228);
nor U10220 (N_10220,N_9864,N_5158);
and U10221 (N_10221,N_8692,N_6845);
nor U10222 (N_10222,N_8948,N_5392);
nor U10223 (N_10223,N_7286,N_7027);
xnor U10224 (N_10224,N_5777,N_6874);
or U10225 (N_10225,N_7799,N_9209);
nor U10226 (N_10226,N_6464,N_9346);
nor U10227 (N_10227,N_6837,N_9438);
and U10228 (N_10228,N_8628,N_5008);
nand U10229 (N_10229,N_5871,N_6455);
and U10230 (N_10230,N_5043,N_7916);
nand U10231 (N_10231,N_6001,N_5198);
nor U10232 (N_10232,N_5369,N_5560);
xnor U10233 (N_10233,N_8629,N_9109);
or U10234 (N_10234,N_9487,N_9428);
or U10235 (N_10235,N_9441,N_6025);
nor U10236 (N_10236,N_8490,N_8057);
nor U10237 (N_10237,N_6694,N_7664);
nor U10238 (N_10238,N_9081,N_5456);
nand U10239 (N_10239,N_9132,N_6787);
nand U10240 (N_10240,N_6062,N_5899);
nand U10241 (N_10241,N_6953,N_8365);
and U10242 (N_10242,N_6557,N_7279);
and U10243 (N_10243,N_5563,N_6945);
and U10244 (N_10244,N_5566,N_8146);
xnor U10245 (N_10245,N_6582,N_5520);
or U10246 (N_10246,N_5374,N_5781);
xor U10247 (N_10247,N_6252,N_6465);
nand U10248 (N_10248,N_7063,N_8547);
or U10249 (N_10249,N_6346,N_6272);
xor U10250 (N_10250,N_5264,N_8564);
xor U10251 (N_10251,N_6867,N_5706);
nor U10252 (N_10252,N_7227,N_6508);
nand U10253 (N_10253,N_7394,N_9085);
nand U10254 (N_10254,N_8296,N_6655);
nand U10255 (N_10255,N_5960,N_6637);
and U10256 (N_10256,N_8616,N_5648);
nor U10257 (N_10257,N_7419,N_7906);
nand U10258 (N_10258,N_9161,N_7330);
or U10259 (N_10259,N_7497,N_9513);
nand U10260 (N_10260,N_8478,N_5303);
nand U10261 (N_10261,N_6639,N_9672);
and U10262 (N_10262,N_7115,N_6826);
nor U10263 (N_10263,N_8226,N_9723);
xnor U10264 (N_10264,N_9077,N_6114);
nand U10265 (N_10265,N_6542,N_5945);
nor U10266 (N_10266,N_8332,N_7877);
xnor U10267 (N_10267,N_6380,N_5173);
and U10268 (N_10268,N_6543,N_5446);
xor U10269 (N_10269,N_6650,N_9596);
xor U10270 (N_10270,N_9601,N_8267);
and U10271 (N_10271,N_6944,N_5006);
nand U10272 (N_10272,N_7844,N_6498);
and U10273 (N_10273,N_8176,N_9360);
or U10274 (N_10274,N_8973,N_5324);
nor U10275 (N_10275,N_8120,N_8260);
nand U10276 (N_10276,N_9405,N_8264);
nor U10277 (N_10277,N_6225,N_7270);
or U10278 (N_10278,N_7182,N_9141);
nand U10279 (N_10279,N_7742,N_8544);
xnor U10280 (N_10280,N_6233,N_9017);
or U10281 (N_10281,N_9073,N_5357);
and U10282 (N_10282,N_7768,N_5635);
or U10283 (N_10283,N_6262,N_9999);
and U10284 (N_10284,N_5274,N_8423);
or U10285 (N_10285,N_5533,N_8297);
xnor U10286 (N_10286,N_6628,N_9230);
xor U10287 (N_10287,N_7300,N_7446);
xnor U10288 (N_10288,N_6361,N_9274);
or U10289 (N_10289,N_6011,N_6427);
nor U10290 (N_10290,N_6173,N_9124);
nor U10291 (N_10291,N_9909,N_7443);
or U10292 (N_10292,N_6856,N_7536);
or U10293 (N_10293,N_6534,N_5812);
xor U10294 (N_10294,N_9744,N_6996);
and U10295 (N_10295,N_7573,N_5375);
xor U10296 (N_10296,N_9968,N_9083);
or U10297 (N_10297,N_5206,N_6468);
nor U10298 (N_10298,N_5544,N_9611);
or U10299 (N_10299,N_9471,N_5823);
or U10300 (N_10300,N_8596,N_6127);
and U10301 (N_10301,N_5559,N_8827);
xnor U10302 (N_10302,N_5199,N_9775);
or U10303 (N_10303,N_9345,N_6827);
xnor U10304 (N_10304,N_7888,N_7592);
or U10305 (N_10305,N_6526,N_5282);
and U10306 (N_10306,N_6315,N_8018);
nand U10307 (N_10307,N_8577,N_5410);
and U10308 (N_10308,N_7902,N_8537);
or U10309 (N_10309,N_6949,N_8412);
nand U10310 (N_10310,N_8923,N_5097);
or U10311 (N_10311,N_8460,N_6558);
nand U10312 (N_10312,N_5619,N_7819);
nand U10313 (N_10313,N_9470,N_9559);
nor U10314 (N_10314,N_8160,N_5108);
nand U10315 (N_10315,N_7483,N_6098);
nor U10316 (N_10316,N_5957,N_5185);
or U10317 (N_10317,N_9571,N_8349);
and U10318 (N_10318,N_8321,N_5513);
or U10319 (N_10319,N_8955,N_9772);
or U10320 (N_10320,N_8485,N_7531);
xnor U10321 (N_10321,N_6685,N_7660);
nor U10322 (N_10322,N_7113,N_6045);
or U10323 (N_10323,N_7407,N_6799);
and U10324 (N_10324,N_9586,N_5952);
or U10325 (N_10325,N_9907,N_8495);
xor U10326 (N_10326,N_5586,N_5644);
nor U10327 (N_10327,N_7647,N_9578);
xor U10328 (N_10328,N_5877,N_8004);
nor U10329 (N_10329,N_7487,N_6288);
nor U10330 (N_10330,N_5072,N_5638);
or U10331 (N_10331,N_5579,N_7107);
nor U10332 (N_10332,N_7489,N_9191);
and U10333 (N_10333,N_9661,N_6450);
and U10334 (N_10334,N_5132,N_9943);
and U10335 (N_10335,N_9227,N_5483);
or U10336 (N_10336,N_7041,N_5679);
nor U10337 (N_10337,N_5067,N_6491);
xnor U10338 (N_10338,N_9323,N_8510);
or U10339 (N_10339,N_5001,N_9366);
nor U10340 (N_10340,N_5930,N_7545);
or U10341 (N_10341,N_8028,N_5540);
and U10342 (N_10342,N_7039,N_7284);
xnor U10343 (N_10343,N_5262,N_9157);
and U10344 (N_10344,N_5980,N_6755);
nand U10345 (N_10345,N_5926,N_9803);
nand U10346 (N_10346,N_6516,N_8023);
or U10347 (N_10347,N_7669,N_9682);
and U10348 (N_10348,N_7519,N_5478);
or U10349 (N_10349,N_7576,N_6675);
or U10350 (N_10350,N_6898,N_8336);
or U10351 (N_10351,N_9128,N_9898);
nor U10352 (N_10352,N_9605,N_8428);
or U10353 (N_10353,N_9619,N_6941);
nand U10354 (N_10354,N_7777,N_7149);
or U10355 (N_10355,N_6019,N_7695);
nor U10356 (N_10356,N_5828,N_5538);
and U10357 (N_10357,N_8752,N_6181);
xor U10358 (N_10358,N_7099,N_6667);
nand U10359 (N_10359,N_8245,N_5451);
nor U10360 (N_10360,N_9699,N_7693);
nor U10361 (N_10361,N_8445,N_6974);
nor U10362 (N_10362,N_9881,N_7396);
and U10363 (N_10363,N_6139,N_8473);
nand U10364 (N_10364,N_7381,N_6219);
nand U10365 (N_10365,N_7741,N_5143);
and U10366 (N_10366,N_5042,N_9052);
and U10367 (N_10367,N_9746,N_8933);
nor U10368 (N_10368,N_6913,N_6903);
nor U10369 (N_10369,N_9374,N_5863);
or U10370 (N_10370,N_9287,N_9096);
or U10371 (N_10371,N_8235,N_6394);
or U10372 (N_10372,N_9508,N_7785);
nor U10373 (N_10373,N_5134,N_6389);
nand U10374 (N_10374,N_6467,N_9215);
nor U10375 (N_10375,N_5229,N_7729);
nor U10376 (N_10376,N_9646,N_6466);
nand U10377 (N_10377,N_7206,N_8090);
and U10378 (N_10378,N_6406,N_5783);
nor U10379 (N_10379,N_7360,N_9084);
nor U10380 (N_10380,N_9544,N_5931);
and U10381 (N_10381,N_8492,N_6412);
nor U10382 (N_10382,N_7312,N_9949);
nand U10383 (N_10383,N_6719,N_9984);
or U10384 (N_10384,N_7872,N_5804);
or U10385 (N_10385,N_6972,N_8359);
or U10386 (N_10386,N_9163,N_7315);
and U10387 (N_10387,N_9613,N_5346);
nor U10388 (N_10388,N_6073,N_6132);
xor U10389 (N_10389,N_7103,N_9190);
nor U10390 (N_10390,N_7431,N_7927);
xor U10391 (N_10391,N_6917,N_5697);
and U10392 (N_10392,N_9540,N_6251);
nor U10393 (N_10393,N_6842,N_5409);
or U10394 (N_10394,N_5779,N_6055);
nand U10395 (N_10395,N_7262,N_5881);
nand U10396 (N_10396,N_9185,N_9843);
nor U10397 (N_10397,N_7224,N_7941);
xnor U10398 (N_10398,N_9890,N_8277);
nand U10399 (N_10399,N_6665,N_8038);
xnor U10400 (N_10400,N_6485,N_6032);
xor U10401 (N_10401,N_9108,N_6854);
and U10402 (N_10402,N_8764,N_8421);
or U10403 (N_10403,N_6072,N_7603);
nand U10404 (N_10404,N_9788,N_7567);
nor U10405 (N_10405,N_6519,N_6656);
nand U10406 (N_10406,N_9368,N_5014);
or U10407 (N_10407,N_8337,N_9742);
or U10408 (N_10408,N_9955,N_5210);
nand U10409 (N_10409,N_9363,N_6638);
or U10410 (N_10410,N_8139,N_7856);
nand U10411 (N_10411,N_9433,N_7009);
or U10412 (N_10412,N_9595,N_6710);
and U10413 (N_10413,N_8292,N_6984);
and U10414 (N_10414,N_9408,N_9871);
nand U10415 (N_10415,N_7170,N_6499);
or U10416 (N_10416,N_8391,N_5834);
or U10417 (N_10417,N_8612,N_8860);
and U10418 (N_10418,N_7173,N_6452);
nand U10419 (N_10419,N_6662,N_5853);
nor U10420 (N_10420,N_5100,N_9616);
nand U10421 (N_10421,N_9306,N_7340);
nor U10422 (N_10422,N_9561,N_8291);
nand U10423 (N_10423,N_8880,N_8103);
nor U10424 (N_10424,N_7415,N_9449);
or U10425 (N_10425,N_9856,N_7874);
xnor U10426 (N_10426,N_9482,N_8530);
nor U10427 (N_10427,N_6549,N_9026);
and U10428 (N_10428,N_6187,N_7342);
xor U10429 (N_10429,N_9067,N_9525);
and U10430 (N_10430,N_6691,N_6163);
or U10431 (N_10431,N_6313,N_6897);
nor U10432 (N_10432,N_5034,N_6523);
xor U10433 (N_10433,N_6443,N_7763);
and U10434 (N_10434,N_8847,N_5186);
and U10435 (N_10435,N_5219,N_7297);
nand U10436 (N_10436,N_6880,N_5182);
or U10437 (N_10437,N_5344,N_7424);
or U10438 (N_10438,N_7550,N_5856);
nor U10439 (N_10439,N_8951,N_8452);
and U10440 (N_10440,N_8471,N_6424);
or U10441 (N_10441,N_6158,N_5806);
or U10442 (N_10442,N_9673,N_8382);
nand U10443 (N_10443,N_9710,N_6037);
nand U10444 (N_10444,N_7862,N_8507);
nand U10445 (N_10445,N_6280,N_8290);
nor U10446 (N_10446,N_6659,N_6309);
and U10447 (N_10447,N_5608,N_8026);
nand U10448 (N_10448,N_6551,N_6050);
and U10449 (N_10449,N_9645,N_6314);
nand U10450 (N_10450,N_5773,N_8775);
nand U10451 (N_10451,N_9959,N_5291);
nor U10452 (N_10452,N_6900,N_7995);
nand U10453 (N_10453,N_9582,N_8774);
nand U10454 (N_10454,N_8192,N_7358);
nor U10455 (N_10455,N_5713,N_6175);
and U10456 (N_10456,N_5507,N_8956);
or U10457 (N_10457,N_5639,N_7163);
or U10458 (N_10458,N_6513,N_9375);
and U10459 (N_10459,N_5464,N_7080);
nor U10460 (N_10460,N_7462,N_6864);
nor U10461 (N_10461,N_8861,N_7701);
nor U10462 (N_10462,N_5824,N_8403);
or U10463 (N_10463,N_8262,N_5663);
and U10464 (N_10464,N_8640,N_8068);
and U10465 (N_10465,N_5036,N_5936);
or U10466 (N_10466,N_5140,N_9804);
or U10467 (N_10467,N_8323,N_8434);
and U10468 (N_10468,N_7070,N_7612);
xnor U10469 (N_10469,N_5028,N_8939);
nand U10470 (N_10470,N_7495,N_9262);
nor U10471 (N_10471,N_6564,N_5434);
and U10472 (N_10472,N_9770,N_9941);
or U10473 (N_10473,N_5855,N_5972);
nor U10474 (N_10474,N_8091,N_7631);
or U10475 (N_10475,N_6714,N_5127);
nor U10476 (N_10476,N_5289,N_8042);
nand U10477 (N_10477,N_5573,N_6322);
or U10478 (N_10478,N_7765,N_8943);
nand U10479 (N_10479,N_8107,N_8055);
or U10480 (N_10480,N_5668,N_7689);
and U10481 (N_10481,N_6382,N_5041);
xor U10482 (N_10482,N_8166,N_5154);
nand U10483 (N_10483,N_9934,N_9461);
nand U10484 (N_10484,N_6728,N_9557);
nand U10485 (N_10485,N_7094,N_9821);
or U10486 (N_10486,N_8259,N_5993);
and U10487 (N_10487,N_9145,N_6716);
nand U10488 (N_10488,N_8531,N_5345);
nand U10489 (N_10489,N_5971,N_9493);
or U10490 (N_10490,N_5523,N_5766);
xnor U10491 (N_10491,N_6112,N_8309);
nand U10492 (N_10492,N_8658,N_8422);
or U10493 (N_10493,N_9151,N_8844);
and U10494 (N_10494,N_9704,N_8871);
nor U10495 (N_10495,N_8261,N_6832);
xor U10496 (N_10496,N_9502,N_8138);
and U10497 (N_10497,N_8858,N_9811);
or U10498 (N_10498,N_8743,N_8551);
and U10499 (N_10499,N_8357,N_7139);
and U10500 (N_10500,N_8493,N_9893);
and U10501 (N_10501,N_9641,N_9312);
nor U10502 (N_10502,N_7326,N_8499);
and U10503 (N_10503,N_7002,N_8486);
or U10504 (N_10504,N_8824,N_5576);
nor U10505 (N_10505,N_5797,N_8716);
or U10506 (N_10506,N_8416,N_8430);
nand U10507 (N_10507,N_7374,N_9240);
or U10508 (N_10508,N_6666,N_5164);
xor U10509 (N_10509,N_5712,N_6835);
and U10510 (N_10510,N_8745,N_7440);
xor U10511 (N_10511,N_9279,N_6152);
xor U10512 (N_10512,N_7373,N_7316);
or U10513 (N_10513,N_8699,N_5907);
nand U10514 (N_10514,N_9629,N_6844);
or U10515 (N_10515,N_6615,N_9402);
xor U10516 (N_10516,N_8545,N_6866);
xnor U10517 (N_10517,N_7514,N_5735);
or U10518 (N_10518,N_7551,N_7835);
and U10519 (N_10519,N_8831,N_7155);
nand U10520 (N_10520,N_6544,N_6236);
xnor U10521 (N_10521,N_9019,N_5528);
nor U10522 (N_10522,N_9178,N_6124);
or U10523 (N_10523,N_7252,N_9299);
and U10524 (N_10524,N_7736,N_7337);
or U10525 (N_10525,N_7480,N_6919);
xnor U10526 (N_10526,N_5013,N_8301);
xnor U10527 (N_10527,N_7171,N_9718);
and U10528 (N_10528,N_8538,N_9436);
xnor U10529 (N_10529,N_6318,N_9919);
or U10530 (N_10530,N_9040,N_8051);
and U10531 (N_10531,N_8191,N_5471);
nor U10532 (N_10532,N_8010,N_8254);
xor U10533 (N_10533,N_9877,N_9497);
nor U10534 (N_10534,N_5818,N_6609);
or U10535 (N_10535,N_5238,N_5935);
or U10536 (N_10536,N_7533,N_5423);
xor U10537 (N_10537,N_7684,N_9874);
or U10538 (N_10538,N_5671,N_9338);
or U10539 (N_10539,N_6680,N_7005);
or U10540 (N_10540,N_6889,N_8676);
nand U10541 (N_10541,N_6372,N_6237);
nand U10542 (N_10542,N_8735,N_7818);
nand U10543 (N_10543,N_5597,N_9863);
xor U10544 (N_10544,N_6853,N_6447);
or U10545 (N_10545,N_7083,N_6244);
or U10546 (N_10546,N_6363,N_8184);
nor U10547 (N_10547,N_8685,N_8795);
xor U10548 (N_10548,N_8317,N_7164);
or U10549 (N_10549,N_6922,N_7242);
and U10550 (N_10550,N_6568,N_6621);
or U10551 (N_10551,N_7518,N_9575);
and U10552 (N_10552,N_8624,N_8447);
nor U10553 (N_10553,N_9822,N_7556);
nand U10554 (N_10554,N_7380,N_8002);
or U10555 (N_10555,N_7096,N_5277);
nand U10556 (N_10556,N_5843,N_8073);
and U10557 (N_10557,N_9149,N_5077);
or U10558 (N_10558,N_5778,N_9305);
and U10559 (N_10559,N_6925,N_8926);
nand U10560 (N_10560,N_9213,N_5854);
or U10561 (N_10561,N_9325,N_7889);
nor U10562 (N_10562,N_9272,N_6802);
nand U10563 (N_10563,N_6267,N_5156);
nor U10564 (N_10564,N_7375,N_9476);
nor U10565 (N_10565,N_7507,N_9071);
or U10566 (N_10566,N_7175,N_7199);
nor U10567 (N_10567,N_5819,N_8766);
nand U10568 (N_10568,N_8124,N_5599);
nand U10569 (N_10569,N_9315,N_7321);
or U10570 (N_10570,N_8060,N_6764);
or U10571 (N_10571,N_9351,N_5406);
nor U10572 (N_10572,N_8084,N_5403);
nor U10573 (N_10573,N_8121,N_7053);
and U10574 (N_10574,N_6384,N_5519);
nor U10575 (N_10575,N_9730,N_7225);
xnor U10576 (N_10576,N_9278,N_7918);
nor U10577 (N_10577,N_9635,N_8976);
nand U10578 (N_10578,N_6198,N_5352);
and U10579 (N_10579,N_8830,N_6242);
nor U10580 (N_10580,N_7437,N_9386);
and U10581 (N_10581,N_9808,N_8101);
nor U10582 (N_10582,N_6287,N_7882);
and U10583 (N_10583,N_7453,N_5733);
or U10584 (N_10584,N_8189,N_9813);
nand U10585 (N_10585,N_6554,N_8704);
nor U10586 (N_10586,N_5726,N_9411);
or U10587 (N_10587,N_5602,N_7403);
and U10588 (N_10588,N_5356,N_8278);
nor U10589 (N_10589,N_8032,N_6520);
or U10590 (N_10590,N_8649,N_9923);
or U10591 (N_10591,N_6071,N_9130);
or U10592 (N_10592,N_7410,N_9535);
and U10593 (N_10593,N_5376,N_7616);
or U10594 (N_10594,N_7447,N_9565);
nand U10595 (N_10595,N_8177,N_5521);
and U10596 (N_10596,N_5688,N_8950);
nand U10597 (N_10597,N_7848,N_6319);
nor U10598 (N_10598,N_9445,N_9027);
and U10599 (N_10599,N_6119,N_5798);
xnor U10600 (N_10600,N_6275,N_9329);
nor U10601 (N_10601,N_5115,N_8781);
and U10602 (N_10602,N_6747,N_5799);
xor U10603 (N_10603,N_7857,N_8575);
xnor U10604 (N_10604,N_5394,N_9424);
nand U10605 (N_10605,N_9537,N_5050);
nand U10606 (N_10606,N_9643,N_8912);
nor U10607 (N_10607,N_7618,N_6702);
nand U10608 (N_10608,N_8878,N_8513);
or U10609 (N_10609,N_5672,N_8307);
xor U10610 (N_10610,N_8663,N_7580);
or U10611 (N_10611,N_9127,N_6556);
or U10612 (N_10612,N_7351,N_8818);
nor U10613 (N_10613,N_6671,N_6147);
nand U10614 (N_10614,N_6308,N_9666);
and U10615 (N_10615,N_5367,N_6954);
nor U10616 (N_10616,N_8753,N_6773);
and U10617 (N_10617,N_9846,N_6358);
and U10618 (N_10618,N_7824,N_5358);
or U10619 (N_10619,N_5941,N_5477);
nand U10620 (N_10620,N_9324,N_8911);
nand U10621 (N_10621,N_5338,N_9456);
nand U10622 (N_10622,N_6053,N_8364);
xnor U10623 (N_10623,N_5107,N_5467);
nor U10624 (N_10624,N_6461,N_8936);
nand U10625 (N_10625,N_6028,N_6463);
nand U10626 (N_10626,N_9486,N_7681);
and U10627 (N_10627,N_5204,N_5074);
nand U10628 (N_10628,N_6197,N_6950);
and U10629 (N_10629,N_7244,N_5947);
nand U10630 (N_10630,N_8895,N_5331);
nor U10631 (N_10631,N_6988,N_8610);
nor U10632 (N_10632,N_7277,N_8082);
or U10633 (N_10633,N_6739,N_8197);
nand U10634 (N_10634,N_5400,N_6370);
nand U10635 (N_10635,N_6786,N_7678);
or U10636 (N_10636,N_7049,N_8572);
nand U10637 (N_10637,N_7696,N_5235);
and U10638 (N_10638,N_5552,N_5151);
and U10639 (N_10639,N_5840,N_9975);
nand U10640 (N_10640,N_8708,N_6732);
nor U10641 (N_10641,N_5801,N_5103);
nor U10642 (N_10642,N_8645,N_6125);
nand U10643 (N_10643,N_6006,N_7555);
xor U10644 (N_10644,N_5073,N_9511);
xnor U10645 (N_10645,N_9033,N_9815);
or U10646 (N_10646,N_5141,N_6238);
or U10647 (N_10647,N_5079,N_5859);
or U10648 (N_10648,N_9838,N_6102);
nand U10649 (N_10649,N_6352,N_7031);
or U10650 (N_10650,N_8093,N_5414);
nand U10651 (N_10651,N_7583,N_7132);
or U10652 (N_10652,N_6231,N_8893);
and U10653 (N_10653,N_7963,N_7931);
nand U10654 (N_10654,N_9121,N_8335);
nand U10655 (N_10655,N_9088,N_6075);
nor U10656 (N_10656,N_8386,N_5710);
nor U10657 (N_10657,N_5592,N_9852);
nor U10658 (N_10658,N_8457,N_7935);
or U10659 (N_10659,N_9798,N_8968);
and U10660 (N_10660,N_5913,N_9844);
nor U10661 (N_10661,N_8990,N_7750);
nand U10662 (N_10662,N_7356,N_9113);
nand U10663 (N_10663,N_6869,N_9009);
nand U10664 (N_10664,N_7448,N_9369);
nand U10665 (N_10665,N_8437,N_8883);
or U10666 (N_10666,N_6942,N_8137);
and U10667 (N_10667,N_6839,N_7416);
xor U10668 (N_10668,N_6597,N_6715);
or U10669 (N_10669,N_8435,N_5526);
nand U10670 (N_10670,N_7746,N_9285);
nand U10671 (N_10671,N_8310,N_7087);
or U10672 (N_10672,N_9779,N_5380);
nand U10673 (N_10673,N_7558,N_7030);
and U10674 (N_10674,N_9897,N_5694);
nor U10675 (N_10675,N_8402,N_5665);
nand U10676 (N_10676,N_8731,N_6970);
xnor U10677 (N_10677,N_7275,N_6976);
and U10678 (N_10678,N_7529,N_8302);
or U10679 (N_10679,N_6403,N_9122);
or U10680 (N_10680,N_5049,N_6518);
and U10681 (N_10681,N_5354,N_7698);
or U10682 (N_10682,N_6497,N_9654);
nand U10683 (N_10683,N_7295,N_5420);
nor U10684 (N_10684,N_9668,N_5894);
nor U10685 (N_10685,N_7100,N_6397);
xnor U10686 (N_10686,N_9412,N_9906);
or U10687 (N_10687,N_7760,N_8127);
nor U10688 (N_10688,N_7738,N_7359);
and U10689 (N_10689,N_8590,N_5581);
or U10690 (N_10690,N_5588,N_5243);
nand U10691 (N_10691,N_6501,N_7353);
or U10692 (N_10692,N_7659,N_5769);
and U10693 (N_10693,N_6565,N_8850);
or U10694 (N_10694,N_7051,N_7870);
xor U10695 (N_10695,N_6029,N_9875);
and U10696 (N_10696,N_8656,N_8031);
nor U10697 (N_10697,N_7201,N_6122);
xor U10698 (N_10698,N_7137,N_8392);
nor U10699 (N_10699,N_7409,N_6687);
and U10700 (N_10700,N_5377,N_5983);
or U10701 (N_10701,N_6256,N_5280);
and U10702 (N_10702,N_6340,N_7193);
and U10703 (N_10703,N_9824,N_9165);
nor U10704 (N_10704,N_5450,N_6535);
nor U10705 (N_10705,N_9452,N_9933);
nor U10706 (N_10706,N_7413,N_6788);
or U10707 (N_10707,N_7088,N_5172);
or U10708 (N_10708,N_6642,N_8020);
xnor U10709 (N_10709,N_7500,N_7781);
nand U10710 (N_10710,N_7989,N_6830);
nand U10711 (N_10711,N_9685,N_8982);
nor U10712 (N_10712,N_6806,N_6378);
nor U10713 (N_10713,N_6088,N_5977);
or U10714 (N_10714,N_9733,N_6066);
or U10715 (N_10715,N_8836,N_8546);
nand U10716 (N_10716,N_5738,N_5387);
nand U10717 (N_10717,N_7718,N_7455);
nor U10718 (N_10718,N_9726,N_8440);
and U10719 (N_10719,N_7176,N_7811);
nand U10720 (N_10720,N_7801,N_8952);
xor U10721 (N_10721,N_8355,N_5342);
or U10722 (N_10722,N_7217,N_8196);
and U10723 (N_10723,N_8294,N_9328);
nand U10724 (N_10724,N_5833,N_9812);
nor U10725 (N_10725,N_6961,N_6817);
nand U10726 (N_10726,N_8181,N_6706);
or U10727 (N_10727,N_7178,N_5722);
nand U10728 (N_10728,N_6815,N_8770);
and U10729 (N_10729,N_5270,N_8342);
and U10730 (N_10730,N_9103,N_9018);
nor U10731 (N_10731,N_5200,N_9659);
and U10732 (N_10732,N_8219,N_6921);
or U10733 (N_10733,N_7930,N_5562);
or U10734 (N_10734,N_6575,N_5921);
nand U10735 (N_10735,N_6263,N_6417);
or U10736 (N_10736,N_7007,N_6209);
and U10737 (N_10737,N_9316,N_6545);
or U10738 (N_10738,N_6813,N_7951);
nand U10739 (N_10739,N_7761,N_9795);
nor U10740 (N_10740,N_9840,N_5780);
nand U10741 (N_10741,N_7328,N_9477);
and U10742 (N_10742,N_8049,N_6916);
nor U10743 (N_10743,N_5438,N_8037);
nand U10744 (N_10744,N_5391,N_6305);
nor U10745 (N_10745,N_6044,N_8243);
nor U10746 (N_10746,N_7895,N_7749);
nor U10747 (N_10747,N_9917,N_9848);
and U10748 (N_10748,N_6335,N_8475);
nand U10749 (N_10749,N_8899,N_7880);
and U10750 (N_10750,N_9070,N_5750);
nand U10751 (N_10751,N_8543,N_7734);
nand U10752 (N_10752,N_9357,N_8665);
nor U10753 (N_10753,N_5703,N_8750);
and U10754 (N_10754,N_7828,N_9766);
and U10755 (N_10755,N_7059,N_9205);
nor U10756 (N_10756,N_9690,N_9998);
and U10757 (N_10757,N_7274,N_9223);
or U10758 (N_10758,N_7796,N_6861);
or U10759 (N_10759,N_7968,N_9886);
nor U10760 (N_10760,N_6192,N_7855);
and U10761 (N_10761,N_7656,N_6034);
nand U10762 (N_10762,N_9398,N_9232);
nor U10763 (N_10763,N_7630,N_8756);
xnor U10764 (N_10764,N_6993,N_6550);
and U10765 (N_10765,N_5236,N_9131);
xor U10766 (N_10766,N_5417,N_6803);
nand U10767 (N_10767,N_6800,N_8109);
and U10768 (N_10768,N_6631,N_7762);
or U10769 (N_10769,N_9800,N_6172);
and U10770 (N_10770,N_8886,N_7683);
and U10771 (N_10771,N_5618,N_5904);
nand U10772 (N_10772,N_7363,N_8857);
xor U10773 (N_10773,N_7649,N_9610);
or U10774 (N_10774,N_8761,N_7491);
nor U10775 (N_10775,N_9280,N_5918);
nor U10776 (N_10776,N_9761,N_9140);
xor U10777 (N_10777,N_5335,N_7952);
or U10778 (N_10778,N_8864,N_6868);
or U10779 (N_10779,N_9958,N_6428);
xor U10780 (N_10780,N_6548,N_5476);
xor U10781 (N_10781,N_5418,N_8144);
or U10782 (N_10782,N_9114,N_7865);
xnor U10783 (N_10783,N_6614,N_6477);
and U10784 (N_10784,N_8525,N_8651);
xor U10785 (N_10785,N_6940,N_8723);
or U10786 (N_10786,N_7853,N_5981);
nand U10787 (N_10787,N_7691,N_7061);
and U10788 (N_10788,N_7702,N_6250);
or U10789 (N_10789,N_9664,N_8622);
or U10790 (N_10790,N_5922,N_5992);
nand U10791 (N_10791,N_9029,N_9677);
nor U10792 (N_10792,N_8164,N_5516);
and U10793 (N_10793,N_7680,N_8081);
xnor U10794 (N_10794,N_7093,N_9931);
or U10795 (N_10795,N_8885,N_8187);
nand U10796 (N_10796,N_5130,N_7344);
nand U10797 (N_10797,N_6199,N_7081);
nand U10798 (N_10798,N_8581,N_8154);
nor U10799 (N_10799,N_6713,N_5426);
and U10800 (N_10800,N_5098,N_8644);
nand U10801 (N_10801,N_9391,N_9987);
and U10802 (N_10802,N_5985,N_7299);
xnor U10803 (N_10803,N_5176,N_9095);
nand U10804 (N_10804,N_5616,N_5178);
xnor U10805 (N_10805,N_5019,N_5975);
or U10806 (N_10806,N_6323,N_7584);
and U10807 (N_10807,N_8040,N_6183);
nand U10808 (N_10808,N_6436,N_7281);
nand U10809 (N_10809,N_8691,N_9001);
and U10810 (N_10810,N_6184,N_7532);
nor U10811 (N_10811,N_9400,N_8275);
and U10812 (N_10812,N_6731,N_8125);
or U10813 (N_10813,N_6161,N_6529);
and U10814 (N_10814,N_5099,N_8902);
nor U10815 (N_10815,N_7074,N_9276);
or U10816 (N_10816,N_7044,N_9882);
or U10817 (N_10817,N_6555,N_6357);
and U10818 (N_10818,N_8683,N_5740);
and U10819 (N_10819,N_8152,N_5543);
nand U10820 (N_10820,N_5782,N_5561);
nand U10821 (N_10821,N_9080,N_5973);
nor U10822 (N_10822,N_7538,N_5306);
nor U10823 (N_10823,N_9731,N_6681);
and U10824 (N_10824,N_8347,N_9162);
nor U10825 (N_10825,N_9182,N_7641);
and U10826 (N_10826,N_5846,N_6824);
nand U10827 (N_10827,N_5118,N_5060);
and U10828 (N_10828,N_7513,N_5880);
nand U10829 (N_10829,N_5872,N_7127);
and U10830 (N_10830,N_6052,N_6255);
nand U10831 (N_10831,N_8334,N_7613);
nor U10832 (N_10832,N_5775,N_6999);
and U10833 (N_10833,N_6368,N_5944);
nor U10834 (N_10834,N_9776,N_9164);
nand U10835 (N_10835,N_5878,N_6076);
or U10836 (N_10836,N_8727,N_8512);
and U10837 (N_10837,N_7391,N_6276);
nand U10838 (N_10838,N_7219,N_5168);
or U10839 (N_10839,N_6528,N_9443);
xnor U10840 (N_10840,N_5258,N_8767);
xor U10841 (N_10841,N_9762,N_9694);
nand U10842 (N_10842,N_8961,N_9588);
or U10843 (N_10843,N_8837,N_9168);
or U10844 (N_10844,N_6517,N_8806);
and U10845 (N_10845,N_7629,N_8374);
nand U10846 (N_10846,N_5989,N_8242);
nand U10847 (N_10847,N_5844,N_9284);
and U10848 (N_10848,N_5626,N_7350);
nand U10849 (N_10849,N_5961,N_9064);
nand U10850 (N_10850,N_7587,N_9252);
nor U10851 (N_10851,N_8027,N_6456);
and U10852 (N_10852,N_5368,N_7456);
nor U10853 (N_10853,N_8305,N_5084);
and U10854 (N_10854,N_7162,N_8937);
nor U10855 (N_10855,N_7308,N_8589);
nand U10856 (N_10856,N_6195,N_7815);
or U10857 (N_10857,N_9501,N_6855);
nor U10858 (N_10858,N_7999,N_6629);
nor U10859 (N_10859,N_6757,N_8805);
and U10860 (N_10860,N_8870,N_6581);
or U10861 (N_10861,N_8945,N_9965);
nor U10862 (N_10862,N_9066,N_9700);
or U10863 (N_10863,N_5911,N_7073);
xor U10864 (N_10864,N_5691,N_9003);
nor U10865 (N_10865,N_5257,N_9826);
nor U10866 (N_10866,N_8295,N_9636);
nor U10867 (N_10867,N_9175,N_8520);
nor U10868 (N_10868,N_8832,N_9377);
xor U10869 (N_10869,N_9167,N_8971);
and U10870 (N_10870,N_8464,N_8463);
nor U10871 (N_10871,N_5407,N_7091);
nor U10872 (N_10872,N_7898,N_6481);
nor U10873 (N_10873,N_7471,N_9900);
and U10874 (N_10874,N_5585,N_5399);
or U10875 (N_10875,N_5987,N_7920);
nor U10876 (N_10876,N_6469,N_7384);
nand U10877 (N_10877,N_9002,N_9717);
nand U10878 (N_10878,N_8225,N_7046);
or U10879 (N_10879,N_9333,N_5009);
xnor U10880 (N_10880,N_6785,N_8088);
nor U10881 (N_10881,N_6310,N_9505);
or U10882 (N_10882,N_7177,N_8396);
or U10883 (N_10883,N_9609,N_7967);
nand U10884 (N_10884,N_8696,N_9942);
and U10885 (N_10885,N_7622,N_6249);
nor U10886 (N_10886,N_9354,N_5969);
or U10887 (N_10887,N_5615,N_9010);
nor U10888 (N_10888,N_8062,N_7530);
and U10889 (N_10889,N_5033,N_9392);
nor U10890 (N_10890,N_7594,N_9286);
nor U10891 (N_10891,N_7737,N_9519);
or U10892 (N_10892,N_7636,N_5574);
nand U10893 (N_10893,N_5505,N_9991);
or U10894 (N_10894,N_7564,N_5040);
or U10895 (N_10895,N_9133,N_6129);
nor U10896 (N_10896,N_6381,N_7581);
or U10897 (N_10897,N_6277,N_8618);
and U10898 (N_10898,N_7745,N_5756);
nor U10899 (N_10899,N_6507,N_7134);
and U10900 (N_10900,N_9792,N_6511);
nand U10901 (N_10901,N_7897,N_6364);
or U10902 (N_10902,N_9466,N_7065);
or U10903 (N_10903,N_9962,N_9410);
nand U10904 (N_10904,N_9913,N_8855);
nor U10905 (N_10905,N_8198,N_5590);
nor U10906 (N_10906,N_6644,N_5541);
nand U10907 (N_10907,N_8419,N_7304);
and U10908 (N_10908,N_7012,N_6095);
and U10909 (N_10909,N_9255,N_6645);
nand U10910 (N_10910,N_6008,N_6435);
nand U10911 (N_10911,N_7884,N_5617);
and U10912 (N_10912,N_5734,N_7667);
or U10913 (N_10913,N_5545,N_9522);
nor U10914 (N_10914,N_5546,N_9058);
nor U10915 (N_10915,N_8360,N_6718);
and U10916 (N_10916,N_8033,N_9036);
or U10917 (N_10917,N_7687,N_6777);
nor U10918 (N_10918,N_7960,N_9359);
or U10919 (N_10919,N_6349,N_8670);
and U10920 (N_10920,N_6030,N_7582);
nor U10921 (N_10921,N_9094,N_7003);
or U10922 (N_10922,N_9459,N_7314);
nand U10923 (N_10923,N_6261,N_7976);
nor U10924 (N_10924,N_5923,N_8248);
nand U10925 (N_10925,N_6847,N_8401);
and U10926 (N_10926,N_9399,N_6320);
nor U10927 (N_10927,N_6791,N_7621);
nand U10928 (N_10928,N_9434,N_5916);
or U10929 (N_10929,N_9835,N_6343);
or U10930 (N_10930,N_8778,N_6760);
xnor U10931 (N_10931,N_6711,N_7451);
and U10932 (N_10932,N_5056,N_5379);
and U10933 (N_10933,N_6943,N_6010);
nor U10934 (N_10934,N_5658,N_7331);
or U10935 (N_10935,N_8250,N_5976);
or U10936 (N_10936,N_7609,N_5070);
nor U10937 (N_10937,N_6617,N_6478);
nor U10938 (N_10938,N_7317,N_5611);
and U10939 (N_10939,N_6783,N_6218);
xor U10940 (N_10940,N_8536,N_9834);
or U10941 (N_10941,N_6206,N_8045);
nand U10942 (N_10942,N_9830,N_9488);
xor U10943 (N_10943,N_8110,N_6273);
xnor U10944 (N_10944,N_7934,N_5194);
xnor U10945 (N_10945,N_5002,N_8773);
nor U10946 (N_10946,N_7982,N_8720);
or U10947 (N_10947,N_8442,N_7473);
or U10948 (N_10948,N_7540,N_7959);
nor U10949 (N_10949,N_7614,N_9339);
nand U10950 (N_10950,N_6657,N_9725);
or U10951 (N_10951,N_7548,N_8263);
and U10952 (N_10952,N_9208,N_7140);
nand U10953 (N_10953,N_9905,N_6598);
and U10954 (N_10954,N_8299,N_7639);
or U10955 (N_10955,N_9341,N_6312);
nor U10956 (N_10956,N_9604,N_8015);
nor U10957 (N_10957,N_9684,N_7377);
and U10958 (N_10958,N_5083,N_7642);
nor U10959 (N_10959,N_6690,N_9118);
nor U10960 (N_10960,N_9777,N_8280);
or U10961 (N_10961,N_9515,N_8568);
nand U10962 (N_10962,N_9396,N_6248);
and U10963 (N_10963,N_9174,N_8992);
nand U10964 (N_10964,N_5498,N_8598);
nand U10965 (N_10965,N_9817,N_8733);
and U10966 (N_10966,N_5920,N_8799);
nor U10967 (N_10967,N_5101,N_9220);
nand U10968 (N_10968,N_9880,N_6373);
nor U10969 (N_10969,N_9764,N_5312);
and U10970 (N_10970,N_6220,N_7910);
nor U10971 (N_10971,N_8671,N_7984);
nand U10972 (N_10972,N_9883,N_9181);
nor U10973 (N_10973,N_9720,N_7633);
or U10974 (N_10974,N_9687,N_5512);
nand U10975 (N_10975,N_6822,N_6259);
nor U10976 (N_10976,N_5152,N_5102);
nor U10977 (N_10977,N_9797,N_8287);
or U10978 (N_10978,N_9602,N_8013);
nor U10979 (N_10979,N_8056,N_9554);
and U10980 (N_10980,N_5772,N_9137);
and U10981 (N_10981,N_8344,N_5517);
or U10982 (N_10982,N_7623,N_5385);
nor U10983 (N_10983,N_7611,N_8080);
nand U10984 (N_10984,N_9946,N_6333);
or U10985 (N_10985,N_8601,N_9136);
nand U10986 (N_10986,N_5316,N_6138);
nand U10987 (N_10987,N_5054,N_6487);
nand U10988 (N_10988,N_7912,N_5903);
and U10989 (N_10989,N_7238,N_7549);
nor U10990 (N_10990,N_9606,N_6510);
nand U10991 (N_10991,N_7338,N_7154);
nor U10992 (N_10992,N_5116,N_5869);
and U10993 (N_10993,N_9148,N_8570);
nor U10994 (N_10994,N_6063,N_9981);
and U10995 (N_10995,N_6896,N_9891);
or U10996 (N_10996,N_5327,N_8779);
or U10997 (N_10997,N_9598,N_6560);
nand U10998 (N_10998,N_6586,N_5605);
and U10999 (N_10999,N_5317,N_5660);
or U11000 (N_11000,N_7833,N_8472);
nand U11001 (N_11001,N_8150,N_7893);
nand U11002 (N_11002,N_5589,N_5181);
xnor U11003 (N_11003,N_6438,N_7841);
nand U11004 (N_11004,N_5187,N_7435);
nor U11005 (N_11005,N_9712,N_8095);
and U11006 (N_11006,N_5578,N_6230);
nand U11007 (N_11007,N_9825,N_5440);
or U11008 (N_11008,N_9929,N_9472);
or U11009 (N_11009,N_8318,N_6770);
nand U11010 (N_11010,N_7349,N_8489);
nand U11011 (N_11011,N_5765,N_7879);
and U11012 (N_11012,N_9986,N_8350);
nand U11013 (N_11013,N_9539,N_5527);
or U11014 (N_11014,N_6239,N_9748);
nand U11015 (N_11015,N_9980,N_9600);
nor U11016 (N_11016,N_7405,N_8098);
nand U11017 (N_11017,N_7645,N_7704);
nand U11018 (N_11018,N_7804,N_7842);
nor U11019 (N_11019,N_6298,N_8652);
and U11020 (N_11020,N_8052,N_7037);
nand U11021 (N_11021,N_5020,N_5419);
nor U11022 (N_11022,N_7652,N_9526);
or U11023 (N_11023,N_6633,N_5847);
nand U11024 (N_11024,N_8910,N_9016);
or U11025 (N_11025,N_9166,N_6771);
or U11026 (N_11026,N_6794,N_7624);
or U11027 (N_11027,N_9403,N_6336);
nor U11028 (N_11028,N_8385,N_5582);
xor U11029 (N_11029,N_6326,N_7301);
nor U11030 (N_11030,N_6143,N_5248);
nor U11031 (N_11031,N_9628,N_6292);
nand U11032 (N_11032,N_8409,N_6243);
and U11033 (N_11033,N_7539,N_7599);
nand U11034 (N_11034,N_6882,N_9427);
nor U11035 (N_11035,N_5239,N_8237);
or U11036 (N_11036,N_7235,N_7060);
or U11037 (N_11037,N_7216,N_6174);
or U11038 (N_11038,N_9633,N_7180);
or U11039 (N_11039,N_7387,N_8988);
and U11040 (N_11040,N_7501,N_9912);
and U11041 (N_11041,N_6672,N_6514);
and U11042 (N_11042,N_8194,N_7896);
nor U11043 (N_11043,N_5122,N_8717);
xnor U11044 (N_11044,N_5089,N_8388);
and U11045 (N_11045,N_8588,N_5888);
nand U11046 (N_11046,N_8389,N_6746);
nand U11047 (N_11047,N_5537,N_5988);
or U11048 (N_11048,N_5479,N_6991);
and U11049 (N_11049,N_7032,N_8579);
or U11050 (N_11050,N_8592,N_7574);
nor U11051 (N_11051,N_5736,N_6330);
nand U11052 (N_11052,N_6960,N_9925);
and U11053 (N_11053,N_8025,N_5723);
xor U11054 (N_11054,N_5979,N_8814);
or U11055 (N_11055,N_8675,N_9469);
or U11056 (N_11056,N_8705,N_8311);
and U11057 (N_11057,N_7554,N_6068);
nor U11058 (N_11058,N_6439,N_6587);
nor U11059 (N_11059,N_5080,N_8690);
nand U11060 (N_11060,N_9679,N_9037);
nand U11061 (N_11061,N_5365,N_9736);
and U11062 (N_11062,N_6966,N_7064);
nor U11063 (N_11063,N_9224,N_6360);
nand U11064 (N_11064,N_7475,N_5313);
or U11065 (N_11065,N_8079,N_6332);
nand U11066 (N_11066,N_8892,N_6580);
and U11067 (N_11067,N_5384,N_6170);
nor U11068 (N_11068,N_7146,N_5484);
nand U11069 (N_11069,N_5603,N_9101);
and U11070 (N_11070,N_9806,N_9523);
nor U11071 (N_11071,N_7106,N_8063);
nor U11072 (N_11072,N_6805,N_8784);
or U11073 (N_11073,N_9454,N_5052);
or U11074 (N_11074,N_7917,N_7675);
xor U11075 (N_11075,N_5684,N_5536);
nor U11076 (N_11076,N_6084,N_5458);
and U11077 (N_11077,N_7082,N_5216);
nor U11078 (N_11078,N_6067,N_7499);
xor U11079 (N_11079,N_7016,N_8458);
and U11080 (N_11080,N_6257,N_6254);
and U11081 (N_11081,N_9885,N_6484);
nand U11082 (N_11082,N_5751,N_9150);
and U11083 (N_11083,N_9384,N_5790);
xor U11084 (N_11084,N_5305,N_8635);
and U11085 (N_11085,N_9416,N_8252);
xnor U11086 (N_11086,N_9888,N_7213);
nand U11087 (N_11087,N_8839,N_5431);
or U11088 (N_11088,N_5929,N_5207);
and U11089 (N_11089,N_8229,N_5093);
nand U11090 (N_11090,N_8474,N_7670);
nor U11091 (N_11091,N_7204,N_5336);
and U11092 (N_11092,N_7825,N_5934);
or U11093 (N_11093,N_7586,N_7682);
and U11094 (N_11094,N_7309,N_7426);
or U11095 (N_11095,N_5791,N_5412);
nor U11096 (N_11096,N_8749,N_5104);
and U11097 (N_11097,N_9335,N_7778);
xor U11098 (N_11098,N_9079,N_5725);
nor U11099 (N_11099,N_5378,N_5076);
or U11100 (N_11100,N_9681,N_8970);
nand U11101 (N_11101,N_5136,N_9358);
nand U11102 (N_11102,N_6362,N_5622);
nand U11103 (N_11103,N_8739,N_8114);
or U11104 (N_11104,N_9550,N_6599);
xnor U11105 (N_11105,N_8375,N_7537);
and U11106 (N_11106,N_9978,N_6836);
nand U11107 (N_11107,N_7123,N_5776);
and U11108 (N_11108,N_6038,N_9431);
and U11109 (N_11109,N_8072,N_9741);
or U11110 (N_11110,N_8657,N_7245);
or U11111 (N_11111,N_5329,N_6415);
and U11112 (N_11112,N_9518,N_7354);
or U11113 (N_11113,N_5860,N_7157);
and U11114 (N_11114,N_9310,N_5943);
nor U11115 (N_11115,N_8835,N_6105);
or U11116 (N_11116,N_8216,N_6080);
nor U11117 (N_11117,N_5850,N_9207);
xnor U11118 (N_11118,N_6325,N_7610);
nand U11119 (N_11119,N_7043,N_5731);
nor U11120 (N_11120,N_8978,N_8660);
nor U11121 (N_11121,N_7940,N_8210);
nor U11122 (N_11122,N_8158,N_9290);
or U11123 (N_11123,N_5900,N_5237);
nor U11124 (N_11124,N_5595,N_7969);
or U11125 (N_11125,N_9615,N_5647);
and U11126 (N_11126,N_7229,N_5755);
and U11127 (N_11127,N_7109,N_8625);
nand U11128 (N_11128,N_8776,N_6608);
nand U11129 (N_11129,N_7887,N_9928);
nor U11130 (N_11130,N_5792,N_6393);
nand U11131 (N_11131,N_7436,N_8387);
or U11132 (N_11132,N_9382,N_9649);
nand U11133 (N_11133,N_7942,N_6094);
nor U11134 (N_11134,N_9850,N_9063);
nor U11135 (N_11135,N_9738,N_9939);
and U11136 (N_11136,N_7677,N_9444);
nand U11137 (N_11137,N_6647,N_9196);
nor U11138 (N_11138,N_9617,N_6379);
nor U11139 (N_11139,N_7595,N_7932);
nor U11140 (N_11140,N_7753,N_7863);
nor U11141 (N_11141,N_7339,N_8284);
nand U11142 (N_11142,N_5686,N_6353);
or U11143 (N_11143,N_8964,N_9231);
and U11144 (N_11144,N_6562,N_6046);
or U11145 (N_11145,N_6938,N_9862);
nand U11146 (N_11146,N_9510,N_9246);
or U11147 (N_11147,N_6753,N_8600);
nor U11148 (N_11148,N_9895,N_7395);
nand U11149 (N_11149,N_5311,N_6890);
or U11150 (N_11150,N_6395,N_9785);
nor U11151 (N_11151,N_9495,N_8372);
nor U11152 (N_11152,N_7803,N_6420);
and U11153 (N_11153,N_6111,N_5836);
nor U11154 (N_11154,N_6057,N_5816);
and U11155 (N_11155,N_9969,N_7869);
xnor U11156 (N_11156,N_6521,N_9670);
or U11157 (N_11157,N_9831,N_6533);
xnor U11158 (N_11158,N_9091,N_8997);
and U11159 (N_11159,N_5746,N_8783);
nand U11160 (N_11160,N_7846,N_5494);
or U11161 (N_11161,N_7161,N_6658);
and U11162 (N_11162,N_8306,N_7757);
or U11163 (N_11163,N_8759,N_7291);
xnor U11164 (N_11164,N_6914,N_6693);
and U11165 (N_11165,N_8074,N_5430);
xor U11166 (N_11166,N_7441,N_8859);
and U11167 (N_11167,N_7679,N_8041);
nor U11168 (N_11168,N_7055,N_9851);
or U11169 (N_11169,N_7784,N_6494);
xor U11170 (N_11170,N_5572,N_9119);
and U11171 (N_11171,N_8340,N_7755);
nor U11172 (N_11172,N_8980,N_8233);
or U11173 (N_11173,N_7364,N_5701);
nand U11174 (N_11174,N_8597,N_7197);
nor U11175 (N_11175,N_7790,N_6997);
or U11176 (N_11176,N_5905,N_9407);
nor U11177 (N_11177,N_9144,N_9724);
and U11178 (N_11178,N_5474,N_5596);
nor U11179 (N_11179,N_5716,N_5753);
or U11180 (N_11180,N_5302,N_8561);
and U11181 (N_11181,N_5055,N_7020);
nor U11182 (N_11182,N_6405,N_8071);
xor U11183 (N_11183,N_5010,N_8965);
or U11184 (N_11184,N_5999,N_6559);
nand U11185 (N_11185,N_5743,N_8741);
nand U11186 (N_11186,N_8438,N_6144);
nor U11187 (N_11187,N_8810,N_9217);
nor U11188 (N_11188,N_9714,N_9827);
nor U11189 (N_11189,N_7265,N_7923);
or U11190 (N_11190,N_9035,N_5299);
nand U11191 (N_11191,N_8722,N_9479);
nor U11192 (N_11192,N_7598,N_6857);
nor U11193 (N_11193,N_6725,N_6451);
nand U11194 (N_11194,N_6100,N_7988);
nand U11195 (N_11195,N_9061,N_6592);
nand U11196 (N_11196,N_7367,N_5473);
nor U11197 (N_11197,N_9632,N_5179);
nand U11198 (N_11198,N_7600,N_6936);
nand U11199 (N_11199,N_5424,N_8368);
nor U11200 (N_11200,N_7185,N_5045);
and U11201 (N_11201,N_8742,N_7089);
nor U11202 (N_11202,N_9833,N_5112);
or U11203 (N_11203,N_6371,N_7634);
nor U11204 (N_11204,N_7929,N_8792);
nand U11205 (N_11205,N_6021,N_9006);
and U11206 (N_11206,N_9050,N_7943);
nand U11207 (N_11207,N_5883,N_7194);
nand U11208 (N_11208,N_9049,N_8481);
nand U11209 (N_11209,N_6081,N_6977);
nor U11210 (N_11210,N_9532,N_9865);
nand U11211 (N_11211,N_7119,N_6337);
and U11212 (N_11212,N_8411,N_6223);
xnor U11213 (N_11213,N_5752,N_8681);
and U11214 (N_11214,N_7223,N_9799);
and U11215 (N_11215,N_6894,N_5714);
or U11216 (N_11216,N_6795,N_5057);
or U11217 (N_11217,N_9536,N_6872);
and U11218 (N_11218,N_9849,N_8215);
or U11219 (N_11219,N_5832,N_7775);
or U11220 (N_11220,N_8362,N_8163);
nor U11221 (N_11221,N_6493,N_8414);
nand U11222 (N_11222,N_9216,N_5048);
nor U11223 (N_11223,N_6512,N_9675);
nand U11224 (N_11224,N_8257,N_6221);
nand U11225 (N_11225,N_9747,N_8083);
and U11226 (N_11226,N_5225,N_7477);
nor U11227 (N_11227,N_6180,N_7970);
xor U11228 (N_11228,N_8270,N_6522);
nand U11229 (N_11229,N_5260,N_7752);
or U11230 (N_11230,N_8608,N_7939);
nand U11231 (N_11231,N_9915,N_5664);
nand U11232 (N_11232,N_8130,N_5004);
nor U11233 (N_11233,N_8035,N_9387);
nand U11234 (N_11234,N_6858,N_7481);
and U11235 (N_11235,N_8554,N_8142);
or U11236 (N_11236,N_9911,N_5144);
nand U11237 (N_11237,N_6085,N_8793);
nand U11238 (N_11238,N_7520,N_7744);
and U11239 (N_11239,N_7280,N_5214);
nand U11240 (N_11240,N_5030,N_5709);
and U11241 (N_11241,N_8755,N_7571);
or U11242 (N_11242,N_6775,N_6214);
or U11243 (N_11243,N_6348,N_5623);
nor U11244 (N_11244,N_9309,N_5320);
nand U11245 (N_11245,N_5139,N_5593);
nor U11246 (N_11246,N_5811,N_6031);
xnor U11247 (N_11247,N_7467,N_5974);
nor U11248 (N_11248,N_9755,N_5296);
and U11249 (N_11249,N_7780,N_5459);
nand U11250 (N_11250,N_6643,N_6091);
and U11251 (N_11251,N_7503,N_8889);
nand U11252 (N_11252,N_9993,N_5220);
nand U11253 (N_11253,N_7544,N_9771);
nor U11254 (N_11254,N_9861,N_8322);
or U11255 (N_11255,N_6885,N_7504);
nand U11256 (N_11256,N_7875,N_7607);
xor U11257 (N_11257,N_8915,N_8427);
nand U11258 (N_11258,N_7390,N_6437);
and U11259 (N_11259,N_7992,N_8574);
and U11260 (N_11260,N_7258,N_9689);
nor U11261 (N_11261,N_6449,N_5402);
and U11262 (N_11262,N_5770,N_8667);
nor U11263 (N_11263,N_5271,N_6086);
and U11264 (N_11264,N_5690,N_6390);
or U11265 (N_11265,N_9090,N_8153);
nor U11266 (N_11266,N_6594,N_7058);
and U11267 (N_11267,N_6388,N_6400);
nand U11268 (N_11268,N_5124,N_9179);
and U11269 (N_11269,N_6804,N_5645);
nand U11270 (N_11270,N_8816,N_7866);
nor U11271 (N_11271,N_5675,N_7240);
nand U11272 (N_11272,N_8221,N_6937);
nand U11273 (N_11273,N_9184,N_6553);
or U11274 (N_11274,N_7883,N_9810);
nor U11275 (N_11275,N_5007,N_9364);
and U11276 (N_11276,N_6488,N_7247);
nor U11277 (N_11277,N_5347,N_8132);
nand U11278 (N_11278,N_8787,N_5227);
nor U11279 (N_11279,N_8934,N_9765);
or U11280 (N_11280,N_9383,N_6923);
or U11281 (N_11281,N_8630,N_7805);
nand U11282 (N_11282,N_8175,N_5965);
nor U11283 (N_11283,N_7019,N_7911);
xor U11284 (N_11284,N_6476,N_5276);
or U11285 (N_11285,N_6920,N_5191);
nor U11286 (N_11286,N_7608,N_6374);
or U11287 (N_11287,N_7015,N_8637);
nor U11288 (N_11288,N_6082,N_8381);
or U11289 (N_11289,N_7807,N_5455);
or U11290 (N_11290,N_8746,N_7283);
xnor U11291 (N_11291,N_9884,N_6660);
nor U11292 (N_11292,N_7836,N_7071);
or U11293 (N_11293,N_9078,N_9648);
xnor U11294 (N_11294,N_6089,N_7459);
and U11295 (N_11295,N_9361,N_9952);
or U11296 (N_11296,N_9206,N_7822);
nor U11297 (N_11297,N_9597,N_5475);
nor U11298 (N_11298,N_8959,N_8431);
or U11299 (N_11299,N_5065,N_5642);
or U11300 (N_11300,N_9878,N_8505);
xor U11301 (N_11301,N_6840,N_9521);
and U11302 (N_11302,N_6016,N_7957);
xnor U11303 (N_11303,N_5386,N_8882);
or U11304 (N_11304,N_8736,N_6524);
and U11305 (N_11305,N_9022,N_8604);
or U11306 (N_11306,N_8527,N_5805);
or U11307 (N_11307,N_7086,N_5457);
nor U11308 (N_11308,N_8953,N_9961);
and U11309 (N_11309,N_7509,N_5940);
or U11310 (N_11310,N_5253,N_6064);
or U11311 (N_11311,N_6232,N_9592);
nand U11312 (N_11312,N_8123,N_7516);
nor U11313 (N_11313,N_5404,N_7808);
xor U11314 (N_11314,N_6809,N_8748);
and U11315 (N_11315,N_7135,N_7189);
nor U11316 (N_11316,N_7813,N_7936);
nand U11317 (N_11317,N_9680,N_9583);
nor U11318 (N_11318,N_5201,N_7191);
xnor U11319 (N_11319,N_7136,N_7215);
nand U11320 (N_11320,N_5870,N_5997);
or U11321 (N_11321,N_7018,N_8788);
or U11322 (N_11322,N_6169,N_9086);
nand U11323 (N_11323,N_8212,N_8854);
and U11324 (N_11324,N_6538,N_5339);
nor U11325 (N_11325,N_7913,N_6618);
or U11326 (N_11326,N_5205,N_6846);
or U11327 (N_11327,N_7269,N_7493);
nor U11328 (N_11328,N_8206,N_5531);
nand U11329 (N_11329,N_9120,N_8754);
nor U11330 (N_11330,N_9807,N_7035);
or U11331 (N_11331,N_5502,N_7526);
nor U11332 (N_11332,N_9620,N_9839);
nor U11333 (N_11333,N_9264,N_5436);
and U11334 (N_11334,N_9977,N_5432);
or U11335 (N_11335,N_6994,N_8983);
or U11336 (N_11336,N_8920,N_7408);
nor U11337 (N_11337,N_8201,N_5937);
nor U11338 (N_11338,N_8274,N_8789);
or U11339 (N_11339,N_8535,N_8719);
or U11340 (N_11340,N_9572,N_6022);
nor U11341 (N_11341,N_5086,N_7042);
or U11342 (N_11342,N_9529,N_5401);
nor U11343 (N_11343,N_9918,N_9988);
nand U11344 (N_11344,N_6156,N_6007);
xor U11345 (N_11345,N_5948,N_7404);
nand U11346 (N_11346,N_7129,N_6342);
nor U11347 (N_11347,N_6796,N_5069);
xnor U11348 (N_11348,N_9790,N_8655);
or U11349 (N_11349,N_7797,N_8841);
nor U11350 (N_11350,N_5986,N_6446);
or U11351 (N_11351,N_7648,N_6579);
nor U11352 (N_11352,N_7143,N_7288);
or U11353 (N_11353,N_8066,N_8896);
nand U11354 (N_11354,N_7014,N_6475);
nand U11355 (N_11355,N_5395,N_6178);
nor U11356 (N_11356,N_7774,N_7821);
xnor U11357 (N_11357,N_9030,N_7056);
xnor U11358 (N_11358,N_7452,N_5398);
and U11359 (N_11359,N_8703,N_9254);
xnor U11360 (N_11360,N_8715,N_8917);
xnor U11361 (N_11361,N_8030,N_6445);
nor U11362 (N_11362,N_9562,N_5362);
and U11363 (N_11363,N_8484,N_8514);
and U11364 (N_11364,N_5128,N_8613);
or U11365 (N_11365,N_8931,N_9551);
and U11366 (N_11366,N_8740,N_9054);
and U11367 (N_11367,N_7726,N_5366);
nor U11368 (N_11368,N_5068,N_6176);
xor U11369 (N_11369,N_5953,N_6736);
nand U11370 (N_11370,N_7820,N_7133);
and U11371 (N_11371,N_6430,N_7938);
nand U11372 (N_11372,N_9809,N_9421);
nand U11373 (N_11373,N_9187,N_7908);
or U11374 (N_11374,N_5875,N_6536);
or U11375 (N_11375,N_9543,N_5197);
and U11376 (N_11376,N_6578,N_6762);
or U11377 (N_11377,N_8508,N_8863);
and U11378 (N_11378,N_5482,N_5075);
or U11379 (N_11379,N_5785,N_5023);
nand U11380 (N_11380,N_7429,N_6653);
or U11381 (N_11381,N_5463,N_5550);
or U11382 (N_11382,N_7789,N_7457);
or U11383 (N_11383,N_6459,N_8092);
xnor U11384 (N_11384,N_9966,N_7830);
nor U11385 (N_11385,N_9112,N_9496);
nand U11386 (N_11386,N_7560,N_7023);
and U11387 (N_11387,N_6473,N_7166);
nand U11388 (N_11388,N_7717,N_8744);
xor U11389 (N_11389,N_6224,N_8845);
nand U11390 (N_11390,N_6967,N_6193);
nand U11391 (N_11391,N_7772,N_8455);
or U11392 (N_11392,N_6772,N_8320);
xnor U11393 (N_11393,N_7925,N_5025);
nand U11394 (N_11394,N_6284,N_8413);
and U11395 (N_11395,N_5890,N_9927);
nand U11396 (N_11396,N_5382,N_9549);
and U11397 (N_11397,N_9491,N_5272);
xnor U11398 (N_11398,N_8012,N_5893);
and U11399 (N_11399,N_9288,N_6848);
or U11400 (N_11400,N_5000,N_7771);
nand U11401 (N_11401,N_7476,N_5032);
or U11402 (N_11402,N_6059,N_6392);
xnor U11403 (N_11403,N_5610,N_6712);
xor U11404 (N_11404,N_6282,N_8583);
or U11405 (N_11405,N_8024,N_9473);
nand U11406 (N_11406,N_5222,N_6703);
or U11407 (N_11407,N_6118,N_8751);
nand U11408 (N_11408,N_7187,N_7221);
or U11409 (N_11409,N_5437,N_5470);
nand U11410 (N_11410,N_6149,N_6123);
nand U11411 (N_11411,N_9490,N_6005);
nand U11412 (N_11412,N_8687,N_6810);
and U11413 (N_11413,N_5211,N_6992);
xnor U11414 (N_11414,N_8476,N_9478);
nand U11415 (N_11415,N_6167,N_8884);
nor U11416 (N_11416,N_5958,N_6935);
nor U11417 (N_11417,N_8480,N_9716);
xor U11418 (N_11418,N_8099,N_7522);
and U11419 (N_11419,N_7210,N_7954);
nand U11420 (N_11420,N_5506,N_7710);
nor U11421 (N_11421,N_7523,N_9111);
xnor U11422 (N_11422,N_5629,N_9212);
nand U11423 (N_11423,N_6211,N_9916);
and U11424 (N_11424,N_9773,N_5825);
nand U11425 (N_11425,N_9282,N_7876);
nor U11426 (N_11426,N_6661,N_6958);
nand U11427 (N_11427,N_5646,N_9457);
and U11428 (N_11428,N_7036,N_7222);
and U11429 (N_11429,N_8341,N_6668);
and U11430 (N_11430,N_7078,N_5481);
nand U11431 (N_11431,N_7468,N_9055);
nor U11432 (N_11432,N_7130,N_8865);
and U11433 (N_11433,N_6222,N_8738);
nor U11434 (N_11434,N_6408,N_8417);
nand U11435 (N_11435,N_6130,N_9053);
and U11436 (N_11436,N_7546,N_6627);
and U11437 (N_11437,N_5175,N_9347);
nor U11438 (N_11438,N_6471,N_8479);
nor U11439 (N_11439,N_5547,N_6733);
or U11440 (N_11440,N_7651,N_6200);
xnor U11441 (N_11441,N_6744,N_6838);
nand U11442 (N_11442,N_8526,N_6194);
nor U11443 (N_11443,N_7508,N_6525);
or U11444 (N_11444,N_8539,N_6041);
nor U11445 (N_11445,N_8256,N_8343);
nor U11446 (N_11446,N_9910,N_7079);
nand U11447 (N_11447,N_8714,N_7008);
xnor U11448 (N_11448,N_8569,N_7852);
nor U11449 (N_11449,N_5865,N_7454);
or U11450 (N_11450,N_5241,N_9499);
nor U11451 (N_11451,N_7254,N_9763);
and U11452 (N_11452,N_6012,N_8969);
and U11453 (N_11453,N_8182,N_6327);
nor U11454 (N_11454,N_5165,N_8981);
and U11455 (N_11455,N_5942,N_8281);
or U11456 (N_11456,N_7249,N_7703);
and U11457 (N_11457,N_7422,N_8075);
and U11458 (N_11458,N_8211,N_8168);
and U11459 (N_11459,N_8097,N_6724);
or U11460 (N_11460,N_8769,N_5634);
nand U11461 (N_11461,N_8621,N_5990);
nor U11462 (N_11462,N_7720,N_6610);
and U11463 (N_11463,N_8482,N_8815);
nor U11464 (N_11464,N_9298,N_7542);
and U11465 (N_11465,N_7336,N_7890);
xor U11466 (N_11466,N_9676,N_6604);
nand U11467 (N_11467,N_6566,N_8555);
xor U11468 (N_11468,N_7728,N_5109);
nand U11469 (N_11469,N_8894,N_5886);
or U11470 (N_11470,N_7577,N_5295);
nor U11471 (N_11471,N_5933,N_9709);
and U11472 (N_11472,N_9300,N_7156);
or U11473 (N_11473,N_6730,N_8966);
nor U11474 (N_11474,N_6679,N_6689);
and U11475 (N_11475,N_5687,N_6607);
nand U11476 (N_11476,N_6134,N_7914);
nor U11477 (N_11477,N_7371,N_8087);
or U11478 (N_11478,N_5820,N_8410);
and U11479 (N_11479,N_8533,N_5939);
nor U11480 (N_11480,N_5837,N_5571);
and U11481 (N_11481,N_7759,N_7228);
nand U11482 (N_11482,N_9801,N_9218);
nand U11483 (N_11483,N_5428,N_9908);
and U11484 (N_11484,N_6801,N_8140);
or U11485 (N_11485,N_8901,N_5307);
or U11486 (N_11486,N_9805,N_6241);
nor U11487 (N_11487,N_6413,N_6852);
and U11488 (N_11488,N_9524,N_8638);
and U11489 (N_11489,N_5529,N_6301);
and U11490 (N_11490,N_9932,N_6932);
nand U11491 (N_11491,N_7212,N_9705);
nor U11492 (N_11492,N_5281,N_8053);
and U11493 (N_11493,N_6203,N_9527);
or U11494 (N_11494,N_7165,N_6264);
and U11495 (N_11495,N_7153,N_9062);
nand U11496 (N_11496,N_5692,N_9415);
nand U11497 (N_11497,N_7947,N_6573);
nor U11498 (N_11498,N_8185,N_5293);
or U11499 (N_11499,N_6763,N_7432);
xnor U11500 (N_11500,N_7640,N_7263);
xor U11501 (N_11501,N_8797,N_9171);
nor U11502 (N_11502,N_8429,N_9039);
and U11503 (N_11503,N_6624,N_8765);
and U11504 (N_11504,N_6302,N_5821);
nor U11505 (N_11505,N_7983,N_7926);
or U11506 (N_11506,N_9201,N_6245);
xnor U11507 (N_11507,N_6831,N_5902);
or U11508 (N_11508,N_8677,N_9222);
xor U11509 (N_11509,N_5290,N_8418);
nand U11510 (N_11510,N_6294,N_6911);
or U11511 (N_11511,N_9198,N_8851);
or U11512 (N_11512,N_8366,N_8180);
nor U11513 (N_11513,N_6886,N_9563);
or U11514 (N_11514,N_9301,N_6486);
and U11515 (N_11515,N_9344,N_8136);
nand U11516 (N_11516,N_8205,N_7692);
and U11517 (N_11517,N_5294,N_9652);
or U11518 (N_11518,N_8231,N_9608);
and U11519 (N_11519,N_7389,N_6017);
or U11520 (N_11520,N_6696,N_7903);
nor U11521 (N_11521,N_6918,N_6584);
and U11522 (N_11522,N_9092,N_9173);
and U11523 (N_11523,N_7625,N_5633);
or U11524 (N_11524,N_9651,N_7346);
nor U11525 (N_11525,N_7798,N_8825);
nand U11526 (N_11526,N_8488,N_8369);
or U11527 (N_11527,N_6591,N_5096);
nor U11528 (N_11528,N_5480,N_9051);
or U11529 (N_11529,N_7891,N_5278);
and U11530 (N_11530,N_8540,N_7643);
and U11531 (N_11531,N_7838,N_7593);
nand U11532 (N_11532,N_5415,N_9013);
nor U11533 (N_11533,N_6155,N_8159);
or U11534 (N_11534,N_8193,N_9156);
xor U11535 (N_11535,N_5994,N_7383);
nor U11536 (N_11536,N_5508,N_9458);
xnor U11537 (N_11537,N_7248,N_6416);
or U11538 (N_11538,N_8454,N_5898);
or U11539 (N_11539,N_7068,N_6054);
nand U11540 (N_11540,N_5510,N_8077);
or U11541 (N_11541,N_6979,N_6410);
and U11542 (N_11542,N_9484,N_8987);
or U11543 (N_11543,N_6646,N_5569);
nor U11544 (N_11544,N_7033,N_5465);
nand U11545 (N_11545,N_9041,N_9789);
and U11546 (N_11546,N_8560,N_5640);
nor U11547 (N_11547,N_6344,N_9560);
and U11548 (N_11548,N_5405,N_6834);
and U11549 (N_11549,N_8826,N_7697);
and U11550 (N_11550,N_6157,N_5741);
xor U11551 (N_11551,N_8813,N_7905);
nor U11552 (N_11552,N_8712,N_6506);
nand U11553 (N_11553,N_7329,N_8006);
nor U11554 (N_11554,N_6009,N_8047);
and U11555 (N_11555,N_5803,N_8316);
nor U11556 (N_11556,N_5082,N_6329);
nand U11557 (N_11557,N_9782,N_5628);
nand U11558 (N_11558,N_5732,N_8995);
nand U11559 (N_11559,N_7098,N_8989);
nand U11560 (N_11560,N_5244,N_6721);
and U11561 (N_11561,N_8232,N_5234);
or U11562 (N_11562,N_6300,N_7711);
nand U11563 (N_11563,N_9451,N_6641);
nand U11564 (N_11564,N_9331,N_6583);
and U11565 (N_11565,N_7725,N_9430);
nand U11566 (N_11566,N_9371,N_5925);
nor U11567 (N_11567,N_5839,N_7596);
xnor U11568 (N_11568,N_8661,N_8634);
and U11569 (N_11569,N_5247,N_6457);
nand U11570 (N_11570,N_7590,N_8718);
nand U11571 (N_11571,N_8379,N_7355);
or U11572 (N_11572,N_9350,N_7421);
nand U11573 (N_11573,N_8487,N_8958);
nor U11574 (N_11574,N_8566,N_8315);
or U11575 (N_11575,N_6602,N_9422);
xor U11576 (N_11576,N_5444,N_8286);
xor U11577 (N_11577,N_7800,N_7707);
nand U11578 (N_11578,N_9200,N_9695);
nand U11579 (N_11579,N_5209,N_9007);
nand U11580 (N_11580,N_7502,N_8822);
or U11581 (N_11581,N_9585,N_8550);
nand U11582 (N_11582,N_8162,N_7186);
or U11583 (N_11583,N_6695,N_7816);
or U11584 (N_11584,N_8021,N_6432);
and U11585 (N_11585,N_9334,N_8448);
and U11586 (N_11586,N_8288,N_8272);
and U11587 (N_11587,N_6998,N_9780);
or U11588 (N_11588,N_9533,N_9732);
or U11589 (N_11589,N_6503,N_6387);
xnor U11590 (N_11590,N_9409,N_7671);
nand U11591 (N_11591,N_5612,N_7547);
nor U11592 (N_11592,N_8803,N_7289);
xnor U11593 (N_11593,N_8567,N_8469);
nand U11594 (N_11594,N_7449,N_6092);
and U11595 (N_11595,N_5435,N_5763);
and U11596 (N_11596,N_5802,N_5817);
nor U11597 (N_11597,N_8728,N_5742);
nand U11598 (N_11598,N_7748,N_5606);
or U11599 (N_11599,N_5252,N_7779);
nand U11600 (N_11600,N_7980,N_9100);
and U11601 (N_11601,N_8707,N_6908);
nand U11602 (N_11602,N_9203,N_6887);
xnor U11603 (N_11603,N_5636,N_5183);
nor U11604 (N_11604,N_5493,N_6440);
and U11605 (N_11605,N_6058,N_7241);
nand U11606 (N_11606,N_6281,N_8085);
and U11607 (N_11607,N_7188,N_6216);
nand U11608 (N_11608,N_9507,N_6448);
xnor U11609 (N_11609,N_6723,N_6818);
and U11610 (N_11610,N_6289,N_9870);
and U11611 (N_11611,N_5879,N_8112);
nand U11612 (N_11612,N_6117,N_5285);
or U11613 (N_11613,N_9727,N_8466);
nor U11614 (N_11614,N_7251,N_8200);
or U11615 (N_11615,N_6065,N_7428);
nor U11616 (N_11616,N_9311,N_6701);
nand U11617 (N_11617,N_8820,N_7672);
and U11618 (N_11618,N_5739,N_6571);
and U11619 (N_11619,N_8941,N_9921);
nand U11620 (N_11620,N_9832,N_8405);
and U11621 (N_11621,N_6109,N_5788);
nor U11622 (N_11622,N_9634,N_5427);
and U11623 (N_11623,N_8078,N_6906);
xnor U11624 (N_11624,N_5466,N_6350);
nor U11625 (N_11625,N_7069,N_5246);
or U11626 (N_11626,N_8397,N_5749);
or U11627 (N_11627,N_7287,N_8812);
nor U11628 (N_11628,N_5111,N_9260);
nand U11629 (N_11629,N_6418,N_7285);
nor U11630 (N_11630,N_5998,N_6907);
nor U11631 (N_11631,N_5885,N_7151);
nor U11632 (N_11632,N_9516,N_8922);
nand U11633 (N_11633,N_5489,N_6626);
xnor U11634 (N_11634,N_6892,N_6480);
nor U11635 (N_11635,N_6910,N_6612);
or U11636 (N_11636,N_9138,N_6875);
nor U11637 (N_11637,N_5433,N_5383);
xor U11638 (N_11638,N_5163,N_5113);
nand U11639 (N_11639,N_5343,N_7972);
nor U11640 (N_11640,N_7430,N_8984);
nor U11641 (N_11641,N_5422,N_6879);
nor U11642 (N_11642,N_6027,N_7243);
nand U11643 (N_11643,N_9065,N_6849);
nand U11644 (N_11644,N_6212,N_5826);
or U11645 (N_11645,N_9876,N_7267);
or U11646 (N_11646,N_6931,N_8603);
or U11647 (N_11647,N_6004,N_7834);
or U11648 (N_11648,N_7840,N_9169);
or U11649 (N_11649,N_8131,N_5212);
nand U11650 (N_11650,N_9068,N_6927);
nand U11651 (N_11651,N_7849,N_6000);
or U11652 (N_11652,N_8253,N_7705);
nand U11653 (N_11653,N_5718,N_5724);
nand U11654 (N_11654,N_8446,N_9711);
and U11655 (N_11655,N_5838,N_5577);
nand U11656 (N_11656,N_9158,N_7921);
nor U11657 (N_11657,N_5353,N_7323);
nand U11658 (N_11658,N_7721,N_7147);
nand U11659 (N_11659,N_8408,N_5325);
and U11660 (N_11660,N_5012,N_9059);
nand U11661 (N_11661,N_5852,N_6002);
or U11662 (N_11662,N_9378,N_9413);
xnor U11663 (N_11663,N_5641,N_7688);
nor U11664 (N_11664,N_7739,N_8157);
nand U11665 (N_11665,N_6460,N_8089);
xnor U11666 (N_11666,N_6359,N_8133);
and U11667 (N_11667,N_9669,N_5174);
xnor U11668 (N_11668,N_8326,N_7334);
xnor U11669 (N_11669,N_5254,N_6722);
xor U11670 (N_11670,N_8891,N_6678);
or U11671 (N_11671,N_6324,N_7343);
and U11672 (N_11672,N_8034,N_7361);
nand U11673 (N_11673,N_8399,N_5259);
and U11674 (N_11674,N_7296,N_5411);
nand U11675 (N_11675,N_5021,N_6097);
xnor U11676 (N_11676,N_5565,N_8044);
nor U11677 (N_11677,N_8390,N_7110);
or U11678 (N_11678,N_7535,N_5652);
nand U11679 (N_11679,N_9370,N_5771);
xor U11680 (N_11680,N_9214,N_8496);
xor U11681 (N_11681,N_7054,N_6404);
or U11682 (N_11682,N_7205,N_9197);
and U11683 (N_11683,N_5230,N_8207);
nand U11684 (N_11684,N_9044,N_9380);
nor U11685 (N_11685,N_9297,N_6228);
nand U11686 (N_11686,N_8467,N_8149);
and U11687 (N_11687,N_6700,N_7723);
or U11688 (N_11688,N_7237,N_8217);
and U11689 (N_11689,N_7208,N_9355);
and U11690 (N_11690,N_8086,N_7474);
and U11691 (N_11691,N_5737,N_7646);
nand U11692 (N_11692,N_6283,N_7946);
or U11693 (N_11693,N_8919,N_6268);
nor U11694 (N_11694,N_6651,N_9859);
xnor U11695 (N_11695,N_8117,N_6191);
and U11696 (N_11696,N_6120,N_8178);
or U11697 (N_11697,N_6093,N_8866);
nor U11698 (N_11698,N_6177,N_5631);
and U11699 (N_11699,N_7203,N_5728);
nor U11700 (N_11700,N_8003,N_7104);
nor U11701 (N_11701,N_5786,N_5268);
nor U11702 (N_11702,N_9995,N_5515);
nand U11703 (N_11703,N_7709,N_5223);
xnor U11704 (N_11704,N_9922,N_5372);
and U11705 (N_11705,N_9448,N_6962);
nor U11706 (N_11706,N_7563,N_7769);
and U11707 (N_11707,N_5332,N_9304);
nand U11708 (N_11708,N_7568,N_8606);
nor U11709 (N_11709,N_7017,N_9253);
nor U11710 (N_11710,N_5575,N_6311);
and U11711 (N_11711,N_7515,N_6789);
or U11712 (N_11712,N_7817,N_9199);
and U11713 (N_11713,N_7788,N_6738);
nor U11714 (N_11714,N_8979,N_5105);
nand U11715 (N_11715,N_5567,N_5698);
or U11716 (N_11716,N_6391,N_9574);
xnor U11717 (N_11717,N_7303,N_9944);
nand U11718 (N_11718,N_6101,N_6168);
nand U11719 (N_11719,N_8991,N_8623);
nand U11720 (N_11720,N_9432,N_9069);
and U11721 (N_11721,N_6605,N_5318);
nor U11722 (N_11722,N_7011,N_9453);
nand U11723 (N_11723,N_7319,N_7365);
and U11724 (N_11724,N_6258,N_5180);
or U11725 (N_11725,N_8105,N_9275);
or U11726 (N_11726,N_7482,N_8611);
nor U11727 (N_11727,N_6589,N_6698);
and U11728 (N_11728,N_8516,N_5809);
and U11729 (N_11729,N_7527,N_7324);
nor U11730 (N_11730,N_9935,N_6227);
nand U11731 (N_11731,N_8562,N_6213);
and U11732 (N_11732,N_7052,N_8925);
nand U11733 (N_11733,N_7458,N_7747);
and U11734 (N_11734,N_7382,N_6188);
or U11735 (N_11735,N_7557,N_5518);
xor U11736 (N_11736,N_6240,N_6606);
nor U11737 (N_11737,N_8433,N_5162);
xnor U11738 (N_11738,N_9662,N_8000);
and U11739 (N_11739,N_6765,N_5486);
and U11740 (N_11740,N_8747,N_8898);
nor U11741 (N_11741,N_8873,N_8963);
or U11742 (N_11742,N_9406,N_6729);
nand U11743 (N_11743,N_7272,N_6402);
and U11744 (N_11744,N_7266,N_7028);
nor U11745 (N_11745,N_5530,N_5570);
and U11746 (N_11746,N_8224,N_6107);
nor U11747 (N_11747,N_8398,N_9219);
nor U11748 (N_11748,N_9056,N_6740);
or U11749 (N_11749,N_8394,N_7486);
nor U11750 (N_11750,N_8313,N_6865);
nor U11751 (N_11751,N_8669,N_7714);
nand U11752 (N_11752,N_5917,N_8678);
or U11753 (N_11753,N_8314,N_9481);
nand U11754 (N_11754,N_8328,N_5966);
or U11755 (N_11755,N_8578,N_5928);
and U11756 (N_11756,N_8862,N_9743);
or U11757 (N_11757,N_5919,N_5721);
nand U11758 (N_11758,N_8524,N_8646);
xnor U11759 (N_11759,N_6928,N_8209);
and U11760 (N_11760,N_7067,N_9972);
or U11761 (N_11761,N_8528,N_8573);
or U11762 (N_11762,N_8734,N_7758);
and U11763 (N_11763,N_9245,N_8393);
or U11764 (N_11764,N_9631,N_9060);
nor U11765 (N_11765,N_8096,N_6776);
nor U11766 (N_11766,N_8102,N_7615);
nor U11767 (N_11767,N_9074,N_5190);
nor U11768 (N_11768,N_8449,N_7167);
or U11769 (N_11769,N_6816,N_6014);
and U11770 (N_11770,N_8094,N_9951);
and U11771 (N_11771,N_9251,N_7510);
and U11772 (N_11772,N_5814,N_5584);
xor U11773 (N_11773,N_8840,N_5594);
xor U11774 (N_11774,N_6593,N_7924);
nand U11775 (N_11775,N_7776,N_7207);
or U11776 (N_11776,N_9268,N_9020);
or U11777 (N_11777,N_7756,N_9774);
and U11778 (N_11778,N_8702,N_9483);
and U11779 (N_11779,N_9340,N_5166);
or U11780 (N_11780,N_5309,N_9990);
and U11781 (N_11781,N_7125,N_6304);
and U11782 (N_11782,N_9837,N_8227);
or U11783 (N_11783,N_9901,N_5609);
nand U11784 (N_11784,N_7878,N_9116);
and U11785 (N_11785,N_9023,N_9750);
and U11786 (N_11786,N_6622,N_5643);
nor U11787 (N_11787,N_6474,N_8147);
and U11788 (N_11788,N_7712,N_7953);
or U11789 (N_11789,N_8867,N_9390);
xor U11790 (N_11790,N_9170,N_7386);
or U11791 (N_11791,N_6973,N_7699);
and U11792 (N_11792,N_7521,N_9867);
and U11793 (N_11793,N_6265,N_5218);
nand U11794 (N_11794,N_8298,N_9924);
nand U11795 (N_11795,N_9015,N_6981);
and U11796 (N_11796,N_8602,N_7907);
nor U11797 (N_11797,N_6208,N_5250);
xor U11798 (N_11798,N_6150,N_7685);
nand U11799 (N_11799,N_6116,N_8145);
or U11800 (N_11800,N_7831,N_7958);
nor U11801 (N_11801,N_7322,N_7786);
and U11802 (N_11802,N_6290,N_8960);
or U11803 (N_11803,N_9362,N_7620);
or U11804 (N_11804,N_7388,N_6726);
nand U11805 (N_11805,N_5310,N_9429);
and U11806 (N_11806,N_9688,N_8972);
xor U11807 (N_11807,N_8269,N_7635);
xor U11808 (N_11808,N_6201,N_9313);
xor U11809 (N_11809,N_6328,N_5159);
nand U11810 (N_11810,N_8019,N_9153);
and U11811 (N_11811,N_9318,N_5439);
and U11812 (N_11812,N_5717,N_5669);
nor U11813 (N_11813,N_9446,N_9159);
or U11814 (N_11814,N_9353,N_7066);
nand U11815 (N_11815,N_5873,N_6160);
xor U11816 (N_11816,N_8807,N_5720);
nor U11817 (N_11817,N_9042,N_5059);
or U11818 (N_11818,N_9435,N_5157);
nand U11819 (N_11819,N_8587,N_9671);
or U11820 (N_11820,N_5729,N_7809);
or U11821 (N_11821,N_8230,N_6654);
xnor U11822 (N_11822,N_9577,N_7292);
and U11823 (N_11823,N_7470,N_8801);
nor U11824 (N_11824,N_7121,N_5831);
nand U11825 (N_11825,N_9587,N_5689);
nand U11826 (N_11826,N_8856,N_5037);
nand U11827 (N_11827,N_8370,N_7400);
xor U11828 (N_11828,N_6968,N_5123);
or U11829 (N_11829,N_5171,N_5719);
nand U11830 (N_11830,N_8929,N_9657);
or U11831 (N_11831,N_5955,N_8684);
nor U11832 (N_11832,N_8383,N_9647);
or U11833 (N_11833,N_7282,N_7966);
nor U11834 (N_11834,N_5866,N_5696);
nand U11835 (N_11835,N_8330,N_6934);
or U11836 (N_11836,N_8954,N_6768);
nand U11837 (N_11837,N_5315,N_5956);
or U11838 (N_11838,N_6018,N_5213);
nand U11839 (N_11839,N_9693,N_6686);
nand U11840 (N_11840,N_9000,N_9896);
and U11841 (N_11841,N_8762,N_6396);
nand U11842 (N_11842,N_6185,N_5487);
nand U11843 (N_11843,N_6532,N_7412);
or U11844 (N_11844,N_8659,N_5388);
nand U11845 (N_11845,N_9642,N_6490);
nor U11846 (N_11846,N_6383,N_5147);
nor U11847 (N_11847,N_9997,N_8680);
and U11848 (N_11848,N_5555,N_7485);
or U11849 (N_11849,N_5767,N_6083);
nand U11850 (N_11850,N_7949,N_8522);
or U11851 (N_11851,N_6623,N_7812);
or U11852 (N_11852,N_5359,N_9678);
nand U11853 (N_11853,N_7362,N_6133);
nor U11854 (N_11854,N_6630,N_8058);
nand U11855 (N_11855,N_7694,N_6504);
and U11856 (N_11856,N_6215,N_7152);
and U11857 (N_11857,N_7000,N_5429);
nor U11858 (N_11858,N_8265,N_9425);
or U11859 (N_11859,N_6670,N_6717);
and U11860 (N_11860,N_5700,N_5620);
nand U11861 (N_11861,N_6087,N_8509);
or U11862 (N_11862,N_8171,N_5233);
nand U11863 (N_11863,N_6819,N_5762);
nor U11864 (N_11864,N_5492,N_9879);
nor U11865 (N_11865,N_9263,N_9697);
or U11866 (N_11866,N_5849,N_5857);
nand U11867 (N_11867,N_9147,N_6769);
nor U11868 (N_11868,N_5685,N_7010);
xor U11869 (N_11869,N_6113,N_8713);
or U11870 (N_11870,N_9098,N_9192);
nand U11871 (N_11871,N_8641,N_6426);
or U11872 (N_11872,N_7766,N_7802);
and U11873 (N_11873,N_8639,N_8444);
nand U11874 (N_11874,N_8014,N_6792);
nor U11875 (N_11875,N_9142,N_6790);
nor U11876 (N_11876,N_9503,N_9273);
nor U11877 (N_11877,N_9468,N_7655);
or U11878 (N_11878,N_7886,N_9530);
nor U11879 (N_11879,N_6509,N_5413);
nor U11880 (N_11880,N_7845,N_9623);
xor U11881 (N_11881,N_5659,N_5120);
xnor U11882 (N_11882,N_9420,N_9847);
nand U11883 (N_11883,N_9757,N_5408);
nor U11884 (N_11884,N_6479,N_9655);
and U11885 (N_11885,N_8011,N_8470);
nand U11886 (N_11886,N_9914,N_5524);
and U11887 (N_11887,N_6444,N_8852);
or U11888 (N_11888,N_9994,N_6570);
and U11889 (N_11889,N_7575,N_8909);
nand U11890 (N_11890,N_8371,N_5630);
and U11891 (N_11891,N_6234,N_8693);
nand U11892 (N_11892,N_6613,N_7994);
or U11893 (N_11893,N_5625,N_8949);
nand U11894 (N_11894,N_8331,N_5654);
nor U11895 (N_11895,N_5275,N_9902);
nor U11896 (N_11896,N_9234,N_9134);
and U11897 (N_11897,N_8338,N_8594);
and U11898 (N_11898,N_6926,N_9754);
and U11899 (N_11899,N_7313,N_8582);
and U11900 (N_11900,N_8875,N_6975);
or U11901 (N_11901,N_6964,N_6619);
or U11902 (N_11902,N_8615,N_5532);
nor U11903 (N_11903,N_6616,N_5085);
and U11904 (N_11904,N_9841,N_9749);
nand U11905 (N_11905,N_7524,N_5554);
nor U11906 (N_11906,N_6767,N_7843);
xor U11907 (N_11907,N_5764,N_6043);
and U11908 (N_11908,N_6376,N_8005);
nand U11909 (N_11909,N_6367,N_6951);
or U11910 (N_11910,N_5064,N_9653);
nand U11911 (N_11911,N_6737,N_6939);
or U11912 (N_11912,N_7378,N_7965);
or U11913 (N_11913,N_5815,N_9233);
and U11914 (N_11914,N_8016,N_6851);
xnor U11915 (N_11915,N_5047,N_9404);
and U11916 (N_11916,N_8106,N_9450);
xnor U11917 (N_11917,N_6260,N_5758);
nand U11918 (N_11918,N_6692,N_6688);
nor U11919 (N_11919,N_8595,N_8353);
or U11920 (N_11920,N_7479,N_5340);
and U11921 (N_11921,N_6850,N_6434);
nor U11922 (N_11922,N_7666,N_7347);
and U11923 (N_11923,N_5461,N_6142);
or U11924 (N_11924,N_9954,N_6338);
or U11925 (N_11925,N_6285,N_8763);
nor U11926 (N_11926,N_7085,N_7638);
nand U11927 (N_11927,N_9660,N_8947);
or U11928 (N_11928,N_8165,N_9460);
nand U11929 (N_11929,N_5708,N_9696);
nand U11930 (N_11930,N_8768,N_5226);
nor U11931 (N_11931,N_5924,N_8378);
xnor U11932 (N_11932,N_9904,N_8279);
nand U11933 (N_11933,N_7981,N_6572);
and U11934 (N_11934,N_7105,N_5497);
or U11935 (N_11935,N_5774,N_7990);
or U11936 (N_11936,N_8151,N_8070);
or U11937 (N_11937,N_9204,N_7209);
nor U11938 (N_11938,N_5126,N_9580);
nand U11939 (N_11939,N_5864,N_7159);
nor U11940 (N_11940,N_7261,N_5707);
and U11941 (N_11941,N_9745,N_5051);
nand U11942 (N_11942,N_6588,N_5656);
nand U11943 (N_11943,N_8905,N_9485);
and U11944 (N_11944,N_9249,N_6603);
and U11945 (N_11945,N_8115,N_7200);
nand U11946 (N_11946,N_7626,N_7740);
and U11947 (N_11947,N_9708,N_5283);
nand U11948 (N_11948,N_7122,N_8946);
or U11949 (N_11949,N_7767,N_8940);
or U11950 (N_11950,N_9135,N_8468);
and U11951 (N_11951,N_9872,N_6422);
nor U11952 (N_11952,N_7120,N_7743);
and U11953 (N_11953,N_6299,N_5195);
xnor U11954 (N_11954,N_9920,N_8689);
or U11955 (N_11955,N_7604,N_6409);
nor U11956 (N_11956,N_5355,N_7829);
or U11957 (N_11957,N_5835,N_8190);
xor U11958 (N_11958,N_7653,N_7944);
xnor U11959 (N_11959,N_8786,N_6751);
nand U11960 (N_11960,N_8710,N_9936);
nor U11961 (N_11961,N_9106,N_7978);
xnor U11962 (N_11962,N_9787,N_6590);
or U11963 (N_11963,N_6136,N_6140);
or U11964 (N_11964,N_6807,N_8549);
or U11965 (N_11965,N_6135,N_6893);
nand U11966 (N_11966,N_7090,N_9004);
xor U11967 (N_11967,N_6279,N_8913);
nor U11968 (N_11968,N_5715,N_6625);
nor U11969 (N_11969,N_6750,N_9210);
and U11970 (N_11970,N_5078,N_6070);
and U11971 (N_11971,N_8135,N_6902);
and U11972 (N_11972,N_6049,N_9034);
and U11973 (N_11973,N_8204,N_8642);
and U11974 (N_11974,N_8007,N_7256);
and U11975 (N_11975,N_6697,N_8975);
nor U11976 (N_11976,N_6766,N_9439);
xnor U11977 (N_11977,N_7158,N_5670);
nand U11978 (N_11978,N_7904,N_6956);
and U11979 (N_11979,N_8796,N_5308);
or U11980 (N_11980,N_5133,N_6339);
nand U11981 (N_11981,N_9024,N_6761);
nor U11982 (N_11982,N_9547,N_7566);
and U11983 (N_11983,N_5830,N_8619);
and U11984 (N_11984,N_9352,N_6316);
and U11985 (N_11985,N_8188,N_5794);
and U11986 (N_11986,N_9394,N_6742);
and U11987 (N_11987,N_9964,N_7260);
nor U11988 (N_11988,N_9960,N_9569);
nor U11989 (N_11989,N_5514,N_5727);
nor U11990 (N_11990,N_7172,N_8921);
nand U11991 (N_11991,N_7439,N_6720);
nand U11992 (N_11992,N_7783,N_5348);
and U11993 (N_11993,N_5906,N_7922);
nor U11994 (N_11994,N_8100,N_6899);
xor U11995 (N_11995,N_8195,N_9967);
nor U11996 (N_11996,N_8918,N_7494);
or U11997 (N_11997,N_8271,N_7814);
and U11998 (N_11998,N_8067,N_6385);
nor U11999 (N_11999,N_6500,N_9105);
nor U12000 (N_12000,N_8156,N_9292);
nor U12001 (N_12001,N_9332,N_7668);
nand U12002 (N_12002,N_9395,N_9752);
and U12003 (N_12003,N_9248,N_9531);
or U12004 (N_12004,N_9570,N_5148);
nand U12005 (N_12005,N_7427,N_8790);
or U12006 (N_12006,N_6539,N_7589);
nand U12007 (N_12007,N_7715,N_8817);
nor U12008 (N_12008,N_5748,N_9075);
and U12009 (N_12009,N_9143,N_8868);
nor U12010 (N_12010,N_9665,N_7562);
and U12011 (N_12011,N_9307,N_7465);
xnor U12012 (N_12012,N_8126,N_9258);
xor U12013 (N_12013,N_9970,N_6266);
nand U12014 (N_12014,N_5202,N_6752);
nand U12015 (N_12015,N_7561,N_7271);
nor U12016 (N_12016,N_8932,N_9414);
and U12017 (N_12017,N_9591,N_8273);
and U12018 (N_12018,N_6930,N_5255);
nand U12019 (N_12019,N_8737,N_6904);
nand U12020 (N_12020,N_6781,N_6347);
or U12021 (N_12021,N_7823,N_5416);
nor U12022 (N_12022,N_6246,N_8698);
nand U12023 (N_12023,N_7632,N_9265);
and U12024 (N_12024,N_9889,N_8333);
nand U12025 (N_12025,N_5228,N_7442);
or U12026 (N_12026,N_6179,N_6407);
nand U12027 (N_12027,N_6321,N_5397);
nor U12028 (N_12028,N_7810,N_9656);
xnor U12029 (N_12029,N_9160,N_8874);
nand U12030 (N_12030,N_6153,N_8439);
nand U12031 (N_12031,N_9618,N_5876);
nor U12032 (N_12032,N_9025,N_7937);
nand U12033 (N_12033,N_9177,N_5754);
nor U12034 (N_12034,N_8203,N_6253);
nor U12035 (N_12035,N_5598,N_9235);
xnor U12036 (N_12036,N_5674,N_7528);
or U12037 (N_12037,N_8048,N_6186);
nand U12038 (N_12038,N_8186,N_8802);
nor U12039 (N_12039,N_7142,N_5251);
xnor U12040 (N_12040,N_8377,N_7348);
or U12041 (N_12041,N_5003,N_8022);
nand U12042 (N_12042,N_9823,N_8161);
nor U12043 (N_12043,N_5909,N_8285);
and U12044 (N_12044,N_7851,N_7541);
and U12045 (N_12045,N_6386,N_5768);
and U12046 (N_12046,N_8283,N_8730);
xor U12047 (N_12047,N_5745,N_5695);
xor U12048 (N_12048,N_8654,N_6269);
or U12049 (N_12049,N_9956,N_9221);
nor U12050 (N_12050,N_9032,N_6341);
and U12051 (N_12051,N_7864,N_7644);
nor U12052 (N_12052,N_7900,N_6708);
nand U12053 (N_12053,N_6377,N_8268);
or U12054 (N_12054,N_6600,N_6020);
nand U12055 (N_12055,N_6812,N_9463);
and U12056 (N_12056,N_5927,N_5131);
or U12057 (N_12057,N_9494,N_5895);
nor U12058 (N_12058,N_6577,N_9940);
nand U12059 (N_12059,N_7393,N_9739);
or U12060 (N_12060,N_7047,N_6901);
nor U12061 (N_12061,N_7955,N_9321);
nor U12062 (N_12062,N_7724,N_6891);
nand U12063 (N_12063,N_5949,N_8532);
or U12064 (N_12064,N_9567,N_6983);
and U12065 (N_12065,N_7433,N_6863);
and U12066 (N_12066,N_7276,N_7333);
and U12067 (N_12067,N_6780,N_7174);
and U12068 (N_12068,N_8064,N_5449);
nor U12069 (N_12069,N_7320,N_8636);
nand U12070 (N_12070,N_5360,N_9293);
nor U12071 (N_12071,N_6502,N_8724);
and U12072 (N_12072,N_7579,N_8780);
nand U12073 (N_12073,N_8556,N_7236);
or U12074 (N_12074,N_9261,N_7973);
and U12075 (N_12075,N_5011,N_8453);
or U12076 (N_12076,N_8432,N_9326);
nand U12077 (N_12077,N_7445,N_5910);
and U12078 (N_12078,N_8208,N_6673);
nand U12079 (N_12079,N_9686,N_7602);
nor U12080 (N_12080,N_8916,N_9319);
nand U12081 (N_12081,N_8924,N_6286);
nand U12082 (N_12082,N_9658,N_7202);
or U12083 (N_12083,N_7327,N_6756);
and U12084 (N_12084,N_5583,N_8557);
nand U12085 (N_12085,N_9625,N_9014);
xnor U12086 (N_12086,N_6207,N_7559);
nand U12087 (N_12087,N_9728,N_5114);
or U12088 (N_12088,N_9869,N_7345);
nand U12089 (N_12089,N_5787,N_7179);
and U12090 (N_12090,N_8834,N_9985);
nor U12091 (N_12091,N_9873,N_9637);
and U12092 (N_12092,N_7418,N_8721);
xor U12093 (N_12093,N_6820,N_5029);
and U12094 (N_12094,N_9517,N_7827);
and U12095 (N_12095,N_9418,N_6210);
nand U12096 (N_12096,N_6980,N_8523);
and U12097 (N_12097,N_5661,N_8008);
nor U12098 (N_12098,N_5288,N_8571);
nand U12099 (N_12099,N_7357,N_7901);
or U12100 (N_12100,N_6204,N_7072);
and U12101 (N_12101,N_7469,N_7022);
or U12102 (N_12102,N_6069,N_5188);
and U12103 (N_12103,N_9857,N_9342);
or U12104 (N_12104,N_9072,N_5682);
and U12105 (N_12105,N_7792,N_7004);
and U12106 (N_12106,N_6741,N_6047);
nor U12107 (N_12107,N_7956,N_7024);
nor U12108 (N_12108,N_9520,N_5963);
xnor U12109 (N_12109,N_5110,N_7306);
and U12110 (N_12110,N_7399,N_6828);
nor U12111 (N_12111,N_7945,N_7782);
nand U12112 (N_12112,N_6905,N_5038);
or U12113 (N_12113,N_5503,N_8994);
nor U12114 (N_12114,N_8686,N_7722);
nand U12115 (N_12115,N_9947,N_9534);
nand U12116 (N_12116,N_8173,N_8241);
and U12117 (N_12117,N_6745,N_7674);
or U12118 (N_12118,N_7506,N_7657);
nor U12119 (N_12119,N_5169,N_7311);
xor U12120 (N_12120,N_7588,N_9250);
and U12121 (N_12121,N_8938,N_7214);
nand U12122 (N_12122,N_5447,N_8303);
and U12123 (N_12123,N_5496,N_5265);
nor U12124 (N_12124,N_8758,N_9475);
and U12125 (N_12125,N_5604,N_5912);
nand U12126 (N_12126,N_7986,N_8304);
or U12127 (N_12127,N_9437,N_9819);
nand U12128 (N_12128,N_5094,N_6978);
nand U12129 (N_12129,N_7601,N_7126);
nor U12130 (N_12130,N_7826,N_5263);
nor U12131 (N_12131,N_8356,N_9729);
nor U12132 (N_12132,N_8709,N_7376);
and U12133 (N_12133,N_8238,N_7850);
or U12134 (N_12134,N_5092,N_6151);
xor U12135 (N_12135,N_7716,N_5221);
and U12136 (N_12136,N_9048,N_5509);
nand U12137 (N_12137,N_5297,N_9894);
nand U12138 (N_12138,N_9087,N_6462);
nand U12139 (N_12139,N_5155,N_6965);
and U12140 (N_12140,N_7234,N_9548);
and U12141 (N_12141,N_9269,N_9247);
or U12142 (N_12142,N_9474,N_9129);
nor U12143 (N_12143,N_9974,N_5485);
nor U12144 (N_12144,N_8517,N_9447);
or U12145 (N_12145,N_5373,N_6355);
xor U12146 (N_12146,N_6841,N_9506);
and U12147 (N_12147,N_8726,N_9899);
nand U12148 (N_12148,N_9624,N_9667);
nor U12149 (N_12149,N_5657,N_7466);
and U12150 (N_12150,N_9266,N_6096);
and U12151 (N_12151,N_5469,N_6957);
xor U12152 (N_12152,N_8999,N_5286);
xor U12153 (N_12153,N_5017,N_6877);
nor U12154 (N_12154,N_6990,N_5677);
nand U12155 (N_12155,N_9028,N_7731);
or U12156 (N_12156,N_9573,N_9125);
nand U12157 (N_12157,N_9154,N_9887);
or U12158 (N_12158,N_9322,N_8881);
nand U12159 (N_12159,N_7414,N_7962);
xnor U12160 (N_12160,N_7183,N_8906);
and U12161 (N_12161,N_8361,N_5970);
nand U12162 (N_12162,N_9706,N_9640);
nand U12163 (N_12163,N_8400,N_6229);
nand U12164 (N_12164,N_9854,N_8155);
nor U12165 (N_12165,N_9021,N_9480);
nor U12166 (N_12166,N_8515,N_5627);
and U12167 (N_12167,N_5269,N_8593);
nand U12168 (N_12168,N_7858,N_7919);
and U12169 (N_12169,N_8869,N_7686);
or U12170 (N_12170,N_9556,N_6196);
xor U12171 (N_12171,N_7084,N_6079);
or U12172 (N_12172,N_5142,N_9211);
and U12173 (N_12173,N_7572,N_8065);
nand U12174 (N_12174,N_9796,N_8511);
or U12175 (N_12175,N_6531,N_9612);
and U12176 (N_12176,N_9330,N_8497);
nor U12177 (N_12177,N_7128,N_5676);
xnor U12178 (N_12178,N_7732,N_7097);
xnor U12179 (N_12179,N_9528,N_9858);
nor U12180 (N_12180,N_6121,N_9270);
nand U12181 (N_12181,N_9379,N_8017);
or U12182 (N_12182,N_6909,N_8491);
xor U12183 (N_12183,N_5887,N_6141);
nand U12184 (N_12184,N_8477,N_9781);
and U12185 (N_12185,N_7794,N_5557);
xnor U12186 (N_12186,N_7993,N_7293);
nor U12187 (N_12187,N_7461,N_6749);
and U12188 (N_12188,N_5441,N_6470);
nand U12189 (N_12189,N_5119,N_6585);
or U12190 (N_12190,N_8794,N_9926);
and U12191 (N_12191,N_6664,N_7933);
or U12192 (N_12192,N_5035,N_7211);
nand U12193 (N_12193,N_5649,N_6595);
nor U12194 (N_12194,N_9950,N_5245);
nand U12195 (N_12195,N_8633,N_8348);
or U12196 (N_12196,N_6955,N_8777);
and U12197 (N_12197,N_6883,N_7979);
or U12198 (N_12198,N_7332,N_8407);
nor U12199 (N_12199,N_9845,N_8312);
nor U12200 (N_12200,N_6411,N_8942);
and U12201 (N_12201,N_6546,N_6056);
nand U12202 (N_12202,N_6821,N_6036);
or U12203 (N_12203,N_6782,N_6735);
or U12204 (N_12204,N_6483,N_7310);
nor U12205 (N_12205,N_8129,N_5501);
nand U12206 (N_12206,N_9257,N_7478);
nor U12207 (N_12207,N_5951,N_6365);
and U12208 (N_12208,N_5892,N_9188);
nand U12209 (N_12209,N_5600,N_9514);
nand U12210 (N_12210,N_6205,N_5196);
or U12211 (N_12211,N_6442,N_8552);
nor U12212 (N_12212,N_9228,N_5192);
or U12213 (N_12213,N_9365,N_5301);
and U12214 (N_12214,N_8036,N_5326);
or U12215 (N_12215,N_6859,N_9172);
nand U12216 (N_12216,N_5146,N_6023);
or U12217 (N_12217,N_8218,N_5614);
or U12218 (N_12218,N_6823,N_5744);
and U12219 (N_12219,N_6527,N_8563);
or U12220 (N_12220,N_8872,N_7553);
and U12221 (N_12221,N_7144,N_8846);
or U12222 (N_12222,N_9937,N_5215);
nor U12223 (N_12223,N_5699,N_5328);
nor U12224 (N_12224,N_9097,N_5095);
nor U12225 (N_12225,N_6103,N_9104);
or U12226 (N_12226,N_5938,N_7192);
nor U12227 (N_12227,N_5031,N_9650);
or U12228 (N_12228,N_9462,N_9638);
nand U12229 (N_12229,N_9903,N_5333);
or U12230 (N_12230,N_6366,N_9836);
and U12231 (N_12231,N_6423,N_7961);
xnor U12232 (N_12232,N_7250,N_6015);
xor U12233 (N_12233,N_7434,N_8172);
and U12234 (N_12234,N_9193,N_9734);
nand U12235 (N_12235,N_6873,N_5704);
or U12236 (N_12236,N_9291,N_6676);
or U12237 (N_12237,N_7305,N_5504);
nor U12238 (N_12238,N_7294,N_6345);
xor U12239 (N_12239,N_8247,N_6472);
or U12240 (N_12240,N_9740,N_7095);
nor U12241 (N_12241,N_8591,N_6419);
nand U12242 (N_12242,N_9707,N_8169);
xor U12243 (N_12243,N_5015,N_7764);
or U12244 (N_12244,N_7597,N_8725);
xnor U12245 (N_12245,N_8518,N_9701);
nor U12246 (N_12246,N_6482,N_7706);
or U12247 (N_12247,N_8584,N_6576);
nor U12248 (N_12248,N_9784,N_7727);
or U12249 (N_12249,N_8798,N_6003);
or U12250 (N_12250,N_5189,N_9552);
xor U12251 (N_12251,N_5490,N_7218);
nand U12252 (N_12252,N_5991,N_8255);
or U12253 (N_12253,N_8009,N_8050);
nand U12254 (N_12254,N_7370,N_5621);
and U12255 (N_12255,N_9388,N_8118);
nand U12256 (N_12256,N_5443,N_6870);
or U12257 (N_12257,N_5996,N_8760);
and U12258 (N_12258,N_5897,N_9794);
or U12259 (N_12259,N_9440,N_7663);
and U12260 (N_12260,N_8076,N_5468);
xor U12261 (N_12261,N_7226,N_9674);
and U12262 (N_12262,N_5488,N_8483);
xnor U12263 (N_12263,N_6569,N_9512);
or U12264 (N_12264,N_5371,N_8928);
nor U12265 (N_12265,N_7230,N_6541);
or U12266 (N_12266,N_5705,N_7264);
or U12267 (N_12267,N_5323,N_7255);
nand U12268 (N_12268,N_6074,N_6274);
nand U12269 (N_12269,N_8694,N_5962);
or U12270 (N_12270,N_5548,N_6574);
or U12271 (N_12271,N_8653,N_8904);
nor U12272 (N_12272,N_6933,N_6351);
nand U12273 (N_12273,N_6811,N_9783);
nor U12274 (N_12274,N_9202,N_8711);
xor U12275 (N_12275,N_8785,N_5666);
nor U12276 (N_12276,N_5525,N_8828);
nor U12277 (N_12277,N_9566,N_6669);
nand U12278 (N_12278,N_8732,N_6013);
nor U12279 (N_12279,N_8647,N_8605);
or U12280 (N_12280,N_6146,N_6110);
or U12281 (N_12281,N_7754,N_7402);
and U12282 (N_12282,N_6441,N_5932);
or U12283 (N_12283,N_8436,N_5553);
xnor U12284 (N_12284,N_8223,N_6401);
nor U12285 (N_12285,N_5071,N_6860);
or U12286 (N_12286,N_8354,N_8985);
nor U12287 (N_12287,N_8700,N_9768);
xnor U12288 (N_12288,N_5448,N_5808);
nand U12289 (N_12289,N_9538,N_5499);
nand U12290 (N_12290,N_7198,N_6496);
nor U12291 (N_12291,N_7839,N_5452);
nor U12292 (N_12292,N_9283,N_7998);
nand U12293 (N_12293,N_5613,N_8503);
nand U12294 (N_12294,N_6278,N_8823);
or U12295 (N_12295,N_8501,N_6652);
and U12296 (N_12296,N_6995,N_9953);
and U12297 (N_12297,N_5982,N_7708);
nand U12298 (N_12298,N_9737,N_9930);
nand U12299 (N_12299,N_6425,N_6895);
xnor U12300 (N_12300,N_5730,N_6601);
nand U12301 (N_12301,N_9442,N_8930);
nand U12302 (N_12302,N_9938,N_8293);
xor U12303 (N_12303,N_5005,N_6296);
or U12304 (N_12304,N_9626,N_9401);
nand U12305 (N_12305,N_5757,N_6683);
xor U12306 (N_12306,N_5026,N_6492);
or U12307 (N_12307,N_7045,N_7997);
nand U12308 (N_12308,N_5106,N_5170);
nor U12309 (N_12309,N_9818,N_6649);
nand U12310 (N_12310,N_9590,N_8324);
nand U12311 (N_12311,N_5460,N_6833);
nor U12312 (N_12312,N_6677,N_7496);
and U12313 (N_12313,N_6946,N_9417);
nor U12314 (N_12314,N_8494,N_5650);
nor U12315 (N_12315,N_9996,N_5149);
and U12316 (N_12316,N_9989,N_5249);
nand U12317 (N_12317,N_5161,N_6985);
xnor U12318 (N_12318,N_5046,N_5121);
nand U12319 (N_12319,N_6108,N_5915);
nand U12320 (N_12320,N_5217,N_7733);
and U12321 (N_12321,N_6061,N_7488);
nor U12322 (N_12322,N_9722,N_5117);
nor U12323 (N_12323,N_7181,N_5053);
nor U12324 (N_12324,N_8327,N_5090);
and U12325 (N_12325,N_7075,N_7118);
and U12326 (N_12326,N_8039,N_8141);
or U12327 (N_12327,N_6270,N_9385);
nor U12328 (N_12328,N_6707,N_6705);
xnor U12329 (N_12329,N_5304,N_5807);
nor U12330 (N_12330,N_6959,N_6843);
nand U12331 (N_12331,N_6399,N_5829);
and U12332 (N_12332,N_5861,N_5370);
nor U12333 (N_12333,N_7145,N_5135);
and U12334 (N_12334,N_6552,N_6829);
nand U12335 (N_12335,N_7860,N_8276);
and U12336 (N_12336,N_6748,N_5066);
or U12337 (N_12337,N_9229,N_5389);
nor U12338 (N_12338,N_8069,N_8043);
nand U12339 (N_12339,N_8249,N_6547);
and U12340 (N_12340,N_9892,N_5138);
and U12341 (N_12341,N_7881,N_8977);
or U12342 (N_12342,N_8214,N_7867);
nand U12343 (N_12343,N_5568,N_7606);
and U12344 (N_12344,N_8519,N_9314);
or U12345 (N_12345,N_8599,N_7116);
or U12346 (N_12346,N_6743,N_7253);
nand U12347 (N_12347,N_8620,N_9542);
nor U12348 (N_12348,N_8529,N_5350);
nand U12349 (N_12349,N_9786,N_5800);
xor U12350 (N_12350,N_9349,N_9303);
nor U12351 (N_12351,N_6779,N_8848);
nor U12352 (N_12352,N_9753,N_8424);
and U12353 (N_12353,N_5889,N_6611);
nor U12354 (N_12354,N_6421,N_8559);
nand U12355 (N_12355,N_8251,N_9855);
nand U12356 (N_12356,N_5810,N_8351);
nor U12357 (N_12357,N_6271,N_7417);
xnor U12358 (N_12358,N_8451,N_7034);
nand U12359 (N_12359,N_5321,N_7379);
nor U12360 (N_12360,N_5208,N_6051);
or U12361 (N_12361,N_7525,N_8534);
nand U12362 (N_12362,N_5535,N_5667);
or U12363 (N_12363,N_9767,N_6042);
and U12364 (N_12364,N_5858,N_9115);
xnor U12365 (N_12365,N_9176,N_7795);
and U12366 (N_12366,N_9639,N_9860);
nand U12367 (N_12367,N_7013,N_5018);
and U12368 (N_12368,N_7974,N_6924);
xor U12369 (N_12369,N_9089,N_9057);
or U12370 (N_12370,N_8993,N_9047);
and U12371 (N_12371,N_5968,N_8804);
or U12372 (N_12372,N_9545,N_7511);
xnor U12373 (N_12373,N_8134,N_7001);
or U12374 (N_12374,N_6778,N_9982);
nor U12375 (N_12375,N_7335,N_7505);
and U12376 (N_12376,N_6871,N_6952);
or U12377 (N_12377,N_7259,N_6888);
and U12378 (N_12378,N_5472,N_7341);
or U12379 (N_12379,N_7038,N_9348);
nor U12380 (N_12380,N_5167,N_8887);
nor U12381 (N_12381,N_5273,N_9621);
nand U12382 (N_12382,N_7025,N_8609);
and U12383 (N_12383,N_9868,N_9829);
nor U12384 (N_12384,N_9110,N_8148);
xor U12385 (N_12385,N_5396,N_5044);
nand U12386 (N_12386,N_5601,N_8900);
nand U12387 (N_12387,N_9381,N_8821);
and U12388 (N_12388,N_8461,N_6596);
or U12389 (N_12389,N_8811,N_5062);
and U12390 (N_12390,N_7793,N_7302);
nor U12391 (N_12391,N_7569,N_5088);
nor U12392 (N_12392,N_7719,N_8998);
nand U12393 (N_12393,N_6040,N_7871);
or U12394 (N_12394,N_9043,N_5591);
or U12395 (N_12395,N_8244,N_9828);
nor U12396 (N_12396,N_5341,N_9259);
nand U12397 (N_12397,N_7658,N_7101);
nand U12398 (N_12398,N_8199,N_6293);
xnor U12399 (N_12399,N_5298,N_8907);
or U12400 (N_12400,N_9005,N_8352);
or U12401 (N_12401,N_9791,N_6971);
or U12402 (N_12402,N_5240,N_9992);
or U12403 (N_12403,N_8576,N_6334);
nand U12404 (N_12404,N_8174,N_5681);
and U12405 (N_12405,N_9721,N_5160);
nand U12406 (N_12406,N_8001,N_9256);
nor U12407 (N_12407,N_5314,N_8319);
or U12408 (N_12408,N_6297,N_6505);
and U12409 (N_12409,N_8183,N_9692);
xnor U12410 (N_12410,N_7676,N_7730);
xnor U12411 (N_12411,N_7735,N_6734);
nand U12412 (N_12412,N_9102,N_9455);
or U12413 (N_12413,N_6912,N_9241);
and U12414 (N_12414,N_5587,N_5967);
nor U12415 (N_12415,N_8914,N_8395);
nor U12416 (N_12416,N_8927,N_6567);
nor U12417 (N_12417,N_7114,N_6291);
nor U12418 (N_12418,N_6793,N_6648);
and U12419 (N_12419,N_6078,N_9195);
nand U12420 (N_12420,N_8500,N_9603);
nor U12421 (N_12421,N_5351,N_9225);
nor U12422 (N_12422,N_8415,N_5442);
nand U12423 (N_12423,N_8308,N_6099);
or U12424 (N_12424,N_6217,N_9715);
nand U12425 (N_12425,N_7662,N_6635);
nand U12426 (N_12426,N_5500,N_9236);
and U12427 (N_12427,N_8441,N_8688);
or U12428 (N_12428,N_7464,N_6798);
or U12429 (N_12429,N_6039,N_9979);
nor U12430 (N_12430,N_6699,N_8695);
or U12431 (N_12431,N_5390,N_7385);
or U12432 (N_12432,N_6620,N_8111);
or U12433 (N_12433,N_5058,N_9194);
and U12434 (N_12434,N_6033,N_6808);
xnor U12435 (N_12435,N_7977,N_8542);
or U12436 (N_12436,N_7290,N_5361);
nor U12437 (N_12437,N_8376,N_9509);
nor U12438 (N_12438,N_7298,N_5231);
or U12439 (N_12439,N_7057,N_8829);
or U12440 (N_12440,N_8833,N_7565);
and U12441 (N_12441,N_7894,N_7006);
or U12442 (N_12442,N_7806,N_7654);
xor U12443 (N_12443,N_5330,N_5145);
nor U12444 (N_12444,N_8061,N_7397);
or U12445 (N_12445,N_9465,N_6634);
xor U12446 (N_12446,N_7307,N_8580);
nand U12447 (N_12447,N_5364,N_5867);
nand U12448 (N_12448,N_5061,N_9793);
and U12449 (N_12449,N_5284,N_8808);
nor U12450 (N_12450,N_9031,N_7423);
nand U12451 (N_12451,N_8673,N_8054);
nor U12452 (N_12452,N_5954,N_5564);
nand U12453 (N_12453,N_9630,N_6182);
nand U12454 (N_12454,N_9281,N_9012);
xnor U12455 (N_12455,N_7928,N_5884);
or U12456 (N_12456,N_9464,N_5950);
and U12457 (N_12457,N_5425,N_9778);
or U12458 (N_12458,N_6104,N_5845);
xnor U12459 (N_12459,N_6530,N_7578);
and U12460 (N_12460,N_8246,N_6915);
or U12461 (N_12461,N_9504,N_9008);
nor U12462 (N_12462,N_6674,N_8363);
nor U12463 (N_12463,N_9046,N_5848);
nand U12464 (N_12464,N_7498,N_6825);
nand U12465 (N_12465,N_6317,N_6982);
nor U12466 (N_12466,N_5662,N_7472);
nand U12467 (N_12467,N_7257,N_7861);
xor U12468 (N_12468,N_8346,N_8443);
nor U12469 (N_12469,N_5789,N_6060);
and U12470 (N_12470,N_7619,N_9107);
nand U12471 (N_12471,N_9426,N_6369);
nor U12472 (N_12472,N_8585,N_5551);
or U12473 (N_12473,N_5747,N_8498);
or U12474 (N_12474,N_8104,N_8380);
xnor U12475 (N_12475,N_6165,N_7650);
or U12476 (N_12476,N_6684,N_6226);
or U12477 (N_12477,N_9576,N_8962);
or U12478 (N_12478,N_9277,N_5868);
nor U12479 (N_12479,N_7492,N_6632);
nand U12480 (N_12480,N_6784,N_8908);
nor U12481 (N_12481,N_6162,N_9180);
nand U12482 (N_12482,N_7169,N_9271);
or U12483 (N_12483,N_5454,N_6561);
or U12484 (N_12484,N_9243,N_5580);
or U12485 (N_12485,N_5842,N_8425);
nand U12486 (N_12486,N_7196,N_8674);
nand U12487 (N_12487,N_8504,N_6537);
nand U12488 (N_12488,N_9735,N_8897);
or U12489 (N_12489,N_7605,N_7517);
nor U12490 (N_12490,N_8849,N_9099);
nor U12491 (N_12491,N_7406,N_9337);
nand U12492 (N_12492,N_8800,N_5184);
and U12493 (N_12493,N_9760,N_6727);
xnor U12494 (N_12494,N_6202,N_9971);
nand U12495 (N_12495,N_9183,N_8548);
nand U12496 (N_12496,N_6884,N_9842);
or U12497 (N_12497,N_8632,N_9343);
and U12498 (N_12498,N_5637,N_9419);
and U12499 (N_12499,N_7971,N_5334);
xnor U12500 (N_12500,N_9125,N_8097);
or U12501 (N_12501,N_6508,N_8698);
nor U12502 (N_12502,N_6800,N_5399);
xnor U12503 (N_12503,N_9663,N_7622);
nor U12504 (N_12504,N_6083,N_5554);
or U12505 (N_12505,N_9146,N_6360);
and U12506 (N_12506,N_9021,N_6271);
and U12507 (N_12507,N_9072,N_6017);
and U12508 (N_12508,N_7226,N_6482);
nor U12509 (N_12509,N_5534,N_8618);
nor U12510 (N_12510,N_5591,N_7911);
or U12511 (N_12511,N_9926,N_7384);
nand U12512 (N_12512,N_7671,N_6807);
or U12513 (N_12513,N_7896,N_8010);
nand U12514 (N_12514,N_5707,N_6480);
or U12515 (N_12515,N_9466,N_9972);
nand U12516 (N_12516,N_7471,N_5357);
or U12517 (N_12517,N_8351,N_6021);
and U12518 (N_12518,N_9067,N_6674);
or U12519 (N_12519,N_5751,N_8669);
nor U12520 (N_12520,N_6969,N_9094);
or U12521 (N_12521,N_5847,N_5114);
nand U12522 (N_12522,N_5075,N_8197);
and U12523 (N_12523,N_7319,N_9335);
nand U12524 (N_12524,N_9385,N_7345);
or U12525 (N_12525,N_5500,N_6610);
nor U12526 (N_12526,N_9716,N_8936);
and U12527 (N_12527,N_7647,N_5413);
and U12528 (N_12528,N_6286,N_5023);
and U12529 (N_12529,N_6462,N_7995);
xor U12530 (N_12530,N_5754,N_8739);
or U12531 (N_12531,N_6389,N_7114);
or U12532 (N_12532,N_5697,N_6202);
nor U12533 (N_12533,N_9226,N_7690);
nand U12534 (N_12534,N_5255,N_5297);
nand U12535 (N_12535,N_7592,N_6317);
nor U12536 (N_12536,N_8884,N_5453);
nand U12537 (N_12537,N_6654,N_8570);
nand U12538 (N_12538,N_9054,N_6188);
nor U12539 (N_12539,N_8710,N_6604);
and U12540 (N_12540,N_9590,N_6602);
xnor U12541 (N_12541,N_9006,N_9377);
nor U12542 (N_12542,N_9422,N_8567);
nand U12543 (N_12543,N_9080,N_7382);
and U12544 (N_12544,N_8407,N_9375);
nand U12545 (N_12545,N_5012,N_7744);
nor U12546 (N_12546,N_8274,N_6419);
nor U12547 (N_12547,N_5257,N_6426);
or U12548 (N_12548,N_5866,N_6407);
and U12549 (N_12549,N_9338,N_7448);
and U12550 (N_12550,N_8159,N_9564);
nand U12551 (N_12551,N_8467,N_8036);
or U12552 (N_12552,N_6201,N_5558);
nor U12553 (N_12553,N_5224,N_5235);
nor U12554 (N_12554,N_7367,N_5126);
xor U12555 (N_12555,N_7750,N_7140);
or U12556 (N_12556,N_5129,N_8145);
nor U12557 (N_12557,N_7163,N_7209);
and U12558 (N_12558,N_5470,N_8786);
and U12559 (N_12559,N_8458,N_5540);
xor U12560 (N_12560,N_6921,N_9996);
and U12561 (N_12561,N_9390,N_7668);
nor U12562 (N_12562,N_7451,N_8667);
nor U12563 (N_12563,N_9746,N_7680);
or U12564 (N_12564,N_5925,N_7571);
nand U12565 (N_12565,N_8884,N_6834);
nor U12566 (N_12566,N_9953,N_5117);
nor U12567 (N_12567,N_8875,N_7138);
or U12568 (N_12568,N_8568,N_7326);
and U12569 (N_12569,N_8595,N_7465);
or U12570 (N_12570,N_5469,N_7199);
nor U12571 (N_12571,N_9442,N_6882);
or U12572 (N_12572,N_7006,N_8462);
nor U12573 (N_12573,N_8274,N_5642);
xnor U12574 (N_12574,N_8950,N_5076);
or U12575 (N_12575,N_9019,N_5443);
or U12576 (N_12576,N_8092,N_6732);
and U12577 (N_12577,N_7751,N_9695);
or U12578 (N_12578,N_7526,N_5607);
and U12579 (N_12579,N_5812,N_5711);
nand U12580 (N_12580,N_5333,N_7601);
nand U12581 (N_12581,N_7596,N_9203);
nor U12582 (N_12582,N_6633,N_9386);
nor U12583 (N_12583,N_8612,N_7597);
nor U12584 (N_12584,N_9095,N_6169);
or U12585 (N_12585,N_5467,N_8839);
or U12586 (N_12586,N_5105,N_8748);
or U12587 (N_12587,N_9130,N_9906);
nor U12588 (N_12588,N_9177,N_9459);
nand U12589 (N_12589,N_7006,N_7724);
xor U12590 (N_12590,N_5332,N_5761);
or U12591 (N_12591,N_7412,N_7953);
or U12592 (N_12592,N_8304,N_5592);
and U12593 (N_12593,N_8172,N_5235);
nand U12594 (N_12594,N_5038,N_6243);
nor U12595 (N_12595,N_6736,N_5787);
nand U12596 (N_12596,N_5666,N_7543);
nand U12597 (N_12597,N_8126,N_7959);
nand U12598 (N_12598,N_9508,N_7905);
nand U12599 (N_12599,N_5121,N_6204);
xor U12600 (N_12600,N_5240,N_6322);
or U12601 (N_12601,N_8011,N_6541);
xor U12602 (N_12602,N_8446,N_9457);
xor U12603 (N_12603,N_6856,N_6073);
and U12604 (N_12604,N_9476,N_5704);
nand U12605 (N_12605,N_9876,N_7977);
and U12606 (N_12606,N_8851,N_7747);
or U12607 (N_12607,N_9448,N_5808);
or U12608 (N_12608,N_8755,N_8022);
nor U12609 (N_12609,N_6430,N_9593);
nor U12610 (N_12610,N_5057,N_8332);
nor U12611 (N_12611,N_5132,N_6291);
and U12612 (N_12612,N_5743,N_5541);
nor U12613 (N_12613,N_9504,N_9212);
or U12614 (N_12614,N_9917,N_9335);
xnor U12615 (N_12615,N_5698,N_8110);
or U12616 (N_12616,N_6020,N_7420);
or U12617 (N_12617,N_9096,N_8675);
nand U12618 (N_12618,N_7156,N_9668);
nand U12619 (N_12619,N_6152,N_9413);
or U12620 (N_12620,N_5321,N_8619);
nand U12621 (N_12621,N_6130,N_6028);
or U12622 (N_12622,N_9622,N_6337);
or U12623 (N_12623,N_6806,N_6773);
and U12624 (N_12624,N_6466,N_5036);
nor U12625 (N_12625,N_9903,N_6064);
or U12626 (N_12626,N_6125,N_5093);
and U12627 (N_12627,N_7367,N_7226);
and U12628 (N_12628,N_5525,N_9853);
nand U12629 (N_12629,N_7343,N_8288);
and U12630 (N_12630,N_8552,N_8699);
nor U12631 (N_12631,N_9866,N_8892);
nand U12632 (N_12632,N_6008,N_6596);
nand U12633 (N_12633,N_8455,N_6213);
or U12634 (N_12634,N_8788,N_9288);
and U12635 (N_12635,N_9823,N_7477);
or U12636 (N_12636,N_7402,N_7196);
nand U12637 (N_12637,N_8498,N_8133);
nor U12638 (N_12638,N_5570,N_6713);
nor U12639 (N_12639,N_8291,N_7795);
and U12640 (N_12640,N_5780,N_5030);
and U12641 (N_12641,N_5096,N_6856);
nand U12642 (N_12642,N_5231,N_7713);
and U12643 (N_12643,N_8756,N_7791);
nor U12644 (N_12644,N_5236,N_6260);
nand U12645 (N_12645,N_5617,N_6163);
nor U12646 (N_12646,N_6427,N_9510);
or U12647 (N_12647,N_6453,N_6392);
and U12648 (N_12648,N_6667,N_6976);
and U12649 (N_12649,N_5718,N_7011);
nand U12650 (N_12650,N_7146,N_7416);
nor U12651 (N_12651,N_5648,N_9965);
nor U12652 (N_12652,N_6331,N_7516);
or U12653 (N_12653,N_8958,N_8554);
or U12654 (N_12654,N_9474,N_9910);
nand U12655 (N_12655,N_5316,N_9908);
nand U12656 (N_12656,N_9687,N_6491);
nand U12657 (N_12657,N_8266,N_8118);
nand U12658 (N_12658,N_8836,N_7772);
or U12659 (N_12659,N_9992,N_7990);
and U12660 (N_12660,N_8907,N_5520);
nor U12661 (N_12661,N_7291,N_5183);
nor U12662 (N_12662,N_9817,N_6455);
nor U12663 (N_12663,N_6535,N_9935);
nor U12664 (N_12664,N_5528,N_5647);
and U12665 (N_12665,N_6970,N_8924);
nor U12666 (N_12666,N_7386,N_9007);
nand U12667 (N_12667,N_5419,N_7981);
xnor U12668 (N_12668,N_9431,N_8159);
or U12669 (N_12669,N_5638,N_8988);
and U12670 (N_12670,N_6292,N_6268);
and U12671 (N_12671,N_5822,N_6766);
and U12672 (N_12672,N_7431,N_8831);
nor U12673 (N_12673,N_8963,N_8623);
nor U12674 (N_12674,N_7165,N_8696);
and U12675 (N_12675,N_7875,N_6832);
nor U12676 (N_12676,N_6720,N_6409);
nor U12677 (N_12677,N_6533,N_6884);
xor U12678 (N_12678,N_5315,N_6446);
xnor U12679 (N_12679,N_8701,N_7961);
xor U12680 (N_12680,N_7582,N_7935);
and U12681 (N_12681,N_8506,N_5479);
or U12682 (N_12682,N_7680,N_8543);
nor U12683 (N_12683,N_6701,N_8379);
nor U12684 (N_12684,N_9495,N_7798);
nand U12685 (N_12685,N_9429,N_9109);
or U12686 (N_12686,N_7200,N_7219);
nor U12687 (N_12687,N_5355,N_5536);
nand U12688 (N_12688,N_6689,N_8107);
and U12689 (N_12689,N_8783,N_6825);
nand U12690 (N_12690,N_6860,N_9828);
nand U12691 (N_12691,N_6649,N_5306);
or U12692 (N_12692,N_7410,N_9903);
and U12693 (N_12693,N_9145,N_6798);
nor U12694 (N_12694,N_7017,N_6853);
nor U12695 (N_12695,N_5649,N_9905);
xor U12696 (N_12696,N_8152,N_5186);
nand U12697 (N_12697,N_8764,N_9616);
or U12698 (N_12698,N_8633,N_9206);
nand U12699 (N_12699,N_6725,N_6729);
nand U12700 (N_12700,N_8900,N_9312);
nand U12701 (N_12701,N_9480,N_9268);
and U12702 (N_12702,N_6786,N_5778);
xnor U12703 (N_12703,N_6672,N_5690);
nor U12704 (N_12704,N_8792,N_6966);
or U12705 (N_12705,N_7676,N_9334);
nor U12706 (N_12706,N_7318,N_8459);
or U12707 (N_12707,N_8687,N_8196);
and U12708 (N_12708,N_8835,N_9552);
nor U12709 (N_12709,N_7307,N_6884);
nor U12710 (N_12710,N_9792,N_8914);
or U12711 (N_12711,N_9244,N_6457);
or U12712 (N_12712,N_7291,N_6155);
nor U12713 (N_12713,N_6732,N_9525);
or U12714 (N_12714,N_6942,N_5401);
or U12715 (N_12715,N_7935,N_6786);
or U12716 (N_12716,N_6919,N_6891);
or U12717 (N_12717,N_9579,N_9486);
or U12718 (N_12718,N_5275,N_8688);
xnor U12719 (N_12719,N_5071,N_8008);
or U12720 (N_12720,N_5594,N_6926);
or U12721 (N_12721,N_8532,N_5098);
or U12722 (N_12722,N_6936,N_6922);
or U12723 (N_12723,N_5413,N_9332);
or U12724 (N_12724,N_6272,N_5292);
nor U12725 (N_12725,N_9364,N_6570);
and U12726 (N_12726,N_9397,N_9822);
nor U12727 (N_12727,N_5793,N_8190);
xnor U12728 (N_12728,N_9753,N_5598);
and U12729 (N_12729,N_7430,N_5305);
nand U12730 (N_12730,N_6725,N_7767);
nand U12731 (N_12731,N_7975,N_7668);
and U12732 (N_12732,N_6808,N_8868);
nand U12733 (N_12733,N_5567,N_7066);
or U12734 (N_12734,N_8005,N_6257);
or U12735 (N_12735,N_7632,N_8990);
nor U12736 (N_12736,N_8440,N_5156);
and U12737 (N_12737,N_7858,N_8211);
nand U12738 (N_12738,N_6568,N_9009);
and U12739 (N_12739,N_7892,N_9153);
and U12740 (N_12740,N_9685,N_7180);
and U12741 (N_12741,N_9753,N_7834);
or U12742 (N_12742,N_5657,N_5560);
nand U12743 (N_12743,N_6108,N_8145);
nand U12744 (N_12744,N_6652,N_8669);
nand U12745 (N_12745,N_9487,N_9877);
or U12746 (N_12746,N_5968,N_9100);
xnor U12747 (N_12747,N_7254,N_8437);
nand U12748 (N_12748,N_7202,N_9541);
nand U12749 (N_12749,N_9908,N_5213);
xor U12750 (N_12750,N_9372,N_7597);
nor U12751 (N_12751,N_8195,N_9975);
or U12752 (N_12752,N_6838,N_5649);
and U12753 (N_12753,N_6885,N_7873);
and U12754 (N_12754,N_7581,N_9811);
or U12755 (N_12755,N_6307,N_6915);
and U12756 (N_12756,N_7583,N_7998);
or U12757 (N_12757,N_8936,N_8384);
xnor U12758 (N_12758,N_7468,N_7041);
nor U12759 (N_12759,N_6359,N_8426);
or U12760 (N_12760,N_9479,N_7919);
or U12761 (N_12761,N_6530,N_8732);
nor U12762 (N_12762,N_7949,N_6932);
nand U12763 (N_12763,N_8802,N_5271);
and U12764 (N_12764,N_8163,N_8982);
nand U12765 (N_12765,N_9280,N_6421);
or U12766 (N_12766,N_8084,N_7167);
or U12767 (N_12767,N_5979,N_8466);
nor U12768 (N_12768,N_7118,N_9993);
and U12769 (N_12769,N_6728,N_5011);
nor U12770 (N_12770,N_9434,N_5485);
xnor U12771 (N_12771,N_6160,N_9134);
xor U12772 (N_12772,N_6546,N_6717);
nand U12773 (N_12773,N_7053,N_9104);
nand U12774 (N_12774,N_6042,N_6470);
or U12775 (N_12775,N_8674,N_5372);
xnor U12776 (N_12776,N_6965,N_8750);
and U12777 (N_12777,N_6303,N_7597);
or U12778 (N_12778,N_9042,N_7166);
or U12779 (N_12779,N_5605,N_6126);
or U12780 (N_12780,N_9409,N_9430);
nand U12781 (N_12781,N_6726,N_9801);
and U12782 (N_12782,N_8831,N_6980);
or U12783 (N_12783,N_6330,N_7666);
or U12784 (N_12784,N_5983,N_8459);
and U12785 (N_12785,N_9963,N_6302);
nand U12786 (N_12786,N_8328,N_9668);
and U12787 (N_12787,N_7077,N_5299);
or U12788 (N_12788,N_5655,N_7892);
or U12789 (N_12789,N_5866,N_9388);
and U12790 (N_12790,N_5771,N_6923);
xnor U12791 (N_12791,N_8298,N_7432);
or U12792 (N_12792,N_7355,N_6347);
or U12793 (N_12793,N_7910,N_6878);
nand U12794 (N_12794,N_8952,N_6636);
nor U12795 (N_12795,N_5159,N_5690);
nand U12796 (N_12796,N_9765,N_7128);
nand U12797 (N_12797,N_8756,N_7969);
xor U12798 (N_12798,N_6617,N_9488);
nand U12799 (N_12799,N_9825,N_8466);
or U12800 (N_12800,N_7055,N_8198);
nor U12801 (N_12801,N_6123,N_5482);
or U12802 (N_12802,N_8496,N_8909);
or U12803 (N_12803,N_9921,N_5520);
and U12804 (N_12804,N_8645,N_9065);
or U12805 (N_12805,N_8224,N_5791);
nor U12806 (N_12806,N_6584,N_5344);
or U12807 (N_12807,N_8041,N_6473);
xnor U12808 (N_12808,N_8219,N_9911);
or U12809 (N_12809,N_7825,N_8505);
nor U12810 (N_12810,N_8138,N_9795);
or U12811 (N_12811,N_8793,N_5867);
nand U12812 (N_12812,N_9088,N_9332);
nor U12813 (N_12813,N_7952,N_8365);
nor U12814 (N_12814,N_6325,N_7242);
nand U12815 (N_12815,N_5615,N_5520);
nor U12816 (N_12816,N_6164,N_8002);
nand U12817 (N_12817,N_5360,N_6522);
nor U12818 (N_12818,N_8490,N_6262);
nand U12819 (N_12819,N_6040,N_8441);
nor U12820 (N_12820,N_6262,N_6733);
or U12821 (N_12821,N_9503,N_8097);
nand U12822 (N_12822,N_6249,N_8005);
or U12823 (N_12823,N_7917,N_6133);
nand U12824 (N_12824,N_7939,N_9085);
nand U12825 (N_12825,N_7291,N_8908);
nor U12826 (N_12826,N_8578,N_8183);
xor U12827 (N_12827,N_6963,N_6576);
and U12828 (N_12828,N_5956,N_8399);
or U12829 (N_12829,N_5224,N_5290);
nor U12830 (N_12830,N_6201,N_8234);
or U12831 (N_12831,N_6803,N_8027);
or U12832 (N_12832,N_9533,N_9554);
or U12833 (N_12833,N_7618,N_6018);
and U12834 (N_12834,N_5764,N_8222);
and U12835 (N_12835,N_6796,N_8888);
nand U12836 (N_12836,N_7533,N_8471);
or U12837 (N_12837,N_6803,N_8522);
nor U12838 (N_12838,N_7770,N_6303);
xnor U12839 (N_12839,N_6877,N_7315);
or U12840 (N_12840,N_9793,N_9888);
or U12841 (N_12841,N_8601,N_6336);
nand U12842 (N_12842,N_5747,N_5987);
and U12843 (N_12843,N_5563,N_7390);
nor U12844 (N_12844,N_7691,N_9994);
nor U12845 (N_12845,N_9979,N_8838);
nor U12846 (N_12846,N_9613,N_9022);
and U12847 (N_12847,N_8483,N_7143);
and U12848 (N_12848,N_5957,N_5774);
nand U12849 (N_12849,N_8765,N_8891);
nand U12850 (N_12850,N_7171,N_5669);
or U12851 (N_12851,N_5151,N_6626);
xor U12852 (N_12852,N_6646,N_9416);
nand U12853 (N_12853,N_8411,N_6006);
and U12854 (N_12854,N_5275,N_8575);
and U12855 (N_12855,N_6376,N_9446);
xor U12856 (N_12856,N_6950,N_8556);
and U12857 (N_12857,N_5127,N_5510);
or U12858 (N_12858,N_7087,N_8741);
nor U12859 (N_12859,N_9052,N_9114);
nor U12860 (N_12860,N_9918,N_6191);
or U12861 (N_12861,N_5547,N_5522);
xnor U12862 (N_12862,N_7491,N_9145);
or U12863 (N_12863,N_5059,N_5481);
nand U12864 (N_12864,N_8146,N_5231);
xnor U12865 (N_12865,N_8879,N_6673);
nand U12866 (N_12866,N_9560,N_8850);
and U12867 (N_12867,N_8011,N_8218);
xnor U12868 (N_12868,N_9039,N_8132);
and U12869 (N_12869,N_9750,N_6592);
and U12870 (N_12870,N_8202,N_7296);
nor U12871 (N_12871,N_7931,N_9201);
and U12872 (N_12872,N_9982,N_8774);
or U12873 (N_12873,N_7413,N_8814);
or U12874 (N_12874,N_6325,N_8569);
and U12875 (N_12875,N_8701,N_7577);
or U12876 (N_12876,N_5146,N_6701);
or U12877 (N_12877,N_6617,N_6105);
and U12878 (N_12878,N_9415,N_8272);
and U12879 (N_12879,N_7214,N_5054);
or U12880 (N_12880,N_8566,N_6242);
nand U12881 (N_12881,N_8858,N_6297);
nand U12882 (N_12882,N_5478,N_5642);
nand U12883 (N_12883,N_9755,N_8490);
xor U12884 (N_12884,N_8177,N_7629);
nand U12885 (N_12885,N_9447,N_6591);
or U12886 (N_12886,N_7586,N_7958);
and U12887 (N_12887,N_5396,N_5849);
or U12888 (N_12888,N_6124,N_6664);
nand U12889 (N_12889,N_9615,N_8458);
nor U12890 (N_12890,N_8230,N_5803);
nand U12891 (N_12891,N_8769,N_9056);
xor U12892 (N_12892,N_9473,N_6544);
or U12893 (N_12893,N_7786,N_8739);
and U12894 (N_12894,N_5953,N_9319);
and U12895 (N_12895,N_7194,N_5703);
or U12896 (N_12896,N_9358,N_5885);
nand U12897 (N_12897,N_6198,N_6479);
nand U12898 (N_12898,N_8499,N_6799);
nand U12899 (N_12899,N_7510,N_5217);
nand U12900 (N_12900,N_7489,N_7291);
xnor U12901 (N_12901,N_9685,N_6984);
xor U12902 (N_12902,N_8591,N_7415);
nor U12903 (N_12903,N_9430,N_8155);
nand U12904 (N_12904,N_8367,N_6595);
nor U12905 (N_12905,N_5867,N_7566);
or U12906 (N_12906,N_5909,N_6453);
and U12907 (N_12907,N_8516,N_7862);
xnor U12908 (N_12908,N_8457,N_8845);
and U12909 (N_12909,N_8583,N_6494);
or U12910 (N_12910,N_8115,N_5995);
or U12911 (N_12911,N_8501,N_9489);
nor U12912 (N_12912,N_8418,N_8383);
nor U12913 (N_12913,N_8966,N_8516);
nand U12914 (N_12914,N_7963,N_5287);
nand U12915 (N_12915,N_9049,N_5889);
xor U12916 (N_12916,N_5541,N_8490);
or U12917 (N_12917,N_6812,N_6799);
nand U12918 (N_12918,N_9394,N_7871);
or U12919 (N_12919,N_6552,N_5967);
or U12920 (N_12920,N_7612,N_6489);
nor U12921 (N_12921,N_9411,N_7661);
nand U12922 (N_12922,N_6888,N_5635);
nand U12923 (N_12923,N_9454,N_8882);
and U12924 (N_12924,N_7869,N_5340);
nor U12925 (N_12925,N_9863,N_8050);
or U12926 (N_12926,N_5170,N_8381);
xnor U12927 (N_12927,N_8072,N_5315);
nor U12928 (N_12928,N_5905,N_7941);
nor U12929 (N_12929,N_7903,N_9266);
nand U12930 (N_12930,N_8795,N_6412);
and U12931 (N_12931,N_9262,N_6101);
nor U12932 (N_12932,N_9524,N_6546);
xnor U12933 (N_12933,N_7614,N_9694);
and U12934 (N_12934,N_5435,N_8507);
nor U12935 (N_12935,N_6505,N_8851);
or U12936 (N_12936,N_5561,N_7950);
nor U12937 (N_12937,N_6963,N_9026);
and U12938 (N_12938,N_5900,N_9717);
or U12939 (N_12939,N_9949,N_6281);
and U12940 (N_12940,N_7472,N_9858);
and U12941 (N_12941,N_5553,N_5748);
or U12942 (N_12942,N_7486,N_6825);
nor U12943 (N_12943,N_8189,N_5140);
nand U12944 (N_12944,N_9031,N_7282);
nor U12945 (N_12945,N_5874,N_8804);
xor U12946 (N_12946,N_5140,N_7207);
nand U12947 (N_12947,N_8932,N_8613);
and U12948 (N_12948,N_8938,N_9689);
nor U12949 (N_12949,N_9522,N_9548);
or U12950 (N_12950,N_7025,N_7862);
and U12951 (N_12951,N_7248,N_7635);
or U12952 (N_12952,N_8691,N_9754);
nand U12953 (N_12953,N_9669,N_9372);
xor U12954 (N_12954,N_8367,N_9432);
nand U12955 (N_12955,N_7306,N_9553);
and U12956 (N_12956,N_7170,N_6773);
nand U12957 (N_12957,N_5916,N_6610);
nor U12958 (N_12958,N_8665,N_6014);
xnor U12959 (N_12959,N_7925,N_6084);
and U12960 (N_12960,N_5141,N_7055);
xor U12961 (N_12961,N_5887,N_5566);
and U12962 (N_12962,N_7055,N_5731);
nand U12963 (N_12963,N_9026,N_8009);
nor U12964 (N_12964,N_7512,N_7205);
or U12965 (N_12965,N_7481,N_7367);
nor U12966 (N_12966,N_7891,N_5855);
nor U12967 (N_12967,N_9021,N_8936);
nand U12968 (N_12968,N_9566,N_8419);
or U12969 (N_12969,N_7246,N_8029);
and U12970 (N_12970,N_5254,N_5390);
or U12971 (N_12971,N_8643,N_6250);
or U12972 (N_12972,N_9657,N_8977);
or U12973 (N_12973,N_6062,N_6299);
and U12974 (N_12974,N_6422,N_9479);
nor U12975 (N_12975,N_9109,N_6771);
nand U12976 (N_12976,N_7607,N_8459);
nand U12977 (N_12977,N_9672,N_8749);
xor U12978 (N_12978,N_8870,N_9247);
and U12979 (N_12979,N_5265,N_8370);
nand U12980 (N_12980,N_9279,N_7613);
and U12981 (N_12981,N_7469,N_9562);
nand U12982 (N_12982,N_9770,N_5373);
and U12983 (N_12983,N_8579,N_5882);
or U12984 (N_12984,N_6187,N_7088);
or U12985 (N_12985,N_8396,N_7580);
nand U12986 (N_12986,N_5823,N_6529);
nor U12987 (N_12987,N_7944,N_7847);
nor U12988 (N_12988,N_6849,N_7987);
and U12989 (N_12989,N_9276,N_9203);
nand U12990 (N_12990,N_7184,N_6764);
nand U12991 (N_12991,N_7307,N_5116);
nand U12992 (N_12992,N_9324,N_7226);
or U12993 (N_12993,N_8941,N_7331);
and U12994 (N_12994,N_5955,N_7360);
and U12995 (N_12995,N_8046,N_7358);
nor U12996 (N_12996,N_8197,N_8433);
nor U12997 (N_12997,N_9118,N_5189);
nor U12998 (N_12998,N_6698,N_9603);
nor U12999 (N_12999,N_8391,N_6895);
nor U13000 (N_13000,N_8846,N_6619);
or U13001 (N_13001,N_9383,N_6073);
nor U13002 (N_13002,N_9636,N_6544);
nor U13003 (N_13003,N_8940,N_6140);
xnor U13004 (N_13004,N_9284,N_9225);
nand U13005 (N_13005,N_6847,N_5444);
or U13006 (N_13006,N_6641,N_5696);
nor U13007 (N_13007,N_6219,N_7717);
nor U13008 (N_13008,N_7621,N_8754);
nor U13009 (N_13009,N_9280,N_7962);
or U13010 (N_13010,N_6517,N_8783);
nand U13011 (N_13011,N_9932,N_6599);
nor U13012 (N_13012,N_9450,N_5948);
nand U13013 (N_13013,N_8507,N_7524);
nor U13014 (N_13014,N_5519,N_7464);
or U13015 (N_13015,N_9482,N_6195);
nor U13016 (N_13016,N_7950,N_8863);
and U13017 (N_13017,N_8658,N_7123);
nand U13018 (N_13018,N_6169,N_5177);
nand U13019 (N_13019,N_6701,N_8824);
nand U13020 (N_13020,N_7704,N_8668);
and U13021 (N_13021,N_5812,N_6961);
or U13022 (N_13022,N_6882,N_5210);
nand U13023 (N_13023,N_8437,N_9236);
nor U13024 (N_13024,N_5849,N_5149);
nor U13025 (N_13025,N_7573,N_8242);
nand U13026 (N_13026,N_7028,N_7494);
nor U13027 (N_13027,N_5042,N_5340);
nand U13028 (N_13028,N_7950,N_5123);
nand U13029 (N_13029,N_7310,N_5984);
nand U13030 (N_13030,N_5352,N_6957);
nand U13031 (N_13031,N_8825,N_6712);
xnor U13032 (N_13032,N_5854,N_7852);
or U13033 (N_13033,N_6990,N_6839);
or U13034 (N_13034,N_6335,N_9174);
nor U13035 (N_13035,N_7998,N_7000);
nand U13036 (N_13036,N_6105,N_5859);
xnor U13037 (N_13037,N_6702,N_7602);
and U13038 (N_13038,N_5431,N_6842);
nand U13039 (N_13039,N_6600,N_8487);
and U13040 (N_13040,N_8819,N_8053);
and U13041 (N_13041,N_7869,N_7014);
and U13042 (N_13042,N_5276,N_7251);
nand U13043 (N_13043,N_9068,N_7206);
nand U13044 (N_13044,N_5792,N_7643);
nand U13045 (N_13045,N_8172,N_7472);
nand U13046 (N_13046,N_9522,N_6254);
and U13047 (N_13047,N_6539,N_9292);
nand U13048 (N_13048,N_9499,N_9493);
nor U13049 (N_13049,N_7473,N_6588);
nand U13050 (N_13050,N_7171,N_9458);
and U13051 (N_13051,N_6211,N_6317);
and U13052 (N_13052,N_9211,N_9550);
and U13053 (N_13053,N_7589,N_6504);
nand U13054 (N_13054,N_8766,N_6930);
or U13055 (N_13055,N_9670,N_6320);
nor U13056 (N_13056,N_6528,N_6962);
nor U13057 (N_13057,N_5234,N_8767);
nor U13058 (N_13058,N_8284,N_8332);
or U13059 (N_13059,N_5355,N_9632);
nand U13060 (N_13060,N_8323,N_8631);
or U13061 (N_13061,N_9336,N_6336);
nor U13062 (N_13062,N_8318,N_9484);
or U13063 (N_13063,N_5609,N_7907);
nand U13064 (N_13064,N_8746,N_9737);
and U13065 (N_13065,N_6039,N_6690);
and U13066 (N_13066,N_8815,N_6926);
nor U13067 (N_13067,N_9864,N_5653);
xnor U13068 (N_13068,N_8672,N_5458);
or U13069 (N_13069,N_8983,N_5928);
or U13070 (N_13070,N_6090,N_9555);
nand U13071 (N_13071,N_6545,N_5015);
nor U13072 (N_13072,N_6009,N_5679);
or U13073 (N_13073,N_5712,N_7750);
nor U13074 (N_13074,N_5218,N_8137);
xor U13075 (N_13075,N_8497,N_7687);
and U13076 (N_13076,N_8526,N_8694);
nand U13077 (N_13077,N_8818,N_9950);
nand U13078 (N_13078,N_5541,N_6933);
or U13079 (N_13079,N_5571,N_6051);
nand U13080 (N_13080,N_8608,N_9828);
and U13081 (N_13081,N_9058,N_5311);
nand U13082 (N_13082,N_7829,N_6391);
xnor U13083 (N_13083,N_8891,N_7762);
nand U13084 (N_13084,N_8050,N_5482);
or U13085 (N_13085,N_5364,N_8914);
nand U13086 (N_13086,N_5837,N_7740);
or U13087 (N_13087,N_8443,N_9597);
nand U13088 (N_13088,N_9367,N_8274);
and U13089 (N_13089,N_8392,N_5915);
and U13090 (N_13090,N_6954,N_9178);
and U13091 (N_13091,N_7161,N_9039);
nor U13092 (N_13092,N_6342,N_9157);
xor U13093 (N_13093,N_5128,N_5099);
nor U13094 (N_13094,N_8032,N_7832);
and U13095 (N_13095,N_5053,N_7735);
and U13096 (N_13096,N_6853,N_9103);
or U13097 (N_13097,N_6205,N_6556);
nand U13098 (N_13098,N_6994,N_7632);
nor U13099 (N_13099,N_5237,N_6318);
and U13100 (N_13100,N_8757,N_9570);
xor U13101 (N_13101,N_9655,N_5421);
and U13102 (N_13102,N_5933,N_6945);
and U13103 (N_13103,N_8828,N_6588);
nor U13104 (N_13104,N_8784,N_5325);
and U13105 (N_13105,N_6357,N_9386);
and U13106 (N_13106,N_9774,N_7042);
xnor U13107 (N_13107,N_6723,N_5215);
and U13108 (N_13108,N_9624,N_8461);
xnor U13109 (N_13109,N_6128,N_5450);
nand U13110 (N_13110,N_7165,N_7440);
and U13111 (N_13111,N_9123,N_5742);
or U13112 (N_13112,N_6771,N_6263);
xor U13113 (N_13113,N_5514,N_9862);
nor U13114 (N_13114,N_6501,N_6487);
nor U13115 (N_13115,N_6593,N_9875);
and U13116 (N_13116,N_7076,N_7195);
or U13117 (N_13117,N_9359,N_6304);
xor U13118 (N_13118,N_5490,N_5273);
or U13119 (N_13119,N_7490,N_9694);
xnor U13120 (N_13120,N_9961,N_9285);
or U13121 (N_13121,N_7873,N_7327);
nor U13122 (N_13122,N_6274,N_8559);
nor U13123 (N_13123,N_9588,N_7970);
nand U13124 (N_13124,N_6906,N_8185);
nor U13125 (N_13125,N_6991,N_5596);
nor U13126 (N_13126,N_5240,N_7575);
xnor U13127 (N_13127,N_6437,N_8999);
nand U13128 (N_13128,N_9673,N_7096);
or U13129 (N_13129,N_5391,N_5205);
xnor U13130 (N_13130,N_8686,N_9253);
and U13131 (N_13131,N_5474,N_6030);
nor U13132 (N_13132,N_7997,N_9839);
nor U13133 (N_13133,N_6135,N_5031);
or U13134 (N_13134,N_5187,N_9529);
nand U13135 (N_13135,N_6622,N_5175);
nand U13136 (N_13136,N_5453,N_6942);
and U13137 (N_13137,N_7338,N_9703);
or U13138 (N_13138,N_6373,N_6172);
xnor U13139 (N_13139,N_9632,N_5668);
nor U13140 (N_13140,N_9600,N_7167);
and U13141 (N_13141,N_6370,N_9377);
xnor U13142 (N_13142,N_9366,N_8557);
nor U13143 (N_13143,N_6682,N_6068);
nor U13144 (N_13144,N_5811,N_8916);
and U13145 (N_13145,N_8866,N_6114);
nor U13146 (N_13146,N_6704,N_6759);
nor U13147 (N_13147,N_8296,N_6666);
and U13148 (N_13148,N_9384,N_8284);
nor U13149 (N_13149,N_6353,N_6280);
or U13150 (N_13150,N_8613,N_5363);
or U13151 (N_13151,N_5445,N_8580);
nor U13152 (N_13152,N_6779,N_8243);
nor U13153 (N_13153,N_9527,N_8780);
nand U13154 (N_13154,N_5709,N_6568);
nor U13155 (N_13155,N_6160,N_5370);
or U13156 (N_13156,N_6578,N_5466);
and U13157 (N_13157,N_8505,N_8406);
and U13158 (N_13158,N_8682,N_9799);
nor U13159 (N_13159,N_7208,N_6311);
nor U13160 (N_13160,N_5053,N_6792);
and U13161 (N_13161,N_7833,N_5548);
nor U13162 (N_13162,N_6168,N_5128);
or U13163 (N_13163,N_9103,N_9060);
and U13164 (N_13164,N_8512,N_8484);
and U13165 (N_13165,N_8648,N_7066);
nor U13166 (N_13166,N_5128,N_7651);
xnor U13167 (N_13167,N_8756,N_9116);
nor U13168 (N_13168,N_8985,N_8542);
nor U13169 (N_13169,N_5237,N_5367);
and U13170 (N_13170,N_9476,N_5568);
xor U13171 (N_13171,N_8434,N_6385);
xnor U13172 (N_13172,N_5597,N_9551);
and U13173 (N_13173,N_5233,N_8592);
or U13174 (N_13174,N_9866,N_6571);
and U13175 (N_13175,N_7725,N_5187);
and U13176 (N_13176,N_5203,N_9552);
or U13177 (N_13177,N_9481,N_9400);
and U13178 (N_13178,N_5704,N_7114);
and U13179 (N_13179,N_6007,N_6992);
and U13180 (N_13180,N_7767,N_6755);
nor U13181 (N_13181,N_7563,N_8392);
or U13182 (N_13182,N_9037,N_8701);
and U13183 (N_13183,N_7906,N_8154);
or U13184 (N_13184,N_6287,N_5596);
and U13185 (N_13185,N_7443,N_6736);
nand U13186 (N_13186,N_8084,N_9865);
nor U13187 (N_13187,N_7379,N_7078);
or U13188 (N_13188,N_8213,N_6083);
nor U13189 (N_13189,N_7713,N_5439);
nand U13190 (N_13190,N_6570,N_7715);
or U13191 (N_13191,N_5292,N_5288);
nor U13192 (N_13192,N_6208,N_6611);
xnor U13193 (N_13193,N_5748,N_6437);
nand U13194 (N_13194,N_7933,N_9509);
and U13195 (N_13195,N_9769,N_9531);
nor U13196 (N_13196,N_6180,N_8707);
nor U13197 (N_13197,N_9334,N_6594);
and U13198 (N_13198,N_7864,N_6468);
and U13199 (N_13199,N_6602,N_8990);
nand U13200 (N_13200,N_6208,N_8313);
nor U13201 (N_13201,N_9980,N_5822);
nand U13202 (N_13202,N_9797,N_9589);
nand U13203 (N_13203,N_7445,N_9728);
or U13204 (N_13204,N_6866,N_7983);
xor U13205 (N_13205,N_8081,N_9657);
nand U13206 (N_13206,N_9940,N_8944);
nand U13207 (N_13207,N_8211,N_6339);
nand U13208 (N_13208,N_6012,N_6667);
and U13209 (N_13209,N_9234,N_5964);
or U13210 (N_13210,N_8056,N_9497);
and U13211 (N_13211,N_9097,N_7003);
and U13212 (N_13212,N_7860,N_8237);
nand U13213 (N_13213,N_8621,N_6642);
or U13214 (N_13214,N_7842,N_8245);
nand U13215 (N_13215,N_5338,N_7702);
xor U13216 (N_13216,N_8198,N_8175);
xor U13217 (N_13217,N_6531,N_8601);
nor U13218 (N_13218,N_7849,N_8209);
nor U13219 (N_13219,N_6581,N_7428);
or U13220 (N_13220,N_8164,N_9801);
and U13221 (N_13221,N_6666,N_6873);
and U13222 (N_13222,N_6685,N_6798);
and U13223 (N_13223,N_9914,N_8188);
nand U13224 (N_13224,N_6533,N_5707);
or U13225 (N_13225,N_5734,N_6432);
and U13226 (N_13226,N_7197,N_7917);
nor U13227 (N_13227,N_9895,N_6621);
or U13228 (N_13228,N_9001,N_7388);
nor U13229 (N_13229,N_9139,N_7009);
or U13230 (N_13230,N_9037,N_8247);
and U13231 (N_13231,N_8675,N_8574);
xor U13232 (N_13232,N_9414,N_5115);
and U13233 (N_13233,N_5946,N_5383);
or U13234 (N_13234,N_9677,N_7843);
or U13235 (N_13235,N_7355,N_8419);
or U13236 (N_13236,N_6611,N_5633);
xnor U13237 (N_13237,N_6917,N_7657);
nand U13238 (N_13238,N_6562,N_9090);
nand U13239 (N_13239,N_7316,N_7705);
and U13240 (N_13240,N_7250,N_7546);
nor U13241 (N_13241,N_8057,N_7691);
nor U13242 (N_13242,N_8365,N_9890);
or U13243 (N_13243,N_9030,N_8065);
nor U13244 (N_13244,N_8994,N_7814);
or U13245 (N_13245,N_6519,N_8309);
nor U13246 (N_13246,N_8701,N_5274);
nand U13247 (N_13247,N_7437,N_9817);
xnor U13248 (N_13248,N_8621,N_6846);
nand U13249 (N_13249,N_6734,N_9819);
nor U13250 (N_13250,N_6619,N_7960);
nor U13251 (N_13251,N_8822,N_8383);
or U13252 (N_13252,N_9954,N_5531);
or U13253 (N_13253,N_6578,N_7627);
and U13254 (N_13254,N_8304,N_6492);
nand U13255 (N_13255,N_9598,N_7729);
nand U13256 (N_13256,N_9083,N_9656);
nor U13257 (N_13257,N_6894,N_6720);
nand U13258 (N_13258,N_8076,N_7127);
or U13259 (N_13259,N_8842,N_5290);
nand U13260 (N_13260,N_5662,N_9675);
and U13261 (N_13261,N_6137,N_8134);
xor U13262 (N_13262,N_6598,N_5689);
and U13263 (N_13263,N_6239,N_8840);
nor U13264 (N_13264,N_6201,N_7245);
and U13265 (N_13265,N_8952,N_7236);
or U13266 (N_13266,N_7714,N_7261);
and U13267 (N_13267,N_5214,N_6609);
or U13268 (N_13268,N_8048,N_8769);
nand U13269 (N_13269,N_8018,N_8341);
nor U13270 (N_13270,N_9895,N_9152);
nand U13271 (N_13271,N_7217,N_8594);
and U13272 (N_13272,N_9230,N_9183);
or U13273 (N_13273,N_8872,N_8893);
and U13274 (N_13274,N_9404,N_5435);
or U13275 (N_13275,N_7717,N_9381);
or U13276 (N_13276,N_8688,N_8226);
and U13277 (N_13277,N_6035,N_6353);
and U13278 (N_13278,N_5481,N_6694);
or U13279 (N_13279,N_9782,N_8572);
or U13280 (N_13280,N_9548,N_9309);
and U13281 (N_13281,N_6175,N_8836);
nor U13282 (N_13282,N_6585,N_6134);
nor U13283 (N_13283,N_6757,N_5808);
or U13284 (N_13284,N_7596,N_8566);
nand U13285 (N_13285,N_8385,N_9571);
nand U13286 (N_13286,N_6570,N_6054);
nand U13287 (N_13287,N_7416,N_9188);
xnor U13288 (N_13288,N_9254,N_8232);
nor U13289 (N_13289,N_7262,N_8916);
xor U13290 (N_13290,N_9346,N_8171);
nor U13291 (N_13291,N_5965,N_8094);
or U13292 (N_13292,N_8148,N_6297);
nand U13293 (N_13293,N_6614,N_8087);
nor U13294 (N_13294,N_6529,N_8979);
nor U13295 (N_13295,N_9578,N_5823);
nor U13296 (N_13296,N_6171,N_5987);
xor U13297 (N_13297,N_8855,N_9922);
nor U13298 (N_13298,N_8839,N_9808);
and U13299 (N_13299,N_8394,N_8471);
nand U13300 (N_13300,N_8442,N_6854);
or U13301 (N_13301,N_9636,N_5483);
or U13302 (N_13302,N_8399,N_9395);
or U13303 (N_13303,N_6627,N_7423);
xor U13304 (N_13304,N_5398,N_5292);
and U13305 (N_13305,N_9424,N_8370);
nor U13306 (N_13306,N_6181,N_5326);
nor U13307 (N_13307,N_7487,N_5923);
nand U13308 (N_13308,N_5586,N_7415);
and U13309 (N_13309,N_8064,N_9176);
or U13310 (N_13310,N_8238,N_7491);
nor U13311 (N_13311,N_5067,N_5907);
nand U13312 (N_13312,N_9301,N_9108);
nand U13313 (N_13313,N_8086,N_8329);
nand U13314 (N_13314,N_5639,N_5953);
or U13315 (N_13315,N_9907,N_6167);
and U13316 (N_13316,N_6561,N_8458);
or U13317 (N_13317,N_8713,N_8645);
or U13318 (N_13318,N_5616,N_9393);
and U13319 (N_13319,N_9013,N_7816);
or U13320 (N_13320,N_8545,N_6554);
nor U13321 (N_13321,N_5906,N_7495);
nand U13322 (N_13322,N_7247,N_5141);
nand U13323 (N_13323,N_8644,N_8125);
and U13324 (N_13324,N_8159,N_8042);
xnor U13325 (N_13325,N_5864,N_7177);
or U13326 (N_13326,N_5518,N_9404);
or U13327 (N_13327,N_9529,N_9401);
nor U13328 (N_13328,N_7787,N_7151);
nor U13329 (N_13329,N_6755,N_6247);
nand U13330 (N_13330,N_8263,N_6411);
nor U13331 (N_13331,N_9806,N_5807);
and U13332 (N_13332,N_8819,N_5403);
nand U13333 (N_13333,N_5660,N_7098);
xnor U13334 (N_13334,N_6212,N_8483);
nand U13335 (N_13335,N_5522,N_6078);
nand U13336 (N_13336,N_7159,N_7494);
and U13337 (N_13337,N_6985,N_6922);
nand U13338 (N_13338,N_5255,N_8096);
xor U13339 (N_13339,N_8387,N_9781);
nor U13340 (N_13340,N_6740,N_8469);
and U13341 (N_13341,N_9617,N_7024);
or U13342 (N_13342,N_5570,N_6960);
nand U13343 (N_13343,N_9942,N_6593);
nand U13344 (N_13344,N_9052,N_6937);
nand U13345 (N_13345,N_7580,N_6025);
nand U13346 (N_13346,N_7696,N_7875);
nand U13347 (N_13347,N_9280,N_8853);
or U13348 (N_13348,N_8271,N_7106);
xnor U13349 (N_13349,N_6166,N_9767);
and U13350 (N_13350,N_5880,N_6934);
nor U13351 (N_13351,N_6515,N_9245);
or U13352 (N_13352,N_7865,N_7845);
nand U13353 (N_13353,N_7418,N_6894);
or U13354 (N_13354,N_5879,N_8874);
nor U13355 (N_13355,N_8587,N_6579);
or U13356 (N_13356,N_6781,N_5140);
or U13357 (N_13357,N_6711,N_7522);
xor U13358 (N_13358,N_7701,N_9673);
nand U13359 (N_13359,N_9470,N_6762);
xnor U13360 (N_13360,N_6798,N_5824);
nand U13361 (N_13361,N_5847,N_8703);
nor U13362 (N_13362,N_6338,N_7087);
nand U13363 (N_13363,N_9537,N_7248);
nor U13364 (N_13364,N_5884,N_9191);
and U13365 (N_13365,N_9023,N_8230);
nor U13366 (N_13366,N_8817,N_6447);
and U13367 (N_13367,N_6764,N_9914);
or U13368 (N_13368,N_9323,N_6661);
or U13369 (N_13369,N_9759,N_9068);
nor U13370 (N_13370,N_5706,N_5707);
nand U13371 (N_13371,N_9464,N_5300);
and U13372 (N_13372,N_9161,N_6516);
nand U13373 (N_13373,N_9013,N_9962);
xor U13374 (N_13374,N_8502,N_9921);
and U13375 (N_13375,N_5707,N_6219);
nand U13376 (N_13376,N_6217,N_5336);
xnor U13377 (N_13377,N_7190,N_5358);
nor U13378 (N_13378,N_8411,N_5579);
and U13379 (N_13379,N_6514,N_6070);
nor U13380 (N_13380,N_7367,N_8771);
nor U13381 (N_13381,N_8943,N_8783);
nor U13382 (N_13382,N_6982,N_5428);
nand U13383 (N_13383,N_9274,N_8873);
nand U13384 (N_13384,N_8167,N_8510);
nand U13385 (N_13385,N_7508,N_6302);
nand U13386 (N_13386,N_5191,N_6770);
and U13387 (N_13387,N_8517,N_6281);
nand U13388 (N_13388,N_6188,N_8856);
nor U13389 (N_13389,N_9385,N_8954);
or U13390 (N_13390,N_7036,N_5368);
nand U13391 (N_13391,N_7767,N_7457);
nor U13392 (N_13392,N_5053,N_5908);
nor U13393 (N_13393,N_8485,N_7037);
nor U13394 (N_13394,N_6259,N_6267);
nor U13395 (N_13395,N_8797,N_7100);
or U13396 (N_13396,N_9594,N_8417);
and U13397 (N_13397,N_9398,N_6241);
and U13398 (N_13398,N_5675,N_6800);
and U13399 (N_13399,N_7103,N_5536);
or U13400 (N_13400,N_5501,N_6868);
nor U13401 (N_13401,N_7016,N_9578);
nor U13402 (N_13402,N_6749,N_9250);
or U13403 (N_13403,N_6935,N_9345);
nand U13404 (N_13404,N_9248,N_5135);
or U13405 (N_13405,N_8610,N_7310);
xnor U13406 (N_13406,N_7589,N_7069);
nor U13407 (N_13407,N_7738,N_7496);
or U13408 (N_13408,N_8043,N_8240);
or U13409 (N_13409,N_6233,N_5613);
or U13410 (N_13410,N_8753,N_8531);
xor U13411 (N_13411,N_7401,N_5150);
xnor U13412 (N_13412,N_5284,N_5372);
xnor U13413 (N_13413,N_9073,N_6283);
nor U13414 (N_13414,N_5014,N_8839);
or U13415 (N_13415,N_7540,N_9885);
nor U13416 (N_13416,N_5996,N_8300);
nand U13417 (N_13417,N_6579,N_7938);
or U13418 (N_13418,N_9580,N_9245);
nor U13419 (N_13419,N_5243,N_9228);
nand U13420 (N_13420,N_9798,N_8299);
and U13421 (N_13421,N_7288,N_8993);
nand U13422 (N_13422,N_8713,N_7168);
nor U13423 (N_13423,N_5497,N_7761);
nand U13424 (N_13424,N_9102,N_7632);
xnor U13425 (N_13425,N_9678,N_8233);
and U13426 (N_13426,N_6361,N_9805);
nand U13427 (N_13427,N_7897,N_5399);
or U13428 (N_13428,N_8807,N_8246);
xor U13429 (N_13429,N_5629,N_7546);
or U13430 (N_13430,N_9068,N_8799);
or U13431 (N_13431,N_9705,N_6157);
or U13432 (N_13432,N_7500,N_5787);
and U13433 (N_13433,N_5845,N_9401);
and U13434 (N_13434,N_9722,N_8080);
xnor U13435 (N_13435,N_7983,N_9770);
nand U13436 (N_13436,N_5557,N_6390);
nor U13437 (N_13437,N_8653,N_7936);
or U13438 (N_13438,N_8013,N_9255);
nand U13439 (N_13439,N_7546,N_9980);
nor U13440 (N_13440,N_7863,N_8001);
and U13441 (N_13441,N_7792,N_8384);
nand U13442 (N_13442,N_9368,N_5360);
nor U13443 (N_13443,N_9659,N_9008);
and U13444 (N_13444,N_5474,N_8264);
or U13445 (N_13445,N_6077,N_8513);
or U13446 (N_13446,N_9120,N_6700);
or U13447 (N_13447,N_7946,N_7616);
nand U13448 (N_13448,N_8108,N_7849);
nor U13449 (N_13449,N_5842,N_6237);
nand U13450 (N_13450,N_5018,N_7206);
and U13451 (N_13451,N_6746,N_5351);
and U13452 (N_13452,N_7733,N_7502);
and U13453 (N_13453,N_5958,N_8925);
and U13454 (N_13454,N_5019,N_6184);
or U13455 (N_13455,N_9732,N_9382);
nand U13456 (N_13456,N_7270,N_9679);
nor U13457 (N_13457,N_5422,N_9063);
nor U13458 (N_13458,N_6972,N_6688);
and U13459 (N_13459,N_7854,N_8798);
nand U13460 (N_13460,N_6702,N_6445);
and U13461 (N_13461,N_6536,N_8382);
nor U13462 (N_13462,N_7060,N_6444);
or U13463 (N_13463,N_7205,N_7588);
xor U13464 (N_13464,N_6585,N_8492);
or U13465 (N_13465,N_9510,N_8164);
or U13466 (N_13466,N_6514,N_6854);
nor U13467 (N_13467,N_7201,N_9423);
and U13468 (N_13468,N_5520,N_8521);
nand U13469 (N_13469,N_6281,N_7375);
xor U13470 (N_13470,N_7143,N_5984);
and U13471 (N_13471,N_5440,N_6812);
nand U13472 (N_13472,N_6339,N_6668);
or U13473 (N_13473,N_5034,N_6271);
nand U13474 (N_13474,N_7593,N_9054);
and U13475 (N_13475,N_6196,N_8713);
xor U13476 (N_13476,N_6926,N_9923);
or U13477 (N_13477,N_5050,N_5353);
xor U13478 (N_13478,N_9442,N_8714);
xnor U13479 (N_13479,N_9884,N_8032);
nand U13480 (N_13480,N_6661,N_5093);
and U13481 (N_13481,N_6835,N_5591);
xor U13482 (N_13482,N_7740,N_8359);
nor U13483 (N_13483,N_9862,N_8542);
or U13484 (N_13484,N_5575,N_7518);
or U13485 (N_13485,N_9940,N_9403);
nor U13486 (N_13486,N_8190,N_9787);
nand U13487 (N_13487,N_5231,N_9548);
or U13488 (N_13488,N_8318,N_7125);
or U13489 (N_13489,N_8485,N_6258);
xor U13490 (N_13490,N_8029,N_5753);
nand U13491 (N_13491,N_8243,N_9507);
nand U13492 (N_13492,N_6280,N_5698);
or U13493 (N_13493,N_6075,N_5991);
and U13494 (N_13494,N_9199,N_8708);
nor U13495 (N_13495,N_7186,N_9208);
and U13496 (N_13496,N_5909,N_6838);
nand U13497 (N_13497,N_5926,N_8562);
or U13498 (N_13498,N_5720,N_5263);
xnor U13499 (N_13499,N_8083,N_6985);
or U13500 (N_13500,N_7864,N_5977);
nor U13501 (N_13501,N_7021,N_7979);
xor U13502 (N_13502,N_7920,N_6675);
nor U13503 (N_13503,N_8491,N_5708);
nor U13504 (N_13504,N_7607,N_7626);
or U13505 (N_13505,N_8554,N_5217);
nor U13506 (N_13506,N_9991,N_5370);
or U13507 (N_13507,N_9968,N_7387);
nand U13508 (N_13508,N_9895,N_6740);
or U13509 (N_13509,N_7928,N_7956);
xor U13510 (N_13510,N_5289,N_8635);
or U13511 (N_13511,N_9332,N_7105);
and U13512 (N_13512,N_8018,N_6350);
or U13513 (N_13513,N_6085,N_9367);
and U13514 (N_13514,N_9131,N_7661);
nand U13515 (N_13515,N_9023,N_9731);
nand U13516 (N_13516,N_9092,N_7580);
nand U13517 (N_13517,N_7400,N_9099);
or U13518 (N_13518,N_8845,N_8597);
nor U13519 (N_13519,N_7909,N_8084);
or U13520 (N_13520,N_7866,N_6127);
and U13521 (N_13521,N_6805,N_6900);
or U13522 (N_13522,N_6296,N_5439);
or U13523 (N_13523,N_8319,N_5817);
or U13524 (N_13524,N_9823,N_6252);
nand U13525 (N_13525,N_8377,N_6940);
or U13526 (N_13526,N_8652,N_8957);
or U13527 (N_13527,N_5955,N_6992);
or U13528 (N_13528,N_8945,N_6778);
and U13529 (N_13529,N_5034,N_7837);
nor U13530 (N_13530,N_9636,N_5583);
xor U13531 (N_13531,N_5648,N_5601);
and U13532 (N_13532,N_5782,N_5464);
nor U13533 (N_13533,N_6541,N_6210);
nor U13534 (N_13534,N_9925,N_5762);
nor U13535 (N_13535,N_5789,N_8452);
and U13536 (N_13536,N_8758,N_8333);
or U13537 (N_13537,N_9732,N_9796);
nor U13538 (N_13538,N_6060,N_9013);
nand U13539 (N_13539,N_9926,N_6525);
nor U13540 (N_13540,N_8762,N_7533);
and U13541 (N_13541,N_8320,N_9528);
nor U13542 (N_13542,N_7484,N_8983);
and U13543 (N_13543,N_7999,N_8003);
nor U13544 (N_13544,N_8359,N_7173);
nand U13545 (N_13545,N_9774,N_7919);
and U13546 (N_13546,N_9374,N_7662);
nand U13547 (N_13547,N_9405,N_8371);
nand U13548 (N_13548,N_8106,N_5297);
or U13549 (N_13549,N_5821,N_8936);
and U13550 (N_13550,N_8236,N_9008);
nor U13551 (N_13551,N_5865,N_9524);
nor U13552 (N_13552,N_6773,N_7380);
nand U13553 (N_13553,N_8744,N_7596);
and U13554 (N_13554,N_7436,N_6835);
nand U13555 (N_13555,N_5828,N_5166);
or U13556 (N_13556,N_6327,N_6888);
and U13557 (N_13557,N_8272,N_8040);
nor U13558 (N_13558,N_7043,N_6708);
nand U13559 (N_13559,N_6462,N_5152);
or U13560 (N_13560,N_8441,N_8628);
nand U13561 (N_13561,N_9330,N_8286);
nor U13562 (N_13562,N_5211,N_9390);
nand U13563 (N_13563,N_5951,N_9693);
or U13564 (N_13564,N_6923,N_8010);
or U13565 (N_13565,N_9622,N_7779);
nor U13566 (N_13566,N_7091,N_5619);
nand U13567 (N_13567,N_6936,N_6039);
nor U13568 (N_13568,N_5088,N_7005);
or U13569 (N_13569,N_7149,N_7696);
nand U13570 (N_13570,N_9723,N_5263);
nor U13571 (N_13571,N_5402,N_5092);
and U13572 (N_13572,N_9533,N_7011);
nor U13573 (N_13573,N_5410,N_6828);
and U13574 (N_13574,N_8682,N_9100);
nor U13575 (N_13575,N_7036,N_9040);
or U13576 (N_13576,N_5407,N_6613);
or U13577 (N_13577,N_9604,N_7737);
xor U13578 (N_13578,N_7406,N_8833);
or U13579 (N_13579,N_9059,N_5678);
or U13580 (N_13580,N_8497,N_8909);
nand U13581 (N_13581,N_6178,N_9416);
and U13582 (N_13582,N_7668,N_6116);
or U13583 (N_13583,N_7158,N_9913);
or U13584 (N_13584,N_5778,N_5374);
or U13585 (N_13585,N_5916,N_6752);
xor U13586 (N_13586,N_7954,N_6043);
and U13587 (N_13587,N_8402,N_7945);
or U13588 (N_13588,N_9937,N_6474);
nor U13589 (N_13589,N_9438,N_7210);
and U13590 (N_13590,N_9677,N_6109);
nand U13591 (N_13591,N_7635,N_6805);
nor U13592 (N_13592,N_8399,N_9208);
nand U13593 (N_13593,N_7751,N_6896);
or U13594 (N_13594,N_7321,N_5856);
xor U13595 (N_13595,N_7177,N_7290);
nor U13596 (N_13596,N_5998,N_8453);
or U13597 (N_13597,N_5835,N_8127);
and U13598 (N_13598,N_5853,N_5349);
and U13599 (N_13599,N_5321,N_6334);
xnor U13600 (N_13600,N_7800,N_8706);
nor U13601 (N_13601,N_5018,N_5712);
nand U13602 (N_13602,N_7783,N_7249);
nand U13603 (N_13603,N_7328,N_6809);
or U13604 (N_13604,N_5353,N_9664);
and U13605 (N_13605,N_5209,N_8771);
nor U13606 (N_13606,N_9469,N_8609);
xor U13607 (N_13607,N_8428,N_6845);
or U13608 (N_13608,N_6350,N_5975);
nor U13609 (N_13609,N_6752,N_6908);
and U13610 (N_13610,N_8438,N_8973);
nor U13611 (N_13611,N_9263,N_5173);
and U13612 (N_13612,N_8034,N_8043);
nor U13613 (N_13613,N_5609,N_9607);
or U13614 (N_13614,N_7518,N_9169);
or U13615 (N_13615,N_5891,N_9250);
nand U13616 (N_13616,N_7222,N_5463);
or U13617 (N_13617,N_9016,N_5808);
and U13618 (N_13618,N_5285,N_5842);
nor U13619 (N_13619,N_5309,N_8993);
or U13620 (N_13620,N_8082,N_5123);
nand U13621 (N_13621,N_8826,N_9422);
nand U13622 (N_13622,N_6302,N_6256);
and U13623 (N_13623,N_5738,N_9793);
xor U13624 (N_13624,N_9582,N_5560);
or U13625 (N_13625,N_8573,N_7326);
nand U13626 (N_13626,N_6368,N_7249);
and U13627 (N_13627,N_9796,N_9768);
and U13628 (N_13628,N_9865,N_6185);
and U13629 (N_13629,N_9987,N_9778);
or U13630 (N_13630,N_7386,N_9937);
or U13631 (N_13631,N_6936,N_9226);
or U13632 (N_13632,N_8212,N_6496);
nor U13633 (N_13633,N_7891,N_5985);
nand U13634 (N_13634,N_8285,N_9220);
or U13635 (N_13635,N_5804,N_6600);
nand U13636 (N_13636,N_9408,N_9777);
nor U13637 (N_13637,N_8425,N_8476);
nor U13638 (N_13638,N_8025,N_9502);
or U13639 (N_13639,N_6924,N_8754);
nand U13640 (N_13640,N_8039,N_6494);
nor U13641 (N_13641,N_5276,N_9541);
and U13642 (N_13642,N_5932,N_6930);
nor U13643 (N_13643,N_6290,N_7779);
nor U13644 (N_13644,N_5702,N_8495);
nor U13645 (N_13645,N_9516,N_7937);
or U13646 (N_13646,N_9278,N_9275);
nor U13647 (N_13647,N_5298,N_9231);
or U13648 (N_13648,N_8280,N_6668);
and U13649 (N_13649,N_8677,N_5625);
nand U13650 (N_13650,N_7415,N_7964);
nand U13651 (N_13651,N_5858,N_7269);
or U13652 (N_13652,N_9432,N_6700);
nor U13653 (N_13653,N_9977,N_7513);
nand U13654 (N_13654,N_5280,N_6922);
and U13655 (N_13655,N_8401,N_8591);
and U13656 (N_13656,N_8029,N_9491);
and U13657 (N_13657,N_7973,N_6265);
or U13658 (N_13658,N_9326,N_9530);
and U13659 (N_13659,N_5421,N_6036);
nor U13660 (N_13660,N_6423,N_8458);
and U13661 (N_13661,N_8772,N_6900);
and U13662 (N_13662,N_5728,N_7426);
nor U13663 (N_13663,N_9147,N_5404);
nor U13664 (N_13664,N_6986,N_9187);
nand U13665 (N_13665,N_6723,N_9613);
xor U13666 (N_13666,N_7311,N_5793);
or U13667 (N_13667,N_6380,N_6678);
nand U13668 (N_13668,N_5991,N_5879);
or U13669 (N_13669,N_6076,N_8013);
nand U13670 (N_13670,N_8957,N_7508);
nor U13671 (N_13671,N_6598,N_9390);
or U13672 (N_13672,N_9015,N_9832);
or U13673 (N_13673,N_8963,N_6822);
nor U13674 (N_13674,N_7207,N_7121);
nor U13675 (N_13675,N_5400,N_9762);
xnor U13676 (N_13676,N_6638,N_9835);
nand U13677 (N_13677,N_6705,N_6506);
or U13678 (N_13678,N_5469,N_7260);
xnor U13679 (N_13679,N_8218,N_6171);
nor U13680 (N_13680,N_8324,N_8234);
or U13681 (N_13681,N_6676,N_5478);
nand U13682 (N_13682,N_8835,N_7692);
and U13683 (N_13683,N_7604,N_8039);
nor U13684 (N_13684,N_8031,N_5029);
nand U13685 (N_13685,N_9587,N_6328);
nor U13686 (N_13686,N_7513,N_7380);
and U13687 (N_13687,N_8944,N_8357);
nand U13688 (N_13688,N_9517,N_7033);
nand U13689 (N_13689,N_8008,N_9212);
nor U13690 (N_13690,N_9092,N_9022);
nor U13691 (N_13691,N_6953,N_7053);
and U13692 (N_13692,N_8569,N_9063);
nor U13693 (N_13693,N_6721,N_9110);
nand U13694 (N_13694,N_8660,N_6459);
or U13695 (N_13695,N_8382,N_7072);
or U13696 (N_13696,N_6338,N_7123);
nor U13697 (N_13697,N_7549,N_5356);
nand U13698 (N_13698,N_7937,N_8986);
or U13699 (N_13699,N_8270,N_6010);
nor U13700 (N_13700,N_6168,N_8347);
nand U13701 (N_13701,N_9306,N_8119);
xor U13702 (N_13702,N_5989,N_6143);
nand U13703 (N_13703,N_6573,N_9232);
and U13704 (N_13704,N_9026,N_7538);
and U13705 (N_13705,N_6092,N_6011);
nand U13706 (N_13706,N_7213,N_5562);
xnor U13707 (N_13707,N_6072,N_6668);
or U13708 (N_13708,N_7763,N_9337);
nor U13709 (N_13709,N_7108,N_7051);
and U13710 (N_13710,N_7156,N_7966);
and U13711 (N_13711,N_7743,N_9832);
and U13712 (N_13712,N_5849,N_8579);
nor U13713 (N_13713,N_6559,N_7578);
or U13714 (N_13714,N_9251,N_7438);
or U13715 (N_13715,N_6666,N_7640);
nand U13716 (N_13716,N_5003,N_5135);
nand U13717 (N_13717,N_7637,N_6598);
xor U13718 (N_13718,N_5251,N_7636);
or U13719 (N_13719,N_8154,N_6351);
xnor U13720 (N_13720,N_7930,N_8112);
or U13721 (N_13721,N_6932,N_7392);
nand U13722 (N_13722,N_9009,N_6751);
nor U13723 (N_13723,N_9210,N_8670);
or U13724 (N_13724,N_5155,N_9081);
and U13725 (N_13725,N_5290,N_8959);
and U13726 (N_13726,N_7615,N_6655);
or U13727 (N_13727,N_5555,N_5539);
and U13728 (N_13728,N_6717,N_9649);
and U13729 (N_13729,N_7484,N_9964);
and U13730 (N_13730,N_6516,N_5427);
nand U13731 (N_13731,N_6979,N_5047);
nor U13732 (N_13732,N_7852,N_9743);
nor U13733 (N_13733,N_8167,N_7374);
and U13734 (N_13734,N_9099,N_5560);
nand U13735 (N_13735,N_9838,N_9292);
and U13736 (N_13736,N_5094,N_5585);
or U13737 (N_13737,N_7240,N_6756);
nand U13738 (N_13738,N_8483,N_6261);
or U13739 (N_13739,N_9740,N_9780);
nor U13740 (N_13740,N_9002,N_7164);
nand U13741 (N_13741,N_9615,N_9950);
or U13742 (N_13742,N_6555,N_8004);
nand U13743 (N_13743,N_7203,N_6375);
or U13744 (N_13744,N_5427,N_9260);
and U13745 (N_13745,N_8603,N_6596);
nor U13746 (N_13746,N_6151,N_6023);
or U13747 (N_13747,N_7336,N_6282);
and U13748 (N_13748,N_8585,N_9480);
or U13749 (N_13749,N_8501,N_5185);
nand U13750 (N_13750,N_9231,N_7077);
or U13751 (N_13751,N_7268,N_6976);
or U13752 (N_13752,N_5255,N_9565);
xor U13753 (N_13753,N_7365,N_6020);
xor U13754 (N_13754,N_6368,N_5130);
and U13755 (N_13755,N_7218,N_8544);
nor U13756 (N_13756,N_9698,N_6565);
or U13757 (N_13757,N_6827,N_8960);
and U13758 (N_13758,N_8345,N_5429);
nor U13759 (N_13759,N_6716,N_6147);
nor U13760 (N_13760,N_7948,N_5558);
nor U13761 (N_13761,N_5858,N_6719);
or U13762 (N_13762,N_9986,N_6947);
or U13763 (N_13763,N_8857,N_7405);
or U13764 (N_13764,N_7200,N_5709);
and U13765 (N_13765,N_7847,N_7793);
nand U13766 (N_13766,N_5147,N_5298);
and U13767 (N_13767,N_5612,N_6104);
xnor U13768 (N_13768,N_7872,N_9532);
or U13769 (N_13769,N_6880,N_5478);
and U13770 (N_13770,N_7509,N_7760);
nand U13771 (N_13771,N_6862,N_7659);
or U13772 (N_13772,N_6046,N_5109);
and U13773 (N_13773,N_9713,N_8841);
and U13774 (N_13774,N_5962,N_6795);
nor U13775 (N_13775,N_8995,N_9176);
or U13776 (N_13776,N_9027,N_5201);
nand U13777 (N_13777,N_9722,N_8123);
and U13778 (N_13778,N_6880,N_9288);
nand U13779 (N_13779,N_9971,N_9724);
xor U13780 (N_13780,N_8300,N_6447);
nand U13781 (N_13781,N_7711,N_7120);
xor U13782 (N_13782,N_8264,N_9159);
or U13783 (N_13783,N_9064,N_5130);
nor U13784 (N_13784,N_8143,N_6458);
and U13785 (N_13785,N_8690,N_6878);
nor U13786 (N_13786,N_9032,N_9267);
or U13787 (N_13787,N_6584,N_8974);
and U13788 (N_13788,N_9674,N_5032);
and U13789 (N_13789,N_7231,N_8386);
and U13790 (N_13790,N_8385,N_7401);
nand U13791 (N_13791,N_5796,N_5201);
and U13792 (N_13792,N_7287,N_5308);
xnor U13793 (N_13793,N_9148,N_8683);
nor U13794 (N_13794,N_7014,N_8486);
or U13795 (N_13795,N_9918,N_7683);
xor U13796 (N_13796,N_5356,N_8043);
or U13797 (N_13797,N_7167,N_9408);
or U13798 (N_13798,N_8327,N_5282);
nand U13799 (N_13799,N_8959,N_7308);
xnor U13800 (N_13800,N_6422,N_5693);
or U13801 (N_13801,N_8636,N_9364);
xnor U13802 (N_13802,N_7563,N_9768);
nand U13803 (N_13803,N_5153,N_6040);
nand U13804 (N_13804,N_6613,N_9477);
and U13805 (N_13805,N_5391,N_9525);
xor U13806 (N_13806,N_9980,N_7895);
and U13807 (N_13807,N_5473,N_5378);
and U13808 (N_13808,N_7438,N_9239);
or U13809 (N_13809,N_9118,N_6521);
xnor U13810 (N_13810,N_9923,N_9930);
xor U13811 (N_13811,N_6467,N_7614);
xnor U13812 (N_13812,N_9063,N_6612);
nand U13813 (N_13813,N_5457,N_9054);
xnor U13814 (N_13814,N_5356,N_6258);
xor U13815 (N_13815,N_8150,N_7477);
nand U13816 (N_13816,N_9043,N_7879);
nand U13817 (N_13817,N_7128,N_8790);
nor U13818 (N_13818,N_6163,N_8477);
nand U13819 (N_13819,N_9873,N_9623);
and U13820 (N_13820,N_5099,N_7104);
nor U13821 (N_13821,N_7120,N_6823);
nor U13822 (N_13822,N_8460,N_9137);
and U13823 (N_13823,N_8506,N_6849);
or U13824 (N_13824,N_7089,N_5791);
nor U13825 (N_13825,N_8598,N_6841);
xor U13826 (N_13826,N_9303,N_8710);
nor U13827 (N_13827,N_6096,N_8475);
or U13828 (N_13828,N_9712,N_9692);
nand U13829 (N_13829,N_9159,N_6559);
nand U13830 (N_13830,N_8783,N_8668);
nand U13831 (N_13831,N_9110,N_5391);
nand U13832 (N_13832,N_7122,N_9436);
and U13833 (N_13833,N_5318,N_9260);
and U13834 (N_13834,N_5277,N_9623);
nand U13835 (N_13835,N_5271,N_6922);
nand U13836 (N_13836,N_7899,N_8589);
or U13837 (N_13837,N_8062,N_8661);
nor U13838 (N_13838,N_8861,N_7484);
or U13839 (N_13839,N_9408,N_7249);
xnor U13840 (N_13840,N_9635,N_9044);
or U13841 (N_13841,N_9878,N_7781);
and U13842 (N_13842,N_9004,N_8118);
or U13843 (N_13843,N_9271,N_7188);
and U13844 (N_13844,N_5409,N_9878);
nand U13845 (N_13845,N_7653,N_5562);
and U13846 (N_13846,N_9150,N_5389);
and U13847 (N_13847,N_6437,N_5696);
or U13848 (N_13848,N_6632,N_5001);
nor U13849 (N_13849,N_7593,N_8533);
or U13850 (N_13850,N_8759,N_8743);
nor U13851 (N_13851,N_6470,N_6991);
nand U13852 (N_13852,N_7466,N_7317);
or U13853 (N_13853,N_7020,N_7639);
nor U13854 (N_13854,N_7665,N_9938);
nor U13855 (N_13855,N_7428,N_6635);
nor U13856 (N_13856,N_6356,N_9989);
and U13857 (N_13857,N_9709,N_6217);
and U13858 (N_13858,N_5188,N_6622);
or U13859 (N_13859,N_7984,N_8302);
and U13860 (N_13860,N_6932,N_6197);
nand U13861 (N_13861,N_6900,N_6989);
xor U13862 (N_13862,N_5039,N_7540);
or U13863 (N_13863,N_5270,N_5348);
and U13864 (N_13864,N_8794,N_8205);
and U13865 (N_13865,N_8643,N_7587);
nand U13866 (N_13866,N_5838,N_8844);
and U13867 (N_13867,N_7751,N_5975);
and U13868 (N_13868,N_7702,N_8726);
nand U13869 (N_13869,N_5453,N_6352);
nand U13870 (N_13870,N_9078,N_5938);
nand U13871 (N_13871,N_9422,N_7881);
and U13872 (N_13872,N_9862,N_8371);
nand U13873 (N_13873,N_5187,N_8352);
nand U13874 (N_13874,N_9811,N_9914);
nor U13875 (N_13875,N_5814,N_5369);
nand U13876 (N_13876,N_8708,N_9543);
nand U13877 (N_13877,N_9952,N_5133);
nand U13878 (N_13878,N_8200,N_6530);
nor U13879 (N_13879,N_6207,N_6009);
and U13880 (N_13880,N_8368,N_5679);
nor U13881 (N_13881,N_9317,N_7384);
nand U13882 (N_13882,N_5316,N_6294);
or U13883 (N_13883,N_5349,N_5197);
and U13884 (N_13884,N_9978,N_9916);
nor U13885 (N_13885,N_9895,N_8392);
or U13886 (N_13886,N_8333,N_8076);
nor U13887 (N_13887,N_9581,N_7424);
and U13888 (N_13888,N_6905,N_9897);
nor U13889 (N_13889,N_7691,N_6357);
and U13890 (N_13890,N_7406,N_5766);
nor U13891 (N_13891,N_7873,N_5201);
or U13892 (N_13892,N_7933,N_8887);
or U13893 (N_13893,N_7465,N_6372);
nor U13894 (N_13894,N_5222,N_7727);
nand U13895 (N_13895,N_9522,N_8759);
or U13896 (N_13896,N_6674,N_6488);
and U13897 (N_13897,N_6348,N_6247);
or U13898 (N_13898,N_7237,N_5845);
xnor U13899 (N_13899,N_8572,N_5389);
nand U13900 (N_13900,N_7789,N_6642);
and U13901 (N_13901,N_8288,N_5143);
nor U13902 (N_13902,N_6475,N_9622);
nand U13903 (N_13903,N_8854,N_9084);
nor U13904 (N_13904,N_9274,N_9028);
or U13905 (N_13905,N_6658,N_7961);
xnor U13906 (N_13906,N_5629,N_6157);
and U13907 (N_13907,N_8599,N_5484);
nand U13908 (N_13908,N_6719,N_8003);
and U13909 (N_13909,N_6989,N_7180);
nor U13910 (N_13910,N_6373,N_8575);
or U13911 (N_13911,N_5481,N_8783);
and U13912 (N_13912,N_6130,N_9940);
xor U13913 (N_13913,N_9487,N_7167);
nor U13914 (N_13914,N_8318,N_9252);
and U13915 (N_13915,N_9970,N_5298);
nand U13916 (N_13916,N_5387,N_8371);
nor U13917 (N_13917,N_7197,N_9137);
nand U13918 (N_13918,N_5216,N_5493);
and U13919 (N_13919,N_8737,N_9918);
nor U13920 (N_13920,N_9368,N_7026);
nor U13921 (N_13921,N_8857,N_7175);
or U13922 (N_13922,N_7735,N_9530);
nand U13923 (N_13923,N_8030,N_9850);
nor U13924 (N_13924,N_7755,N_6593);
nor U13925 (N_13925,N_6386,N_7461);
nor U13926 (N_13926,N_8924,N_6479);
nor U13927 (N_13927,N_9227,N_6084);
and U13928 (N_13928,N_6420,N_7247);
nor U13929 (N_13929,N_7006,N_6660);
nor U13930 (N_13930,N_6254,N_9049);
and U13931 (N_13931,N_8150,N_8686);
or U13932 (N_13932,N_9976,N_5461);
nand U13933 (N_13933,N_8801,N_8660);
nand U13934 (N_13934,N_9136,N_6911);
xnor U13935 (N_13935,N_6847,N_8151);
or U13936 (N_13936,N_8189,N_8797);
nand U13937 (N_13937,N_7889,N_7207);
or U13938 (N_13938,N_9359,N_9612);
nand U13939 (N_13939,N_5461,N_6758);
or U13940 (N_13940,N_9246,N_8863);
or U13941 (N_13941,N_9330,N_9738);
or U13942 (N_13942,N_5581,N_5418);
nand U13943 (N_13943,N_5412,N_6910);
or U13944 (N_13944,N_9119,N_6524);
nor U13945 (N_13945,N_8930,N_6440);
nand U13946 (N_13946,N_9227,N_5016);
nor U13947 (N_13947,N_8290,N_8840);
and U13948 (N_13948,N_8725,N_6201);
and U13949 (N_13949,N_7244,N_9559);
nor U13950 (N_13950,N_6551,N_7074);
or U13951 (N_13951,N_7118,N_9413);
and U13952 (N_13952,N_8216,N_8070);
or U13953 (N_13953,N_7186,N_8844);
nor U13954 (N_13954,N_9912,N_7342);
nor U13955 (N_13955,N_7944,N_9582);
and U13956 (N_13956,N_7165,N_8949);
nand U13957 (N_13957,N_8128,N_9649);
xor U13958 (N_13958,N_5682,N_8599);
xnor U13959 (N_13959,N_7185,N_7916);
nand U13960 (N_13960,N_7201,N_5254);
nor U13961 (N_13961,N_8082,N_5130);
or U13962 (N_13962,N_8565,N_6073);
and U13963 (N_13963,N_7073,N_8539);
or U13964 (N_13964,N_7964,N_9594);
and U13965 (N_13965,N_6253,N_6362);
or U13966 (N_13966,N_7579,N_9835);
nor U13967 (N_13967,N_9890,N_9202);
or U13968 (N_13968,N_5402,N_5449);
or U13969 (N_13969,N_6028,N_7206);
or U13970 (N_13970,N_5028,N_8210);
xnor U13971 (N_13971,N_5882,N_7388);
nor U13972 (N_13972,N_9488,N_9124);
nor U13973 (N_13973,N_7437,N_5950);
and U13974 (N_13974,N_7881,N_9107);
nor U13975 (N_13975,N_8035,N_8057);
or U13976 (N_13976,N_6416,N_8137);
and U13977 (N_13977,N_7859,N_9575);
nand U13978 (N_13978,N_5770,N_6866);
and U13979 (N_13979,N_6630,N_9241);
nand U13980 (N_13980,N_6742,N_9880);
or U13981 (N_13981,N_5205,N_9730);
and U13982 (N_13982,N_5287,N_8480);
or U13983 (N_13983,N_7093,N_7143);
nor U13984 (N_13984,N_5796,N_6657);
and U13985 (N_13985,N_6539,N_7558);
or U13986 (N_13986,N_9888,N_5029);
and U13987 (N_13987,N_6680,N_5488);
nor U13988 (N_13988,N_9044,N_9352);
or U13989 (N_13989,N_6697,N_7769);
or U13990 (N_13990,N_5122,N_5551);
and U13991 (N_13991,N_6268,N_9335);
nor U13992 (N_13992,N_6129,N_7695);
nor U13993 (N_13993,N_8899,N_6287);
and U13994 (N_13994,N_8639,N_6248);
nor U13995 (N_13995,N_5450,N_9302);
nand U13996 (N_13996,N_8259,N_6519);
xor U13997 (N_13997,N_7398,N_6746);
xnor U13998 (N_13998,N_6816,N_6930);
nand U13999 (N_13999,N_8869,N_6212);
nand U14000 (N_14000,N_9436,N_7558);
xnor U14001 (N_14001,N_7637,N_6918);
and U14002 (N_14002,N_7813,N_5201);
nand U14003 (N_14003,N_5280,N_5966);
nand U14004 (N_14004,N_7226,N_6955);
xnor U14005 (N_14005,N_7442,N_6504);
nand U14006 (N_14006,N_5018,N_7513);
and U14007 (N_14007,N_8081,N_8357);
nor U14008 (N_14008,N_9178,N_7692);
and U14009 (N_14009,N_6858,N_6385);
xor U14010 (N_14010,N_9537,N_5455);
or U14011 (N_14011,N_6004,N_9925);
and U14012 (N_14012,N_5883,N_7881);
nand U14013 (N_14013,N_7919,N_7031);
or U14014 (N_14014,N_6193,N_9803);
or U14015 (N_14015,N_7668,N_8729);
nor U14016 (N_14016,N_8071,N_6938);
and U14017 (N_14017,N_7450,N_7185);
nor U14018 (N_14018,N_8311,N_9222);
nand U14019 (N_14019,N_9985,N_9413);
or U14020 (N_14020,N_5331,N_9153);
nor U14021 (N_14021,N_5664,N_9356);
and U14022 (N_14022,N_8847,N_6115);
xor U14023 (N_14023,N_9623,N_8161);
nor U14024 (N_14024,N_6015,N_9432);
nor U14025 (N_14025,N_5141,N_8234);
nand U14026 (N_14026,N_6000,N_6599);
and U14027 (N_14027,N_7571,N_7490);
nor U14028 (N_14028,N_9269,N_6699);
nand U14029 (N_14029,N_5355,N_8361);
nand U14030 (N_14030,N_5116,N_9471);
nand U14031 (N_14031,N_8241,N_7598);
nand U14032 (N_14032,N_7923,N_6206);
and U14033 (N_14033,N_7846,N_7653);
nand U14034 (N_14034,N_5344,N_7749);
nand U14035 (N_14035,N_5864,N_6034);
xor U14036 (N_14036,N_5087,N_6258);
nand U14037 (N_14037,N_8453,N_5309);
nor U14038 (N_14038,N_7877,N_6091);
nor U14039 (N_14039,N_8430,N_8449);
and U14040 (N_14040,N_9736,N_6917);
nor U14041 (N_14041,N_5024,N_5238);
xor U14042 (N_14042,N_8232,N_8393);
nand U14043 (N_14043,N_8059,N_8510);
xor U14044 (N_14044,N_8806,N_5399);
or U14045 (N_14045,N_5960,N_6820);
and U14046 (N_14046,N_7821,N_6580);
xnor U14047 (N_14047,N_9442,N_6171);
and U14048 (N_14048,N_9622,N_7156);
or U14049 (N_14049,N_9721,N_9567);
xnor U14050 (N_14050,N_5596,N_5969);
and U14051 (N_14051,N_5146,N_9318);
nor U14052 (N_14052,N_6479,N_6741);
nand U14053 (N_14053,N_7224,N_6301);
or U14054 (N_14054,N_7991,N_8800);
nor U14055 (N_14055,N_9279,N_9479);
nand U14056 (N_14056,N_9608,N_7664);
or U14057 (N_14057,N_9517,N_7060);
nand U14058 (N_14058,N_6358,N_7106);
nand U14059 (N_14059,N_8518,N_5069);
and U14060 (N_14060,N_5290,N_7702);
xnor U14061 (N_14061,N_7700,N_9750);
and U14062 (N_14062,N_7354,N_8259);
or U14063 (N_14063,N_8589,N_7979);
and U14064 (N_14064,N_7623,N_6014);
nor U14065 (N_14065,N_9065,N_5482);
or U14066 (N_14066,N_7391,N_5888);
nand U14067 (N_14067,N_9955,N_7763);
nand U14068 (N_14068,N_6189,N_6908);
nor U14069 (N_14069,N_7697,N_5547);
nor U14070 (N_14070,N_5066,N_7829);
nand U14071 (N_14071,N_9254,N_6361);
nor U14072 (N_14072,N_8689,N_5320);
and U14073 (N_14073,N_5503,N_7937);
nand U14074 (N_14074,N_8228,N_8071);
and U14075 (N_14075,N_9723,N_7544);
or U14076 (N_14076,N_7566,N_7016);
and U14077 (N_14077,N_5109,N_8525);
or U14078 (N_14078,N_9945,N_8154);
nand U14079 (N_14079,N_5226,N_9709);
nand U14080 (N_14080,N_9013,N_8853);
and U14081 (N_14081,N_6372,N_6556);
and U14082 (N_14082,N_9822,N_6705);
and U14083 (N_14083,N_7769,N_6163);
nor U14084 (N_14084,N_9835,N_9902);
nand U14085 (N_14085,N_8502,N_5555);
or U14086 (N_14086,N_5456,N_9337);
nand U14087 (N_14087,N_6310,N_6380);
or U14088 (N_14088,N_8533,N_7985);
xor U14089 (N_14089,N_5009,N_9402);
or U14090 (N_14090,N_8993,N_8759);
and U14091 (N_14091,N_9670,N_5872);
or U14092 (N_14092,N_6305,N_7168);
nand U14093 (N_14093,N_9712,N_7821);
or U14094 (N_14094,N_8359,N_8924);
xor U14095 (N_14095,N_5460,N_9666);
xnor U14096 (N_14096,N_9985,N_9560);
nor U14097 (N_14097,N_6836,N_7364);
or U14098 (N_14098,N_5998,N_9180);
nor U14099 (N_14099,N_8657,N_8952);
nand U14100 (N_14100,N_6710,N_6546);
and U14101 (N_14101,N_6370,N_8979);
or U14102 (N_14102,N_7097,N_7189);
nand U14103 (N_14103,N_5483,N_9222);
nand U14104 (N_14104,N_7237,N_7949);
or U14105 (N_14105,N_7003,N_6280);
nand U14106 (N_14106,N_9408,N_8871);
and U14107 (N_14107,N_5940,N_6897);
and U14108 (N_14108,N_5094,N_8763);
and U14109 (N_14109,N_6897,N_9932);
and U14110 (N_14110,N_5080,N_7794);
or U14111 (N_14111,N_6187,N_8200);
or U14112 (N_14112,N_7834,N_8402);
xor U14113 (N_14113,N_7854,N_8000);
nor U14114 (N_14114,N_6561,N_9893);
or U14115 (N_14115,N_8028,N_8773);
and U14116 (N_14116,N_7388,N_9966);
or U14117 (N_14117,N_5459,N_5254);
or U14118 (N_14118,N_7005,N_7453);
and U14119 (N_14119,N_5338,N_5744);
nor U14120 (N_14120,N_8548,N_8997);
or U14121 (N_14121,N_6540,N_9612);
nand U14122 (N_14122,N_5219,N_5666);
or U14123 (N_14123,N_7020,N_6692);
nand U14124 (N_14124,N_6452,N_7293);
and U14125 (N_14125,N_5251,N_7927);
or U14126 (N_14126,N_6563,N_5776);
nand U14127 (N_14127,N_5198,N_5606);
and U14128 (N_14128,N_9298,N_6449);
and U14129 (N_14129,N_7968,N_8520);
and U14130 (N_14130,N_9804,N_5463);
and U14131 (N_14131,N_5290,N_9709);
and U14132 (N_14132,N_8641,N_9708);
or U14133 (N_14133,N_5978,N_8734);
xor U14134 (N_14134,N_9228,N_7206);
nand U14135 (N_14135,N_9380,N_5870);
or U14136 (N_14136,N_8207,N_6608);
and U14137 (N_14137,N_9136,N_6201);
and U14138 (N_14138,N_7148,N_5192);
and U14139 (N_14139,N_7903,N_7581);
nor U14140 (N_14140,N_8093,N_5881);
nor U14141 (N_14141,N_7626,N_6735);
and U14142 (N_14142,N_9811,N_5360);
nand U14143 (N_14143,N_8210,N_5283);
nand U14144 (N_14144,N_6164,N_8093);
xnor U14145 (N_14145,N_9228,N_9924);
nand U14146 (N_14146,N_9404,N_7116);
and U14147 (N_14147,N_9892,N_9587);
or U14148 (N_14148,N_7906,N_8873);
and U14149 (N_14149,N_8862,N_9427);
nand U14150 (N_14150,N_5374,N_7103);
or U14151 (N_14151,N_5259,N_6804);
or U14152 (N_14152,N_7585,N_5771);
xnor U14153 (N_14153,N_5537,N_5840);
nor U14154 (N_14154,N_9060,N_7943);
and U14155 (N_14155,N_9319,N_6231);
or U14156 (N_14156,N_5930,N_5085);
and U14157 (N_14157,N_9843,N_6404);
nor U14158 (N_14158,N_5217,N_5042);
and U14159 (N_14159,N_5443,N_7242);
and U14160 (N_14160,N_7450,N_5920);
nor U14161 (N_14161,N_7279,N_7656);
xnor U14162 (N_14162,N_5975,N_9799);
or U14163 (N_14163,N_7889,N_5843);
xnor U14164 (N_14164,N_8829,N_9125);
nor U14165 (N_14165,N_6621,N_9476);
and U14166 (N_14166,N_5717,N_6119);
nor U14167 (N_14167,N_6368,N_8842);
or U14168 (N_14168,N_5320,N_6601);
nand U14169 (N_14169,N_8915,N_9705);
and U14170 (N_14170,N_6238,N_7404);
or U14171 (N_14171,N_9852,N_7628);
nor U14172 (N_14172,N_5274,N_8370);
nor U14173 (N_14173,N_7992,N_7915);
and U14174 (N_14174,N_8771,N_7890);
and U14175 (N_14175,N_5101,N_5215);
xor U14176 (N_14176,N_7818,N_5621);
and U14177 (N_14177,N_6371,N_9047);
nand U14178 (N_14178,N_8054,N_9894);
or U14179 (N_14179,N_6453,N_5441);
nand U14180 (N_14180,N_8333,N_6658);
nand U14181 (N_14181,N_9212,N_5218);
xor U14182 (N_14182,N_7331,N_9646);
nand U14183 (N_14183,N_5489,N_8970);
or U14184 (N_14184,N_6882,N_7748);
xor U14185 (N_14185,N_8297,N_5972);
or U14186 (N_14186,N_6453,N_9741);
nor U14187 (N_14187,N_9928,N_7827);
and U14188 (N_14188,N_6279,N_6946);
and U14189 (N_14189,N_7945,N_5993);
nand U14190 (N_14190,N_5700,N_5728);
xnor U14191 (N_14191,N_6319,N_8126);
nor U14192 (N_14192,N_6402,N_9626);
xnor U14193 (N_14193,N_7709,N_6401);
nor U14194 (N_14194,N_8793,N_8041);
nor U14195 (N_14195,N_9764,N_7161);
or U14196 (N_14196,N_8224,N_8326);
nand U14197 (N_14197,N_8025,N_8561);
or U14198 (N_14198,N_8053,N_7588);
nor U14199 (N_14199,N_6369,N_5500);
xor U14200 (N_14200,N_8191,N_6899);
xnor U14201 (N_14201,N_9537,N_6209);
or U14202 (N_14202,N_6124,N_8091);
or U14203 (N_14203,N_6328,N_8011);
nand U14204 (N_14204,N_8618,N_6184);
and U14205 (N_14205,N_9648,N_8195);
and U14206 (N_14206,N_9234,N_5985);
nor U14207 (N_14207,N_7046,N_7102);
nand U14208 (N_14208,N_5476,N_6718);
or U14209 (N_14209,N_6357,N_6902);
and U14210 (N_14210,N_9519,N_9675);
nand U14211 (N_14211,N_7973,N_8190);
nor U14212 (N_14212,N_5541,N_7305);
and U14213 (N_14213,N_7393,N_5699);
and U14214 (N_14214,N_7975,N_7055);
nor U14215 (N_14215,N_7318,N_8398);
nand U14216 (N_14216,N_5232,N_5089);
and U14217 (N_14217,N_7257,N_6083);
nand U14218 (N_14218,N_7870,N_6144);
nor U14219 (N_14219,N_7321,N_7543);
or U14220 (N_14220,N_6266,N_5793);
or U14221 (N_14221,N_6167,N_8185);
nand U14222 (N_14222,N_5311,N_7959);
nor U14223 (N_14223,N_7333,N_7014);
or U14224 (N_14224,N_8632,N_9246);
nand U14225 (N_14225,N_9583,N_9720);
and U14226 (N_14226,N_7438,N_5410);
xnor U14227 (N_14227,N_9519,N_9183);
or U14228 (N_14228,N_9633,N_6402);
and U14229 (N_14229,N_7611,N_9677);
nand U14230 (N_14230,N_6974,N_5331);
nand U14231 (N_14231,N_7624,N_8732);
nand U14232 (N_14232,N_5611,N_8327);
or U14233 (N_14233,N_5187,N_8424);
or U14234 (N_14234,N_5666,N_7737);
nor U14235 (N_14235,N_6102,N_6939);
nand U14236 (N_14236,N_6363,N_9083);
or U14237 (N_14237,N_5613,N_5080);
and U14238 (N_14238,N_6916,N_6305);
and U14239 (N_14239,N_5038,N_8862);
nand U14240 (N_14240,N_9317,N_9177);
nand U14241 (N_14241,N_9057,N_9604);
and U14242 (N_14242,N_7214,N_8443);
or U14243 (N_14243,N_5200,N_9402);
and U14244 (N_14244,N_6453,N_9962);
and U14245 (N_14245,N_5475,N_6203);
and U14246 (N_14246,N_7871,N_6465);
and U14247 (N_14247,N_5153,N_7071);
or U14248 (N_14248,N_7075,N_9024);
nand U14249 (N_14249,N_7107,N_8728);
nor U14250 (N_14250,N_8705,N_8601);
nand U14251 (N_14251,N_6654,N_6939);
nor U14252 (N_14252,N_8167,N_8148);
nor U14253 (N_14253,N_6438,N_6656);
nor U14254 (N_14254,N_9259,N_5418);
nor U14255 (N_14255,N_7446,N_5720);
and U14256 (N_14256,N_5722,N_9435);
xor U14257 (N_14257,N_8656,N_5871);
and U14258 (N_14258,N_5241,N_6935);
nor U14259 (N_14259,N_5768,N_8570);
nor U14260 (N_14260,N_9210,N_5935);
and U14261 (N_14261,N_5946,N_9783);
nand U14262 (N_14262,N_8079,N_5249);
or U14263 (N_14263,N_8770,N_7320);
nor U14264 (N_14264,N_6896,N_6636);
and U14265 (N_14265,N_8739,N_8924);
nand U14266 (N_14266,N_5566,N_8575);
or U14267 (N_14267,N_6190,N_6793);
and U14268 (N_14268,N_8973,N_6544);
and U14269 (N_14269,N_9344,N_7423);
or U14270 (N_14270,N_9775,N_7297);
and U14271 (N_14271,N_6086,N_6222);
nor U14272 (N_14272,N_8575,N_7669);
or U14273 (N_14273,N_6545,N_8321);
or U14274 (N_14274,N_8162,N_9402);
nor U14275 (N_14275,N_6351,N_7094);
xor U14276 (N_14276,N_9729,N_5932);
or U14277 (N_14277,N_8160,N_5415);
nand U14278 (N_14278,N_9913,N_8554);
or U14279 (N_14279,N_5900,N_7944);
and U14280 (N_14280,N_8369,N_7871);
or U14281 (N_14281,N_7905,N_9240);
nor U14282 (N_14282,N_7669,N_7395);
nand U14283 (N_14283,N_6118,N_6977);
and U14284 (N_14284,N_9378,N_9629);
nor U14285 (N_14285,N_5471,N_6928);
and U14286 (N_14286,N_6150,N_5543);
or U14287 (N_14287,N_8407,N_8886);
or U14288 (N_14288,N_8073,N_8396);
nand U14289 (N_14289,N_8492,N_9326);
nand U14290 (N_14290,N_9055,N_9844);
nor U14291 (N_14291,N_6503,N_5980);
nor U14292 (N_14292,N_5009,N_9610);
nand U14293 (N_14293,N_5795,N_6853);
xnor U14294 (N_14294,N_9656,N_8291);
xnor U14295 (N_14295,N_7258,N_7833);
and U14296 (N_14296,N_7983,N_9539);
nor U14297 (N_14297,N_7833,N_9473);
nand U14298 (N_14298,N_6542,N_9778);
or U14299 (N_14299,N_8048,N_8064);
nor U14300 (N_14300,N_8462,N_7377);
nand U14301 (N_14301,N_7816,N_5194);
and U14302 (N_14302,N_9517,N_6215);
and U14303 (N_14303,N_9408,N_6774);
nor U14304 (N_14304,N_5826,N_5685);
nand U14305 (N_14305,N_5925,N_8609);
or U14306 (N_14306,N_8776,N_5861);
and U14307 (N_14307,N_6084,N_9474);
or U14308 (N_14308,N_6970,N_7816);
nand U14309 (N_14309,N_7224,N_9399);
nand U14310 (N_14310,N_9706,N_7432);
nand U14311 (N_14311,N_8769,N_8612);
and U14312 (N_14312,N_5177,N_5769);
nand U14313 (N_14313,N_7727,N_7634);
or U14314 (N_14314,N_7793,N_9476);
nand U14315 (N_14315,N_9686,N_6279);
nor U14316 (N_14316,N_6427,N_8719);
nor U14317 (N_14317,N_7111,N_9076);
and U14318 (N_14318,N_6487,N_9283);
or U14319 (N_14319,N_7682,N_7860);
nand U14320 (N_14320,N_5700,N_9946);
and U14321 (N_14321,N_9903,N_5807);
and U14322 (N_14322,N_7877,N_8205);
nor U14323 (N_14323,N_9931,N_9144);
and U14324 (N_14324,N_7959,N_9585);
or U14325 (N_14325,N_6747,N_6104);
xnor U14326 (N_14326,N_5374,N_7241);
or U14327 (N_14327,N_6828,N_9542);
and U14328 (N_14328,N_7203,N_5014);
nor U14329 (N_14329,N_8613,N_9630);
or U14330 (N_14330,N_8657,N_7106);
or U14331 (N_14331,N_8073,N_5351);
and U14332 (N_14332,N_6936,N_7512);
nand U14333 (N_14333,N_7944,N_9825);
and U14334 (N_14334,N_6791,N_5488);
nand U14335 (N_14335,N_7796,N_6942);
and U14336 (N_14336,N_8888,N_9589);
nor U14337 (N_14337,N_9115,N_5560);
nor U14338 (N_14338,N_5431,N_5433);
nand U14339 (N_14339,N_7061,N_7081);
nand U14340 (N_14340,N_7427,N_5868);
nor U14341 (N_14341,N_7934,N_8265);
nor U14342 (N_14342,N_6001,N_7362);
and U14343 (N_14343,N_7646,N_5473);
nor U14344 (N_14344,N_7499,N_5417);
or U14345 (N_14345,N_7903,N_5012);
and U14346 (N_14346,N_6005,N_9827);
nor U14347 (N_14347,N_7404,N_9371);
nor U14348 (N_14348,N_7794,N_5741);
nor U14349 (N_14349,N_9210,N_5902);
or U14350 (N_14350,N_7696,N_9841);
nand U14351 (N_14351,N_8083,N_6571);
nand U14352 (N_14352,N_8050,N_8289);
nor U14353 (N_14353,N_5325,N_6159);
nor U14354 (N_14354,N_7135,N_7541);
or U14355 (N_14355,N_8267,N_8860);
or U14356 (N_14356,N_9284,N_5721);
and U14357 (N_14357,N_8874,N_8736);
nor U14358 (N_14358,N_5950,N_8411);
nand U14359 (N_14359,N_5004,N_8335);
nand U14360 (N_14360,N_6544,N_9659);
and U14361 (N_14361,N_9291,N_8709);
nor U14362 (N_14362,N_8938,N_6211);
xnor U14363 (N_14363,N_9394,N_8496);
nand U14364 (N_14364,N_6996,N_5312);
or U14365 (N_14365,N_7917,N_8183);
nor U14366 (N_14366,N_6449,N_7017);
nand U14367 (N_14367,N_6778,N_6600);
nor U14368 (N_14368,N_6379,N_5792);
and U14369 (N_14369,N_7588,N_6500);
nor U14370 (N_14370,N_5212,N_9607);
nor U14371 (N_14371,N_7126,N_7892);
nor U14372 (N_14372,N_6243,N_6829);
nand U14373 (N_14373,N_8743,N_5360);
and U14374 (N_14374,N_7441,N_9625);
or U14375 (N_14375,N_7799,N_9719);
or U14376 (N_14376,N_8346,N_8784);
or U14377 (N_14377,N_5281,N_5492);
nor U14378 (N_14378,N_7034,N_5760);
or U14379 (N_14379,N_6852,N_5251);
nor U14380 (N_14380,N_6151,N_9776);
nand U14381 (N_14381,N_5722,N_9100);
or U14382 (N_14382,N_9446,N_5466);
or U14383 (N_14383,N_6673,N_9496);
or U14384 (N_14384,N_6663,N_6072);
or U14385 (N_14385,N_8915,N_5918);
nor U14386 (N_14386,N_5627,N_7121);
or U14387 (N_14387,N_7722,N_9475);
nor U14388 (N_14388,N_9742,N_8338);
or U14389 (N_14389,N_6056,N_5373);
nor U14390 (N_14390,N_6008,N_5652);
or U14391 (N_14391,N_5082,N_5065);
nand U14392 (N_14392,N_9816,N_5590);
or U14393 (N_14393,N_9180,N_5819);
nand U14394 (N_14394,N_7450,N_8265);
and U14395 (N_14395,N_5428,N_5320);
nor U14396 (N_14396,N_7184,N_7462);
nand U14397 (N_14397,N_9625,N_5134);
and U14398 (N_14398,N_8490,N_7718);
or U14399 (N_14399,N_6177,N_9824);
and U14400 (N_14400,N_8487,N_9901);
and U14401 (N_14401,N_9136,N_7983);
xor U14402 (N_14402,N_5530,N_6509);
nor U14403 (N_14403,N_5876,N_8241);
nand U14404 (N_14404,N_7508,N_5959);
and U14405 (N_14405,N_8723,N_6977);
nor U14406 (N_14406,N_6254,N_5282);
and U14407 (N_14407,N_8501,N_8140);
nor U14408 (N_14408,N_6963,N_9415);
nand U14409 (N_14409,N_6747,N_8830);
xor U14410 (N_14410,N_8851,N_9012);
and U14411 (N_14411,N_7667,N_8315);
or U14412 (N_14412,N_7033,N_8448);
or U14413 (N_14413,N_9174,N_7460);
xor U14414 (N_14414,N_6935,N_5045);
or U14415 (N_14415,N_5405,N_6988);
nand U14416 (N_14416,N_9962,N_8975);
or U14417 (N_14417,N_8066,N_5361);
xnor U14418 (N_14418,N_7331,N_5777);
and U14419 (N_14419,N_6006,N_5159);
xor U14420 (N_14420,N_7782,N_6591);
nor U14421 (N_14421,N_9187,N_8949);
nor U14422 (N_14422,N_9003,N_6950);
nor U14423 (N_14423,N_5804,N_9573);
nand U14424 (N_14424,N_5115,N_5330);
nand U14425 (N_14425,N_9772,N_8722);
nand U14426 (N_14426,N_9617,N_6893);
nor U14427 (N_14427,N_8702,N_5718);
nor U14428 (N_14428,N_6061,N_6475);
nand U14429 (N_14429,N_6372,N_8490);
and U14430 (N_14430,N_7379,N_5754);
and U14431 (N_14431,N_6146,N_8811);
nor U14432 (N_14432,N_7907,N_9148);
and U14433 (N_14433,N_5859,N_7491);
and U14434 (N_14434,N_6579,N_6120);
or U14435 (N_14435,N_8467,N_6937);
and U14436 (N_14436,N_9771,N_8027);
or U14437 (N_14437,N_5163,N_8732);
or U14438 (N_14438,N_8307,N_6372);
nor U14439 (N_14439,N_9765,N_5021);
and U14440 (N_14440,N_9613,N_6203);
nor U14441 (N_14441,N_7789,N_6144);
xnor U14442 (N_14442,N_7480,N_8661);
or U14443 (N_14443,N_6332,N_9493);
nand U14444 (N_14444,N_8943,N_5596);
and U14445 (N_14445,N_7618,N_7980);
nor U14446 (N_14446,N_5373,N_5757);
nand U14447 (N_14447,N_7200,N_5431);
nand U14448 (N_14448,N_5977,N_6572);
nor U14449 (N_14449,N_9480,N_6660);
nand U14450 (N_14450,N_6957,N_9563);
nand U14451 (N_14451,N_6764,N_8241);
or U14452 (N_14452,N_6613,N_9239);
or U14453 (N_14453,N_9387,N_8016);
nor U14454 (N_14454,N_7905,N_5153);
or U14455 (N_14455,N_7976,N_7044);
xnor U14456 (N_14456,N_8171,N_8059);
xnor U14457 (N_14457,N_8976,N_8919);
nor U14458 (N_14458,N_5663,N_8288);
and U14459 (N_14459,N_9825,N_9334);
nor U14460 (N_14460,N_5129,N_5497);
nor U14461 (N_14461,N_7068,N_7156);
or U14462 (N_14462,N_5364,N_9283);
or U14463 (N_14463,N_6915,N_5829);
nor U14464 (N_14464,N_7025,N_7588);
or U14465 (N_14465,N_7765,N_9209);
and U14466 (N_14466,N_8201,N_8363);
or U14467 (N_14467,N_7624,N_8554);
or U14468 (N_14468,N_8329,N_5095);
nor U14469 (N_14469,N_8341,N_5682);
nand U14470 (N_14470,N_5740,N_6554);
or U14471 (N_14471,N_9027,N_9710);
nor U14472 (N_14472,N_5639,N_5672);
and U14473 (N_14473,N_8371,N_9799);
and U14474 (N_14474,N_5362,N_5032);
xor U14475 (N_14475,N_8201,N_6136);
nor U14476 (N_14476,N_5916,N_5751);
and U14477 (N_14477,N_9265,N_7384);
nand U14478 (N_14478,N_5778,N_9197);
xor U14479 (N_14479,N_6785,N_6269);
and U14480 (N_14480,N_8495,N_5957);
or U14481 (N_14481,N_8889,N_5151);
or U14482 (N_14482,N_6406,N_8776);
and U14483 (N_14483,N_7015,N_7868);
or U14484 (N_14484,N_5272,N_8979);
and U14485 (N_14485,N_8106,N_5341);
nor U14486 (N_14486,N_6052,N_6146);
nor U14487 (N_14487,N_6026,N_8375);
or U14488 (N_14488,N_7097,N_7221);
or U14489 (N_14489,N_7498,N_6633);
or U14490 (N_14490,N_5161,N_5174);
xnor U14491 (N_14491,N_7564,N_9698);
nand U14492 (N_14492,N_7242,N_6865);
nor U14493 (N_14493,N_5363,N_9440);
and U14494 (N_14494,N_5527,N_6126);
or U14495 (N_14495,N_5278,N_5565);
or U14496 (N_14496,N_9601,N_6430);
or U14497 (N_14497,N_9426,N_8765);
or U14498 (N_14498,N_6606,N_9597);
nand U14499 (N_14499,N_5641,N_7951);
xnor U14500 (N_14500,N_7070,N_7429);
and U14501 (N_14501,N_5540,N_5320);
nor U14502 (N_14502,N_8211,N_6920);
nand U14503 (N_14503,N_8058,N_7177);
or U14504 (N_14504,N_5311,N_8318);
nand U14505 (N_14505,N_8970,N_7156);
nor U14506 (N_14506,N_8191,N_6657);
and U14507 (N_14507,N_6048,N_5515);
nand U14508 (N_14508,N_7452,N_8561);
nand U14509 (N_14509,N_9895,N_6505);
nand U14510 (N_14510,N_6390,N_7748);
or U14511 (N_14511,N_5565,N_8899);
and U14512 (N_14512,N_6965,N_8932);
or U14513 (N_14513,N_8477,N_7001);
and U14514 (N_14514,N_8176,N_7866);
or U14515 (N_14515,N_8713,N_5907);
or U14516 (N_14516,N_8842,N_5533);
or U14517 (N_14517,N_5334,N_7418);
and U14518 (N_14518,N_6808,N_7443);
or U14519 (N_14519,N_9944,N_5129);
nand U14520 (N_14520,N_9455,N_8152);
or U14521 (N_14521,N_6328,N_9178);
or U14522 (N_14522,N_9937,N_5809);
and U14523 (N_14523,N_6676,N_5656);
nand U14524 (N_14524,N_8844,N_7036);
nand U14525 (N_14525,N_9425,N_5742);
or U14526 (N_14526,N_8485,N_8966);
nand U14527 (N_14527,N_8440,N_9373);
nand U14528 (N_14528,N_9939,N_7139);
and U14529 (N_14529,N_5286,N_7465);
nand U14530 (N_14530,N_8030,N_9031);
and U14531 (N_14531,N_9125,N_8045);
nor U14532 (N_14532,N_6998,N_5128);
and U14533 (N_14533,N_9955,N_6745);
and U14534 (N_14534,N_8829,N_8431);
nand U14535 (N_14535,N_5358,N_7431);
or U14536 (N_14536,N_8584,N_9422);
and U14537 (N_14537,N_7184,N_8704);
or U14538 (N_14538,N_5201,N_5831);
nand U14539 (N_14539,N_6559,N_9220);
nand U14540 (N_14540,N_8040,N_5407);
and U14541 (N_14541,N_9353,N_7108);
and U14542 (N_14542,N_7910,N_7590);
xor U14543 (N_14543,N_7382,N_7610);
and U14544 (N_14544,N_9720,N_9798);
xor U14545 (N_14545,N_6705,N_7310);
nor U14546 (N_14546,N_5020,N_8089);
xor U14547 (N_14547,N_7595,N_5674);
nor U14548 (N_14548,N_7753,N_5755);
xnor U14549 (N_14549,N_9418,N_9936);
nor U14550 (N_14550,N_5867,N_9905);
or U14551 (N_14551,N_7675,N_9429);
xor U14552 (N_14552,N_8422,N_9127);
xnor U14553 (N_14553,N_9444,N_6061);
nor U14554 (N_14554,N_8395,N_7331);
or U14555 (N_14555,N_6916,N_8240);
and U14556 (N_14556,N_5198,N_5239);
nor U14557 (N_14557,N_9478,N_8718);
nand U14558 (N_14558,N_9430,N_7610);
and U14559 (N_14559,N_6146,N_7746);
nand U14560 (N_14560,N_5785,N_7850);
and U14561 (N_14561,N_9122,N_7946);
and U14562 (N_14562,N_8675,N_7394);
xnor U14563 (N_14563,N_5009,N_5844);
nand U14564 (N_14564,N_8602,N_6744);
and U14565 (N_14565,N_6698,N_5271);
and U14566 (N_14566,N_5834,N_8541);
or U14567 (N_14567,N_9869,N_6573);
and U14568 (N_14568,N_6875,N_6830);
nand U14569 (N_14569,N_8255,N_6242);
nor U14570 (N_14570,N_9160,N_5637);
and U14571 (N_14571,N_9737,N_6876);
nor U14572 (N_14572,N_5475,N_9099);
xnor U14573 (N_14573,N_6024,N_7785);
nor U14574 (N_14574,N_7684,N_6361);
or U14575 (N_14575,N_8933,N_6933);
and U14576 (N_14576,N_8236,N_6372);
and U14577 (N_14577,N_5789,N_7919);
nand U14578 (N_14578,N_7867,N_5254);
nor U14579 (N_14579,N_9758,N_9116);
nand U14580 (N_14580,N_5461,N_8536);
nand U14581 (N_14581,N_5335,N_5345);
or U14582 (N_14582,N_8667,N_9949);
nor U14583 (N_14583,N_8935,N_9837);
and U14584 (N_14584,N_7460,N_5624);
or U14585 (N_14585,N_9860,N_7681);
and U14586 (N_14586,N_8702,N_8596);
or U14587 (N_14587,N_7406,N_8154);
xor U14588 (N_14588,N_9093,N_9794);
nand U14589 (N_14589,N_8313,N_9505);
or U14590 (N_14590,N_5061,N_8607);
or U14591 (N_14591,N_7559,N_9808);
nand U14592 (N_14592,N_9628,N_9958);
nand U14593 (N_14593,N_5640,N_8177);
and U14594 (N_14594,N_7109,N_9876);
nand U14595 (N_14595,N_9526,N_9632);
or U14596 (N_14596,N_9065,N_8657);
and U14597 (N_14597,N_6775,N_9993);
and U14598 (N_14598,N_5227,N_8741);
nor U14599 (N_14599,N_8178,N_7501);
nand U14600 (N_14600,N_8770,N_6667);
nand U14601 (N_14601,N_5012,N_8685);
and U14602 (N_14602,N_7049,N_6192);
and U14603 (N_14603,N_7267,N_6346);
nand U14604 (N_14604,N_6115,N_8554);
nor U14605 (N_14605,N_5418,N_7772);
nand U14606 (N_14606,N_8156,N_6361);
and U14607 (N_14607,N_6346,N_8734);
and U14608 (N_14608,N_6804,N_7648);
or U14609 (N_14609,N_7690,N_7934);
xor U14610 (N_14610,N_6808,N_6964);
and U14611 (N_14611,N_7750,N_5374);
or U14612 (N_14612,N_7196,N_7245);
nor U14613 (N_14613,N_8832,N_5519);
nand U14614 (N_14614,N_9351,N_7871);
xor U14615 (N_14615,N_6325,N_9097);
and U14616 (N_14616,N_9434,N_9588);
xor U14617 (N_14617,N_7233,N_5687);
nor U14618 (N_14618,N_6673,N_7119);
nor U14619 (N_14619,N_9097,N_7030);
or U14620 (N_14620,N_8121,N_6112);
and U14621 (N_14621,N_7130,N_7359);
nand U14622 (N_14622,N_9690,N_5613);
and U14623 (N_14623,N_8517,N_6183);
nor U14624 (N_14624,N_5753,N_9151);
xnor U14625 (N_14625,N_9499,N_5174);
or U14626 (N_14626,N_8037,N_9544);
or U14627 (N_14627,N_7783,N_7329);
and U14628 (N_14628,N_7907,N_7718);
nand U14629 (N_14629,N_5459,N_7474);
and U14630 (N_14630,N_6907,N_5548);
and U14631 (N_14631,N_8467,N_7666);
nand U14632 (N_14632,N_7335,N_6507);
or U14633 (N_14633,N_8747,N_6045);
nor U14634 (N_14634,N_7922,N_6716);
and U14635 (N_14635,N_6887,N_7171);
or U14636 (N_14636,N_8035,N_6762);
or U14637 (N_14637,N_5081,N_9250);
nor U14638 (N_14638,N_6246,N_6124);
and U14639 (N_14639,N_9144,N_8899);
nor U14640 (N_14640,N_7324,N_6748);
nand U14641 (N_14641,N_6776,N_6040);
nand U14642 (N_14642,N_7037,N_8799);
nand U14643 (N_14643,N_6834,N_5279);
or U14644 (N_14644,N_7328,N_7821);
nand U14645 (N_14645,N_7438,N_5028);
or U14646 (N_14646,N_9430,N_6850);
nand U14647 (N_14647,N_8478,N_6450);
nand U14648 (N_14648,N_6559,N_9939);
nand U14649 (N_14649,N_8792,N_7547);
xnor U14650 (N_14650,N_7442,N_7340);
or U14651 (N_14651,N_6699,N_5516);
and U14652 (N_14652,N_7794,N_6125);
and U14653 (N_14653,N_8603,N_9505);
nor U14654 (N_14654,N_7400,N_8151);
and U14655 (N_14655,N_5371,N_6877);
nand U14656 (N_14656,N_6282,N_6907);
and U14657 (N_14657,N_5201,N_6210);
and U14658 (N_14658,N_5501,N_5238);
and U14659 (N_14659,N_8077,N_5105);
nand U14660 (N_14660,N_8164,N_5287);
or U14661 (N_14661,N_5559,N_6646);
nand U14662 (N_14662,N_8559,N_6915);
nor U14663 (N_14663,N_9706,N_8146);
nand U14664 (N_14664,N_7268,N_8172);
xor U14665 (N_14665,N_5409,N_5949);
and U14666 (N_14666,N_6738,N_7991);
or U14667 (N_14667,N_9284,N_9584);
and U14668 (N_14668,N_7625,N_5729);
nor U14669 (N_14669,N_7095,N_9963);
nor U14670 (N_14670,N_7667,N_6910);
or U14671 (N_14671,N_7658,N_9445);
or U14672 (N_14672,N_9298,N_8914);
xnor U14673 (N_14673,N_5208,N_9345);
nor U14674 (N_14674,N_5069,N_7333);
and U14675 (N_14675,N_8513,N_5208);
nand U14676 (N_14676,N_6357,N_5465);
nor U14677 (N_14677,N_5247,N_7202);
nand U14678 (N_14678,N_5438,N_9546);
and U14679 (N_14679,N_7648,N_6592);
and U14680 (N_14680,N_7469,N_9655);
and U14681 (N_14681,N_5296,N_8226);
and U14682 (N_14682,N_6133,N_7480);
nor U14683 (N_14683,N_8387,N_5527);
nand U14684 (N_14684,N_5141,N_5820);
nand U14685 (N_14685,N_5496,N_7182);
or U14686 (N_14686,N_7601,N_9904);
nor U14687 (N_14687,N_9350,N_9287);
or U14688 (N_14688,N_8873,N_9259);
or U14689 (N_14689,N_8344,N_9739);
xor U14690 (N_14690,N_6261,N_6791);
nor U14691 (N_14691,N_5319,N_8967);
nor U14692 (N_14692,N_5571,N_5143);
nor U14693 (N_14693,N_5733,N_8493);
and U14694 (N_14694,N_6221,N_5631);
and U14695 (N_14695,N_9968,N_7013);
nor U14696 (N_14696,N_5825,N_6586);
or U14697 (N_14697,N_5362,N_8911);
nand U14698 (N_14698,N_7858,N_7145);
or U14699 (N_14699,N_9200,N_7711);
nand U14700 (N_14700,N_5865,N_7153);
or U14701 (N_14701,N_7885,N_6575);
nand U14702 (N_14702,N_7060,N_8295);
xor U14703 (N_14703,N_9948,N_9477);
or U14704 (N_14704,N_9916,N_8964);
or U14705 (N_14705,N_9302,N_7878);
and U14706 (N_14706,N_7650,N_9200);
or U14707 (N_14707,N_7958,N_6563);
nand U14708 (N_14708,N_5858,N_7804);
xor U14709 (N_14709,N_7884,N_5261);
and U14710 (N_14710,N_6693,N_9180);
or U14711 (N_14711,N_8683,N_9086);
and U14712 (N_14712,N_8411,N_5469);
and U14713 (N_14713,N_7963,N_6686);
or U14714 (N_14714,N_9234,N_5695);
nor U14715 (N_14715,N_6797,N_7901);
nand U14716 (N_14716,N_8166,N_8944);
and U14717 (N_14717,N_5218,N_8923);
nand U14718 (N_14718,N_5784,N_8396);
nand U14719 (N_14719,N_7393,N_9272);
nand U14720 (N_14720,N_8021,N_6831);
or U14721 (N_14721,N_5308,N_7415);
nor U14722 (N_14722,N_5763,N_5292);
xor U14723 (N_14723,N_6987,N_5798);
xor U14724 (N_14724,N_5889,N_6444);
nor U14725 (N_14725,N_6886,N_5431);
nor U14726 (N_14726,N_5383,N_5164);
or U14727 (N_14727,N_5368,N_8813);
nand U14728 (N_14728,N_8325,N_9999);
nor U14729 (N_14729,N_8365,N_6691);
nor U14730 (N_14730,N_6321,N_6219);
nand U14731 (N_14731,N_5983,N_8750);
xnor U14732 (N_14732,N_5352,N_6132);
and U14733 (N_14733,N_6125,N_6733);
nand U14734 (N_14734,N_7732,N_9081);
or U14735 (N_14735,N_5584,N_5876);
and U14736 (N_14736,N_6595,N_5713);
nand U14737 (N_14737,N_9058,N_5536);
nand U14738 (N_14738,N_9561,N_7388);
xor U14739 (N_14739,N_7644,N_6575);
and U14740 (N_14740,N_6003,N_6130);
nand U14741 (N_14741,N_7148,N_5942);
xor U14742 (N_14742,N_8508,N_5970);
and U14743 (N_14743,N_5250,N_6119);
xor U14744 (N_14744,N_8300,N_7789);
and U14745 (N_14745,N_5123,N_7749);
nand U14746 (N_14746,N_6706,N_6070);
or U14747 (N_14747,N_6622,N_7783);
nand U14748 (N_14748,N_9049,N_6251);
nand U14749 (N_14749,N_7316,N_9999);
nand U14750 (N_14750,N_5910,N_6765);
xnor U14751 (N_14751,N_6385,N_7483);
xor U14752 (N_14752,N_5263,N_9188);
nand U14753 (N_14753,N_7255,N_6223);
or U14754 (N_14754,N_5118,N_6675);
nand U14755 (N_14755,N_7043,N_5844);
nor U14756 (N_14756,N_5538,N_8535);
or U14757 (N_14757,N_7789,N_8153);
and U14758 (N_14758,N_8823,N_8957);
or U14759 (N_14759,N_9358,N_7285);
nand U14760 (N_14760,N_7500,N_8497);
nand U14761 (N_14761,N_6964,N_6698);
and U14762 (N_14762,N_7674,N_7865);
nand U14763 (N_14763,N_6450,N_6886);
nor U14764 (N_14764,N_7744,N_6248);
or U14765 (N_14765,N_8693,N_6693);
nor U14766 (N_14766,N_9220,N_6096);
nand U14767 (N_14767,N_9777,N_9352);
nand U14768 (N_14768,N_6131,N_6635);
nand U14769 (N_14769,N_7529,N_7223);
or U14770 (N_14770,N_7683,N_9866);
and U14771 (N_14771,N_5064,N_5471);
nor U14772 (N_14772,N_6714,N_8430);
nand U14773 (N_14773,N_9786,N_5273);
or U14774 (N_14774,N_7670,N_8542);
and U14775 (N_14775,N_6775,N_9291);
and U14776 (N_14776,N_7032,N_9044);
or U14777 (N_14777,N_5369,N_7656);
or U14778 (N_14778,N_9715,N_8941);
and U14779 (N_14779,N_6110,N_7607);
or U14780 (N_14780,N_5894,N_8481);
or U14781 (N_14781,N_9929,N_7956);
nor U14782 (N_14782,N_7895,N_8332);
and U14783 (N_14783,N_8216,N_9144);
and U14784 (N_14784,N_6252,N_6209);
nor U14785 (N_14785,N_6668,N_6556);
nor U14786 (N_14786,N_7287,N_9003);
nand U14787 (N_14787,N_6041,N_8054);
or U14788 (N_14788,N_8085,N_5943);
xnor U14789 (N_14789,N_9405,N_5396);
nand U14790 (N_14790,N_7966,N_5724);
or U14791 (N_14791,N_6343,N_8235);
and U14792 (N_14792,N_6628,N_9132);
or U14793 (N_14793,N_7512,N_9858);
and U14794 (N_14794,N_6337,N_7169);
nor U14795 (N_14795,N_8355,N_6647);
and U14796 (N_14796,N_6526,N_6019);
nor U14797 (N_14797,N_9277,N_6867);
or U14798 (N_14798,N_8023,N_9517);
and U14799 (N_14799,N_5565,N_7530);
nor U14800 (N_14800,N_5641,N_9199);
xor U14801 (N_14801,N_6821,N_5618);
xor U14802 (N_14802,N_7702,N_7565);
or U14803 (N_14803,N_5361,N_9803);
xor U14804 (N_14804,N_5861,N_6145);
or U14805 (N_14805,N_8187,N_9062);
and U14806 (N_14806,N_8489,N_9244);
or U14807 (N_14807,N_5080,N_7241);
or U14808 (N_14808,N_8039,N_5214);
or U14809 (N_14809,N_8728,N_6746);
and U14810 (N_14810,N_9390,N_6659);
nand U14811 (N_14811,N_7892,N_9087);
nor U14812 (N_14812,N_9890,N_5535);
nor U14813 (N_14813,N_6649,N_8827);
and U14814 (N_14814,N_5185,N_8632);
and U14815 (N_14815,N_5099,N_9473);
nor U14816 (N_14816,N_7406,N_5209);
and U14817 (N_14817,N_9085,N_6146);
and U14818 (N_14818,N_5693,N_8735);
or U14819 (N_14819,N_8883,N_5900);
nor U14820 (N_14820,N_8003,N_7161);
nand U14821 (N_14821,N_6136,N_5962);
or U14822 (N_14822,N_6377,N_7967);
nor U14823 (N_14823,N_6778,N_8356);
or U14824 (N_14824,N_8705,N_6942);
and U14825 (N_14825,N_8607,N_7774);
and U14826 (N_14826,N_5116,N_8736);
and U14827 (N_14827,N_6921,N_6964);
nand U14828 (N_14828,N_9820,N_8691);
or U14829 (N_14829,N_6628,N_9847);
nor U14830 (N_14830,N_9856,N_6548);
nor U14831 (N_14831,N_9658,N_8620);
and U14832 (N_14832,N_6353,N_6309);
nand U14833 (N_14833,N_8249,N_9777);
or U14834 (N_14834,N_9521,N_6167);
or U14835 (N_14835,N_8343,N_8928);
or U14836 (N_14836,N_9455,N_7718);
nor U14837 (N_14837,N_9291,N_5275);
nand U14838 (N_14838,N_9407,N_8467);
or U14839 (N_14839,N_5781,N_7928);
or U14840 (N_14840,N_5592,N_9784);
nor U14841 (N_14841,N_7677,N_5917);
xnor U14842 (N_14842,N_8719,N_6880);
and U14843 (N_14843,N_8868,N_6413);
and U14844 (N_14844,N_5989,N_5541);
and U14845 (N_14845,N_9960,N_8599);
or U14846 (N_14846,N_7242,N_6553);
nand U14847 (N_14847,N_5619,N_7492);
nand U14848 (N_14848,N_8455,N_9731);
nand U14849 (N_14849,N_9241,N_9647);
and U14850 (N_14850,N_5451,N_6120);
and U14851 (N_14851,N_6786,N_9058);
and U14852 (N_14852,N_5804,N_9845);
nor U14853 (N_14853,N_9149,N_6052);
or U14854 (N_14854,N_8825,N_9786);
nor U14855 (N_14855,N_6319,N_7978);
nand U14856 (N_14856,N_6960,N_5623);
nor U14857 (N_14857,N_5433,N_5824);
and U14858 (N_14858,N_9531,N_7212);
xnor U14859 (N_14859,N_5605,N_8943);
nand U14860 (N_14860,N_9438,N_8910);
nand U14861 (N_14861,N_5198,N_8604);
and U14862 (N_14862,N_6112,N_8021);
nand U14863 (N_14863,N_5608,N_7955);
nor U14864 (N_14864,N_7602,N_5779);
or U14865 (N_14865,N_7512,N_5344);
or U14866 (N_14866,N_6702,N_8787);
or U14867 (N_14867,N_6517,N_5671);
and U14868 (N_14868,N_5637,N_5145);
xor U14869 (N_14869,N_5806,N_8458);
nand U14870 (N_14870,N_5396,N_9770);
nor U14871 (N_14871,N_8500,N_7560);
nand U14872 (N_14872,N_8551,N_8558);
xnor U14873 (N_14873,N_7179,N_5053);
or U14874 (N_14874,N_7890,N_8522);
nor U14875 (N_14875,N_9848,N_6305);
nor U14876 (N_14876,N_9208,N_5699);
and U14877 (N_14877,N_6467,N_9827);
nand U14878 (N_14878,N_8597,N_5819);
nand U14879 (N_14879,N_8551,N_8650);
nand U14880 (N_14880,N_9190,N_6418);
nand U14881 (N_14881,N_5781,N_5581);
and U14882 (N_14882,N_8768,N_7682);
and U14883 (N_14883,N_7673,N_8357);
and U14884 (N_14884,N_8156,N_5744);
nor U14885 (N_14885,N_5168,N_5115);
nand U14886 (N_14886,N_9791,N_6464);
or U14887 (N_14887,N_5859,N_9794);
nand U14888 (N_14888,N_6206,N_8067);
or U14889 (N_14889,N_7244,N_7153);
or U14890 (N_14890,N_7090,N_6471);
and U14891 (N_14891,N_8660,N_8448);
nor U14892 (N_14892,N_7193,N_8902);
or U14893 (N_14893,N_6690,N_8807);
or U14894 (N_14894,N_6172,N_5722);
nor U14895 (N_14895,N_5912,N_8274);
or U14896 (N_14896,N_8502,N_7896);
nand U14897 (N_14897,N_9244,N_6162);
nor U14898 (N_14898,N_6582,N_8342);
nand U14899 (N_14899,N_7874,N_6731);
nand U14900 (N_14900,N_5458,N_7450);
xor U14901 (N_14901,N_8577,N_6125);
nand U14902 (N_14902,N_5148,N_6131);
nand U14903 (N_14903,N_8620,N_8191);
nor U14904 (N_14904,N_8683,N_8906);
nand U14905 (N_14905,N_5549,N_6615);
or U14906 (N_14906,N_5536,N_5466);
nand U14907 (N_14907,N_5471,N_6489);
and U14908 (N_14908,N_5581,N_6924);
and U14909 (N_14909,N_5032,N_6848);
and U14910 (N_14910,N_7996,N_9476);
nor U14911 (N_14911,N_5313,N_8388);
and U14912 (N_14912,N_8591,N_9911);
nor U14913 (N_14913,N_8771,N_5917);
or U14914 (N_14914,N_7561,N_9057);
xor U14915 (N_14915,N_8025,N_9541);
nor U14916 (N_14916,N_7436,N_8416);
and U14917 (N_14917,N_7261,N_8601);
and U14918 (N_14918,N_8657,N_5011);
or U14919 (N_14919,N_7100,N_5160);
nand U14920 (N_14920,N_8212,N_6455);
and U14921 (N_14921,N_8105,N_9593);
or U14922 (N_14922,N_8387,N_5046);
or U14923 (N_14923,N_5546,N_5574);
xnor U14924 (N_14924,N_9480,N_5931);
or U14925 (N_14925,N_5652,N_9284);
nand U14926 (N_14926,N_6800,N_6287);
and U14927 (N_14927,N_6691,N_6081);
nor U14928 (N_14928,N_5901,N_8297);
and U14929 (N_14929,N_9395,N_7852);
nand U14930 (N_14930,N_8074,N_7501);
and U14931 (N_14931,N_9509,N_6417);
nor U14932 (N_14932,N_8451,N_9786);
and U14933 (N_14933,N_5092,N_9918);
or U14934 (N_14934,N_5839,N_8260);
nand U14935 (N_14935,N_9770,N_5993);
nand U14936 (N_14936,N_7300,N_7453);
and U14937 (N_14937,N_9630,N_7472);
xnor U14938 (N_14938,N_9557,N_8899);
or U14939 (N_14939,N_8367,N_5028);
nor U14940 (N_14940,N_9660,N_8673);
nor U14941 (N_14941,N_9909,N_9783);
or U14942 (N_14942,N_9565,N_6634);
nand U14943 (N_14943,N_6321,N_8267);
nand U14944 (N_14944,N_6376,N_7282);
and U14945 (N_14945,N_5898,N_5473);
and U14946 (N_14946,N_9025,N_6324);
and U14947 (N_14947,N_9938,N_8346);
and U14948 (N_14948,N_9831,N_8097);
and U14949 (N_14949,N_6678,N_7150);
xnor U14950 (N_14950,N_7493,N_7635);
and U14951 (N_14951,N_7615,N_7541);
or U14952 (N_14952,N_8499,N_8692);
nor U14953 (N_14953,N_6068,N_6008);
nor U14954 (N_14954,N_7451,N_6791);
or U14955 (N_14955,N_8819,N_5012);
nor U14956 (N_14956,N_9970,N_8007);
nand U14957 (N_14957,N_5898,N_7831);
nand U14958 (N_14958,N_5947,N_7828);
and U14959 (N_14959,N_9865,N_6103);
nor U14960 (N_14960,N_7792,N_9431);
nand U14961 (N_14961,N_7792,N_8585);
or U14962 (N_14962,N_6784,N_7894);
nand U14963 (N_14963,N_9491,N_8640);
or U14964 (N_14964,N_8656,N_6656);
xor U14965 (N_14965,N_9746,N_7765);
and U14966 (N_14966,N_7426,N_6032);
or U14967 (N_14967,N_8653,N_5232);
nor U14968 (N_14968,N_8840,N_7438);
nor U14969 (N_14969,N_7527,N_9035);
or U14970 (N_14970,N_7665,N_8488);
and U14971 (N_14971,N_8184,N_9613);
or U14972 (N_14972,N_8125,N_8195);
xnor U14973 (N_14973,N_5266,N_7182);
nand U14974 (N_14974,N_8982,N_6286);
and U14975 (N_14975,N_5415,N_9713);
or U14976 (N_14976,N_6224,N_9386);
xor U14977 (N_14977,N_5918,N_8780);
nor U14978 (N_14978,N_8840,N_8393);
nand U14979 (N_14979,N_8831,N_8574);
nor U14980 (N_14980,N_8849,N_6388);
nand U14981 (N_14981,N_6696,N_9906);
or U14982 (N_14982,N_7238,N_9649);
xor U14983 (N_14983,N_5434,N_6830);
or U14984 (N_14984,N_9033,N_7650);
xnor U14985 (N_14985,N_7700,N_7547);
or U14986 (N_14986,N_6791,N_9582);
nor U14987 (N_14987,N_8784,N_7296);
nand U14988 (N_14988,N_7473,N_9288);
or U14989 (N_14989,N_5728,N_5498);
nand U14990 (N_14990,N_6459,N_7412);
nand U14991 (N_14991,N_6781,N_6068);
or U14992 (N_14992,N_9544,N_5135);
and U14993 (N_14993,N_9310,N_9674);
nand U14994 (N_14994,N_8018,N_7785);
nor U14995 (N_14995,N_6553,N_7795);
and U14996 (N_14996,N_6154,N_6562);
nor U14997 (N_14997,N_5330,N_7399);
nand U14998 (N_14998,N_6227,N_9464);
nor U14999 (N_14999,N_7236,N_5715);
or U15000 (N_15000,N_12916,N_13702);
nor U15001 (N_15001,N_12804,N_13810);
nand U15002 (N_15002,N_12920,N_10898);
and U15003 (N_15003,N_11871,N_14410);
nor U15004 (N_15004,N_12973,N_14103);
or U15005 (N_15005,N_12358,N_14953);
and U15006 (N_15006,N_10552,N_10750);
nor U15007 (N_15007,N_14077,N_14520);
or U15008 (N_15008,N_11611,N_13803);
nor U15009 (N_15009,N_11863,N_14177);
nand U15010 (N_15010,N_14459,N_10733);
and U15011 (N_15011,N_10369,N_14059);
or U15012 (N_15012,N_10061,N_13392);
or U15013 (N_15013,N_13209,N_12837);
nand U15014 (N_15014,N_10368,N_12775);
nor U15015 (N_15015,N_13764,N_11614);
and U15016 (N_15016,N_14833,N_14875);
and U15017 (N_15017,N_10423,N_13102);
nor U15018 (N_15018,N_12158,N_10753);
xor U15019 (N_15019,N_12546,N_10103);
or U15020 (N_15020,N_14386,N_12796);
or U15021 (N_15021,N_13233,N_12406);
nand U15022 (N_15022,N_14905,N_14295);
nand U15023 (N_15023,N_10667,N_12567);
nand U15024 (N_15024,N_14142,N_12516);
nor U15025 (N_15025,N_10772,N_13585);
nand U15026 (N_15026,N_12642,N_14268);
nor U15027 (N_15027,N_12093,N_13431);
nand U15028 (N_15028,N_14493,N_12986);
or U15029 (N_15029,N_14932,N_13680);
nor U15030 (N_15030,N_13313,N_11452);
or U15031 (N_15031,N_11372,N_11536);
or U15032 (N_15032,N_12416,N_12123);
nand U15033 (N_15033,N_10383,N_13359);
or U15034 (N_15034,N_12352,N_13440);
nand U15035 (N_15035,N_11719,N_13698);
nand U15036 (N_15036,N_14563,N_14720);
nand U15037 (N_15037,N_14117,N_14707);
nor U15038 (N_15038,N_11784,N_13593);
nor U15039 (N_15039,N_13166,N_11996);
nand U15040 (N_15040,N_13528,N_12253);
nand U15041 (N_15041,N_12731,N_13920);
or U15042 (N_15042,N_13616,N_10145);
nand U15043 (N_15043,N_12592,N_13965);
nand U15044 (N_15044,N_12934,N_12995);
and U15045 (N_15045,N_10946,N_12395);
nor U15046 (N_15046,N_11338,N_13605);
nor U15047 (N_15047,N_14831,N_11744);
nor U15048 (N_15048,N_10333,N_12559);
xnor U15049 (N_15049,N_12381,N_13922);
or U15050 (N_15050,N_13078,N_14682);
nand U15051 (N_15051,N_13257,N_13817);
nand U15052 (N_15052,N_11770,N_11115);
and U15053 (N_15053,N_11938,N_10764);
nor U15054 (N_15054,N_14503,N_14975);
nor U15055 (N_15055,N_12797,N_11028);
nand U15056 (N_15056,N_14791,N_11976);
nand U15057 (N_15057,N_10325,N_11239);
xor U15058 (N_15058,N_13406,N_13564);
nand U15059 (N_15059,N_10550,N_12952);
xnor U15060 (N_15060,N_10362,N_13594);
nor U15061 (N_15061,N_13513,N_11844);
nand U15062 (N_15062,N_10602,N_14065);
nor U15063 (N_15063,N_11812,N_10076);
and U15064 (N_15064,N_12700,N_10889);
and U15065 (N_15065,N_14502,N_10166);
nor U15066 (N_15066,N_14464,N_10332);
and U15067 (N_15067,N_14475,N_14613);
xnor U15068 (N_15068,N_14909,N_12247);
nand U15069 (N_15069,N_14958,N_11796);
or U15070 (N_15070,N_11586,N_10818);
nand U15071 (N_15071,N_14238,N_11691);
or U15072 (N_15072,N_13197,N_13608);
nor U15073 (N_15073,N_12023,N_14895);
and U15074 (N_15074,N_10460,N_14869);
or U15075 (N_15075,N_10807,N_13609);
nand U15076 (N_15076,N_10473,N_13100);
nand U15077 (N_15077,N_13548,N_13498);
nand U15078 (N_15078,N_14823,N_13047);
nand U15079 (N_15079,N_14190,N_12701);
nand U15080 (N_15080,N_11205,N_10715);
xor U15081 (N_15081,N_13301,N_13921);
and U15082 (N_15082,N_10371,N_13021);
xor U15083 (N_15083,N_10612,N_12538);
nor U15084 (N_15084,N_13410,N_13016);
nand U15085 (N_15085,N_10739,N_11663);
nand U15086 (N_15086,N_12122,N_13540);
nand U15087 (N_15087,N_12029,N_13270);
nand U15088 (N_15088,N_10238,N_12010);
nand U15089 (N_15089,N_14181,N_12765);
or U15090 (N_15090,N_13550,N_10420);
xnor U15091 (N_15091,N_11135,N_12204);
xnor U15092 (N_15092,N_14279,N_11179);
nor U15093 (N_15093,N_11085,N_13177);
or U15094 (N_15094,N_10707,N_11108);
xnor U15095 (N_15095,N_13829,N_11383);
or U15096 (N_15096,N_13806,N_12771);
nor U15097 (N_15097,N_13141,N_11072);
nor U15098 (N_15098,N_12981,N_14023);
and U15099 (N_15099,N_10669,N_13750);
xor U15100 (N_15100,N_12600,N_14094);
nor U15101 (N_15101,N_10598,N_14834);
nor U15102 (N_15102,N_10497,N_13252);
and U15103 (N_15103,N_13723,N_10948);
and U15104 (N_15104,N_11813,N_11762);
and U15105 (N_15105,N_13394,N_12280);
nand U15106 (N_15106,N_13751,N_10636);
nor U15107 (N_15107,N_12593,N_14830);
and U15108 (N_15108,N_13875,N_14818);
nor U15109 (N_15109,N_14570,N_13876);
and U15110 (N_15110,N_12457,N_14485);
or U15111 (N_15111,N_10815,N_13289);
and U15112 (N_15112,N_11106,N_14028);
and U15113 (N_15113,N_10915,N_13898);
xor U15114 (N_15114,N_14015,N_14242);
nand U15115 (N_15115,N_13891,N_11385);
xnor U15116 (N_15116,N_11349,N_11743);
nand U15117 (N_15117,N_12534,N_11170);
xor U15118 (N_15118,N_11978,N_10743);
or U15119 (N_15119,N_12794,N_12662);
and U15120 (N_15120,N_14110,N_13388);
nand U15121 (N_15121,N_11504,N_12954);
and U15122 (N_15122,N_14771,N_12484);
nor U15123 (N_15123,N_14797,N_13283);
nor U15124 (N_15124,N_11169,N_11622);
xor U15125 (N_15125,N_10248,N_12378);
nor U15126 (N_15126,N_12753,N_11080);
and U15127 (N_15127,N_11985,N_12800);
and U15128 (N_15128,N_12273,N_14221);
nor U15129 (N_15129,N_14335,N_11369);
nor U15130 (N_15130,N_11667,N_13588);
and U15131 (N_15131,N_13162,N_10846);
and U15132 (N_15132,N_12054,N_12186);
nand U15133 (N_15133,N_14179,N_14285);
nor U15134 (N_15134,N_11840,N_12555);
nand U15135 (N_15135,N_14385,N_11275);
and U15136 (N_15136,N_14135,N_10624);
or U15137 (N_15137,N_11470,N_10956);
or U15138 (N_15138,N_13692,N_11451);
nor U15139 (N_15139,N_13424,N_10949);
and U15140 (N_15140,N_11050,N_13816);
and U15141 (N_15141,N_14315,N_13995);
and U15142 (N_15142,N_11416,N_12919);
or U15143 (N_15143,N_13731,N_14750);
and U15144 (N_15144,N_12941,N_10126);
nor U15145 (N_15145,N_10806,N_11725);
or U15146 (N_15146,N_10731,N_11260);
xnor U15147 (N_15147,N_13774,N_11285);
xnor U15148 (N_15148,N_12754,N_11315);
nor U15149 (N_15149,N_10840,N_10400);
nand U15150 (N_15150,N_13826,N_13568);
nand U15151 (N_15151,N_14603,N_12821);
nor U15152 (N_15152,N_11103,N_13583);
nor U15153 (N_15153,N_11186,N_13142);
or U15154 (N_15154,N_13862,N_13469);
nand U15155 (N_15155,N_13989,N_13369);
and U15156 (N_15156,N_14164,N_12672);
nor U15157 (N_15157,N_11312,N_13940);
and U15158 (N_15158,N_11727,N_12887);
and U15159 (N_15159,N_13978,N_10802);
nand U15160 (N_15160,N_11419,N_11728);
or U15161 (N_15161,N_14388,N_14754);
nor U15162 (N_15162,N_11867,N_13835);
and U15163 (N_15163,N_11478,N_11534);
or U15164 (N_15164,N_12624,N_12831);
nor U15165 (N_15165,N_13587,N_11579);
nor U15166 (N_15166,N_10797,N_10107);
nand U15167 (N_15167,N_11776,N_10877);
or U15168 (N_15168,N_10466,N_10240);
nor U15169 (N_15169,N_11927,N_13353);
nand U15170 (N_15170,N_12177,N_12166);
nor U15171 (N_15171,N_14924,N_10077);
nor U15172 (N_15172,N_12570,N_11956);
nand U15173 (N_15173,N_12188,N_11032);
or U15174 (N_15174,N_13765,N_12854);
nand U15175 (N_15175,N_13178,N_10892);
and U15176 (N_15176,N_10385,N_11629);
nor U15177 (N_15177,N_10441,N_10099);
nand U15178 (N_15178,N_10523,N_13517);
nand U15179 (N_15179,N_11191,N_13506);
or U15180 (N_15180,N_11695,N_14524);
or U15181 (N_15181,N_10329,N_13983);
and U15182 (N_15182,N_12580,N_12793);
nand U15183 (N_15183,N_14546,N_14427);
or U15184 (N_15184,N_14558,N_10630);
and U15185 (N_15185,N_12152,N_13813);
xnor U15186 (N_15186,N_11301,N_10509);
nand U15187 (N_15187,N_14235,N_11146);
nand U15188 (N_15188,N_14165,N_11900);
or U15189 (N_15189,N_13733,N_11136);
or U15190 (N_15190,N_12888,N_12153);
xor U15191 (N_15191,N_13244,N_10520);
or U15192 (N_15192,N_12175,N_13012);
and U15193 (N_15193,N_10834,N_10457);
or U15194 (N_15194,N_12034,N_13944);
nand U15195 (N_15195,N_12875,N_12084);
nand U15196 (N_15196,N_12129,N_11559);
or U15197 (N_15197,N_10737,N_13542);
nor U15198 (N_15198,N_11111,N_10256);
and U15199 (N_15199,N_13781,N_11530);
and U15200 (N_15200,N_10983,N_14918);
and U15201 (N_15201,N_12865,N_10507);
xor U15202 (N_15202,N_11417,N_13055);
nor U15203 (N_15203,N_11401,N_14844);
and U15204 (N_15204,N_12703,N_10088);
and U15205 (N_15205,N_10249,N_11428);
nand U15206 (N_15206,N_10295,N_10012);
or U15207 (N_15207,N_14597,N_10535);
and U15208 (N_15208,N_10018,N_13734);
nand U15209 (N_15209,N_12761,N_12266);
nand U15210 (N_15210,N_14821,N_14945);
nand U15211 (N_15211,N_13551,N_10471);
or U15212 (N_15212,N_10866,N_12623);
or U15213 (N_15213,N_14217,N_14614);
nor U15214 (N_15214,N_10968,N_10283);
xnor U15215 (N_15215,N_10639,N_14031);
nand U15216 (N_15216,N_10578,N_11462);
nor U15217 (N_15217,N_13398,N_10851);
nor U15218 (N_15218,N_14726,N_12557);
nand U15219 (N_15219,N_14659,N_11858);
and U15220 (N_15220,N_10594,N_10773);
or U15221 (N_15221,N_10068,N_12150);
nor U15222 (N_15222,N_14311,N_13547);
and U15223 (N_15223,N_12808,N_13490);
nor U15224 (N_15224,N_11857,N_14532);
or U15225 (N_15225,N_14262,N_10048);
nand U15226 (N_15226,N_12597,N_10264);
nand U15227 (N_15227,N_13671,N_11198);
nand U15228 (N_15228,N_12673,N_14930);
nor U15229 (N_15229,N_14319,N_12544);
nor U15230 (N_15230,N_12383,N_12421);
and U15231 (N_15231,N_14215,N_10341);
nor U15232 (N_15232,N_13356,N_11522);
and U15233 (N_15233,N_11099,N_13138);
nand U15234 (N_15234,N_11658,N_10627);
and U15235 (N_15235,N_11873,N_13226);
or U15236 (N_15236,N_14965,N_12418);
and U15237 (N_15237,N_11351,N_10486);
nand U15238 (N_15238,N_14521,N_13526);
and U15239 (N_15239,N_12047,N_13673);
and U15240 (N_15240,N_13237,N_11003);
and U15241 (N_15241,N_11131,N_13215);
nand U15242 (N_15242,N_13465,N_14928);
or U15243 (N_15243,N_14974,N_14528);
nor U15244 (N_15244,N_12107,N_14606);
nand U15245 (N_15245,N_14740,N_10501);
nor U15246 (N_15246,N_11091,N_14798);
nand U15247 (N_15247,N_11196,N_14715);
and U15248 (N_15248,N_10318,N_10051);
and U15249 (N_15249,N_13699,N_10752);
or U15250 (N_15250,N_10290,N_10237);
nand U15251 (N_15251,N_10962,N_12869);
nor U15252 (N_15252,N_12721,N_12227);
nand U15253 (N_15253,N_14902,N_11688);
xnor U15254 (N_15254,N_13372,N_10830);
and U15255 (N_15255,N_13689,N_12246);
nand U15256 (N_15256,N_11690,N_12659);
nand U15257 (N_15257,N_10786,N_11891);
or U15258 (N_15258,N_12530,N_14397);
or U15259 (N_15259,N_13397,N_12776);
nor U15260 (N_15260,N_10440,N_13456);
or U15261 (N_15261,N_13326,N_11255);
and U15262 (N_15262,N_13874,N_12654);
or U15263 (N_15263,N_14363,N_11204);
nand U15264 (N_15264,N_11447,N_12684);
or U15265 (N_15265,N_11782,N_13620);
nand U15266 (N_15266,N_10175,N_11684);
nand U15267 (N_15267,N_11082,N_14991);
and U15268 (N_15268,N_14002,N_13163);
nor U15269 (N_15269,N_10601,N_14371);
nor U15270 (N_15270,N_10692,N_14781);
or U15271 (N_15271,N_11702,N_11811);
xor U15272 (N_15272,N_12782,N_12582);
or U15273 (N_15273,N_14938,N_11889);
nor U15274 (N_15274,N_11963,N_13277);
nor U15275 (N_15275,N_10093,N_10222);
or U15276 (N_15276,N_10364,N_11113);
or U15277 (N_15277,N_13943,N_10734);
and U15278 (N_15278,N_13098,N_12361);
xnor U15279 (N_15279,N_12543,N_11737);
and U15280 (N_15280,N_11547,N_11377);
and U15281 (N_15281,N_12250,N_11306);
or U15282 (N_15282,N_13837,N_11937);
nand U15283 (N_15283,N_10888,N_13065);
nand U15284 (N_15284,N_11843,N_13343);
or U15285 (N_15285,N_11642,N_10268);
nand U15286 (N_15286,N_13499,N_10749);
or U15287 (N_15287,N_14862,N_10589);
or U15288 (N_15288,N_14312,N_10309);
and U15289 (N_15289,N_12167,N_11414);
nor U15290 (N_15290,N_11537,N_12518);
or U15291 (N_15291,N_10990,N_12482);
xor U15292 (N_15292,N_13436,N_14592);
xnor U15293 (N_15293,N_14583,N_11760);
nand U15294 (N_15294,N_10174,N_12252);
nand U15295 (N_15295,N_13648,N_12602);
or U15296 (N_15296,N_10035,N_11914);
nor U15297 (N_15297,N_10540,N_13981);
nand U15298 (N_15298,N_13555,N_12675);
nor U15299 (N_15299,N_12090,N_14741);
nor U15300 (N_15300,N_14112,N_11183);
xor U15301 (N_15301,N_14073,N_10817);
and U15302 (N_15302,N_10875,N_11321);
nor U15303 (N_15303,N_12350,N_10482);
nand U15304 (N_15304,N_10695,N_10262);
nand U15305 (N_15305,N_13064,N_14751);
nand U15306 (N_15306,N_13076,N_10529);
and U15307 (N_15307,N_13766,N_10156);
or U15308 (N_15308,N_10849,N_13683);
nor U15309 (N_15309,N_10814,N_10542);
and U15310 (N_15310,N_11201,N_12314);
or U15311 (N_15311,N_12898,N_12044);
and U15312 (N_15312,N_13953,N_10213);
nor U15313 (N_15313,N_12211,N_11977);
or U15314 (N_15314,N_10186,N_12907);
or U15315 (N_15315,N_13979,N_14555);
xor U15316 (N_15316,N_11326,N_12131);
nand U15317 (N_15317,N_13948,N_11550);
nor U15318 (N_15318,N_11849,N_14591);
nor U15319 (N_15319,N_12610,N_11793);
nand U15320 (N_15320,N_10785,N_12665);
and U15321 (N_15321,N_13621,N_14430);
nand U15322 (N_15322,N_14208,N_11124);
or U15323 (N_15323,N_13808,N_12994);
or U15324 (N_15324,N_11410,N_11680);
or U15325 (N_15325,N_13366,N_10719);
and U15326 (N_15326,N_12181,N_11525);
and U15327 (N_15327,N_11772,N_13515);
nor U15328 (N_15328,N_13224,N_13463);
nor U15329 (N_15329,N_11731,N_10910);
and U15330 (N_15330,N_14318,N_12363);
and U15331 (N_15331,N_14403,N_11778);
xor U15332 (N_15332,N_14025,N_12144);
nand U15333 (N_15333,N_13668,N_13095);
nand U15334 (N_15334,N_13002,N_13543);
nand U15335 (N_15335,N_12539,N_11049);
nand U15336 (N_15336,N_13791,N_11546);
nor U15337 (N_15337,N_10592,N_10660);
nor U15338 (N_15338,N_14894,N_10472);
nand U15339 (N_15339,N_14661,N_12850);
or U15340 (N_15340,N_11999,N_12730);
or U15341 (N_15341,N_10299,N_14137);
or U15342 (N_15342,N_13273,N_14647);
or U15343 (N_15343,N_14738,N_12745);
or U15344 (N_15344,N_11519,N_10958);
nand U15345 (N_15345,N_11258,N_11804);
nor U15346 (N_15346,N_12588,N_10326);
or U15347 (N_15347,N_10885,N_14163);
nor U15348 (N_15348,N_12005,N_13975);
nand U15349 (N_15349,N_11521,N_11502);
xnor U15350 (N_15350,N_14589,N_11624);
and U15351 (N_15351,N_10841,N_14406);
nand U15352 (N_15352,N_11398,N_11162);
and U15353 (N_15353,N_12022,N_14899);
nor U15354 (N_15354,N_10596,N_10146);
nor U15355 (N_15355,N_11267,N_10928);
xnor U15356 (N_15356,N_11141,N_14944);
and U15357 (N_15357,N_12728,N_11304);
or U15358 (N_15358,N_13715,N_14625);
nand U15359 (N_15359,N_12976,N_14541);
nor U15360 (N_15360,N_10223,N_14799);
nand U15361 (N_15361,N_11668,N_14472);
nand U15362 (N_15362,N_14256,N_12750);
nor U15363 (N_15363,N_11545,N_10813);
nand U15364 (N_15364,N_11700,N_11669);
or U15365 (N_15365,N_13425,N_10997);
and U15366 (N_15366,N_10470,N_11166);
and U15367 (N_15367,N_11942,N_11666);
and U15368 (N_15368,N_14193,N_13763);
or U15369 (N_15369,N_11472,N_11563);
nand U15370 (N_15370,N_11202,N_14153);
nand U15371 (N_15371,N_11588,N_14402);
or U15372 (N_15372,N_12709,N_11792);
nor U15373 (N_15373,N_10285,N_12851);
nand U15374 (N_15374,N_11216,N_10409);
and U15375 (N_15375,N_12717,N_10679);
nor U15376 (N_15376,N_13822,N_14843);
nor U15377 (N_15377,N_12359,N_14828);
nand U15378 (N_15378,N_14340,N_12064);
nand U15379 (N_15379,N_13558,N_12112);
and U15380 (N_15380,N_11043,N_13576);
or U15381 (N_15381,N_13007,N_13591);
or U15382 (N_15382,N_14617,N_13112);
and U15383 (N_15383,N_13695,N_12748);
or U15384 (N_15384,N_12053,N_10393);
nand U15385 (N_15385,N_10573,N_11568);
xor U15386 (N_15386,N_10190,N_11980);
and U15387 (N_15387,N_12103,N_11655);
xor U15388 (N_15388,N_14616,N_14205);
xor U15389 (N_15389,N_13081,N_14483);
nand U15390 (N_15390,N_11151,N_10780);
nor U15391 (N_15391,N_10908,N_10343);
xor U15392 (N_15392,N_10685,N_10887);
nor U15393 (N_15393,N_13537,N_13453);
xor U15394 (N_15394,N_10407,N_13416);
nor U15395 (N_15395,N_10917,N_12269);
nand U15396 (N_15396,N_10244,N_13139);
nand U15397 (N_15397,N_13200,N_14228);
nor U15398 (N_15398,N_11697,N_13900);
and U15399 (N_15399,N_12162,N_13861);
nand U15400 (N_15400,N_13871,N_11987);
nand U15401 (N_15401,N_14452,N_14444);
and U15402 (N_15402,N_14784,N_14016);
or U15403 (N_15403,N_10419,N_11748);
nor U15404 (N_15404,N_13522,N_10622);
nor U15405 (N_15405,N_11011,N_14687);
nand U15406 (N_15406,N_11030,N_14789);
and U15407 (N_15407,N_12724,N_13739);
and U15408 (N_15408,N_12468,N_12220);
and U15409 (N_15409,N_12500,N_10706);
and U15410 (N_15410,N_13208,N_14013);
nor U15411 (N_15411,N_11223,N_12294);
nand U15412 (N_15412,N_13128,N_13386);
and U15413 (N_15413,N_12943,N_14018);
nor U15414 (N_15414,N_14087,N_13033);
or U15415 (N_15415,N_10004,N_14681);
nor U15416 (N_15416,N_11562,N_11088);
nor U15417 (N_15417,N_13685,N_14816);
or U15418 (N_15418,N_13667,N_13529);
nand U15419 (N_15419,N_13061,N_12649);
nor U15420 (N_15420,N_11592,N_11484);
and U15421 (N_15421,N_11694,N_12531);
and U15422 (N_15422,N_12276,N_12692);
and U15423 (N_15423,N_13996,N_11104);
nand U15424 (N_15424,N_12806,N_12075);
nor U15425 (N_15425,N_10163,N_13134);
nand U15426 (N_15426,N_13470,N_10454);
xor U15427 (N_15427,N_13484,N_12407);
nor U15428 (N_15428,N_11286,N_11848);
and U15429 (N_15429,N_12141,N_14936);
nand U15430 (N_15430,N_11047,N_14979);
xnor U15431 (N_15431,N_13473,N_11715);
nor U15432 (N_15432,N_11529,N_13236);
or U15433 (N_15433,N_10561,N_12392);
and U15434 (N_15434,N_11635,N_13973);
and U15435 (N_15435,N_14382,N_14404);
nand U15436 (N_15436,N_11826,N_14694);
nor U15437 (N_15437,N_11459,N_11660);
or U15438 (N_15438,N_11145,N_12763);
nand U15439 (N_15439,N_11872,N_11855);
and U15440 (N_15440,N_12296,N_10297);
nand U15441 (N_15441,N_14511,N_10425);
or U15442 (N_15442,N_10778,N_14904);
or U15443 (N_15443,N_14693,N_11167);
nor U15444 (N_15444,N_10006,N_10179);
nor U15445 (N_15445,N_14166,N_10744);
and U15446 (N_15446,N_11945,N_14516);
and U15447 (N_15447,N_10476,N_10762);
xnor U15448 (N_15448,N_11965,N_14032);
nor U15449 (N_15449,N_14739,N_13881);
and U15450 (N_15450,N_13486,N_14674);
or U15451 (N_15451,N_11064,N_10923);
and U15452 (N_15452,N_14450,N_11653);
or U15453 (N_15453,N_11055,N_10090);
nor U15454 (N_15454,N_12671,N_12133);
or U15455 (N_15455,N_11314,N_11387);
or U15456 (N_15456,N_14539,N_14728);
and U15457 (N_15457,N_14272,N_10097);
nand U15458 (N_15458,N_14253,N_12825);
nand U15459 (N_15459,N_12680,N_13815);
or U15460 (N_15460,N_13274,N_10347);
nand U15461 (N_15461,N_14229,N_14615);
xnor U15462 (N_15462,N_14586,N_13253);
and U15463 (N_15463,N_11226,N_13909);
and U15464 (N_15464,N_14239,N_12801);
nor U15465 (N_15465,N_12982,N_13193);
and U15466 (N_15466,N_11445,N_13084);
or U15467 (N_15467,N_14527,N_11422);
nand U15468 (N_15468,N_14961,N_14246);
nor U15469 (N_15469,N_13120,N_11723);
and U15470 (N_15470,N_12494,N_10953);
nand U15471 (N_15471,N_14759,N_14811);
nand U15472 (N_15472,N_13746,N_14994);
or U15473 (N_15473,N_11676,N_12751);
nor U15474 (N_15474,N_12959,N_10714);
and U15475 (N_15475,N_10172,N_10634);
xnor U15476 (N_15476,N_10867,N_14220);
nand U15477 (N_15477,N_14841,N_12423);
xor U15478 (N_15478,N_14884,N_14897);
nand U15479 (N_15479,N_10835,N_13612);
nand U15480 (N_15480,N_14986,N_11625);
or U15481 (N_15481,N_10137,N_12562);
nand U15482 (N_15482,N_11902,N_11059);
or U15483 (N_15483,N_10129,N_14438);
or U15484 (N_15484,N_13468,N_10979);
or U15485 (N_15485,N_10502,N_10847);
and U15486 (N_15486,N_14775,N_12503);
or U15487 (N_15487,N_14443,N_12370);
nand U15488 (N_15488,N_11297,N_10965);
xor U15489 (N_15489,N_12304,N_12702);
or U15490 (N_15490,N_13234,N_14104);
nand U15491 (N_15491,N_14982,N_14927);
nand U15492 (N_15492,N_11037,N_11527);
and U15493 (N_15493,N_12931,N_10996);
xor U15494 (N_15494,N_14251,N_14805);
or U15495 (N_15495,N_14413,N_12430);
nor U15496 (N_15496,N_12611,N_13866);
nand U15497 (N_15497,N_10683,N_14736);
or U15498 (N_15498,N_14676,N_10865);
or U15499 (N_15499,N_13483,N_10581);
and U15500 (N_15500,N_10620,N_14960);
xor U15501 (N_15501,N_12146,N_14442);
nand U15502 (N_15502,N_12891,N_12573);
xnor U15503 (N_15503,N_13938,N_14298);
nor U15504 (N_15504,N_10494,N_10618);
nand U15505 (N_15505,N_14287,N_14180);
and U15506 (N_15506,N_11777,N_13319);
and U15507 (N_15507,N_14892,N_14639);
xor U15508 (N_15508,N_14425,N_13172);
nand U15509 (N_15509,N_11986,N_11988);
and U15510 (N_15510,N_13851,N_13652);
nor U15511 (N_15511,N_13789,N_13503);
or U15512 (N_15512,N_13895,N_12087);
nand U15513 (N_15513,N_11160,N_10666);
nor U15514 (N_15514,N_10593,N_13005);
or U15515 (N_15515,N_14230,N_12061);
nand U15516 (N_15516,N_13085,N_10989);
nor U15517 (N_15517,N_11069,N_13291);
xor U15518 (N_15518,N_12527,N_10652);
nand U15519 (N_15519,N_14602,N_11325);
nor U15520 (N_15520,N_14412,N_11973);
nor U15521 (N_15521,N_11802,N_13014);
nand U15522 (N_15522,N_13083,N_12130);
nor U15523 (N_15523,N_11294,N_14522);
xnor U15524 (N_15524,N_13176,N_14192);
nand U15525 (N_15525,N_11713,N_13454);
nand U15526 (N_15526,N_11117,N_11931);
nand U15527 (N_15527,N_14695,N_13097);
and U15528 (N_15528,N_10196,N_11841);
and U15529 (N_15529,N_10049,N_14317);
xor U15530 (N_15530,N_13164,N_10100);
and U15531 (N_15531,N_12605,N_10243);
xor U15532 (N_15532,N_10522,N_14236);
xnor U15533 (N_15533,N_11954,N_12293);
or U15534 (N_15534,N_13328,N_13525);
or U15535 (N_15535,N_13057,N_10247);
or U15536 (N_15536,N_13309,N_11820);
and U15537 (N_15537,N_10736,N_14313);
nor U15538 (N_15538,N_13906,N_14118);
and U15539 (N_15539,N_14632,N_10200);
nor U15540 (N_15540,N_14574,N_13778);
or U15541 (N_15541,N_14326,N_11153);
and U15542 (N_15542,N_10763,N_12996);
xnor U15543 (N_15543,N_13022,N_11610);
nor U15544 (N_15544,N_14568,N_10735);
nand U15545 (N_15545,N_14601,N_11704);
nor U15546 (N_15546,N_12414,N_10907);
nor U15547 (N_15547,N_14610,N_10113);
or U15548 (N_15548,N_10199,N_14124);
xnor U15549 (N_15549,N_12125,N_10217);
or U15550 (N_15550,N_10884,N_13256);
nand U15551 (N_15551,N_12584,N_14301);
or U15552 (N_15552,N_11184,N_11121);
nor U15553 (N_15553,N_12532,N_11075);
nor U15554 (N_15554,N_12848,N_13000);
nand U15555 (N_15555,N_10862,N_10526);
nand U15556 (N_15556,N_11359,N_13074);
nor U15557 (N_15557,N_13316,N_10779);
xor U15558 (N_15558,N_10135,N_12553);
or U15559 (N_15559,N_10165,N_13240);
nor U15560 (N_15560,N_12290,N_12741);
and U15561 (N_15561,N_12343,N_10022);
or U15562 (N_15562,N_13346,N_10389);
and U15563 (N_15563,N_14379,N_12020);
nand U15564 (N_15564,N_14045,N_12102);
nor U15565 (N_15565,N_14453,N_14972);
nor U15566 (N_15566,N_13170,N_12758);
nor U15567 (N_15567,N_12085,N_11982);
or U15568 (N_15568,N_11701,N_12161);
and U15569 (N_15569,N_11555,N_13939);
and U15570 (N_15570,N_10663,N_10748);
and U15571 (N_15571,N_14063,N_10251);
nand U15572 (N_15572,N_11433,N_12729);
nor U15573 (N_15573,N_10798,N_14030);
or U15574 (N_15574,N_10294,N_14393);
or U15575 (N_15575,N_10260,N_11180);
or U15576 (N_15576,N_11495,N_13839);
nand U15577 (N_15577,N_13205,N_10205);
and U15578 (N_15578,N_12134,N_10911);
or U15579 (N_15579,N_10906,N_13415);
xor U15580 (N_15580,N_11287,N_11094);
and U15581 (N_15581,N_11950,N_12802);
or U15582 (N_15582,N_12393,N_13444);
nor U15583 (N_15583,N_10081,N_14992);
and U15584 (N_15584,N_14766,N_11218);
xor U15585 (N_15585,N_14121,N_12055);
nand U15586 (N_15586,N_11961,N_12657);
and U15587 (N_15587,N_10690,N_11974);
or U15588 (N_15588,N_10342,N_10653);
nand U15589 (N_15589,N_14552,N_10599);
nand U15590 (N_15590,N_14874,N_10373);
nand U15591 (N_15591,N_13155,N_13282);
nand U15592 (N_15592,N_12045,N_14569);
nor U15593 (N_15593,N_11152,N_10929);
nand U15594 (N_15594,N_10276,N_14641);
nand U15595 (N_15595,N_14489,N_12194);
nand U15596 (N_15596,N_11161,N_14173);
or U15597 (N_15597,N_12501,N_13717);
nor U15598 (N_15598,N_13811,N_11118);
and U15599 (N_15599,N_12510,N_14649);
nor U15600 (N_15600,N_10269,N_13538);
nand U15601 (N_15601,N_10991,N_13242);
and U15602 (N_15602,N_10073,N_14638);
nand U15603 (N_15603,N_12958,N_12024);
nor U15604 (N_15604,N_14501,N_12226);
nor U15605 (N_15605,N_11157,N_12576);
or U15606 (N_15606,N_12424,N_10582);
and U15607 (N_15607,N_13455,N_11021);
and U15608 (N_15608,N_14596,N_12988);
nor U15609 (N_15609,N_13009,N_10859);
xnor U15610 (N_15610,N_12128,N_12645);
xnor U15611 (N_15611,N_13625,N_13669);
nand U15612 (N_15612,N_13131,N_12245);
nand U15613 (N_15613,N_10607,N_11042);
nor U15614 (N_15614,N_10032,N_14545);
nand U15615 (N_15615,N_12136,N_13570);
nand U15616 (N_15616,N_12279,N_10350);
nand U15617 (N_15617,N_13091,N_11946);
nand U15618 (N_15618,N_14530,N_13044);
or U15619 (N_15619,N_14291,N_12078);
or U15620 (N_15620,N_12324,N_10795);
xnor U15621 (N_15621,N_13169,N_10994);
xnor U15622 (N_15622,N_13559,N_10033);
xor U15623 (N_15623,N_13694,N_11120);
and U15624 (N_15624,N_13451,N_11716);
and U15625 (N_15625,N_11262,N_11320);
nor U15626 (N_15626,N_14700,N_14162);
nor U15627 (N_15627,N_11324,N_10136);
nor U15628 (N_15628,N_10754,N_13660);
and U15629 (N_15629,N_13367,N_14713);
and U15630 (N_15630,N_13927,N_10345);
or U15631 (N_15631,N_14009,N_14624);
nand U15632 (N_15632,N_11573,N_11541);
xnor U15633 (N_15633,N_10632,N_14692);
nor U15634 (N_15634,N_14551,N_11040);
and U15635 (N_15635,N_12864,N_11966);
nand U15636 (N_15636,N_10919,N_12617);
nor U15637 (N_15637,N_11925,N_10431);
or U15638 (N_15638,N_12953,N_11093);
or U15639 (N_15639,N_11019,N_12036);
xnor U15640 (N_15640,N_14499,N_10209);
nor U15641 (N_15641,N_11808,N_10822);
and U15642 (N_15642,N_10610,N_13028);
and U15643 (N_15643,N_10278,N_11698);
or U15644 (N_15644,N_13883,N_10459);
nor U15645 (N_15645,N_11584,N_13776);
nor U15646 (N_15646,N_13032,N_10864);
or U15647 (N_15647,N_10487,N_10360);
nor U15648 (N_15648,N_14881,N_11430);
nand U15649 (N_15649,N_11063,N_10936);
nor U15650 (N_15650,N_14108,N_14196);
and U15651 (N_15651,N_10788,N_12376);
and U15652 (N_15652,N_10918,N_11076);
nand U15653 (N_15653,N_12372,N_14926);
xnor U15654 (N_15654,N_13168,N_11269);
nor U15655 (N_15655,N_10204,N_14648);
xor U15656 (N_15656,N_14222,N_11879);
nor U15657 (N_15657,N_13510,N_11006);
or U15658 (N_15658,N_13382,N_13935);
and U15659 (N_15659,N_14353,N_12714);
nor U15660 (N_15660,N_14640,N_12639);
or U15661 (N_15661,N_12690,N_10571);
or U15662 (N_15662,N_12799,N_13575);
or U15663 (N_15663,N_10484,N_14361);
nand U15664 (N_15664,N_11060,N_14460);
nor U15665 (N_15665,N_11752,N_10852);
nand U15666 (N_15666,N_14915,N_12096);
or U15667 (N_15667,N_10128,N_12051);
and U15668 (N_15668,N_14174,N_12968);
nor U15669 (N_15669,N_13719,N_13914);
nand U15670 (N_15670,N_13872,N_12525);
xnor U15671 (N_15671,N_14655,N_13655);
nand U15672 (N_15672,N_10316,N_10547);
nand U15673 (N_15673,N_13565,N_11257);
nand U15674 (N_15674,N_11865,N_11730);
or U15675 (N_15675,N_10930,N_11307);
nor U15676 (N_15676,N_11847,N_13725);
and U15677 (N_15677,N_13650,N_12732);
and U15678 (N_15678,N_10207,N_10434);
or U15679 (N_15679,N_12322,N_12619);
xnor U15680 (N_15680,N_11092,N_14396);
nor U15681 (N_15681,N_13630,N_14167);
or U15682 (N_15682,N_12676,N_10397);
xor U15683 (N_15683,N_12081,N_14814);
and U15684 (N_15684,N_12990,N_12083);
or U15685 (N_15685,N_10686,N_13846);
nor U15686 (N_15686,N_10966,N_14742);
or U15687 (N_15687,N_11585,N_13365);
and U15688 (N_15688,N_13879,N_14967);
or U15689 (N_15689,N_14860,N_13476);
nor U15690 (N_15690,N_11794,N_10104);
nor U15691 (N_15691,N_11413,N_12019);
nand U15692 (N_15692,N_12192,N_10349);
or U15693 (N_15693,N_12403,N_11732);
and U15694 (N_15694,N_13693,N_14725);
nand U15695 (N_15695,N_12258,N_11356);
nor U15696 (N_15696,N_12149,N_12739);
nor U15697 (N_15697,N_11290,N_11944);
nor U15698 (N_15698,N_13614,N_14010);
or U15699 (N_15699,N_14303,N_10312);
nand U15700 (N_15700,N_14977,N_10258);
or U15701 (N_15701,N_14098,N_10062);
nor U15702 (N_15702,N_10893,N_12989);
nor U15703 (N_15703,N_10271,N_13401);
and U15704 (N_15704,N_12678,N_11237);
or U15705 (N_15705,N_14809,N_12367);
or U15706 (N_15706,N_13368,N_10564);
nor U15707 (N_15707,N_13578,N_10323);
or U15708 (N_15708,N_12809,N_14200);
nand U15709 (N_15709,N_13726,N_11600);
and U15710 (N_15710,N_14055,N_14468);
nor U15711 (N_15711,N_13105,N_11630);
nand U15712 (N_15712,N_10406,N_14330);
or U15713 (N_15713,N_13714,N_14758);
or U15714 (N_15714,N_11390,N_14628);
nand U15715 (N_15715,N_11594,N_10514);
nand U15716 (N_15716,N_13754,N_14399);
nand U15717 (N_15717,N_12734,N_12275);
or U15718 (N_15718,N_14407,N_11122);
or U15719 (N_15719,N_12569,N_12781);
and U15720 (N_15720,N_11787,N_10254);
or U15721 (N_15721,N_14755,N_14553);
and U15722 (N_15722,N_14415,N_11225);
nand U15723 (N_15723,N_10334,N_10468);
or U15724 (N_15724,N_11846,N_10909);
nor U15725 (N_15725,N_11391,N_12330);
nand U15726 (N_15726,N_14067,N_13755);
or U15727 (N_15727,N_12077,N_14749);
nand U15728 (N_15728,N_14622,N_14983);
and U15729 (N_15729,N_11714,N_14278);
and U15730 (N_15730,N_13651,N_12178);
and U15731 (N_15731,N_10916,N_10895);
xor U15732 (N_15732,N_10960,N_13532);
nand U15733 (N_15733,N_10825,N_12306);
and U15734 (N_15734,N_11564,N_14060);
and U15735 (N_15735,N_14029,N_12321);
nand U15736 (N_15736,N_10151,N_14544);
or U15737 (N_15737,N_12613,N_13321);
or U15738 (N_15738,N_14886,N_10436);
nor U15739 (N_15739,N_12609,N_11031);
nand U15740 (N_15740,N_10045,N_14658);
nand U15741 (N_15741,N_10981,N_13481);
or U15742 (N_15742,N_13482,N_14389);
and U15743 (N_15743,N_11922,N_13435);
nor U15744 (N_15744,N_10595,N_13023);
nand U15745 (N_15745,N_12859,N_11612);
or U15746 (N_15746,N_12522,N_10633);
and U15747 (N_15747,N_10413,N_14289);
nor U15748 (N_15748,N_14584,N_10988);
nor U15749 (N_15749,N_10315,N_11511);
and U15750 (N_15750,N_14409,N_14734);
nor U15751 (N_15751,N_14269,N_12193);
and U15752 (N_15752,N_14537,N_10234);
or U15753 (N_15753,N_12116,N_10381);
nand U15754 (N_15754,N_10040,N_13315);
and U15755 (N_15755,N_10000,N_12271);
xor U15756 (N_15756,N_12663,N_12011);
nor U15757 (N_15757,N_10713,N_12176);
nor U15758 (N_15758,N_10827,N_14411);
or U15759 (N_15759,N_10304,N_14297);
or U15760 (N_15760,N_11556,N_12882);
nand U15761 (N_15761,N_10584,N_11177);
nor U15762 (N_15762,N_12300,N_13779);
nand U15763 (N_15763,N_10106,N_10421);
and U15764 (N_15764,N_13188,N_10046);
or U15765 (N_15765,N_11253,N_13682);
and U15766 (N_15766,N_11249,N_12190);
or U15767 (N_15767,N_13659,N_14366);
or U15768 (N_15768,N_14150,N_10451);
nor U15769 (N_15769,N_10649,N_12550);
or U15770 (N_15770,N_10955,N_11366);
nand U15771 (N_15771,N_11831,N_14733);
nand U15772 (N_15772,N_10828,N_14364);
nor U15773 (N_15773,N_12590,N_10503);
nand U15774 (N_15774,N_14391,N_12681);
or U15775 (N_15775,N_14946,N_10896);
nand U15776 (N_15776,N_13136,N_12938);
or U15777 (N_15777,N_10286,N_13957);
and U15778 (N_15778,N_11247,N_10709);
or U15779 (N_15779,N_13017,N_10267);
nand U15780 (N_15780,N_12264,N_11951);
and U15781 (N_15781,N_12236,N_10944);
xor U15782 (N_15782,N_13267,N_11213);
xnor U15783 (N_15783,N_14859,N_12533);
xnor U15784 (N_15784,N_13512,N_14684);
nand U15785 (N_15785,N_13687,N_11215);
nand U15786 (N_15786,N_13831,N_14817);
nand U15787 (N_15787,N_14931,N_14145);
nor U15788 (N_15788,N_12400,N_12453);
and U15789 (N_15789,N_11952,N_14996);
and U15790 (N_15790,N_13104,N_14822);
nand U15791 (N_15791,N_13579,N_14469);
and U15792 (N_15792,N_14140,N_10941);
and U15793 (N_15793,N_14835,N_12098);
xnor U15794 (N_15794,N_14111,N_10094);
xnor U15795 (N_15795,N_10390,N_10102);
or U15796 (N_15796,N_14020,N_12050);
nand U15797 (N_15797,N_13094,N_12991);
or U15798 (N_15798,N_13337,N_14350);
xor U15799 (N_15799,N_14158,N_13589);
nand U15800 (N_15800,N_12351,N_13183);
and U15801 (N_15801,N_14046,N_12390);
and U15802 (N_15802,N_13067,N_10467);
nand U15803 (N_15803,N_10266,N_12923);
or U15804 (N_15804,N_12641,N_14322);
nor U15805 (N_15805,N_11397,N_10432);
and U15806 (N_15806,N_14360,N_13849);
xnor U15807 (N_15807,N_11886,N_12230);
nor U15808 (N_15808,N_11012,N_10771);
and U15809 (N_15809,N_10590,N_11148);
nand U15810 (N_15810,N_11708,N_12257);
nor U15811 (N_15811,N_12104,N_12479);
nor U15812 (N_15812,N_12863,N_14921);
or U15813 (N_15813,N_10543,N_10038);
or U15814 (N_15814,N_11673,N_14605);
or U15815 (N_15815,N_10202,N_11751);
nand U15816 (N_15816,N_12097,N_14051);
nor U15817 (N_15817,N_10296,N_13046);
nand U15818 (N_15818,N_10148,N_13031);
xnor U15819 (N_15819,N_11916,N_12946);
nand U15820 (N_15820,N_12375,N_10481);
nand U15821 (N_15821,N_11979,N_13533);
and U15822 (N_15822,N_13768,N_10089);
nand U15823 (N_15823,N_12621,N_12151);
nor U15824 (N_15824,N_11178,N_12379);
and U15825 (N_15825,N_11551,N_14963);
or U15826 (N_15826,N_10095,N_10659);
and U15827 (N_15827,N_12297,N_13824);
xnor U15828 (N_15828,N_12398,N_14998);
or U15829 (N_15829,N_10986,N_11581);
or U15830 (N_15830,N_10319,N_10579);
and U15831 (N_15831,N_14666,N_10116);
nor U15832 (N_15832,N_14084,N_14891);
and U15833 (N_15833,N_11211,N_13096);
nand U15834 (N_15834,N_12466,N_12594);
nor U15835 (N_15835,N_10324,N_12032);
xor U15836 (N_15836,N_10671,N_12373);
and U15837 (N_15837,N_11374,N_12285);
nor U15838 (N_15838,N_10745,N_13960);
nand U15839 (N_15839,N_14334,N_13487);
or U15840 (N_15840,N_14710,N_12858);
xnor U15841 (N_15841,N_12435,N_11523);
nor U15842 (N_15842,N_13281,N_14600);
xor U15843 (N_15843,N_13239,N_12670);
xnor U15844 (N_15844,N_12857,N_10496);
nand U15845 (N_15845,N_12819,N_12225);
nor U15846 (N_15846,N_12224,N_12726);
nor U15847 (N_15847,N_11962,N_14260);
and U15848 (N_15848,N_11469,N_10740);
or U15849 (N_15849,N_13192,N_13361);
or U15850 (N_15850,N_14284,N_11955);
nand U15851 (N_15851,N_13250,N_10812);
and U15852 (N_15852,N_11765,N_14827);
or U15853 (N_15853,N_12807,N_14542);
nor U15854 (N_15854,N_13677,N_11302);
or U15855 (N_15855,N_11605,N_12815);
and U15856 (N_15856,N_11566,N_12489);
xor U15857 (N_15857,N_14760,N_12944);
nand U15858 (N_15858,N_14593,N_12267);
nor U15859 (N_15859,N_12334,N_10870);
nand U15860 (N_15860,N_10305,N_10352);
nor U15861 (N_15861,N_13211,N_13295);
nor U15862 (N_15862,N_13936,N_11412);
or U15863 (N_15863,N_14776,N_13611);
and U15864 (N_15864,N_13986,N_14631);
or U15865 (N_15865,N_10015,N_10242);
xor U15866 (N_15866,N_13834,N_11100);
and U15867 (N_15867,N_13247,N_11233);
or U15868 (N_15868,N_10220,N_12422);
nand U15869 (N_15869,N_11721,N_14968);
nand U15870 (N_15870,N_10387,N_12326);
nor U15871 (N_15871,N_13446,N_14850);
and U15872 (N_15872,N_13864,N_12928);
and U15873 (N_15873,N_12535,N_13039);
nor U15874 (N_15874,N_10699,N_14747);
nand U15875 (N_15875,N_14134,N_10873);
nand U15876 (N_15876,N_14347,N_12743);
and U15877 (N_15877,N_12327,N_13101);
nor U15878 (N_15878,N_12028,N_13632);
or U15879 (N_15879,N_10722,N_12841);
nand U15880 (N_15880,N_11814,N_14688);
xor U15881 (N_15881,N_13496,N_10154);
nor U15882 (N_15882,N_12091,N_14114);
nor U15883 (N_15883,N_10741,N_11923);
and U15884 (N_15884,N_10008,N_10905);
nand U15885 (N_15885,N_12459,N_13788);
nand U15886 (N_15886,N_10328,N_10580);
and U15887 (N_15887,N_13951,N_10108);
and U15888 (N_15888,N_14696,N_10838);
and U15889 (N_15889,N_10606,N_12607);
nor U15890 (N_15890,N_10569,N_12564);
nor U15891 (N_15891,N_13624,N_14405);
and U15892 (N_15892,N_12221,N_13320);
or U15893 (N_15893,N_11318,N_10011);
xnor U15894 (N_15894,N_11128,N_10019);
or U15895 (N_15895,N_11785,N_10411);
or U15896 (N_15896,N_14496,N_13607);
and U15897 (N_15897,N_10039,N_13210);
nor U15898 (N_15898,N_13549,N_10755);
nand U15899 (N_15899,N_14240,N_12999);
nor U15900 (N_15900,N_13910,N_12317);
nand U15901 (N_15901,N_12312,N_13730);
xor U15902 (N_15902,N_13150,N_14348);
nor U15903 (N_15903,N_13812,N_13912);
nand U15904 (N_15904,N_11885,N_10167);
or U15905 (N_15905,N_11678,N_14316);
nor U15906 (N_15906,N_14941,N_13795);
xnor U15907 (N_15907,N_12961,N_10545);
nand U15908 (N_15908,N_13474,N_12138);
and U15909 (N_15909,N_11364,N_13852);
and U15910 (N_15910,N_12249,N_14455);
and U15911 (N_15911,N_12719,N_13413);
nor U15912 (N_15912,N_11877,N_10353);
and U15913 (N_15913,N_12514,N_11633);
nand U15914 (N_15914,N_14088,N_14148);
xnor U15915 (N_15915,N_11488,N_11358);
xnor U15916 (N_15916,N_13818,N_14727);
nor U15917 (N_15917,N_14557,N_14564);
or U15918 (N_15918,N_13407,N_12214);
or U15919 (N_15919,N_12325,N_11819);
and U15920 (N_15920,N_12437,N_12402);
xnor U15921 (N_15921,N_12599,N_12242);
xor U15922 (N_15922,N_14608,N_10758);
nor U15923 (N_15923,N_11899,N_12766);
and U15924 (N_15924,N_10574,N_11450);
or U15925 (N_15925,N_12356,N_10513);
or U15926 (N_15926,N_10003,N_11907);
nand U15927 (N_15927,N_10900,N_12552);
or U15928 (N_15928,N_14730,N_12828);
or U15929 (N_15929,N_11685,N_10952);
and U15930 (N_15930,N_14743,N_10796);
nor U15931 (N_15931,N_11582,N_11056);
nor U15932 (N_15932,N_11775,N_10191);
and U15933 (N_15933,N_10392,N_11067);
nor U15934 (N_15934,N_10831,N_13300);
xor U15935 (N_15935,N_12388,N_13298);
and U15936 (N_15936,N_13043,N_12282);
nand U15937 (N_15937,N_10098,N_11371);
xor U15938 (N_15938,N_12608,N_10184);
nor U15939 (N_15939,N_10897,N_14369);
nand U15940 (N_15940,N_12823,N_13422);
nor U15941 (N_15941,N_14290,N_13877);
nand U15942 (N_15942,N_10087,N_12345);
or U15943 (N_15943,N_13450,N_14487);
or U15944 (N_15944,N_13229,N_10394);
nor U15945 (N_15945,N_11327,N_11540);
or U15946 (N_15946,N_12777,N_11005);
or U15947 (N_15947,N_10357,N_10677);
nand U15948 (N_15948,N_14128,N_12886);
nand U15949 (N_15949,N_12126,N_10358);
or U15950 (N_15950,N_14266,N_10558);
nor U15951 (N_15951,N_11825,N_12759);
xor U15952 (N_15952,N_10330,N_13460);
nand U15953 (N_15953,N_14197,N_10193);
and U15954 (N_15954,N_12086,N_12065);
or U15955 (N_15955,N_13732,N_12760);
nor U15956 (N_15956,N_10114,N_12906);
and U15957 (N_15957,N_10970,N_14250);
or U15958 (N_15958,N_13508,N_13329);
or U15959 (N_15959,N_12512,N_14143);
xnor U15960 (N_15960,N_14952,N_14133);
nand U15961 (N_15961,N_13926,N_14156);
or U15962 (N_15962,N_11228,N_12547);
nand U15963 (N_15963,N_10541,N_13740);
xor U15964 (N_15964,N_14380,N_13327);
xor U15965 (N_15965,N_13182,N_13175);
and U15966 (N_15966,N_10404,N_11227);
nand U15967 (N_15967,N_11437,N_13899);
xnor U15968 (N_15968,N_13246,N_10790);
and U15969 (N_15969,N_10321,N_11388);
xor U15970 (N_15970,N_14398,N_14234);
or U15971 (N_15971,N_10054,N_13322);
and U15972 (N_15972,N_11278,N_12115);
and U15973 (N_15973,N_12786,N_11027);
and U15974 (N_15974,N_13118,N_11376);
nand U15975 (N_15975,N_14939,N_14122);
nand U15976 (N_15976,N_10977,N_11615);
nor U15977 (N_15977,N_14554,N_14997);
xnor U15978 (N_15978,N_14085,N_13582);
or U15979 (N_15979,N_12215,N_12089);
nand U15980 (N_15980,N_11908,N_10566);
nor U15981 (N_15981,N_11500,N_14779);
nand U15982 (N_15982,N_12283,N_13001);
or U15983 (N_15983,N_14356,N_12894);
or U15984 (N_15984,N_13459,N_14774);
nand U15985 (N_15985,N_10693,N_11339);
xor U15986 (N_15986,N_11342,N_12066);
nor U15987 (N_15987,N_11114,N_14130);
xor U15988 (N_15988,N_13019,N_10776);
or U15989 (N_15989,N_10475,N_10224);
and U15990 (N_15990,N_13443,N_14066);
or U15991 (N_15991,N_12561,N_13006);
xor U15992 (N_15992,N_10625,N_13785);
or U15993 (N_15993,N_14672,N_13264);
nor U15994 (N_15994,N_13331,N_10469);
and U15995 (N_15995,N_10465,N_14604);
and U15996 (N_15996,N_11507,N_13154);
nor U15997 (N_15997,N_10065,N_12747);
nand U15998 (N_15998,N_10942,N_12521);
and U15999 (N_15999,N_14908,N_12528);
xor U16000 (N_16000,N_13857,N_10074);
nand U16001 (N_16001,N_12174,N_10554);
nand U16002 (N_16002,N_11332,N_14717);
nand U16003 (N_16003,N_13674,N_14999);
xor U16004 (N_16004,N_13762,N_12674);
nor U16005 (N_16005,N_12222,N_10613);
or U16006 (N_16006,N_10871,N_11061);
xor U16007 (N_16007,N_13130,N_11073);
nand U16008 (N_16008,N_10142,N_13584);
nand U16009 (N_16009,N_11222,N_12643);
and U16010 (N_16010,N_10804,N_13544);
or U16011 (N_16011,N_11953,N_10506);
xor U16012 (N_16012,N_13681,N_10386);
and U16013 (N_16013,N_11786,N_12788);
or U16014 (N_16014,N_13964,N_12789);
and U16015 (N_16015,N_13511,N_10853);
and U16016 (N_16016,N_10879,N_14204);
and U16017 (N_16017,N_11593,N_14376);
xnor U16018 (N_16018,N_11870,N_11859);
and U16019 (N_16019,N_12866,N_12099);
or U16020 (N_16020,N_13952,N_11830);
and U16021 (N_16021,N_14257,N_14769);
and U16022 (N_16022,N_11874,N_11531);
nor U16023 (N_16023,N_13196,N_11757);
xor U16024 (N_16024,N_13354,N_14903);
and U16025 (N_16025,N_11189,N_13949);
nand U16026 (N_16026,N_14500,N_13052);
and U16027 (N_16027,N_10585,N_11574);
nand U16028 (N_16028,N_10770,N_13086);
or U16029 (N_16029,N_13801,N_13775);
xnor U16030 (N_16030,N_13077,N_14351);
xnor U16031 (N_16031,N_14517,N_11471);
nand U16032 (N_16032,N_11755,N_13827);
nor U16033 (N_16033,N_14510,N_11435);
nand U16034 (N_16034,N_10259,N_14323);
and U16035 (N_16035,N_13545,N_13823);
xor U16036 (N_16036,N_14152,N_14949);
and U16037 (N_16037,N_10931,N_14346);
nor U16038 (N_16038,N_11078,N_14169);
nand U16039 (N_16039,N_12892,N_11749);
nand U16040 (N_16040,N_11350,N_13254);
nand U16041 (N_16041,N_12187,N_10516);
and U16042 (N_16042,N_12454,N_10396);
or U16043 (N_16043,N_14962,N_14585);
nand U16044 (N_16044,N_14480,N_11242);
or U16045 (N_16045,N_11608,N_14854);
or U16046 (N_16046,N_13618,N_12628);
and U16047 (N_16047,N_14697,N_11947);
or U16048 (N_16048,N_13380,N_13362);
nand U16049 (N_16049,N_12101,N_11295);
nor U16050 (N_16050,N_10056,N_12270);
nand U16051 (N_16051,N_11429,N_14913);
and U16052 (N_16052,N_13179,N_12713);
nor U16053 (N_16053,N_13712,N_11466);
nor U16054 (N_16054,N_14461,N_12653);
nand U16055 (N_16055,N_13048,N_11798);
nand U16056 (N_16056,N_13276,N_11648);
and U16057 (N_16057,N_11616,N_14701);
nor U16058 (N_16058,N_14325,N_10366);
or U16059 (N_16059,N_14254,N_12113);
or U16060 (N_16060,N_13708,N_10401);
and U16061 (N_16061,N_11268,N_14214);
nand U16062 (N_16062,N_12408,N_10303);
xnor U16063 (N_16063,N_10241,N_11461);
or U16064 (N_16064,N_10072,N_10723);
nand U16065 (N_16065,N_14650,N_12767);
or U16066 (N_16066,N_12856,N_14328);
or U16067 (N_16067,N_14095,N_10805);
xnor U16068 (N_16068,N_14764,N_12419);
and U16069 (N_16069,N_10143,N_11203);
and U16070 (N_16070,N_12936,N_13753);
and U16071 (N_16071,N_13931,N_11533);
and U16072 (N_16072,N_13050,N_12448);
or U16073 (N_16073,N_13439,N_11045);
xnor U16074 (N_16074,N_11706,N_14074);
and U16075 (N_16075,N_13679,N_14852);
or U16076 (N_16076,N_10257,N_14478);
nor U16077 (N_16077,N_14582,N_10617);
and U16078 (N_16078,N_11904,N_12591);
and U16079 (N_16079,N_10063,N_11212);
and U16080 (N_16080,N_13627,N_14699);
and U16081 (N_16081,N_10899,N_11448);
nand U16082 (N_16082,N_13235,N_12526);
or U16083 (N_16083,N_12704,N_13160);
or U16084 (N_16084,N_13203,N_11964);
nor U16085 (N_16085,N_14218,N_10891);
or U16086 (N_16086,N_12947,N_13505);
nand U16087 (N_16087,N_10055,N_14079);
or U16088 (N_16088,N_12362,N_12725);
or U16089 (N_16089,N_12316,N_11096);
and U16090 (N_16090,N_14575,N_14426);
nor U16091 (N_16091,N_14993,N_10650);
or U16092 (N_16092,N_13769,N_11657);
nor U16093 (N_16093,N_12816,N_11720);
nor U16094 (N_16094,N_12572,N_10203);
or U16095 (N_16095,N_11217,N_11016);
nand U16096 (N_16096,N_11526,N_14954);
nand U16097 (N_16097,N_12637,N_10631);
and U16098 (N_16098,N_10085,N_13114);
and U16099 (N_16099,N_14675,N_14531);
nand U16100 (N_16100,N_12861,N_12646);
and U16101 (N_16101,N_13675,N_11520);
and U16102 (N_16102,N_10020,N_11659);
nor U16103 (N_16103,N_12897,N_14548);
and U16104 (N_16104,N_12933,N_12432);
and U16105 (N_16105,N_10122,N_12905);
or U16106 (N_16106,N_11766,N_14870);
nor U16107 (N_16107,N_12474,N_14748);
nand U16108 (N_16108,N_12967,N_10053);
xnor U16109 (N_16109,N_10537,N_11509);
or U16110 (N_16110,N_12001,N_10201);
and U16111 (N_16111,N_14049,N_12191);
or U16112 (N_16112,N_10182,N_13820);
and U16113 (N_16113,N_10359,N_11062);
nor U16114 (N_16114,N_11754,N_14825);
or U16115 (N_16115,N_12007,N_10858);
xor U16116 (N_16116,N_13355,N_11906);
nor U16117 (N_16117,N_10351,N_10079);
or U16118 (N_16118,N_10533,N_14950);
nor U16119 (N_16119,N_13342,N_10576);
nor U16120 (N_16120,N_13133,N_10518);
or U16121 (N_16121,N_12829,N_14183);
nand U16122 (N_16122,N_13814,N_14685);
nor U16123 (N_16123,N_12467,N_11421);
nor U16124 (N_16124,N_10876,N_13310);
xnor U16125 (N_16125,N_14595,N_13489);
and U16126 (N_16126,N_13491,N_10575);
or U16127 (N_16127,N_11769,N_10532);
nor U16128 (N_16128,N_12744,N_12733);
or U16129 (N_16129,N_12004,N_11617);
and U16130 (N_16130,N_14957,N_13971);
nand U16131 (N_16131,N_10002,N_14670);
nand U16132 (N_16132,N_12868,N_11905);
nand U16133 (N_16133,N_10803,N_11868);
and U16134 (N_16134,N_10288,N_12446);
or U16135 (N_16135,N_14906,N_12048);
or U16136 (N_16136,N_12710,N_14392);
xnor U16137 (N_16137,N_14115,N_10808);
nand U16138 (N_16138,N_13780,N_13956);
nand U16139 (N_16139,N_12901,N_13873);
or U16140 (N_16140,N_14829,N_13445);
nand U16141 (N_16141,N_12735,N_13111);
xor U16142 (N_16142,N_13595,N_10416);
and U16143 (N_16143,N_12630,N_13718);
or U16144 (N_16144,N_11197,N_10626);
nor U16145 (N_16145,N_14856,N_13008);
nor U16146 (N_16146,N_13110,N_13187);
nor U16147 (N_16147,N_10031,N_13970);
nor U16148 (N_16148,N_11403,N_10560);
nor U16149 (N_16149,N_14280,N_14509);
or U16150 (N_16150,N_10078,N_13984);
nor U16151 (N_16151,N_10218,N_11822);
nand U16152 (N_16152,N_11866,N_11845);
nand U16153 (N_16153,N_14807,N_12420);
nor U16154 (N_16154,N_13859,N_14381);
nor U16155 (N_16155,N_12650,N_14634);
nand U16156 (N_16156,N_14249,N_10384);
nor U16157 (N_16157,N_13408,N_10415);
xor U16158 (N_16158,N_11499,N_13026);
nand U16159 (N_16159,N_10837,N_10605);
nor U16160 (N_16160,N_13686,N_10057);
nor U16161 (N_16161,N_13600,N_13099);
nor U16162 (N_16162,N_13610,N_14802);
nor U16163 (N_16163,N_12568,N_14866);
and U16164 (N_16164,N_12814,N_11774);
nand U16165 (N_16165,N_14105,N_10971);
nand U16166 (N_16166,N_11839,N_11674);
nand U16167 (N_16167,N_10854,N_13279);
or U16168 (N_16168,N_11601,N_11010);
nor U16169 (N_16169,N_11767,N_10498);
nand U16170 (N_16170,N_10101,N_10177);
nor U16171 (N_16171,N_10742,N_11123);
nand U16172 (N_16172,N_14873,N_11959);
nor U16173 (N_16173,N_10338,N_10133);
and U16174 (N_16174,N_12014,N_13619);
xor U16175 (N_16175,N_10775,N_14598);
nand U16176 (N_16176,N_10314,N_12778);
nand U16177 (N_16177,N_12292,N_11396);
and U16178 (N_16178,N_14454,N_11970);
nand U16179 (N_16179,N_12159,N_11367);
nor U16180 (N_16180,N_14724,N_13041);
nor U16181 (N_16181,N_13546,N_10252);
xor U16182 (N_16182,N_10214,N_13942);
nand U16183 (N_16183,N_13773,N_13161);
xnor U16184 (N_16184,N_12656,N_12339);
or U16185 (N_16185,N_14901,N_14099);
nand U16186 (N_16186,N_12855,N_11453);
and U16187 (N_16187,N_14559,N_10824);
and U16188 (N_16188,N_12094,N_11360);
nor U16189 (N_16189,N_11296,N_10604);
or U16190 (N_16190,N_11883,N_13004);
or U16191 (N_16191,N_14090,N_10024);
nor U16192 (N_16192,N_13384,N_10855);
nand U16193 (N_16193,N_13848,N_10013);
and U16194 (N_16194,N_10784,N_13807);
and U16195 (N_16195,N_10327,N_10525);
nor U16196 (N_16196,N_13999,N_12301);
or U16197 (N_16197,N_12440,N_12930);
and U16198 (N_16198,N_12371,N_10975);
xnor U16199 (N_16199,N_11434,N_14770);
or U16200 (N_16200,N_11515,N_11098);
xnor U16201 (N_16201,N_12357,N_13903);
or U16202 (N_16202,N_13389,N_11707);
or U16203 (N_16203,N_13603,N_13409);
xnor U16204 (N_16204,N_13402,N_11806);
and U16205 (N_16205,N_14263,N_14656);
xnor U16206 (N_16206,N_12922,N_10422);
or U16207 (N_16207,N_14744,N_11252);
xor U16208 (N_16208,N_13783,N_10120);
or U16209 (N_16209,N_14458,N_14535);
or U16210 (N_16210,N_12870,N_14100);
or U16211 (N_16211,N_13143,N_12218);
and U16212 (N_16212,N_14058,N_10230);
or U16213 (N_16213,N_14893,N_11572);
or U16214 (N_16214,N_12415,N_11195);
xor U16215 (N_16215,N_13212,N_12889);
nor U16216 (N_16216,N_14048,N_14491);
and U16217 (N_16217,N_14080,N_11194);
nor U16218 (N_16218,N_11365,N_10681);
nor U16219 (N_16219,N_13592,N_11949);
nand U16220 (N_16220,N_10280,N_11109);
nor U16221 (N_16221,N_12634,N_10208);
nor U16222 (N_16222,N_14421,N_12520);
nor U16223 (N_16223,N_11014,N_14698);
or U16224 (N_16224,N_14806,N_12168);
xnor U16225 (N_16225,N_14508,N_14007);
or U16226 (N_16226,N_12473,N_14429);
or U16227 (N_16227,N_14035,N_13638);
nor U16228 (N_16228,N_13615,N_12900);
nand U16229 (N_16229,N_12813,N_14925);
nand U16230 (N_16230,N_10974,N_12993);
nor U16231 (N_16231,N_12977,N_14576);
nor U16232 (N_16232,N_14307,N_10495);
nand U16233 (N_16233,N_12265,N_11780);
nand U16234 (N_16234,N_13438,N_13158);
and U16235 (N_16235,N_13666,N_11570);
nand U16236 (N_16236,N_14062,N_11932);
or U16237 (N_16237,N_14004,N_14437);
nor U16238 (N_16238,N_14507,N_14333);
and U16239 (N_16239,N_10082,N_10781);
and U16240 (N_16240,N_11957,N_10682);
nor U16241 (N_16241,N_14026,N_13629);
and U16242 (N_16242,N_12832,N_13982);
or U16243 (N_16243,N_11913,N_11683);
nand U16244 (N_16244,N_14910,N_11164);
or U16245 (N_16245,N_11958,N_11411);
or U16246 (N_16246,N_12200,N_12844);
or U16247 (N_16247,N_11276,N_13850);
or U16248 (N_16248,N_11210,N_10751);
or U16249 (N_16249,N_10490,N_10430);
or U16250 (N_16250,N_13037,N_13946);
nand U16251 (N_16251,N_10211,N_11323);
nor U16252 (N_16252,N_10801,N_11155);
nor U16253 (N_16253,N_13894,N_14547);
and U16254 (N_16254,N_12405,N_14832);
or U16255 (N_16255,N_10379,N_14027);
nand U16256 (N_16256,N_10361,N_12549);
or U16257 (N_16257,N_13285,N_11524);
nand U16258 (N_16258,N_11590,N_14446);
nor U16259 (N_16259,N_10150,N_13420);
nor U16260 (N_16260,N_11102,N_11686);
nor U16261 (N_16261,N_12737,N_11053);
nand U16262 (N_16262,N_13441,N_11129);
nor U16263 (N_16263,N_13370,N_11463);
and U16264 (N_16264,N_10583,N_11881);
and U16265 (N_16265,N_11580,N_13393);
nor U16266 (N_16266,N_13063,N_10935);
and U16267 (N_16267,N_11291,N_13889);
or U16268 (N_16268,N_11703,N_11036);
xor U16269 (N_16269,N_10823,N_11569);
nand U16270 (N_16270,N_10548,N_11571);
or U16271 (N_16271,N_11854,N_10839);
nor U16272 (N_16272,N_12201,N_12720);
or U16273 (N_16273,N_11347,N_11090);
xnor U16274 (N_16274,N_13516,N_13479);
nand U16275 (N_16275,N_10703,N_12606);
nand U16276 (N_16276,N_13972,N_14536);
nor U16277 (N_16277,N_12043,N_11020);
or U16278 (N_16278,N_14645,N_12287);
nand U16279 (N_16279,N_14024,N_10921);
and U16280 (N_16280,N_10308,N_11741);
and U16281 (N_16281,N_11934,N_10424);
or U16282 (N_16282,N_12052,N_12499);
nor U16283 (N_16283,N_13628,N_14276);
nor U16284 (N_16284,N_10782,N_11441);
or U16285 (N_16285,N_13070,N_11370);
and U16286 (N_16286,N_11476,N_10449);
nor U16287 (N_16287,N_12320,N_12059);
nand U16288 (N_16288,N_14785,N_14711);
or U16289 (N_16289,N_10992,N_14447);
nor U16290 (N_16290,N_11548,N_12723);
nand U16291 (N_16291,N_13985,N_11638);
nor U16292 (N_16292,N_12240,N_11596);
and U16293 (N_16293,N_10645,N_11809);
and U16294 (N_16294,N_13204,N_12386);
nand U16295 (N_16295,N_11518,N_14042);
or U16296 (N_16296,N_14401,N_13863);
xnor U16297 (N_16297,N_14003,N_12315);
xor U16298 (N_16298,N_13375,N_12504);
nand U16299 (N_16299,N_13577,N_13855);
nor U16300 (N_16300,N_10757,N_13294);
and U16301 (N_16301,N_10793,N_13238);
or U16302 (N_16302,N_10872,N_13390);
nor U16303 (N_16303,N_13049,N_13925);
nand U16304 (N_16304,N_14056,N_10139);
nand U16305 (N_16305,N_10984,N_14414);
xnor U16306 (N_16306,N_12696,N_11439);
nand U16307 (N_16307,N_14435,N_11661);
or U16308 (N_16308,N_13290,N_12329);
nor U16309 (N_16309,N_11143,N_10322);
or U16310 (N_16310,N_11856,N_14096);
or U16311 (N_16311,N_13560,N_12987);
nor U16312 (N_16312,N_14224,N_10967);
nand U16313 (N_16313,N_14824,N_10732);
and U16314 (N_16314,N_14341,N_10608);
nand U16315 (N_16315,N_12677,N_10192);
or U16316 (N_16316,N_10842,N_12711);
nor U16317 (N_16317,N_12160,N_12434);
or U16318 (N_16318,N_14621,N_12417);
or U16319 (N_16319,N_11289,N_11079);
and U16320 (N_16320,N_13606,N_11230);
or U16321 (N_16321,N_14078,N_10043);
xor U16322 (N_16322,N_11631,N_13056);
or U16323 (N_16323,N_13195,N_14933);
nand U16324 (N_16324,N_12651,N_14283);
and U16325 (N_16325,N_13232,N_12295);
nor U16326 (N_16326,N_12978,N_13153);
nand U16327 (N_16327,N_12049,N_11554);
or U16328 (N_16328,N_12697,N_12574);
xor U16329 (N_16329,N_10704,N_14168);
nor U16330 (N_16330,N_10950,N_14686);
or U16331 (N_16331,N_14657,N_10920);
nor U16332 (N_16332,N_10718,N_11311);
and U16333 (N_16333,N_10152,N_11229);
or U16334 (N_16334,N_10993,N_14231);
and U16335 (N_16335,N_14209,N_13434);
and U16336 (N_16336,N_12585,N_10253);
nor U16337 (N_16337,N_10881,N_13278);
and U16338 (N_16338,N_14947,N_11309);
nor U16339 (N_16339,N_12496,N_13721);
or U16340 (N_16340,N_13901,N_12833);
or U16341 (N_16341,N_12860,N_11948);
and U16342 (N_16342,N_10067,N_11788);
or U16343 (N_16343,N_14432,N_11071);
xor U16344 (N_16344,N_14691,N_10696);
and U16345 (N_16345,N_13561,N_11116);
or U16346 (N_16346,N_11599,N_14064);
nand U16347 (N_16347,N_12604,N_14838);
or U16348 (N_16348,N_12348,N_14187);
and U16349 (N_16349,N_12843,N_14370);
nand U16350 (N_16350,N_13379,N_14723);
or U16351 (N_16351,N_12385,N_14803);
nand U16352 (N_16352,N_12366,N_10075);
nand U16353 (N_16353,N_13643,N_13417);
and U16354 (N_16354,N_13213,N_10391);
or U16355 (N_16355,N_10037,N_12955);
nor U16356 (N_16356,N_13412,N_12950);
or U16357 (N_16357,N_14206,N_12918);
nand U16358 (N_16358,N_12180,N_11022);
or U16359 (N_16359,N_13284,N_11864);
and U16360 (N_16360,N_14885,N_14660);
or U16361 (N_16361,N_14937,N_10761);
nor U16362 (N_16362,N_11639,N_12756);
nor U16363 (N_16363,N_10378,N_10447);
nor U16364 (N_16364,N_14332,N_14194);
nor U16365 (N_16365,N_11832,N_10477);
or U16366 (N_16366,N_10816,N_10246);
or U16367 (N_16367,N_10125,N_13804);
nor U16368 (N_16368,N_12438,N_11756);
nor U16369 (N_16369,N_14567,N_11975);
nand U16370 (N_16370,N_10310,N_10957);
nand U16371 (N_16371,N_13363,N_11912);
nand U16372 (N_16372,N_10164,N_13330);
nand U16373 (N_16373,N_10829,N_12288);
and U16374 (N_16374,N_14395,N_11044);
nand U16375 (N_16375,N_14043,N_10016);
nand U16376 (N_16376,N_12635,N_13830);
and U16377 (N_16377,N_12686,N_11054);
or U16378 (N_16378,N_11960,N_11455);
nor U16379 (N_16379,N_10245,N_14144);
nor U16380 (N_16380,N_12309,N_12495);
xnor U16381 (N_16381,N_12394,N_12027);
and U16382 (N_16382,N_12927,N_10500);
nor U16383 (N_16383,N_13360,N_14106);
and U16384 (N_16384,N_11647,N_12262);
nor U16385 (N_16385,N_11941,N_13639);
or U16386 (N_16386,N_11329,N_14188);
nand U16387 (N_16387,N_13312,N_14182);
nor U16388 (N_16388,N_12506,N_10227);
xor U16389 (N_16389,N_14966,N_13225);
nand U16390 (N_16390,N_11898,N_13466);
nor U16391 (N_16391,N_12699,N_13847);
nor U16392 (N_16392,N_14956,N_11712);
or U16393 (N_16393,N_12631,N_10765);
or U16394 (N_16394,N_12970,N_10689);
or U16395 (N_16395,N_14768,N_11758);
and U16396 (N_16396,N_12511,N_10947);
nand U16397 (N_16397,N_14792,N_14988);
nor U16398 (N_16398,N_13633,N_10302);
nand U16399 (N_16399,N_13171,N_11407);
and U16400 (N_16400,N_11984,N_14336);
or U16401 (N_16401,N_14155,N_11368);
or U16402 (N_16402,N_12349,N_11933);
xnor U16403 (N_16403,N_10044,N_14384);
and U16404 (N_16404,N_14879,N_13869);
or U16405 (N_16405,N_14057,N_12203);
nand U16406 (N_16406,N_14462,N_12640);
and U16407 (N_16407,N_13010,N_10614);
and U16408 (N_16408,N_10756,N_14457);
or U16409 (N_16409,N_10843,N_14609);
nand U16410 (N_16410,N_11127,N_13787);
xnor U16411 (N_16411,N_13932,N_11968);
and U16412 (N_16412,N_14107,N_14372);
nor U16413 (N_16413,N_12475,N_14034);
and U16414 (N_16414,N_12013,N_12332);
and U16415 (N_16415,N_10091,N_10367);
nand U16416 (N_16416,N_12998,N_10344);
and U16417 (N_16417,N_14922,N_11498);
and U16418 (N_16418,N_10226,N_13868);
nor U16419 (N_16419,N_10536,N_11763);
nand U16420 (N_16420,N_11651,N_13488);
nor U16421 (N_16421,N_12017,N_10648);
and U16422 (N_16422,N_12205,N_11207);
nor U16423 (N_16423,N_13581,N_10664);
and U16424 (N_16424,N_10886,N_10691);
nand U16425 (N_16425,N_11836,N_12037);
nor U16426 (N_16426,N_11543,N_11834);
xnor U16427 (N_16427,N_11671,N_11303);
and U16428 (N_16428,N_14244,N_11168);
nor U16429 (N_16429,N_12683,N_13941);
and U16430 (N_16430,N_14871,N_14119);
nor U16431 (N_16431,N_12117,N_11850);
nor U16432 (N_16432,N_10932,N_11375);
nor U16433 (N_16433,N_12945,N_12707);
or U16434 (N_16434,N_10291,N_11083);
and U16435 (N_16435,N_12110,N_10029);
nor U16436 (N_16436,N_13758,N_13073);
nand U16437 (N_16437,N_14091,N_12563);
nand U16438 (N_16438,N_13075,N_14219);
nand U16439 (N_16439,N_14959,N_13649);
nor U16440 (N_16440,N_14044,N_13376);
and U16441 (N_16441,N_13042,N_10320);
and U16442 (N_16442,N_12755,N_14786);
and U16443 (N_16443,N_13945,N_12565);
and U16444 (N_16444,N_11181,N_10287);
or U16445 (N_16445,N_13809,N_11487);
or U16446 (N_16446,N_10215,N_12715);
nand U16447 (N_16447,N_14149,N_13571);
or U16448 (N_16448,N_11623,N_12880);
nand U16449 (N_16449,N_14305,N_14304);
nor U16450 (N_16450,N_13794,N_13223);
or U16451 (N_16451,N_10030,N_13790);
and U16452 (N_16452,N_14790,N_13703);
and U16453 (N_16453,N_12620,N_12067);
nand U16454 (N_16454,N_13756,N_11801);
nor U16455 (N_16455,N_13201,N_12769);
nor U16456 (N_16456,N_12913,N_14185);
and U16457 (N_16457,N_10933,N_12951);
or U16458 (N_16458,N_14052,N_13152);
nand U16459 (N_16459,N_14793,N_11940);
nand U16460 (N_16460,N_10729,N_10964);
or U16461 (N_16461,N_14678,N_12693);
and U16462 (N_16462,N_11057,N_10282);
nor U16463 (N_16463,N_10456,N_12155);
or U16464 (N_16464,N_10809,N_11807);
nand U16465 (N_16465,N_14671,N_13523);
nand U16466 (N_16466,N_13108,N_14612);
nor U16467 (N_16467,N_14428,N_14264);
or U16468 (N_16468,N_14796,N_13860);
and U16469 (N_16469,N_11627,N_12626);
nand U16470 (N_16470,N_14842,N_11259);
or U16471 (N_16471,N_10034,N_10275);
or U16472 (N_16472,N_13770,N_13963);
or U16473 (N_16473,N_11017,N_12118);
nand U16474 (N_16474,N_10370,N_10811);
nor U16475 (N_16475,N_14006,N_14136);
and U16476 (N_16476,N_13107,N_14514);
nor U16477 (N_16477,N_13457,N_12812);
xor U16478 (N_16478,N_10728,N_12042);
nand U16479 (N_16479,N_12612,N_12601);
xnor U16480 (N_16480,N_14038,N_14172);
and U16481 (N_16481,N_13165,N_11282);
nand U16482 (N_16482,N_11281,N_11283);
nand U16483 (N_16483,N_10643,N_14157);
xnor U16484 (N_16484,N_10157,N_11994);
or U16485 (N_16485,N_12073,N_12433);
or U16486 (N_16486,N_13631,N_13024);
or U16487 (N_16487,N_13317,N_14810);
nor U16488 (N_16488,N_12202,N_11382);
and U16489 (N_16489,N_12305,N_13514);
and U16490 (N_16490,N_14549,N_12638);
nor U16491 (N_16491,N_14756,N_11838);
or U16492 (N_16492,N_10675,N_12030);
nor U16493 (N_16493,N_12121,N_14418);
or U16494 (N_16494,N_12015,N_11491);
or U16495 (N_16495,N_13387,N_12337);
and U16496 (N_16496,N_13333,N_14248);
nand U16497 (N_16497,N_10963,N_13303);
and U16498 (N_16498,N_14419,N_12867);
nor U16499 (N_16499,N_14940,N_10339);
and U16500 (N_16500,N_11528,N_13590);
nand U16501 (N_16501,N_10769,N_12274);
and U16502 (N_16502,N_14573,N_11119);
xnor U16503 (N_16503,N_14765,N_13475);
and U16504 (N_16504,N_12509,N_12229);
nand U16505 (N_16505,N_13888,N_11936);
nand U16506 (N_16506,N_11454,N_13399);
xnor U16507 (N_16507,N_14973,N_11693);
nor U16508 (N_16508,N_11709,N_11009);
and U16509 (N_16509,N_13626,N_13882);
nand U16510 (N_16510,N_11101,N_14787);
and U16511 (N_16511,N_13262,N_13261);
nor U16512 (N_16512,N_13858,N_12255);
nand U16513 (N_16513,N_13364,N_10973);
and U16514 (N_16514,N_11219,N_10587);
nor U16515 (N_16515,N_13886,N_13258);
nor U16516 (N_16516,N_10747,N_12876);
nor U16517 (N_16517,N_13106,N_12722);
nor U16518 (N_16518,N_13828,N_11652);
nand U16519 (N_16519,N_11875,N_11672);
and U16520 (N_16520,N_14683,N_12063);
xor U16521 (N_16521,N_14761,N_12040);
or U16522 (N_16522,N_14308,N_12256);
and U16523 (N_16523,N_12820,N_14890);
nor U16524 (N_16524,N_13950,N_13711);
nand U16525 (N_16525,N_12445,N_11284);
nand U16526 (N_16526,N_10438,N_14021);
nand U16527 (N_16527,N_14889,N_13013);
nor U16528 (N_16528,N_14513,N_11248);
nor U16529 (N_16529,N_13478,N_13249);
nand U16530 (N_16530,N_11165,N_10382);
and U16531 (N_16531,N_10195,N_12145);
nand U16532 (N_16532,N_11200,N_14131);
nor U16533 (N_16533,N_11173,N_11609);
nand U16534 (N_16534,N_14092,N_10132);
and U16535 (N_16535,N_13381,N_10922);
nor U16536 (N_16536,N_14365,N_13663);
xnor U16537 (N_16537,N_10160,N_13036);
or U16538 (N_16538,N_11159,N_11636);
nor U16539 (N_16539,N_12746,N_11261);
nand U16540 (N_16540,N_11399,N_11742);
and U16541 (N_16541,N_14677,N_12985);
or U16542 (N_16542,N_10913,N_11035);
xnor U16543 (N_16543,N_10721,N_11024);
nand U16544 (N_16544,N_12234,N_13697);
and U16545 (N_16545,N_13745,N_12197);
xor U16546 (N_16546,N_12877,N_12243);
xor U16547 (N_16547,N_14951,N_14390);
nor U16548 (N_16548,N_10437,N_13821);
nand U16549 (N_16549,N_11926,N_11052);
nor U16550 (N_16550,N_13411,N_10565);
nor U16551 (N_16551,N_10799,N_10444);
nand U16552 (N_16552,N_12439,N_12542);
nand U16553 (N_16553,N_14296,N_10221);
nor U16554 (N_16554,N_13396,N_11510);
xor U16555 (N_16555,N_14225,N_11389);
nor U16556 (N_16556,N_12387,N_13458);
or U16557 (N_16557,N_11733,N_10446);
xor U16558 (N_16558,N_12908,N_11626);
nand U16559 (N_16559,N_14923,N_14243);
nand U16560 (N_16560,N_14587,N_12932);
nand U16561 (N_16561,N_14232,N_10307);
nor U16562 (N_16562,N_11634,N_14579);
nor U16563 (N_16563,N_13214,N_14619);
and U16564 (N_16564,N_10483,N_13035);
and U16565 (N_16565,N_14995,N_12142);
nand U16566 (N_16566,N_11992,N_13378);
xor U16567 (N_16567,N_11039,N_12100);
or U16568 (N_16568,N_13743,N_13658);
and U16569 (N_16569,N_10534,N_11810);
xnor U16570 (N_16570,N_11352,N_11710);
xor U16571 (N_16571,N_12431,N_12971);
nand U16572 (N_16572,N_12384,N_10448);
nand U16573 (N_16573,N_12694,N_12893);
and U16574 (N_16574,N_10376,N_14495);
or U16575 (N_16575,N_12780,N_10080);
nand U16576 (N_16576,N_14314,N_11538);
and U16577 (N_16577,N_13706,N_10712);
or U16578 (N_16578,N_12536,N_12299);
nor U16579 (N_16579,N_10130,N_14689);
nand U16580 (N_16580,N_12791,N_12632);
nand U16581 (N_16581,N_12772,N_12033);
or U16582 (N_16582,N_10959,N_12695);
nand U16583 (N_16583,N_12910,N_14800);
and U16584 (N_16584,N_12452,N_10883);
nand U16585 (N_16585,N_11458,N_13887);
and U16586 (N_16586,N_11910,N_10414);
and U16587 (N_16587,N_11722,N_12935);
nor U16588 (N_16588,N_13245,N_11823);
nor U16589 (N_16589,N_12137,N_12328);
nor U16590 (N_16590,N_11613,N_13199);
nand U16591 (N_16591,N_12554,N_12154);
nand U16592 (N_16592,N_12057,N_12354);
or U16593 (N_16593,N_12508,N_13524);
xnor U16594 (N_16594,N_10042,N_13071);
nor U16595 (N_16595,N_12957,N_10646);
nor U16596 (N_16596,N_14293,N_10489);
or U16597 (N_16597,N_14729,N_10635);
nor U16598 (N_16598,N_13403,N_13645);
or U16599 (N_16599,N_11717,N_14718);
nand U16600 (N_16600,N_10701,N_11065);
nand U16601 (N_16601,N_10462,N_12924);
xor U16602 (N_16602,N_12338,N_13093);
nand U16603 (N_16603,N_12839,N_10281);
nand U16604 (N_16604,N_11193,N_12235);
nand U16605 (N_16605,N_10894,N_12556);
nand U16606 (N_16606,N_14920,N_14213);
nand U16607 (N_16607,N_13427,N_13259);
and U16608 (N_16608,N_14093,N_14561);
and U16609 (N_16609,N_10857,N_12241);
or U16610 (N_16610,N_11015,N_10549);
and U16611 (N_16611,N_13287,N_14431);
nand U16612 (N_16612,N_10555,N_12964);
nor U16613 (N_16613,N_13961,N_13720);
nor U16614 (N_16614,N_12548,N_12333);
and U16615 (N_16615,N_10119,N_12463);
or U16616 (N_16616,N_11764,N_13159);
nand U16617 (N_16617,N_13678,N_11750);
nor U16618 (N_16618,N_14329,N_13967);
nor U16619 (N_16619,N_14989,N_13832);
nand U16620 (N_16620,N_13642,N_14097);
and U16621 (N_16621,N_12805,N_10363);
nand U16622 (N_16622,N_14858,N_13089);
or U16623 (N_16623,N_13980,N_13304);
xnor U16624 (N_16624,N_10206,N_11415);
or U16625 (N_16625,N_12682,N_13374);
and U16626 (N_16626,N_11983,N_14358);
nand U16627 (N_16627,N_10052,N_13344);
or U16628 (N_16628,N_11163,N_13027);
nand U16629 (N_16629,N_10336,N_11274);
nor U16630 (N_16630,N_11379,N_12849);
or U16631 (N_16631,N_14083,N_10187);
nand U16632 (N_16632,N_12302,N_13728);
and U16633 (N_16633,N_10768,N_12974);
or U16634 (N_16634,N_13404,N_10428);
or U16635 (N_16635,N_10255,N_11263);
nor U16636 (N_16636,N_12470,N_11095);
nand U16637 (N_16637,N_14565,N_11409);
and U16638 (N_16638,N_11621,N_11154);
or U16639 (N_16639,N_12196,N_11969);
and U16640 (N_16640,N_10118,N_10418);
and U16641 (N_16641,N_12904,N_11465);
and U16642 (N_16642,N_10528,N_13167);
nand U16643 (N_16643,N_14076,N_11892);
xor U16644 (N_16644,N_10229,N_14857);
nand U16645 (N_16645,N_10982,N_10109);
nand U16646 (N_16646,N_11280,N_11300);
nor U16647 (N_16647,N_12840,N_12109);
or U16648 (N_16648,N_10273,N_10313);
or U16649 (N_16649,N_10939,N_10181);
nand U16650 (N_16650,N_13020,N_10178);
or U16651 (N_16651,N_13218,N_11400);
and U16652 (N_16652,N_14572,N_10642);
and U16653 (N_16653,N_13933,N_10640);
and U16654 (N_16654,N_11643,N_10702);
nor U16655 (N_16655,N_12401,N_13307);
nand U16656 (N_16656,N_14721,N_12966);
nor U16657 (N_16657,N_14441,N_13748);
or U16658 (N_16658,N_14865,N_14292);
nor U16659 (N_16659,N_11243,N_13437);
nor U16660 (N_16660,N_12231,N_13248);
and U16661 (N_16661,N_11783,N_10272);
or U16662 (N_16662,N_11597,N_13896);
nor U16663 (N_16663,N_13230,N_13348);
or U16664 (N_16664,N_12486,N_14847);
nand U16665 (N_16665,N_14408,N_10007);
or U16666 (N_16666,N_10517,N_11254);
nor U16667 (N_16667,N_14848,N_14864);
nand U16668 (N_16668,N_13969,N_13622);
nand U16669 (N_16669,N_14017,N_13461);
nand U16670 (N_16670,N_10521,N_12031);
or U16671 (N_16671,N_12578,N_11386);
or U16672 (N_16672,N_14160,N_13586);
and U16673 (N_16673,N_11381,N_13987);
nor U16674 (N_16674,N_14722,N_11884);
xnor U16675 (N_16675,N_13976,N_13916);
nor U16676 (N_16676,N_11561,N_14479);
nor U16677 (N_16677,N_11607,N_14519);
and U16678 (N_16678,N_10083,N_14302);
nand U16679 (N_16679,N_13149,N_13856);
and U16680 (N_16680,N_13994,N_11589);
and U16681 (N_16681,N_12488,N_10644);
nand U16682 (N_16682,N_11251,N_11084);
and U16683 (N_16683,N_10023,N_12413);
and U16684 (N_16684,N_11142,N_11221);
nor U16685 (N_16685,N_13880,N_12558);
xor U16686 (N_16686,N_11738,N_10355);
and U16687 (N_16687,N_10697,N_12233);
nor U16688 (N_16688,N_13018,N_14161);
nor U16689 (N_16689,N_10236,N_11517);
and U16690 (N_16690,N_13947,N_12827);
nand U16691 (N_16691,N_13297,N_14669);
and U16692 (N_16692,N_14146,N_13184);
and U16693 (N_16693,N_13613,N_13433);
xnor U16694 (N_16694,N_10792,N_13742);
nand U16695 (N_16695,N_12237,N_12428);
nand U16696 (N_16696,N_10559,N_12143);
nand U16697 (N_16697,N_12026,N_12615);
nand U16698 (N_16698,N_10141,N_10479);
nor U16699 (N_16699,N_10621,N_13640);
nand U16700 (N_16700,N_13462,N_14976);
and U16701 (N_16701,N_10064,N_11431);
nand U16702 (N_16702,N_13670,N_13705);
or U16703 (N_16703,N_13636,N_11077);
nand U16704 (N_16704,N_11272,N_12926);
nor U16705 (N_16705,N_14482,N_10402);
nor U16706 (N_16706,N_13534,N_10577);
nand U16707 (N_16707,N_12962,N_14352);
or U16708 (N_16708,N_13771,N_11552);
nand U16709 (N_16709,N_11929,N_11271);
or U16710 (N_16710,N_13217,N_12881);
xor U16711 (N_16711,N_12480,N_10017);
or U16712 (N_16712,N_12360,N_10225);
and U16713 (N_16713,N_14417,N_12636);
nor U16714 (N_16714,N_13991,N_14788);
nor U16715 (N_16715,N_12261,N_10505);
and U16716 (N_16716,N_14345,N_13341);
nor U16717 (N_16717,N_12915,N_10856);
and U16718 (N_16718,N_10674,N_13915);
nor U16719 (N_16719,N_11486,N_13729);
or U16720 (N_16720,N_13219,N_14732);
nand U16721 (N_16721,N_10860,N_11485);
nand U16722 (N_16722,N_12830,N_11565);
nor U16723 (N_16723,N_12443,N_11649);
nand U16724 (N_16724,N_14237,N_13266);
or U16725 (N_16725,N_13129,N_13557);
and U16726 (N_16726,N_14463,N_11544);
xnor U16727 (N_16727,N_11089,N_10284);
or U16728 (N_16728,N_11026,N_14533);
and U16729 (N_16729,N_13793,N_10071);
or U16730 (N_16730,N_13034,N_13127);
or U16731 (N_16731,N_13429,N_12652);
nand U16732 (N_16732,N_11895,N_11664);
xnor U16733 (N_16733,N_11299,N_13572);
nor U16734 (N_16734,N_12377,N_13157);
nor U16735 (N_16735,N_12896,N_14767);
xor U16736 (N_16736,N_10069,N_14274);
nor U16737 (N_16737,N_10435,N_12353);
nor U16738 (N_16738,N_11408,N_11909);
or U16739 (N_16739,N_12658,N_10134);
nand U16740 (N_16740,N_14737,N_14578);
nor U16741 (N_16741,N_12979,N_10388);
nor U16742 (N_16742,N_11781,N_14470);
nand U16743 (N_16743,N_10563,N_11214);
and U16744 (N_16744,N_14022,N_12975);
and U16745 (N_16745,N_14310,N_13738);
and U16746 (N_16746,N_11105,N_10115);
xor U16747 (N_16747,N_12074,N_13122);
nor U16748 (N_16748,N_12135,N_10787);
nand U16749 (N_16749,N_11241,N_12268);
and U16750 (N_16750,N_13800,N_13352);
nand U16751 (N_16751,N_12210,N_11789);
xnor U16752 (N_16752,N_10239,N_10869);
nand U16753 (N_16753,N_13492,N_12165);
nor U16754 (N_16754,N_13617,N_10374);
nand U16755 (N_16755,N_13569,N_10551);
nor U16756 (N_16756,N_14102,N_14752);
nor U16757 (N_16757,N_11833,N_11490);
nor U16758 (N_16758,N_12076,N_11816);
nor U16759 (N_16759,N_12478,N_14481);
nand U16760 (N_16760,N_10270,N_13784);
or U16761 (N_16761,N_13977,N_12972);
or U16762 (N_16762,N_11805,N_10600);
or U16763 (N_16763,N_12477,N_13371);
nand U16764 (N_16764,N_12263,N_11475);
and U16765 (N_16765,N_12513,N_12310);
or U16766 (N_16766,N_12427,N_14070);
and U16767 (N_16767,N_13448,N_14324);
and U16768 (N_16768,N_10050,N_14277);
or U16769 (N_16769,N_12627,N_12698);
and U16770 (N_16770,N_12119,N_11346);
xor U16771 (N_16771,N_12021,N_11126);
nand U16772 (N_16772,N_14086,N_13554);
or U16773 (N_16773,N_14037,N_14929);
xnor U16774 (N_16774,N_14980,N_12523);
nor U16775 (N_16775,N_13657,N_13339);
or U16776 (N_16776,N_14178,N_10789);
xnor U16777 (N_16777,N_14211,N_10059);
or U16778 (N_16778,N_14375,N_11943);
nor U16779 (N_16779,N_11513,N_14488);
nand U16780 (N_16780,N_13156,N_11395);
and U16781 (N_16781,N_12560,N_11348);
or U16782 (N_16782,N_11319,N_13798);
xor U16783 (N_16783,N_14955,N_12069);
nor U16784 (N_16784,N_11288,N_13318);
and U16785 (N_16785,N_12156,N_11483);
nand U16786 (N_16786,N_13493,N_14863);
nor U16787 (N_16787,N_10228,N_14286);
and U16788 (N_16788,N_14008,N_14653);
nor U16789 (N_16789,N_10925,N_12541);
nand U16790 (N_16790,N_13351,N_10662);
nor U16791 (N_16791,N_14819,N_14195);
or U16792 (N_16792,N_10711,N_12948);
nor U16793 (N_16793,N_10688,N_11644);
or U16794 (N_16794,N_11602,N_13480);
nor U16795 (N_16795,N_14036,N_14377);
and U16796 (N_16796,N_11901,N_10372);
nor U16797 (N_16797,N_12842,N_14914);
nand U16798 (N_16798,N_10527,N_10399);
nor U16799 (N_16799,N_14970,N_11595);
or U16800 (N_16800,N_11279,N_13350);
and U16801 (N_16801,N_12397,N_14378);
nor U16802 (N_16802,N_13527,N_10331);
nor U16803 (N_16803,N_14777,N_10924);
nor U16804 (N_16804,N_14373,N_13186);
nor U16805 (N_16805,N_11670,N_14900);
nor U16806 (N_16806,N_10036,N_10375);
and U16807 (N_16807,N_14878,N_12212);
xnor U16808 (N_16808,N_10980,N_11646);
nor U16809 (N_16809,N_14849,N_10445);
nor U16810 (N_16810,N_14141,N_11328);
nor U16811 (N_16811,N_11232,N_10417);
nor U16812 (N_16812,N_11739,N_12346);
and U16813 (N_16813,N_13260,N_13897);
nand U16814 (N_16814,N_12507,N_12727);
nor U16815 (N_16815,N_12476,N_12217);
nand U16816 (N_16816,N_11797,N_13228);
nor U16817 (N_16817,N_13216,N_12284);
nor U16818 (N_16818,N_14189,N_11505);
and U16819 (N_16819,N_12862,N_14186);
nor U16820 (N_16820,N_12000,N_12449);
nor U16821 (N_16821,N_14227,N_14665);
or U16822 (N_16822,N_12826,N_12259);
nand U16823 (N_16823,N_14081,N_14226);
and U16824 (N_16824,N_12308,N_12062);
nand U16825 (N_16825,N_12016,N_11308);
and U16826 (N_16826,N_13324,N_13959);
and U16827 (N_16827,N_11344,N_13314);
or U16828 (N_16828,N_12025,N_13357);
or U16829 (N_16829,N_14139,N_14299);
or U16830 (N_16830,N_10619,N_12369);
or U16831 (N_16831,N_11149,N_14247);
or U16832 (N_16832,N_12182,N_13383);
and U16833 (N_16833,N_12497,N_12519);
nor U16834 (N_16834,N_14636,N_14309);
nor U16835 (N_16835,N_12757,N_11144);
nor U16836 (N_16836,N_10759,N_11008);
xnor U16837 (N_16837,N_12277,N_11199);
xnor U16838 (N_16838,N_11110,N_14203);
nor U16839 (N_16839,N_13082,N_11424);
xnor U16840 (N_16840,N_10538,N_14868);
nand U16841 (N_16841,N_12942,N_14985);
xnor U16842 (N_16842,N_13015,N_11341);
nand U16843 (N_16843,N_14590,N_13759);
nor U16844 (N_16844,N_13418,N_13124);
and U16845 (N_16845,N_11583,N_13345);
and U16846 (N_16846,N_14434,N_10112);
or U16847 (N_16847,N_12879,N_13323);
xor U16848 (N_16848,N_14132,N_11393);
and U16849 (N_16849,N_13761,N_10567);
or U16850 (N_16850,N_12616,N_13904);
xnor U16851 (N_16851,N_12742,N_14534);
xnor U16852 (N_16852,N_14607,N_13865);
or U16853 (N_16853,N_14069,N_10623);
xnor U16854 (N_16854,N_11467,N_10553);
nand U16855 (N_16855,N_11736,N_12685);
and U16856 (N_16856,N_13206,N_11023);
and U16857 (N_16857,N_10562,N_12335);
nor U16858 (N_16858,N_14794,N_12529);
nand U16859 (N_16859,N_14877,N_10452);
xor U16860 (N_16860,N_14644,N_14846);
and U16861 (N_16861,N_13623,N_11637);
and U16862 (N_16862,N_14159,N_10405);
or U16863 (N_16863,N_10493,N_10277);
xnor U16864 (N_16864,N_12895,N_13347);
nand U16865 (N_16865,N_10508,N_12071);
nor U16866 (N_16866,N_12251,N_10173);
nor U16867 (N_16867,N_14492,N_13562);
nor U16868 (N_16868,N_10833,N_12492);
and U16869 (N_16869,N_10684,N_12364);
or U16870 (N_16870,N_13038,N_12762);
xor U16871 (N_16871,N_12644,N_11587);
or U16872 (N_16872,N_13521,N_10261);
nand U16873 (N_16873,N_10488,N_11147);
and U16874 (N_16874,N_12164,N_12382);
and U16875 (N_16875,N_13596,N_11489);
nand U16876 (N_16876,N_14518,N_11333);
or U16877 (N_16877,N_11172,N_13421);
nand U16878 (N_16878,N_14129,N_13221);
nand U16879 (N_16879,N_10180,N_10458);
xnor U16880 (N_16880,N_12003,N_10557);
and U16881 (N_16881,N_13385,N_13825);
and U16882 (N_16882,N_13145,N_14705);
and U16883 (N_16883,N_11185,N_12307);
nand U16884 (N_16884,N_14367,N_12505);
or U16885 (N_16885,N_11837,N_13426);
nor U16886 (N_16886,N_10844,N_11890);
nand U16887 (N_16887,N_11687,N_10194);
nor U16888 (N_16888,N_13432,N_10868);
nor U16889 (N_16889,N_13690,N_14259);
and U16890 (N_16890,N_12885,N_13772);
and U16891 (N_16891,N_14000,N_13395);
nor U16892 (N_16892,N_11174,N_14261);
or U16893 (N_16893,N_12460,N_14882);
xnor U16894 (N_16894,N_14731,N_13059);
xnor U16895 (N_16895,N_14887,N_10162);
nor U16896 (N_16896,N_10767,N_12706);
or U16897 (N_16897,N_13268,N_14763);
or U16898 (N_16898,N_11330,N_12465);
nor U16899 (N_16899,N_14948,N_12195);
nor U16900 (N_16900,N_11705,N_10716);
xor U16901 (N_16901,N_10638,N_10439);
or U16902 (N_16902,N_14538,N_11007);
nand U16903 (N_16903,N_13552,N_13325);
xnor U16904 (N_16904,N_12272,N_11208);
or U16905 (N_16905,N_14422,N_12441);
nand U16906 (N_16906,N_12365,N_14815);
and U16907 (N_16907,N_12577,N_11336);
nor U16908 (N_16908,N_12822,N_11558);
nor U16909 (N_16909,N_12254,N_11967);
nor U16910 (N_16910,N_11603,N_13722);
or U16911 (N_16911,N_12515,N_11818);
nand U16912 (N_16912,N_12009,N_13092);
and U16913 (N_16913,N_13974,N_10819);
and U16914 (N_16914,N_14337,N_11464);
and U16915 (N_16915,N_14529,N_14523);
nor U16916 (N_16916,N_12545,N_14184);
nor U16917 (N_16917,N_13519,N_14919);
nor U16918 (N_16918,N_10426,N_14898);
and U16919 (N_16919,N_10861,N_11231);
nand U16920 (N_16920,N_13684,N_13707);
nand U16921 (N_16921,N_10306,N_14837);
xnor U16922 (N_16922,N_12426,N_10628);
or U16923 (N_16923,N_12391,N_12169);
or U16924 (N_16924,N_11449,N_14706);
nor U16925 (N_16925,N_12689,N_14716);
or U16926 (N_16926,N_12738,N_10783);
nor U16927 (N_16927,N_10656,N_13255);
and U16928 (N_16928,N_11405,N_11514);
nor U16929 (N_16929,N_11480,N_12785);
nor U16930 (N_16930,N_12716,N_10161);
nor U16931 (N_16931,N_13296,N_10027);
xor U16932 (N_16932,N_13911,N_13334);
xor U16933 (N_16933,N_12803,N_11138);
and U16934 (N_16934,N_12331,N_13634);
and U16935 (N_16935,N_10826,N_11175);
nand U16936 (N_16936,N_14588,N_11423);
nor U16937 (N_16937,N_14876,N_10943);
and U16938 (N_16938,N_13653,N_14387);
nor U16939 (N_16939,N_12106,N_14663);
nand U16940 (N_16940,N_14652,N_14907);
nand U16941 (N_16941,N_12487,N_14525);
or U16942 (N_16942,N_10800,N_13292);
nand U16943 (N_16943,N_13495,N_11991);
or U16944 (N_16944,N_10147,N_11803);
nor U16945 (N_16945,N_13069,N_13928);
nand U16946 (N_16946,N_13786,N_12784);
or U16947 (N_16947,N_11496,N_13471);
and U16948 (N_16948,N_10708,N_10086);
and U16949 (N_16949,N_13716,N_10730);
and U16950 (N_16950,N_12679,N_11492);
nor U16951 (N_16951,N_10531,N_12798);
or U16952 (N_16952,N_11606,N_10198);
or U16953 (N_16953,N_11112,N_13647);
or U16954 (N_16954,N_14916,N_11591);
nand U16955 (N_16955,N_12206,N_12111);
nor U16956 (N_16956,N_13040,N_11444);
xnor U16957 (N_16957,N_12566,N_13485);
nand U16958 (N_16958,N_12949,N_14252);
and U16959 (N_16959,N_11139,N_12498);
and U16960 (N_16960,N_13430,N_11058);
nand U16961 (N_16961,N_12291,N_14147);
or U16962 (N_16962,N_11427,N_13799);
xnor U16963 (N_16963,N_12583,N_14033);
nor U16964 (N_16964,N_14571,N_10665);
and U16965 (N_16965,N_14420,N_11270);
xor U16966 (N_16966,N_10111,N_11654);
and U16967 (N_16967,N_11795,N_12997);
nor U16968 (N_16968,N_14466,N_13767);
xnor U16969 (N_16969,N_11619,N_14845);
nand U16970 (N_16970,N_10572,N_11876);
xor U16971 (N_16971,N_13400,N_12002);
or U16972 (N_16972,N_13135,N_12929);
and U16973 (N_16973,N_11256,N_11501);
nor U16974 (N_16974,N_12157,N_14594);
nand U16975 (N_16975,N_11740,N_11824);
xor U16976 (N_16976,N_14011,N_14368);
and U16977 (N_16977,N_10774,N_14984);
nor U16978 (N_16978,N_12909,N_11888);
and U16979 (N_16979,N_13567,N_13391);
nor U16980 (N_16980,N_13836,N_13054);
nand U16981 (N_16981,N_10189,N_13749);
nor U16982 (N_16982,N_11539,N_12660);
or U16983 (N_16983,N_14072,N_10250);
or U16984 (N_16984,N_11406,N_10127);
or U16985 (N_16985,N_11068,N_10410);
or U16986 (N_16986,N_10461,N_14019);
or U16987 (N_16987,N_10850,N_13113);
and U16988 (N_16988,N_14753,N_12874);
or U16989 (N_16989,N_11425,N_14176);
or U16990 (N_16990,N_11894,N_12228);
nor U16991 (N_16991,N_12311,N_13472);
nand U16992 (N_16992,N_14050,N_10836);
nand U16993 (N_16993,N_14577,N_11418);
and U16994 (N_16994,N_13890,N_10710);
or U16995 (N_16995,N_11851,N_11337);
and U16996 (N_16996,N_10060,N_10969);
and U16997 (N_16997,N_11553,N_12471);
nand U16998 (N_16998,N_12079,N_10233);
nand U16999 (N_16999,N_12540,N_13843);
nand U17000 (N_17000,N_14990,N_12108);
or U17001 (N_17001,N_13918,N_14808);
and U17002 (N_17002,N_14005,N_12347);
nor U17003 (N_17003,N_12399,N_12018);
nor U17004 (N_17004,N_12219,N_10335);
nand U17005 (N_17005,N_11735,N_12444);
nand U17006 (N_17006,N_12980,N_11930);
or U17007 (N_17007,N_14971,N_11436);
xnor U17008 (N_17008,N_10544,N_12389);
or U17009 (N_17009,N_11277,N_13088);
xnor U17010 (N_17010,N_14075,N_14526);
nor U17011 (N_17011,N_14445,N_10183);
nor U17012 (N_17012,N_12589,N_13541);
nor U17013 (N_17013,N_14339,N_14210);
or U17014 (N_17014,N_13604,N_11681);
nand U17015 (N_17015,N_11000,N_13173);
or U17016 (N_17016,N_14294,N_14199);
or U17017 (N_17017,N_12853,N_14964);
nand U17018 (N_17018,N_12795,N_11771);
or U17019 (N_17019,N_12687,N_13635);
and U17020 (N_17020,N_10676,N_10464);
nor U17021 (N_17021,N_12409,N_11699);
nor U17022 (N_17022,N_14448,N_14629);
nor U17023 (N_17023,N_14651,N_12783);
nor U17024 (N_17024,N_11481,N_13741);
nand U17025 (N_17025,N_12380,N_10629);
nor U17026 (N_17026,N_11245,N_13202);
or U17027 (N_17027,N_11567,N_12688);
nor U17028 (N_17028,N_10092,N_13993);
and U17029 (N_17029,N_12216,N_12586);
nand U17030 (N_17030,N_11862,N_10903);
nor U17031 (N_17031,N_14757,N_12396);
or U17032 (N_17032,N_12058,N_13053);
xor U17033 (N_17033,N_13306,N_13428);
nor U17034 (N_17034,N_14981,N_10961);
nor U17035 (N_17035,N_10586,N_13700);
nand U17036 (N_17036,N_12668,N_13280);
and U17037 (N_17037,N_12852,N_13744);
nand U17038 (N_17038,N_13227,N_12914);
and U17039 (N_17039,N_10380,N_13536);
nor U17040 (N_17040,N_14198,N_10429);
and U17041 (N_17041,N_13087,N_14424);
nand U17042 (N_17042,N_11074,N_12925);
or U17043 (N_17043,N_11404,N_11696);
and U17044 (N_17044,N_14911,N_10216);
nand U17045 (N_17045,N_13275,N_13335);
or U17046 (N_17046,N_12207,N_13116);
and U17047 (N_17047,N_13646,N_14245);
nand U17048 (N_17048,N_14151,N_14804);
and U17049 (N_17049,N_14826,N_14113);
nand U17050 (N_17050,N_13752,N_14288);
nor U17051 (N_17051,N_10354,N_11835);
nor U17052 (N_17052,N_13338,N_10904);
xor U17053 (N_17053,N_12035,N_13998);
or U17054 (N_17054,N_14101,N_13151);
or U17055 (N_17055,N_10680,N_13251);
or U17056 (N_17056,N_11392,N_13535);
xnor U17057 (N_17057,N_10159,N_10546);
and U17058 (N_17058,N_11107,N_12238);
or U17059 (N_17059,N_13029,N_13222);
nand U17060 (N_17060,N_11620,N_10047);
or U17061 (N_17061,N_10153,N_14888);
nor U17062 (N_17062,N_10717,N_14762);
or U17063 (N_17063,N_13782,N_12902);
or U17064 (N_17064,N_11250,N_10530);
nand U17065 (N_17065,N_14120,N_10443);
or U17066 (N_17066,N_13672,N_10058);
or U17067 (N_17067,N_10874,N_14170);
nor U17068 (N_17068,N_13696,N_13181);
nor U17069 (N_17069,N_11734,N_13293);
and U17070 (N_17070,N_10616,N_12039);
and U17071 (N_17071,N_11882,N_10066);
and U17072 (N_17072,N_11048,N_12451);
nand U17073 (N_17073,N_11493,N_11361);
nor U17074 (N_17074,N_12983,N_10021);
or U17075 (N_17075,N_13414,N_10289);
or U17076 (N_17076,N_12462,N_10821);
or U17077 (N_17077,N_13340,N_11897);
nor U17078 (N_17078,N_11903,N_10455);
and U17079 (N_17079,N_11440,N_13045);
or U17080 (N_17080,N_12490,N_12595);
nor U17081 (N_17081,N_12184,N_14667);
nand U17082 (N_17082,N_13853,N_11516);
and U17083 (N_17083,N_13747,N_13068);
or U17084 (N_17084,N_10954,N_11692);
or U17085 (N_17085,N_11679,N_13709);
or U17086 (N_17086,N_11041,N_13190);
xnor U17087 (N_17087,N_11761,N_13710);
xor U17088 (N_17088,N_10197,N_14343);
nand U17089 (N_17089,N_13185,N_10927);
and U17090 (N_17090,N_11033,N_11264);
or U17091 (N_17091,N_10725,N_14354);
nor U17092 (N_17092,N_11542,N_11628);
nand U17093 (N_17093,N_14306,N_12596);
nand U17094 (N_17094,N_12410,N_11998);
or U17095 (N_17095,N_12173,N_12223);
and U17096 (N_17096,N_12006,N_14562);
or U17097 (N_17097,N_14207,N_10492);
or U17098 (N_17098,N_12068,N_12817);
and U17099 (N_17099,N_13802,N_10658);
xnor U17100 (N_17100,N_10673,N_12172);
or U17101 (N_17101,N_12836,N_12323);
nor U17102 (N_17102,N_12764,N_14047);
nand U17103 (N_17103,N_10615,N_10028);
nor U17104 (N_17104,N_13805,N_10433);
nand U17105 (N_17105,N_11087,N_10597);
xnor U17106 (N_17106,N_10651,N_10832);
nand U17107 (N_17107,N_13452,N_12056);
nand U17108 (N_17108,N_10096,N_12740);
nand U17109 (N_17109,N_12903,N_14265);
or U17110 (N_17110,N_14867,N_14690);
nand U17111 (N_17111,N_12239,N_14175);
xor U17112 (N_17112,N_11745,N_12340);
xnor U17113 (N_17113,N_11001,N_14191);
and U17114 (N_17114,N_11997,N_12209);
nor U17115 (N_17115,N_10657,N_10914);
nor U17116 (N_17116,N_13243,N_12458);
nor U17117 (N_17117,N_12939,N_14202);
and U17118 (N_17118,N_12114,N_12911);
and U17119 (N_17119,N_14556,N_14855);
nor U17120 (N_17120,N_11086,N_12260);
or U17121 (N_17121,N_10427,N_10698);
or U17122 (N_17122,N_14255,N_13757);
or U17123 (N_17123,N_14853,N_14416);
and U17124 (N_17124,N_11773,N_14978);
nor U17125 (N_17125,N_14662,N_11675);
and U17126 (N_17126,N_12450,N_14813);
nor U17127 (N_17127,N_11503,N_11918);
xor U17128 (N_17128,N_13220,N_12088);
and U17129 (N_17129,N_13442,N_13072);
nand U17130 (N_17130,N_11896,N_10863);
nor U17131 (N_17131,N_12303,N_13602);
nor U17132 (N_17132,N_12412,N_11917);
and U17133 (N_17133,N_12669,N_11331);
or U17134 (N_17134,N_12198,N_13854);
nor U17135 (N_17135,N_10110,N_12140);
nor U17136 (N_17136,N_14626,N_14812);
xnor U17137 (N_17137,N_12374,N_11340);
nor U17138 (N_17138,N_13119,N_12183);
nand U17139 (N_17139,N_13231,N_14780);
and U17140 (N_17140,N_12622,N_14349);
nor U17141 (N_17141,N_10026,N_12517);
nand U17142 (N_17142,N_14331,N_11137);
or U17143 (N_17143,N_10746,N_10123);
or U17144 (N_17144,N_13556,N_12625);
xnor U17145 (N_17145,N_11746,N_12425);
xor U17146 (N_17146,N_11893,N_13907);
nor U17147 (N_17147,N_11240,N_14512);
xnor U17148 (N_17148,N_11156,N_11512);
nand U17149 (N_17149,N_10263,N_14359);
nor U17150 (N_17150,N_13566,N_13844);
nor U17151 (N_17151,N_14473,N_14709);
or U17152 (N_17152,N_14355,N_11234);
nor U17153 (N_17153,N_14171,N_11853);
or U17154 (N_17154,N_12718,N_14880);
nor U17155 (N_17155,N_11373,N_12041);
nand U17156 (N_17156,N_11791,N_14883);
nand U17157 (N_17157,N_14917,N_13966);
and U17158 (N_17158,N_10987,N_12811);
and U17159 (N_17159,N_13937,N_12940);
or U17160 (N_17160,N_10539,N_12921);
xor U17161 (N_17161,N_12779,N_14082);
nand U17162 (N_17162,N_14836,N_12661);
nor U17163 (N_17163,N_14801,N_11313);
nand U17164 (N_17164,N_12493,N_14451);
nand U17165 (N_17165,N_14618,N_14362);
and U17166 (N_17166,N_12092,N_14795);
xor U17167 (N_17167,N_13656,N_11353);
or U17168 (N_17168,N_13644,N_10591);
and U17169 (N_17169,N_11753,N_11273);
and U17170 (N_17170,N_11640,N_13423);
and U17171 (N_17171,N_10934,N_12342);
nor U17172 (N_17172,N_12712,N_12139);
or U17173 (N_17173,N_13058,N_14270);
nand U17174 (N_17174,N_10408,N_11442);
xor U17175 (N_17175,N_10232,N_10485);
and U17176 (N_17176,N_13051,N_11482);
xnor U17177 (N_17177,N_13539,N_11378);
nand U17178 (N_17178,N_11911,N_13126);
xor U17179 (N_17179,N_13060,N_12244);
nand U17180 (N_17180,N_12899,N_12598);
and U17181 (N_17181,N_14275,N_13958);
nand U17182 (N_17182,N_12752,N_11575);
or U17183 (N_17183,N_10504,N_14127);
nor U17184 (N_17184,N_10976,N_10395);
nor U17185 (N_17185,N_10588,N_11235);
xor U17186 (N_17186,N_11446,N_10014);
or U17187 (N_17187,N_14772,N_12965);
nand U17188 (N_17188,N_14896,N_13011);
nor U17189 (N_17189,N_11443,N_11632);
nor U17190 (N_17190,N_11310,N_12818);
nand U17191 (N_17191,N_10300,N_10301);
xor U17192 (N_17192,N_13819,N_14477);
nand U17193 (N_17193,N_14394,N_11206);
nor U17194 (N_17194,N_12579,N_14515);
nor U17195 (N_17195,N_11004,N_14282);
or U17196 (N_17196,N_13117,N_13180);
or U17197 (N_17197,N_12960,N_10641);
nor U17198 (N_17198,N_12464,N_13988);
nor U17199 (N_17199,N_11677,N_14851);
and U17200 (N_17200,N_13509,N_12120);
or U17201 (N_17201,N_10678,N_12963);
nor U17202 (N_17202,N_10009,N_11438);
and U17203 (N_17203,N_13191,N_11034);
or U17204 (N_17204,N_10365,N_12481);
and U17205 (N_17205,N_13599,N_10945);
xnor U17206 (N_17206,N_12469,N_12105);
nand U17207 (N_17207,N_11799,N_14498);
or U17208 (N_17208,N_14861,N_12189);
or U17209 (N_17209,N_10274,N_13840);
nand U17210 (N_17210,N_14433,N_13500);
or U17211 (N_17211,N_14273,N_10499);
and U17212 (N_17212,N_11134,N_12456);
nand U17213 (N_17213,N_14001,N_12046);
xnor U17214 (N_17214,N_14061,N_10317);
nand U17215 (N_17215,N_12341,N_10926);
or U17216 (N_17216,N_11993,N_10463);
nand U17217 (N_17217,N_14637,N_10512);
or U17218 (N_17218,N_11246,N_10070);
nor U17219 (N_17219,N_11815,N_13265);
and U17220 (N_17220,N_12502,N_11187);
nand U17221 (N_17221,N_11394,N_12883);
and U17222 (N_17222,N_12012,N_13735);
or U17223 (N_17223,N_14680,N_11662);
nand U17224 (N_17224,N_12319,N_13504);
or U17225 (N_17225,N_13207,N_11682);
or U17226 (N_17226,N_11508,N_13833);
xor U17227 (N_17227,N_12411,N_14109);
or U17228 (N_17228,N_13502,N_13867);
nand U17229 (N_17229,N_14611,N_10998);
and U17230 (N_17230,N_11549,N_10687);
and U17231 (N_17231,N_11729,N_13737);
and U17232 (N_17232,N_10999,N_13917);
nor U17233 (N_17233,N_14327,N_10356);
and U17234 (N_17234,N_12132,N_11176);
and U17235 (N_17235,N_11576,N_14633);
nand U17236 (N_17236,N_11689,N_13597);
or U17237 (N_17237,N_10978,N_14223);
nand U17238 (N_17238,N_12917,N_13148);
and U17239 (N_17239,N_10346,N_13796);
or U17240 (N_17240,N_13598,N_13563);
xnor U17241 (N_17241,N_10570,N_13893);
or U17242 (N_17242,N_13286,N_11013);
or U17243 (N_17243,N_10169,N_12984);
and U17244 (N_17244,N_13518,N_12170);
nand U17245 (N_17245,N_10398,N_11829);
and U17246 (N_17246,N_11209,N_11779);
nor U17247 (N_17247,N_13736,N_10912);
nor U17248 (N_17248,N_14773,N_14089);
or U17249 (N_17249,N_13902,N_13377);
or U17250 (N_17250,N_13934,N_10185);
nand U17251 (N_17251,N_14374,N_12286);
or U17252 (N_17252,N_10705,N_12355);
nor U17253 (N_17253,N_13913,N_14467);
nor U17254 (N_17254,N_11292,N_10442);
or U17255 (N_17255,N_10670,N_11497);
or U17256 (N_17256,N_10170,N_13676);
or U17257 (N_17257,N_10231,N_11972);
nor U17258 (N_17258,N_11935,N_11384);
nand U17259 (N_17259,N_10672,N_14241);
nor U17260 (N_17260,N_12810,N_13241);
nor U17261 (N_17261,N_12873,N_11598);
and U17262 (N_17262,N_10453,N_10158);
nor U17263 (N_17263,N_14735,N_13030);
xnor U17264 (N_17264,N_10694,N_14935);
and U17265 (N_17265,N_13713,N_11494);
and U17266 (N_17266,N_13090,N_12436);
or U17267 (N_17267,N_14476,N_10882);
or U17268 (N_17268,N_14840,N_10820);
nor U17269 (N_17269,N_11343,N_14719);
and U17270 (N_17270,N_14599,N_13109);
nand U17271 (N_17271,N_14344,N_12344);
nand U17272 (N_17272,N_10901,N_14943);
xor U17273 (N_17273,N_13507,N_12847);
nand U17274 (N_17274,N_14987,N_12845);
and U17275 (N_17275,N_13530,N_14673);
and U17276 (N_17276,N_10720,N_10845);
nand U17277 (N_17277,N_12787,N_14703);
or U17278 (N_17278,N_10138,N_11357);
nand U17279 (N_17279,N_11002,N_12969);
nor U17280 (N_17280,N_10005,N_10337);
or U17281 (N_17281,N_11817,N_13288);
nand U17282 (N_17282,N_11305,N_11711);
nor U17283 (N_17283,N_13662,N_10760);
and U17284 (N_17284,N_13760,N_12691);
and U17285 (N_17285,N_10726,N_12318);
or U17286 (N_17286,N_11828,N_11532);
xor U17287 (N_17287,N_12648,N_11981);
and U17288 (N_17288,N_14212,N_12551);
nor U17289 (N_17289,N_10188,N_12890);
xnor U17290 (N_17290,N_13792,N_11029);
xnor U17291 (N_17291,N_10311,N_12871);
or U17292 (N_17292,N_12749,N_11989);
or U17293 (N_17293,N_13123,N_10609);
or U17294 (N_17294,N_10603,N_12666);
and U17295 (N_17295,N_11921,N_13271);
nand U17296 (N_17296,N_14630,N_12912);
and U17297 (N_17297,N_11578,N_13062);
nand U17298 (N_17298,N_14654,N_12618);
and U17299 (N_17299,N_14039,N_11724);
nand U17300 (N_17300,N_10940,N_12633);
and U17301 (N_17301,N_11171,N_11266);
nand U17302 (N_17302,N_10121,N_11018);
nor U17303 (N_17303,N_13997,N_10480);
nand U17304 (N_17304,N_13701,N_12368);
and U17305 (N_17305,N_12773,N_12603);
nor U17306 (N_17306,N_11915,N_13930);
nand U17307 (N_17307,N_11038,N_12587);
and U17308 (N_17308,N_10293,N_14745);
or U17309 (N_17309,N_14116,N_14041);
and U17310 (N_17310,N_13332,N_13477);
xnor U17311 (N_17311,N_13884,N_11479);
nor U17312 (N_17312,N_14281,N_13664);
nor U17313 (N_17313,N_13870,N_10292);
nor U17314 (N_17314,N_12834,N_14126);
and U17315 (N_17315,N_13637,N_13311);
nor U17316 (N_17316,N_11316,N_11293);
nor U17317 (N_17317,N_12082,N_11457);
nand U17318 (N_17318,N_13924,N_10235);
or U17319 (N_17319,N_11473,N_10654);
and U17320 (N_17320,N_11939,N_10298);
and U17321 (N_17321,N_10265,N_14154);
xnor U17322 (N_17322,N_14504,N_11759);
and U17323 (N_17323,N_12127,N_11046);
nand U17324 (N_17324,N_12667,N_11971);
nand U17325 (N_17325,N_10724,N_13447);
and U17326 (N_17326,N_11192,N_14942);
and U17327 (N_17327,N_11650,N_11362);
nor U17328 (N_17328,N_13146,N_13641);
or U17329 (N_17329,N_12232,N_14704);
nand U17330 (N_17330,N_11188,N_11190);
nor U17331 (N_17331,N_11460,N_11224);
and U17332 (N_17332,N_10010,N_12447);
nand U17333 (N_17333,N_11322,N_14300);
nand U17334 (N_17334,N_11878,N_12072);
nor U17335 (N_17335,N_14712,N_10637);
and U17336 (N_17336,N_13308,N_12524);
nor U17337 (N_17337,N_13724,N_12080);
or U17338 (N_17338,N_10700,N_10144);
nand U17339 (N_17339,N_13025,N_14271);
and U17340 (N_17340,N_10279,N_12060);
or U17341 (N_17341,N_11334,N_13121);
and U17342 (N_17342,N_12095,N_11133);
and U17343 (N_17343,N_12937,N_10647);
and U17344 (N_17344,N_12213,N_13144);
nand U17345 (N_17345,N_10668,N_12992);
nor U17346 (N_17346,N_14123,N_14436);
nand U17347 (N_17347,N_11335,N_13838);
nand U17348 (N_17348,N_11265,N_13929);
xor U17349 (N_17349,N_10511,N_12148);
and U17350 (N_17350,N_10972,N_13841);
or U17351 (N_17351,N_13580,N_12537);
xor U17352 (N_17352,N_12163,N_11821);
and U17353 (N_17353,N_14839,N_14623);
and U17354 (N_17354,N_11150,N_14465);
and U17355 (N_17355,N_12248,N_12768);
nand U17356 (N_17356,N_10655,N_10171);
and U17357 (N_17357,N_12770,N_14456);
or U17358 (N_17358,N_10568,N_11158);
nand U17359 (N_17359,N_13654,N_13373);
and U17360 (N_17360,N_11051,N_13137);
nor U17361 (N_17361,N_13992,N_14054);
nand U17362 (N_17362,N_14783,N_10791);
nand U17363 (N_17363,N_11920,N_12278);
xnor U17364 (N_17364,N_10140,N_12614);
and U17365 (N_17365,N_12313,N_13336);
or U17366 (N_17366,N_10210,N_12647);
nand U17367 (N_17367,N_13797,N_12774);
or U17368 (N_17368,N_12185,N_14505);
or U17369 (N_17369,N_11928,N_13140);
and U17370 (N_17370,N_10938,N_13688);
nand U17371 (N_17371,N_14040,N_14068);
or U17372 (N_17372,N_13842,N_13704);
or U17373 (N_17373,N_13405,N_14471);
and U17374 (N_17374,N_10025,N_11432);
nand U17375 (N_17375,N_14357,N_14012);
xnor U17376 (N_17376,N_12884,N_14400);
and U17377 (N_17377,N_10131,N_11140);
nor U17378 (N_17378,N_12835,N_11025);
nand U17379 (N_17379,N_11880,N_12878);
and U17380 (N_17380,N_11995,N_12655);
or U17381 (N_17381,N_14490,N_14440);
and U17382 (N_17382,N_13079,N_13147);
and U17383 (N_17383,N_14233,N_14778);
nand U17384 (N_17384,N_13349,N_13494);
and U17385 (N_17385,N_12208,N_10340);
or U17386 (N_17386,N_11402,N_14540);
nor U17387 (N_17387,N_10041,N_13691);
nor U17388 (N_17388,N_10117,N_13467);
nand U17389 (N_17389,N_11641,N_14912);
xor U17390 (N_17390,N_11130,N_13174);
or U17391 (N_17391,N_13305,N_10176);
xnor U17392 (N_17392,N_14627,N_10519);
nand U17393 (N_17393,N_13501,N_13885);
or U17394 (N_17394,N_12571,N_12461);
or U17395 (N_17395,N_10880,N_11420);
and U17396 (N_17396,N_14543,N_10937);
or U17397 (N_17397,N_13302,N_13665);
nand U17398 (N_17398,N_11869,N_11852);
xor U17399 (N_17399,N_10611,N_11577);
and U17400 (N_17400,N_11656,N_14321);
xnor U17401 (N_17401,N_13845,N_10794);
nand U17402 (N_17402,N_14338,N_10124);
nor U17403 (N_17403,N_11506,N_12455);
or U17404 (N_17404,N_10219,N_11860);
and U17405 (N_17405,N_11645,N_11560);
nand U17406 (N_17406,N_10878,N_11298);
or U17407 (N_17407,N_13449,N_13727);
or U17408 (N_17408,N_14581,N_10168);
nand U17409 (N_17409,N_10902,N_10412);
or U17410 (N_17410,N_13272,N_14934);
or U17411 (N_17411,N_12070,N_12581);
and U17412 (N_17412,N_10001,N_11244);
or U17413 (N_17413,N_10212,N_10848);
nor U17414 (N_17414,N_11718,N_10478);
nand U17415 (N_17415,N_14714,N_11097);
nor U17416 (N_17416,N_13601,N_12824);
nand U17417 (N_17417,N_10995,N_14506);
or U17418 (N_17418,N_13269,N_12429);
or U17419 (N_17419,N_11535,N_14138);
nand U17420 (N_17420,N_14258,N_10951);
nor U17421 (N_17421,N_12575,N_11604);
nor U17422 (N_17422,N_14635,N_13531);
nor U17423 (N_17423,N_10738,N_10084);
nor U17424 (N_17424,N_12199,N_14474);
or U17425 (N_17425,N_12846,N_11768);
and U17426 (N_17426,N_14449,N_14872);
or U17427 (N_17427,N_10377,N_13299);
nor U17428 (N_17428,N_14550,N_13194);
or U17429 (N_17429,N_12491,N_14646);
nor U17430 (N_17430,N_11827,N_11477);
nor U17431 (N_17431,N_11345,N_13080);
nor U17432 (N_17432,N_11066,N_13115);
nand U17433 (N_17433,N_12838,N_14702);
xor U17434 (N_17434,N_13573,N_12664);
and U17435 (N_17435,N_13954,N_10149);
nor U17436 (N_17436,N_11456,N_11887);
or U17437 (N_17437,N_11317,N_11468);
and U17438 (N_17438,N_14014,N_12790);
nor U17439 (N_17439,N_11790,N_11355);
and U17440 (N_17440,N_10515,N_11990);
and U17441 (N_17441,N_13661,N_12708);
or U17442 (N_17442,N_14320,N_12124);
or U17443 (N_17443,N_10155,N_14643);
or U17444 (N_17444,N_12629,N_12485);
and U17445 (N_17445,N_13520,N_13892);
and U17446 (N_17446,N_11380,N_14664);
nor U17447 (N_17447,N_13464,N_10348);
nand U17448 (N_17448,N_10890,N_10810);
nand U17449 (N_17449,N_14782,N_12008);
or U17450 (N_17450,N_14267,N_13553);
nor U17451 (N_17451,N_10727,N_14620);
nor U17452 (N_17452,N_14053,N_13962);
nand U17453 (N_17453,N_12872,N_11236);
nor U17454 (N_17454,N_12289,N_13955);
or U17455 (N_17455,N_14342,N_14497);
nand U17456 (N_17456,N_12956,N_13003);
and U17457 (N_17457,N_10105,N_10524);
or U17458 (N_17458,N_10777,N_10450);
nand U17459 (N_17459,N_13923,N_12281);
and U17460 (N_17460,N_11924,N_11125);
nor U17461 (N_17461,N_10556,N_11919);
or U17462 (N_17462,N_11354,N_10985);
or U17463 (N_17463,N_14668,N_11132);
or U17464 (N_17464,N_14439,N_11842);
and U17465 (N_17465,N_11665,N_11861);
or U17466 (N_17466,N_10491,N_12147);
or U17467 (N_17467,N_14820,N_12792);
and U17468 (N_17468,N_12404,N_11426);
and U17469 (N_17469,N_14125,N_13990);
nand U17470 (N_17470,N_10474,N_14071);
nand U17471 (N_17471,N_14216,N_13263);
nor U17472 (N_17472,N_12483,N_13497);
or U17473 (N_17473,N_13878,N_11182);
and U17474 (N_17474,N_12472,N_14494);
nand U17475 (N_17475,N_11800,N_12705);
or U17476 (N_17476,N_12171,N_11557);
and U17477 (N_17477,N_12298,N_10766);
nand U17478 (N_17478,N_14201,N_11726);
nand U17479 (N_17479,N_13066,N_14423);
nand U17480 (N_17480,N_13198,N_13419);
nor U17481 (N_17481,N_12179,N_13103);
and U17482 (N_17482,N_14969,N_12038);
xnor U17483 (N_17483,N_11618,N_14679);
nor U17484 (N_17484,N_14566,N_14580);
and U17485 (N_17485,N_13189,N_12736);
nand U17486 (N_17486,N_14383,N_11070);
xnor U17487 (N_17487,N_13777,N_14560);
nand U17488 (N_17488,N_14746,N_13905);
xor U17489 (N_17489,N_13358,N_13908);
nor U17490 (N_17490,N_11747,N_11220);
and U17491 (N_17491,N_12336,N_13132);
nand U17492 (N_17492,N_14642,N_14484);
xnor U17493 (N_17493,N_13125,N_10403);
and U17494 (N_17494,N_14486,N_11363);
nor U17495 (N_17495,N_13574,N_13968);
and U17496 (N_17496,N_10510,N_10661);
and U17497 (N_17497,N_12442,N_11081);
nand U17498 (N_17498,N_13919,N_11238);
nand U17499 (N_17499,N_11474,N_14708);
and U17500 (N_17500,N_13172,N_12545);
xnor U17501 (N_17501,N_10595,N_10475);
nor U17502 (N_17502,N_10387,N_14902);
or U17503 (N_17503,N_12620,N_10544);
and U17504 (N_17504,N_14439,N_13155);
nor U17505 (N_17505,N_13055,N_12250);
nand U17506 (N_17506,N_14127,N_12976);
nand U17507 (N_17507,N_11475,N_14806);
nor U17508 (N_17508,N_14560,N_11585);
nor U17509 (N_17509,N_14893,N_14386);
xor U17510 (N_17510,N_13832,N_13642);
nor U17511 (N_17511,N_12318,N_14857);
xnor U17512 (N_17512,N_11825,N_14636);
nor U17513 (N_17513,N_10911,N_13475);
or U17514 (N_17514,N_12405,N_14145);
nor U17515 (N_17515,N_14205,N_12191);
or U17516 (N_17516,N_14637,N_10896);
xnor U17517 (N_17517,N_10795,N_11122);
and U17518 (N_17518,N_11565,N_12222);
nor U17519 (N_17519,N_11060,N_11478);
and U17520 (N_17520,N_10624,N_10701);
and U17521 (N_17521,N_14990,N_12678);
nand U17522 (N_17522,N_14826,N_13592);
and U17523 (N_17523,N_14268,N_11564);
nand U17524 (N_17524,N_13944,N_12514);
or U17525 (N_17525,N_13342,N_14044);
nand U17526 (N_17526,N_13270,N_12444);
and U17527 (N_17527,N_11415,N_13158);
nor U17528 (N_17528,N_11815,N_11048);
or U17529 (N_17529,N_13757,N_13887);
nor U17530 (N_17530,N_11336,N_13279);
nand U17531 (N_17531,N_10444,N_13386);
nor U17532 (N_17532,N_10498,N_14814);
xor U17533 (N_17533,N_14554,N_13397);
or U17534 (N_17534,N_14518,N_14958);
or U17535 (N_17535,N_14788,N_12886);
nand U17536 (N_17536,N_12695,N_12092);
nand U17537 (N_17537,N_10563,N_14575);
nor U17538 (N_17538,N_14648,N_13083);
and U17539 (N_17539,N_12018,N_12492);
nor U17540 (N_17540,N_10791,N_11039);
nor U17541 (N_17541,N_10504,N_14900);
and U17542 (N_17542,N_12570,N_14630);
nor U17543 (N_17543,N_14264,N_14407);
and U17544 (N_17544,N_11276,N_10450);
and U17545 (N_17545,N_12469,N_14908);
xnor U17546 (N_17546,N_12942,N_13014);
and U17547 (N_17547,N_13613,N_10757);
nand U17548 (N_17548,N_12101,N_10793);
nand U17549 (N_17549,N_13365,N_14043);
nand U17550 (N_17550,N_11339,N_10718);
or U17551 (N_17551,N_10272,N_11391);
or U17552 (N_17552,N_12267,N_13850);
nand U17553 (N_17553,N_13989,N_13723);
nor U17554 (N_17554,N_10130,N_13877);
nor U17555 (N_17555,N_12721,N_11683);
nand U17556 (N_17556,N_13160,N_13332);
and U17557 (N_17557,N_14020,N_12486);
nor U17558 (N_17558,N_14270,N_14294);
nor U17559 (N_17559,N_13325,N_12496);
nor U17560 (N_17560,N_12215,N_11519);
or U17561 (N_17561,N_14793,N_10490);
and U17562 (N_17562,N_10114,N_13840);
nand U17563 (N_17563,N_10293,N_12366);
xnor U17564 (N_17564,N_13741,N_14040);
nand U17565 (N_17565,N_10789,N_11952);
xor U17566 (N_17566,N_10368,N_10479);
nor U17567 (N_17567,N_12873,N_11222);
nor U17568 (N_17568,N_11586,N_11680);
or U17569 (N_17569,N_12887,N_11132);
xnor U17570 (N_17570,N_13795,N_14636);
or U17571 (N_17571,N_13797,N_13812);
nand U17572 (N_17572,N_10005,N_10244);
and U17573 (N_17573,N_13194,N_14466);
or U17574 (N_17574,N_11474,N_12689);
and U17575 (N_17575,N_14180,N_10693);
xor U17576 (N_17576,N_14476,N_14269);
or U17577 (N_17577,N_14833,N_12326);
nor U17578 (N_17578,N_12833,N_14891);
or U17579 (N_17579,N_12739,N_14147);
xnor U17580 (N_17580,N_10117,N_13610);
nand U17581 (N_17581,N_14240,N_14092);
xor U17582 (N_17582,N_14322,N_11237);
nor U17583 (N_17583,N_10896,N_10012);
or U17584 (N_17584,N_14886,N_12429);
nor U17585 (N_17585,N_14691,N_10505);
or U17586 (N_17586,N_12483,N_12679);
and U17587 (N_17587,N_14340,N_11567);
or U17588 (N_17588,N_13363,N_10274);
or U17589 (N_17589,N_12138,N_14007);
or U17590 (N_17590,N_11456,N_10670);
xnor U17591 (N_17591,N_12935,N_12293);
xnor U17592 (N_17592,N_14866,N_11194);
or U17593 (N_17593,N_13196,N_12917);
nand U17594 (N_17594,N_11031,N_12894);
and U17595 (N_17595,N_13202,N_13785);
and U17596 (N_17596,N_13218,N_14005);
and U17597 (N_17597,N_14605,N_13348);
and U17598 (N_17598,N_10413,N_10206);
or U17599 (N_17599,N_11104,N_10170);
nand U17600 (N_17600,N_14286,N_11132);
or U17601 (N_17601,N_14511,N_14166);
or U17602 (N_17602,N_10801,N_13401);
xnor U17603 (N_17603,N_13154,N_12883);
xnor U17604 (N_17604,N_10632,N_11441);
nor U17605 (N_17605,N_13550,N_13021);
and U17606 (N_17606,N_11291,N_13260);
nor U17607 (N_17607,N_11712,N_13738);
or U17608 (N_17608,N_11977,N_13725);
nor U17609 (N_17609,N_10583,N_14822);
nor U17610 (N_17610,N_14684,N_13692);
nand U17611 (N_17611,N_11514,N_11228);
nor U17612 (N_17612,N_13801,N_10073);
and U17613 (N_17613,N_13342,N_10679);
xor U17614 (N_17614,N_10354,N_11920);
and U17615 (N_17615,N_14785,N_11682);
xnor U17616 (N_17616,N_12619,N_13511);
nand U17617 (N_17617,N_11859,N_12699);
nor U17618 (N_17618,N_13025,N_11210);
or U17619 (N_17619,N_10044,N_14707);
or U17620 (N_17620,N_12979,N_13203);
nand U17621 (N_17621,N_13307,N_13970);
nor U17622 (N_17622,N_11286,N_10252);
nor U17623 (N_17623,N_10374,N_11975);
and U17624 (N_17624,N_11871,N_14611);
or U17625 (N_17625,N_13541,N_13328);
or U17626 (N_17626,N_14688,N_14887);
nor U17627 (N_17627,N_12894,N_11178);
nand U17628 (N_17628,N_11294,N_14365);
or U17629 (N_17629,N_10767,N_13022);
and U17630 (N_17630,N_12987,N_11668);
nand U17631 (N_17631,N_10923,N_11682);
nor U17632 (N_17632,N_14593,N_12856);
nor U17633 (N_17633,N_11448,N_11900);
or U17634 (N_17634,N_11073,N_11172);
and U17635 (N_17635,N_11197,N_10638);
nor U17636 (N_17636,N_14739,N_14348);
and U17637 (N_17637,N_13661,N_10278);
or U17638 (N_17638,N_12986,N_10027);
nor U17639 (N_17639,N_13383,N_10017);
xor U17640 (N_17640,N_13153,N_10273);
nor U17641 (N_17641,N_14442,N_10964);
and U17642 (N_17642,N_10140,N_14006);
and U17643 (N_17643,N_14640,N_12593);
nand U17644 (N_17644,N_10163,N_10921);
or U17645 (N_17645,N_12330,N_14050);
and U17646 (N_17646,N_11675,N_13875);
and U17647 (N_17647,N_13830,N_12973);
xnor U17648 (N_17648,N_13348,N_12369);
or U17649 (N_17649,N_14157,N_10158);
xnor U17650 (N_17650,N_12905,N_13124);
xnor U17651 (N_17651,N_14644,N_12124);
nand U17652 (N_17652,N_11466,N_13839);
nand U17653 (N_17653,N_11842,N_11459);
nor U17654 (N_17654,N_14972,N_10115);
or U17655 (N_17655,N_11300,N_10849);
nor U17656 (N_17656,N_14514,N_11948);
and U17657 (N_17657,N_11387,N_12958);
nand U17658 (N_17658,N_14084,N_10810);
nand U17659 (N_17659,N_11540,N_11217);
nand U17660 (N_17660,N_12529,N_14046);
nor U17661 (N_17661,N_14264,N_13523);
and U17662 (N_17662,N_12719,N_10044);
xor U17663 (N_17663,N_13965,N_12678);
nand U17664 (N_17664,N_13539,N_10564);
nor U17665 (N_17665,N_10103,N_14169);
xor U17666 (N_17666,N_12711,N_14461);
nor U17667 (N_17667,N_13861,N_11094);
and U17668 (N_17668,N_11966,N_14765);
xnor U17669 (N_17669,N_11820,N_10367);
and U17670 (N_17670,N_11783,N_11299);
nor U17671 (N_17671,N_12632,N_12268);
and U17672 (N_17672,N_11807,N_14222);
or U17673 (N_17673,N_10266,N_12755);
and U17674 (N_17674,N_14120,N_11543);
or U17675 (N_17675,N_12859,N_11811);
or U17676 (N_17676,N_13278,N_11160);
nand U17677 (N_17677,N_13335,N_14361);
and U17678 (N_17678,N_13361,N_12829);
nand U17679 (N_17679,N_11038,N_13268);
and U17680 (N_17680,N_11860,N_10446);
and U17681 (N_17681,N_14308,N_13709);
and U17682 (N_17682,N_11947,N_11850);
or U17683 (N_17683,N_11481,N_13845);
and U17684 (N_17684,N_11979,N_13891);
and U17685 (N_17685,N_12315,N_14302);
nand U17686 (N_17686,N_14409,N_10330);
or U17687 (N_17687,N_14691,N_13204);
nor U17688 (N_17688,N_12945,N_14246);
or U17689 (N_17689,N_10648,N_13914);
or U17690 (N_17690,N_14407,N_11978);
xnor U17691 (N_17691,N_11621,N_12350);
nor U17692 (N_17692,N_11048,N_14949);
nand U17693 (N_17693,N_12106,N_11775);
nand U17694 (N_17694,N_11341,N_14957);
and U17695 (N_17695,N_14278,N_13132);
nor U17696 (N_17696,N_11944,N_14666);
nor U17697 (N_17697,N_10090,N_11152);
and U17698 (N_17698,N_12947,N_13085);
and U17699 (N_17699,N_10791,N_10707);
and U17700 (N_17700,N_14788,N_13422);
or U17701 (N_17701,N_11831,N_11944);
nor U17702 (N_17702,N_11396,N_12023);
nand U17703 (N_17703,N_11793,N_14644);
and U17704 (N_17704,N_11278,N_11120);
nand U17705 (N_17705,N_10396,N_14013);
xnor U17706 (N_17706,N_13204,N_12550);
and U17707 (N_17707,N_10037,N_13501);
nand U17708 (N_17708,N_11806,N_14493);
xor U17709 (N_17709,N_10698,N_10453);
nand U17710 (N_17710,N_11855,N_13251);
nand U17711 (N_17711,N_14305,N_13176);
and U17712 (N_17712,N_14227,N_11061);
nand U17713 (N_17713,N_12856,N_13111);
nor U17714 (N_17714,N_13433,N_10793);
nand U17715 (N_17715,N_10489,N_13444);
or U17716 (N_17716,N_14965,N_12044);
nor U17717 (N_17717,N_11038,N_13172);
nor U17718 (N_17718,N_10779,N_10174);
nand U17719 (N_17719,N_13323,N_11399);
nor U17720 (N_17720,N_13863,N_13928);
and U17721 (N_17721,N_12238,N_10488);
nor U17722 (N_17722,N_14496,N_12528);
nor U17723 (N_17723,N_13765,N_12706);
nor U17724 (N_17724,N_12813,N_12442);
and U17725 (N_17725,N_12398,N_12169);
xor U17726 (N_17726,N_12240,N_11766);
nand U17727 (N_17727,N_12073,N_10626);
and U17728 (N_17728,N_14653,N_12705);
or U17729 (N_17729,N_13561,N_10812);
xor U17730 (N_17730,N_10313,N_14620);
nor U17731 (N_17731,N_14870,N_11447);
nand U17732 (N_17732,N_11011,N_12432);
or U17733 (N_17733,N_10687,N_12821);
nor U17734 (N_17734,N_13719,N_14014);
and U17735 (N_17735,N_10504,N_14514);
nor U17736 (N_17736,N_13845,N_11241);
nor U17737 (N_17737,N_13636,N_12679);
and U17738 (N_17738,N_12100,N_14289);
and U17739 (N_17739,N_10459,N_11648);
or U17740 (N_17740,N_12860,N_14991);
nor U17741 (N_17741,N_14848,N_11508);
nor U17742 (N_17742,N_11533,N_10033);
nand U17743 (N_17743,N_14405,N_14617);
and U17744 (N_17744,N_10331,N_10197);
and U17745 (N_17745,N_11224,N_14807);
or U17746 (N_17746,N_10300,N_12032);
nand U17747 (N_17747,N_10990,N_10198);
nand U17748 (N_17748,N_10452,N_13283);
nand U17749 (N_17749,N_14503,N_14259);
and U17750 (N_17750,N_13093,N_10028);
or U17751 (N_17751,N_13753,N_13470);
or U17752 (N_17752,N_10338,N_11465);
or U17753 (N_17753,N_12200,N_13302);
or U17754 (N_17754,N_13046,N_10122);
xor U17755 (N_17755,N_12349,N_10598);
or U17756 (N_17756,N_12467,N_12972);
or U17757 (N_17757,N_11945,N_13066);
and U17758 (N_17758,N_13960,N_13829);
and U17759 (N_17759,N_12586,N_12846);
or U17760 (N_17760,N_13909,N_10754);
nand U17761 (N_17761,N_12913,N_12680);
and U17762 (N_17762,N_13209,N_13911);
nand U17763 (N_17763,N_12494,N_13981);
or U17764 (N_17764,N_13312,N_14482);
or U17765 (N_17765,N_14201,N_12127);
and U17766 (N_17766,N_12706,N_10401);
or U17767 (N_17767,N_13835,N_11670);
nand U17768 (N_17768,N_14471,N_13958);
nand U17769 (N_17769,N_10373,N_13070);
or U17770 (N_17770,N_10902,N_14677);
nand U17771 (N_17771,N_13799,N_11047);
nor U17772 (N_17772,N_11779,N_14036);
or U17773 (N_17773,N_13942,N_10402);
or U17774 (N_17774,N_11415,N_11597);
or U17775 (N_17775,N_10553,N_12728);
xor U17776 (N_17776,N_11572,N_12380);
nand U17777 (N_17777,N_14575,N_14000);
nand U17778 (N_17778,N_10800,N_11601);
nand U17779 (N_17779,N_13296,N_12261);
or U17780 (N_17780,N_11652,N_14432);
nor U17781 (N_17781,N_14247,N_14682);
nand U17782 (N_17782,N_10973,N_13846);
nand U17783 (N_17783,N_11746,N_13268);
and U17784 (N_17784,N_13281,N_10868);
nand U17785 (N_17785,N_10166,N_11353);
or U17786 (N_17786,N_13311,N_14092);
nand U17787 (N_17787,N_10400,N_12796);
and U17788 (N_17788,N_12959,N_11968);
nand U17789 (N_17789,N_12675,N_11479);
nand U17790 (N_17790,N_13923,N_13941);
nand U17791 (N_17791,N_12297,N_14126);
and U17792 (N_17792,N_13976,N_10460);
or U17793 (N_17793,N_10705,N_14650);
nand U17794 (N_17794,N_11241,N_13663);
nor U17795 (N_17795,N_10496,N_13011);
nand U17796 (N_17796,N_12822,N_10345);
nand U17797 (N_17797,N_10292,N_13665);
nor U17798 (N_17798,N_12473,N_12720);
and U17799 (N_17799,N_11591,N_10538);
nor U17800 (N_17800,N_14544,N_13942);
nor U17801 (N_17801,N_12912,N_13622);
xor U17802 (N_17802,N_11478,N_10675);
and U17803 (N_17803,N_12069,N_12790);
or U17804 (N_17804,N_14876,N_13630);
and U17805 (N_17805,N_12284,N_11834);
nand U17806 (N_17806,N_10973,N_10430);
or U17807 (N_17807,N_11318,N_13114);
and U17808 (N_17808,N_12607,N_10900);
or U17809 (N_17809,N_12068,N_13240);
or U17810 (N_17810,N_12659,N_12986);
xnor U17811 (N_17811,N_14179,N_10741);
nor U17812 (N_17812,N_12460,N_10649);
and U17813 (N_17813,N_10433,N_13896);
and U17814 (N_17814,N_11433,N_13522);
and U17815 (N_17815,N_12422,N_11812);
and U17816 (N_17816,N_12918,N_11283);
or U17817 (N_17817,N_11593,N_12892);
xor U17818 (N_17818,N_14214,N_14422);
and U17819 (N_17819,N_14137,N_13954);
nand U17820 (N_17820,N_10753,N_10018);
and U17821 (N_17821,N_11514,N_13149);
nand U17822 (N_17822,N_12623,N_11048);
and U17823 (N_17823,N_11046,N_10604);
or U17824 (N_17824,N_12596,N_14140);
nand U17825 (N_17825,N_14203,N_13443);
nand U17826 (N_17826,N_12772,N_12272);
nand U17827 (N_17827,N_11583,N_13543);
nor U17828 (N_17828,N_11906,N_12832);
nand U17829 (N_17829,N_12418,N_10102);
nand U17830 (N_17830,N_14259,N_13239);
or U17831 (N_17831,N_12267,N_10457);
nor U17832 (N_17832,N_10939,N_13501);
nor U17833 (N_17833,N_13920,N_13489);
xor U17834 (N_17834,N_13664,N_10937);
nand U17835 (N_17835,N_14162,N_14285);
nor U17836 (N_17836,N_13839,N_14031);
or U17837 (N_17837,N_11498,N_14781);
nand U17838 (N_17838,N_12261,N_10943);
and U17839 (N_17839,N_14295,N_12073);
xnor U17840 (N_17840,N_14474,N_13827);
nor U17841 (N_17841,N_10515,N_10044);
nor U17842 (N_17842,N_12930,N_10537);
nand U17843 (N_17843,N_14818,N_10985);
or U17844 (N_17844,N_11942,N_13903);
or U17845 (N_17845,N_13175,N_14587);
nand U17846 (N_17846,N_12678,N_14639);
and U17847 (N_17847,N_12929,N_13161);
and U17848 (N_17848,N_10095,N_11169);
and U17849 (N_17849,N_11428,N_13483);
and U17850 (N_17850,N_11914,N_10775);
nand U17851 (N_17851,N_10810,N_11697);
and U17852 (N_17852,N_12909,N_12908);
xnor U17853 (N_17853,N_10869,N_13967);
nor U17854 (N_17854,N_13083,N_10555);
and U17855 (N_17855,N_12063,N_12944);
nand U17856 (N_17856,N_13580,N_12203);
and U17857 (N_17857,N_13776,N_14537);
nor U17858 (N_17858,N_11759,N_11888);
nand U17859 (N_17859,N_14450,N_11234);
nand U17860 (N_17860,N_11884,N_14266);
nor U17861 (N_17861,N_14500,N_14305);
or U17862 (N_17862,N_13725,N_10102);
nand U17863 (N_17863,N_13149,N_10739);
nor U17864 (N_17864,N_13008,N_13415);
or U17865 (N_17865,N_13385,N_13752);
nor U17866 (N_17866,N_13413,N_10146);
xor U17867 (N_17867,N_10494,N_11729);
nor U17868 (N_17868,N_10884,N_11278);
and U17869 (N_17869,N_13029,N_13060);
or U17870 (N_17870,N_11356,N_12902);
and U17871 (N_17871,N_14380,N_14372);
or U17872 (N_17872,N_12533,N_14537);
and U17873 (N_17873,N_13733,N_11014);
and U17874 (N_17874,N_11188,N_11511);
and U17875 (N_17875,N_13245,N_11456);
nand U17876 (N_17876,N_13670,N_10385);
xor U17877 (N_17877,N_13202,N_11072);
nor U17878 (N_17878,N_11008,N_13222);
nand U17879 (N_17879,N_10787,N_14487);
nor U17880 (N_17880,N_10057,N_10637);
nand U17881 (N_17881,N_13332,N_12456);
nor U17882 (N_17882,N_13509,N_11887);
or U17883 (N_17883,N_13099,N_11296);
and U17884 (N_17884,N_14700,N_14268);
or U17885 (N_17885,N_13101,N_14879);
and U17886 (N_17886,N_13801,N_10676);
nand U17887 (N_17887,N_10876,N_11182);
nor U17888 (N_17888,N_14904,N_12646);
xor U17889 (N_17889,N_13985,N_13304);
nor U17890 (N_17890,N_11528,N_10950);
nor U17891 (N_17891,N_14765,N_10415);
nand U17892 (N_17892,N_14160,N_10390);
and U17893 (N_17893,N_14385,N_14738);
nand U17894 (N_17894,N_14366,N_11421);
nor U17895 (N_17895,N_10519,N_10170);
and U17896 (N_17896,N_12701,N_10208);
and U17897 (N_17897,N_11509,N_12148);
nor U17898 (N_17898,N_14251,N_14478);
and U17899 (N_17899,N_12414,N_14476);
nand U17900 (N_17900,N_14451,N_12708);
nor U17901 (N_17901,N_13726,N_13753);
xnor U17902 (N_17902,N_12015,N_11866);
and U17903 (N_17903,N_10875,N_11720);
or U17904 (N_17904,N_14842,N_14924);
or U17905 (N_17905,N_14160,N_10566);
xnor U17906 (N_17906,N_14093,N_13713);
nor U17907 (N_17907,N_14761,N_12252);
and U17908 (N_17908,N_11461,N_12111);
or U17909 (N_17909,N_14806,N_10655);
xor U17910 (N_17910,N_14765,N_13886);
nor U17911 (N_17911,N_14352,N_10518);
and U17912 (N_17912,N_12788,N_14262);
and U17913 (N_17913,N_12416,N_13253);
nor U17914 (N_17914,N_12471,N_10759);
xnor U17915 (N_17915,N_14206,N_12383);
and U17916 (N_17916,N_12330,N_10847);
or U17917 (N_17917,N_12788,N_14784);
nor U17918 (N_17918,N_12547,N_13895);
or U17919 (N_17919,N_13077,N_12050);
and U17920 (N_17920,N_12593,N_12337);
nor U17921 (N_17921,N_14120,N_10937);
nand U17922 (N_17922,N_13519,N_11732);
or U17923 (N_17923,N_13985,N_11338);
nand U17924 (N_17924,N_14786,N_14603);
nand U17925 (N_17925,N_12894,N_12893);
or U17926 (N_17926,N_12489,N_10216);
and U17927 (N_17927,N_12118,N_10532);
nand U17928 (N_17928,N_14649,N_14769);
nor U17929 (N_17929,N_10848,N_14199);
nor U17930 (N_17930,N_12696,N_11633);
and U17931 (N_17931,N_11999,N_13796);
nand U17932 (N_17932,N_14657,N_11340);
and U17933 (N_17933,N_12650,N_10559);
xnor U17934 (N_17934,N_12904,N_14643);
nor U17935 (N_17935,N_12371,N_10417);
nand U17936 (N_17936,N_11958,N_10056);
nor U17937 (N_17937,N_14343,N_14620);
or U17938 (N_17938,N_14721,N_11138);
xnor U17939 (N_17939,N_13461,N_11594);
nor U17940 (N_17940,N_10545,N_13947);
nor U17941 (N_17941,N_12847,N_14280);
nand U17942 (N_17942,N_13267,N_10801);
or U17943 (N_17943,N_13521,N_10872);
nand U17944 (N_17944,N_11899,N_11935);
xnor U17945 (N_17945,N_12911,N_12467);
or U17946 (N_17946,N_12754,N_13743);
and U17947 (N_17947,N_11484,N_10358);
xnor U17948 (N_17948,N_13715,N_14315);
or U17949 (N_17949,N_14206,N_11479);
nor U17950 (N_17950,N_13197,N_11686);
nor U17951 (N_17951,N_12069,N_10346);
xnor U17952 (N_17952,N_12063,N_13271);
nand U17953 (N_17953,N_10108,N_10190);
nor U17954 (N_17954,N_13296,N_11295);
and U17955 (N_17955,N_11794,N_10403);
nor U17956 (N_17956,N_13048,N_10588);
nor U17957 (N_17957,N_13392,N_12744);
or U17958 (N_17958,N_12737,N_13384);
and U17959 (N_17959,N_13830,N_13588);
and U17960 (N_17960,N_12118,N_13721);
and U17961 (N_17961,N_13959,N_12790);
and U17962 (N_17962,N_10209,N_13353);
or U17963 (N_17963,N_12287,N_14822);
nand U17964 (N_17964,N_11780,N_10368);
and U17965 (N_17965,N_12576,N_14603);
and U17966 (N_17966,N_12775,N_13473);
nand U17967 (N_17967,N_10279,N_14112);
nand U17968 (N_17968,N_13106,N_10151);
nand U17969 (N_17969,N_12103,N_10946);
and U17970 (N_17970,N_13449,N_10937);
nor U17971 (N_17971,N_11451,N_14635);
nand U17972 (N_17972,N_10517,N_11555);
nand U17973 (N_17973,N_10474,N_12296);
or U17974 (N_17974,N_13397,N_13439);
nor U17975 (N_17975,N_12654,N_10468);
and U17976 (N_17976,N_13361,N_14426);
nor U17977 (N_17977,N_11733,N_14251);
or U17978 (N_17978,N_11206,N_11604);
nor U17979 (N_17979,N_13075,N_13422);
nand U17980 (N_17980,N_10015,N_10750);
nand U17981 (N_17981,N_12614,N_10854);
xor U17982 (N_17982,N_11245,N_10275);
and U17983 (N_17983,N_14513,N_10617);
nor U17984 (N_17984,N_14823,N_14259);
or U17985 (N_17985,N_11230,N_14486);
or U17986 (N_17986,N_10118,N_11576);
or U17987 (N_17987,N_14922,N_10976);
xnor U17988 (N_17988,N_12688,N_10365);
xnor U17989 (N_17989,N_13254,N_11358);
nor U17990 (N_17990,N_13064,N_13572);
or U17991 (N_17991,N_13788,N_11239);
or U17992 (N_17992,N_13716,N_13901);
and U17993 (N_17993,N_13645,N_14994);
xor U17994 (N_17994,N_13894,N_11059);
nand U17995 (N_17995,N_11750,N_14544);
xnor U17996 (N_17996,N_12167,N_14775);
or U17997 (N_17997,N_11508,N_14520);
nor U17998 (N_17998,N_13813,N_13417);
or U17999 (N_17999,N_13628,N_14376);
or U18000 (N_18000,N_11763,N_12829);
nand U18001 (N_18001,N_11443,N_11541);
xnor U18002 (N_18002,N_14815,N_10245);
and U18003 (N_18003,N_13756,N_10690);
xor U18004 (N_18004,N_12071,N_13800);
nor U18005 (N_18005,N_10010,N_11963);
or U18006 (N_18006,N_10482,N_13056);
and U18007 (N_18007,N_11977,N_14838);
nand U18008 (N_18008,N_14170,N_13747);
nor U18009 (N_18009,N_11991,N_12604);
or U18010 (N_18010,N_10897,N_10562);
nand U18011 (N_18011,N_12767,N_13007);
nor U18012 (N_18012,N_11784,N_14645);
nand U18013 (N_18013,N_13860,N_12384);
and U18014 (N_18014,N_12195,N_13975);
nand U18015 (N_18015,N_14728,N_13404);
or U18016 (N_18016,N_13165,N_13203);
nor U18017 (N_18017,N_10657,N_10362);
or U18018 (N_18018,N_11763,N_11215);
nor U18019 (N_18019,N_12345,N_11354);
nor U18020 (N_18020,N_12447,N_12764);
nor U18021 (N_18021,N_11416,N_14163);
and U18022 (N_18022,N_14733,N_12808);
nand U18023 (N_18023,N_11147,N_10333);
or U18024 (N_18024,N_14267,N_14364);
and U18025 (N_18025,N_13469,N_13849);
and U18026 (N_18026,N_11671,N_10890);
nor U18027 (N_18027,N_14486,N_10442);
nand U18028 (N_18028,N_12984,N_14026);
nor U18029 (N_18029,N_10452,N_13678);
nand U18030 (N_18030,N_13282,N_12212);
nor U18031 (N_18031,N_10702,N_11041);
nand U18032 (N_18032,N_13286,N_10987);
nand U18033 (N_18033,N_14311,N_13596);
nor U18034 (N_18034,N_11746,N_14755);
nand U18035 (N_18035,N_11174,N_14610);
nand U18036 (N_18036,N_10924,N_12145);
or U18037 (N_18037,N_10641,N_11757);
xor U18038 (N_18038,N_11102,N_13948);
and U18039 (N_18039,N_13679,N_13696);
xnor U18040 (N_18040,N_14056,N_10033);
nor U18041 (N_18041,N_13300,N_11530);
nand U18042 (N_18042,N_14451,N_11742);
xnor U18043 (N_18043,N_12797,N_10707);
and U18044 (N_18044,N_13744,N_10545);
nand U18045 (N_18045,N_10359,N_12728);
xor U18046 (N_18046,N_12184,N_11439);
nor U18047 (N_18047,N_12527,N_13660);
or U18048 (N_18048,N_13526,N_12254);
xor U18049 (N_18049,N_10844,N_11112);
nor U18050 (N_18050,N_13224,N_11755);
or U18051 (N_18051,N_12902,N_13609);
nor U18052 (N_18052,N_14475,N_10950);
or U18053 (N_18053,N_12836,N_10608);
or U18054 (N_18054,N_11648,N_11214);
nand U18055 (N_18055,N_11844,N_12057);
or U18056 (N_18056,N_14016,N_14785);
and U18057 (N_18057,N_12795,N_11647);
xnor U18058 (N_18058,N_12787,N_10932);
or U18059 (N_18059,N_12078,N_13210);
or U18060 (N_18060,N_12217,N_12514);
nand U18061 (N_18061,N_11613,N_12091);
xor U18062 (N_18062,N_13704,N_11242);
and U18063 (N_18063,N_11430,N_10150);
nor U18064 (N_18064,N_14683,N_10088);
or U18065 (N_18065,N_11847,N_10576);
nand U18066 (N_18066,N_12684,N_13035);
and U18067 (N_18067,N_10380,N_12437);
nand U18068 (N_18068,N_10007,N_13074);
nor U18069 (N_18069,N_11370,N_13758);
and U18070 (N_18070,N_12207,N_14587);
and U18071 (N_18071,N_12562,N_12332);
and U18072 (N_18072,N_12576,N_14791);
nand U18073 (N_18073,N_12810,N_11979);
nand U18074 (N_18074,N_13859,N_12050);
nand U18075 (N_18075,N_12419,N_11505);
or U18076 (N_18076,N_11548,N_14864);
nand U18077 (N_18077,N_10362,N_13950);
and U18078 (N_18078,N_12684,N_14943);
xor U18079 (N_18079,N_14630,N_12813);
nor U18080 (N_18080,N_12130,N_10888);
xor U18081 (N_18081,N_14815,N_11755);
nor U18082 (N_18082,N_12871,N_10617);
and U18083 (N_18083,N_11025,N_10395);
nor U18084 (N_18084,N_12096,N_11239);
or U18085 (N_18085,N_12210,N_12638);
xnor U18086 (N_18086,N_13473,N_13829);
or U18087 (N_18087,N_14541,N_10339);
xor U18088 (N_18088,N_12741,N_11529);
and U18089 (N_18089,N_12109,N_13052);
nand U18090 (N_18090,N_10815,N_11322);
and U18091 (N_18091,N_14257,N_10245);
xor U18092 (N_18092,N_12762,N_14184);
and U18093 (N_18093,N_12730,N_13985);
nand U18094 (N_18094,N_12603,N_12058);
or U18095 (N_18095,N_10694,N_14538);
nor U18096 (N_18096,N_11913,N_13000);
nor U18097 (N_18097,N_13179,N_12874);
or U18098 (N_18098,N_13477,N_10742);
nand U18099 (N_18099,N_11746,N_10125);
nor U18100 (N_18100,N_11921,N_10419);
xnor U18101 (N_18101,N_14908,N_10104);
nor U18102 (N_18102,N_13144,N_11186);
or U18103 (N_18103,N_14613,N_12315);
nor U18104 (N_18104,N_10856,N_10888);
nand U18105 (N_18105,N_10923,N_13622);
and U18106 (N_18106,N_11002,N_10230);
and U18107 (N_18107,N_14770,N_13356);
nor U18108 (N_18108,N_11908,N_13406);
nand U18109 (N_18109,N_12709,N_11448);
nor U18110 (N_18110,N_14150,N_12477);
and U18111 (N_18111,N_11104,N_11246);
nor U18112 (N_18112,N_12118,N_13578);
or U18113 (N_18113,N_12283,N_10623);
nor U18114 (N_18114,N_13663,N_11334);
nand U18115 (N_18115,N_10471,N_10174);
nand U18116 (N_18116,N_10509,N_10607);
nand U18117 (N_18117,N_13387,N_12040);
and U18118 (N_18118,N_14927,N_10644);
nand U18119 (N_18119,N_10492,N_14623);
xor U18120 (N_18120,N_14208,N_12196);
and U18121 (N_18121,N_10876,N_14982);
and U18122 (N_18122,N_12275,N_11576);
nor U18123 (N_18123,N_11757,N_13051);
nand U18124 (N_18124,N_14858,N_11376);
and U18125 (N_18125,N_13621,N_14374);
or U18126 (N_18126,N_10833,N_11689);
nand U18127 (N_18127,N_11444,N_12866);
nor U18128 (N_18128,N_10981,N_12643);
nor U18129 (N_18129,N_13454,N_10476);
nand U18130 (N_18130,N_11531,N_11864);
or U18131 (N_18131,N_13787,N_10083);
or U18132 (N_18132,N_10642,N_14340);
and U18133 (N_18133,N_11920,N_11106);
nor U18134 (N_18134,N_12933,N_13618);
nand U18135 (N_18135,N_12990,N_11809);
nor U18136 (N_18136,N_13575,N_12924);
nand U18137 (N_18137,N_12546,N_12796);
xor U18138 (N_18138,N_14546,N_11685);
nor U18139 (N_18139,N_11110,N_12222);
nor U18140 (N_18140,N_10005,N_12264);
and U18141 (N_18141,N_12677,N_11428);
nand U18142 (N_18142,N_13816,N_14233);
or U18143 (N_18143,N_10231,N_11163);
nor U18144 (N_18144,N_10331,N_12648);
and U18145 (N_18145,N_11089,N_13440);
nor U18146 (N_18146,N_13615,N_13501);
nand U18147 (N_18147,N_10801,N_14783);
or U18148 (N_18148,N_11804,N_14667);
and U18149 (N_18149,N_11380,N_10293);
nor U18150 (N_18150,N_11243,N_12986);
nand U18151 (N_18151,N_12400,N_12803);
nand U18152 (N_18152,N_11807,N_10653);
and U18153 (N_18153,N_14395,N_11498);
and U18154 (N_18154,N_12055,N_12324);
xnor U18155 (N_18155,N_11114,N_14515);
nand U18156 (N_18156,N_10654,N_10441);
and U18157 (N_18157,N_10510,N_13506);
or U18158 (N_18158,N_13125,N_11018);
or U18159 (N_18159,N_14836,N_10640);
and U18160 (N_18160,N_12860,N_10575);
nand U18161 (N_18161,N_12682,N_10529);
nor U18162 (N_18162,N_14103,N_12648);
nor U18163 (N_18163,N_12678,N_13476);
and U18164 (N_18164,N_11989,N_13443);
nand U18165 (N_18165,N_12196,N_12814);
xnor U18166 (N_18166,N_13186,N_14245);
nor U18167 (N_18167,N_13569,N_11228);
nor U18168 (N_18168,N_11309,N_12652);
or U18169 (N_18169,N_10695,N_11945);
or U18170 (N_18170,N_12266,N_11243);
nand U18171 (N_18171,N_14212,N_13950);
nor U18172 (N_18172,N_11604,N_11674);
nor U18173 (N_18173,N_12245,N_10746);
nand U18174 (N_18174,N_11161,N_14615);
or U18175 (N_18175,N_10119,N_14224);
or U18176 (N_18176,N_13203,N_11623);
nand U18177 (N_18177,N_12471,N_12971);
or U18178 (N_18178,N_10081,N_10139);
nor U18179 (N_18179,N_13282,N_14231);
xor U18180 (N_18180,N_13348,N_10511);
or U18181 (N_18181,N_14150,N_12629);
nand U18182 (N_18182,N_12211,N_14671);
nor U18183 (N_18183,N_11183,N_11235);
nand U18184 (N_18184,N_11268,N_11481);
xor U18185 (N_18185,N_12273,N_14191);
or U18186 (N_18186,N_11639,N_11398);
nand U18187 (N_18187,N_11574,N_14592);
and U18188 (N_18188,N_12348,N_13459);
or U18189 (N_18189,N_11313,N_13179);
nor U18190 (N_18190,N_13654,N_14751);
nand U18191 (N_18191,N_12785,N_10401);
and U18192 (N_18192,N_12191,N_14497);
nor U18193 (N_18193,N_12660,N_10728);
nand U18194 (N_18194,N_10961,N_14073);
nand U18195 (N_18195,N_10927,N_12843);
nor U18196 (N_18196,N_10503,N_13802);
or U18197 (N_18197,N_14023,N_11745);
or U18198 (N_18198,N_14909,N_11445);
and U18199 (N_18199,N_12775,N_14056);
and U18200 (N_18200,N_11221,N_10903);
nand U18201 (N_18201,N_13362,N_14552);
xnor U18202 (N_18202,N_13385,N_11757);
and U18203 (N_18203,N_14154,N_14751);
nand U18204 (N_18204,N_12344,N_12342);
and U18205 (N_18205,N_14141,N_14496);
nor U18206 (N_18206,N_11682,N_10593);
nand U18207 (N_18207,N_12300,N_12994);
and U18208 (N_18208,N_12041,N_11444);
nand U18209 (N_18209,N_10852,N_13924);
and U18210 (N_18210,N_10495,N_12146);
nand U18211 (N_18211,N_11879,N_12451);
nand U18212 (N_18212,N_10511,N_11350);
xor U18213 (N_18213,N_13737,N_13151);
nand U18214 (N_18214,N_13249,N_12607);
nand U18215 (N_18215,N_14391,N_13504);
or U18216 (N_18216,N_10750,N_10315);
or U18217 (N_18217,N_11643,N_10563);
and U18218 (N_18218,N_12051,N_11594);
and U18219 (N_18219,N_11128,N_12025);
xnor U18220 (N_18220,N_13808,N_10643);
xnor U18221 (N_18221,N_14445,N_10340);
or U18222 (N_18222,N_12213,N_10637);
nor U18223 (N_18223,N_13978,N_11517);
nand U18224 (N_18224,N_11412,N_11528);
nand U18225 (N_18225,N_10493,N_14115);
xor U18226 (N_18226,N_12517,N_13240);
and U18227 (N_18227,N_12021,N_10006);
nor U18228 (N_18228,N_13207,N_14299);
and U18229 (N_18229,N_10972,N_12711);
and U18230 (N_18230,N_14286,N_13682);
or U18231 (N_18231,N_13718,N_10419);
and U18232 (N_18232,N_13699,N_13779);
nand U18233 (N_18233,N_10374,N_13366);
nand U18234 (N_18234,N_10251,N_11083);
and U18235 (N_18235,N_11245,N_10650);
or U18236 (N_18236,N_13646,N_11124);
or U18237 (N_18237,N_10303,N_13690);
nand U18238 (N_18238,N_12991,N_12857);
and U18239 (N_18239,N_11852,N_10008);
nor U18240 (N_18240,N_10063,N_12311);
or U18241 (N_18241,N_11551,N_14297);
nand U18242 (N_18242,N_11711,N_13075);
and U18243 (N_18243,N_14685,N_14402);
nor U18244 (N_18244,N_10103,N_13454);
and U18245 (N_18245,N_11115,N_13847);
or U18246 (N_18246,N_14659,N_14981);
nand U18247 (N_18247,N_10611,N_14811);
nor U18248 (N_18248,N_12811,N_14112);
nand U18249 (N_18249,N_13675,N_12529);
nor U18250 (N_18250,N_14845,N_14594);
nor U18251 (N_18251,N_14000,N_14479);
and U18252 (N_18252,N_10818,N_12042);
nor U18253 (N_18253,N_11510,N_13604);
nand U18254 (N_18254,N_10435,N_10874);
or U18255 (N_18255,N_12642,N_14614);
or U18256 (N_18256,N_12627,N_10984);
xnor U18257 (N_18257,N_14803,N_11347);
and U18258 (N_18258,N_11102,N_13848);
or U18259 (N_18259,N_12052,N_11934);
or U18260 (N_18260,N_13842,N_10285);
or U18261 (N_18261,N_13923,N_10339);
nand U18262 (N_18262,N_13334,N_11285);
and U18263 (N_18263,N_14358,N_11725);
or U18264 (N_18264,N_13354,N_14650);
and U18265 (N_18265,N_11543,N_14035);
xnor U18266 (N_18266,N_12852,N_14568);
nor U18267 (N_18267,N_13176,N_13704);
nand U18268 (N_18268,N_11092,N_12050);
nand U18269 (N_18269,N_14416,N_10167);
and U18270 (N_18270,N_13891,N_14047);
nor U18271 (N_18271,N_14927,N_11896);
nand U18272 (N_18272,N_12575,N_11633);
and U18273 (N_18273,N_11452,N_11512);
xnor U18274 (N_18274,N_14058,N_12085);
nand U18275 (N_18275,N_12474,N_14725);
xor U18276 (N_18276,N_14363,N_12560);
nor U18277 (N_18277,N_11265,N_13453);
and U18278 (N_18278,N_11332,N_13493);
nor U18279 (N_18279,N_14402,N_13838);
nand U18280 (N_18280,N_14369,N_11262);
nor U18281 (N_18281,N_11188,N_13640);
and U18282 (N_18282,N_14457,N_13766);
or U18283 (N_18283,N_13858,N_10657);
nor U18284 (N_18284,N_11536,N_12290);
and U18285 (N_18285,N_12154,N_11698);
nand U18286 (N_18286,N_14077,N_10860);
nand U18287 (N_18287,N_10569,N_14752);
nand U18288 (N_18288,N_12882,N_11651);
or U18289 (N_18289,N_12085,N_12102);
or U18290 (N_18290,N_10307,N_13153);
or U18291 (N_18291,N_13013,N_14433);
nor U18292 (N_18292,N_12456,N_13340);
nor U18293 (N_18293,N_13457,N_11537);
or U18294 (N_18294,N_11406,N_13719);
nand U18295 (N_18295,N_12775,N_12465);
or U18296 (N_18296,N_13713,N_12417);
nor U18297 (N_18297,N_14498,N_14743);
or U18298 (N_18298,N_13023,N_12481);
nand U18299 (N_18299,N_10808,N_10903);
or U18300 (N_18300,N_11170,N_10328);
nor U18301 (N_18301,N_14868,N_11501);
nor U18302 (N_18302,N_10361,N_14235);
xnor U18303 (N_18303,N_11204,N_12707);
nor U18304 (N_18304,N_10866,N_10253);
or U18305 (N_18305,N_14038,N_12232);
nor U18306 (N_18306,N_12209,N_13124);
xor U18307 (N_18307,N_10975,N_10093);
or U18308 (N_18308,N_11894,N_13578);
nor U18309 (N_18309,N_12891,N_11438);
xor U18310 (N_18310,N_14878,N_11229);
nor U18311 (N_18311,N_14280,N_12781);
or U18312 (N_18312,N_11727,N_14286);
or U18313 (N_18313,N_10691,N_10720);
and U18314 (N_18314,N_10148,N_13830);
nand U18315 (N_18315,N_12603,N_13870);
nand U18316 (N_18316,N_12685,N_13485);
nor U18317 (N_18317,N_11366,N_10855);
nand U18318 (N_18318,N_13239,N_11058);
nand U18319 (N_18319,N_11163,N_12627);
nand U18320 (N_18320,N_12298,N_10542);
nor U18321 (N_18321,N_14719,N_13983);
nand U18322 (N_18322,N_13295,N_14295);
xnor U18323 (N_18323,N_13219,N_11890);
nand U18324 (N_18324,N_12674,N_10289);
xor U18325 (N_18325,N_11488,N_10188);
or U18326 (N_18326,N_14114,N_11320);
or U18327 (N_18327,N_13680,N_11316);
nor U18328 (N_18328,N_12102,N_14766);
and U18329 (N_18329,N_10982,N_10062);
nor U18330 (N_18330,N_13975,N_14067);
nor U18331 (N_18331,N_11470,N_11173);
or U18332 (N_18332,N_11895,N_14469);
and U18333 (N_18333,N_11245,N_13461);
xor U18334 (N_18334,N_12514,N_11476);
nor U18335 (N_18335,N_11932,N_14185);
or U18336 (N_18336,N_14468,N_11040);
nand U18337 (N_18337,N_10336,N_12087);
or U18338 (N_18338,N_14321,N_10683);
or U18339 (N_18339,N_10974,N_12428);
nand U18340 (N_18340,N_12570,N_12389);
nor U18341 (N_18341,N_11203,N_12309);
and U18342 (N_18342,N_12217,N_11616);
nand U18343 (N_18343,N_12193,N_10970);
and U18344 (N_18344,N_10054,N_14448);
xnor U18345 (N_18345,N_11776,N_13640);
and U18346 (N_18346,N_13396,N_11904);
nand U18347 (N_18347,N_14423,N_13918);
xnor U18348 (N_18348,N_10039,N_11617);
xor U18349 (N_18349,N_11850,N_10494);
or U18350 (N_18350,N_12856,N_11235);
nor U18351 (N_18351,N_11807,N_13580);
nor U18352 (N_18352,N_13637,N_13236);
nor U18353 (N_18353,N_12552,N_12271);
nor U18354 (N_18354,N_13878,N_11444);
nor U18355 (N_18355,N_13094,N_13720);
nor U18356 (N_18356,N_12531,N_14345);
or U18357 (N_18357,N_12835,N_11120);
or U18358 (N_18358,N_13860,N_13174);
and U18359 (N_18359,N_11933,N_14554);
and U18360 (N_18360,N_10146,N_12104);
nor U18361 (N_18361,N_12367,N_11347);
and U18362 (N_18362,N_10703,N_12044);
nor U18363 (N_18363,N_12693,N_12247);
and U18364 (N_18364,N_13873,N_10307);
and U18365 (N_18365,N_14169,N_10578);
nand U18366 (N_18366,N_13791,N_12891);
xor U18367 (N_18367,N_12502,N_12103);
or U18368 (N_18368,N_13417,N_13068);
and U18369 (N_18369,N_10660,N_14526);
nor U18370 (N_18370,N_11107,N_12391);
and U18371 (N_18371,N_13336,N_13199);
nand U18372 (N_18372,N_13739,N_11346);
and U18373 (N_18373,N_14655,N_12459);
nand U18374 (N_18374,N_11025,N_11880);
and U18375 (N_18375,N_13501,N_14740);
nand U18376 (N_18376,N_12325,N_10644);
xor U18377 (N_18377,N_10024,N_13445);
and U18378 (N_18378,N_13522,N_10091);
and U18379 (N_18379,N_10208,N_11271);
and U18380 (N_18380,N_10877,N_12827);
or U18381 (N_18381,N_10489,N_14039);
or U18382 (N_18382,N_11932,N_12756);
xor U18383 (N_18383,N_14449,N_12524);
nand U18384 (N_18384,N_14030,N_13941);
or U18385 (N_18385,N_10681,N_14150);
and U18386 (N_18386,N_13446,N_11216);
or U18387 (N_18387,N_14838,N_11668);
or U18388 (N_18388,N_10566,N_12612);
and U18389 (N_18389,N_13042,N_11141);
nand U18390 (N_18390,N_12169,N_12890);
and U18391 (N_18391,N_11012,N_12542);
nand U18392 (N_18392,N_14855,N_12851);
or U18393 (N_18393,N_10887,N_10979);
and U18394 (N_18394,N_14637,N_14721);
and U18395 (N_18395,N_13468,N_13300);
and U18396 (N_18396,N_10612,N_10688);
and U18397 (N_18397,N_10755,N_13548);
or U18398 (N_18398,N_13602,N_12425);
nand U18399 (N_18399,N_12606,N_14991);
or U18400 (N_18400,N_10404,N_10494);
or U18401 (N_18401,N_12703,N_10461);
or U18402 (N_18402,N_12102,N_10844);
xor U18403 (N_18403,N_12577,N_14581);
or U18404 (N_18404,N_13459,N_12899);
nand U18405 (N_18405,N_11519,N_13160);
nand U18406 (N_18406,N_11311,N_13863);
nand U18407 (N_18407,N_10864,N_10297);
and U18408 (N_18408,N_10237,N_14988);
nand U18409 (N_18409,N_12642,N_10909);
nor U18410 (N_18410,N_11435,N_13796);
and U18411 (N_18411,N_11031,N_14339);
or U18412 (N_18412,N_10244,N_10946);
nand U18413 (N_18413,N_13734,N_11618);
nand U18414 (N_18414,N_11740,N_11434);
or U18415 (N_18415,N_13777,N_13111);
or U18416 (N_18416,N_12662,N_11821);
and U18417 (N_18417,N_14091,N_11521);
nand U18418 (N_18418,N_14418,N_13119);
nand U18419 (N_18419,N_13462,N_10079);
or U18420 (N_18420,N_13551,N_11792);
nand U18421 (N_18421,N_10757,N_13132);
and U18422 (N_18422,N_14364,N_10244);
and U18423 (N_18423,N_12837,N_14168);
nand U18424 (N_18424,N_12010,N_12891);
nor U18425 (N_18425,N_11957,N_13140);
and U18426 (N_18426,N_11966,N_13259);
nor U18427 (N_18427,N_10120,N_11015);
nor U18428 (N_18428,N_10926,N_12637);
nand U18429 (N_18429,N_12297,N_14278);
and U18430 (N_18430,N_13742,N_12262);
nand U18431 (N_18431,N_11966,N_11719);
or U18432 (N_18432,N_10877,N_11531);
nor U18433 (N_18433,N_10383,N_11630);
nor U18434 (N_18434,N_12275,N_10609);
and U18435 (N_18435,N_12357,N_13771);
and U18436 (N_18436,N_11092,N_11292);
and U18437 (N_18437,N_12002,N_11347);
and U18438 (N_18438,N_11286,N_12268);
nor U18439 (N_18439,N_14277,N_10267);
or U18440 (N_18440,N_12104,N_11125);
nor U18441 (N_18441,N_10358,N_10338);
or U18442 (N_18442,N_10075,N_14070);
and U18443 (N_18443,N_10275,N_13972);
or U18444 (N_18444,N_11415,N_13364);
and U18445 (N_18445,N_14685,N_10740);
nor U18446 (N_18446,N_11653,N_10520);
nor U18447 (N_18447,N_11938,N_12923);
xnor U18448 (N_18448,N_12669,N_13998);
xor U18449 (N_18449,N_14213,N_10150);
xnor U18450 (N_18450,N_10452,N_14858);
nand U18451 (N_18451,N_14726,N_14929);
or U18452 (N_18452,N_10576,N_11373);
nand U18453 (N_18453,N_12990,N_13787);
nand U18454 (N_18454,N_10482,N_13804);
nand U18455 (N_18455,N_10697,N_12515);
or U18456 (N_18456,N_13623,N_10849);
nor U18457 (N_18457,N_12539,N_13975);
or U18458 (N_18458,N_10945,N_11081);
or U18459 (N_18459,N_14025,N_11618);
nand U18460 (N_18460,N_12132,N_14847);
and U18461 (N_18461,N_10450,N_13674);
or U18462 (N_18462,N_14830,N_14259);
nand U18463 (N_18463,N_10777,N_10536);
and U18464 (N_18464,N_11615,N_10273);
nor U18465 (N_18465,N_11521,N_14937);
and U18466 (N_18466,N_13595,N_13096);
and U18467 (N_18467,N_10638,N_10721);
and U18468 (N_18468,N_10425,N_11812);
or U18469 (N_18469,N_11136,N_14331);
and U18470 (N_18470,N_11062,N_12466);
xnor U18471 (N_18471,N_10337,N_10783);
and U18472 (N_18472,N_12866,N_13783);
nand U18473 (N_18473,N_14702,N_11641);
and U18474 (N_18474,N_14289,N_13816);
nand U18475 (N_18475,N_11707,N_14501);
nor U18476 (N_18476,N_13873,N_13816);
nand U18477 (N_18477,N_11743,N_10128);
nand U18478 (N_18478,N_14620,N_14821);
and U18479 (N_18479,N_10657,N_11381);
nor U18480 (N_18480,N_10464,N_10369);
or U18481 (N_18481,N_11843,N_10377);
and U18482 (N_18482,N_12041,N_14169);
and U18483 (N_18483,N_10642,N_11497);
xnor U18484 (N_18484,N_11978,N_10385);
or U18485 (N_18485,N_12111,N_13964);
nand U18486 (N_18486,N_11291,N_13390);
nand U18487 (N_18487,N_11487,N_10827);
and U18488 (N_18488,N_11207,N_12301);
and U18489 (N_18489,N_14278,N_13978);
nor U18490 (N_18490,N_12201,N_11935);
and U18491 (N_18491,N_13051,N_13481);
xnor U18492 (N_18492,N_10373,N_10537);
or U18493 (N_18493,N_11613,N_13264);
nand U18494 (N_18494,N_13408,N_13130);
nand U18495 (N_18495,N_10965,N_14813);
or U18496 (N_18496,N_10855,N_13525);
and U18497 (N_18497,N_11095,N_12398);
and U18498 (N_18498,N_11378,N_10645);
or U18499 (N_18499,N_14852,N_10610);
nand U18500 (N_18500,N_13865,N_12223);
nor U18501 (N_18501,N_14953,N_12985);
nor U18502 (N_18502,N_12283,N_10675);
or U18503 (N_18503,N_10825,N_12582);
and U18504 (N_18504,N_11658,N_11970);
nor U18505 (N_18505,N_10180,N_13534);
nand U18506 (N_18506,N_10375,N_13934);
nor U18507 (N_18507,N_14731,N_11727);
xnor U18508 (N_18508,N_10288,N_12991);
or U18509 (N_18509,N_13068,N_13017);
nor U18510 (N_18510,N_14056,N_11872);
and U18511 (N_18511,N_12445,N_11312);
xnor U18512 (N_18512,N_13186,N_14557);
nor U18513 (N_18513,N_10971,N_12917);
nor U18514 (N_18514,N_14175,N_13556);
and U18515 (N_18515,N_12388,N_13496);
and U18516 (N_18516,N_13321,N_12168);
or U18517 (N_18517,N_12893,N_14183);
nand U18518 (N_18518,N_10446,N_14413);
nor U18519 (N_18519,N_10474,N_10230);
and U18520 (N_18520,N_14979,N_11204);
or U18521 (N_18521,N_10233,N_11310);
xnor U18522 (N_18522,N_13044,N_13195);
nand U18523 (N_18523,N_14012,N_12575);
nand U18524 (N_18524,N_13886,N_13068);
nand U18525 (N_18525,N_13830,N_12608);
nand U18526 (N_18526,N_14531,N_11614);
nor U18527 (N_18527,N_10703,N_13221);
nor U18528 (N_18528,N_14602,N_10209);
or U18529 (N_18529,N_12080,N_10154);
and U18530 (N_18530,N_12177,N_14211);
nor U18531 (N_18531,N_13467,N_12107);
or U18532 (N_18532,N_10552,N_12666);
and U18533 (N_18533,N_10339,N_11309);
nand U18534 (N_18534,N_13278,N_13935);
nand U18535 (N_18535,N_11917,N_13789);
nor U18536 (N_18536,N_12324,N_14930);
xor U18537 (N_18537,N_14070,N_14605);
or U18538 (N_18538,N_13773,N_14746);
nand U18539 (N_18539,N_10483,N_13849);
or U18540 (N_18540,N_12506,N_12678);
nand U18541 (N_18541,N_11942,N_13549);
or U18542 (N_18542,N_13740,N_10508);
and U18543 (N_18543,N_14770,N_12989);
nor U18544 (N_18544,N_10406,N_12367);
or U18545 (N_18545,N_10519,N_12259);
nand U18546 (N_18546,N_14930,N_13036);
or U18547 (N_18547,N_13742,N_11272);
nand U18548 (N_18548,N_11501,N_10922);
nor U18549 (N_18549,N_11556,N_10782);
nand U18550 (N_18550,N_12197,N_11471);
nor U18551 (N_18551,N_14876,N_13488);
or U18552 (N_18552,N_11906,N_14851);
nor U18553 (N_18553,N_10353,N_14937);
nand U18554 (N_18554,N_14345,N_12931);
nor U18555 (N_18555,N_10197,N_10061);
nor U18556 (N_18556,N_13638,N_11245);
nand U18557 (N_18557,N_11884,N_10116);
or U18558 (N_18558,N_12492,N_13082);
and U18559 (N_18559,N_13596,N_14555);
xor U18560 (N_18560,N_14856,N_14305);
xor U18561 (N_18561,N_10592,N_11551);
and U18562 (N_18562,N_14675,N_11758);
or U18563 (N_18563,N_10531,N_14481);
and U18564 (N_18564,N_12967,N_11507);
or U18565 (N_18565,N_11313,N_10468);
and U18566 (N_18566,N_12706,N_10766);
nand U18567 (N_18567,N_11101,N_13777);
and U18568 (N_18568,N_12735,N_14951);
and U18569 (N_18569,N_12847,N_11552);
nor U18570 (N_18570,N_12679,N_13018);
xnor U18571 (N_18571,N_10864,N_14574);
xnor U18572 (N_18572,N_11431,N_14276);
and U18573 (N_18573,N_14856,N_10329);
or U18574 (N_18574,N_11390,N_12287);
nor U18575 (N_18575,N_14021,N_12905);
nor U18576 (N_18576,N_14428,N_10552);
nand U18577 (N_18577,N_10863,N_13018);
nor U18578 (N_18578,N_11428,N_12778);
or U18579 (N_18579,N_11454,N_12936);
or U18580 (N_18580,N_12699,N_13481);
or U18581 (N_18581,N_11001,N_13400);
nand U18582 (N_18582,N_14303,N_12357);
nand U18583 (N_18583,N_13668,N_13935);
and U18584 (N_18584,N_12661,N_11549);
nand U18585 (N_18585,N_13685,N_13009);
and U18586 (N_18586,N_14069,N_12447);
and U18587 (N_18587,N_10996,N_10406);
nor U18588 (N_18588,N_10371,N_14812);
nor U18589 (N_18589,N_12997,N_13091);
xor U18590 (N_18590,N_13724,N_10954);
xnor U18591 (N_18591,N_11113,N_12195);
nand U18592 (N_18592,N_11375,N_14966);
nor U18593 (N_18593,N_12113,N_10036);
xnor U18594 (N_18594,N_10111,N_10348);
and U18595 (N_18595,N_13149,N_14723);
nand U18596 (N_18596,N_14473,N_10837);
or U18597 (N_18597,N_10107,N_13855);
and U18598 (N_18598,N_10672,N_14131);
or U18599 (N_18599,N_14362,N_13298);
nor U18600 (N_18600,N_11634,N_12460);
nand U18601 (N_18601,N_14023,N_11117);
and U18602 (N_18602,N_10836,N_12913);
nor U18603 (N_18603,N_12812,N_12283);
and U18604 (N_18604,N_13045,N_10249);
nand U18605 (N_18605,N_14588,N_10382);
and U18606 (N_18606,N_11624,N_13357);
nand U18607 (N_18607,N_14305,N_11722);
xnor U18608 (N_18608,N_12137,N_10526);
nor U18609 (N_18609,N_13477,N_11642);
nand U18610 (N_18610,N_11094,N_10649);
nand U18611 (N_18611,N_14579,N_11186);
nand U18612 (N_18612,N_13564,N_13325);
nand U18613 (N_18613,N_14477,N_13226);
and U18614 (N_18614,N_10227,N_14179);
and U18615 (N_18615,N_14085,N_11822);
or U18616 (N_18616,N_12226,N_13485);
and U18617 (N_18617,N_13947,N_10126);
xor U18618 (N_18618,N_13800,N_13310);
and U18619 (N_18619,N_14241,N_14281);
nor U18620 (N_18620,N_14510,N_10425);
nor U18621 (N_18621,N_10170,N_10929);
nor U18622 (N_18622,N_13786,N_10614);
nor U18623 (N_18623,N_10190,N_12552);
xor U18624 (N_18624,N_10350,N_10978);
nor U18625 (N_18625,N_10003,N_11466);
and U18626 (N_18626,N_11190,N_12943);
nand U18627 (N_18627,N_14001,N_14695);
nand U18628 (N_18628,N_12728,N_14919);
and U18629 (N_18629,N_12596,N_14445);
nand U18630 (N_18630,N_14705,N_14513);
nand U18631 (N_18631,N_12452,N_14606);
and U18632 (N_18632,N_11148,N_10681);
nor U18633 (N_18633,N_13908,N_14298);
nand U18634 (N_18634,N_13419,N_11504);
nor U18635 (N_18635,N_10039,N_12220);
and U18636 (N_18636,N_12368,N_12990);
nor U18637 (N_18637,N_10312,N_12669);
nand U18638 (N_18638,N_14432,N_13856);
nand U18639 (N_18639,N_11040,N_10270);
and U18640 (N_18640,N_10138,N_14958);
and U18641 (N_18641,N_10955,N_10424);
nand U18642 (N_18642,N_12653,N_11795);
xor U18643 (N_18643,N_11073,N_12449);
or U18644 (N_18644,N_13249,N_13835);
xor U18645 (N_18645,N_14836,N_10473);
and U18646 (N_18646,N_14388,N_11503);
xnor U18647 (N_18647,N_11687,N_13422);
xnor U18648 (N_18648,N_12296,N_12724);
nor U18649 (N_18649,N_10045,N_10859);
nor U18650 (N_18650,N_11351,N_11740);
and U18651 (N_18651,N_14633,N_14169);
nor U18652 (N_18652,N_10432,N_14064);
nor U18653 (N_18653,N_11862,N_14205);
nand U18654 (N_18654,N_10958,N_11843);
nand U18655 (N_18655,N_11227,N_14828);
and U18656 (N_18656,N_13092,N_13268);
or U18657 (N_18657,N_12423,N_11975);
nor U18658 (N_18658,N_11102,N_14937);
nor U18659 (N_18659,N_13060,N_13807);
and U18660 (N_18660,N_13078,N_11877);
nand U18661 (N_18661,N_11227,N_13697);
nor U18662 (N_18662,N_10101,N_11197);
xor U18663 (N_18663,N_10221,N_14730);
or U18664 (N_18664,N_13263,N_14697);
and U18665 (N_18665,N_14208,N_10813);
nor U18666 (N_18666,N_11645,N_10411);
or U18667 (N_18667,N_11716,N_12692);
nand U18668 (N_18668,N_13512,N_12570);
and U18669 (N_18669,N_14377,N_11826);
nand U18670 (N_18670,N_12770,N_12801);
xor U18671 (N_18671,N_12697,N_11341);
xnor U18672 (N_18672,N_12885,N_12775);
nor U18673 (N_18673,N_10266,N_10342);
nor U18674 (N_18674,N_13654,N_14006);
or U18675 (N_18675,N_13885,N_14982);
and U18676 (N_18676,N_12684,N_13556);
or U18677 (N_18677,N_10421,N_13899);
or U18678 (N_18678,N_13480,N_10700);
or U18679 (N_18679,N_11129,N_14339);
xor U18680 (N_18680,N_14523,N_12318);
xor U18681 (N_18681,N_14639,N_14430);
or U18682 (N_18682,N_13136,N_13270);
and U18683 (N_18683,N_14836,N_14246);
nand U18684 (N_18684,N_10997,N_13781);
nand U18685 (N_18685,N_14152,N_10747);
or U18686 (N_18686,N_10753,N_13102);
or U18687 (N_18687,N_10090,N_11734);
nand U18688 (N_18688,N_12784,N_11932);
nor U18689 (N_18689,N_14767,N_14310);
or U18690 (N_18690,N_13771,N_10777);
or U18691 (N_18691,N_11818,N_12947);
nor U18692 (N_18692,N_12678,N_12981);
xnor U18693 (N_18693,N_12298,N_11517);
or U18694 (N_18694,N_12651,N_14959);
nand U18695 (N_18695,N_14214,N_14748);
nand U18696 (N_18696,N_14766,N_10548);
and U18697 (N_18697,N_13371,N_11806);
or U18698 (N_18698,N_10892,N_11401);
and U18699 (N_18699,N_13266,N_10751);
nand U18700 (N_18700,N_11693,N_13837);
nor U18701 (N_18701,N_12527,N_14924);
xor U18702 (N_18702,N_14491,N_14712);
and U18703 (N_18703,N_10144,N_13656);
and U18704 (N_18704,N_10889,N_10663);
nor U18705 (N_18705,N_11429,N_14973);
and U18706 (N_18706,N_11757,N_11066);
nand U18707 (N_18707,N_10230,N_13619);
or U18708 (N_18708,N_14325,N_14142);
xor U18709 (N_18709,N_11110,N_14597);
nor U18710 (N_18710,N_13348,N_14126);
xor U18711 (N_18711,N_14714,N_14710);
nand U18712 (N_18712,N_14649,N_12781);
nor U18713 (N_18713,N_11209,N_13617);
or U18714 (N_18714,N_14191,N_11421);
nor U18715 (N_18715,N_13546,N_11997);
or U18716 (N_18716,N_14007,N_14025);
or U18717 (N_18717,N_14019,N_14336);
or U18718 (N_18718,N_12393,N_11869);
nor U18719 (N_18719,N_11987,N_13631);
or U18720 (N_18720,N_11937,N_14750);
nor U18721 (N_18721,N_12060,N_13914);
or U18722 (N_18722,N_13849,N_10737);
or U18723 (N_18723,N_10674,N_13631);
nor U18724 (N_18724,N_10292,N_14257);
and U18725 (N_18725,N_13575,N_13506);
nand U18726 (N_18726,N_14765,N_13017);
or U18727 (N_18727,N_12724,N_14127);
nand U18728 (N_18728,N_11948,N_11267);
or U18729 (N_18729,N_12511,N_13428);
or U18730 (N_18730,N_14396,N_13361);
nand U18731 (N_18731,N_12198,N_11857);
or U18732 (N_18732,N_10213,N_11892);
or U18733 (N_18733,N_13310,N_11050);
nor U18734 (N_18734,N_13572,N_14612);
or U18735 (N_18735,N_10652,N_13954);
nand U18736 (N_18736,N_12721,N_13969);
nor U18737 (N_18737,N_13873,N_13613);
and U18738 (N_18738,N_13170,N_14201);
or U18739 (N_18739,N_11340,N_14198);
and U18740 (N_18740,N_10474,N_11276);
or U18741 (N_18741,N_11650,N_14448);
and U18742 (N_18742,N_14910,N_11797);
nand U18743 (N_18743,N_14164,N_13861);
nand U18744 (N_18744,N_12491,N_14743);
nand U18745 (N_18745,N_14729,N_11997);
nand U18746 (N_18746,N_12568,N_13758);
nand U18747 (N_18747,N_11945,N_12159);
and U18748 (N_18748,N_10700,N_11218);
nand U18749 (N_18749,N_10364,N_10821);
nand U18750 (N_18750,N_13357,N_13151);
xnor U18751 (N_18751,N_13415,N_10002);
or U18752 (N_18752,N_13932,N_11064);
nand U18753 (N_18753,N_14066,N_12934);
nor U18754 (N_18754,N_12353,N_11590);
xor U18755 (N_18755,N_12660,N_12442);
nor U18756 (N_18756,N_13717,N_11400);
and U18757 (N_18757,N_11288,N_10046);
nand U18758 (N_18758,N_12063,N_12031);
or U18759 (N_18759,N_14529,N_12869);
nor U18760 (N_18760,N_12282,N_14854);
nor U18761 (N_18761,N_11574,N_13981);
and U18762 (N_18762,N_14991,N_10424);
or U18763 (N_18763,N_13819,N_13440);
nor U18764 (N_18764,N_13979,N_14217);
and U18765 (N_18765,N_13210,N_13960);
nor U18766 (N_18766,N_10291,N_14067);
or U18767 (N_18767,N_14193,N_11697);
nand U18768 (N_18768,N_13601,N_14280);
or U18769 (N_18769,N_14841,N_14608);
nand U18770 (N_18770,N_14882,N_14185);
or U18771 (N_18771,N_10827,N_14549);
nand U18772 (N_18772,N_14610,N_11165);
or U18773 (N_18773,N_12905,N_14450);
and U18774 (N_18774,N_12124,N_13535);
nor U18775 (N_18775,N_11616,N_13818);
or U18776 (N_18776,N_13138,N_14375);
or U18777 (N_18777,N_12030,N_13921);
nor U18778 (N_18778,N_14997,N_14836);
nand U18779 (N_18779,N_11037,N_12015);
xnor U18780 (N_18780,N_12092,N_13546);
nand U18781 (N_18781,N_11550,N_12653);
or U18782 (N_18782,N_14214,N_13393);
and U18783 (N_18783,N_13640,N_13592);
nand U18784 (N_18784,N_13915,N_11303);
and U18785 (N_18785,N_11289,N_13432);
and U18786 (N_18786,N_12344,N_11984);
and U18787 (N_18787,N_11162,N_13658);
xnor U18788 (N_18788,N_10668,N_14645);
and U18789 (N_18789,N_13313,N_13996);
and U18790 (N_18790,N_13675,N_10557);
and U18791 (N_18791,N_10822,N_13700);
nand U18792 (N_18792,N_10326,N_12810);
or U18793 (N_18793,N_11755,N_12442);
and U18794 (N_18794,N_14965,N_13233);
or U18795 (N_18795,N_12073,N_10536);
nand U18796 (N_18796,N_11119,N_10770);
xnor U18797 (N_18797,N_13885,N_14033);
and U18798 (N_18798,N_10539,N_12266);
nand U18799 (N_18799,N_10592,N_10008);
and U18800 (N_18800,N_10177,N_10897);
nand U18801 (N_18801,N_10883,N_10985);
and U18802 (N_18802,N_14534,N_12486);
or U18803 (N_18803,N_11045,N_10150);
xor U18804 (N_18804,N_14360,N_13120);
nand U18805 (N_18805,N_11402,N_12794);
or U18806 (N_18806,N_10807,N_12193);
xor U18807 (N_18807,N_11384,N_11094);
xnor U18808 (N_18808,N_13246,N_14441);
xnor U18809 (N_18809,N_10334,N_13549);
nand U18810 (N_18810,N_14826,N_12978);
nor U18811 (N_18811,N_14116,N_12206);
nand U18812 (N_18812,N_12629,N_14323);
nand U18813 (N_18813,N_12430,N_12138);
or U18814 (N_18814,N_12097,N_10383);
or U18815 (N_18815,N_14717,N_14833);
nand U18816 (N_18816,N_14767,N_11234);
and U18817 (N_18817,N_12327,N_14414);
and U18818 (N_18818,N_11478,N_10993);
nor U18819 (N_18819,N_12464,N_11362);
and U18820 (N_18820,N_14341,N_10822);
nor U18821 (N_18821,N_14095,N_12230);
or U18822 (N_18822,N_13006,N_12134);
nand U18823 (N_18823,N_13314,N_11456);
nor U18824 (N_18824,N_14743,N_14872);
or U18825 (N_18825,N_11104,N_11126);
and U18826 (N_18826,N_12955,N_10937);
or U18827 (N_18827,N_12191,N_10362);
nand U18828 (N_18828,N_12337,N_10222);
xnor U18829 (N_18829,N_10360,N_14852);
xor U18830 (N_18830,N_11205,N_14594);
or U18831 (N_18831,N_10832,N_10436);
nand U18832 (N_18832,N_13173,N_13686);
nor U18833 (N_18833,N_11264,N_12145);
and U18834 (N_18834,N_12650,N_13572);
or U18835 (N_18835,N_10419,N_14602);
and U18836 (N_18836,N_13529,N_14760);
nand U18837 (N_18837,N_14272,N_13458);
xor U18838 (N_18838,N_12233,N_10749);
and U18839 (N_18839,N_11365,N_13112);
nor U18840 (N_18840,N_10703,N_11363);
and U18841 (N_18841,N_11672,N_14149);
nor U18842 (N_18842,N_11465,N_14144);
nand U18843 (N_18843,N_14237,N_10544);
nor U18844 (N_18844,N_10292,N_12376);
and U18845 (N_18845,N_12747,N_12069);
or U18846 (N_18846,N_10812,N_12963);
nor U18847 (N_18847,N_11957,N_13821);
xnor U18848 (N_18848,N_10876,N_11451);
and U18849 (N_18849,N_11615,N_14997);
or U18850 (N_18850,N_14742,N_13432);
nor U18851 (N_18851,N_14128,N_14255);
or U18852 (N_18852,N_13130,N_10144);
or U18853 (N_18853,N_12752,N_13679);
nor U18854 (N_18854,N_13606,N_11812);
and U18855 (N_18855,N_11403,N_10744);
nor U18856 (N_18856,N_11042,N_14037);
nand U18857 (N_18857,N_14918,N_11979);
nand U18858 (N_18858,N_10290,N_11188);
or U18859 (N_18859,N_13076,N_10258);
or U18860 (N_18860,N_10774,N_13582);
nand U18861 (N_18861,N_13788,N_10267);
xnor U18862 (N_18862,N_10160,N_14968);
nor U18863 (N_18863,N_10801,N_14250);
or U18864 (N_18864,N_11074,N_12701);
nand U18865 (N_18865,N_10927,N_13661);
nand U18866 (N_18866,N_11490,N_12502);
and U18867 (N_18867,N_12078,N_10199);
or U18868 (N_18868,N_13559,N_14685);
nand U18869 (N_18869,N_12485,N_13420);
nor U18870 (N_18870,N_13553,N_14824);
and U18871 (N_18871,N_13569,N_13111);
xnor U18872 (N_18872,N_11320,N_11506);
nor U18873 (N_18873,N_11872,N_10405);
nand U18874 (N_18874,N_11224,N_10796);
nand U18875 (N_18875,N_11871,N_11574);
nor U18876 (N_18876,N_12476,N_13674);
nand U18877 (N_18877,N_14666,N_11604);
xor U18878 (N_18878,N_10473,N_11118);
or U18879 (N_18879,N_12360,N_10843);
or U18880 (N_18880,N_12372,N_12360);
nand U18881 (N_18881,N_10302,N_10630);
or U18882 (N_18882,N_11653,N_14237);
nor U18883 (N_18883,N_14247,N_13708);
nor U18884 (N_18884,N_14049,N_14487);
and U18885 (N_18885,N_12335,N_10687);
nand U18886 (N_18886,N_13773,N_11751);
and U18887 (N_18887,N_14292,N_10287);
xnor U18888 (N_18888,N_12828,N_10694);
or U18889 (N_18889,N_10304,N_10749);
nor U18890 (N_18890,N_10777,N_10656);
nor U18891 (N_18891,N_13058,N_13623);
xor U18892 (N_18892,N_14907,N_14299);
xnor U18893 (N_18893,N_13880,N_14131);
nand U18894 (N_18894,N_14390,N_14743);
or U18895 (N_18895,N_14041,N_12115);
and U18896 (N_18896,N_12941,N_11540);
nand U18897 (N_18897,N_10679,N_12422);
nand U18898 (N_18898,N_10091,N_13399);
or U18899 (N_18899,N_13289,N_14123);
and U18900 (N_18900,N_11145,N_12919);
nor U18901 (N_18901,N_14353,N_14049);
nand U18902 (N_18902,N_11528,N_10129);
and U18903 (N_18903,N_14760,N_14820);
xor U18904 (N_18904,N_12359,N_13181);
and U18905 (N_18905,N_13610,N_10201);
nor U18906 (N_18906,N_10984,N_10397);
nor U18907 (N_18907,N_13143,N_11987);
nand U18908 (N_18908,N_13324,N_10211);
and U18909 (N_18909,N_12583,N_13224);
xnor U18910 (N_18910,N_12832,N_11769);
nand U18911 (N_18911,N_14925,N_11816);
nand U18912 (N_18912,N_13108,N_11690);
nor U18913 (N_18913,N_13335,N_14857);
or U18914 (N_18914,N_10326,N_11578);
or U18915 (N_18915,N_11068,N_14228);
nor U18916 (N_18916,N_10981,N_12025);
nand U18917 (N_18917,N_14217,N_11945);
nor U18918 (N_18918,N_13569,N_12906);
nor U18919 (N_18919,N_11946,N_11708);
or U18920 (N_18920,N_12701,N_12403);
nor U18921 (N_18921,N_11684,N_10550);
and U18922 (N_18922,N_11949,N_14835);
and U18923 (N_18923,N_13295,N_11790);
and U18924 (N_18924,N_10297,N_14780);
nand U18925 (N_18925,N_12919,N_12834);
nand U18926 (N_18926,N_13954,N_12085);
nor U18927 (N_18927,N_13020,N_11899);
nand U18928 (N_18928,N_11692,N_12635);
xor U18929 (N_18929,N_14909,N_10727);
nor U18930 (N_18930,N_13090,N_14014);
nor U18931 (N_18931,N_11924,N_13391);
nor U18932 (N_18932,N_13018,N_10658);
or U18933 (N_18933,N_13392,N_12993);
nand U18934 (N_18934,N_13983,N_14071);
or U18935 (N_18935,N_12431,N_12897);
and U18936 (N_18936,N_10815,N_11492);
and U18937 (N_18937,N_12187,N_11678);
nand U18938 (N_18938,N_11193,N_14360);
xor U18939 (N_18939,N_12204,N_12854);
nor U18940 (N_18940,N_13969,N_10371);
nand U18941 (N_18941,N_10398,N_12021);
nand U18942 (N_18942,N_10957,N_10379);
or U18943 (N_18943,N_12342,N_13354);
nand U18944 (N_18944,N_11740,N_12262);
or U18945 (N_18945,N_12918,N_13011);
and U18946 (N_18946,N_13719,N_13148);
nand U18947 (N_18947,N_11263,N_13342);
or U18948 (N_18948,N_10447,N_10317);
or U18949 (N_18949,N_14816,N_10129);
or U18950 (N_18950,N_10913,N_13797);
xor U18951 (N_18951,N_11643,N_10134);
and U18952 (N_18952,N_11599,N_10787);
and U18953 (N_18953,N_12104,N_13954);
xor U18954 (N_18954,N_14403,N_13095);
and U18955 (N_18955,N_11029,N_12045);
nor U18956 (N_18956,N_11981,N_12901);
or U18957 (N_18957,N_13558,N_11134);
nand U18958 (N_18958,N_13496,N_14400);
nor U18959 (N_18959,N_13818,N_14172);
nor U18960 (N_18960,N_14564,N_12971);
nand U18961 (N_18961,N_12297,N_12969);
nand U18962 (N_18962,N_13380,N_10147);
or U18963 (N_18963,N_14540,N_11662);
nor U18964 (N_18964,N_12499,N_12985);
nor U18965 (N_18965,N_14475,N_13913);
and U18966 (N_18966,N_12986,N_11642);
nor U18967 (N_18967,N_12465,N_10745);
nor U18968 (N_18968,N_10368,N_12145);
and U18969 (N_18969,N_14128,N_12942);
or U18970 (N_18970,N_11089,N_13221);
or U18971 (N_18971,N_12517,N_10121);
nor U18972 (N_18972,N_12776,N_14024);
or U18973 (N_18973,N_14892,N_14337);
and U18974 (N_18974,N_12732,N_12795);
or U18975 (N_18975,N_13387,N_14213);
and U18976 (N_18976,N_13795,N_10156);
nand U18977 (N_18977,N_14417,N_11527);
and U18978 (N_18978,N_12885,N_12935);
xor U18979 (N_18979,N_11018,N_11082);
nand U18980 (N_18980,N_13986,N_11833);
and U18981 (N_18981,N_12104,N_11330);
and U18982 (N_18982,N_12366,N_13059);
or U18983 (N_18983,N_14203,N_11399);
or U18984 (N_18984,N_10337,N_13086);
or U18985 (N_18985,N_12606,N_11113);
nand U18986 (N_18986,N_13476,N_11695);
nand U18987 (N_18987,N_12103,N_11217);
or U18988 (N_18988,N_14279,N_14216);
and U18989 (N_18989,N_10204,N_11616);
and U18990 (N_18990,N_11831,N_12670);
nor U18991 (N_18991,N_10642,N_14054);
or U18992 (N_18992,N_10301,N_14101);
and U18993 (N_18993,N_11978,N_14449);
nor U18994 (N_18994,N_14397,N_14811);
nor U18995 (N_18995,N_14648,N_14100);
and U18996 (N_18996,N_12929,N_11640);
or U18997 (N_18997,N_14705,N_10362);
xnor U18998 (N_18998,N_11382,N_13410);
and U18999 (N_18999,N_14329,N_12857);
xor U19000 (N_19000,N_14915,N_14601);
nand U19001 (N_19001,N_11933,N_12783);
or U19002 (N_19002,N_13580,N_10032);
xnor U19003 (N_19003,N_14591,N_13990);
nand U19004 (N_19004,N_13898,N_14609);
and U19005 (N_19005,N_14570,N_13821);
or U19006 (N_19006,N_13703,N_11764);
and U19007 (N_19007,N_11550,N_11878);
and U19008 (N_19008,N_10316,N_11788);
nor U19009 (N_19009,N_14946,N_14026);
nand U19010 (N_19010,N_14055,N_14358);
or U19011 (N_19011,N_14957,N_14134);
or U19012 (N_19012,N_13415,N_12958);
xnor U19013 (N_19013,N_14606,N_13875);
or U19014 (N_19014,N_10597,N_14173);
nor U19015 (N_19015,N_12727,N_13329);
or U19016 (N_19016,N_11134,N_11293);
nand U19017 (N_19017,N_10767,N_14098);
nor U19018 (N_19018,N_14231,N_12920);
nor U19019 (N_19019,N_14447,N_13782);
and U19020 (N_19020,N_10749,N_10524);
or U19021 (N_19021,N_14494,N_12357);
or U19022 (N_19022,N_13554,N_11465);
nor U19023 (N_19023,N_12110,N_12713);
nand U19024 (N_19024,N_12500,N_12754);
xor U19025 (N_19025,N_13528,N_11049);
xnor U19026 (N_19026,N_11394,N_10311);
nor U19027 (N_19027,N_13320,N_14119);
or U19028 (N_19028,N_11134,N_10680);
and U19029 (N_19029,N_11251,N_12190);
and U19030 (N_19030,N_10477,N_14924);
or U19031 (N_19031,N_10567,N_11313);
nand U19032 (N_19032,N_12454,N_13621);
and U19033 (N_19033,N_13471,N_10554);
nand U19034 (N_19034,N_10755,N_13706);
xor U19035 (N_19035,N_13003,N_14548);
or U19036 (N_19036,N_14243,N_11659);
or U19037 (N_19037,N_14657,N_13561);
and U19038 (N_19038,N_10287,N_11362);
or U19039 (N_19039,N_11857,N_11752);
nor U19040 (N_19040,N_11245,N_13645);
nand U19041 (N_19041,N_14133,N_12508);
nand U19042 (N_19042,N_10617,N_11140);
and U19043 (N_19043,N_12685,N_10168);
nand U19044 (N_19044,N_14703,N_11083);
nor U19045 (N_19045,N_10415,N_10678);
nor U19046 (N_19046,N_13717,N_10004);
or U19047 (N_19047,N_10520,N_14237);
and U19048 (N_19048,N_10683,N_13397);
and U19049 (N_19049,N_10279,N_14686);
or U19050 (N_19050,N_10598,N_10839);
or U19051 (N_19051,N_14864,N_11632);
nor U19052 (N_19052,N_13229,N_13268);
nand U19053 (N_19053,N_11811,N_10892);
nor U19054 (N_19054,N_10522,N_13789);
nand U19055 (N_19055,N_14239,N_10705);
nor U19056 (N_19056,N_10322,N_14820);
or U19057 (N_19057,N_11564,N_10434);
and U19058 (N_19058,N_10973,N_12942);
or U19059 (N_19059,N_13995,N_14340);
and U19060 (N_19060,N_14020,N_13604);
and U19061 (N_19061,N_11747,N_10183);
nor U19062 (N_19062,N_12858,N_14916);
xnor U19063 (N_19063,N_11943,N_14437);
xnor U19064 (N_19064,N_12421,N_13801);
nor U19065 (N_19065,N_13811,N_11700);
nor U19066 (N_19066,N_10710,N_13723);
nor U19067 (N_19067,N_13790,N_14692);
and U19068 (N_19068,N_14433,N_13354);
nand U19069 (N_19069,N_10034,N_10294);
nor U19070 (N_19070,N_12681,N_11380);
nand U19071 (N_19071,N_11158,N_10910);
nand U19072 (N_19072,N_13052,N_10974);
xor U19073 (N_19073,N_14271,N_14632);
nand U19074 (N_19074,N_10751,N_10713);
nand U19075 (N_19075,N_13557,N_10981);
nand U19076 (N_19076,N_12805,N_11930);
nor U19077 (N_19077,N_11860,N_14312);
nor U19078 (N_19078,N_10650,N_11302);
nor U19079 (N_19079,N_12272,N_14560);
nor U19080 (N_19080,N_11603,N_10446);
or U19081 (N_19081,N_13761,N_12663);
nor U19082 (N_19082,N_10650,N_10830);
nor U19083 (N_19083,N_10874,N_12131);
or U19084 (N_19084,N_10507,N_10514);
and U19085 (N_19085,N_12809,N_13380);
or U19086 (N_19086,N_11995,N_13681);
or U19087 (N_19087,N_12438,N_10892);
xor U19088 (N_19088,N_14772,N_13253);
nor U19089 (N_19089,N_11559,N_13527);
and U19090 (N_19090,N_11274,N_10161);
or U19091 (N_19091,N_11189,N_12860);
nand U19092 (N_19092,N_12129,N_11387);
or U19093 (N_19093,N_11045,N_13865);
and U19094 (N_19094,N_14328,N_10458);
nand U19095 (N_19095,N_11792,N_12129);
xnor U19096 (N_19096,N_10972,N_11470);
or U19097 (N_19097,N_12671,N_11906);
nor U19098 (N_19098,N_13671,N_12494);
nand U19099 (N_19099,N_13914,N_13641);
or U19100 (N_19100,N_14563,N_10971);
nor U19101 (N_19101,N_11033,N_14219);
nand U19102 (N_19102,N_10981,N_10395);
nand U19103 (N_19103,N_10090,N_13419);
nor U19104 (N_19104,N_14928,N_10032);
or U19105 (N_19105,N_12904,N_13010);
and U19106 (N_19106,N_13533,N_11310);
nand U19107 (N_19107,N_13292,N_12397);
or U19108 (N_19108,N_13056,N_13806);
or U19109 (N_19109,N_10525,N_13949);
or U19110 (N_19110,N_10155,N_13848);
nand U19111 (N_19111,N_10683,N_11904);
or U19112 (N_19112,N_13580,N_11273);
and U19113 (N_19113,N_11619,N_13834);
or U19114 (N_19114,N_12058,N_10862);
or U19115 (N_19115,N_13863,N_11085);
nor U19116 (N_19116,N_12982,N_10139);
nor U19117 (N_19117,N_13634,N_14063);
nand U19118 (N_19118,N_14347,N_13249);
or U19119 (N_19119,N_10944,N_10318);
or U19120 (N_19120,N_10806,N_12371);
and U19121 (N_19121,N_13094,N_13550);
nand U19122 (N_19122,N_10149,N_11330);
nand U19123 (N_19123,N_13442,N_12647);
or U19124 (N_19124,N_13737,N_12077);
and U19125 (N_19125,N_11496,N_10276);
nor U19126 (N_19126,N_14376,N_14287);
xor U19127 (N_19127,N_10361,N_10953);
nor U19128 (N_19128,N_13283,N_10617);
and U19129 (N_19129,N_12996,N_10029);
nand U19130 (N_19130,N_13137,N_12982);
or U19131 (N_19131,N_12249,N_14132);
and U19132 (N_19132,N_11320,N_14036);
nand U19133 (N_19133,N_11187,N_13861);
xnor U19134 (N_19134,N_13326,N_14492);
or U19135 (N_19135,N_11078,N_14515);
xnor U19136 (N_19136,N_14168,N_14721);
nand U19137 (N_19137,N_12450,N_12385);
and U19138 (N_19138,N_14288,N_13248);
or U19139 (N_19139,N_11844,N_11956);
and U19140 (N_19140,N_13843,N_12798);
or U19141 (N_19141,N_11312,N_13131);
or U19142 (N_19142,N_10959,N_13578);
xnor U19143 (N_19143,N_11898,N_14476);
and U19144 (N_19144,N_10243,N_11892);
or U19145 (N_19145,N_10857,N_11974);
or U19146 (N_19146,N_13523,N_13078);
and U19147 (N_19147,N_11236,N_11797);
xnor U19148 (N_19148,N_11518,N_12516);
nor U19149 (N_19149,N_11536,N_10787);
and U19150 (N_19150,N_10822,N_12856);
nand U19151 (N_19151,N_10700,N_13691);
nor U19152 (N_19152,N_12419,N_10140);
nand U19153 (N_19153,N_12996,N_10884);
nor U19154 (N_19154,N_10375,N_13137);
or U19155 (N_19155,N_14112,N_14525);
and U19156 (N_19156,N_11066,N_11081);
and U19157 (N_19157,N_13803,N_14639);
nand U19158 (N_19158,N_12938,N_14120);
nand U19159 (N_19159,N_13683,N_14438);
nor U19160 (N_19160,N_11499,N_11265);
nand U19161 (N_19161,N_12121,N_10189);
and U19162 (N_19162,N_13366,N_10526);
xnor U19163 (N_19163,N_14070,N_11638);
nand U19164 (N_19164,N_11798,N_13240);
nor U19165 (N_19165,N_11025,N_13166);
nor U19166 (N_19166,N_11676,N_12910);
or U19167 (N_19167,N_13326,N_13116);
nor U19168 (N_19168,N_11720,N_12730);
xor U19169 (N_19169,N_11159,N_14737);
or U19170 (N_19170,N_13823,N_14747);
nand U19171 (N_19171,N_13537,N_12691);
and U19172 (N_19172,N_13650,N_10146);
xnor U19173 (N_19173,N_11905,N_11287);
nor U19174 (N_19174,N_11217,N_11799);
or U19175 (N_19175,N_13086,N_14281);
nor U19176 (N_19176,N_14148,N_10266);
nand U19177 (N_19177,N_10539,N_13567);
nor U19178 (N_19178,N_11021,N_13323);
and U19179 (N_19179,N_13328,N_11538);
and U19180 (N_19180,N_13285,N_14946);
nor U19181 (N_19181,N_13914,N_14145);
or U19182 (N_19182,N_10584,N_11654);
and U19183 (N_19183,N_14190,N_14737);
xnor U19184 (N_19184,N_14082,N_14660);
xor U19185 (N_19185,N_14961,N_12833);
nand U19186 (N_19186,N_11915,N_14519);
or U19187 (N_19187,N_11585,N_12453);
xnor U19188 (N_19188,N_11815,N_10707);
and U19189 (N_19189,N_13260,N_14120);
and U19190 (N_19190,N_10105,N_12980);
and U19191 (N_19191,N_13958,N_12652);
or U19192 (N_19192,N_14681,N_11078);
nor U19193 (N_19193,N_13972,N_14135);
and U19194 (N_19194,N_11884,N_13229);
or U19195 (N_19195,N_10908,N_12152);
or U19196 (N_19196,N_10260,N_12032);
or U19197 (N_19197,N_14805,N_11089);
or U19198 (N_19198,N_10313,N_10494);
and U19199 (N_19199,N_11973,N_10312);
nor U19200 (N_19200,N_11459,N_11181);
or U19201 (N_19201,N_13149,N_14381);
and U19202 (N_19202,N_13259,N_11385);
or U19203 (N_19203,N_13006,N_10222);
nor U19204 (N_19204,N_13745,N_13165);
and U19205 (N_19205,N_10676,N_11244);
or U19206 (N_19206,N_11177,N_11878);
nor U19207 (N_19207,N_12265,N_11831);
nor U19208 (N_19208,N_14580,N_11065);
and U19209 (N_19209,N_13486,N_10654);
and U19210 (N_19210,N_13332,N_14446);
xor U19211 (N_19211,N_11163,N_10397);
nor U19212 (N_19212,N_12287,N_13544);
nor U19213 (N_19213,N_11333,N_13362);
nand U19214 (N_19214,N_13219,N_10501);
and U19215 (N_19215,N_13036,N_10227);
nor U19216 (N_19216,N_10507,N_12362);
nor U19217 (N_19217,N_12787,N_13355);
and U19218 (N_19218,N_12040,N_12140);
nor U19219 (N_19219,N_14542,N_12053);
and U19220 (N_19220,N_14716,N_11519);
or U19221 (N_19221,N_10887,N_11978);
or U19222 (N_19222,N_14375,N_10924);
nor U19223 (N_19223,N_14852,N_11155);
or U19224 (N_19224,N_14521,N_13063);
nor U19225 (N_19225,N_14260,N_13371);
nor U19226 (N_19226,N_13102,N_10699);
nor U19227 (N_19227,N_14265,N_11175);
or U19228 (N_19228,N_12098,N_10513);
nand U19229 (N_19229,N_12026,N_12967);
nor U19230 (N_19230,N_12571,N_12582);
and U19231 (N_19231,N_13324,N_14397);
and U19232 (N_19232,N_13324,N_12928);
and U19233 (N_19233,N_10417,N_12296);
xor U19234 (N_19234,N_14385,N_11083);
and U19235 (N_19235,N_12612,N_14168);
nor U19236 (N_19236,N_12069,N_12990);
nor U19237 (N_19237,N_14868,N_13891);
or U19238 (N_19238,N_13429,N_14531);
and U19239 (N_19239,N_13199,N_10739);
nand U19240 (N_19240,N_12016,N_10495);
or U19241 (N_19241,N_10759,N_12669);
or U19242 (N_19242,N_12494,N_10192);
or U19243 (N_19243,N_11259,N_13142);
nor U19244 (N_19244,N_11524,N_12539);
nand U19245 (N_19245,N_11402,N_10687);
nand U19246 (N_19246,N_10870,N_11186);
nor U19247 (N_19247,N_12282,N_12404);
nand U19248 (N_19248,N_14387,N_13668);
nand U19249 (N_19249,N_11017,N_12681);
or U19250 (N_19250,N_10576,N_11947);
or U19251 (N_19251,N_13518,N_13242);
nor U19252 (N_19252,N_11054,N_10321);
and U19253 (N_19253,N_10984,N_13086);
nor U19254 (N_19254,N_10050,N_13294);
nor U19255 (N_19255,N_11151,N_10929);
nand U19256 (N_19256,N_10068,N_14672);
and U19257 (N_19257,N_12788,N_13464);
nor U19258 (N_19258,N_10636,N_12098);
nand U19259 (N_19259,N_13872,N_14863);
nor U19260 (N_19260,N_11521,N_14201);
nand U19261 (N_19261,N_11344,N_12023);
xor U19262 (N_19262,N_13045,N_12898);
nor U19263 (N_19263,N_12402,N_10573);
or U19264 (N_19264,N_13423,N_10938);
nor U19265 (N_19265,N_12226,N_11328);
or U19266 (N_19266,N_12964,N_11966);
nand U19267 (N_19267,N_11602,N_14548);
and U19268 (N_19268,N_14030,N_14139);
nand U19269 (N_19269,N_12455,N_12284);
or U19270 (N_19270,N_14567,N_10688);
nor U19271 (N_19271,N_13214,N_11655);
or U19272 (N_19272,N_10510,N_10508);
nor U19273 (N_19273,N_11571,N_10361);
and U19274 (N_19274,N_10205,N_14006);
and U19275 (N_19275,N_13654,N_11687);
and U19276 (N_19276,N_12435,N_11792);
and U19277 (N_19277,N_11052,N_11232);
or U19278 (N_19278,N_14261,N_14561);
nor U19279 (N_19279,N_13650,N_11256);
nor U19280 (N_19280,N_12186,N_14968);
or U19281 (N_19281,N_11527,N_10921);
nor U19282 (N_19282,N_10049,N_14389);
and U19283 (N_19283,N_14100,N_13494);
nor U19284 (N_19284,N_12417,N_10598);
or U19285 (N_19285,N_12794,N_11005);
or U19286 (N_19286,N_11995,N_13900);
xnor U19287 (N_19287,N_14692,N_14448);
and U19288 (N_19288,N_11218,N_13305);
xnor U19289 (N_19289,N_10250,N_11776);
nand U19290 (N_19290,N_11846,N_14629);
and U19291 (N_19291,N_14948,N_10604);
or U19292 (N_19292,N_11536,N_11641);
nor U19293 (N_19293,N_11751,N_11624);
nor U19294 (N_19294,N_13346,N_13222);
nor U19295 (N_19295,N_12749,N_14798);
and U19296 (N_19296,N_11411,N_11030);
and U19297 (N_19297,N_14737,N_11271);
or U19298 (N_19298,N_14657,N_14271);
nor U19299 (N_19299,N_12056,N_13219);
nand U19300 (N_19300,N_11539,N_10091);
nand U19301 (N_19301,N_11417,N_11381);
or U19302 (N_19302,N_10908,N_10901);
nor U19303 (N_19303,N_12523,N_11232);
nand U19304 (N_19304,N_12642,N_14121);
or U19305 (N_19305,N_13970,N_12660);
and U19306 (N_19306,N_11326,N_12038);
and U19307 (N_19307,N_14735,N_11792);
or U19308 (N_19308,N_12936,N_10163);
or U19309 (N_19309,N_13445,N_13732);
and U19310 (N_19310,N_14038,N_11427);
or U19311 (N_19311,N_11900,N_12757);
or U19312 (N_19312,N_14142,N_14809);
and U19313 (N_19313,N_14080,N_14750);
xnor U19314 (N_19314,N_10352,N_14770);
nand U19315 (N_19315,N_11672,N_12367);
or U19316 (N_19316,N_12262,N_11030);
nand U19317 (N_19317,N_10252,N_12187);
or U19318 (N_19318,N_10613,N_12637);
nand U19319 (N_19319,N_14570,N_13773);
and U19320 (N_19320,N_14079,N_14187);
nand U19321 (N_19321,N_14285,N_13669);
or U19322 (N_19322,N_12871,N_12220);
or U19323 (N_19323,N_14603,N_14399);
or U19324 (N_19324,N_13294,N_10984);
or U19325 (N_19325,N_13890,N_11241);
xor U19326 (N_19326,N_11505,N_10434);
or U19327 (N_19327,N_14864,N_10526);
and U19328 (N_19328,N_14816,N_11165);
nor U19329 (N_19329,N_12175,N_13777);
nand U19330 (N_19330,N_13922,N_14486);
nand U19331 (N_19331,N_11446,N_10450);
nand U19332 (N_19332,N_12113,N_14157);
and U19333 (N_19333,N_12406,N_10292);
or U19334 (N_19334,N_13105,N_14091);
or U19335 (N_19335,N_12812,N_12711);
nand U19336 (N_19336,N_14704,N_11341);
and U19337 (N_19337,N_13201,N_11997);
nand U19338 (N_19338,N_13862,N_11510);
nor U19339 (N_19339,N_10558,N_12373);
or U19340 (N_19340,N_10952,N_12965);
nand U19341 (N_19341,N_11278,N_10510);
nand U19342 (N_19342,N_12801,N_14615);
nor U19343 (N_19343,N_10040,N_11964);
nand U19344 (N_19344,N_10922,N_12648);
xor U19345 (N_19345,N_13055,N_10363);
and U19346 (N_19346,N_14554,N_13328);
or U19347 (N_19347,N_14459,N_10655);
or U19348 (N_19348,N_10340,N_14531);
and U19349 (N_19349,N_14251,N_14584);
nand U19350 (N_19350,N_14100,N_11069);
nor U19351 (N_19351,N_13190,N_12998);
nand U19352 (N_19352,N_11927,N_13932);
or U19353 (N_19353,N_11000,N_14365);
or U19354 (N_19354,N_12230,N_11977);
or U19355 (N_19355,N_11202,N_12696);
xor U19356 (N_19356,N_10491,N_13244);
xnor U19357 (N_19357,N_11790,N_10748);
nand U19358 (N_19358,N_12093,N_11538);
or U19359 (N_19359,N_14922,N_10962);
nand U19360 (N_19360,N_10717,N_10923);
nand U19361 (N_19361,N_12679,N_14532);
xor U19362 (N_19362,N_12757,N_13836);
and U19363 (N_19363,N_12547,N_10359);
nand U19364 (N_19364,N_13009,N_13707);
xnor U19365 (N_19365,N_13141,N_12824);
and U19366 (N_19366,N_14537,N_14695);
nor U19367 (N_19367,N_11070,N_13183);
or U19368 (N_19368,N_12280,N_14040);
or U19369 (N_19369,N_10024,N_13423);
and U19370 (N_19370,N_13722,N_13517);
and U19371 (N_19371,N_14769,N_12693);
and U19372 (N_19372,N_11941,N_14204);
nor U19373 (N_19373,N_11112,N_12206);
nor U19374 (N_19374,N_12863,N_10863);
or U19375 (N_19375,N_12535,N_11147);
nand U19376 (N_19376,N_10943,N_12121);
nor U19377 (N_19377,N_12111,N_10693);
or U19378 (N_19378,N_10102,N_14169);
nand U19379 (N_19379,N_10695,N_11086);
nand U19380 (N_19380,N_13827,N_13757);
nor U19381 (N_19381,N_11316,N_10947);
nand U19382 (N_19382,N_10752,N_13308);
and U19383 (N_19383,N_12381,N_10887);
or U19384 (N_19384,N_11424,N_13486);
nand U19385 (N_19385,N_14606,N_13932);
and U19386 (N_19386,N_12692,N_13779);
or U19387 (N_19387,N_11974,N_12050);
nand U19388 (N_19388,N_14270,N_10769);
nand U19389 (N_19389,N_10819,N_14553);
nor U19390 (N_19390,N_13068,N_12659);
or U19391 (N_19391,N_13889,N_12122);
nand U19392 (N_19392,N_14856,N_12504);
nor U19393 (N_19393,N_10620,N_11409);
and U19394 (N_19394,N_13422,N_14315);
and U19395 (N_19395,N_11152,N_13226);
nand U19396 (N_19396,N_14906,N_13098);
and U19397 (N_19397,N_10579,N_14432);
and U19398 (N_19398,N_10000,N_13521);
xnor U19399 (N_19399,N_12268,N_11289);
xnor U19400 (N_19400,N_11683,N_14022);
or U19401 (N_19401,N_12011,N_11021);
nor U19402 (N_19402,N_13678,N_14881);
or U19403 (N_19403,N_13397,N_13637);
and U19404 (N_19404,N_11710,N_14446);
nand U19405 (N_19405,N_11675,N_14927);
and U19406 (N_19406,N_13232,N_14368);
nand U19407 (N_19407,N_13845,N_13891);
nand U19408 (N_19408,N_11413,N_13360);
or U19409 (N_19409,N_12142,N_11182);
or U19410 (N_19410,N_14880,N_13271);
xor U19411 (N_19411,N_11358,N_13662);
nand U19412 (N_19412,N_14610,N_11620);
or U19413 (N_19413,N_12240,N_10920);
nor U19414 (N_19414,N_11407,N_13557);
or U19415 (N_19415,N_10512,N_12108);
nor U19416 (N_19416,N_13663,N_11218);
or U19417 (N_19417,N_10701,N_12897);
and U19418 (N_19418,N_11267,N_12640);
nor U19419 (N_19419,N_13776,N_12152);
nand U19420 (N_19420,N_12667,N_12134);
or U19421 (N_19421,N_10889,N_10483);
nand U19422 (N_19422,N_12549,N_10837);
xor U19423 (N_19423,N_14481,N_14692);
nor U19424 (N_19424,N_14005,N_11972);
nand U19425 (N_19425,N_11578,N_13436);
nor U19426 (N_19426,N_13979,N_12917);
xnor U19427 (N_19427,N_12489,N_11256);
nor U19428 (N_19428,N_14240,N_10658);
or U19429 (N_19429,N_12389,N_14738);
and U19430 (N_19430,N_14433,N_12047);
and U19431 (N_19431,N_11112,N_10383);
xor U19432 (N_19432,N_10332,N_13117);
and U19433 (N_19433,N_10160,N_10866);
nand U19434 (N_19434,N_10197,N_14698);
and U19435 (N_19435,N_13886,N_11106);
xnor U19436 (N_19436,N_12401,N_13033);
nor U19437 (N_19437,N_12230,N_12434);
or U19438 (N_19438,N_12941,N_13606);
nand U19439 (N_19439,N_13715,N_10566);
nand U19440 (N_19440,N_14759,N_10472);
nand U19441 (N_19441,N_10934,N_11173);
and U19442 (N_19442,N_13596,N_10154);
nor U19443 (N_19443,N_14652,N_10997);
xor U19444 (N_19444,N_10396,N_10029);
nand U19445 (N_19445,N_11245,N_12751);
xnor U19446 (N_19446,N_11830,N_14331);
xnor U19447 (N_19447,N_10234,N_10920);
or U19448 (N_19448,N_13240,N_10763);
nand U19449 (N_19449,N_11039,N_11142);
and U19450 (N_19450,N_13632,N_13697);
and U19451 (N_19451,N_14958,N_11742);
or U19452 (N_19452,N_14506,N_12079);
xor U19453 (N_19453,N_14943,N_14026);
and U19454 (N_19454,N_11874,N_11224);
or U19455 (N_19455,N_14840,N_11931);
nor U19456 (N_19456,N_14091,N_12211);
and U19457 (N_19457,N_11975,N_11331);
and U19458 (N_19458,N_11158,N_11009);
or U19459 (N_19459,N_12262,N_10319);
or U19460 (N_19460,N_14142,N_11728);
and U19461 (N_19461,N_13778,N_11921);
or U19462 (N_19462,N_14043,N_13804);
or U19463 (N_19463,N_12242,N_12120);
nor U19464 (N_19464,N_12656,N_13822);
and U19465 (N_19465,N_10747,N_14577);
nand U19466 (N_19466,N_14877,N_10838);
xnor U19467 (N_19467,N_14001,N_10942);
and U19468 (N_19468,N_14656,N_14865);
nand U19469 (N_19469,N_13302,N_14587);
nor U19470 (N_19470,N_14055,N_10317);
xnor U19471 (N_19471,N_14840,N_13592);
or U19472 (N_19472,N_11019,N_14392);
nand U19473 (N_19473,N_10199,N_10170);
nand U19474 (N_19474,N_14808,N_11937);
nand U19475 (N_19475,N_12927,N_14656);
nor U19476 (N_19476,N_12093,N_10772);
or U19477 (N_19477,N_11904,N_12850);
and U19478 (N_19478,N_14333,N_11622);
and U19479 (N_19479,N_14504,N_14302);
or U19480 (N_19480,N_14005,N_14196);
or U19481 (N_19481,N_11458,N_13768);
xor U19482 (N_19482,N_10726,N_11196);
nor U19483 (N_19483,N_12053,N_10552);
or U19484 (N_19484,N_12917,N_12497);
nor U19485 (N_19485,N_14678,N_12783);
nand U19486 (N_19486,N_13009,N_11095);
nand U19487 (N_19487,N_14110,N_10993);
nor U19488 (N_19488,N_13506,N_10041);
nor U19489 (N_19489,N_14801,N_14703);
and U19490 (N_19490,N_11396,N_10111);
nand U19491 (N_19491,N_14872,N_10447);
xor U19492 (N_19492,N_11585,N_13204);
and U19493 (N_19493,N_12793,N_11751);
nor U19494 (N_19494,N_10044,N_10186);
nor U19495 (N_19495,N_12824,N_13641);
and U19496 (N_19496,N_13096,N_11128);
and U19497 (N_19497,N_14163,N_12282);
or U19498 (N_19498,N_13629,N_10281);
xor U19499 (N_19499,N_13444,N_11589);
and U19500 (N_19500,N_14152,N_10095);
xnor U19501 (N_19501,N_11141,N_11055);
nand U19502 (N_19502,N_12499,N_10760);
xnor U19503 (N_19503,N_13512,N_10290);
or U19504 (N_19504,N_13884,N_12674);
or U19505 (N_19505,N_13491,N_13152);
nor U19506 (N_19506,N_13484,N_10858);
nand U19507 (N_19507,N_13169,N_14783);
and U19508 (N_19508,N_14934,N_12508);
or U19509 (N_19509,N_12732,N_12208);
nor U19510 (N_19510,N_10256,N_12579);
or U19511 (N_19511,N_11279,N_13031);
nand U19512 (N_19512,N_13701,N_14934);
xnor U19513 (N_19513,N_11715,N_13735);
nand U19514 (N_19514,N_12155,N_10758);
or U19515 (N_19515,N_12555,N_10321);
xor U19516 (N_19516,N_10713,N_12242);
nor U19517 (N_19517,N_13065,N_12496);
nand U19518 (N_19518,N_13787,N_13101);
xnor U19519 (N_19519,N_12158,N_12173);
or U19520 (N_19520,N_11384,N_12201);
and U19521 (N_19521,N_13358,N_14928);
or U19522 (N_19522,N_10386,N_13137);
or U19523 (N_19523,N_12739,N_12477);
or U19524 (N_19524,N_13413,N_12490);
or U19525 (N_19525,N_13801,N_10797);
nor U19526 (N_19526,N_12754,N_11339);
nand U19527 (N_19527,N_12911,N_10107);
nand U19528 (N_19528,N_14677,N_12835);
nor U19529 (N_19529,N_11076,N_10282);
nor U19530 (N_19530,N_11783,N_11059);
xnor U19531 (N_19531,N_13048,N_11911);
and U19532 (N_19532,N_14040,N_14139);
or U19533 (N_19533,N_10159,N_13444);
nor U19534 (N_19534,N_13372,N_12952);
nor U19535 (N_19535,N_14180,N_11290);
or U19536 (N_19536,N_11879,N_11915);
nor U19537 (N_19537,N_12951,N_12753);
or U19538 (N_19538,N_11187,N_10787);
or U19539 (N_19539,N_12194,N_11613);
nand U19540 (N_19540,N_12024,N_10935);
or U19541 (N_19541,N_10637,N_11175);
nand U19542 (N_19542,N_13943,N_14231);
or U19543 (N_19543,N_13349,N_13119);
nand U19544 (N_19544,N_12251,N_14375);
xor U19545 (N_19545,N_12891,N_12136);
nor U19546 (N_19546,N_10502,N_13424);
nor U19547 (N_19547,N_10691,N_10755);
or U19548 (N_19548,N_11783,N_14758);
and U19549 (N_19549,N_13972,N_14387);
and U19550 (N_19550,N_14956,N_10945);
and U19551 (N_19551,N_10294,N_13325);
xnor U19552 (N_19552,N_14396,N_14170);
and U19553 (N_19553,N_13894,N_14556);
nor U19554 (N_19554,N_11089,N_10681);
or U19555 (N_19555,N_11512,N_12823);
and U19556 (N_19556,N_11761,N_13228);
xnor U19557 (N_19557,N_12861,N_11198);
nor U19558 (N_19558,N_12892,N_11505);
xor U19559 (N_19559,N_10999,N_11302);
nand U19560 (N_19560,N_11258,N_14538);
or U19561 (N_19561,N_12679,N_12100);
and U19562 (N_19562,N_13276,N_10342);
nor U19563 (N_19563,N_12387,N_10450);
or U19564 (N_19564,N_11432,N_10948);
nand U19565 (N_19565,N_10902,N_11284);
nand U19566 (N_19566,N_10906,N_11699);
nor U19567 (N_19567,N_13063,N_13707);
or U19568 (N_19568,N_11027,N_10678);
nor U19569 (N_19569,N_10543,N_12115);
and U19570 (N_19570,N_11502,N_12167);
nor U19571 (N_19571,N_12999,N_11770);
and U19572 (N_19572,N_13187,N_12708);
and U19573 (N_19573,N_12713,N_10901);
or U19574 (N_19574,N_10766,N_13523);
or U19575 (N_19575,N_14665,N_10235);
nand U19576 (N_19576,N_13960,N_14643);
nor U19577 (N_19577,N_11632,N_14568);
and U19578 (N_19578,N_14512,N_14005);
nor U19579 (N_19579,N_12921,N_11322);
nor U19580 (N_19580,N_12669,N_12531);
nand U19581 (N_19581,N_10978,N_14149);
or U19582 (N_19582,N_10665,N_10554);
and U19583 (N_19583,N_14597,N_12668);
nor U19584 (N_19584,N_13171,N_12041);
xnor U19585 (N_19585,N_10937,N_11715);
xnor U19586 (N_19586,N_12558,N_10423);
and U19587 (N_19587,N_12856,N_13151);
and U19588 (N_19588,N_13197,N_11863);
or U19589 (N_19589,N_10292,N_11319);
nor U19590 (N_19590,N_11207,N_14249);
and U19591 (N_19591,N_14800,N_12958);
or U19592 (N_19592,N_11467,N_11566);
and U19593 (N_19593,N_10311,N_12128);
nand U19594 (N_19594,N_10169,N_14586);
and U19595 (N_19595,N_14196,N_10065);
nor U19596 (N_19596,N_11884,N_13684);
and U19597 (N_19597,N_10459,N_14989);
nor U19598 (N_19598,N_10241,N_12925);
and U19599 (N_19599,N_11655,N_11606);
nand U19600 (N_19600,N_12390,N_13972);
nor U19601 (N_19601,N_13188,N_13617);
or U19602 (N_19602,N_12707,N_11990);
nand U19603 (N_19603,N_13449,N_13204);
and U19604 (N_19604,N_13300,N_10787);
nand U19605 (N_19605,N_14039,N_11713);
nor U19606 (N_19606,N_10602,N_13624);
nand U19607 (N_19607,N_13194,N_13182);
and U19608 (N_19608,N_14576,N_12635);
or U19609 (N_19609,N_14734,N_13399);
or U19610 (N_19610,N_12011,N_14528);
and U19611 (N_19611,N_11137,N_11883);
and U19612 (N_19612,N_10773,N_12879);
and U19613 (N_19613,N_14904,N_14845);
xor U19614 (N_19614,N_13905,N_13923);
or U19615 (N_19615,N_10715,N_10427);
nand U19616 (N_19616,N_11786,N_13490);
or U19617 (N_19617,N_11609,N_13309);
nand U19618 (N_19618,N_11707,N_12303);
xnor U19619 (N_19619,N_14322,N_11733);
nor U19620 (N_19620,N_14867,N_11521);
nor U19621 (N_19621,N_13890,N_13689);
or U19622 (N_19622,N_10109,N_13560);
or U19623 (N_19623,N_10752,N_10667);
and U19624 (N_19624,N_10586,N_14212);
and U19625 (N_19625,N_10205,N_12164);
xor U19626 (N_19626,N_10582,N_13807);
nor U19627 (N_19627,N_13414,N_14747);
and U19628 (N_19628,N_11820,N_12083);
nand U19629 (N_19629,N_11772,N_12680);
nor U19630 (N_19630,N_11160,N_11948);
or U19631 (N_19631,N_10514,N_13401);
nor U19632 (N_19632,N_10104,N_12151);
or U19633 (N_19633,N_13944,N_12230);
nand U19634 (N_19634,N_13072,N_11386);
xnor U19635 (N_19635,N_11832,N_13138);
nor U19636 (N_19636,N_14934,N_13726);
or U19637 (N_19637,N_13736,N_12543);
nor U19638 (N_19638,N_12221,N_12294);
and U19639 (N_19639,N_12590,N_14263);
nor U19640 (N_19640,N_14427,N_14682);
nor U19641 (N_19641,N_12221,N_10655);
nand U19642 (N_19642,N_11356,N_12801);
nand U19643 (N_19643,N_11776,N_11113);
nor U19644 (N_19644,N_14179,N_12838);
xor U19645 (N_19645,N_14118,N_13050);
or U19646 (N_19646,N_10361,N_12579);
or U19647 (N_19647,N_11584,N_11327);
and U19648 (N_19648,N_13651,N_11312);
nand U19649 (N_19649,N_12922,N_12626);
nand U19650 (N_19650,N_11494,N_10862);
nor U19651 (N_19651,N_11348,N_13790);
and U19652 (N_19652,N_13128,N_14091);
nand U19653 (N_19653,N_10072,N_11960);
and U19654 (N_19654,N_12020,N_13680);
nor U19655 (N_19655,N_12182,N_13565);
nand U19656 (N_19656,N_14853,N_11665);
nand U19657 (N_19657,N_10914,N_13906);
nor U19658 (N_19658,N_12185,N_13471);
nand U19659 (N_19659,N_12318,N_13880);
or U19660 (N_19660,N_10448,N_11319);
xnor U19661 (N_19661,N_13911,N_11884);
nand U19662 (N_19662,N_13842,N_13659);
nand U19663 (N_19663,N_11611,N_14411);
nand U19664 (N_19664,N_13910,N_12395);
or U19665 (N_19665,N_11630,N_11978);
or U19666 (N_19666,N_12540,N_11005);
or U19667 (N_19667,N_12740,N_11232);
and U19668 (N_19668,N_10921,N_11261);
and U19669 (N_19669,N_11210,N_11155);
xnor U19670 (N_19670,N_11590,N_11878);
or U19671 (N_19671,N_13246,N_10816);
nand U19672 (N_19672,N_10813,N_10367);
nand U19673 (N_19673,N_12453,N_13177);
nor U19674 (N_19674,N_13886,N_11438);
and U19675 (N_19675,N_12029,N_10548);
nor U19676 (N_19676,N_13397,N_12859);
or U19677 (N_19677,N_12005,N_11361);
xnor U19678 (N_19678,N_14588,N_12137);
nand U19679 (N_19679,N_12418,N_14165);
xor U19680 (N_19680,N_13694,N_11511);
nand U19681 (N_19681,N_10024,N_12455);
or U19682 (N_19682,N_14575,N_12605);
nand U19683 (N_19683,N_11503,N_13159);
or U19684 (N_19684,N_14835,N_14506);
nor U19685 (N_19685,N_11945,N_12731);
nand U19686 (N_19686,N_11281,N_12257);
and U19687 (N_19687,N_12845,N_11484);
nor U19688 (N_19688,N_13089,N_11252);
and U19689 (N_19689,N_11509,N_14806);
and U19690 (N_19690,N_12273,N_11304);
nor U19691 (N_19691,N_11541,N_13109);
nor U19692 (N_19692,N_13661,N_11099);
nor U19693 (N_19693,N_10947,N_10420);
and U19694 (N_19694,N_13719,N_11070);
and U19695 (N_19695,N_10247,N_12764);
and U19696 (N_19696,N_11795,N_13191);
nor U19697 (N_19697,N_13895,N_13179);
or U19698 (N_19698,N_12890,N_11816);
nor U19699 (N_19699,N_13002,N_14417);
nand U19700 (N_19700,N_11045,N_14125);
xor U19701 (N_19701,N_11102,N_13994);
xnor U19702 (N_19702,N_10126,N_11122);
and U19703 (N_19703,N_13649,N_12474);
xnor U19704 (N_19704,N_11982,N_11471);
nand U19705 (N_19705,N_11571,N_10703);
nor U19706 (N_19706,N_14629,N_12149);
nand U19707 (N_19707,N_12053,N_11712);
nor U19708 (N_19708,N_12166,N_10838);
nor U19709 (N_19709,N_14439,N_12882);
or U19710 (N_19710,N_13383,N_10867);
or U19711 (N_19711,N_10856,N_10318);
nor U19712 (N_19712,N_11518,N_11867);
xor U19713 (N_19713,N_10349,N_12627);
xnor U19714 (N_19714,N_13104,N_10817);
nand U19715 (N_19715,N_10355,N_12972);
and U19716 (N_19716,N_12978,N_11051);
nor U19717 (N_19717,N_11110,N_14090);
xor U19718 (N_19718,N_11291,N_13988);
nor U19719 (N_19719,N_13040,N_14439);
nand U19720 (N_19720,N_12317,N_10241);
nand U19721 (N_19721,N_13885,N_13595);
nand U19722 (N_19722,N_11264,N_13494);
or U19723 (N_19723,N_14392,N_10071);
and U19724 (N_19724,N_13903,N_14118);
and U19725 (N_19725,N_14331,N_11253);
nor U19726 (N_19726,N_13951,N_13002);
nor U19727 (N_19727,N_14348,N_12952);
nand U19728 (N_19728,N_12336,N_10552);
or U19729 (N_19729,N_13167,N_13523);
or U19730 (N_19730,N_10860,N_12167);
xor U19731 (N_19731,N_13502,N_13831);
nor U19732 (N_19732,N_11685,N_10626);
xor U19733 (N_19733,N_10979,N_13470);
nand U19734 (N_19734,N_10488,N_12891);
or U19735 (N_19735,N_11725,N_12075);
and U19736 (N_19736,N_14610,N_10667);
xor U19737 (N_19737,N_11649,N_12747);
or U19738 (N_19738,N_12718,N_11778);
nand U19739 (N_19739,N_11737,N_14832);
and U19740 (N_19740,N_10209,N_10358);
nor U19741 (N_19741,N_14657,N_10839);
or U19742 (N_19742,N_12670,N_12822);
nor U19743 (N_19743,N_11742,N_11346);
nand U19744 (N_19744,N_12493,N_14844);
xnor U19745 (N_19745,N_13574,N_11378);
nand U19746 (N_19746,N_13316,N_12761);
or U19747 (N_19747,N_11837,N_10702);
and U19748 (N_19748,N_12592,N_11043);
and U19749 (N_19749,N_10652,N_12681);
and U19750 (N_19750,N_13728,N_12517);
and U19751 (N_19751,N_14949,N_13258);
nor U19752 (N_19752,N_14536,N_11074);
nor U19753 (N_19753,N_13517,N_10346);
nor U19754 (N_19754,N_12784,N_10363);
xor U19755 (N_19755,N_11732,N_12214);
and U19756 (N_19756,N_13256,N_11496);
nor U19757 (N_19757,N_12259,N_12749);
nor U19758 (N_19758,N_10629,N_11064);
or U19759 (N_19759,N_12511,N_11613);
nand U19760 (N_19760,N_14691,N_11587);
nand U19761 (N_19761,N_10868,N_12237);
or U19762 (N_19762,N_13402,N_11530);
or U19763 (N_19763,N_11208,N_11582);
nor U19764 (N_19764,N_13690,N_14136);
nand U19765 (N_19765,N_11011,N_11128);
or U19766 (N_19766,N_12320,N_12108);
and U19767 (N_19767,N_13485,N_10730);
nand U19768 (N_19768,N_11071,N_12209);
nand U19769 (N_19769,N_13474,N_10950);
nand U19770 (N_19770,N_14207,N_13502);
nor U19771 (N_19771,N_12330,N_12060);
or U19772 (N_19772,N_13090,N_13668);
nand U19773 (N_19773,N_13202,N_13308);
xnor U19774 (N_19774,N_10624,N_10283);
or U19775 (N_19775,N_13539,N_10527);
xor U19776 (N_19776,N_11682,N_13422);
nor U19777 (N_19777,N_11715,N_12461);
xor U19778 (N_19778,N_11721,N_12343);
or U19779 (N_19779,N_13869,N_13144);
or U19780 (N_19780,N_12172,N_12067);
or U19781 (N_19781,N_11080,N_13906);
or U19782 (N_19782,N_10963,N_12621);
and U19783 (N_19783,N_11744,N_12027);
nand U19784 (N_19784,N_12640,N_13460);
nor U19785 (N_19785,N_10851,N_12448);
nor U19786 (N_19786,N_11817,N_10936);
nor U19787 (N_19787,N_12025,N_11982);
or U19788 (N_19788,N_10029,N_14292);
and U19789 (N_19789,N_11587,N_14451);
and U19790 (N_19790,N_14506,N_14507);
nand U19791 (N_19791,N_13256,N_13813);
or U19792 (N_19792,N_11729,N_14583);
nor U19793 (N_19793,N_10175,N_10076);
nor U19794 (N_19794,N_11969,N_13717);
nand U19795 (N_19795,N_13194,N_11641);
and U19796 (N_19796,N_14292,N_13520);
nand U19797 (N_19797,N_11673,N_10800);
or U19798 (N_19798,N_13700,N_14062);
nor U19799 (N_19799,N_11350,N_10463);
or U19800 (N_19800,N_12830,N_11157);
xnor U19801 (N_19801,N_11022,N_10060);
xnor U19802 (N_19802,N_13571,N_13128);
and U19803 (N_19803,N_13558,N_11561);
nor U19804 (N_19804,N_13928,N_10435);
nand U19805 (N_19805,N_10405,N_12482);
and U19806 (N_19806,N_13906,N_11413);
or U19807 (N_19807,N_14410,N_11166);
or U19808 (N_19808,N_13428,N_10835);
nor U19809 (N_19809,N_10461,N_12463);
nor U19810 (N_19810,N_14872,N_10782);
and U19811 (N_19811,N_14330,N_13180);
nor U19812 (N_19812,N_11076,N_10233);
nor U19813 (N_19813,N_11044,N_10658);
xor U19814 (N_19814,N_12283,N_14305);
or U19815 (N_19815,N_13113,N_14515);
or U19816 (N_19816,N_11832,N_12673);
nor U19817 (N_19817,N_10530,N_13190);
and U19818 (N_19818,N_12612,N_10007);
or U19819 (N_19819,N_14245,N_14677);
or U19820 (N_19820,N_12301,N_10853);
nor U19821 (N_19821,N_14072,N_14402);
nor U19822 (N_19822,N_13945,N_14929);
or U19823 (N_19823,N_11110,N_10099);
nor U19824 (N_19824,N_12760,N_14543);
or U19825 (N_19825,N_12645,N_12879);
nor U19826 (N_19826,N_13112,N_14042);
or U19827 (N_19827,N_12664,N_10343);
and U19828 (N_19828,N_13037,N_13453);
or U19829 (N_19829,N_10132,N_13497);
and U19830 (N_19830,N_10291,N_11819);
or U19831 (N_19831,N_13336,N_12977);
or U19832 (N_19832,N_10041,N_11922);
nor U19833 (N_19833,N_11174,N_11052);
and U19834 (N_19834,N_10489,N_10663);
nor U19835 (N_19835,N_10450,N_13991);
nor U19836 (N_19836,N_12880,N_13015);
or U19837 (N_19837,N_10953,N_10074);
and U19838 (N_19838,N_14031,N_13148);
or U19839 (N_19839,N_13294,N_13941);
or U19840 (N_19840,N_11064,N_12352);
nor U19841 (N_19841,N_11827,N_10630);
or U19842 (N_19842,N_10669,N_13314);
nor U19843 (N_19843,N_11780,N_10987);
xor U19844 (N_19844,N_12772,N_12429);
nor U19845 (N_19845,N_11148,N_14897);
or U19846 (N_19846,N_14745,N_11478);
and U19847 (N_19847,N_11721,N_10841);
and U19848 (N_19848,N_12794,N_13894);
nor U19849 (N_19849,N_14728,N_13125);
xnor U19850 (N_19850,N_13433,N_10133);
and U19851 (N_19851,N_14457,N_12017);
nor U19852 (N_19852,N_10018,N_11003);
nor U19853 (N_19853,N_10953,N_13582);
xnor U19854 (N_19854,N_13108,N_10703);
nand U19855 (N_19855,N_12159,N_14568);
and U19856 (N_19856,N_10434,N_14369);
nand U19857 (N_19857,N_13271,N_11680);
nand U19858 (N_19858,N_11409,N_13908);
and U19859 (N_19859,N_12970,N_11284);
nand U19860 (N_19860,N_13706,N_12025);
nand U19861 (N_19861,N_14359,N_14291);
and U19862 (N_19862,N_12821,N_14763);
nand U19863 (N_19863,N_12123,N_13600);
xor U19864 (N_19864,N_10487,N_12218);
nor U19865 (N_19865,N_11613,N_13806);
nor U19866 (N_19866,N_11033,N_14068);
or U19867 (N_19867,N_14740,N_12755);
xor U19868 (N_19868,N_13396,N_13649);
or U19869 (N_19869,N_13292,N_13177);
nor U19870 (N_19870,N_11119,N_10479);
or U19871 (N_19871,N_10879,N_13332);
and U19872 (N_19872,N_10152,N_12996);
or U19873 (N_19873,N_11892,N_11066);
and U19874 (N_19874,N_12403,N_11337);
and U19875 (N_19875,N_12466,N_11408);
and U19876 (N_19876,N_12775,N_13629);
nor U19877 (N_19877,N_11473,N_11583);
nor U19878 (N_19878,N_11301,N_11230);
nor U19879 (N_19879,N_14775,N_14256);
and U19880 (N_19880,N_11434,N_12570);
or U19881 (N_19881,N_13795,N_10862);
nor U19882 (N_19882,N_12519,N_11235);
nand U19883 (N_19883,N_12064,N_13160);
nor U19884 (N_19884,N_13458,N_13042);
nand U19885 (N_19885,N_14960,N_14129);
nand U19886 (N_19886,N_14160,N_13125);
and U19887 (N_19887,N_10810,N_14359);
or U19888 (N_19888,N_11259,N_14236);
nand U19889 (N_19889,N_14126,N_14691);
nand U19890 (N_19890,N_13882,N_10905);
nor U19891 (N_19891,N_12695,N_14468);
nand U19892 (N_19892,N_10363,N_11958);
xor U19893 (N_19893,N_12598,N_11969);
nand U19894 (N_19894,N_14850,N_12244);
or U19895 (N_19895,N_14883,N_14967);
nor U19896 (N_19896,N_14410,N_11514);
nor U19897 (N_19897,N_12241,N_14459);
nor U19898 (N_19898,N_11571,N_14446);
xor U19899 (N_19899,N_13769,N_11574);
or U19900 (N_19900,N_14960,N_13338);
and U19901 (N_19901,N_14009,N_14064);
nor U19902 (N_19902,N_10687,N_11962);
and U19903 (N_19903,N_12666,N_10602);
and U19904 (N_19904,N_12212,N_10758);
or U19905 (N_19905,N_13867,N_11814);
xor U19906 (N_19906,N_13758,N_12975);
or U19907 (N_19907,N_11277,N_13843);
and U19908 (N_19908,N_12388,N_14453);
nand U19909 (N_19909,N_12077,N_13604);
and U19910 (N_19910,N_10212,N_14355);
or U19911 (N_19911,N_10657,N_12272);
and U19912 (N_19912,N_14230,N_13099);
nor U19913 (N_19913,N_12386,N_11850);
or U19914 (N_19914,N_13518,N_10936);
and U19915 (N_19915,N_14804,N_14901);
nand U19916 (N_19916,N_10112,N_12488);
nand U19917 (N_19917,N_13550,N_11693);
nor U19918 (N_19918,N_12548,N_10702);
nor U19919 (N_19919,N_14833,N_13579);
and U19920 (N_19920,N_13279,N_14097);
nand U19921 (N_19921,N_11266,N_12678);
nor U19922 (N_19922,N_13368,N_14345);
nand U19923 (N_19923,N_14007,N_12314);
or U19924 (N_19924,N_11146,N_10343);
nor U19925 (N_19925,N_12050,N_11295);
or U19926 (N_19926,N_13001,N_11401);
and U19927 (N_19927,N_14018,N_14841);
nor U19928 (N_19928,N_14231,N_13474);
or U19929 (N_19929,N_12244,N_13023);
nand U19930 (N_19930,N_12918,N_13664);
and U19931 (N_19931,N_13817,N_13540);
nor U19932 (N_19932,N_12000,N_14043);
or U19933 (N_19933,N_13015,N_11894);
or U19934 (N_19934,N_12763,N_14990);
and U19935 (N_19935,N_13040,N_11883);
nand U19936 (N_19936,N_13738,N_10682);
and U19937 (N_19937,N_12028,N_13636);
and U19938 (N_19938,N_13729,N_10776);
and U19939 (N_19939,N_12497,N_13220);
nor U19940 (N_19940,N_11866,N_14123);
nand U19941 (N_19941,N_12778,N_10282);
nand U19942 (N_19942,N_11983,N_11704);
nand U19943 (N_19943,N_14441,N_13050);
xor U19944 (N_19944,N_13360,N_14319);
or U19945 (N_19945,N_11621,N_11650);
and U19946 (N_19946,N_13555,N_12759);
nand U19947 (N_19947,N_13505,N_11007);
and U19948 (N_19948,N_10063,N_10352);
and U19949 (N_19949,N_10206,N_14943);
and U19950 (N_19950,N_12075,N_11944);
nand U19951 (N_19951,N_12941,N_12525);
nand U19952 (N_19952,N_14711,N_14533);
nand U19953 (N_19953,N_14310,N_10430);
nor U19954 (N_19954,N_13226,N_10042);
and U19955 (N_19955,N_12139,N_10504);
or U19956 (N_19956,N_14470,N_13854);
nand U19957 (N_19957,N_14846,N_13675);
or U19958 (N_19958,N_14050,N_13950);
xnor U19959 (N_19959,N_14580,N_12352);
nand U19960 (N_19960,N_10848,N_11386);
nand U19961 (N_19961,N_14902,N_12524);
nand U19962 (N_19962,N_13918,N_14777);
nor U19963 (N_19963,N_13586,N_14463);
nand U19964 (N_19964,N_10798,N_13682);
nand U19965 (N_19965,N_11737,N_11529);
nand U19966 (N_19966,N_11674,N_10042);
or U19967 (N_19967,N_14268,N_11338);
nand U19968 (N_19968,N_12631,N_10407);
nor U19969 (N_19969,N_13936,N_13382);
nor U19970 (N_19970,N_14893,N_14703);
or U19971 (N_19971,N_10674,N_14314);
and U19972 (N_19972,N_11228,N_10042);
nand U19973 (N_19973,N_10119,N_12506);
or U19974 (N_19974,N_11282,N_13828);
nor U19975 (N_19975,N_11579,N_13810);
or U19976 (N_19976,N_13311,N_10834);
and U19977 (N_19977,N_12097,N_11137);
or U19978 (N_19978,N_10690,N_13226);
nor U19979 (N_19979,N_11722,N_12262);
or U19980 (N_19980,N_11701,N_13591);
nand U19981 (N_19981,N_14566,N_13168);
xnor U19982 (N_19982,N_12044,N_10722);
and U19983 (N_19983,N_12381,N_14371);
nand U19984 (N_19984,N_10049,N_14915);
nor U19985 (N_19985,N_11665,N_12330);
or U19986 (N_19986,N_14731,N_13945);
nand U19987 (N_19987,N_12745,N_13791);
or U19988 (N_19988,N_12422,N_14763);
and U19989 (N_19989,N_11527,N_13575);
and U19990 (N_19990,N_11543,N_13088);
or U19991 (N_19991,N_12325,N_12688);
and U19992 (N_19992,N_10807,N_10715);
xnor U19993 (N_19993,N_12122,N_11519);
nand U19994 (N_19994,N_10510,N_13306);
nor U19995 (N_19995,N_11687,N_13845);
nor U19996 (N_19996,N_12392,N_10104);
nand U19997 (N_19997,N_12469,N_12098);
nand U19998 (N_19998,N_13523,N_14170);
xor U19999 (N_19999,N_14201,N_10690);
or UO_0 (O_0,N_15457,N_17208);
or UO_1 (O_1,N_15605,N_19142);
nor UO_2 (O_2,N_19486,N_19890);
nand UO_3 (O_3,N_17964,N_15108);
nand UO_4 (O_4,N_16275,N_19513);
xnor UO_5 (O_5,N_15553,N_16906);
nor UO_6 (O_6,N_15573,N_15741);
nand UO_7 (O_7,N_18156,N_17275);
nor UO_8 (O_8,N_18751,N_16018);
nand UO_9 (O_9,N_16369,N_19241);
nor UO_10 (O_10,N_18676,N_18986);
nor UO_11 (O_11,N_17393,N_17899);
nor UO_12 (O_12,N_19076,N_15054);
nand UO_13 (O_13,N_17390,N_18848);
or UO_14 (O_14,N_19406,N_17292);
and UO_15 (O_15,N_17141,N_18446);
nor UO_16 (O_16,N_15044,N_15890);
or UO_17 (O_17,N_18534,N_15239);
nand UO_18 (O_18,N_17860,N_15430);
nand UO_19 (O_19,N_15823,N_16184);
or UO_20 (O_20,N_17590,N_15319);
and UO_21 (O_21,N_17652,N_16991);
xor UO_22 (O_22,N_16070,N_18095);
xor UO_23 (O_23,N_18933,N_15226);
and UO_24 (O_24,N_15874,N_16979);
or UO_25 (O_25,N_18993,N_18880);
nand UO_26 (O_26,N_15110,N_17391);
nand UO_27 (O_27,N_16605,N_15956);
xnor UO_28 (O_28,N_15900,N_15832);
nor UO_29 (O_29,N_18757,N_16085);
and UO_30 (O_30,N_15973,N_18407);
and UO_31 (O_31,N_18711,N_19074);
nor UO_32 (O_32,N_19280,N_18208);
or UO_33 (O_33,N_18712,N_19430);
or UO_34 (O_34,N_19049,N_15174);
or UO_35 (O_35,N_19887,N_16058);
nor UO_36 (O_36,N_17161,N_18469);
xor UO_37 (O_37,N_15760,N_19741);
and UO_38 (O_38,N_15439,N_18530);
nor UO_39 (O_39,N_16022,N_19427);
and UO_40 (O_40,N_15467,N_18588);
nor UO_41 (O_41,N_15841,N_15342);
nand UO_42 (O_42,N_15733,N_18009);
or UO_43 (O_43,N_16782,N_17126);
nand UO_44 (O_44,N_17955,N_19946);
and UO_45 (O_45,N_15462,N_17140);
or UO_46 (O_46,N_15887,N_17113);
nor UO_47 (O_47,N_18758,N_18778);
xor UO_48 (O_48,N_17884,N_16598);
or UO_49 (O_49,N_18051,N_15525);
nand UO_50 (O_50,N_19010,N_17686);
nor UO_51 (O_51,N_15512,N_15953);
nor UO_52 (O_52,N_15100,N_15707);
nand UO_53 (O_53,N_18125,N_19967);
and UO_54 (O_54,N_19623,N_19933);
and UO_55 (O_55,N_19817,N_17895);
or UO_56 (O_56,N_19019,N_15798);
nor UO_57 (O_57,N_16017,N_16749);
and UO_58 (O_58,N_18226,N_15781);
or UO_59 (O_59,N_16786,N_16137);
or UO_60 (O_60,N_15807,N_15433);
nor UO_61 (O_61,N_19526,N_18411);
nor UO_62 (O_62,N_19233,N_18982);
and UO_63 (O_63,N_16948,N_17909);
and UO_64 (O_64,N_19336,N_17672);
nor UO_65 (O_65,N_17482,N_19458);
or UO_66 (O_66,N_16042,N_19463);
nand UO_67 (O_67,N_19337,N_18936);
nor UO_68 (O_68,N_16169,N_17935);
nor UO_69 (O_69,N_18533,N_15192);
and UO_70 (O_70,N_19878,N_16514);
and UO_71 (O_71,N_18216,N_17684);
nor UO_72 (O_72,N_18867,N_19418);
and UO_73 (O_73,N_18419,N_18200);
or UO_74 (O_74,N_17312,N_16316);
nand UO_75 (O_75,N_17748,N_18395);
nor UO_76 (O_76,N_18769,N_16958);
nor UO_77 (O_77,N_15928,N_18231);
nand UO_78 (O_78,N_16265,N_17134);
nand UO_79 (O_79,N_18700,N_18238);
and UO_80 (O_80,N_15301,N_16073);
or UO_81 (O_81,N_19966,N_15107);
xnor UO_82 (O_82,N_15762,N_15412);
and UO_83 (O_83,N_16315,N_15620);
and UO_84 (O_84,N_17417,N_17387);
and UO_85 (O_85,N_18034,N_15895);
nand UO_86 (O_86,N_19766,N_18295);
nor UO_87 (O_87,N_16756,N_19979);
nand UO_88 (O_88,N_16268,N_16325);
or UO_89 (O_89,N_16513,N_18330);
and UO_90 (O_90,N_17398,N_18389);
nor UO_91 (O_91,N_16375,N_19532);
and UO_92 (O_92,N_15509,N_15492);
nand UO_93 (O_93,N_19941,N_17222);
nand UO_94 (O_94,N_19928,N_15809);
nor UO_95 (O_95,N_15775,N_15323);
nand UO_96 (O_96,N_15254,N_18709);
nand UO_97 (O_97,N_15036,N_18786);
and UO_98 (O_98,N_16394,N_17264);
and UO_99 (O_99,N_16269,N_19291);
nor UO_100 (O_100,N_15668,N_19365);
xor UO_101 (O_101,N_19052,N_15094);
nand UO_102 (O_102,N_18574,N_19309);
nor UO_103 (O_103,N_17130,N_15117);
or UO_104 (O_104,N_18043,N_16060);
nand UO_105 (O_105,N_17095,N_17146);
and UO_106 (O_106,N_18459,N_16811);
nand UO_107 (O_107,N_15383,N_17936);
or UO_108 (O_108,N_17086,N_15950);
nor UO_109 (O_109,N_19923,N_17494);
nor UO_110 (O_110,N_18193,N_17712);
or UO_111 (O_111,N_16779,N_18843);
nor UO_112 (O_112,N_16495,N_19625);
or UO_113 (O_113,N_18468,N_17976);
nand UO_114 (O_114,N_15691,N_19642);
and UO_115 (O_115,N_16228,N_19410);
or UO_116 (O_116,N_17252,N_18635);
nand UO_117 (O_117,N_15768,N_16446);
or UO_118 (O_118,N_15600,N_19891);
nor UO_119 (O_119,N_16416,N_17347);
or UO_120 (O_120,N_17553,N_16839);
or UO_121 (O_121,N_18979,N_15750);
or UO_122 (O_122,N_17947,N_17226);
nor UO_123 (O_123,N_16898,N_17806);
and UO_124 (O_124,N_19604,N_15275);
and UO_125 (O_125,N_17675,N_16908);
nor UO_126 (O_126,N_19544,N_18178);
and UO_127 (O_127,N_19898,N_16101);
or UO_128 (O_128,N_17516,N_16214);
or UO_129 (O_129,N_16038,N_16652);
and UO_130 (O_130,N_18710,N_15150);
nand UO_131 (O_131,N_16133,N_18144);
or UO_132 (O_132,N_17693,N_18575);
and UO_133 (O_133,N_16925,N_19438);
nor UO_134 (O_134,N_15073,N_17442);
or UO_135 (O_135,N_15134,N_15951);
nand UO_136 (O_136,N_17106,N_18341);
nor UO_137 (O_137,N_17598,N_18854);
or UO_138 (O_138,N_16213,N_18770);
and UO_139 (O_139,N_18728,N_19730);
or UO_140 (O_140,N_17413,N_18823);
nor UO_141 (O_141,N_15247,N_16428);
nand UO_142 (O_142,N_19476,N_16143);
and UO_143 (O_143,N_15386,N_16603);
nand UO_144 (O_144,N_19515,N_18706);
and UO_145 (O_145,N_18492,N_18600);
and UO_146 (O_146,N_18098,N_19094);
nand UO_147 (O_147,N_16094,N_17316);
nor UO_148 (O_148,N_17338,N_19750);
nor UO_149 (O_149,N_16482,N_19763);
and UO_150 (O_150,N_15853,N_17439);
nand UO_151 (O_151,N_16784,N_18572);
or UO_152 (O_152,N_15542,N_18374);
nor UO_153 (O_153,N_19705,N_19151);
nand UO_154 (O_154,N_19688,N_17622);
and UO_155 (O_155,N_18458,N_17758);
xor UO_156 (O_156,N_18528,N_17389);
and UO_157 (O_157,N_19170,N_15485);
nor UO_158 (O_158,N_19183,N_19072);
nor UO_159 (O_159,N_16453,N_19379);
and UO_160 (O_160,N_17081,N_18957);
and UO_161 (O_161,N_18460,N_19847);
nand UO_162 (O_162,N_17096,N_15850);
and UO_163 (O_163,N_15541,N_19453);
or UO_164 (O_164,N_19912,N_16934);
nor UO_165 (O_165,N_15612,N_16668);
nor UO_166 (O_166,N_18427,N_18303);
and UO_167 (O_167,N_18324,N_16945);
xnor UO_168 (O_168,N_19452,N_15451);
or UO_169 (O_169,N_18820,N_19185);
or UO_170 (O_170,N_17714,N_18525);
and UO_171 (O_171,N_15112,N_17650);
xor UO_172 (O_172,N_19601,N_18570);
xnor UO_173 (O_173,N_17193,N_16760);
nand UO_174 (O_174,N_16575,N_17489);
nand UO_175 (O_175,N_17968,N_18452);
or UO_176 (O_176,N_18931,N_18124);
or UO_177 (O_177,N_16506,N_19570);
or UO_178 (O_178,N_17916,N_17454);
nor UO_179 (O_179,N_15714,N_16167);
nor UO_180 (O_180,N_15375,N_15622);
nand UO_181 (O_181,N_17566,N_19609);
xnor UO_182 (O_182,N_19004,N_15593);
or UO_183 (O_183,N_17372,N_17979);
nand UO_184 (O_184,N_18423,N_19612);
or UO_185 (O_185,N_18204,N_16004);
xnor UO_186 (O_186,N_16966,N_18404);
nor UO_187 (O_187,N_15436,N_16984);
nand UO_188 (O_188,N_17245,N_19543);
nand UO_189 (O_189,N_18559,N_18142);
nand UO_190 (O_190,N_16700,N_15458);
nand UO_191 (O_191,N_18059,N_15629);
and UO_192 (O_192,N_16472,N_15828);
nand UO_193 (O_193,N_19779,N_18531);
and UO_194 (O_194,N_17846,N_18775);
and UO_195 (O_195,N_16821,N_17696);
and UO_196 (O_196,N_18798,N_15425);
nor UO_197 (O_197,N_15012,N_16914);
xnor UO_198 (O_198,N_19533,N_16009);
nand UO_199 (O_199,N_15394,N_19769);
and UO_200 (O_200,N_18271,N_18762);
nor UO_201 (O_201,N_15734,N_19082);
nand UO_202 (O_202,N_17896,N_17573);
or UO_203 (O_203,N_19103,N_16666);
or UO_204 (O_204,N_17395,N_17400);
xnor UO_205 (O_205,N_18319,N_18234);
xor UO_206 (O_206,N_16347,N_15329);
or UO_207 (O_207,N_15912,N_18147);
nor UO_208 (O_208,N_19501,N_15062);
nand UO_209 (O_209,N_18510,N_19125);
or UO_210 (O_210,N_18593,N_16067);
or UO_211 (O_211,N_16551,N_18129);
nor UO_212 (O_212,N_15043,N_17240);
nand UO_213 (O_213,N_16146,N_16541);
or UO_214 (O_214,N_18214,N_18385);
nor UO_215 (O_215,N_15392,N_19836);
xor UO_216 (O_216,N_19765,N_16826);
or UO_217 (O_217,N_18900,N_15308);
nand UO_218 (O_218,N_15606,N_19484);
or UO_219 (O_219,N_16783,N_17263);
nand UO_220 (O_220,N_19767,N_16404);
nor UO_221 (O_221,N_19641,N_15754);
nand UO_222 (O_222,N_16522,N_19386);
nor UO_223 (O_223,N_18477,N_17565);
nor UO_224 (O_224,N_15182,N_17753);
nor UO_225 (O_225,N_19648,N_16650);
nor UO_226 (O_226,N_17967,N_19305);
xnor UO_227 (O_227,N_15670,N_17910);
nor UO_228 (O_228,N_17772,N_19083);
nand UO_229 (O_229,N_16647,N_19711);
and UO_230 (O_230,N_15241,N_19924);
nor UO_231 (O_231,N_15642,N_16903);
xnor UO_232 (O_232,N_16419,N_16496);
nor UO_233 (O_233,N_16261,N_19855);
nor UO_234 (O_234,N_18225,N_15789);
and UO_235 (O_235,N_19640,N_19186);
nand UO_236 (O_236,N_18978,N_17776);
nor UO_237 (O_237,N_18096,N_15786);
nand UO_238 (O_238,N_16855,N_19347);
and UO_239 (O_239,N_16828,N_16562);
and UO_240 (O_240,N_17645,N_16528);
nor UO_241 (O_241,N_19917,N_16020);
or UO_242 (O_242,N_16103,N_15369);
nor UO_243 (O_243,N_15030,N_18674);
nand UO_244 (O_244,N_15989,N_18479);
nor UO_245 (O_245,N_16178,N_16462);
xor UO_246 (O_246,N_18307,N_18306);
nor UO_247 (O_247,N_19279,N_18425);
nor UO_248 (O_248,N_19736,N_17254);
nor UO_249 (O_249,N_15290,N_19393);
nor UO_250 (O_250,N_16356,N_15501);
nand UO_251 (O_251,N_16871,N_19586);
or UO_252 (O_252,N_17288,N_17717);
or UO_253 (O_253,N_15505,N_15376);
or UO_254 (O_254,N_16362,N_17517);
nand UO_255 (O_255,N_15400,N_19576);
nor UO_256 (O_256,N_18045,N_15128);
nor UO_257 (O_257,N_15005,N_17195);
nor UO_258 (O_258,N_16186,N_16113);
nand UO_259 (O_259,N_17500,N_15996);
or UO_260 (O_260,N_18401,N_16770);
or UO_261 (O_261,N_15384,N_15413);
or UO_262 (O_262,N_16217,N_18015);
and UO_263 (O_263,N_15255,N_18007);
and UO_264 (O_264,N_15923,N_17690);
nand UO_265 (O_265,N_16274,N_17027);
nor UO_266 (O_266,N_15669,N_16011);
nor UO_267 (O_267,N_16919,N_16245);
nor UO_268 (O_268,N_17983,N_16753);
nor UO_269 (O_269,N_17302,N_16258);
nor UO_270 (O_270,N_17041,N_17019);
nand UO_271 (O_271,N_16249,N_17278);
nand UO_272 (O_272,N_16985,N_16293);
nor UO_273 (O_273,N_15237,N_15114);
xnor UO_274 (O_274,N_18000,N_16606);
or UO_275 (O_275,N_15124,N_15328);
nor UO_276 (O_276,N_15561,N_17354);
or UO_277 (O_277,N_19949,N_19588);
and UO_278 (O_278,N_15157,N_15017);
or UO_279 (O_279,N_18365,N_18328);
nand UO_280 (O_280,N_18772,N_18785);
xnor UO_281 (O_281,N_16659,N_19193);
nor UO_282 (O_282,N_18236,N_16092);
or UO_283 (O_283,N_19230,N_17416);
and UO_284 (O_284,N_15105,N_19323);
nand UO_285 (O_285,N_15565,N_15686);
or UO_286 (O_286,N_16181,N_18373);
and UO_287 (O_287,N_17341,N_18199);
or UO_288 (O_288,N_16664,N_19038);
nor UO_289 (O_289,N_16790,N_19413);
xor UO_290 (O_290,N_19714,N_16165);
nand UO_291 (O_291,N_16492,N_16736);
or UO_292 (O_292,N_15398,N_15722);
and UO_293 (O_293,N_17887,N_15886);
or UO_294 (O_294,N_18230,N_17861);
and UO_295 (O_295,N_18987,N_19455);
xor UO_296 (O_296,N_15528,N_15904);
nor UO_297 (O_297,N_16709,N_17411);
or UO_298 (O_298,N_16118,N_17966);
nor UO_299 (O_299,N_16987,N_16380);
nor UO_300 (O_300,N_16024,N_19169);
nor UO_301 (O_301,N_15966,N_17954);
or UO_302 (O_302,N_19590,N_16333);
nand UO_303 (O_303,N_16577,N_18431);
xnor UO_304 (O_304,N_15003,N_17602);
or UO_305 (O_305,N_15067,N_18849);
and UO_306 (O_306,N_16954,N_18722);
or UO_307 (O_307,N_17745,N_16532);
and UO_308 (O_308,N_16277,N_19848);
nor UO_309 (O_309,N_15470,N_17939);
nor UO_310 (O_310,N_18585,N_16629);
nor UO_311 (O_311,N_19360,N_16849);
nor UO_312 (O_312,N_17178,N_15184);
and UO_313 (O_313,N_17784,N_17535);
and UO_314 (O_314,N_19519,N_15305);
nor UO_315 (O_315,N_19416,N_16051);
and UO_316 (O_316,N_16007,N_15295);
nor UO_317 (O_317,N_16690,N_16632);
and UO_318 (O_318,N_15637,N_15998);
xnor UO_319 (O_319,N_18551,N_16438);
and UO_320 (O_320,N_15427,N_17202);
and UO_321 (O_321,N_16158,N_18002);
or UO_322 (O_322,N_15995,N_19464);
xor UO_323 (O_323,N_15796,N_16711);
nor UO_324 (O_324,N_17660,N_19180);
or UO_325 (O_325,N_16157,N_17459);
nand UO_326 (O_326,N_19943,N_18629);
nand UO_327 (O_327,N_18241,N_16595);
or UO_328 (O_328,N_17682,N_18380);
and UO_329 (O_329,N_16076,N_18447);
nand UO_330 (O_330,N_15264,N_18504);
nor UO_331 (O_331,N_15939,N_19270);
nor UO_332 (O_332,N_16266,N_15937);
nand UO_333 (O_333,N_15719,N_16408);
nor UO_334 (O_334,N_18871,N_15534);
nand UO_335 (O_335,N_18121,N_18542);
nor UO_336 (O_336,N_18801,N_17345);
or UO_337 (O_337,N_18143,N_19035);
and UO_338 (O_338,N_16893,N_18515);
nand UO_339 (O_339,N_15898,N_19794);
or UO_340 (O_340,N_16122,N_15683);
nor UO_341 (O_341,N_16489,N_17749);
and UO_342 (O_342,N_19733,N_16470);
nand UO_343 (O_343,N_15663,N_18347);
and UO_344 (O_344,N_17546,N_16992);
and UO_345 (O_345,N_18195,N_19080);
nor UO_346 (O_346,N_15658,N_19175);
and UO_347 (O_347,N_17754,N_16069);
xor UO_348 (O_348,N_18004,N_19036);
nand UO_349 (O_349,N_16973,N_17706);
nand UO_350 (O_350,N_19111,N_16995);
nand UO_351 (O_351,N_16110,N_16799);
xnor UO_352 (O_352,N_16808,N_18461);
nor UO_353 (O_353,N_17577,N_17528);
xor UO_354 (O_354,N_19530,N_17775);
or UO_355 (O_355,N_16542,N_15782);
or UO_356 (O_356,N_18298,N_17642);
and UO_357 (O_357,N_15679,N_19317);
or UO_358 (O_358,N_16128,N_17656);
or UO_359 (O_359,N_16511,N_18716);
or UO_360 (O_360,N_16382,N_16993);
nand UO_361 (O_361,N_16504,N_16791);
nor UO_362 (O_362,N_18284,N_15818);
nor UO_363 (O_363,N_15917,N_19339);
nor UO_364 (O_364,N_15446,N_16544);
or UO_365 (O_365,N_18450,N_19746);
or UO_366 (O_366,N_15300,N_19177);
xnor UO_367 (O_367,N_19579,N_18437);
nand UO_368 (O_368,N_15029,N_17687);
nand UO_369 (O_369,N_15071,N_16980);
nand UO_370 (O_370,N_19137,N_19838);
or UO_371 (O_371,N_18120,N_18929);
and UO_372 (O_372,N_19292,N_18311);
nor UO_373 (O_373,N_17209,N_16454);
or UO_374 (O_374,N_15849,N_17467);
nor UO_375 (O_375,N_17369,N_19349);
or UO_376 (O_376,N_19271,N_19422);
xnor UO_377 (O_377,N_19277,N_18289);
nor UO_378 (O_378,N_16106,N_19974);
or UO_379 (O_379,N_19600,N_19716);
or UO_380 (O_380,N_17107,N_18262);
nand UO_381 (O_381,N_18731,N_18787);
nor UO_382 (O_382,N_19404,N_16895);
and UO_383 (O_383,N_17931,N_15048);
or UO_384 (O_384,N_17904,N_19626);
nor UO_385 (O_385,N_18997,N_18272);
or UO_386 (O_386,N_17621,N_19272);
and UO_387 (O_387,N_19665,N_17868);
and UO_388 (O_388,N_15449,N_18906);
nand UO_389 (O_389,N_18249,N_18872);
nor UO_390 (O_390,N_19099,N_18680);
or UO_391 (O_391,N_15066,N_19918);
or UO_392 (O_392,N_15142,N_18985);
or UO_393 (O_393,N_15438,N_17762);
nand UO_394 (O_394,N_16918,N_19163);
or UO_395 (O_395,N_15033,N_17938);
nor UO_396 (O_396,N_19583,N_16003);
or UO_397 (O_397,N_17587,N_19995);
nor UO_398 (O_398,N_19408,N_18500);
nor UO_399 (O_399,N_17972,N_16148);
or UO_400 (O_400,N_17453,N_16349);
nor UO_401 (O_401,N_19247,N_16256);
nand UO_402 (O_402,N_15655,N_17928);
or UO_403 (O_403,N_19265,N_18133);
nor UO_404 (O_404,N_15881,N_19773);
nand UO_405 (O_405,N_17379,N_16057);
or UO_406 (O_406,N_19031,N_18304);
and UO_407 (O_407,N_16874,N_16398);
nor UO_408 (O_408,N_17492,N_15633);
nor UO_409 (O_409,N_19929,N_18153);
and UO_410 (O_410,N_16593,N_15316);
nand UO_411 (O_411,N_18718,N_16396);
or UO_412 (O_412,N_17797,N_15894);
or UO_413 (O_413,N_19011,N_16225);
and UO_414 (O_414,N_15169,N_15601);
nand UO_415 (O_415,N_17985,N_17215);
or UO_416 (O_416,N_16538,N_17958);
nand UO_417 (O_417,N_19024,N_19826);
nor UO_418 (O_418,N_17483,N_19800);
nor UO_419 (O_419,N_19694,N_16040);
or UO_420 (O_420,N_19028,N_19092);
or UO_421 (O_421,N_16109,N_15829);
nor UO_422 (O_422,N_19203,N_15050);
or UO_423 (O_423,N_16765,N_19692);
xnor UO_424 (O_424,N_16121,N_19657);
nor UO_425 (O_425,N_15190,N_19584);
or UO_426 (O_426,N_15483,N_16221);
nor UO_427 (O_427,N_19109,N_15877);
or UO_428 (O_428,N_15479,N_15672);
nor UO_429 (O_429,N_19511,N_18959);
nor UO_430 (O_430,N_17310,N_19234);
nor UO_431 (O_431,N_19454,N_19402);
and UO_432 (O_432,N_17863,N_19059);
or UO_433 (O_433,N_15282,N_18232);
nor UO_434 (O_434,N_18387,N_19598);
nand UO_435 (O_435,N_17282,N_17343);
and UO_436 (O_436,N_17079,N_18821);
nand UO_437 (O_437,N_18875,N_15311);
xor UO_438 (O_438,N_19118,N_17231);
xnor UO_439 (O_439,N_18091,N_17153);
nor UO_440 (O_440,N_19421,N_16884);
or UO_441 (O_441,N_18526,N_19482);
nor UO_442 (O_442,N_18081,N_17190);
and UO_443 (O_443,N_19362,N_18818);
or UO_444 (O_444,N_17789,N_18806);
nand UO_445 (O_445,N_15559,N_19479);
nand UO_446 (O_446,N_18683,N_19263);
xnor UO_447 (O_447,N_15721,N_18615);
nand UO_448 (O_448,N_18784,N_16055);
nand UO_449 (O_449,N_16230,N_19034);
nand UO_450 (O_450,N_15034,N_16655);
nand UO_451 (O_451,N_18565,N_17234);
xnor UO_452 (O_452,N_18248,N_19715);
nand UO_453 (O_453,N_15560,N_19162);
or UO_454 (O_454,N_17920,N_19131);
nand UO_455 (O_455,N_15803,N_18960);
nand UO_456 (O_456,N_16291,N_15374);
nand UO_457 (O_457,N_19329,N_19245);
nor UO_458 (O_458,N_17230,N_17544);
xor UO_459 (O_459,N_18989,N_17760);
and UO_460 (O_460,N_18625,N_17606);
nand UO_461 (O_461,N_16235,N_17647);
or UO_462 (O_462,N_17834,N_19850);
xor UO_463 (O_463,N_18323,N_19723);
and UO_464 (O_464,N_15138,N_16490);
nand UO_465 (O_465,N_19948,N_19123);
or UO_466 (O_466,N_18894,N_16570);
nor UO_467 (O_467,N_18107,N_16077);
and UO_468 (O_468,N_17104,N_19889);
xnor UO_469 (O_469,N_17249,N_15661);
or UO_470 (O_470,N_15699,N_18422);
or UO_471 (O_471,N_16427,N_17375);
and UO_472 (O_472,N_18383,N_17255);
nor UO_473 (O_473,N_15429,N_16145);
nor UO_474 (O_474,N_15580,N_19026);
nor UO_475 (O_475,N_19631,N_16292);
and UO_476 (O_476,N_18354,N_17550);
and UO_477 (O_477,N_15656,N_17114);
and UO_478 (O_478,N_18840,N_16284);
xnor UO_479 (O_479,N_19150,N_18973);
and UO_480 (O_480,N_16034,N_17225);
nor UO_481 (O_481,N_18630,N_16717);
nor UO_482 (O_482,N_16176,N_15246);
or UO_483 (O_483,N_16188,N_15968);
nor UO_484 (O_484,N_16124,N_19105);
nand UO_485 (O_485,N_17363,N_15481);
nor UO_486 (O_486,N_17262,N_17362);
nor UO_487 (O_487,N_19507,N_18657);
nand UO_488 (O_488,N_19450,N_19108);
or UO_489 (O_489,N_19634,N_16545);
nor UO_490 (O_490,N_18981,N_15940);
xor UO_491 (O_491,N_16326,N_17638);
or UO_492 (O_492,N_19961,N_18339);
or UO_493 (O_493,N_18218,N_16212);
and UO_494 (O_494,N_16373,N_19469);
and UO_495 (O_495,N_18123,N_16000);
or UO_496 (O_496,N_18656,N_17791);
xnor UO_497 (O_497,N_18317,N_15727);
nand UO_498 (O_498,N_17608,N_19156);
nand UO_499 (O_499,N_16957,N_19729);
and UO_500 (O_500,N_16848,N_17946);
nor UO_501 (O_501,N_17876,N_16521);
and UO_502 (O_502,N_18435,N_16015);
nor UO_503 (O_503,N_19471,N_19549);
xnor UO_504 (O_504,N_17893,N_18895);
xnor UO_505 (O_505,N_18448,N_19431);
or UO_506 (O_506,N_17232,N_15931);
nor UO_507 (O_507,N_19468,N_16758);
nor UO_508 (O_508,N_16132,N_15028);
nor UO_509 (O_509,N_15903,N_19037);
xnor UO_510 (O_510,N_16503,N_17468);
nand UO_511 (O_511,N_18223,N_19005);
nand UO_512 (O_512,N_17816,N_18267);
nor UO_513 (O_513,N_19216,N_17881);
nor UO_514 (O_514,N_15706,N_15567);
nor UO_515 (O_515,N_17429,N_18742);
nand UO_516 (O_516,N_17378,N_17061);
and UO_517 (O_517,N_16889,N_16456);
or UO_518 (O_518,N_17640,N_16519);
nor UO_519 (O_519,N_19493,N_19359);
nor UO_520 (O_520,N_15546,N_17512);
nor UO_521 (O_521,N_15570,N_17891);
nand UO_522 (O_522,N_17785,N_19983);
or UO_523 (O_523,N_18412,N_16680);
or UO_524 (O_524,N_19330,N_18527);
xnor UO_525 (O_525,N_16968,N_16752);
nor UO_526 (O_526,N_19089,N_17037);
and UO_527 (O_527,N_16805,N_19223);
nand UO_528 (O_528,N_17307,N_18835);
and UO_529 (O_529,N_17488,N_18647);
and UO_530 (O_530,N_15231,N_19592);
or UO_531 (O_531,N_19646,N_17381);
or UO_532 (O_532,N_19409,N_19555);
nand UO_533 (O_533,N_18508,N_19157);
nor UO_534 (O_534,N_19888,N_19407);
nand UO_535 (O_535,N_15868,N_15964);
nor UO_536 (O_536,N_15098,N_16278);
nand UO_537 (O_537,N_15822,N_19435);
or UO_538 (O_538,N_15675,N_15920);
or UO_539 (O_539,N_18512,N_17470);
or UO_540 (O_540,N_17836,N_19858);
or UO_541 (O_541,N_15576,N_18663);
xnor UO_542 (O_542,N_17874,N_15678);
and UO_543 (O_543,N_15445,N_19557);
nor UO_544 (O_544,N_16243,N_19066);
or UO_545 (O_545,N_17408,N_16164);
and UO_546 (O_546,N_19202,N_17164);
and UO_547 (O_547,N_19232,N_15957);
or UO_548 (O_548,N_17698,N_18109);
nand UO_549 (O_549,N_18345,N_17591);
nand UO_550 (O_550,N_19577,N_17907);
nor UO_551 (O_551,N_18740,N_15696);
nor UO_552 (O_552,N_19085,N_16241);
nor UO_553 (O_553,N_18012,N_17093);
or UO_554 (O_554,N_18598,N_19167);
nor UO_555 (O_555,N_16442,N_19251);
and UO_556 (O_556,N_18294,N_17770);
and UO_557 (O_557,N_18761,N_15636);
nor UO_558 (O_558,N_16327,N_19816);
nor UO_559 (O_559,N_17685,N_15245);
nor UO_560 (O_560,N_19905,N_17905);
and UO_561 (O_561,N_16719,N_19593);
or UO_562 (O_562,N_18472,N_15417);
or UO_563 (O_563,N_15702,N_19972);
nand UO_564 (O_564,N_16913,N_17665);
or UO_565 (O_565,N_15981,N_19211);
nand UO_566 (O_566,N_18242,N_17619);
or UO_567 (O_567,N_15503,N_17561);
and UO_568 (O_568,N_17455,N_16702);
or UO_569 (O_569,N_17197,N_15393);
xnor UO_570 (O_570,N_19116,N_17253);
or UO_571 (O_571,N_17039,N_18976);
nand UO_572 (O_572,N_19938,N_15103);
nand UO_573 (O_573,N_18372,N_19776);
or UO_574 (O_574,N_18163,N_18170);
and UO_575 (O_575,N_17515,N_16182);
nand UO_576 (O_576,N_17035,N_15586);
or UO_577 (O_577,N_16673,N_18613);
nor UO_578 (O_578,N_17036,N_15059);
or UO_579 (O_579,N_15910,N_17060);
xnor UO_580 (O_580,N_18224,N_15487);
nand UO_581 (O_581,N_15836,N_18974);
nor UO_582 (O_582,N_18569,N_15557);
xor UO_583 (O_583,N_15709,N_15327);
and UO_584 (O_584,N_18019,N_18776);
or UO_585 (O_585,N_18865,N_15880);
and UO_586 (O_586,N_17601,N_16645);
or UO_587 (O_587,N_15424,N_18078);
nand UO_588 (O_588,N_19445,N_17290);
nand UO_589 (O_589,N_15990,N_17563);
and UO_590 (O_590,N_19048,N_15397);
or UO_591 (O_591,N_16836,N_17653);
nand UO_592 (O_592,N_19664,N_16204);
nor UO_593 (O_593,N_15960,N_16086);
nand UO_594 (O_594,N_18364,N_15211);
xor UO_595 (O_595,N_16052,N_18501);
nand UO_596 (O_596,N_15974,N_19927);
nor UO_597 (O_597,N_16642,N_18049);
or UO_598 (O_598,N_18975,N_15891);
nand UO_599 (O_599,N_16232,N_16596);
and UO_600 (O_600,N_15725,N_16377);
or UO_601 (O_601,N_19171,N_19346);
or UO_602 (O_602,N_17809,N_15843);
nor UO_603 (O_603,N_17593,N_15623);
and UO_604 (O_604,N_19496,N_16295);
nor UO_605 (O_605,N_18090,N_19456);
nand UO_606 (O_606,N_18587,N_15813);
or UO_607 (O_607,N_17630,N_17751);
and UO_608 (O_608,N_15145,N_17300);
and UO_609 (O_609,N_17764,N_18075);
or UO_610 (O_610,N_18602,N_19206);
or UO_611 (O_611,N_18333,N_15293);
nor UO_612 (O_612,N_15025,N_16683);
nor UO_613 (O_613,N_16621,N_17995);
nor UO_614 (O_614,N_16728,N_19808);
nand UO_615 (O_615,N_15665,N_19267);
nor UO_616 (O_616,N_17547,N_15262);
or UO_617 (O_617,N_18607,N_19481);
xnor UO_618 (O_618,N_17298,N_16072);
and UO_619 (O_619,N_18273,N_15482);
nand UO_620 (O_620,N_16097,N_17847);
xor UO_621 (O_621,N_15892,N_16977);
nand UO_622 (O_622,N_19757,N_17668);
nor UO_623 (O_623,N_19785,N_17212);
nor UO_624 (O_624,N_17978,N_16566);
or UO_625 (O_625,N_15102,N_18868);
and UO_626 (O_626,N_18064,N_19227);
nor UO_627 (O_627,N_17756,N_16437);
xnor UO_628 (O_628,N_15188,N_16071);
nor UO_629 (O_629,N_19522,N_19260);
nor UO_630 (O_630,N_18650,N_17138);
nand UO_631 (O_631,N_16952,N_15224);
and UO_632 (O_632,N_15140,N_19119);
nand UO_633 (O_633,N_18111,N_16956);
nand UO_634 (O_634,N_15615,N_19742);
or UO_635 (O_635,N_19751,N_18521);
nor UO_636 (O_636,N_18669,N_19671);
nor UO_637 (O_637,N_18118,N_18922);
or UO_638 (O_638,N_15947,N_16107);
xor UO_639 (O_639,N_16580,N_19325);
xnor UO_640 (O_640,N_18055,N_17508);
and UO_641 (O_641,N_17157,N_16986);
and UO_642 (O_642,N_15022,N_15191);
nor UO_643 (O_643,N_15302,N_15074);
or UO_644 (O_644,N_15092,N_19636);
or UO_645 (O_645,N_17004,N_19397);
nand UO_646 (O_646,N_18148,N_16065);
and UO_647 (O_647,N_18950,N_16486);
or UO_648 (O_648,N_16411,N_18554);
xor UO_649 (O_649,N_18314,N_19965);
nor UO_650 (O_650,N_16131,N_16798);
xor UO_651 (O_651,N_16775,N_15893);
and UO_652 (O_652,N_18595,N_17128);
nand UO_653 (O_653,N_16878,N_17103);
or UO_654 (O_654,N_16318,N_17094);
nor UO_655 (O_655,N_15391,N_17926);
and UO_656 (O_656,N_16413,N_16981);
xor UO_657 (O_657,N_16117,N_19134);
or UO_658 (O_658,N_16731,N_15196);
or UO_659 (O_659,N_17915,N_16620);
or UO_660 (O_660,N_18637,N_18139);
or UO_661 (O_661,N_16426,N_18949);
xor UO_662 (O_662,N_15513,N_15827);
nor UO_663 (O_663,N_17330,N_19148);
and UO_664 (O_664,N_15530,N_19718);
nor UO_665 (O_665,N_15288,N_18890);
nor UO_666 (O_666,N_19000,N_18540);
or UO_667 (O_667,N_18882,N_18523);
nand UO_668 (O_668,N_19192,N_19815);
nand UO_669 (O_669,N_17664,N_16890);
nand UO_670 (O_670,N_16355,N_16524);
nand UO_671 (O_671,N_17367,N_15592);
and UO_672 (O_672,N_17089,N_19936);
nor UO_673 (O_673,N_19115,N_15144);
nand UO_674 (O_674,N_19906,N_16397);
nand UO_675 (O_675,N_19663,N_15403);
or UO_676 (O_676,N_18379,N_16090);
or UO_677 (O_677,N_19225,N_17855);
nand UO_678 (O_678,N_16194,N_17883);
nor UO_679 (O_679,N_15654,N_17718);
or UO_680 (O_680,N_15765,N_16806);
nor UO_681 (O_681,N_16942,N_18621);
and UO_682 (O_682,N_17047,N_19401);
nor UO_683 (O_683,N_16520,N_16894);
nand UO_684 (O_684,N_16592,N_19320);
and UO_685 (O_685,N_15421,N_19176);
nor UO_686 (O_686,N_18037,N_17236);
or UO_687 (O_687,N_17496,N_15621);
nand UO_688 (O_688,N_16646,N_18888);
and UO_689 (O_689,N_15283,N_15504);
nor UO_690 (O_690,N_15626,N_18320);
or UO_691 (O_691,N_19789,N_19285);
or UO_692 (O_692,N_16321,N_18903);
nor UO_693 (O_693,N_16403,N_16788);
or UO_694 (O_694,N_16559,N_15348);
or UO_695 (O_695,N_17139,N_18179);
and UO_696 (O_696,N_16634,N_17497);
or UO_697 (O_697,N_19166,N_15006);
nand UO_698 (O_698,N_17447,N_15724);
or UO_699 (O_699,N_15506,N_16483);
nor UO_700 (O_700,N_19508,N_15200);
nand UO_701 (O_701,N_17180,N_16587);
nand UO_702 (O_702,N_19467,N_16643);
xnor UO_703 (O_703,N_18842,N_19568);
xnor UO_704 (O_704,N_16846,N_19348);
nand UO_705 (O_705,N_17850,N_15862);
nand UO_706 (O_706,N_15676,N_18632);
nor UO_707 (O_707,N_17703,N_19683);
or UO_708 (O_708,N_17010,N_16313);
or UO_709 (O_709,N_16179,N_19315);
nand UO_710 (O_710,N_16390,N_19686);
and UO_711 (O_711,N_15780,N_16727);
and UO_712 (O_712,N_17360,N_19740);
or UO_713 (O_713,N_18817,N_18047);
or UO_714 (O_714,N_16105,N_19212);
and UO_715 (O_715,N_17988,N_19158);
xnor UO_716 (O_716,N_17299,N_18485);
nand UO_717 (O_717,N_17530,N_16191);
or UO_718 (O_718,N_15396,N_17799);
or UO_719 (O_719,N_18863,N_16560);
nand UO_720 (O_720,N_19253,N_17989);
or UO_721 (O_721,N_18287,N_15091);
or UO_722 (O_722,N_16762,N_16341);
and UO_723 (O_723,N_15607,N_19529);
nor UO_724 (O_724,N_19316,N_16801);
and UO_725 (O_725,N_15173,N_17617);
nor UO_726 (O_726,N_17308,N_18074);
or UO_727 (O_727,N_15065,N_15550);
xor UO_728 (O_728,N_17551,N_16661);
nor UO_729 (O_729,N_15236,N_15548);
and UO_730 (O_730,N_17506,N_17571);
nand UO_731 (O_731,N_18968,N_16967);
or UO_732 (O_732,N_18507,N_19968);
nand UO_733 (O_733,N_19812,N_17048);
and UO_734 (O_734,N_17585,N_16363);
nor UO_735 (O_735,N_18829,N_15058);
nor UO_736 (O_736,N_15440,N_17366);
or UO_737 (O_737,N_19676,N_18773);
nor UO_738 (O_738,N_15465,N_17805);
and UO_739 (O_739,N_19033,N_17404);
nand UO_740 (O_740,N_18760,N_15463);
or UO_741 (O_741,N_15363,N_15007);
nor UO_742 (O_742,N_16084,N_18874);
nor UO_743 (O_743,N_15355,N_19231);
xor UO_744 (O_744,N_16556,N_16787);
nor UO_745 (O_745,N_18748,N_15153);
nor UO_746 (O_746,N_18308,N_18297);
or UO_747 (O_747,N_16924,N_17445);
xor UO_748 (O_748,N_15377,N_19086);
and UO_749 (O_749,N_16971,N_19633);
and UO_750 (O_750,N_18063,N_16493);
nor UO_751 (O_751,N_15866,N_18207);
or UO_752 (O_752,N_19298,N_17111);
and UO_753 (O_753,N_19728,N_15705);
nand UO_754 (O_754,N_18567,N_18264);
nand UO_755 (O_755,N_15106,N_15326);
nor UO_756 (O_756,N_17440,N_19674);
and UO_757 (O_757,N_19964,N_16869);
and UO_758 (O_758,N_17773,N_16155);
and UO_759 (O_759,N_19226,N_19606);
or UO_760 (O_760,N_15619,N_18336);
or UO_761 (O_761,N_19615,N_16112);
nor UO_762 (O_762,N_19335,N_17574);
or UO_763 (O_763,N_19067,N_17109);
nor UO_764 (O_764,N_16508,N_15013);
and UO_765 (O_765,N_15962,N_15484);
xor UO_766 (O_766,N_18687,N_19284);
nand UO_767 (O_767,N_16755,N_17092);
or UO_768 (O_768,N_17737,N_16299);
nand UO_769 (O_769,N_16424,N_17374);
nand UO_770 (O_770,N_16348,N_16725);
or UO_771 (O_771,N_17556,N_17852);
nand UO_772 (O_772,N_16843,N_16006);
and UO_773 (O_773,N_19910,N_15825);
nor UO_774 (O_774,N_19350,N_18781);
xor UO_775 (O_775,N_16116,N_15121);
nor UO_776 (O_776,N_19425,N_17521);
nand UO_777 (O_777,N_17067,N_16102);
nor UO_778 (O_778,N_17560,N_18789);
nand UO_779 (O_779,N_17123,N_17464);
nor UO_780 (O_780,N_16088,N_16491);
or UO_781 (O_781,N_17370,N_18266);
nor UO_782 (O_782,N_18348,N_15164);
nor UO_783 (O_783,N_18549,N_17023);
and UO_784 (O_784,N_19863,N_16674);
and UO_785 (O_785,N_15076,N_18334);
nor UO_786 (O_786,N_15921,N_16754);
and UO_787 (O_787,N_19516,N_19744);
and UO_788 (O_788,N_17151,N_17851);
nand UO_789 (O_789,N_16166,N_16063);
or UO_790 (O_790,N_17662,N_15332);
nand UO_791 (O_791,N_16921,N_19935);
nor UO_792 (O_792,N_17604,N_16091);
xor UO_793 (O_793,N_15464,N_16053);
xor UO_794 (O_794,N_15432,N_15373);
or UO_795 (O_795,N_16792,N_15867);
nor UO_796 (O_796,N_16608,N_16074);
and UO_797 (O_797,N_19960,N_19210);
and UO_798 (O_798,N_15052,N_15284);
or UO_799 (O_799,N_17819,N_18503);
and UO_800 (O_800,N_15072,N_19217);
nand UO_801 (O_801,N_18725,N_19919);
and UO_802 (O_802,N_19573,N_15993);
nor UO_803 (O_803,N_17879,N_17481);
and UO_804 (O_804,N_18827,N_19874);
xnor UO_805 (O_805,N_19145,N_17539);
xor UO_806 (O_806,N_16582,N_15268);
xor UO_807 (O_807,N_15078,N_19687);
or UO_808 (O_808,N_16343,N_15292);
nand UO_809 (O_809,N_18794,N_15564);
nor UO_810 (O_810,N_17627,N_18171);
nand UO_811 (O_811,N_18001,N_18733);
and UO_812 (O_812,N_18877,N_17732);
nor UO_813 (O_813,N_17336,N_19191);
xor UO_814 (O_814,N_15337,N_17063);
xnor UO_815 (O_815,N_15405,N_19510);
xor UO_816 (O_816,N_16854,N_18227);
or UO_817 (O_817,N_16211,N_17382);
or UO_818 (O_818,N_15791,N_15717);
nand UO_819 (O_819,N_15450,N_16601);
and UO_820 (O_820,N_17200,N_17596);
or UO_821 (O_821,N_15589,N_18029);
nand UO_822 (O_822,N_18858,N_17554);
or UO_823 (O_823,N_19956,N_17844);
nand UO_824 (O_824,N_18646,N_15831);
nor UO_825 (O_825,N_19102,N_18648);
and UO_826 (O_826,N_16134,N_16441);
xor UO_827 (O_827,N_19739,N_16622);
and UO_828 (O_828,N_16026,N_18579);
nand UO_829 (O_829,N_17268,N_18730);
xnor UO_830 (O_830,N_16715,N_18855);
nand UO_831 (O_831,N_17942,N_17043);
xnor UO_832 (O_832,N_17320,N_16774);
nand UO_833 (O_833,N_19238,N_17011);
and UO_834 (O_834,N_16420,N_18359);
nor UO_835 (O_835,N_17294,N_15596);
or UO_836 (O_836,N_17396,N_15587);
or UO_837 (O_837,N_18860,N_16247);
nor UO_838 (O_838,N_18482,N_19797);
nor UO_839 (O_839,N_18788,N_15399);
or UO_840 (O_840,N_16618,N_18653);
xnor UO_841 (O_841,N_17803,N_19509);
or UO_842 (O_842,N_16803,N_19250);
and UO_843 (O_843,N_17716,N_19473);
nor UO_844 (O_844,N_17314,N_16163);
nor UO_845 (O_845,N_15581,N_19857);
and UO_846 (O_846,N_15520,N_16050);
and UO_847 (O_847,N_19822,N_19294);
xor UO_848 (O_848,N_18038,N_17948);
or UO_849 (O_849,N_18209,N_16461);
xor UO_850 (O_850,N_19930,N_15120);
or UO_851 (O_851,N_17295,N_17826);
or UO_852 (O_852,N_18131,N_17297);
nand UO_853 (O_853,N_18488,N_16130);
nor UO_854 (O_854,N_16807,N_18424);
xor UO_855 (O_855,N_19945,N_18927);
nor UO_856 (O_856,N_16336,N_18830);
nor UO_857 (O_857,N_17735,N_18189);
xnor UO_858 (O_858,N_18157,N_17975);
nor UO_859 (O_859,N_19539,N_19023);
nor UO_860 (O_860,N_17499,N_19220);
nor UO_861 (O_861,N_18753,N_17356);
or UO_862 (O_862,N_15963,N_18191);
or UO_863 (O_863,N_18105,N_16525);
nand UO_864 (O_864,N_18259,N_17158);
and UO_865 (O_865,N_15135,N_17015);
nand UO_866 (O_866,N_16307,N_18764);
or UO_867 (O_867,N_15784,N_18357);
nor UO_868 (O_868,N_19065,N_19524);
nand UO_869 (O_869,N_17634,N_19061);
or UO_870 (O_870,N_19367,N_18318);
and UO_871 (O_871,N_19057,N_16431);
xor UO_872 (O_872,N_15583,N_17418);
and UO_873 (O_873,N_19400,N_17446);
and UO_874 (O_874,N_19534,N_17765);
or UO_875 (O_875,N_18432,N_15997);
or UO_876 (O_876,N_16160,N_19160);
and UO_877 (O_877,N_15815,N_19578);
and UO_878 (O_878,N_16820,N_17070);
nor UO_879 (O_879,N_17796,N_19190);
nor UO_880 (O_880,N_19942,N_18697);
or UO_881 (O_881,N_18429,N_18035);
and UO_882 (O_882,N_17423,N_17631);
or UO_883 (O_883,N_18161,N_15020);
or UO_884 (O_884,N_15959,N_19370);
nor UO_885 (O_885,N_16033,N_19461);
or UO_886 (O_886,N_18353,N_17977);
or UO_887 (O_887,N_16460,N_18441);
and UO_888 (O_888,N_18752,N_19764);
and UO_889 (O_889,N_19321,N_19293);
nor UO_890 (O_890,N_19900,N_17051);
and UO_891 (O_891,N_16471,N_18165);
nor UO_892 (O_892,N_18253,N_19278);
and UO_893 (O_893,N_16534,N_15662);
or UO_894 (O_894,N_18793,N_18137);
nor UO_895 (O_895,N_17425,N_17313);
nor UO_896 (O_896,N_16005,N_19499);
nand UO_897 (O_897,N_18636,N_17137);
or UO_898 (O_898,N_17100,N_17527);
nor UO_899 (O_899,N_16218,N_18456);
and UO_900 (O_900,N_16638,N_19628);
nand UO_901 (O_901,N_15228,N_19699);
nand UO_902 (O_902,N_18668,N_15788);
nand UO_903 (O_903,N_15004,N_18463);
xnor UO_904 (O_904,N_18282,N_18106);
xor UO_905 (O_905,N_16694,N_15353);
nand UO_906 (O_906,N_16422,N_16150);
xor UO_907 (O_907,N_19882,N_15069);
nand UO_908 (O_908,N_17925,N_17045);
nand UO_909 (O_909,N_16126,N_15588);
or UO_910 (O_910,N_18739,N_19433);
and UO_911 (O_911,N_19922,N_19915);
nor UO_912 (O_912,N_17734,N_18594);
or UO_913 (O_913,N_17502,N_18491);
nor UO_914 (O_914,N_16429,N_15875);
nor UO_915 (O_915,N_17414,N_17992);
nand UO_916 (O_916,N_16750,N_15086);
or UO_917 (O_917,N_16553,N_17655);
nor UO_918 (O_918,N_16741,N_17085);
or UO_919 (O_919,N_16975,N_18892);
xnor UO_920 (O_920,N_19090,N_19853);
or UO_921 (O_921,N_16350,N_18634);
and UO_922 (O_922,N_16724,N_15130);
nor UO_923 (O_923,N_17584,N_17962);
nor UO_924 (O_924,N_19006,N_16543);
or UO_925 (O_925,N_15242,N_16565);
or UO_926 (O_926,N_17882,N_15848);
or UO_927 (O_927,N_17001,N_17575);
and UO_928 (O_928,N_18146,N_18692);
nor UO_929 (O_929,N_19485,N_18483);
xnor UO_930 (O_930,N_17034,N_17615);
nand UO_931 (O_931,N_16746,N_18809);
and UO_932 (O_932,N_17933,N_19442);
and UO_933 (O_933,N_18493,N_17607);
and UO_934 (O_934,N_17339,N_18813);
nor UO_935 (O_935,N_18834,N_16533);
nor UO_936 (O_936,N_17802,N_18768);
nor UO_937 (O_937,N_17538,N_16947);
nor UO_938 (O_938,N_17579,N_16781);
or UO_939 (O_939,N_17635,N_15175);
nor UO_940 (O_940,N_17471,N_18344);
or UO_941 (O_941,N_16047,N_19351);
nand UO_942 (O_942,N_15949,N_15810);
nor UO_943 (O_943,N_18149,N_19824);
nand UO_944 (O_944,N_17133,N_18726);
nor UO_945 (O_945,N_19703,N_15422);
and UO_946 (O_946,N_19777,N_19492);
nor UO_947 (O_947,N_18396,N_18377);
or UO_948 (O_948,N_17583,N_16494);
and UO_949 (O_949,N_17451,N_19635);
or UO_950 (O_950,N_19772,N_19383);
nor UO_951 (O_951,N_15743,N_17392);
or UO_952 (O_952,N_17219,N_15214);
nor UO_953 (O_953,N_17963,N_17941);
nor UO_954 (O_954,N_19864,N_16714);
nor UO_955 (O_955,N_16328,N_17557);
or UO_956 (O_956,N_16433,N_19165);
nor UO_957 (O_957,N_15770,N_18859);
nand UO_958 (O_958,N_18831,N_15179);
xnor UO_959 (O_959,N_18067,N_15569);
or UO_960 (O_960,N_17610,N_17174);
or UO_961 (O_961,N_19605,N_19846);
and UO_962 (O_962,N_17049,N_17007);
nand UO_963 (O_963,N_19060,N_19643);
nor UO_964 (O_964,N_16505,N_15240);
nor UO_965 (O_965,N_17659,N_16285);
nand UO_966 (O_966,N_18360,N_15842);
or UO_967 (O_967,N_18351,N_18322);
nand UO_968 (O_968,N_17289,N_16823);
nand UO_969 (O_969,N_18198,N_15334);
and UO_970 (O_970,N_19376,N_15899);
nor UO_971 (O_971,N_15523,N_18946);
nor UO_972 (O_972,N_17752,N_19075);
nand UO_973 (O_973,N_18196,N_15933);
nand UO_974 (O_974,N_16999,N_16850);
nand UO_975 (O_975,N_19446,N_16928);
or UO_976 (O_976,N_15468,N_17820);
and UO_977 (O_977,N_19803,N_17325);
xnor UO_978 (O_978,N_15088,N_16537);
nand UO_979 (O_979,N_15010,N_17628);
nand UO_980 (O_980,N_15361,N_19290);
xnor UO_981 (O_981,N_15497,N_16962);
nor UO_982 (O_982,N_19312,N_16193);
nor UO_983 (O_983,N_17449,N_18961);
and UO_984 (O_984,N_15772,N_15518);
and UO_985 (O_985,N_17889,N_19861);
nand UO_986 (O_986,N_17731,N_19457);
nor UO_987 (O_987,N_17000,N_17726);
and UO_988 (O_988,N_16466,N_15143);
nor UO_989 (O_989,N_16574,N_16036);
or UO_990 (O_990,N_16457,N_18547);
nand UO_991 (O_991,N_15119,N_18673);
nor UO_992 (O_992,N_18679,N_16704);
or UO_993 (O_993,N_17217,N_18678);
nor UO_994 (O_994,N_19707,N_18027);
nor UO_995 (O_995,N_18086,N_17709);
or UO_996 (O_996,N_16360,N_19712);
and UO_997 (O_997,N_16367,N_19748);
and UO_998 (O_998,N_15732,N_17597);
or UO_999 (O_999,N_17576,N_19639);
or UO_1000 (O_1000,N_19107,N_17677);
or UO_1001 (O_1001,N_17285,N_15641);
or UO_1002 (O_1002,N_16851,N_18591);
nor UO_1003 (O_1003,N_16941,N_15800);
and UO_1004 (O_1004,N_16757,N_18543);
or UO_1005 (O_1005,N_19303,N_16387);
or UO_1006 (O_1006,N_18754,N_19443);
nor UO_1007 (O_1007,N_19068,N_18802);
and UO_1008 (O_1008,N_16794,N_18022);
or UO_1009 (O_1009,N_18281,N_16936);
nand UO_1010 (O_1010,N_15820,N_16766);
and UO_1011 (O_1011,N_15783,N_19262);
nand UO_1012 (O_1012,N_16391,N_17503);
or UO_1013 (O_1013,N_15994,N_17062);
nand UO_1014 (O_1014,N_19690,N_17402);
nor UO_1015 (O_1015,N_16064,N_19423);
nor UO_1016 (O_1016,N_16742,N_16663);
or UO_1017 (O_1017,N_18623,N_15016);
and UO_1018 (O_1018,N_19710,N_19021);
xnor UO_1019 (O_1019,N_17082,N_15423);
nor UO_1020 (O_1020,N_17064,N_18203);
xnor UO_1021 (O_1021,N_15320,N_16240);
xor UO_1022 (O_1022,N_17038,N_17629);
nor UO_1023 (O_1023,N_17519,N_17435);
nor UO_1024 (O_1024,N_17148,N_15935);
nor UO_1025 (O_1025,N_17867,N_19432);
or UO_1026 (O_1026,N_19113,N_16865);
or UO_1027 (O_1027,N_18449,N_15250);
nand UO_1028 (O_1028,N_16312,N_18369);
or UO_1029 (O_1029,N_16726,N_16469);
nand UO_1030 (O_1030,N_17112,N_19375);
nand UO_1031 (O_1031,N_16059,N_18428);
nand UO_1032 (O_1032,N_18136,N_17397);
nor UO_1033 (O_1033,N_16901,N_15793);
nand UO_1034 (O_1034,N_17875,N_19571);
and UO_1035 (O_1035,N_15046,N_15985);
and UO_1036 (O_1036,N_16099,N_19804);
and UO_1037 (O_1037,N_17129,N_17781);
nand UO_1038 (O_1038,N_18263,N_18972);
and UO_1039 (O_1039,N_17578,N_18392);
or UO_1040 (O_1040,N_18454,N_17999);
or UO_1041 (O_1041,N_16845,N_16628);
or UO_1042 (O_1042,N_19895,N_16374);
and UO_1043 (O_1043,N_15955,N_19384);
nor UO_1044 (O_1044,N_19440,N_18069);
nand UO_1045 (O_1045,N_18642,N_17040);
nand UO_1046 (O_1046,N_17534,N_16436);
and UO_1047 (O_1047,N_18073,N_16793);
nand UO_1048 (O_1048,N_15751,N_15161);
nand UO_1049 (O_1049,N_16693,N_15176);
nand UO_1050 (O_1050,N_17594,N_15922);
nor UO_1051 (O_1051,N_18708,N_19219);
nor UO_1052 (O_1052,N_15752,N_18928);
and UO_1053 (O_1053,N_16847,N_16206);
or UO_1054 (O_1054,N_18268,N_16909);
or UO_1055 (O_1055,N_18803,N_15763);
or UO_1056 (O_1056,N_18502,N_15296);
or UO_1057 (O_1057,N_19542,N_17746);
xor UO_1058 (O_1058,N_18278,N_15608);
or UO_1059 (O_1059,N_18332,N_16115);
nand UO_1060 (O_1060,N_15193,N_16951);
and UO_1061 (O_1061,N_16888,N_19693);
nor UO_1062 (O_1062,N_18750,N_15049);
and UO_1063 (O_1063,N_17960,N_18965);
or UO_1064 (O_1064,N_19719,N_19518);
and UO_1065 (O_1065,N_17211,N_16215);
xnor UO_1066 (O_1066,N_17885,N_19448);
nor UO_1067 (O_1067,N_19369,N_17415);
xor UO_1068 (O_1068,N_16242,N_15343);
nor UO_1069 (O_1069,N_19269,N_18342);
nand UO_1070 (O_1070,N_17996,N_16651);
xnor UO_1071 (O_1071,N_15766,N_18220);
or UO_1072 (O_1072,N_18291,N_19702);
and UO_1073 (O_1073,N_17147,N_15204);
and UO_1074 (O_1074,N_16859,N_17700);
nor UO_1075 (O_1075,N_15604,N_15159);
or UO_1076 (O_1076,N_15566,N_17272);
or UO_1077 (O_1077,N_15444,N_15729);
and UO_1078 (O_1078,N_18796,N_15324);
or UO_1079 (O_1079,N_18846,N_17306);
nor UO_1080 (O_1080,N_17877,N_18084);
or UO_1081 (O_1081,N_16777,N_19827);
and UO_1082 (O_1082,N_16804,N_17788);
nor UO_1083 (O_1083,N_16744,N_18919);
xor UO_1084 (O_1084,N_15806,N_19672);
and UO_1085 (O_1085,N_19428,N_16597);
nor UO_1086 (O_1086,N_15992,N_18519);
nor UO_1087 (O_1087,N_19319,N_19079);
or UO_1088 (O_1088,N_16929,N_15395);
nand UO_1089 (O_1089,N_19441,N_19398);
or UO_1090 (O_1090,N_15286,N_16208);
and UO_1091 (O_1091,N_15499,N_19288);
nand UO_1092 (O_1092,N_16546,N_19944);
or UO_1093 (O_1093,N_15748,N_15666);
or UO_1094 (O_1094,N_18436,N_16459);
and UO_1095 (O_1095,N_19371,N_16079);
or UO_1096 (O_1096,N_16236,N_18413);
or UO_1097 (O_1097,N_18116,N_15402);
and UO_1098 (O_1098,N_18013,N_15488);
nor UO_1099 (O_1099,N_18478,N_17216);
nand UO_1100 (O_1100,N_16319,N_17871);
or UO_1101 (O_1101,N_19993,N_16818);
nand UO_1102 (O_1102,N_16671,N_15716);
nor UO_1103 (O_1103,N_19698,N_17757);
nand UO_1104 (O_1104,N_18720,N_18765);
and UO_1105 (O_1105,N_15897,N_16961);
and UO_1106 (O_1106,N_15206,N_19830);
or UO_1107 (O_1107,N_16607,N_19331);
nand UO_1108 (O_1108,N_16282,N_15199);
nor UO_1109 (O_1109,N_19523,N_16061);
or UO_1110 (O_1110,N_17763,N_18996);
xor UO_1111 (O_1111,N_17825,N_15009);
and UO_1112 (O_1112,N_17465,N_17206);
nor UO_1113 (O_1113,N_17152,N_17088);
nor UO_1114 (O_1114,N_19405,N_19261);
and UO_1115 (O_1115,N_18685,N_16233);
or UO_1116 (O_1116,N_15744,N_17132);
nand UO_1117 (O_1117,N_16227,N_18942);
xnor UO_1118 (O_1118,N_16586,N_19437);
nand UO_1119 (O_1119,N_15253,N_19056);
nor UO_1120 (O_1120,N_17667,N_19904);
or UO_1121 (O_1121,N_16324,N_19194);
nand UO_1122 (O_1122,N_17839,N_17150);
nor UO_1123 (O_1123,N_15410,N_15238);
xnor UO_1124 (O_1124,N_19558,N_18115);
nand UO_1125 (O_1125,N_17993,N_15533);
nand UO_1126 (O_1126,N_18062,N_15147);
or UO_1127 (O_1127,N_16376,N_15599);
nand UO_1128 (O_1128,N_17108,N_15322);
xnor UO_1129 (O_1129,N_18935,N_18050);
nand UO_1130 (O_1130,N_16138,N_17097);
nand UO_1131 (O_1131,N_17845,N_15539);
and UO_1132 (O_1132,N_17678,N_15019);
and UO_1133 (O_1133,N_18522,N_18415);
xnor UO_1134 (O_1134,N_15790,N_19950);
and UO_1135 (O_1135,N_15988,N_17555);
nor UO_1136 (O_1136,N_19809,N_16281);
and UO_1137 (O_1137,N_19536,N_17279);
nand UO_1138 (O_1138,N_17328,N_17116);
nand UO_1139 (O_1139,N_15624,N_19870);
or UO_1140 (O_1140,N_16263,N_15041);
nor UO_1141 (O_1141,N_15370,N_18807);
nand UO_1142 (O_1142,N_19495,N_17600);
nor UO_1143 (O_1143,N_16738,N_19806);
and UO_1144 (O_1144,N_15111,N_16978);
nor UO_1145 (O_1145,N_16583,N_18884);
and UO_1146 (O_1146,N_18723,N_17405);
nand UO_1147 (O_1147,N_17463,N_19801);
or UO_1148 (O_1148,N_17319,N_17029);
and UO_1149 (O_1149,N_15312,N_17854);
and UO_1150 (O_1150,N_17075,N_19791);
or UO_1151 (O_1151,N_15180,N_16448);
and UO_1152 (O_1152,N_18573,N_15808);
nand UO_1153 (O_1153,N_17729,N_18640);
nor UO_1154 (O_1154,N_15170,N_17927);
or UO_1155 (O_1155,N_19382,N_17428);
nor UO_1156 (O_1156,N_15701,N_17741);
and UO_1157 (O_1157,N_19128,N_17124);
xor UO_1158 (O_1158,N_15115,N_15687);
or UO_1159 (O_1159,N_16648,N_15371);
nand UO_1160 (O_1160,N_15532,N_16173);
xnor UO_1161 (O_1161,N_18717,N_15409);
xor UO_1162 (O_1162,N_16156,N_15080);
or UO_1163 (O_1163,N_17203,N_16300);
and UO_1164 (O_1164,N_16008,N_19133);
xnor UO_1165 (O_1165,N_18228,N_16698);
or UO_1166 (O_1166,N_18024,N_15500);
and UO_1167 (O_1167,N_18983,N_17853);
nand UO_1168 (O_1168,N_16435,N_15930);
nor UO_1169 (O_1169,N_17115,N_17970);
xnor UO_1170 (O_1170,N_19095,N_17857);
and UO_1171 (O_1171,N_16665,N_18826);
nor UO_1172 (O_1172,N_17056,N_15256);
and UO_1173 (O_1173,N_16010,N_16778);
nand UO_1174 (O_1174,N_19998,N_19475);
and UO_1175 (O_1175,N_18538,N_17251);
or UO_1176 (O_1176,N_15306,N_15517);
or UO_1177 (O_1177,N_19894,N_17870);
nand UO_1178 (O_1178,N_15977,N_17783);
or UO_1179 (O_1179,N_18470,N_18026);
xor UO_1180 (O_1180,N_18953,N_19091);
and UO_1181 (O_1181,N_18897,N_17837);
nor UO_1182 (O_1182,N_16922,N_18744);
or UO_1183 (O_1183,N_15667,N_17017);
or UO_1184 (O_1184,N_17510,N_19680);
nor UO_1185 (O_1185,N_19093,N_19252);
nand UO_1186 (O_1186,N_19301,N_16672);
nand UO_1187 (O_1187,N_15737,N_18932);
and UO_1188 (O_1188,N_17727,N_19342);
or UO_1189 (O_1189,N_15330,N_19695);
or UO_1190 (O_1190,N_18883,N_15611);
nand UO_1191 (O_1191,N_17894,N_17768);
nor UO_1192 (O_1192,N_19761,N_18544);
nor UO_1193 (O_1193,N_18652,N_15015);
nor UO_1194 (O_1194,N_17177,N_17790);
nor UO_1195 (O_1195,N_15210,N_18280);
nor UO_1196 (O_1196,N_15753,N_18651);
nand UO_1197 (O_1197,N_18481,N_19268);
nand UO_1198 (O_1198,N_19621,N_15510);
xnor UO_1199 (O_1199,N_18495,N_19255);
nor UO_1200 (O_1200,N_17105,N_15053);
xor UO_1201 (O_1201,N_16151,N_17214);
nand UO_1202 (O_1202,N_17266,N_15694);
and UO_1203 (O_1203,N_17207,N_15040);
nor UO_1204 (O_1204,N_18173,N_15833);
and UO_1205 (O_1205,N_19627,N_17744);
nor UO_1206 (O_1206,N_16677,N_15978);
and UO_1207 (O_1207,N_18732,N_18923);
nor UO_1208 (O_1208,N_15919,N_19651);
or UO_1209 (O_1209,N_15133,N_17611);
or UO_1210 (O_1210,N_17616,N_16926);
nor UO_1211 (O_1211,N_19537,N_17163);
nand UO_1212 (O_1212,N_17848,N_16001);
and UO_1213 (O_1213,N_19784,N_16844);
nand UO_1214 (O_1214,N_17318,N_19281);
or UO_1215 (O_1215,N_15938,N_18202);
or UO_1216 (O_1216,N_15644,N_19975);
nor UO_1217 (O_1217,N_19417,N_18638);
nor UO_1218 (O_1218,N_15154,N_17076);
and UO_1219 (O_1219,N_19911,N_19146);
nand UO_1220 (O_1220,N_17472,N_15056);
nor UO_1221 (O_1221,N_19982,N_19720);
nor UO_1222 (O_1222,N_15442,N_16357);
nor UO_1223 (O_1223,N_15755,N_17474);
or UO_1224 (O_1224,N_17077,N_19130);
and UO_1225 (O_1225,N_17974,N_16654);
nor UO_1226 (O_1226,N_19015,N_17823);
nand UO_1227 (O_1227,N_15258,N_19554);
and UO_1228 (O_1228,N_18934,N_17688);
xnor UO_1229 (O_1229,N_16168,N_16624);
or UO_1230 (O_1230,N_17456,N_19009);
and UO_1231 (O_1231,N_18584,N_15884);
nor UO_1232 (O_1232,N_16915,N_17273);
and UO_1233 (O_1233,N_16644,N_17943);
or UO_1234 (O_1234,N_17198,N_18506);
and UO_1235 (O_1235,N_15958,N_15364);
or UO_1236 (O_1236,N_18182,N_18140);
or UO_1237 (O_1237,N_17903,N_15857);
and UO_1238 (O_1238,N_18735,N_15008);
and UO_1239 (O_1239,N_17689,N_17427);
and UO_1240 (O_1240,N_19700,N_17241);
or UO_1241 (O_1241,N_17856,N_18462);
and UO_1242 (O_1242,N_15645,N_15954);
nor UO_1243 (O_1243,N_17980,N_19527);
nor UO_1244 (O_1244,N_16370,N_15340);
and UO_1245 (O_1245,N_15673,N_18285);
or UO_1246 (O_1246,N_19849,N_19840);
or UO_1247 (O_1247,N_16197,N_18690);
nor UO_1248 (O_1248,N_15720,N_16389);
nor UO_1249 (O_1249,N_17589,N_18671);
and UO_1250 (O_1250,N_19209,N_15965);
nor UO_1251 (O_1251,N_15378,N_19833);
or UO_1252 (O_1252,N_18517,N_19834);
nand UO_1253 (O_1253,N_18609,N_18780);
and UO_1254 (O_1254,N_16885,N_17026);
nand UO_1255 (O_1255,N_15183,N_18245);
xor UO_1256 (O_1256,N_19616,N_19283);
nor UO_1257 (O_1257,N_19738,N_17176);
and UO_1258 (O_1258,N_16231,N_19472);
nand UO_1259 (O_1259,N_16479,N_17412);
or UO_1260 (O_1260,N_17277,N_18382);
xor UO_1261 (O_1261,N_15982,N_19896);
or UO_1262 (O_1262,N_18274,N_17432);
and UO_1263 (O_1263,N_15869,N_18618);
nor UO_1264 (O_1264,N_17779,N_19856);
or UO_1265 (O_1265,N_17121,N_19465);
nor UO_1266 (O_1266,N_19637,N_18896);
nor UO_1267 (O_1267,N_17008,N_19396);
or UO_1268 (O_1268,N_15149,N_18782);
nor UO_1269 (O_1269,N_19050,N_18524);
nand UO_1270 (O_1270,N_17537,N_17702);
or UO_1271 (O_1271,N_16619,N_18005);
and UO_1272 (O_1272,N_17003,N_19796);
or UO_1273 (O_1273,N_19673,N_18498);
nand UO_1274 (O_1274,N_17491,N_15494);
and UO_1275 (O_1275,N_16450,N_19820);
and UO_1276 (O_1276,N_18008,N_17167);
xor UO_1277 (O_1277,N_15230,N_18684);
nand UO_1278 (O_1278,N_17859,N_17592);
and UO_1279 (O_1279,N_19868,N_17201);
nand UO_1280 (O_1280,N_16515,N_19899);
or UO_1281 (O_1281,N_18590,N_15814);
xnor UO_1282 (O_1282,N_15812,N_15064);
and UO_1283 (O_1283,N_19914,N_18747);
xnor UO_1284 (O_1284,N_15554,N_18141);
and UO_1285 (O_1285,N_16280,N_16838);
nor UO_1286 (O_1286,N_18925,N_15671);
and UO_1287 (O_1287,N_16623,N_19828);
nand UO_1288 (O_1288,N_17971,N_18641);
nor UO_1289 (O_1289,N_17487,N_15475);
nand UO_1290 (O_1290,N_17466,N_19768);
nor UO_1291 (O_1291,N_19124,N_15801);
nor UO_1292 (O_1292,N_17728,N_17326);
and UO_1293 (O_1293,N_18518,N_16095);
nand UO_1294 (O_1294,N_15616,N_19322);
nand UO_1295 (O_1295,N_17156,N_15244);
or UO_1296 (O_1296,N_18406,N_15591);
and UO_1297 (O_1297,N_16418,N_18962);
and UO_1298 (O_1298,N_15168,N_17849);
nand UO_1299 (O_1299,N_15618,N_17738);
nand UO_1300 (O_1300,N_18913,N_17169);
and UO_1301 (O_1301,N_15469,N_19514);
and UO_1302 (O_1302,N_17961,N_17676);
nor UO_1303 (O_1303,N_18601,N_15381);
and UO_1304 (O_1304,N_15201,N_18824);
or UO_1305 (O_1305,N_17352,N_15767);
nor UO_1306 (O_1306,N_15203,N_16686);
nand UO_1307 (O_1307,N_19017,N_16816);
nor UO_1308 (O_1308,N_18099,N_18056);
nor UO_1309 (O_1309,N_15331,N_17238);
nand UO_1310 (O_1310,N_17213,N_18666);
nor UO_1311 (O_1311,N_18219,N_16254);
or UO_1312 (O_1312,N_15146,N_18489);
nor UO_1313 (O_1313,N_15453,N_16517);
nand UO_1314 (O_1314,N_18104,N_19439);
or UO_1315 (O_1315,N_18955,N_18475);
nor UO_1316 (O_1316,N_19737,N_18135);
or UO_1317 (O_1317,N_18023,N_19307);
and UO_1318 (O_1318,N_16861,N_18183);
and UO_1319 (O_1319,N_19244,N_16402);
nand UO_1320 (O_1320,N_17358,N_15804);
xnor UO_1321 (O_1321,N_17452,N_15847);
and UO_1322 (O_1322,N_17691,N_18102);
or UO_1323 (O_1323,N_16641,N_18321);
or UO_1324 (O_1324,N_19556,N_16771);
nor UO_1325 (O_1325,N_16558,N_17531);
and UO_1326 (O_1326,N_16640,N_17329);
or UO_1327 (O_1327,N_18018,N_15055);
nand UO_1328 (O_1328,N_15365,N_16887);
or UO_1329 (O_1329,N_15740,N_19242);
nor UO_1330 (O_1330,N_15289,N_16440);
and UO_1331 (O_1331,N_17543,N_18631);
nand UO_1332 (O_1332,N_15024,N_18172);
and UO_1333 (O_1333,N_16571,N_16497);
and UO_1334 (O_1334,N_17618,N_17191);
and UO_1335 (O_1335,N_18292,N_15927);
nor UO_1336 (O_1336,N_18152,N_17256);
or UO_1337 (O_1337,N_18958,N_19925);
xnor UO_1338 (O_1338,N_15220,N_15684);
nand UO_1339 (O_1339,N_19781,N_19184);
nand UO_1340 (O_1340,N_17069,N_16381);
nand UO_1341 (O_1341,N_17247,N_15426);
nand UO_1342 (O_1342,N_18201,N_19591);
and UO_1343 (O_1343,N_15480,N_18856);
nand UO_1344 (O_1344,N_15795,N_16633);
xnor UO_1345 (O_1345,N_16021,N_18658);
nor UO_1346 (O_1346,N_15042,N_18822);
nor UO_1347 (O_1347,N_15126,N_15051);
nand UO_1348 (O_1348,N_19679,N_17457);
nor UO_1349 (O_1349,N_15372,N_15625);
nor UO_1350 (O_1350,N_18520,N_17821);
nor UO_1351 (O_1351,N_19994,N_17654);
xnor UO_1352 (O_1352,N_18066,N_16388);
nand UO_1353 (O_1353,N_19153,N_16780);
nor UO_1354 (O_1354,N_15495,N_15197);
and UO_1355 (O_1355,N_17649,N_16678);
nand UO_1356 (O_1356,N_17952,N_17866);
xnor UO_1357 (O_1357,N_19014,N_19388);
nor UO_1358 (O_1358,N_18190,N_19835);
or UO_1359 (O_1359,N_19565,N_15359);
and UO_1360 (O_1360,N_16563,N_18627);
xnor UO_1361 (O_1361,N_15032,N_18644);
nor UO_1362 (O_1362,N_17545,N_18006);
and UO_1363 (O_1363,N_18476,N_17359);
nand UO_1364 (O_1364,N_16526,N_15858);
or UO_1365 (O_1365,N_15333,N_18496);
and UO_1366 (O_1366,N_19563,N_15307);
or UO_1367 (O_1367,N_18952,N_19147);
nand UO_1368 (O_1368,N_16449,N_19344);
or UO_1369 (O_1369,N_17549,N_19020);
or UO_1370 (O_1370,N_16867,N_18368);
and UO_1371 (O_1371,N_18017,N_15252);
or UO_1372 (O_1372,N_16997,N_15650);
and UO_1373 (O_1373,N_15578,N_19814);
xor UO_1374 (O_1374,N_17692,N_17959);
or UO_1375 (O_1375,N_17812,N_15908);
nand UO_1376 (O_1376,N_17708,N_15896);
nand UO_1377 (O_1377,N_19841,N_17430);
nor UO_1378 (O_1378,N_15093,N_17187);
and UO_1379 (O_1379,N_19903,N_15911);
xor UO_1380 (O_1380,N_18032,N_16953);
nor UO_1381 (O_1381,N_17376,N_15360);
xnor UO_1382 (O_1382,N_18580,N_15718);
or UO_1383 (O_1383,N_19547,N_15545);
or UO_1384 (O_1384,N_16049,N_18819);
xor UO_1385 (O_1385,N_18239,N_15659);
and UO_1386 (O_1386,N_19470,N_18724);
and UO_1387 (O_1387,N_17101,N_18675);
or UO_1388 (O_1388,N_19897,N_16557);
nor UO_1389 (O_1389,N_16548,N_18400);
or UO_1390 (O_1390,N_15350,N_19875);
and UO_1391 (O_1391,N_15027,N_19860);
and UO_1392 (O_1392,N_18366,N_15999);
or UO_1393 (O_1393,N_19978,N_15486);
xnor UO_1394 (O_1394,N_17872,N_18659);
and UO_1395 (O_1395,N_19161,N_18046);
or UO_1396 (O_1396,N_19051,N_15131);
or UO_1397 (O_1397,N_19984,N_18310);
or UO_1398 (O_1398,N_17674,N_17924);
and UO_1399 (O_1399,N_19743,N_16879);
nand UO_1400 (O_1400,N_17997,N_15826);
nor UO_1401 (O_1401,N_16739,N_19753);
nor UO_1402 (O_1402,N_16378,N_15651);
or UO_1403 (O_1403,N_18541,N_17725);
nor UO_1404 (O_1404,N_17644,N_19871);
and UO_1405 (O_1405,N_18681,N_19535);
nand UO_1406 (O_1406,N_16414,N_15278);
nor UO_1407 (O_1407,N_18560,N_17340);
nand UO_1408 (O_1408,N_15389,N_19243);
or UO_1409 (O_1409,N_16251,N_16905);
and UO_1410 (O_1410,N_16860,N_17074);
nor UO_1411 (O_1411,N_17721,N_16881);
or UO_1412 (O_1412,N_17033,N_18837);
or UO_1413 (O_1413,N_15021,N_19372);
or UO_1414 (O_1414,N_17183,N_15603);
and UO_1415 (O_1415,N_15266,N_19582);
nand UO_1416 (O_1416,N_16322,N_18564);
or UO_1417 (O_1417,N_15026,N_16244);
nor UO_1418 (O_1418,N_19614,N_16656);
and UO_1419 (O_1419,N_19264,N_17437);
nor UO_1420 (O_1420,N_18622,N_17016);
xnor UO_1421 (O_1421,N_16023,N_19538);
nand UO_1422 (O_1422,N_16837,N_17154);
nand UO_1423 (O_1423,N_18577,N_16226);
and UO_1424 (O_1424,N_16104,N_16795);
nor UO_1425 (O_1425,N_15834,N_17042);
or UO_1426 (O_1426,N_19881,N_19466);
and UO_1427 (O_1427,N_16189,N_18606);
xnor UO_1428 (O_1428,N_19682,N_16972);
nor UO_1429 (O_1429,N_19937,N_17188);
or UO_1430 (O_1430,N_16864,N_16569);
nand UO_1431 (O_1431,N_19669,N_18869);
and UO_1432 (O_1432,N_17353,N_19168);
or UO_1433 (O_1433,N_17663,N_15171);
and UO_1434 (O_1434,N_19363,N_16386);
nand UO_1435 (O_1435,N_17581,N_15527);
or UO_1436 (O_1436,N_19818,N_19201);
nor UO_1437 (O_1437,N_18355,N_16809);
nand UO_1438 (O_1438,N_15194,N_19624);
or UO_1439 (O_1439,N_19462,N_15356);
or UO_1440 (O_1440,N_16054,N_17605);
and UO_1441 (O_1441,N_15728,N_18068);
and UO_1442 (O_1442,N_19825,N_16359);
or UO_1443 (O_1443,N_17066,N_17934);
nor UO_1444 (O_1444,N_16835,N_18583);
nor UO_1445 (O_1445,N_15217,N_16172);
xor UO_1446 (O_1446,N_15986,N_19724);
nand UO_1447 (O_1447,N_15700,N_17801);
or UO_1448 (O_1448,N_17651,N_18546);
or UO_1449 (O_1449,N_18626,N_17265);
nand UO_1450 (O_1450,N_16311,N_16465);
nand UO_1451 (O_1451,N_17529,N_19063);
nor UO_1452 (O_1452,N_15547,N_15677);
nand UO_1453 (O_1453,N_17831,N_18388);
nand UO_1454 (O_1454,N_15643,N_19996);
and UO_1455 (O_1455,N_15774,N_16502);
or UO_1456 (O_1456,N_18954,N_16393);
and UO_1457 (O_1457,N_16477,N_19353);
or UO_1458 (O_1458,N_15585,N_15163);
and UO_1459 (O_1459,N_18970,N_18349);
nor UO_1460 (O_1460,N_17473,N_19886);
nand UO_1461 (O_1461,N_18457,N_18686);
xnor UO_1462 (O_1462,N_18497,N_18286);
or UO_1463 (O_1463,N_17184,N_18370);
xor UO_1464 (O_1464,N_16573,N_15474);
nand UO_1465 (O_1465,N_17742,N_15889);
nand UO_1466 (O_1466,N_19460,N_15116);
or UO_1467 (O_1467,N_17514,N_15166);
xor UO_1468 (O_1468,N_16555,N_18247);
xnor UO_1469 (O_1469,N_16931,N_17469);
and UO_1470 (O_1470,N_19959,N_17475);
or UO_1471 (O_1471,N_16802,N_17237);
and UO_1472 (O_1472,N_19282,N_15416);
nor UO_1473 (O_1473,N_16016,N_19997);
or UO_1474 (O_1474,N_19040,N_16970);
nand UO_1475 (O_1475,N_16361,N_15693);
nand UO_1476 (O_1476,N_19236,N_16187);
and UO_1477 (O_1477,N_18197,N_18756);
nor UO_1478 (O_1478,N_17046,N_16707);
and UO_1479 (O_1479,N_19608,N_19007);
or UO_1480 (O_1480,N_18887,N_19077);
nor UO_1481 (O_1481,N_16219,N_16345);
nand UO_1482 (O_1482,N_15285,N_18660);
and UO_1483 (O_1483,N_16789,N_16224);
or UO_1484 (O_1484,N_19173,N_15932);
nor UO_1485 (O_1485,N_19585,N_18176);
nand UO_1486 (O_1486,N_18661,N_19136);
nand UO_1487 (O_1487,N_16013,N_15961);
and UO_1488 (O_1488,N_15321,N_17636);
nor UO_1489 (O_1489,N_19934,N_16056);
nor UO_1490 (O_1490,N_16639,N_15272);
nor UO_1491 (O_1491,N_19689,N_18977);
nand UO_1492 (O_1492,N_15674,N_17869);
and UO_1493 (O_1493,N_16175,N_18316);
nand UO_1494 (O_1494,N_17569,N_19951);
nor UO_1495 (O_1495,N_19782,N_17533);
nor UO_1496 (O_1496,N_19747,N_18430);
nand UO_1497 (O_1497,N_16626,N_19505);
and UO_1498 (O_1498,N_18036,N_18254);
or UO_1499 (O_1499,N_16303,N_16549);
nand UO_1500 (O_1500,N_16670,N_17175);
and UO_1501 (O_1501,N_19991,N_16407);
nor UO_1502 (O_1502,N_18514,N_19395);
and UO_1503 (O_1503,N_17648,N_18839);
xor UO_1504 (O_1504,N_16308,N_16237);
nand UO_1505 (O_1505,N_19341,N_15855);
nand UO_1506 (O_1506,N_17377,N_17181);
nor UO_1507 (O_1507,N_16501,N_15038);
or UO_1508 (O_1508,N_17981,N_16098);
xor UO_1509 (O_1509,N_17243,N_16342);
and UO_1510 (O_1510,N_15582,N_19195);
and UO_1511 (O_1511,N_17840,N_17239);
xnor UO_1512 (O_1512,N_15087,N_19678);
and UO_1513 (O_1513,N_15090,N_16950);
or UO_1514 (O_1514,N_15478,N_16445);
nor UO_1515 (O_1515,N_19343,N_15195);
or UO_1516 (O_1516,N_16264,N_15835);
nor UO_1517 (O_1517,N_15864,N_18870);
nor UO_1518 (O_1518,N_15313,N_15865);
and UO_1519 (O_1519,N_16923,N_15708);
and UO_1520 (O_1520,N_17270,N_19480);
and UO_1521 (O_1521,N_15524,N_19304);
and UO_1522 (O_1522,N_19355,N_16068);
and UO_1523 (O_1523,N_19187,N_17509);
and UO_1524 (O_1524,N_18999,N_15924);
nor UO_1525 (O_1525,N_15431,N_16840);
nor UO_1526 (O_1526,N_19078,N_17609);
and UO_1527 (O_1527,N_18548,N_15351);
xnor UO_1528 (O_1528,N_16708,N_17923);
nor UO_1529 (O_1529,N_18040,N_18397);
and UO_1530 (O_1530,N_16041,N_18309);
nor UO_1531 (O_1531,N_18409,N_15344);
nor UO_1532 (O_1532,N_16636,N_16706);
nor UO_1533 (O_1533,N_16882,N_16290);
nand UO_1534 (O_1534,N_15136,N_16613);
and UO_1535 (O_1535,N_19884,N_19378);
nor UO_1536 (O_1536,N_16365,N_19139);
or UO_1537 (O_1537,N_16866,N_17087);
and UO_1538 (O_1538,N_19155,N_17804);
nor UO_1539 (O_1539,N_17006,N_19774);
nand UO_1540 (O_1540,N_19844,N_18229);
nand UO_1541 (O_1541,N_19813,N_16198);
or UO_1542 (O_1542,N_19831,N_17018);
nand UO_1543 (O_1543,N_15473,N_15419);
or UO_1544 (O_1544,N_17291,N_19503);
nand UO_1545 (O_1545,N_17930,N_18589);
and UO_1546 (O_1546,N_19958,N_15698);
nor UO_1547 (O_1547,N_16963,N_17323);
nand UO_1548 (O_1548,N_19385,N_16701);
or UO_1549 (O_1549,N_16142,N_15243);
or UO_1550 (O_1550,N_18028,N_19289);
nand UO_1551 (O_1551,N_16688,N_17280);
xnor UO_1552 (O_1552,N_19755,N_15491);
xnor UO_1553 (O_1553,N_18471,N_17990);
nand UO_1554 (O_1554,N_15742,N_19098);
nand UO_1555 (O_1555,N_15906,N_17009);
or UO_1556 (O_1556,N_17782,N_17274);
nand UO_1557 (O_1557,N_18557,N_18568);
nand UO_1558 (O_1558,N_16899,N_18930);
and UO_1559 (O_1559,N_19727,N_19775);
or UO_1560 (O_1560,N_17305,N_18844);
nor UO_1561 (O_1561,N_17057,N_19667);
nor UO_1562 (O_1562,N_16368,N_19611);
nor UO_1563 (O_1563,N_16484,N_18994);
and UO_1564 (O_1564,N_17073,N_15635);
or UO_1565 (O_1565,N_16028,N_18327);
or UO_1566 (O_1566,N_18331,N_17246);
and UO_1567 (O_1567,N_17625,N_16510);
nor UO_1568 (O_1568,N_16334,N_18335);
nand UO_1569 (O_1569,N_18350,N_17827);
nand UO_1570 (O_1570,N_18597,N_18513);
or UO_1571 (O_1571,N_18619,N_17257);
nand UO_1572 (O_1572,N_16769,N_16043);
nor UO_1573 (O_1573,N_19411,N_15297);
and UO_1574 (O_1574,N_19436,N_18361);
nor UO_1575 (O_1575,N_15514,N_19668);
and UO_1576 (O_1576,N_18180,N_16075);
and UO_1577 (O_1577,N_17493,N_18943);
nor UO_1578 (O_1578,N_16405,N_15148);
and UO_1579 (O_1579,N_19008,N_18014);
nand UO_1580 (O_1580,N_19778,N_16415);
nor UO_1581 (O_1581,N_18800,N_19189);
nor UO_1582 (O_1582,N_16248,N_15660);
xnor UO_1583 (O_1583,N_15141,N_17986);
and UO_1584 (O_1584,N_16352,N_16081);
nor UO_1585 (O_1585,N_16358,N_17832);
nor UO_1586 (O_1586,N_18749,N_18417);
xnor UO_1587 (O_1587,N_19449,N_17624);
and UO_1588 (O_1588,N_16379,N_16539);
and UO_1589 (O_1589,N_15816,N_17536);
nand UO_1590 (O_1590,N_18151,N_18085);
xor UO_1591 (O_1591,N_17024,N_19352);
or UO_1592 (O_1592,N_16679,N_17541);
xnor UO_1593 (O_1593,N_16452,N_17994);
nand UO_1594 (O_1594,N_16203,N_17350);
and UO_1595 (O_1595,N_15279,N_18715);
nor UO_1596 (O_1596,N_16949,N_17317);
nand UO_1597 (O_1597,N_16201,N_18048);
and UO_1598 (O_1598,N_19308,N_16096);
or UO_1599 (O_1599,N_18058,N_15083);
and UO_1600 (O_1600,N_19589,N_17303);
and UO_1601 (O_1601,N_16974,N_16535);
or UO_1602 (O_1602,N_15817,N_17324);
nand UO_1603 (O_1603,N_17444,N_15218);
xor UO_1604 (O_1604,N_15209,N_19842);
and UO_1605 (O_1605,N_18878,N_16960);
or UO_1606 (O_1606,N_19545,N_16576);
nor UO_1607 (O_1607,N_18808,N_18556);
nor UO_1608 (O_1608,N_18312,N_17054);
or UO_1609 (O_1609,N_16703,N_18795);
nand UO_1610 (O_1610,N_19867,N_18921);
or UO_1611 (O_1611,N_17949,N_19823);
nor UO_1612 (O_1612,N_19572,N_18210);
nand UO_1613 (O_1613,N_19380,N_18511);
xor UO_1614 (O_1614,N_18092,N_16530);
nor UO_1615 (O_1615,N_15317,N_18670);
and UO_1616 (O_1616,N_19042,N_18030);
or UO_1617 (O_1617,N_18301,N_18393);
nand UO_1618 (O_1618,N_16712,N_16868);
and UO_1619 (O_1619,N_18122,N_15568);
or UO_1620 (O_1620,N_18578,N_17119);
or UO_1621 (O_1621,N_18969,N_17441);
nand UO_1622 (O_1622,N_15227,N_18777);
nor UO_1623 (O_1623,N_16039,N_16912);
nand UO_1624 (O_1624,N_19596,N_18378);
or UO_1625 (O_1625,N_19810,N_17914);
xor UO_1626 (O_1626,N_19580,N_18707);
xor UO_1627 (O_1627,N_18474,N_16996);
nand UO_1628 (O_1628,N_19392,N_15652);
or UO_1629 (O_1629,N_17633,N_16617);
nand UO_1630 (O_1630,N_16421,N_15151);
nor UO_1631 (O_1631,N_15785,N_17739);
or UO_1632 (O_1632,N_18033,N_19434);
and UO_1633 (O_1633,N_16473,N_16330);
and UO_1634 (O_1634,N_18912,N_15039);
nor UO_1635 (O_1635,N_18184,N_19969);
or UO_1636 (O_1636,N_15944,N_15079);
or UO_1637 (O_1637,N_17131,N_19647);
or UO_1638 (O_1638,N_18362,N_18956);
or UO_1639 (O_1639,N_18167,N_15234);
nand UO_1640 (O_1640,N_16722,N_16939);
or UO_1641 (O_1641,N_18555,N_17937);
and UO_1642 (O_1642,N_15856,N_15118);
nor UO_1643 (O_1643,N_16012,N_19962);
nand UO_1644 (O_1644,N_18984,N_16430);
nand UO_1645 (O_1645,N_16392,N_19708);
nor UO_1646 (O_1646,N_16257,N_19630);
nand UO_1647 (O_1647,N_17118,N_18260);
nor UO_1648 (O_1648,N_19581,N_16455);
or UO_1649 (O_1649,N_19799,N_18159);
or UO_1650 (O_1650,N_19213,N_18258);
nor UO_1651 (O_1651,N_19498,N_18065);
xor UO_1652 (O_1652,N_17144,N_19670);
nor UO_1653 (O_1653,N_19780,N_18375);
nand UO_1654 (O_1654,N_15202,N_19999);
xor UO_1655 (O_1655,N_15844,N_15101);
nor UO_1656 (O_1656,N_16669,N_17520);
nand UO_1657 (O_1657,N_18168,N_16161);
and UO_1658 (O_1658,N_19088,N_18966);
xnor UO_1659 (O_1659,N_17099,N_15089);
and UO_1660 (O_1660,N_16323,N_15761);
nor UO_1661 (O_1661,N_17052,N_19143);
and UO_1662 (O_1662,N_15639,N_15205);
xnor UO_1663 (O_1663,N_18885,N_18279);
and UO_1664 (O_1664,N_19266,N_16830);
nand UO_1665 (O_1665,N_18509,N_17479);
nand UO_1666 (O_1666,N_15281,N_19653);
and UO_1667 (O_1667,N_19762,N_16734);
and UO_1668 (O_1668,N_18025,N_18916);
or UO_1669 (O_1669,N_18633,N_18852);
nand UO_1670 (O_1670,N_17403,N_15713);
and UO_1671 (O_1671,N_16412,N_15824);
xnor UO_1672 (O_1672,N_18358,N_19629);
xor UO_1673 (O_1673,N_16904,N_15682);
nand UO_1674 (O_1674,N_17862,N_18914);
nor UO_1675 (O_1675,N_16748,N_16682);
nand UO_1676 (O_1676,N_16705,N_17258);
and UO_1677 (O_1677,N_19013,N_19575);
and UO_1678 (O_1678,N_17351,N_17906);
nor UO_1679 (O_1679,N_18682,N_18713);
nor UO_1680 (O_1680,N_16317,N_16842);
or UO_1681 (O_1681,N_15000,N_16301);
nor UO_1682 (O_1682,N_18836,N_18410);
nor UO_1683 (O_1683,N_16572,N_15248);
nand UO_1684 (O_1684,N_16474,N_15872);
nor UO_1685 (O_1685,N_19548,N_17586);
nor UO_1686 (O_1686,N_16108,N_19412);
nor UO_1687 (O_1687,N_19569,N_19970);
xnor UO_1688 (O_1688,N_17945,N_18103);
and UO_1689 (O_1689,N_17283,N_19798);
and UO_1690 (O_1690,N_15979,N_16207);
xor UO_1691 (O_1691,N_18898,N_15461);
and UO_1692 (O_1692,N_17614,N_16743);
nor UO_1693 (O_1693,N_18283,N_16564);
nand UO_1694 (O_1694,N_16353,N_15549);
or UO_1695 (O_1695,N_17711,N_16763);
nor UO_1696 (O_1696,N_19414,N_16988);
nor UO_1697 (O_1697,N_16964,N_15936);
or UO_1698 (O_1698,N_18251,N_17793);
nor UO_1699 (O_1699,N_18466,N_19564);
and UO_1700 (O_1700,N_15156,N_19149);
nor UO_1701 (O_1701,N_15314,N_17747);
or UO_1702 (O_1702,N_17084,N_16675);
and UO_1703 (O_1703,N_16695,N_19954);
nor UO_1704 (O_1704,N_19655,N_18980);
nand UO_1705 (O_1705,N_15945,N_19916);
or UO_1706 (O_1706,N_18426,N_16401);
nor UO_1707 (O_1707,N_18093,N_16032);
and UO_1708 (O_1708,N_19259,N_15690);
nor UO_1709 (O_1709,N_17477,N_18714);
or UO_1710 (O_1710,N_16767,N_16443);
or UO_1711 (O_1711,N_19771,N_19829);
and UO_1712 (O_1712,N_15876,N_19986);
nand UO_1713 (O_1713,N_19274,N_17956);
and UO_1714 (O_1714,N_17386,N_15516);
nor UO_1715 (O_1715,N_15730,N_18070);
or UO_1716 (O_1716,N_19058,N_15543);
nor UO_1717 (O_1717,N_16940,N_16529);
nor UO_1718 (O_1718,N_17842,N_17309);
and UO_1719 (O_1719,N_17162,N_19381);
and UO_1720 (O_1720,N_17171,N_17331);
xor UO_1721 (O_1721,N_19327,N_17918);
and UO_1722 (O_1722,N_15584,N_15075);
nor UO_1723 (O_1723,N_18215,N_16764);
nor UO_1724 (O_1724,N_16812,N_16627);
nand UO_1725 (O_1725,N_19374,N_15367);
nor UO_1726 (O_1726,N_18405,N_15870);
xnor UO_1727 (O_1727,N_18743,N_17443);
and UO_1728 (O_1728,N_17271,N_19795);
nor UO_1729 (O_1729,N_16944,N_16933);
or UO_1730 (O_1730,N_17498,N_15181);
nor UO_1731 (O_1731,N_19920,N_15575);
and UO_1732 (O_1732,N_16366,N_18566);
or UO_1733 (O_1733,N_18964,N_18117);
nand UO_1734 (O_1734,N_17022,N_16190);
nand UO_1735 (O_1735,N_16029,N_17755);
nor UO_1736 (O_1736,N_16246,N_18205);
nor UO_1737 (O_1737,N_19659,N_18699);
and UO_1738 (O_1738,N_16488,N_15460);
nand UO_1739 (O_1739,N_15077,N_15466);
nand UO_1740 (O_1740,N_19790,N_18071);
xor UO_1741 (O_1741,N_18486,N_16136);
nor UO_1742 (O_1742,N_16272,N_16932);
or UO_1743 (O_1743,N_15975,N_18603);
nand UO_1744 (O_1744,N_15047,N_17613);
and UO_1745 (O_1745,N_16856,N_17908);
or UO_1746 (O_1746,N_19658,N_16276);
nor UO_1747 (O_1747,N_18302,N_18246);
nand UO_1748 (O_1748,N_17835,N_16657);
nand UO_1749 (O_1749,N_15688,N_16732);
and UO_1750 (O_1750,N_16723,N_15347);
and UO_1751 (O_1751,N_15498,N_15563);
nor UO_1752 (O_1752,N_18945,N_17078);
xor UO_1753 (O_1753,N_16523,N_18550);
nor UO_1754 (O_1754,N_16294,N_17406);
nor UO_1755 (O_1755,N_15980,N_17873);
nor UO_1756 (O_1756,N_18791,N_19311);
and UO_1757 (O_1757,N_15697,N_19027);
and UO_1758 (O_1758,N_17091,N_16447);
nor UO_1759 (O_1759,N_18233,N_18918);
nand UO_1760 (O_1760,N_16468,N_17014);
nand UO_1761 (O_1761,N_18052,N_17922);
or UO_1762 (O_1762,N_19735,N_15577);
xnor UO_1763 (O_1763,N_15926,N_19638);
xor UO_1764 (O_1764,N_17670,N_18356);
xnor UO_1765 (O_1765,N_18832,N_17704);
nor UO_1766 (O_1766,N_19215,N_18611);
nor UO_1767 (O_1767,N_17632,N_18119);
or UO_1768 (O_1768,N_17284,N_19876);
xor UO_1769 (O_1769,N_15861,N_19046);
nand UO_1770 (O_1770,N_16658,N_17286);
nand UO_1771 (O_1771,N_17671,N_19802);
nand UO_1772 (O_1772,N_15792,N_19931);
nor UO_1773 (O_1773,N_18771,N_19087);
or UO_1774 (O_1774,N_16335,N_17552);
xor UO_1775 (O_1775,N_16660,N_15971);
or UO_1776 (O_1776,N_18920,N_19240);
xor UO_1777 (O_1777,N_15515,N_15222);
or UO_1778 (O_1778,N_18833,N_15160);
nor UO_1779 (O_1779,N_19963,N_17568);
nand UO_1780 (O_1780,N_15270,N_18596);
nor UO_1781 (O_1781,N_19805,N_17501);
and UO_1782 (O_1782,N_18790,N_16195);
xnor UO_1783 (O_1783,N_18181,N_18499);
nor UO_1784 (O_1784,N_16302,N_15132);
nor UO_1785 (O_1785,N_16814,N_17365);
or UO_1786 (O_1786,N_19178,N_18021);
xnor UO_1787 (O_1787,N_17787,N_16611);
nor UO_1788 (O_1788,N_17564,N_17267);
xnor UO_1789 (O_1789,N_18089,N_17002);
or UO_1790 (O_1790,N_16114,N_17532);
or UO_1791 (O_1791,N_17218,N_15496);
nor UO_1792 (O_1792,N_16907,N_17221);
or UO_1793 (O_1793,N_15271,N_16139);
and UO_1794 (O_1794,N_17028,N_15315);
or UO_1795 (O_1795,N_19172,N_16111);
and UO_1796 (O_1796,N_16891,N_19373);
nor UO_1797 (O_1797,N_17348,N_17276);
or UO_1798 (O_1798,N_16444,N_16296);
or UO_1799 (O_1799,N_15401,N_15420);
and UO_1800 (O_1800,N_16289,N_15368);
nand UO_1801 (O_1801,N_18816,N_15018);
nor UO_1802 (O_1802,N_17013,N_18164);
or UO_1803 (O_1803,N_19197,N_18891);
nor UO_1804 (O_1804,N_18592,N_19032);
and UO_1805 (O_1805,N_18850,N_15502);
xnor UO_1806 (O_1806,N_19656,N_16872);
or UO_1807 (O_1807,N_18614,N_18275);
and UO_1808 (O_1808,N_17168,N_18031);
and UO_1809 (O_1809,N_19122,N_17186);
or UO_1810 (O_1810,N_18645,N_16588);
and UO_1811 (O_1811,N_17346,N_16171);
nor UO_1812 (O_1812,N_18252,N_19112);
nand UO_1813 (O_1813,N_17562,N_15695);
nor UO_1814 (O_1814,N_15901,N_18845);
xor UO_1815 (O_1815,N_16897,N_19650);
nand UO_1816 (O_1816,N_15212,N_18861);
xnor UO_1817 (O_1817,N_15902,N_19239);
and UO_1818 (O_1818,N_18951,N_17030);
nor UO_1819 (O_1819,N_17917,N_15859);
xor UO_1820 (O_1820,N_17973,N_15726);
nand UO_1821 (O_1821,N_15251,N_15531);
xor UO_1822 (O_1822,N_17987,N_15303);
nor UO_1823 (O_1823,N_17944,N_16699);
or UO_1824 (O_1824,N_16870,N_18113);
or UO_1825 (O_1825,N_16409,N_17843);
or UO_1826 (O_1826,N_17599,N_18293);
nand UO_1827 (O_1827,N_15158,N_17385);
and UO_1828 (O_1828,N_15536,N_15318);
or UO_1829 (O_1829,N_18694,N_18907);
nor UO_1830 (O_1830,N_17815,N_18737);
xnor UO_1831 (O_1831,N_18343,N_19121);
or UO_1832 (O_1832,N_19704,N_16298);
nor UO_1833 (O_1833,N_18003,N_19338);
or UO_1834 (O_1834,N_15223,N_18664);
nor UO_1835 (O_1835,N_16267,N_15613);
or UO_1836 (O_1836,N_17476,N_15617);
or UO_1837 (O_1837,N_16552,N_17841);
nor UO_1838 (O_1838,N_15778,N_16718);
nor UO_1839 (O_1839,N_16223,N_15759);
nand UO_1840 (O_1840,N_16476,N_15261);
xnor UO_1841 (O_1841,N_15537,N_17155);
nor UO_1842 (O_1842,N_18041,N_16853);
and UO_1843 (O_1843,N_15914,N_18296);
nand UO_1844 (O_1844,N_18908,N_15452);
and UO_1845 (O_1845,N_15096,N_15404);
and UO_1846 (O_1846,N_17965,N_19491);
or UO_1847 (O_1847,N_15155,N_19429);
nand UO_1848 (O_1848,N_16832,N_18160);
xor UO_1849 (O_1849,N_19562,N_17921);
nor UO_1850 (O_1850,N_15408,N_15023);
nor UO_1851 (O_1851,N_16500,N_19926);
and UO_1852 (O_1852,N_15165,N_18438);
nor UO_1853 (O_1853,N_15773,N_16458);
and UO_1854 (O_1854,N_15871,N_18691);
nand UO_1855 (O_1855,N_16911,N_16463);
and UO_1856 (O_1856,N_17661,N_15647);
nand UO_1857 (O_1857,N_17880,N_17149);
and UO_1858 (O_1858,N_16080,N_19832);
nand UO_1859 (O_1859,N_17740,N_16205);
or UO_1860 (O_1860,N_18763,N_15925);
and UO_1861 (O_1861,N_15776,N_16720);
and UO_1862 (O_1862,N_15081,N_17957);
nand UO_1863 (O_1863,N_19205,N_19725);
or UO_1864 (O_1864,N_17426,N_19566);
nor UO_1865 (O_1865,N_17523,N_17813);
nor UO_1866 (O_1866,N_15929,N_17818);
and UO_1867 (O_1867,N_16031,N_18276);
nor UO_1868 (O_1868,N_15723,N_15983);
nand UO_1869 (O_1869,N_18381,N_19420);
and UO_1870 (O_1870,N_16990,N_17582);
xor UO_1871 (O_1871,N_16210,N_18698);
nand UO_1872 (O_1872,N_15794,N_15879);
or UO_1873 (O_1873,N_19188,N_18941);
and UO_1874 (O_1874,N_19073,N_18177);
xor UO_1875 (O_1875,N_18083,N_17940);
and UO_1876 (O_1876,N_17233,N_15207);
and UO_1877 (O_1877,N_15325,N_16554);
and UO_1878 (O_1878,N_16423,N_15819);
and UO_1879 (O_1879,N_19332,N_19939);
or UO_1880 (O_1880,N_19661,N_19787);
or UO_1881 (O_1881,N_15437,N_16153);
nand UO_1882 (O_1882,N_16078,N_16222);
and UO_1883 (O_1883,N_18235,N_18617);
nor UO_1884 (O_1884,N_15011,N_17012);
or UO_1885 (O_1885,N_18445,N_19649);
xnor UO_1886 (O_1886,N_15984,N_19235);
and UO_1887 (O_1887,N_19249,N_15758);
nand UO_1888 (O_1888,N_15298,N_15915);
nand UO_1889 (O_1889,N_16250,N_18455);
and UO_1890 (O_1890,N_15456,N_16255);
nor UO_1891 (O_1891,N_15380,N_15127);
or UO_1892 (O_1892,N_17462,N_15265);
and UO_1893 (O_1893,N_17683,N_15362);
nand UO_1894 (O_1894,N_17196,N_17431);
nand UO_1895 (O_1895,N_18346,N_15123);
and UO_1896 (O_1896,N_15139,N_19444);
and UO_1897 (O_1897,N_16220,N_16697);
or UO_1898 (O_1898,N_16089,N_17707);
xnor UO_1899 (O_1899,N_18562,N_18394);
nand UO_1900 (O_1900,N_17559,N_18265);
nand UO_1901 (O_1901,N_17969,N_15779);
and UO_1902 (O_1902,N_16309,N_19500);
xnor UO_1903 (O_1903,N_16174,N_18939);
nor UO_1904 (O_1904,N_15952,N_16875);
nor UO_1905 (O_1905,N_18300,N_16900);
and UO_1906 (O_1906,N_15851,N_19141);
nor UO_1907 (O_1907,N_15863,N_16612);
and UO_1908 (O_1908,N_19770,N_19357);
or UO_1909 (O_1909,N_17071,N_19837);
and UO_1910 (O_1910,N_15358,N_17460);
or UO_1911 (O_1911,N_17461,N_15736);
and UO_1912 (O_1912,N_18904,N_19126);
and UO_1913 (O_1913,N_18677,N_19843);
nor UO_1914 (O_1914,N_17259,N_19550);
and UO_1915 (O_1915,N_18473,N_17892);
or UO_1916 (O_1916,N_19594,N_15511);
and UO_1917 (O_1917,N_18639,N_15014);
and UO_1918 (O_1918,N_17170,N_16692);
and UO_1919 (O_1919,N_17072,N_18166);
nand UO_1920 (O_1920,N_19752,N_18886);
xnor UO_1921 (O_1921,N_18811,N_19001);
and UO_1922 (O_1922,N_19333,N_16509);
or UO_1923 (O_1923,N_19506,N_19909);
or UO_1924 (O_1924,N_18132,N_17743);
or UO_1925 (O_1925,N_16935,N_15529);
and UO_1926 (O_1926,N_18087,N_17368);
or UO_1927 (O_1927,N_18729,N_15057);
nand UO_1928 (O_1928,N_16027,N_16581);
or UO_1929 (O_1929,N_18391,N_16877);
nand UO_1930 (O_1930,N_16135,N_17401);
nor UO_1931 (O_1931,N_15970,N_17032);
nor UO_1932 (O_1932,N_19138,N_15598);
and UO_1933 (O_1933,N_17388,N_17120);
nand UO_1934 (O_1934,N_19039,N_18154);
nand UO_1935 (O_1935,N_19602,N_17838);
and UO_1936 (O_1936,N_19106,N_18044);
nor UO_1937 (O_1937,N_16834,N_17165);
or UO_1938 (O_1938,N_16969,N_16480);
and UO_1939 (O_1939,N_18255,N_16354);
nor UO_1940 (O_1940,N_15263,N_18108);
or UO_1941 (O_1941,N_18539,N_17641);
xor UO_1942 (O_1942,N_17448,N_18010);
nor UO_1943 (O_1943,N_15471,N_19872);
or UO_1944 (O_1944,N_15336,N_17953);
nor UO_1945 (O_1945,N_15631,N_16831);
nand UO_1946 (O_1946,N_17117,N_18876);
and UO_1947 (O_1947,N_15579,N_18315);
or UO_1948 (O_1948,N_18376,N_17311);
nand UO_1949 (O_1949,N_15213,N_17767);
or UO_1950 (O_1950,N_16432,N_18516);
nor UO_1951 (O_1951,N_18060,N_19971);
and UO_1952 (O_1952,N_19296,N_16927);
or UO_1953 (O_1953,N_19254,N_19483);
and UO_1954 (O_1954,N_19685,N_16625);
nor UO_1955 (O_1955,N_18192,N_15441);
and UO_1956 (O_1956,N_15614,N_17710);
xnor UO_1957 (O_1957,N_17774,N_17495);
xnor UO_1958 (O_1958,N_17886,N_19908);
and UO_1959 (O_1959,N_17526,N_17407);
nand UO_1960 (O_1960,N_18881,N_18741);
or UO_1961 (O_1961,N_19610,N_16129);
nand UO_1962 (O_1962,N_16478,N_16614);
nor UO_1963 (O_1963,N_18076,N_19845);
xor UO_1964 (O_1964,N_16635,N_16916);
nor UO_1965 (O_1965,N_15113,N_16883);
and UO_1966 (O_1966,N_19022,N_19567);
or UO_1967 (O_1967,N_15045,N_17090);
nand UO_1968 (O_1968,N_16253,N_18194);
and UO_1969 (O_1969,N_17595,N_15063);
nand UO_1970 (O_1970,N_18608,N_15692);
or UO_1971 (O_1971,N_18244,N_18703);
and UO_1972 (O_1972,N_19029,N_17701);
nand UO_1973 (O_1973,N_16776,N_17127);
nor UO_1974 (O_1974,N_19989,N_19684);
and UO_1975 (O_1975,N_15225,N_18847);
or UO_1976 (O_1976,N_16399,N_15787);
nand UO_1977 (O_1977,N_15346,N_19877);
nor UO_1978 (O_1978,N_18352,N_15976);
and UO_1979 (O_1979,N_15627,N_19559);
nand UO_1980 (O_1980,N_18480,N_16602);
nor UO_1981 (O_1981,N_15746,N_18558);
and UO_1982 (O_1982,N_15969,N_17504);
or UO_1983 (O_1983,N_16384,N_19726);
nand UO_1984 (O_1984,N_18783,N_16594);
nor UO_1985 (O_1985,N_15664,N_17293);
nand UO_1986 (O_1986,N_18150,N_18963);
nand UO_1987 (O_1987,N_15745,N_17420);
and UO_1988 (O_1988,N_15941,N_19717);
xnor UO_1989 (O_1989,N_19016,N_19553);
and UO_1990 (O_1990,N_18443,N_16578);
or UO_1991 (O_1991,N_17204,N_16030);
or UO_1992 (O_1992,N_17637,N_16591);
or UO_1993 (O_1993,N_18444,N_18893);
and UO_1994 (O_1994,N_19358,N_17919);
nand UO_1995 (O_1995,N_16046,N_19018);
nand UO_1996 (O_1996,N_16584,N_17897);
xor UO_1997 (O_1997,N_16481,N_19114);
nand UO_1998 (O_1998,N_15273,N_15991);
or UO_1999 (O_1999,N_17929,N_18505);
nor UO_2000 (O_2000,N_18134,N_19478);
nand UO_2001 (O_2001,N_16516,N_17335);
and UO_2002 (O_2002,N_18313,N_17991);
xor UO_2003 (O_2003,N_16200,N_18269);
and UO_2004 (O_2004,N_19490,N_17135);
nand UO_2005 (O_2005,N_15335,N_16721);
xnor UO_2006 (O_2006,N_18386,N_16045);
nand UO_2007 (O_2007,N_17865,N_18995);
and UO_2008 (O_2008,N_17205,N_18221);
nand UO_2009 (O_2009,N_19459,N_18487);
or UO_2010 (O_2010,N_17145,N_15648);
and UO_2011 (O_2011,N_17733,N_18243);
xor UO_2012 (O_2012,N_16982,N_17657);
and UO_2013 (O_2013,N_18390,N_18186);
or UO_2014 (O_2014,N_15597,N_18213);
nor UO_2015 (O_2015,N_18162,N_19394);
and UO_2016 (O_2016,N_19391,N_16087);
or UO_2017 (O_2017,N_16141,N_16943);
and UO_2018 (O_2018,N_19314,N_15747);
nor UO_2019 (O_2019,N_18605,N_18655);
xnor UO_2020 (O_2020,N_19062,N_17364);
nor UO_2021 (O_2021,N_17044,N_18552);
and UO_2022 (O_2022,N_19977,N_15447);
and UO_2023 (O_2023,N_15522,N_19334);
nor UO_2024 (O_2024,N_15186,N_15172);
and UO_2025 (O_2025,N_17080,N_17567);
nor UO_2026 (O_2026,N_19055,N_17394);
xnor UO_2027 (O_2027,N_15558,N_15097);
xnor UO_2028 (O_2028,N_19697,N_15574);
nor UO_2029 (O_2029,N_15556,N_16858);
or UO_2030 (O_2030,N_17912,N_17344);
or UO_2031 (O_2031,N_18727,N_17792);
and UO_2032 (O_2032,N_15109,N_16649);
nor UO_2033 (O_2033,N_18814,N_17342);
nor UO_2034 (O_2034,N_18371,N_19622);
nand UO_2035 (O_2035,N_16385,N_16498);
or UO_2036 (O_2036,N_15415,N_18250);
and UO_2037 (O_2037,N_19883,N_16938);
nand UO_2038 (O_2038,N_16332,N_16062);
nor UO_2039 (O_2039,N_19045,N_19619);
xnor UO_2040 (O_2040,N_18020,N_18873);
or UO_2041 (O_2041,N_15562,N_17098);
or UO_2042 (O_2042,N_17478,N_17524);
xor UO_2043 (O_2043,N_18915,N_16829);
nand UO_2044 (O_2044,N_18240,N_16761);
and UO_2045 (O_2045,N_15294,N_16337);
nand UO_2046 (O_2046,N_17399,N_17669);
nand UO_2047 (O_2047,N_16616,N_17722);
and UO_2048 (O_2048,N_18695,N_17055);
and UO_2049 (O_2049,N_18665,N_16305);
and UO_2050 (O_2050,N_17814,N_18257);
and UO_2051 (O_2051,N_16014,N_19179);
nand UO_2052 (O_2052,N_17227,N_18442);
or UO_2053 (O_2053,N_18100,N_19345);
or UO_2054 (O_2054,N_19607,N_19980);
nor UO_2055 (O_2055,N_15731,N_15122);
or UO_2056 (O_2056,N_17419,N_19520);
xnor UO_2057 (O_2057,N_17913,N_15434);
or UO_2058 (O_2058,N_16270,N_17383);
nor UO_2059 (O_2059,N_17777,N_19869);
nand UO_2060 (O_2060,N_19140,N_17626);
and UO_2061 (O_2061,N_17800,N_19788);
nor UO_2062 (O_2062,N_19613,N_16824);
nor UO_2063 (O_2063,N_19387,N_17911);
and UO_2064 (O_2064,N_16288,N_18494);
nor UO_2065 (O_2065,N_15287,N_18211);
and UO_2066 (O_2066,N_15454,N_19313);
and UO_2067 (O_2067,N_17433,N_19174);
nor UO_2068 (O_2068,N_15715,N_15338);
nor UO_2069 (O_2069,N_18042,N_19002);
and UO_2070 (O_2070,N_19632,N_16125);
xor UO_2071 (O_2071,N_16464,N_18853);
or UO_2072 (O_2072,N_19732,N_19117);
nand UO_2073 (O_2073,N_15764,N_19759);
and UO_2074 (O_2074,N_15860,N_16066);
xnor UO_2075 (O_2075,N_18237,N_18126);
or UO_2076 (O_2076,N_15821,N_19854);
nor UO_2077 (O_2077,N_18537,N_15411);
nor UO_2078 (O_2078,N_15540,N_16604);
or UO_2079 (O_2079,N_18535,N_15888);
xor UO_2080 (O_2080,N_15710,N_18988);
nor UO_2081 (O_2081,N_17505,N_15680);
and UO_2082 (O_2082,N_15472,N_18905);
nand UO_2083 (O_2083,N_16451,N_16127);
xor UO_2084 (O_2084,N_16862,N_15435);
nand UO_2085 (O_2085,N_17281,N_16600);
nor UO_2086 (O_2086,N_18403,N_17371);
nor UO_2087 (O_2087,N_18947,N_18910);
nand UO_2088 (O_2088,N_15681,N_15232);
or UO_2089 (O_2089,N_19097,N_15738);
nor UO_2090 (O_2090,N_16154,N_16279);
xor UO_2091 (O_2091,N_15477,N_19866);
nand UO_2092 (O_2092,N_17771,N_19198);
nand UO_2093 (O_2093,N_16196,N_17658);
and UO_2094 (O_2094,N_19546,N_16202);
and UO_2095 (O_2095,N_15414,N_17830);
xor UO_2096 (O_2096,N_19044,N_19981);
nor UO_2097 (O_2097,N_17680,N_19811);
nor UO_2098 (O_2098,N_15304,N_19224);
nand UO_2099 (O_2099,N_18971,N_15905);
and UO_2100 (O_2100,N_16093,N_19064);
or UO_2101 (O_2101,N_15878,N_16229);
and UO_2102 (O_2102,N_15277,N_18101);
nor UO_2103 (O_2103,N_16286,N_17699);
nor UO_2104 (O_2104,N_17059,N_19487);
nand UO_2105 (O_2105,N_15229,N_16713);
nand UO_2106 (O_2106,N_16351,N_18805);
nand UO_2107 (O_2107,N_18402,N_16467);
nand UO_2108 (O_2108,N_18054,N_15085);
and UO_2109 (O_2109,N_17110,N_15345);
or UO_2110 (O_2110,N_17192,N_16667);
nor UO_2111 (O_2111,N_19069,N_19955);
nor UO_2112 (O_2112,N_19709,N_19248);
nand UO_2113 (O_2113,N_17058,N_17507);
nand UO_2114 (O_2114,N_18088,N_17623);
xnor UO_2115 (O_2115,N_17296,N_16696);
nand UO_2116 (O_2116,N_15799,N_19786);
and UO_2117 (O_2117,N_16536,N_16400);
and UO_2118 (O_2118,N_19196,N_17322);
nand UO_2119 (O_2119,N_16406,N_17142);
and UO_2120 (O_2120,N_18421,N_17794);
nand UO_2121 (O_2121,N_16994,N_16119);
and UO_2122 (O_2122,N_16512,N_15916);
and UO_2123 (O_2123,N_16531,N_19208);
nand UO_2124 (O_2124,N_16439,N_16873);
or UO_2125 (O_2125,N_18667,N_16083);
nand UO_2126 (O_2126,N_16199,N_19110);
and UO_2127 (O_2127,N_15739,N_16485);
nand UO_2128 (O_2128,N_17901,N_19043);
and UO_2129 (O_2129,N_19913,N_15907);
or UO_2130 (O_2130,N_17224,N_19054);
xor UO_2131 (O_2131,N_18581,N_18612);
nor UO_2132 (O_2132,N_18616,N_19200);
or UO_2133 (O_2133,N_18755,N_17160);
nor UO_2134 (O_2134,N_18080,N_15555);
nor UO_2135 (O_2135,N_16886,N_18451);
and UO_2136 (O_2136,N_19756,N_18967);
nand UO_2137 (O_2137,N_18719,N_16259);
nor UO_2138 (O_2138,N_16372,N_19356);
nor UO_2139 (O_2139,N_16297,N_16527);
nor UO_2140 (O_2140,N_17373,N_19221);
nor UO_2141 (O_2141,N_16002,N_15198);
and UO_2142 (O_2142,N_15385,N_16383);
nor UO_2143 (O_2143,N_19654,N_17890);
nor UO_2144 (O_2144,N_18130,N_15280);
or UO_2145 (O_2145,N_19892,N_18563);
or UO_2146 (O_2146,N_19560,N_19852);
and UO_2147 (O_2147,N_16689,N_18838);
nand UO_2148 (O_2148,N_19070,N_15310);
and UO_2149 (O_2149,N_16329,N_17436);
and UO_2150 (O_2150,N_15455,N_16183);
or UO_2151 (O_2151,N_18899,N_15418);
nand UO_2152 (O_2152,N_16306,N_15387);
nor UO_2153 (O_2153,N_19229,N_17337);
nand UO_2154 (O_2154,N_19662,N_18384);
nand UO_2155 (O_2155,N_15943,N_19164);
or UO_2156 (O_2156,N_15104,N_16331);
nand UO_2157 (O_2157,N_18866,N_17525);
xnor UO_2158 (O_2158,N_15852,N_19100);
nor UO_2159 (O_2159,N_19976,N_15689);
or UO_2160 (O_2160,N_16880,N_18138);
and UO_2161 (O_2161,N_17357,N_18582);
or UO_2162 (O_2162,N_15630,N_17125);
nand UO_2163 (O_2163,N_19152,N_19907);
nand UO_2164 (O_2164,N_16192,N_18948);
and UO_2165 (O_2165,N_19132,N_16946);
xnor UO_2166 (O_2166,N_16547,N_17736);
nor UO_2167 (O_2167,N_16827,N_15777);
nor UO_2168 (O_2168,N_16170,N_19256);
nand UO_2169 (O_2169,N_16304,N_15354);
nand UO_2170 (O_2170,N_16100,N_16338);
nand UO_2171 (O_2171,N_17522,N_18701);
nand UO_2172 (O_2172,N_16609,N_17679);
and UO_2173 (O_2173,N_19144,N_16152);
nor UO_2174 (O_2174,N_19218,N_16800);
xnor UO_2175 (O_2175,N_15521,N_18917);
xor UO_2176 (O_2176,N_19644,N_18702);
or UO_2177 (O_2177,N_16817,N_16273);
nand UO_2178 (O_2178,N_17025,N_15735);
nand UO_2179 (O_2179,N_16716,N_17603);
and UO_2180 (O_2180,N_16589,N_17250);
and UO_2181 (O_2181,N_17223,N_19181);
nand UO_2182 (O_2182,N_15628,N_15152);
xor UO_2183 (O_2183,N_17189,N_18420);
xor UO_2184 (O_2184,N_19985,N_18944);
nor UO_2185 (O_2185,N_19760,N_18576);
xnor UO_2186 (O_2186,N_17666,N_19207);
xnor UO_2187 (O_2187,N_18620,N_17750);
and UO_2188 (O_2188,N_17229,N_19084);
nand UO_2189 (O_2189,N_19415,N_18901);
nand UO_2190 (O_2190,N_19030,N_17759);
or UO_2191 (O_2191,N_19368,N_15703);
and UO_2192 (O_2192,N_18097,N_19696);
or UO_2193 (O_2193,N_15802,N_19987);
and UO_2194 (O_2194,N_18672,N_15489);
and UO_2195 (O_2195,N_16737,N_15946);
or UO_2196 (O_2196,N_15771,N_15037);
nor UO_2197 (O_2197,N_17548,N_16019);
nand UO_2198 (O_2198,N_15519,N_15189);
and UO_2199 (O_2199,N_18408,N_19551);
nand UO_2200 (O_2200,N_19988,N_19318);
nor UO_2201 (O_2201,N_18416,N_15208);
or UO_2202 (O_2202,N_15756,N_17304);
and UO_2203 (O_2203,N_15610,N_19902);
and UO_2204 (O_2204,N_18561,N_19025);
xnor UO_2205 (O_2205,N_19921,N_16735);
nand UO_2206 (O_2206,N_16025,N_19276);
and UO_2207 (O_2207,N_18998,N_17334);
nand UO_2208 (O_2208,N_15646,N_18902);
or UO_2209 (O_2209,N_16747,N_15185);
xor UO_2210 (O_2210,N_15769,N_16499);
or UO_2211 (O_2211,N_16653,N_17242);
or UO_2212 (O_2212,N_15805,N_19783);
nor UO_2213 (O_2213,N_15216,N_15357);
nor UO_2214 (O_2214,N_19792,N_16610);
or UO_2215 (O_2215,N_15811,N_16733);
nand UO_2216 (O_2216,N_17159,N_18799);
nor UO_2217 (O_2217,N_17540,N_15873);
and UO_2218 (O_2218,N_17261,N_19300);
and UO_2219 (O_2219,N_18532,N_15535);
xor UO_2220 (O_2220,N_16037,N_15797);
or UO_2221 (O_2221,N_19540,N_19389);
nand UO_2222 (O_2222,N_19807,N_18270);
nor UO_2223 (O_2223,N_17888,N_17858);
nor UO_2224 (O_2224,N_19713,N_17458);
and UO_2225 (O_2225,N_17705,N_17185);
nor UO_2226 (O_2226,N_15095,N_17761);
xnor UO_2227 (O_2227,N_15552,N_19859);
and UO_2228 (O_2228,N_19645,N_17166);
nor UO_2229 (O_2229,N_17769,N_18185);
nand UO_2230 (O_2230,N_16955,N_17807);
xnor UO_2231 (O_2231,N_17421,N_16252);
nor UO_2232 (O_2232,N_16140,N_16819);
and UO_2233 (O_2233,N_15137,N_19561);
nand UO_2234 (O_2234,N_16902,N_15595);
or UO_2235 (O_2235,N_16815,N_18114);
nor UO_2236 (O_2236,N_15129,N_18610);
or UO_2237 (O_2237,N_15883,N_16216);
and UO_2238 (O_2238,N_16048,N_16417);
nand UO_2239 (O_2239,N_15070,N_18112);
nor UO_2240 (O_2240,N_15657,N_15443);
nand UO_2241 (O_2241,N_19691,N_18792);
or UO_2242 (O_2242,N_18094,N_17713);
nand UO_2243 (O_2243,N_16910,N_16238);
nand UO_2244 (O_2244,N_16339,N_16180);
nor UO_2245 (O_2245,N_16568,N_16785);
and UO_2246 (O_2246,N_15918,N_19328);
or UO_2247 (O_2247,N_19525,N_17244);
and UO_2248 (O_2248,N_15942,N_16983);
or UO_2249 (O_2249,N_16857,N_18586);
or UO_2250 (O_2250,N_16615,N_16567);
nand UO_2251 (O_2251,N_19947,N_16561);
and UO_2252 (O_2252,N_18536,N_16773);
xor UO_2253 (O_2253,N_18774,N_19096);
or UO_2254 (O_2254,N_17932,N_19287);
nor UO_2255 (O_2255,N_16346,N_19104);
nand UO_2256 (O_2256,N_16863,N_18862);
nand UO_2257 (O_2257,N_18992,N_17136);
xnor UO_2258 (O_2258,N_15379,N_15459);
nor UO_2259 (O_2259,N_19901,N_19041);
nor UO_2260 (O_2260,N_17194,N_16082);
nand UO_2261 (O_2261,N_19839,N_17021);
xor UO_2262 (O_2262,N_19722,N_18545);
nand UO_2263 (O_2263,N_15838,N_18016);
nor UO_2264 (O_2264,N_18079,N_18704);
or UO_2265 (O_2265,N_15634,N_17766);
nand UO_2266 (O_2266,N_18039,N_18828);
nor UO_2267 (O_2267,N_15476,N_17572);
nand UO_2268 (O_2268,N_16730,N_15162);
nor UO_2269 (O_2269,N_17982,N_16035);
and UO_2270 (O_2270,N_17050,N_17182);
and UO_2271 (O_2271,N_17984,N_15854);
or UO_2272 (O_2272,N_17695,N_18340);
or UO_2273 (O_2273,N_18453,N_19497);
and UO_2274 (O_2274,N_15167,N_19932);
nand UO_2275 (O_2275,N_19885,N_15649);
and UO_2276 (O_2276,N_17998,N_15538);
and UO_2277 (O_2277,N_17518,N_16976);
or UO_2278 (O_2278,N_16475,N_17349);
nand UO_2279 (O_2279,N_17410,N_19821);
or UO_2280 (O_2280,N_19675,N_16676);
nor UO_2281 (O_2281,N_15339,N_18128);
xor UO_2282 (O_2282,N_17315,N_17422);
xor UO_2283 (O_2283,N_18721,N_19257);
and UO_2284 (O_2284,N_18175,N_16518);
and UO_2285 (O_2285,N_17450,N_19214);
or UO_2286 (O_2286,N_17424,N_16044);
or UO_2287 (O_2287,N_18399,N_19873);
nand UO_2288 (O_2288,N_15390,N_16271);
nand UO_2289 (O_2289,N_18057,N_17053);
or UO_2290 (O_2290,N_16745,N_16822);
nand UO_2291 (O_2291,N_17588,N_19127);
and UO_2292 (O_2292,N_19517,N_16797);
nor UO_2293 (O_2293,N_15845,N_17083);
nand UO_2294 (O_2294,N_19745,N_15846);
and UO_2295 (O_2295,N_17355,N_18155);
nand UO_2296 (O_2296,N_18256,N_16185);
or UO_2297 (O_2297,N_17122,N_16662);
nand UO_2298 (O_2298,N_15602,N_17005);
and UO_2299 (O_2299,N_19879,N_15609);
nor UO_2300 (O_2300,N_17384,N_18857);
nor UO_2301 (O_2301,N_16144,N_16876);
nor UO_2302 (O_2302,N_19618,N_19237);
nand UO_2303 (O_2303,N_19597,N_19793);
nand UO_2304 (O_2304,N_17730,N_15640);
and UO_2305 (O_2305,N_18169,N_19120);
nand UO_2306 (O_2306,N_18628,N_18434);
and UO_2307 (O_2307,N_17542,N_17643);
and UO_2308 (O_2308,N_18490,N_19677);
nor UO_2309 (O_2309,N_17639,N_15757);
nor UO_2310 (O_2310,N_18738,N_16310);
nand UO_2311 (O_2311,N_17409,N_17810);
or UO_2312 (O_2312,N_16710,N_18766);
nor UO_2313 (O_2313,N_16637,N_17719);
xor UO_2314 (O_2314,N_16540,N_18643);
or UO_2315 (O_2315,N_18736,N_17808);
or UO_2316 (O_2316,N_19652,N_19326);
nand UO_2317 (O_2317,N_18571,N_16159);
nor UO_2318 (O_2318,N_18188,N_16989);
nor UO_2319 (O_2319,N_17333,N_15267);
or UO_2320 (O_2320,N_18693,N_18212);
xnor UO_2321 (O_2321,N_19306,N_15837);
nand UO_2322 (O_2322,N_19071,N_16687);
and UO_2323 (O_2323,N_18363,N_18688);
nand UO_2324 (O_2324,N_15125,N_19721);
nor UO_2325 (O_2325,N_17020,N_19734);
nor UO_2326 (O_2326,N_19354,N_15269);
or UO_2327 (O_2327,N_15830,N_17822);
nand UO_2328 (O_2328,N_17511,N_17558);
nand UO_2329 (O_2329,N_18329,N_17321);
and UO_2330 (O_2330,N_19512,N_18467);
nor UO_2331 (O_2331,N_15544,N_19990);
and UO_2332 (O_2332,N_19541,N_15221);
nand UO_2333 (O_2333,N_17786,N_16681);
nand UO_2334 (O_2334,N_19940,N_17780);
or UO_2335 (O_2335,N_17486,N_18864);
or UO_2336 (O_2336,N_16825,N_19599);
nor UO_2337 (O_2337,N_19617,N_16920);
or UO_2338 (O_2338,N_15366,N_18398);
nor UO_2339 (O_2339,N_19228,N_18158);
and UO_2340 (O_2340,N_16550,N_19488);
nor UO_2341 (O_2341,N_15493,N_18649);
nand UO_2342 (O_2342,N_19273,N_17612);
or UO_2343 (O_2343,N_18061,N_19474);
or UO_2344 (O_2344,N_17878,N_19731);
xnor UO_2345 (O_2345,N_15407,N_16234);
and UO_2346 (O_2346,N_16965,N_19952);
and UO_2347 (O_2347,N_16751,N_18825);
nor UO_2348 (O_2348,N_19275,N_16630);
or UO_2349 (O_2349,N_15082,N_18127);
nand UO_2350 (O_2350,N_15590,N_15987);
or UO_2351 (O_2351,N_15507,N_19957);
nor UO_2352 (O_2352,N_17490,N_17480);
nor UO_2353 (O_2353,N_18529,N_16833);
and UO_2354 (O_2354,N_16344,N_19364);
xor UO_2355 (O_2355,N_18187,N_19101);
nor UO_2356 (O_2356,N_19880,N_17361);
nand UO_2357 (O_2357,N_17269,N_15840);
nor UO_2358 (O_2358,N_17210,N_18759);
nor UO_2359 (O_2359,N_19620,N_19701);
nor UO_2360 (O_2360,N_17031,N_15068);
or UO_2361 (O_2361,N_19419,N_16314);
nor UO_2362 (O_2362,N_16340,N_18053);
xnor UO_2363 (O_2363,N_19246,N_15309);
nor UO_2364 (O_2364,N_18662,N_15711);
nor UO_2365 (O_2365,N_18261,N_15749);
nand UO_2366 (O_2366,N_17065,N_18414);
or UO_2367 (O_2367,N_19204,N_16959);
nand UO_2368 (O_2368,N_17301,N_19862);
xnor UO_2369 (O_2369,N_17811,N_15967);
and UO_2370 (O_2370,N_15061,N_15934);
and UO_2371 (O_2371,N_17570,N_17646);
or UO_2372 (O_2372,N_16434,N_17068);
nor UO_2373 (O_2373,N_19390,N_15177);
nor UO_2374 (O_2374,N_19681,N_15406);
and UO_2375 (O_2375,N_16162,N_15712);
and UO_2376 (O_2376,N_18433,N_17248);
and UO_2377 (O_2377,N_16410,N_17580);
xor UO_2378 (O_2378,N_18779,N_19081);
nor UO_2379 (O_2379,N_15948,N_15259);
nand UO_2380 (O_2380,N_15349,N_17327);
and UO_2381 (O_2381,N_15972,N_18484);
and UO_2382 (O_2382,N_19159,N_19603);
and UO_2383 (O_2383,N_18797,N_15352);
or UO_2384 (O_2384,N_15035,N_15257);
nor UO_2385 (O_2385,N_16579,N_19893);
nor UO_2386 (O_2386,N_16691,N_18305);
or UO_2387 (O_2387,N_17829,N_17220);
and UO_2388 (O_2388,N_19003,N_15653);
nand UO_2389 (O_2389,N_17723,N_18082);
nand UO_2390 (O_2390,N_16772,N_16283);
nand UO_2391 (O_2391,N_17950,N_18337);
xor UO_2392 (O_2392,N_19399,N_18734);
xnor UO_2393 (O_2393,N_15187,N_18804);
and UO_2394 (O_2394,N_15428,N_18011);
xnor UO_2395 (O_2395,N_15099,N_19154);
and UO_2396 (O_2396,N_18217,N_18325);
nand UO_2397 (O_2397,N_15388,N_19489);
or UO_2398 (O_2398,N_18926,N_15382);
or UO_2399 (O_2399,N_18689,N_16395);
nor UO_2400 (O_2400,N_19447,N_19426);
nor UO_2401 (O_2401,N_15215,N_18889);
and UO_2402 (O_2402,N_16937,N_16631);
nor UO_2403 (O_2403,N_18991,N_17620);
nor UO_2404 (O_2404,N_15632,N_15178);
or UO_2405 (O_2405,N_19286,N_18924);
nand UO_2406 (O_2406,N_18815,N_18938);
nand UO_2407 (O_2407,N_15260,N_15490);
and UO_2408 (O_2408,N_16147,N_16425);
or UO_2409 (O_2409,N_19135,N_15526);
nand UO_2410 (O_2410,N_19451,N_19012);
xor UO_2411 (O_2411,N_19302,N_17694);
nand UO_2412 (O_2412,N_19973,N_16260);
and UO_2413 (O_2413,N_15594,N_19424);
nor UO_2414 (O_2414,N_18746,N_18604);
and UO_2415 (O_2415,N_16590,N_18440);
nand UO_2416 (O_2416,N_17724,N_15341);
nand UO_2417 (O_2417,N_15233,N_18338);
nand UO_2418 (O_2418,N_19758,N_18145);
xnor UO_2419 (O_2419,N_17778,N_18553);
nor UO_2420 (O_2420,N_17900,N_18367);
nand UO_2421 (O_2421,N_17833,N_18696);
and UO_2422 (O_2422,N_16896,N_19403);
and UO_2423 (O_2423,N_16813,N_18418);
nor UO_2424 (O_2424,N_18290,N_15249);
nand UO_2425 (O_2425,N_17172,N_18851);
or UO_2426 (O_2426,N_17795,N_17434);
nor UO_2427 (O_2427,N_17485,N_17513);
nand UO_2428 (O_2428,N_19587,N_18174);
nand UO_2429 (O_2429,N_19324,N_18599);
and UO_2430 (O_2430,N_17484,N_18937);
nand UO_2431 (O_2431,N_15839,N_19595);
nor UO_2432 (O_2432,N_18879,N_17228);
and UO_2433 (O_2433,N_18326,N_19310);
or UO_2434 (O_2434,N_15060,N_18745);
nand UO_2435 (O_2435,N_19865,N_17715);
nand UO_2436 (O_2436,N_18810,N_15909);
or UO_2437 (O_2437,N_17697,N_18841);
nand UO_2438 (O_2438,N_18911,N_19377);
nor UO_2439 (O_2439,N_15571,N_16364);
or UO_2440 (O_2440,N_16123,N_16796);
nand UO_2441 (O_2441,N_17798,N_17102);
and UO_2442 (O_2442,N_17332,N_19552);
nor UO_2443 (O_2443,N_16841,N_17898);
xor UO_2444 (O_2444,N_16852,N_15002);
nor UO_2445 (O_2445,N_19531,N_15685);
nand UO_2446 (O_2446,N_19953,N_19361);
nor UO_2447 (O_2447,N_17817,N_15551);
nor UO_2448 (O_2448,N_19047,N_19749);
or UO_2449 (O_2449,N_19494,N_16507);
xnor UO_2450 (O_2450,N_18990,N_17143);
and UO_2451 (O_2451,N_18465,N_15031);
or UO_2452 (O_2452,N_19297,N_17720);
or UO_2453 (O_2453,N_16930,N_16892);
nor UO_2454 (O_2454,N_16759,N_19504);
nor UO_2455 (O_2455,N_17864,N_19258);
and UO_2456 (O_2456,N_17438,N_19660);
and UO_2457 (O_2457,N_17951,N_19340);
nor UO_2458 (O_2458,N_19521,N_18277);
nor UO_2459 (O_2459,N_15001,N_19295);
and UO_2460 (O_2460,N_19477,N_16262);
nand UO_2461 (O_2461,N_15219,N_16239);
or UO_2462 (O_2462,N_15704,N_15638);
or UO_2463 (O_2463,N_18222,N_15276);
and UO_2464 (O_2464,N_19754,N_16371);
xnor UO_2465 (O_2465,N_19053,N_19299);
and UO_2466 (O_2466,N_16810,N_16320);
and UO_2467 (O_2467,N_17824,N_19819);
nor UO_2468 (O_2468,N_18439,N_18110);
and UO_2469 (O_2469,N_17179,N_19366);
or UO_2470 (O_2470,N_17199,N_17681);
and UO_2471 (O_2471,N_16209,N_15299);
nand UO_2472 (O_2472,N_19502,N_17380);
and UO_2473 (O_2473,N_18624,N_18288);
and UO_2474 (O_2474,N_18299,N_19199);
and UO_2475 (O_2475,N_18767,N_19129);
xor UO_2476 (O_2476,N_17902,N_19528);
or UO_2477 (O_2477,N_15913,N_16487);
nor UO_2478 (O_2478,N_19574,N_16684);
xor UO_2479 (O_2479,N_16729,N_15291);
nor UO_2480 (O_2480,N_19851,N_17287);
or UO_2481 (O_2481,N_15235,N_16120);
nand UO_2482 (O_2482,N_15508,N_18077);
or UO_2483 (O_2483,N_17260,N_18812);
and UO_2484 (O_2484,N_18654,N_18909);
and UO_2485 (O_2485,N_15885,N_16685);
or UO_2486 (O_2486,N_18464,N_18206);
and UO_2487 (O_2487,N_18072,N_16768);
nor UO_2488 (O_2488,N_17173,N_17673);
nand UO_2489 (O_2489,N_16599,N_16149);
nand UO_2490 (O_2490,N_19706,N_17828);
nand UO_2491 (O_2491,N_19222,N_15572);
and UO_2492 (O_2492,N_15448,N_16585);
nor UO_2493 (O_2493,N_16287,N_19182);
or UO_2494 (O_2494,N_19992,N_15084);
and UO_2495 (O_2495,N_19666,N_15274);
and UO_2496 (O_2496,N_18705,N_18940);
nor UO_2497 (O_2497,N_16177,N_16740);
and UO_2498 (O_2498,N_17235,N_16917);
nand UO_2499 (O_2499,N_16998,N_15882);
endmodule