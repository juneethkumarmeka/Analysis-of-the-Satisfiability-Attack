module basic_1500_15000_2000_5_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1244,In_140);
or U1 (N_1,In_625,In_273);
nand U2 (N_2,In_703,In_370);
nor U3 (N_3,In_1427,In_1192);
or U4 (N_4,In_760,In_1477);
nand U5 (N_5,In_1292,In_1096);
and U6 (N_6,In_1127,In_838);
nand U7 (N_7,In_329,In_559);
nand U8 (N_8,In_157,In_875);
and U9 (N_9,In_1432,In_785);
nor U10 (N_10,In_340,In_1142);
or U11 (N_11,In_1396,In_474);
nand U12 (N_12,In_770,In_587);
nand U13 (N_13,In_17,In_1138);
nor U14 (N_14,In_1483,In_246);
or U15 (N_15,In_364,In_1023);
and U16 (N_16,In_965,In_634);
and U17 (N_17,In_926,In_1337);
nand U18 (N_18,In_1406,In_1106);
or U19 (N_19,In_549,In_462);
or U20 (N_20,In_1336,In_818);
nand U21 (N_21,In_59,In_1391);
nand U22 (N_22,In_663,In_920);
and U23 (N_23,In_1319,In_829);
nand U24 (N_24,In_162,In_1462);
or U25 (N_25,In_626,In_1144);
or U26 (N_26,In_1001,In_566);
or U27 (N_27,In_1496,In_1368);
nand U28 (N_28,In_1194,In_632);
and U29 (N_29,In_48,In_379);
nand U30 (N_30,In_1331,In_235);
nand U31 (N_31,In_1407,In_1400);
or U32 (N_32,In_790,In_1321);
and U33 (N_33,In_660,In_70);
and U34 (N_34,In_1480,In_1146);
nand U35 (N_35,In_464,In_957);
or U36 (N_36,In_1344,In_247);
nand U37 (N_37,In_153,In_1049);
nand U38 (N_38,In_1343,In_569);
nand U39 (N_39,In_1470,In_65);
and U40 (N_40,In_20,In_1082);
nand U41 (N_41,In_540,In_1205);
nor U42 (N_42,In_548,In_145);
nand U43 (N_43,In_557,In_582);
and U44 (N_44,In_114,In_131);
or U45 (N_45,In_953,In_414);
and U46 (N_46,In_1151,In_620);
nand U47 (N_47,In_775,In_107);
nand U48 (N_48,In_1035,In_1311);
or U49 (N_49,In_1453,In_682);
or U50 (N_50,In_215,In_1257);
xnor U51 (N_51,In_46,In_1017);
nand U52 (N_52,In_923,In_482);
and U53 (N_53,In_1000,In_191);
nand U54 (N_54,In_542,In_174);
nand U55 (N_55,In_1121,In_1447);
nor U56 (N_56,In_441,In_948);
nor U57 (N_57,In_1497,In_214);
nand U58 (N_58,In_445,In_997);
nor U59 (N_59,In_406,In_182);
nand U60 (N_60,In_1412,In_1430);
nand U61 (N_61,In_617,In_350);
or U62 (N_62,In_74,In_1189);
nand U63 (N_63,In_10,In_1067);
nand U64 (N_64,In_264,In_1043);
and U65 (N_65,In_972,In_1449);
or U66 (N_66,In_1282,In_995);
nand U67 (N_67,In_1476,In_431);
nor U68 (N_68,In_76,In_1044);
nand U69 (N_69,In_801,In_561);
or U70 (N_70,In_584,In_1385);
nand U71 (N_71,In_26,In_283);
and U72 (N_72,In_1392,In_1165);
and U73 (N_73,In_45,In_423);
and U74 (N_74,In_152,In_1223);
and U75 (N_75,In_978,In_1098);
nand U76 (N_76,In_761,In_156);
and U77 (N_77,In_281,In_15);
nor U78 (N_78,In_1107,In_846);
and U79 (N_79,In_865,In_927);
nor U80 (N_80,In_498,In_823);
and U81 (N_81,In_764,In_41);
nand U82 (N_82,In_507,In_435);
nor U83 (N_83,In_976,In_359);
nor U84 (N_84,In_432,In_677);
nand U85 (N_85,In_741,In_1084);
nand U86 (N_86,In_1118,In_808);
nand U87 (N_87,In_735,In_242);
or U88 (N_88,In_515,In_510);
nor U89 (N_89,In_892,In_766);
nor U90 (N_90,In_335,In_803);
or U91 (N_91,In_492,In_1443);
nand U92 (N_92,In_1079,In_470);
nand U93 (N_93,In_240,In_594);
or U94 (N_94,In_394,In_461);
or U95 (N_95,In_1214,In_168);
and U96 (N_96,In_637,In_1195);
nand U97 (N_97,In_552,In_781);
or U98 (N_98,In_843,In_252);
nand U99 (N_99,In_155,In_720);
xnor U100 (N_100,In_1314,In_993);
or U101 (N_101,In_1366,In_579);
or U102 (N_102,In_1128,In_1081);
and U103 (N_103,In_1372,In_97);
or U104 (N_104,In_630,In_751);
and U105 (N_105,In_377,In_177);
nand U106 (N_106,In_1033,In_138);
nor U107 (N_107,In_125,In_527);
and U108 (N_108,In_1188,In_472);
or U109 (N_109,In_583,In_1219);
nor U110 (N_110,In_621,In_344);
nand U111 (N_111,In_1293,In_66);
or U112 (N_112,In_1078,In_1089);
nand U113 (N_113,In_239,In_1168);
or U114 (N_114,In_267,In_53);
nor U115 (N_115,In_1277,In_1123);
nand U116 (N_116,In_1409,In_1494);
nor U117 (N_117,In_1454,In_907);
and U118 (N_118,In_698,In_1021);
nand U119 (N_119,In_79,In_777);
nand U120 (N_120,In_811,In_969);
and U121 (N_121,In_317,In_25);
or U122 (N_122,In_649,In_124);
or U123 (N_123,In_732,In_608);
nor U124 (N_124,In_736,In_1467);
nand U125 (N_125,In_1299,In_947);
and U126 (N_126,In_639,In_830);
or U127 (N_127,In_1080,In_1369);
nor U128 (N_128,In_734,In_874);
or U129 (N_129,In_565,In_506);
or U130 (N_130,In_450,In_1110);
nand U131 (N_131,In_1442,In_1275);
nor U132 (N_132,In_1008,In_398);
nand U133 (N_133,In_1458,In_1298);
or U134 (N_134,In_648,In_1408);
and U135 (N_135,In_509,In_110);
nor U136 (N_136,In_1295,In_1281);
or U137 (N_137,In_746,In_918);
or U138 (N_138,In_855,In_303);
nand U139 (N_139,In_1358,In_788);
or U140 (N_140,In_1472,In_1076);
nand U141 (N_141,In_712,In_1308);
nand U142 (N_142,In_1426,In_1147);
or U143 (N_143,In_816,In_603);
and U144 (N_144,In_289,In_849);
nor U145 (N_145,In_418,In_684);
and U146 (N_146,In_337,In_109);
nand U147 (N_147,In_1237,In_1352);
or U148 (N_148,In_361,In_609);
nand U149 (N_149,In_478,In_690);
or U150 (N_150,In_1290,In_352);
and U151 (N_151,In_574,In_8);
or U152 (N_152,In_1285,In_1353);
nand U153 (N_153,In_1065,In_845);
and U154 (N_154,In_867,In_1243);
xnor U155 (N_155,In_494,In_1161);
nor U156 (N_156,In_178,In_456);
nor U157 (N_157,In_80,In_419);
or U158 (N_158,In_962,In_534);
nor U159 (N_159,In_334,In_1357);
or U160 (N_160,In_659,In_102);
or U161 (N_161,In_296,In_1163);
xnor U162 (N_162,In_34,In_1029);
and U163 (N_163,In_1238,In_840);
and U164 (N_164,In_1446,In_979);
nand U165 (N_165,In_1016,In_558);
or U166 (N_166,In_413,In_310);
nor U167 (N_167,In_1464,In_856);
and U168 (N_168,In_688,In_287);
nand U169 (N_169,In_1039,In_237);
or U170 (N_170,In_1239,In_1274);
or U171 (N_171,In_1156,In_985);
and U172 (N_172,In_694,In_248);
or U173 (N_173,In_717,In_657);
nor U174 (N_174,In_827,In_297);
nor U175 (N_175,In_1030,In_1145);
and U176 (N_176,In_1071,In_835);
nor U177 (N_177,In_290,In_475);
and U178 (N_178,In_1388,In_384);
and U179 (N_179,In_349,In_1095);
nand U180 (N_180,In_755,In_195);
or U181 (N_181,In_1278,In_817);
and U182 (N_182,In_47,In_716);
or U183 (N_183,In_424,In_750);
nor U184 (N_184,In_1347,In_1460);
nand U185 (N_185,In_51,In_1059);
or U186 (N_186,In_1171,In_1421);
nor U187 (N_187,In_535,In_459);
and U188 (N_188,In_1487,In_792);
or U189 (N_189,In_245,In_932);
nand U190 (N_190,In_911,In_1124);
or U191 (N_191,In_1379,In_1428);
and U192 (N_192,In_854,In_83);
and U193 (N_193,In_1191,In_1270);
and U194 (N_194,In_1361,In_1068);
and U195 (N_195,In_573,In_338);
and U196 (N_196,In_436,In_315);
and U197 (N_197,In_299,In_873);
and U198 (N_198,In_1228,In_841);
or U199 (N_199,In_1032,In_385);
nor U200 (N_200,In_1088,In_1466);
and U201 (N_201,In_1286,In_263);
and U202 (N_202,In_63,In_726);
nor U203 (N_203,In_1420,In_1053);
or U204 (N_204,In_1212,In_699);
nor U205 (N_205,In_1122,In_165);
and U206 (N_206,In_119,In_33);
nand U207 (N_207,In_1309,In_483);
or U208 (N_208,In_1003,In_1063);
or U209 (N_209,In_493,In_199);
nor U210 (N_210,In_807,In_1069);
xor U211 (N_211,In_139,In_987);
nor U212 (N_212,In_782,In_783);
or U213 (N_213,In_280,In_421);
and U214 (N_214,In_925,In_171);
or U215 (N_215,In_1418,In_5);
and U216 (N_216,In_137,In_207);
and U217 (N_217,In_941,In_689);
nor U218 (N_218,In_958,In_67);
nor U219 (N_219,In_345,In_3);
and U220 (N_220,In_251,In_222);
or U221 (N_221,In_667,In_219);
nor U222 (N_222,In_541,In_1026);
nand U223 (N_223,In_860,In_990);
or U224 (N_224,In_791,In_484);
and U225 (N_225,In_402,In_1092);
and U226 (N_226,In_727,In_757);
nand U227 (N_227,In_148,In_709);
or U228 (N_228,In_1208,In_1249);
xor U229 (N_229,In_1135,In_497);
xor U230 (N_230,In_1450,In_1116);
and U231 (N_231,In_311,In_1230);
and U232 (N_232,In_982,In_906);
and U233 (N_233,In_598,In_576);
or U234 (N_234,In_1207,In_651);
nand U235 (N_235,In_44,In_244);
nand U236 (N_236,In_342,In_1371);
or U237 (N_237,In_208,In_82);
and U238 (N_238,In_848,In_730);
nand U239 (N_239,In_852,In_1499);
and U240 (N_240,In_1104,In_1370);
and U241 (N_241,In_1186,In_1258);
or U242 (N_242,In_917,In_1306);
nor U243 (N_243,In_1355,In_711);
and U244 (N_244,In_1444,In_108);
nor U245 (N_245,In_1136,In_793);
nand U246 (N_246,In_1119,In_453);
nor U247 (N_247,In_1125,In_446);
and U248 (N_248,In_449,In_241);
nand U249 (N_249,In_704,In_183);
nand U250 (N_250,In_1280,In_1055);
or U251 (N_251,In_553,In_1302);
and U252 (N_252,In_1229,In_200);
nand U253 (N_253,In_405,In_522);
nand U254 (N_254,In_1325,In_973);
nand U255 (N_255,In_502,In_942);
or U256 (N_256,In_1326,In_547);
nor U257 (N_257,In_756,In_1060);
xnor U258 (N_258,In_851,In_890);
nand U259 (N_259,In_546,In_585);
nand U260 (N_260,In_1172,In_984);
or U261 (N_261,In_1226,In_771);
or U262 (N_262,In_706,In_2);
and U263 (N_263,In_479,In_601);
nand U264 (N_264,In_596,In_1187);
and U265 (N_265,In_1149,In_588);
nand U266 (N_266,In_1108,In_1140);
or U267 (N_267,In_1201,In_320);
nor U268 (N_268,In_1231,In_224);
and U269 (N_269,In_433,In_1261);
nand U270 (N_270,In_531,In_964);
or U271 (N_271,In_939,In_1221);
nand U272 (N_272,In_321,In_440);
nand U273 (N_273,In_123,In_1087);
nor U274 (N_274,In_1439,In_213);
nand U275 (N_275,In_1091,In_1236);
nand U276 (N_276,In_779,In_210);
or U277 (N_277,In_480,In_1143);
nand U278 (N_278,In_575,In_900);
and U279 (N_279,In_197,In_810);
nor U280 (N_280,In_358,In_988);
nor U281 (N_281,In_1036,In_416);
nor U282 (N_282,In_710,In_271);
and U283 (N_283,In_1455,In_1024);
nor U284 (N_284,In_314,In_186);
nor U285 (N_285,In_1064,In_227);
nand U286 (N_286,In_868,In_190);
nor U287 (N_287,In_1083,In_1377);
or U288 (N_288,In_323,In_209);
or U289 (N_289,In_989,In_908);
nor U290 (N_290,In_412,In_913);
and U291 (N_291,In_1493,In_1410);
or U292 (N_292,In_1378,In_376);
nor U293 (N_293,In_28,In_738);
and U294 (N_294,In_1490,In_1090);
nand U295 (N_295,In_1247,In_160);
nor U296 (N_296,In_1203,In_580);
or U297 (N_297,In_869,In_217);
nor U298 (N_298,In_254,In_1101);
or U299 (N_299,In_877,In_753);
nand U300 (N_300,In_1062,In_929);
and U301 (N_301,In_1154,In_255);
nor U302 (N_302,In_13,In_826);
nand U303 (N_303,In_11,In_312);
and U304 (N_304,In_586,In_170);
nand U305 (N_305,In_1041,In_175);
nor U306 (N_306,In_452,In_477);
xnor U307 (N_307,In_1332,In_357);
nand U308 (N_308,In_1485,In_154);
and U309 (N_309,In_1004,In_455);
nand U310 (N_310,In_1448,In_1072);
or U311 (N_311,In_1322,In_212);
nand U312 (N_312,In_686,In_680);
or U313 (N_313,In_1429,In_327);
nor U314 (N_314,In_1375,In_591);
and U315 (N_315,In_322,In_1491);
and U316 (N_316,In_332,In_266);
and U317 (N_317,In_1384,In_1437);
nand U318 (N_318,In_517,In_759);
nand U319 (N_319,In_556,In_970);
or U320 (N_320,In_37,In_539);
nand U321 (N_321,In_318,In_871);
nor U322 (N_322,In_391,In_991);
or U323 (N_323,In_1038,In_380);
nand U324 (N_324,In_604,In_1100);
and U325 (N_325,In_476,In_974);
nor U326 (N_326,In_16,In_1181);
and U327 (N_327,In_328,In_491);
or U328 (N_328,In_86,In_912);
or U329 (N_329,In_950,In_1196);
and U330 (N_330,In_1027,In_279);
nand U331 (N_331,In_363,In_971);
nor U332 (N_332,In_19,In_1020);
nand U333 (N_333,In_1218,In_1433);
nand U334 (N_334,In_687,In_545);
nor U335 (N_335,In_98,In_645);
nand U336 (N_336,In_928,In_1009);
and U337 (N_337,In_487,In_762);
or U338 (N_338,In_383,In_1114);
nand U339 (N_339,In_220,In_812);
or U340 (N_340,In_692,In_886);
or U341 (N_341,In_831,In_1276);
and U342 (N_342,In_1289,In_967);
nor U343 (N_343,In_62,In_1253);
nand U344 (N_344,In_1052,In_146);
nor U345 (N_345,In_1198,In_748);
nand U346 (N_346,In_1073,In_371);
or U347 (N_347,In_336,In_1362);
nand U348 (N_348,In_615,In_650);
or U349 (N_349,In_4,In_503);
or U350 (N_350,In_909,In_1394);
nand U351 (N_351,In_326,In_232);
nand U352 (N_352,In_1297,In_981);
nor U353 (N_353,In_613,In_744);
nor U354 (N_354,In_1050,In_616);
nand U355 (N_355,In_1441,In_422);
and U356 (N_356,In_729,In_367);
nor U357 (N_357,In_333,In_1048);
nor U358 (N_358,In_919,In_1227);
and U359 (N_359,In_270,In_1303);
or U360 (N_360,In_1498,In_1338);
and U361 (N_361,In_43,In_1349);
or U362 (N_362,In_128,In_1011);
nor U363 (N_363,In_940,In_194);
nand U364 (N_364,In_1232,In_316);
nor U365 (N_365,In_158,In_23);
nand U366 (N_366,In_1042,In_903);
nor U367 (N_367,In_313,In_104);
and U368 (N_368,In_1182,In_599);
or U369 (N_369,In_447,In_572);
and U370 (N_370,In_904,In_551);
or U371 (N_371,In_1475,In_1085);
nand U372 (N_372,In_707,In_1376);
or U373 (N_373,In_863,In_309);
or U374 (N_374,In_256,In_400);
nor U375 (N_375,In_977,In_1170);
and U376 (N_376,In_1465,In_1047);
nand U377 (N_377,In_828,In_864);
and U378 (N_378,In_1279,In_758);
nor U379 (N_379,In_887,In_563);
and U380 (N_380,In_205,In_1359);
nand U381 (N_381,In_463,In_1438);
nor U382 (N_382,In_1129,In_204);
nor U383 (N_383,In_268,In_32);
or U384 (N_384,In_882,In_495);
and U385 (N_385,In_1094,In_1382);
or U386 (N_386,In_1199,In_898);
nand U387 (N_387,In_945,In_438);
and U388 (N_388,In_528,In_1294);
nand U389 (N_389,In_1401,In_1463);
or U390 (N_390,In_676,In_1457);
nand U391 (N_391,In_936,In_938);
nor U392 (N_392,In_1474,In_530);
nand U393 (N_393,In_1305,In_1141);
and U394 (N_394,In_428,In_862);
nand U395 (N_395,In_1028,In_1117);
and U396 (N_396,In_532,In_975);
or U397 (N_397,In_633,In_1184);
and U398 (N_398,In_1,In_166);
nor U399 (N_399,In_1296,In_705);
nor U400 (N_400,In_1300,In_101);
or U401 (N_401,In_1393,In_1130);
or U402 (N_402,In_147,In_1111);
nor U403 (N_403,In_40,In_1241);
nor U404 (N_404,In_847,In_1492);
or U405 (N_405,In_1185,In_106);
and U406 (N_406,In_500,In_1225);
and U407 (N_407,In_1350,In_49);
nand U408 (N_408,In_395,In_799);
nand U409 (N_409,In_724,In_1373);
nand U410 (N_410,In_93,In_404);
nand U411 (N_411,In_1031,In_1213);
nand U412 (N_412,In_1160,In_1139);
or U413 (N_413,In_693,In_1074);
nor U414 (N_414,In_1265,In_996);
nand U415 (N_415,In_225,In_1481);
and U416 (N_416,In_804,In_1197);
and U417 (N_417,In_467,In_167);
nand U418 (N_418,In_891,In_276);
nand U419 (N_419,In_1266,In_638);
or U420 (N_420,In_439,In_1200);
xor U421 (N_421,In_824,In_272);
and U422 (N_422,In_765,In_1315);
nand U423 (N_423,In_796,In_577);
nand U424 (N_424,In_844,In_87);
nor U425 (N_425,In_111,In_719);
nor U426 (N_426,In_623,In_1175);
or U427 (N_427,In_381,In_54);
or U428 (N_428,In_922,In_885);
or U429 (N_429,In_1262,In_1415);
nand U430 (N_430,In_115,In_536);
or U431 (N_431,In_1404,In_1133);
nor U432 (N_432,In_902,In_1180);
nor U433 (N_433,In_1288,In_839);
nand U434 (N_434,In_820,In_611);
nand U435 (N_435,In_1177,In_448);
and U436 (N_436,In_425,In_1158);
nand U437 (N_437,In_238,In_81);
and U438 (N_438,In_151,In_35);
or U439 (N_439,In_392,In_259);
and U440 (N_440,In_1399,In_520);
xor U441 (N_441,In_485,In_6);
or U442 (N_442,In_673,In_784);
and U443 (N_443,In_176,In_1380);
nor U444 (N_444,In_728,In_1323);
nand U445 (N_445,In_931,In_504);
and U446 (N_446,In_1166,In_127);
or U447 (N_447,In_443,In_894);
or U448 (N_448,In_1413,In_933);
nor U449 (N_449,In_1105,In_135);
and U450 (N_450,In_21,In_821);
and U451 (N_451,In_451,In_260);
or U452 (N_452,In_1131,In_952);
or U453 (N_453,In_733,In_893);
or U454 (N_454,In_460,In_1287);
nand U455 (N_455,In_399,In_544);
nor U456 (N_456,In_725,In_1179);
nor U457 (N_457,In_30,In_1397);
and U458 (N_458,In_486,In_1473);
nand U459 (N_459,In_206,In_1417);
and U460 (N_460,In_1102,In_1134);
and U461 (N_461,In_880,In_9);
nand U462 (N_462,In_814,In_787);
xnor U463 (N_463,In_597,In_691);
and U464 (N_464,In_1204,In_325);
and U465 (N_465,In_351,In_100);
nand U466 (N_466,In_173,In_136);
or U467 (N_467,In_278,In_560);
nor U468 (N_468,In_1263,In_656);
or U469 (N_469,In_1159,In_1395);
nor U470 (N_470,In_442,In_1220);
nand U471 (N_471,In_1070,In_308);
nand U472 (N_472,In_1153,In_341);
or U473 (N_473,In_678,In_700);
nand U474 (N_474,In_437,In_937);
and U475 (N_475,In_1099,In_878);
or U476 (N_476,In_1251,In_1284);
and U477 (N_477,In_702,In_202);
nand U478 (N_478,In_1206,In_763);
nand U479 (N_479,In_670,In_72);
or U480 (N_480,In_614,In_731);
nand U481 (N_481,In_354,In_387);
or U482 (N_482,In_768,In_1120);
xor U483 (N_483,In_417,In_794);
nor U484 (N_484,In_740,In_905);
and U485 (N_485,In_1310,In_653);
and U486 (N_486,In_1209,In_1045);
and U487 (N_487,In_1093,In_1327);
nor U488 (N_488,In_662,In_538);
or U489 (N_489,In_658,In_1307);
or U490 (N_490,In_181,In_605);
or U491 (N_491,In_189,In_600);
and U492 (N_492,In_275,In_595);
or U493 (N_493,In_1440,In_643);
and U494 (N_494,In_1215,In_473);
or U495 (N_495,In_798,In_961);
nor U496 (N_496,In_90,In_430);
or U497 (N_497,In_681,In_58);
nor U498 (N_498,In_150,In_521);
nand U499 (N_499,In_331,In_18);
nand U500 (N_500,In_723,In_1005);
nor U501 (N_501,In_85,In_1162);
xor U502 (N_502,In_188,In_1489);
and U503 (N_503,In_1240,In_1320);
nor U504 (N_504,In_960,In_130);
nand U505 (N_505,In_1233,In_718);
or U506 (N_506,In_1414,In_899);
and U507 (N_507,In_1012,In_1486);
or U508 (N_508,In_1132,In_866);
and U509 (N_509,In_602,In_554);
nor U510 (N_510,In_832,In_809);
nor U511 (N_511,In_368,In_606);
and U512 (N_512,In_1351,In_1335);
nand U513 (N_513,In_1354,In_1250);
nand U514 (N_514,In_672,In_519);
or U515 (N_515,In_1167,In_1014);
or U516 (N_516,In_50,In_1360);
nor U517 (N_517,In_1173,In_590);
nor U518 (N_518,In_57,In_524);
and U519 (N_519,In_1403,In_96);
or U520 (N_520,In_149,In_665);
and U521 (N_521,In_1435,In_806);
or U522 (N_522,In_411,In_924);
nor U523 (N_523,In_1248,In_1291);
nor U524 (N_524,In_269,In_1015);
and U525 (N_525,In_980,In_288);
nand U526 (N_526,In_525,In_1216);
and U527 (N_527,In_496,In_68);
nor U528 (N_528,In_641,In_29);
nor U529 (N_529,In_752,In_1002);
nand U530 (N_530,In_1313,In_373);
and U531 (N_531,In_876,In_881);
or U532 (N_532,In_112,In_1312);
or U533 (N_533,In_951,In_1150);
and U534 (N_534,In_850,In_1334);
or U535 (N_535,In_1260,In_1183);
and U536 (N_536,In_888,In_822);
or U537 (N_537,In_77,In_388);
nor U538 (N_538,In_282,In_713);
or U539 (N_539,In_537,In_1178);
nor U540 (N_540,In_837,In_427);
nor U541 (N_541,In_795,In_627);
nor U542 (N_542,In_14,In_1423);
nand U543 (N_543,In_697,In_360);
nand U544 (N_544,In_0,In_879);
or U545 (N_545,In_1316,In_1152);
nand U546 (N_546,In_75,In_564);
nand U547 (N_547,In_802,In_1346);
nand U548 (N_548,In_285,In_301);
nor U549 (N_549,In_1019,In_184);
and U550 (N_550,In_526,In_374);
and U551 (N_551,In_1345,In_1222);
or U552 (N_552,In_1324,In_622);
nand U553 (N_553,In_581,In_780);
and U554 (N_554,In_1330,In_1367);
and U555 (N_555,In_306,In_1234);
nor U556 (N_556,In_141,In_578);
or U557 (N_557,In_386,In_819);
and U558 (N_558,In_223,In_568);
and U559 (N_559,In_1267,In_369);
nor U560 (N_560,In_396,In_284);
and U561 (N_561,In_99,In_203);
and U562 (N_562,In_570,In_94);
or U563 (N_563,In_291,In_258);
nand U564 (N_564,In_298,In_1054);
or U565 (N_565,In_1057,In_1456);
nand U566 (N_566,In_571,In_1436);
nor U567 (N_567,In_901,In_39);
and U568 (N_568,In_772,In_1381);
and U569 (N_569,In_444,In_12);
and U570 (N_570,In_959,In_1007);
nand U571 (N_571,In_513,In_1022);
nor U572 (N_572,In_196,In_1339);
or U573 (N_573,In_708,In_1329);
and U574 (N_574,In_382,In_1484);
and U575 (N_575,In_133,In_674);
and U576 (N_576,In_216,In_1273);
nand U577 (N_577,In_356,In_769);
nand U578 (N_578,In_1419,In_1317);
and U579 (N_579,In_465,In_469);
nor U580 (N_580,In_1254,In_1245);
and U581 (N_581,In_915,In_624);
nand U582 (N_582,In_1046,In_198);
and U583 (N_583,In_348,In_671);
nor U584 (N_584,In_518,In_1242);
or U585 (N_585,In_1264,In_7);
nor U586 (N_586,In_1398,In_1075);
nand U587 (N_587,In_661,In_655);
nand U588 (N_588,In_1459,In_31);
xnor U589 (N_589,In_126,In_749);
or U590 (N_590,In_1482,In_389);
and U591 (N_591,In_721,In_1402);
nor U592 (N_592,In_1137,In_679);
or U593 (N_593,In_789,In_408);
nor U594 (N_594,In_636,In_253);
or U595 (N_595,In_1190,In_523);
nand U596 (N_596,In_265,In_499);
nand U597 (N_597,In_555,In_800);
nand U598 (N_598,In_378,In_754);
or U599 (N_599,In_512,In_1425);
and U600 (N_600,In_262,In_236);
and U601 (N_601,In_366,In_1405);
nor U602 (N_602,In_403,In_1445);
and U603 (N_603,In_956,In_52);
or U604 (N_604,In_955,In_946);
nor U605 (N_605,In_1383,In_842);
nand U606 (N_606,In_434,In_896);
nor U607 (N_607,In_353,In_966);
or U608 (N_608,In_797,In_739);
and U609 (N_609,In_629,In_861);
nand U610 (N_610,In_1416,In_963);
nand U611 (N_611,In_91,In_1211);
nor U612 (N_612,In_159,In_420);
and U613 (N_613,In_1488,In_302);
nor U614 (N_614,In_715,In_1066);
or U615 (N_615,In_129,In_1256);
or U616 (N_616,In_1348,In_390);
and U617 (N_617,In_683,In_954);
and U618 (N_618,In_1364,In_231);
nand U619 (N_619,In_1272,In_192);
nand U620 (N_620,In_1269,In_294);
and U621 (N_621,In_1217,In_261);
or U622 (N_622,In_211,In_1268);
and U623 (N_623,In_218,In_833);
and U624 (N_624,In_1058,In_1252);
nor U625 (N_625,In_567,In_116);
nand U626 (N_626,In_375,In_593);
and U627 (N_627,In_857,In_1255);
nor U628 (N_628,In_511,In_1037);
nand U629 (N_629,In_489,In_229);
and U630 (N_630,In_295,In_914);
and U631 (N_631,In_118,In_774);
nor U632 (N_632,In_1356,In_1018);
nor U633 (N_633,In_853,In_1283);
or U634 (N_634,In_934,In_1034);
nor U635 (N_635,In_1365,In_56);
nor U636 (N_636,In_142,In_628);
and U637 (N_637,In_234,In_935);
or U638 (N_638,In_815,In_71);
nand U639 (N_639,In_274,In_610);
or U640 (N_640,In_407,In_488);
nor U641 (N_641,In_1202,In_640);
nand U642 (N_642,In_805,In_501);
nand U643 (N_643,In_543,In_60);
nand U644 (N_644,In_113,In_393);
and U645 (N_645,In_1097,In_921);
nor U646 (N_646,In_172,In_300);
nand U647 (N_647,In_180,In_365);
nor U648 (N_648,In_105,In_27);
and U649 (N_649,In_944,In_836);
or U650 (N_650,In_675,In_1103);
nor U651 (N_651,In_293,In_1164);
nor U652 (N_652,In_562,In_1157);
or U653 (N_653,In_508,In_897);
or U654 (N_654,In_747,In_619);
nor U655 (N_655,In_201,In_1374);
nor U656 (N_656,In_992,In_409);
or U657 (N_657,In_949,In_121);
and U658 (N_658,In_95,In_669);
or U659 (N_659,In_426,In_193);
and U660 (N_660,In_1301,In_859);
nand U661 (N_661,In_968,In_1174);
and U662 (N_662,In_1061,In_773);
and U663 (N_663,In_89,In_346);
nor U664 (N_664,In_1235,In_24);
or U665 (N_665,In_1495,In_233);
or U666 (N_666,In_1115,In_330);
nand U667 (N_667,In_1210,In_696);
and U668 (N_668,In_983,In_362);
nor U669 (N_669,In_607,In_64);
nor U670 (N_670,In_221,In_1246);
nand U671 (N_671,In_307,In_1471);
nand U672 (N_672,In_73,In_910);
nand U673 (N_673,In_1077,In_695);
and U674 (N_674,In_42,In_466);
nor U675 (N_675,In_1176,In_134);
or U676 (N_676,In_132,In_277);
or U677 (N_677,In_187,In_103);
nand U678 (N_678,In_618,In_1479);
and U679 (N_679,In_355,In_743);
and U680 (N_680,In_1468,In_454);
nand U681 (N_681,In_635,In_778);
and U682 (N_682,In_895,In_243);
nand U683 (N_683,In_401,In_185);
and U684 (N_684,In_481,In_1109);
nor U685 (N_685,In_825,In_410);
or U686 (N_686,In_612,In_1390);
nand U687 (N_687,In_1126,In_1025);
or U688 (N_688,In_230,In_529);
or U689 (N_689,In_38,In_1318);
and U690 (N_690,In_664,In_1422);
nand U691 (N_691,In_1169,In_1259);
or U692 (N_692,In_120,In_1434);
nor U693 (N_693,In_1155,In_652);
nand U694 (N_694,In_889,In_457);
nand U695 (N_695,In_1193,In_1148);
nor U696 (N_696,In_516,In_685);
and U697 (N_697,In_813,In_305);
nor U698 (N_698,In_646,In_250);
nor U699 (N_699,In_1006,In_163);
or U700 (N_700,In_1451,In_429);
or U701 (N_701,In_88,In_1333);
nand U702 (N_702,In_767,In_1341);
or U703 (N_703,In_61,In_347);
or U704 (N_704,In_1478,In_589);
nand U705 (N_705,In_372,In_1340);
and U706 (N_706,In_999,In_1040);
xnor U707 (N_707,In_1086,In_468);
nor U708 (N_708,In_286,In_339);
and U709 (N_709,In_36,In_343);
nand U710 (N_710,In_1461,In_319);
nor U711 (N_711,In_144,In_22);
nor U712 (N_712,In_742,In_458);
nand U713 (N_713,In_1013,In_164);
or U714 (N_714,In_78,In_1469);
and U715 (N_715,In_161,In_304);
nor U716 (N_716,In_1452,In_884);
nor U717 (N_717,In_592,In_998);
nor U718 (N_718,In_786,In_722);
nand U719 (N_719,In_292,In_1342);
or U720 (N_720,In_257,In_179);
and U721 (N_721,In_872,In_226);
nand U722 (N_722,In_1051,In_228);
nand U723 (N_723,In_776,In_858);
and U724 (N_724,In_1112,In_514);
nor U725 (N_725,In_1271,In_644);
nand U726 (N_726,In_249,In_490);
nand U727 (N_727,In_1431,In_533);
or U728 (N_728,In_1363,In_943);
or U729 (N_729,In_55,In_916);
nand U730 (N_730,In_745,In_1328);
or U731 (N_731,In_647,In_1056);
or U732 (N_732,In_324,In_642);
or U733 (N_733,In_668,In_654);
or U734 (N_734,In_122,In_69);
nor U735 (N_735,In_1411,In_397);
or U736 (N_736,In_169,In_505);
and U737 (N_737,In_84,In_143);
and U738 (N_738,In_870,In_92);
nor U739 (N_739,In_701,In_1224);
nor U740 (N_740,In_1010,In_1113);
and U741 (N_741,In_550,In_1386);
nand U742 (N_742,In_834,In_1389);
nor U743 (N_743,In_737,In_1304);
nor U744 (N_744,In_883,In_631);
and U745 (N_745,In_471,In_666);
or U746 (N_746,In_986,In_930);
nand U747 (N_747,In_1387,In_994);
and U748 (N_748,In_1424,In_415);
nor U749 (N_749,In_714,In_117);
nand U750 (N_750,In_985,In_312);
or U751 (N_751,In_40,In_671);
nand U752 (N_752,In_1398,In_307);
nand U753 (N_753,In_1001,In_712);
nand U754 (N_754,In_174,In_1397);
nand U755 (N_755,In_1478,In_372);
nand U756 (N_756,In_1076,In_536);
and U757 (N_757,In_517,In_863);
or U758 (N_758,In_284,In_614);
nand U759 (N_759,In_1382,In_1279);
and U760 (N_760,In_1099,In_148);
or U761 (N_761,In_119,In_913);
nor U762 (N_762,In_764,In_295);
or U763 (N_763,In_1385,In_1236);
and U764 (N_764,In_1314,In_43);
or U765 (N_765,In_989,In_1058);
nor U766 (N_766,In_620,In_797);
nand U767 (N_767,In_1397,In_1403);
or U768 (N_768,In_253,In_350);
nor U769 (N_769,In_947,In_92);
nor U770 (N_770,In_145,In_1292);
nand U771 (N_771,In_1041,In_733);
nor U772 (N_772,In_1328,In_872);
nor U773 (N_773,In_922,In_1266);
nor U774 (N_774,In_110,In_591);
nor U775 (N_775,In_1442,In_1220);
or U776 (N_776,In_916,In_1279);
nor U777 (N_777,In_478,In_853);
or U778 (N_778,In_648,In_1377);
nand U779 (N_779,In_448,In_1176);
nor U780 (N_780,In_454,In_879);
and U781 (N_781,In_519,In_942);
or U782 (N_782,In_667,In_478);
or U783 (N_783,In_1377,In_427);
or U784 (N_784,In_1051,In_1273);
or U785 (N_785,In_1226,In_1310);
nor U786 (N_786,In_122,In_1106);
nand U787 (N_787,In_1139,In_1290);
or U788 (N_788,In_1453,In_1120);
or U789 (N_789,In_914,In_36);
and U790 (N_790,In_584,In_909);
and U791 (N_791,In_234,In_1380);
or U792 (N_792,In_728,In_123);
or U793 (N_793,In_989,In_153);
and U794 (N_794,In_1446,In_436);
or U795 (N_795,In_222,In_1376);
and U796 (N_796,In_426,In_369);
or U797 (N_797,In_1138,In_618);
nand U798 (N_798,In_1403,In_454);
and U799 (N_799,In_722,In_617);
nand U800 (N_800,In_473,In_540);
or U801 (N_801,In_1116,In_457);
nor U802 (N_802,In_661,In_453);
and U803 (N_803,In_710,In_505);
and U804 (N_804,In_1216,In_226);
or U805 (N_805,In_1079,In_1434);
and U806 (N_806,In_1311,In_1008);
or U807 (N_807,In_482,In_1213);
or U808 (N_808,In_1384,In_1385);
or U809 (N_809,In_193,In_131);
and U810 (N_810,In_830,In_1237);
or U811 (N_811,In_831,In_32);
nand U812 (N_812,In_1458,In_703);
nand U813 (N_813,In_1127,In_986);
nand U814 (N_814,In_385,In_852);
and U815 (N_815,In_623,In_1416);
nor U816 (N_816,In_421,In_42);
nor U817 (N_817,In_156,In_867);
and U818 (N_818,In_1248,In_610);
or U819 (N_819,In_1189,In_126);
or U820 (N_820,In_475,In_340);
nand U821 (N_821,In_337,In_882);
nor U822 (N_822,In_825,In_1450);
and U823 (N_823,In_1115,In_666);
nor U824 (N_824,In_286,In_1245);
nand U825 (N_825,In_123,In_96);
or U826 (N_826,In_486,In_653);
or U827 (N_827,In_1348,In_997);
nor U828 (N_828,In_1180,In_243);
nor U829 (N_829,In_606,In_461);
or U830 (N_830,In_1336,In_306);
nand U831 (N_831,In_160,In_353);
and U832 (N_832,In_1259,In_1266);
nor U833 (N_833,In_219,In_1486);
nor U834 (N_834,In_1090,In_216);
or U835 (N_835,In_1205,In_840);
nand U836 (N_836,In_621,In_1414);
nand U837 (N_837,In_1286,In_1168);
nor U838 (N_838,In_532,In_1012);
nor U839 (N_839,In_1209,In_668);
or U840 (N_840,In_226,In_263);
nand U841 (N_841,In_569,In_1344);
nand U842 (N_842,In_643,In_407);
nand U843 (N_843,In_894,In_47);
nor U844 (N_844,In_350,In_1218);
and U845 (N_845,In_1002,In_1422);
nand U846 (N_846,In_115,In_593);
or U847 (N_847,In_1042,In_446);
or U848 (N_848,In_1265,In_856);
and U849 (N_849,In_478,In_611);
nand U850 (N_850,In_1254,In_221);
and U851 (N_851,In_1153,In_734);
and U852 (N_852,In_1261,In_1273);
nand U853 (N_853,In_60,In_585);
or U854 (N_854,In_1351,In_1461);
nor U855 (N_855,In_1374,In_1148);
nor U856 (N_856,In_470,In_126);
nand U857 (N_857,In_210,In_1225);
and U858 (N_858,In_460,In_1250);
nand U859 (N_859,In_832,In_196);
nor U860 (N_860,In_945,In_1377);
nand U861 (N_861,In_1419,In_610);
nor U862 (N_862,In_777,In_1348);
or U863 (N_863,In_112,In_766);
or U864 (N_864,In_1363,In_704);
nand U865 (N_865,In_748,In_1053);
or U866 (N_866,In_276,In_794);
nand U867 (N_867,In_559,In_315);
nor U868 (N_868,In_481,In_1469);
and U869 (N_869,In_445,In_256);
nand U870 (N_870,In_1007,In_1107);
or U871 (N_871,In_347,In_1169);
or U872 (N_872,In_381,In_273);
nand U873 (N_873,In_1258,In_1389);
or U874 (N_874,In_590,In_666);
or U875 (N_875,In_1334,In_1197);
or U876 (N_876,In_927,In_1267);
nor U877 (N_877,In_619,In_98);
nor U878 (N_878,In_1368,In_244);
or U879 (N_879,In_916,In_702);
nor U880 (N_880,In_1313,In_625);
or U881 (N_881,In_315,In_115);
nand U882 (N_882,In_1366,In_1301);
and U883 (N_883,In_1443,In_64);
nand U884 (N_884,In_1006,In_466);
or U885 (N_885,In_1441,In_56);
nand U886 (N_886,In_1076,In_402);
and U887 (N_887,In_1386,In_126);
or U888 (N_888,In_1279,In_68);
and U889 (N_889,In_973,In_235);
nand U890 (N_890,In_882,In_109);
or U891 (N_891,In_1361,In_1013);
and U892 (N_892,In_311,In_1321);
or U893 (N_893,In_81,In_165);
or U894 (N_894,In_851,In_581);
nand U895 (N_895,In_778,In_548);
or U896 (N_896,In_748,In_679);
nor U897 (N_897,In_78,In_1146);
and U898 (N_898,In_1346,In_832);
nand U899 (N_899,In_191,In_653);
or U900 (N_900,In_273,In_66);
and U901 (N_901,In_1135,In_1316);
and U902 (N_902,In_1389,In_954);
or U903 (N_903,In_410,In_1153);
nor U904 (N_904,In_664,In_7);
nor U905 (N_905,In_1475,In_331);
or U906 (N_906,In_103,In_1237);
nor U907 (N_907,In_43,In_567);
and U908 (N_908,In_55,In_1393);
or U909 (N_909,In_1251,In_248);
or U910 (N_910,In_761,In_636);
or U911 (N_911,In_1189,In_511);
nor U912 (N_912,In_574,In_1059);
or U913 (N_913,In_1354,In_980);
or U914 (N_914,In_848,In_1419);
and U915 (N_915,In_1479,In_1372);
or U916 (N_916,In_902,In_1076);
nand U917 (N_917,In_88,In_834);
nor U918 (N_918,In_1483,In_1495);
and U919 (N_919,In_315,In_19);
nor U920 (N_920,In_671,In_929);
and U921 (N_921,In_115,In_676);
nor U922 (N_922,In_448,In_458);
nand U923 (N_923,In_760,In_1204);
nand U924 (N_924,In_755,In_1445);
nor U925 (N_925,In_277,In_293);
nand U926 (N_926,In_995,In_1209);
nor U927 (N_927,In_936,In_299);
nand U928 (N_928,In_1474,In_1082);
nand U929 (N_929,In_358,In_1162);
and U930 (N_930,In_903,In_777);
or U931 (N_931,In_1258,In_186);
nor U932 (N_932,In_1376,In_796);
or U933 (N_933,In_864,In_798);
or U934 (N_934,In_216,In_65);
and U935 (N_935,In_1371,In_860);
nand U936 (N_936,In_1284,In_742);
and U937 (N_937,In_282,In_201);
nand U938 (N_938,In_1168,In_1031);
nand U939 (N_939,In_282,In_545);
nor U940 (N_940,In_129,In_349);
and U941 (N_941,In_1053,In_492);
or U942 (N_942,In_366,In_685);
or U943 (N_943,In_695,In_653);
or U944 (N_944,In_1088,In_1264);
nand U945 (N_945,In_1372,In_1324);
nand U946 (N_946,In_1453,In_779);
nor U947 (N_947,In_579,In_12);
or U948 (N_948,In_805,In_1300);
and U949 (N_949,In_1441,In_544);
or U950 (N_950,In_362,In_410);
nor U951 (N_951,In_1151,In_1221);
and U952 (N_952,In_1363,In_1018);
or U953 (N_953,In_955,In_1085);
nor U954 (N_954,In_382,In_521);
or U955 (N_955,In_1161,In_818);
nor U956 (N_956,In_808,In_1074);
and U957 (N_957,In_1499,In_263);
and U958 (N_958,In_1246,In_369);
xnor U959 (N_959,In_576,In_1014);
nor U960 (N_960,In_314,In_92);
nand U961 (N_961,In_211,In_287);
nand U962 (N_962,In_440,In_263);
or U963 (N_963,In_935,In_1446);
or U964 (N_964,In_698,In_152);
and U965 (N_965,In_352,In_943);
nand U966 (N_966,In_930,In_447);
or U967 (N_967,In_1372,In_462);
nor U968 (N_968,In_1059,In_1053);
and U969 (N_969,In_1031,In_1397);
or U970 (N_970,In_308,In_228);
xor U971 (N_971,In_209,In_255);
and U972 (N_972,In_151,In_1220);
and U973 (N_973,In_679,In_309);
or U974 (N_974,In_77,In_37);
nor U975 (N_975,In_7,In_692);
nor U976 (N_976,In_1302,In_1437);
or U977 (N_977,In_943,In_1085);
or U978 (N_978,In_1018,In_336);
nand U979 (N_979,In_1361,In_917);
nand U980 (N_980,In_1034,In_157);
and U981 (N_981,In_933,In_1394);
and U982 (N_982,In_723,In_1308);
nand U983 (N_983,In_1295,In_1394);
or U984 (N_984,In_959,In_736);
and U985 (N_985,In_92,In_808);
nor U986 (N_986,In_184,In_775);
and U987 (N_987,In_75,In_1124);
or U988 (N_988,In_458,In_447);
nor U989 (N_989,In_1315,In_632);
xor U990 (N_990,In_114,In_1475);
nor U991 (N_991,In_1295,In_876);
or U992 (N_992,In_835,In_932);
nand U993 (N_993,In_602,In_344);
xor U994 (N_994,In_273,In_17);
or U995 (N_995,In_850,In_784);
xnor U996 (N_996,In_1383,In_422);
and U997 (N_997,In_256,In_770);
nor U998 (N_998,In_605,In_112);
nand U999 (N_999,In_1153,In_1357);
or U1000 (N_1000,In_737,In_1278);
nor U1001 (N_1001,In_538,In_940);
nor U1002 (N_1002,In_1488,In_1279);
and U1003 (N_1003,In_943,In_87);
and U1004 (N_1004,In_77,In_229);
nor U1005 (N_1005,In_721,In_1370);
and U1006 (N_1006,In_138,In_598);
and U1007 (N_1007,In_52,In_180);
nand U1008 (N_1008,In_710,In_894);
and U1009 (N_1009,In_625,In_1432);
nor U1010 (N_1010,In_1202,In_1209);
nand U1011 (N_1011,In_978,In_701);
and U1012 (N_1012,In_851,In_1215);
or U1013 (N_1013,In_1332,In_218);
nand U1014 (N_1014,In_653,In_685);
nand U1015 (N_1015,In_604,In_882);
nand U1016 (N_1016,In_90,In_315);
or U1017 (N_1017,In_970,In_439);
nor U1018 (N_1018,In_619,In_302);
nor U1019 (N_1019,In_223,In_719);
and U1020 (N_1020,In_435,In_933);
nor U1021 (N_1021,In_1250,In_1056);
nor U1022 (N_1022,In_564,In_12);
or U1023 (N_1023,In_505,In_1178);
or U1024 (N_1024,In_1004,In_138);
nand U1025 (N_1025,In_496,In_1298);
or U1026 (N_1026,In_414,In_526);
and U1027 (N_1027,In_1288,In_1084);
or U1028 (N_1028,In_313,In_145);
and U1029 (N_1029,In_994,In_965);
nor U1030 (N_1030,In_848,In_158);
nor U1031 (N_1031,In_586,In_44);
nand U1032 (N_1032,In_252,In_742);
nor U1033 (N_1033,In_1388,In_960);
xnor U1034 (N_1034,In_1227,In_1274);
or U1035 (N_1035,In_1215,In_836);
and U1036 (N_1036,In_1478,In_598);
and U1037 (N_1037,In_208,In_762);
and U1038 (N_1038,In_838,In_463);
or U1039 (N_1039,In_1405,In_1110);
and U1040 (N_1040,In_1316,In_747);
nor U1041 (N_1041,In_267,In_584);
nor U1042 (N_1042,In_203,In_1188);
and U1043 (N_1043,In_963,In_1438);
nand U1044 (N_1044,In_1414,In_587);
and U1045 (N_1045,In_471,In_805);
and U1046 (N_1046,In_672,In_774);
and U1047 (N_1047,In_386,In_291);
nor U1048 (N_1048,In_158,In_497);
nor U1049 (N_1049,In_1260,In_642);
and U1050 (N_1050,In_815,In_1096);
or U1051 (N_1051,In_773,In_260);
nand U1052 (N_1052,In_18,In_1094);
nand U1053 (N_1053,In_454,In_541);
nand U1054 (N_1054,In_741,In_5);
and U1055 (N_1055,In_849,In_1050);
or U1056 (N_1056,In_1492,In_56);
and U1057 (N_1057,In_245,In_887);
and U1058 (N_1058,In_940,In_1205);
nor U1059 (N_1059,In_643,In_35);
or U1060 (N_1060,In_1227,In_1298);
and U1061 (N_1061,In_337,In_338);
and U1062 (N_1062,In_26,In_1336);
or U1063 (N_1063,In_161,In_595);
and U1064 (N_1064,In_764,In_1458);
nand U1065 (N_1065,In_483,In_1434);
nand U1066 (N_1066,In_842,In_546);
nand U1067 (N_1067,In_366,In_1444);
nor U1068 (N_1068,In_1157,In_145);
or U1069 (N_1069,In_1399,In_860);
nand U1070 (N_1070,In_1280,In_88);
nand U1071 (N_1071,In_1201,In_804);
nand U1072 (N_1072,In_868,In_1299);
nand U1073 (N_1073,In_772,In_920);
nand U1074 (N_1074,In_778,In_649);
nor U1075 (N_1075,In_1114,In_908);
or U1076 (N_1076,In_1045,In_653);
and U1077 (N_1077,In_712,In_1341);
or U1078 (N_1078,In_522,In_9);
nor U1079 (N_1079,In_382,In_154);
nand U1080 (N_1080,In_1466,In_1377);
and U1081 (N_1081,In_1083,In_52);
and U1082 (N_1082,In_178,In_489);
nor U1083 (N_1083,In_1342,In_237);
or U1084 (N_1084,In_229,In_128);
and U1085 (N_1085,In_47,In_245);
xor U1086 (N_1086,In_1185,In_849);
and U1087 (N_1087,In_778,In_6);
or U1088 (N_1088,In_1135,In_81);
and U1089 (N_1089,In_588,In_1040);
or U1090 (N_1090,In_249,In_1287);
or U1091 (N_1091,In_1410,In_281);
and U1092 (N_1092,In_1366,In_847);
nor U1093 (N_1093,In_120,In_125);
nand U1094 (N_1094,In_1124,In_1017);
or U1095 (N_1095,In_1172,In_121);
and U1096 (N_1096,In_361,In_1087);
nor U1097 (N_1097,In_434,In_866);
and U1098 (N_1098,In_965,In_6);
nor U1099 (N_1099,In_1090,In_1016);
nand U1100 (N_1100,In_72,In_2);
and U1101 (N_1101,In_1118,In_739);
nor U1102 (N_1102,In_867,In_550);
nand U1103 (N_1103,In_912,In_660);
nand U1104 (N_1104,In_496,In_342);
or U1105 (N_1105,In_1033,In_217);
nor U1106 (N_1106,In_522,In_1097);
nor U1107 (N_1107,In_1389,In_546);
nand U1108 (N_1108,In_160,In_720);
nor U1109 (N_1109,In_676,In_372);
or U1110 (N_1110,In_908,In_845);
nor U1111 (N_1111,In_1371,In_944);
nor U1112 (N_1112,In_312,In_1246);
and U1113 (N_1113,In_753,In_1488);
or U1114 (N_1114,In_335,In_1333);
or U1115 (N_1115,In_734,In_1393);
nor U1116 (N_1116,In_1338,In_540);
nand U1117 (N_1117,In_749,In_357);
nand U1118 (N_1118,In_451,In_577);
or U1119 (N_1119,In_1004,In_745);
nand U1120 (N_1120,In_1192,In_783);
nand U1121 (N_1121,In_988,In_221);
nand U1122 (N_1122,In_909,In_757);
nand U1123 (N_1123,In_824,In_619);
nand U1124 (N_1124,In_653,In_302);
or U1125 (N_1125,In_117,In_116);
nand U1126 (N_1126,In_1015,In_1040);
or U1127 (N_1127,In_659,In_549);
and U1128 (N_1128,In_1453,In_1114);
nor U1129 (N_1129,In_491,In_1007);
xnor U1130 (N_1130,In_51,In_798);
and U1131 (N_1131,In_748,In_506);
or U1132 (N_1132,In_1107,In_437);
nand U1133 (N_1133,In_229,In_895);
and U1134 (N_1134,In_1035,In_187);
nand U1135 (N_1135,In_1101,In_1488);
nor U1136 (N_1136,In_655,In_1070);
and U1137 (N_1137,In_505,In_413);
and U1138 (N_1138,In_690,In_176);
nor U1139 (N_1139,In_827,In_643);
or U1140 (N_1140,In_111,In_791);
or U1141 (N_1141,In_921,In_278);
and U1142 (N_1142,In_322,In_207);
and U1143 (N_1143,In_450,In_273);
or U1144 (N_1144,In_42,In_503);
and U1145 (N_1145,In_438,In_1053);
nand U1146 (N_1146,In_1113,In_568);
or U1147 (N_1147,In_968,In_801);
nor U1148 (N_1148,In_523,In_1214);
nor U1149 (N_1149,In_1478,In_1205);
and U1150 (N_1150,In_268,In_388);
nand U1151 (N_1151,In_5,In_284);
or U1152 (N_1152,In_1105,In_701);
xor U1153 (N_1153,In_550,In_1095);
nand U1154 (N_1154,In_606,In_1137);
or U1155 (N_1155,In_407,In_752);
and U1156 (N_1156,In_1147,In_1320);
or U1157 (N_1157,In_882,In_1085);
nor U1158 (N_1158,In_152,In_611);
and U1159 (N_1159,In_466,In_641);
nor U1160 (N_1160,In_1232,In_693);
or U1161 (N_1161,In_151,In_1375);
nand U1162 (N_1162,In_630,In_521);
nand U1163 (N_1163,In_1475,In_46);
or U1164 (N_1164,In_917,In_828);
nor U1165 (N_1165,In_1369,In_642);
or U1166 (N_1166,In_322,In_679);
and U1167 (N_1167,In_483,In_849);
nand U1168 (N_1168,In_3,In_767);
and U1169 (N_1169,In_336,In_1148);
or U1170 (N_1170,In_390,In_241);
and U1171 (N_1171,In_837,In_1077);
or U1172 (N_1172,In_1437,In_1063);
nor U1173 (N_1173,In_1386,In_721);
nor U1174 (N_1174,In_1180,In_170);
nor U1175 (N_1175,In_13,In_437);
or U1176 (N_1176,In_1106,In_1281);
and U1177 (N_1177,In_726,In_1201);
nand U1178 (N_1178,In_552,In_519);
nor U1179 (N_1179,In_752,In_514);
and U1180 (N_1180,In_31,In_698);
or U1181 (N_1181,In_880,In_596);
or U1182 (N_1182,In_1498,In_135);
nor U1183 (N_1183,In_922,In_1057);
or U1184 (N_1184,In_819,In_388);
and U1185 (N_1185,In_854,In_1381);
nand U1186 (N_1186,In_1274,In_1106);
nor U1187 (N_1187,In_1280,In_267);
and U1188 (N_1188,In_167,In_1361);
xor U1189 (N_1189,In_433,In_448);
nand U1190 (N_1190,In_152,In_1278);
xnor U1191 (N_1191,In_101,In_1464);
and U1192 (N_1192,In_438,In_1267);
or U1193 (N_1193,In_951,In_575);
nand U1194 (N_1194,In_119,In_1114);
or U1195 (N_1195,In_270,In_1037);
and U1196 (N_1196,In_546,In_137);
nor U1197 (N_1197,In_621,In_337);
or U1198 (N_1198,In_1444,In_279);
or U1199 (N_1199,In_1071,In_1011);
or U1200 (N_1200,In_604,In_497);
nand U1201 (N_1201,In_1184,In_1014);
nand U1202 (N_1202,In_1423,In_15);
nand U1203 (N_1203,In_841,In_580);
nand U1204 (N_1204,In_428,In_628);
or U1205 (N_1205,In_1368,In_838);
xor U1206 (N_1206,In_232,In_681);
nand U1207 (N_1207,In_778,In_330);
nand U1208 (N_1208,In_1405,In_1457);
nor U1209 (N_1209,In_906,In_684);
or U1210 (N_1210,In_1364,In_1029);
or U1211 (N_1211,In_812,In_781);
nand U1212 (N_1212,In_1324,In_51);
nor U1213 (N_1213,In_1253,In_401);
nand U1214 (N_1214,In_1122,In_59);
nand U1215 (N_1215,In_1093,In_1176);
nor U1216 (N_1216,In_1081,In_871);
and U1217 (N_1217,In_1327,In_23);
nor U1218 (N_1218,In_1105,In_356);
nand U1219 (N_1219,In_292,In_1407);
nor U1220 (N_1220,In_1334,In_614);
nand U1221 (N_1221,In_1439,In_1441);
nor U1222 (N_1222,In_611,In_306);
nand U1223 (N_1223,In_358,In_1248);
nand U1224 (N_1224,In_670,In_163);
or U1225 (N_1225,In_1020,In_1226);
nand U1226 (N_1226,In_604,In_806);
nand U1227 (N_1227,In_688,In_212);
nor U1228 (N_1228,In_806,In_301);
nand U1229 (N_1229,In_1231,In_1368);
nand U1230 (N_1230,In_1181,In_411);
or U1231 (N_1231,In_554,In_428);
nor U1232 (N_1232,In_36,In_1214);
nor U1233 (N_1233,In_854,In_374);
nand U1234 (N_1234,In_1104,In_61);
or U1235 (N_1235,In_1309,In_346);
nand U1236 (N_1236,In_366,In_901);
nor U1237 (N_1237,In_630,In_535);
nor U1238 (N_1238,In_1255,In_1157);
nor U1239 (N_1239,In_220,In_39);
nand U1240 (N_1240,In_1298,In_633);
nand U1241 (N_1241,In_967,In_309);
nand U1242 (N_1242,In_173,In_147);
and U1243 (N_1243,In_78,In_1223);
nand U1244 (N_1244,In_61,In_241);
nor U1245 (N_1245,In_569,In_1056);
and U1246 (N_1246,In_1353,In_1076);
or U1247 (N_1247,In_573,In_43);
or U1248 (N_1248,In_105,In_488);
or U1249 (N_1249,In_1318,In_800);
or U1250 (N_1250,In_892,In_1242);
or U1251 (N_1251,In_439,In_521);
nand U1252 (N_1252,In_1287,In_621);
nand U1253 (N_1253,In_1269,In_345);
or U1254 (N_1254,In_0,In_658);
nor U1255 (N_1255,In_505,In_1310);
nor U1256 (N_1256,In_1277,In_556);
nor U1257 (N_1257,In_852,In_792);
and U1258 (N_1258,In_1287,In_837);
or U1259 (N_1259,In_98,In_794);
or U1260 (N_1260,In_323,In_799);
and U1261 (N_1261,In_1131,In_468);
or U1262 (N_1262,In_1227,In_939);
nand U1263 (N_1263,In_1034,In_1196);
nand U1264 (N_1264,In_1411,In_1499);
or U1265 (N_1265,In_863,In_208);
and U1266 (N_1266,In_113,In_250);
and U1267 (N_1267,In_67,In_1001);
nor U1268 (N_1268,In_638,In_189);
nor U1269 (N_1269,In_763,In_731);
and U1270 (N_1270,In_561,In_186);
and U1271 (N_1271,In_231,In_292);
or U1272 (N_1272,In_294,In_1231);
or U1273 (N_1273,In_353,In_861);
nand U1274 (N_1274,In_281,In_1311);
xnor U1275 (N_1275,In_76,In_933);
and U1276 (N_1276,In_1238,In_843);
nand U1277 (N_1277,In_475,In_1258);
or U1278 (N_1278,In_1460,In_795);
nand U1279 (N_1279,In_1489,In_1147);
nor U1280 (N_1280,In_985,In_1161);
or U1281 (N_1281,In_15,In_903);
and U1282 (N_1282,In_460,In_1495);
nand U1283 (N_1283,In_755,In_895);
nand U1284 (N_1284,In_1318,In_1157);
and U1285 (N_1285,In_541,In_841);
or U1286 (N_1286,In_1079,In_26);
or U1287 (N_1287,In_1492,In_690);
or U1288 (N_1288,In_1266,In_478);
and U1289 (N_1289,In_518,In_668);
or U1290 (N_1290,In_810,In_758);
and U1291 (N_1291,In_1478,In_403);
and U1292 (N_1292,In_203,In_842);
nor U1293 (N_1293,In_1257,In_794);
and U1294 (N_1294,In_1119,In_751);
and U1295 (N_1295,In_902,In_1127);
and U1296 (N_1296,In_987,In_233);
and U1297 (N_1297,In_446,In_1339);
nor U1298 (N_1298,In_1157,In_1256);
and U1299 (N_1299,In_45,In_527);
nand U1300 (N_1300,In_1208,In_1151);
nand U1301 (N_1301,In_1452,In_1148);
or U1302 (N_1302,In_64,In_1401);
nand U1303 (N_1303,In_1451,In_727);
nor U1304 (N_1304,In_819,In_1406);
nor U1305 (N_1305,In_174,In_79);
or U1306 (N_1306,In_1194,In_575);
nor U1307 (N_1307,In_433,In_682);
xnor U1308 (N_1308,In_1410,In_14);
nand U1309 (N_1309,In_1154,In_65);
and U1310 (N_1310,In_1023,In_1440);
or U1311 (N_1311,In_233,In_844);
nor U1312 (N_1312,In_370,In_1489);
nor U1313 (N_1313,In_923,In_1445);
and U1314 (N_1314,In_1038,In_586);
nand U1315 (N_1315,In_1178,In_790);
or U1316 (N_1316,In_1348,In_119);
and U1317 (N_1317,In_393,In_1039);
or U1318 (N_1318,In_50,In_428);
and U1319 (N_1319,In_220,In_880);
xnor U1320 (N_1320,In_859,In_713);
and U1321 (N_1321,In_224,In_232);
and U1322 (N_1322,In_69,In_1404);
nor U1323 (N_1323,In_579,In_1006);
nand U1324 (N_1324,In_1269,In_657);
or U1325 (N_1325,In_772,In_979);
nor U1326 (N_1326,In_945,In_148);
and U1327 (N_1327,In_764,In_772);
nand U1328 (N_1328,In_83,In_765);
or U1329 (N_1329,In_66,In_1344);
nor U1330 (N_1330,In_1107,In_373);
nand U1331 (N_1331,In_1227,In_137);
and U1332 (N_1332,In_44,In_414);
nand U1333 (N_1333,In_1317,In_375);
and U1334 (N_1334,In_13,In_1148);
or U1335 (N_1335,In_1075,In_1240);
or U1336 (N_1336,In_514,In_1180);
or U1337 (N_1337,In_127,In_952);
xor U1338 (N_1338,In_10,In_1026);
or U1339 (N_1339,In_958,In_1118);
nor U1340 (N_1340,In_399,In_764);
nand U1341 (N_1341,In_487,In_374);
and U1342 (N_1342,In_1324,In_1414);
nor U1343 (N_1343,In_1315,In_753);
or U1344 (N_1344,In_911,In_1346);
and U1345 (N_1345,In_288,In_1462);
or U1346 (N_1346,In_837,In_166);
or U1347 (N_1347,In_1390,In_700);
or U1348 (N_1348,In_1436,In_614);
or U1349 (N_1349,In_382,In_741);
nand U1350 (N_1350,In_202,In_304);
nand U1351 (N_1351,In_422,In_1013);
or U1352 (N_1352,In_1415,In_189);
nand U1353 (N_1353,In_695,In_788);
nand U1354 (N_1354,In_1160,In_371);
and U1355 (N_1355,In_1221,In_1359);
and U1356 (N_1356,In_1475,In_946);
or U1357 (N_1357,In_992,In_1161);
nor U1358 (N_1358,In_808,In_1393);
or U1359 (N_1359,In_1375,In_1003);
and U1360 (N_1360,In_1437,In_1176);
nand U1361 (N_1361,In_941,In_84);
and U1362 (N_1362,In_1305,In_830);
or U1363 (N_1363,In_254,In_1237);
nand U1364 (N_1364,In_1187,In_415);
or U1365 (N_1365,In_174,In_668);
nor U1366 (N_1366,In_95,In_774);
nor U1367 (N_1367,In_203,In_370);
nor U1368 (N_1368,In_1281,In_304);
nand U1369 (N_1369,In_146,In_1136);
or U1370 (N_1370,In_1170,In_123);
nor U1371 (N_1371,In_590,In_1022);
nor U1372 (N_1372,In_752,In_1101);
nor U1373 (N_1373,In_356,In_56);
and U1374 (N_1374,In_949,In_970);
and U1375 (N_1375,In_749,In_1434);
nand U1376 (N_1376,In_1288,In_583);
nand U1377 (N_1377,In_154,In_723);
or U1378 (N_1378,In_178,In_1122);
nand U1379 (N_1379,In_242,In_184);
nand U1380 (N_1380,In_191,In_250);
nor U1381 (N_1381,In_756,In_931);
nor U1382 (N_1382,In_1267,In_360);
nand U1383 (N_1383,In_1032,In_898);
nand U1384 (N_1384,In_649,In_846);
and U1385 (N_1385,In_1257,In_876);
nor U1386 (N_1386,In_673,In_388);
and U1387 (N_1387,In_1334,In_1346);
nor U1388 (N_1388,In_1111,In_450);
nor U1389 (N_1389,In_1099,In_543);
nor U1390 (N_1390,In_483,In_202);
nand U1391 (N_1391,In_773,In_18);
nor U1392 (N_1392,In_207,In_1455);
nand U1393 (N_1393,In_950,In_580);
nand U1394 (N_1394,In_720,In_119);
nand U1395 (N_1395,In_603,In_135);
or U1396 (N_1396,In_634,In_188);
and U1397 (N_1397,In_1422,In_398);
nand U1398 (N_1398,In_111,In_907);
or U1399 (N_1399,In_336,In_968);
nand U1400 (N_1400,In_601,In_245);
nor U1401 (N_1401,In_965,In_803);
nand U1402 (N_1402,In_1456,In_217);
and U1403 (N_1403,In_1127,In_1321);
and U1404 (N_1404,In_1403,In_809);
and U1405 (N_1405,In_973,In_1420);
and U1406 (N_1406,In_845,In_322);
nor U1407 (N_1407,In_1350,In_450);
nand U1408 (N_1408,In_120,In_1458);
nor U1409 (N_1409,In_1416,In_636);
nand U1410 (N_1410,In_47,In_1377);
nor U1411 (N_1411,In_595,In_1014);
and U1412 (N_1412,In_656,In_769);
nand U1413 (N_1413,In_908,In_977);
and U1414 (N_1414,In_1343,In_543);
and U1415 (N_1415,In_558,In_941);
and U1416 (N_1416,In_486,In_69);
nand U1417 (N_1417,In_117,In_952);
nor U1418 (N_1418,In_246,In_943);
and U1419 (N_1419,In_667,In_1108);
nand U1420 (N_1420,In_900,In_1326);
nor U1421 (N_1421,In_221,In_476);
or U1422 (N_1422,In_330,In_1162);
nor U1423 (N_1423,In_972,In_209);
nor U1424 (N_1424,In_1369,In_870);
and U1425 (N_1425,In_1495,In_1095);
or U1426 (N_1426,In_1098,In_228);
and U1427 (N_1427,In_297,In_151);
nor U1428 (N_1428,In_1430,In_456);
nand U1429 (N_1429,In_1454,In_1175);
nor U1430 (N_1430,In_700,In_925);
nor U1431 (N_1431,In_86,In_1328);
or U1432 (N_1432,In_1271,In_157);
nand U1433 (N_1433,In_1397,In_1369);
nor U1434 (N_1434,In_440,In_251);
nor U1435 (N_1435,In_167,In_445);
nand U1436 (N_1436,In_1462,In_383);
and U1437 (N_1437,In_755,In_1380);
nor U1438 (N_1438,In_237,In_456);
xnor U1439 (N_1439,In_760,In_734);
or U1440 (N_1440,In_154,In_46);
nor U1441 (N_1441,In_738,In_1417);
nor U1442 (N_1442,In_648,In_71);
nor U1443 (N_1443,In_1199,In_1427);
and U1444 (N_1444,In_1203,In_84);
or U1445 (N_1445,In_1365,In_979);
nor U1446 (N_1446,In_732,In_1301);
nor U1447 (N_1447,In_1347,In_796);
or U1448 (N_1448,In_342,In_212);
and U1449 (N_1449,In_1295,In_957);
nor U1450 (N_1450,In_898,In_1484);
or U1451 (N_1451,In_1373,In_697);
nor U1452 (N_1452,In_1037,In_106);
or U1453 (N_1453,In_1233,In_158);
nand U1454 (N_1454,In_808,In_517);
nor U1455 (N_1455,In_1011,In_1426);
or U1456 (N_1456,In_570,In_531);
and U1457 (N_1457,In_997,In_1401);
nor U1458 (N_1458,In_1383,In_608);
nor U1459 (N_1459,In_260,In_1213);
nand U1460 (N_1460,In_713,In_1);
or U1461 (N_1461,In_332,In_1207);
nor U1462 (N_1462,In_503,In_553);
nand U1463 (N_1463,In_992,In_475);
and U1464 (N_1464,In_6,In_829);
nor U1465 (N_1465,In_635,In_842);
nor U1466 (N_1466,In_582,In_785);
nand U1467 (N_1467,In_1284,In_522);
or U1468 (N_1468,In_952,In_1019);
or U1469 (N_1469,In_872,In_957);
nor U1470 (N_1470,In_359,In_1461);
nor U1471 (N_1471,In_367,In_1214);
nand U1472 (N_1472,In_173,In_1070);
nand U1473 (N_1473,In_164,In_941);
and U1474 (N_1474,In_42,In_102);
and U1475 (N_1475,In_1167,In_31);
nor U1476 (N_1476,In_775,In_136);
and U1477 (N_1477,In_410,In_136);
nand U1478 (N_1478,In_956,In_313);
or U1479 (N_1479,In_193,In_100);
or U1480 (N_1480,In_204,In_1325);
and U1481 (N_1481,In_1062,In_1094);
or U1482 (N_1482,In_391,In_269);
nor U1483 (N_1483,In_488,In_936);
nor U1484 (N_1484,In_626,In_502);
and U1485 (N_1485,In_461,In_1475);
nor U1486 (N_1486,In_605,In_234);
nor U1487 (N_1487,In_1262,In_653);
nor U1488 (N_1488,In_1261,In_802);
nand U1489 (N_1489,In_744,In_410);
nor U1490 (N_1490,In_1015,In_1457);
nand U1491 (N_1491,In_26,In_1030);
nor U1492 (N_1492,In_93,In_96);
nand U1493 (N_1493,In_824,In_1016);
or U1494 (N_1494,In_328,In_1487);
nor U1495 (N_1495,In_314,In_1017);
or U1496 (N_1496,In_1257,In_87);
and U1497 (N_1497,In_1314,In_1332);
nor U1498 (N_1498,In_702,In_1493);
or U1499 (N_1499,In_1499,In_573);
nand U1500 (N_1500,In_1340,In_1217);
or U1501 (N_1501,In_45,In_186);
and U1502 (N_1502,In_160,In_632);
nor U1503 (N_1503,In_143,In_1468);
and U1504 (N_1504,In_1080,In_1254);
nand U1505 (N_1505,In_1242,In_739);
or U1506 (N_1506,In_75,In_371);
nand U1507 (N_1507,In_270,In_834);
and U1508 (N_1508,In_1118,In_1419);
nand U1509 (N_1509,In_122,In_879);
or U1510 (N_1510,In_291,In_1349);
or U1511 (N_1511,In_497,In_1025);
nor U1512 (N_1512,In_934,In_286);
and U1513 (N_1513,In_274,In_642);
nand U1514 (N_1514,In_1214,In_1329);
and U1515 (N_1515,In_110,In_1303);
nor U1516 (N_1516,In_88,In_995);
and U1517 (N_1517,In_1162,In_1345);
and U1518 (N_1518,In_796,In_1424);
or U1519 (N_1519,In_509,In_525);
and U1520 (N_1520,In_630,In_1199);
and U1521 (N_1521,In_581,In_44);
and U1522 (N_1522,In_178,In_1261);
or U1523 (N_1523,In_591,In_1437);
or U1524 (N_1524,In_257,In_955);
nand U1525 (N_1525,In_1272,In_39);
nor U1526 (N_1526,In_997,In_61);
xor U1527 (N_1527,In_278,In_787);
or U1528 (N_1528,In_1256,In_426);
nand U1529 (N_1529,In_1141,In_1367);
nor U1530 (N_1530,In_1266,In_496);
nor U1531 (N_1531,In_186,In_1060);
xnor U1532 (N_1532,In_1016,In_375);
nand U1533 (N_1533,In_869,In_889);
nor U1534 (N_1534,In_381,In_1045);
and U1535 (N_1535,In_481,In_991);
nor U1536 (N_1536,In_247,In_1072);
and U1537 (N_1537,In_58,In_499);
and U1538 (N_1538,In_353,In_815);
nand U1539 (N_1539,In_1141,In_1238);
and U1540 (N_1540,In_662,In_1437);
or U1541 (N_1541,In_521,In_775);
or U1542 (N_1542,In_504,In_1082);
nand U1543 (N_1543,In_204,In_236);
nand U1544 (N_1544,In_1249,In_1052);
nor U1545 (N_1545,In_6,In_1208);
nand U1546 (N_1546,In_1078,In_559);
nand U1547 (N_1547,In_1400,In_344);
and U1548 (N_1548,In_1277,In_171);
nor U1549 (N_1549,In_761,In_281);
or U1550 (N_1550,In_1316,In_46);
nand U1551 (N_1551,In_1134,In_1426);
or U1552 (N_1552,In_274,In_1184);
nor U1553 (N_1553,In_590,In_282);
or U1554 (N_1554,In_1022,In_1117);
or U1555 (N_1555,In_792,In_310);
nor U1556 (N_1556,In_970,In_1207);
or U1557 (N_1557,In_44,In_625);
and U1558 (N_1558,In_453,In_1394);
and U1559 (N_1559,In_1310,In_827);
or U1560 (N_1560,In_1457,In_328);
or U1561 (N_1561,In_267,In_1113);
or U1562 (N_1562,In_434,In_1086);
and U1563 (N_1563,In_46,In_1022);
nor U1564 (N_1564,In_1158,In_534);
nand U1565 (N_1565,In_566,In_1298);
nand U1566 (N_1566,In_1191,In_566);
nand U1567 (N_1567,In_21,In_569);
nor U1568 (N_1568,In_1067,In_822);
or U1569 (N_1569,In_1205,In_628);
and U1570 (N_1570,In_1116,In_539);
or U1571 (N_1571,In_41,In_654);
nor U1572 (N_1572,In_989,In_388);
and U1573 (N_1573,In_74,In_1019);
or U1574 (N_1574,In_1000,In_813);
nor U1575 (N_1575,In_412,In_851);
nand U1576 (N_1576,In_284,In_546);
nor U1577 (N_1577,In_168,In_91);
and U1578 (N_1578,In_1040,In_1386);
nor U1579 (N_1579,In_19,In_444);
or U1580 (N_1580,In_569,In_671);
or U1581 (N_1581,In_1417,In_817);
or U1582 (N_1582,In_320,In_809);
or U1583 (N_1583,In_405,In_879);
nor U1584 (N_1584,In_598,In_1070);
nand U1585 (N_1585,In_1315,In_395);
or U1586 (N_1586,In_282,In_1092);
nor U1587 (N_1587,In_1178,In_123);
nand U1588 (N_1588,In_2,In_901);
nor U1589 (N_1589,In_1227,In_193);
nand U1590 (N_1590,In_799,In_377);
xor U1591 (N_1591,In_898,In_1182);
and U1592 (N_1592,In_472,In_164);
nor U1593 (N_1593,In_477,In_1236);
nand U1594 (N_1594,In_171,In_257);
nor U1595 (N_1595,In_14,In_260);
nor U1596 (N_1596,In_698,In_767);
or U1597 (N_1597,In_905,In_1328);
nand U1598 (N_1598,In_713,In_922);
or U1599 (N_1599,In_619,In_1221);
and U1600 (N_1600,In_1287,In_1281);
and U1601 (N_1601,In_1120,In_1256);
nor U1602 (N_1602,In_237,In_733);
or U1603 (N_1603,In_1147,In_375);
and U1604 (N_1604,In_503,In_873);
xnor U1605 (N_1605,In_1219,In_592);
nor U1606 (N_1606,In_514,In_421);
or U1607 (N_1607,In_1126,In_737);
nor U1608 (N_1608,In_78,In_1042);
nand U1609 (N_1609,In_1484,In_1128);
nor U1610 (N_1610,In_461,In_78);
nor U1611 (N_1611,In_1140,In_425);
nand U1612 (N_1612,In_577,In_447);
or U1613 (N_1613,In_112,In_1078);
nand U1614 (N_1614,In_235,In_649);
and U1615 (N_1615,In_1222,In_591);
and U1616 (N_1616,In_129,In_257);
nor U1617 (N_1617,In_944,In_864);
and U1618 (N_1618,In_679,In_132);
or U1619 (N_1619,In_1020,In_992);
nand U1620 (N_1620,In_1295,In_674);
nor U1621 (N_1621,In_728,In_765);
xor U1622 (N_1622,In_26,In_1088);
or U1623 (N_1623,In_1150,In_751);
and U1624 (N_1624,In_1116,In_1436);
nand U1625 (N_1625,In_411,In_568);
nand U1626 (N_1626,In_819,In_1328);
and U1627 (N_1627,In_1051,In_234);
nand U1628 (N_1628,In_277,In_100);
or U1629 (N_1629,In_69,In_180);
xor U1630 (N_1630,In_495,In_579);
nor U1631 (N_1631,In_595,In_762);
nor U1632 (N_1632,In_634,In_1484);
or U1633 (N_1633,In_1478,In_360);
or U1634 (N_1634,In_868,In_1143);
and U1635 (N_1635,In_1449,In_1400);
nand U1636 (N_1636,In_335,In_498);
nand U1637 (N_1637,In_1319,In_411);
nor U1638 (N_1638,In_1151,In_11);
nor U1639 (N_1639,In_605,In_1252);
nand U1640 (N_1640,In_774,In_1177);
nand U1641 (N_1641,In_616,In_1377);
nand U1642 (N_1642,In_412,In_402);
nand U1643 (N_1643,In_1483,In_99);
or U1644 (N_1644,In_262,In_1256);
nand U1645 (N_1645,In_800,In_1387);
or U1646 (N_1646,In_1385,In_37);
or U1647 (N_1647,In_501,In_1127);
and U1648 (N_1648,In_716,In_1169);
or U1649 (N_1649,In_218,In_1188);
nor U1650 (N_1650,In_351,In_1054);
nand U1651 (N_1651,In_157,In_703);
or U1652 (N_1652,In_1322,In_957);
or U1653 (N_1653,In_80,In_225);
and U1654 (N_1654,In_244,In_819);
nor U1655 (N_1655,In_1473,In_577);
nor U1656 (N_1656,In_558,In_586);
and U1657 (N_1657,In_318,In_1246);
and U1658 (N_1658,In_147,In_1404);
nor U1659 (N_1659,In_184,In_760);
nor U1660 (N_1660,In_1288,In_1032);
nor U1661 (N_1661,In_1099,In_1130);
and U1662 (N_1662,In_435,In_1081);
nor U1663 (N_1663,In_974,In_792);
and U1664 (N_1664,In_817,In_380);
nand U1665 (N_1665,In_956,In_504);
and U1666 (N_1666,In_243,In_1349);
nor U1667 (N_1667,In_325,In_595);
or U1668 (N_1668,In_366,In_489);
nand U1669 (N_1669,In_941,In_275);
and U1670 (N_1670,In_300,In_1129);
nor U1671 (N_1671,In_870,In_1206);
or U1672 (N_1672,In_87,In_1453);
and U1673 (N_1673,In_1444,In_1494);
nand U1674 (N_1674,In_324,In_1256);
nor U1675 (N_1675,In_1063,In_1062);
nand U1676 (N_1676,In_343,In_747);
and U1677 (N_1677,In_659,In_879);
nand U1678 (N_1678,In_1458,In_793);
nor U1679 (N_1679,In_312,In_1298);
nand U1680 (N_1680,In_671,In_24);
or U1681 (N_1681,In_1214,In_1437);
and U1682 (N_1682,In_1357,In_900);
nand U1683 (N_1683,In_381,In_27);
and U1684 (N_1684,In_1188,In_812);
or U1685 (N_1685,In_231,In_1146);
nand U1686 (N_1686,In_885,In_380);
nor U1687 (N_1687,In_1187,In_383);
nor U1688 (N_1688,In_406,In_232);
nor U1689 (N_1689,In_1135,In_1225);
nand U1690 (N_1690,In_486,In_582);
and U1691 (N_1691,In_136,In_1379);
nand U1692 (N_1692,In_977,In_860);
nor U1693 (N_1693,In_443,In_378);
or U1694 (N_1694,In_666,In_1201);
nor U1695 (N_1695,In_53,In_985);
nor U1696 (N_1696,In_1192,In_156);
nand U1697 (N_1697,In_658,In_248);
and U1698 (N_1698,In_1462,In_1098);
or U1699 (N_1699,In_764,In_868);
and U1700 (N_1700,In_1324,In_879);
or U1701 (N_1701,In_822,In_640);
and U1702 (N_1702,In_575,In_307);
or U1703 (N_1703,In_1188,In_842);
nor U1704 (N_1704,In_1378,In_1425);
nor U1705 (N_1705,In_94,In_826);
nor U1706 (N_1706,In_263,In_984);
and U1707 (N_1707,In_339,In_386);
nand U1708 (N_1708,In_1353,In_745);
nand U1709 (N_1709,In_312,In_188);
nor U1710 (N_1710,In_352,In_24);
and U1711 (N_1711,In_563,In_1127);
and U1712 (N_1712,In_730,In_495);
or U1713 (N_1713,In_501,In_1334);
and U1714 (N_1714,In_292,In_1295);
or U1715 (N_1715,In_168,In_1229);
nand U1716 (N_1716,In_926,In_638);
nand U1717 (N_1717,In_525,In_711);
or U1718 (N_1718,In_1411,In_201);
nand U1719 (N_1719,In_538,In_1005);
and U1720 (N_1720,In_23,In_7);
xnor U1721 (N_1721,In_909,In_390);
nor U1722 (N_1722,In_1053,In_158);
nor U1723 (N_1723,In_613,In_353);
and U1724 (N_1724,In_573,In_523);
nand U1725 (N_1725,In_1287,In_1260);
nand U1726 (N_1726,In_175,In_874);
nand U1727 (N_1727,In_256,In_157);
nand U1728 (N_1728,In_185,In_1358);
or U1729 (N_1729,In_1054,In_1356);
nand U1730 (N_1730,In_452,In_451);
nand U1731 (N_1731,In_315,In_537);
nand U1732 (N_1732,In_274,In_260);
and U1733 (N_1733,In_1064,In_642);
nor U1734 (N_1734,In_1312,In_1440);
and U1735 (N_1735,In_1432,In_1113);
xnor U1736 (N_1736,In_690,In_286);
and U1737 (N_1737,In_1224,In_349);
nor U1738 (N_1738,In_624,In_1032);
and U1739 (N_1739,In_779,In_1013);
nand U1740 (N_1740,In_1346,In_780);
or U1741 (N_1741,In_319,In_69);
nand U1742 (N_1742,In_113,In_11);
nand U1743 (N_1743,In_414,In_479);
nor U1744 (N_1744,In_1132,In_193);
and U1745 (N_1745,In_455,In_1214);
or U1746 (N_1746,In_199,In_1027);
or U1747 (N_1747,In_372,In_890);
nand U1748 (N_1748,In_696,In_1331);
nor U1749 (N_1749,In_1181,In_1019);
nand U1750 (N_1750,In_960,In_1229);
nor U1751 (N_1751,In_1391,In_814);
or U1752 (N_1752,In_813,In_884);
or U1753 (N_1753,In_1409,In_906);
and U1754 (N_1754,In_272,In_1492);
nand U1755 (N_1755,In_1230,In_643);
nand U1756 (N_1756,In_599,In_1396);
or U1757 (N_1757,In_485,In_184);
and U1758 (N_1758,In_756,In_179);
nand U1759 (N_1759,In_1492,In_418);
nor U1760 (N_1760,In_298,In_224);
nor U1761 (N_1761,In_656,In_941);
nand U1762 (N_1762,In_76,In_910);
nor U1763 (N_1763,In_950,In_544);
or U1764 (N_1764,In_288,In_439);
xnor U1765 (N_1765,In_1361,In_213);
or U1766 (N_1766,In_411,In_1000);
or U1767 (N_1767,In_1190,In_251);
and U1768 (N_1768,In_410,In_779);
or U1769 (N_1769,In_1384,In_53);
nor U1770 (N_1770,In_441,In_884);
nor U1771 (N_1771,In_511,In_190);
or U1772 (N_1772,In_638,In_677);
nand U1773 (N_1773,In_134,In_1383);
or U1774 (N_1774,In_621,In_567);
or U1775 (N_1775,In_846,In_410);
nor U1776 (N_1776,In_1120,In_1346);
nand U1777 (N_1777,In_1496,In_1090);
nand U1778 (N_1778,In_226,In_780);
or U1779 (N_1779,In_1298,In_268);
or U1780 (N_1780,In_677,In_907);
nand U1781 (N_1781,In_1021,In_1296);
or U1782 (N_1782,In_1116,In_400);
nor U1783 (N_1783,In_55,In_993);
or U1784 (N_1784,In_639,In_443);
nor U1785 (N_1785,In_848,In_1140);
or U1786 (N_1786,In_105,In_1201);
xnor U1787 (N_1787,In_1054,In_276);
or U1788 (N_1788,In_911,In_689);
and U1789 (N_1789,In_1316,In_128);
nor U1790 (N_1790,In_382,In_701);
nand U1791 (N_1791,In_671,In_817);
or U1792 (N_1792,In_1388,In_1347);
nand U1793 (N_1793,In_789,In_768);
nor U1794 (N_1794,In_1146,In_25);
nor U1795 (N_1795,In_429,In_295);
nor U1796 (N_1796,In_424,In_529);
or U1797 (N_1797,In_210,In_950);
or U1798 (N_1798,In_633,In_1043);
and U1799 (N_1799,In_1007,In_520);
nor U1800 (N_1800,In_1184,In_373);
and U1801 (N_1801,In_470,In_480);
nand U1802 (N_1802,In_1248,In_882);
nor U1803 (N_1803,In_82,In_1096);
nand U1804 (N_1804,In_1255,In_697);
or U1805 (N_1805,In_122,In_126);
and U1806 (N_1806,In_941,In_1484);
and U1807 (N_1807,In_1173,In_245);
and U1808 (N_1808,In_248,In_1073);
nor U1809 (N_1809,In_1057,In_1352);
or U1810 (N_1810,In_180,In_585);
nand U1811 (N_1811,In_298,In_1306);
or U1812 (N_1812,In_1003,In_880);
nand U1813 (N_1813,In_1093,In_770);
and U1814 (N_1814,In_202,In_35);
nand U1815 (N_1815,In_1404,In_936);
nand U1816 (N_1816,In_335,In_36);
and U1817 (N_1817,In_1000,In_938);
nand U1818 (N_1818,In_784,In_365);
or U1819 (N_1819,In_692,In_1388);
nand U1820 (N_1820,In_1169,In_1017);
nor U1821 (N_1821,In_1141,In_909);
xor U1822 (N_1822,In_712,In_1220);
and U1823 (N_1823,In_917,In_511);
nand U1824 (N_1824,In_161,In_129);
and U1825 (N_1825,In_10,In_1378);
or U1826 (N_1826,In_553,In_321);
and U1827 (N_1827,In_597,In_996);
nor U1828 (N_1828,In_698,In_1416);
or U1829 (N_1829,In_1497,In_290);
nand U1830 (N_1830,In_906,In_234);
and U1831 (N_1831,In_170,In_951);
nor U1832 (N_1832,In_66,In_1352);
nand U1833 (N_1833,In_1005,In_243);
or U1834 (N_1834,In_467,In_1433);
nor U1835 (N_1835,In_142,In_1032);
or U1836 (N_1836,In_1287,In_1454);
nand U1837 (N_1837,In_535,In_100);
nor U1838 (N_1838,In_827,In_40);
nand U1839 (N_1839,In_197,In_828);
and U1840 (N_1840,In_891,In_740);
nor U1841 (N_1841,In_1260,In_186);
and U1842 (N_1842,In_129,In_287);
or U1843 (N_1843,In_369,In_1374);
and U1844 (N_1844,In_815,In_1249);
and U1845 (N_1845,In_1039,In_443);
nor U1846 (N_1846,In_324,In_801);
nand U1847 (N_1847,In_636,In_321);
and U1848 (N_1848,In_625,In_1220);
nand U1849 (N_1849,In_1133,In_583);
or U1850 (N_1850,In_1492,In_680);
nand U1851 (N_1851,In_1142,In_375);
nand U1852 (N_1852,In_598,In_1413);
and U1853 (N_1853,In_669,In_750);
and U1854 (N_1854,In_301,In_1229);
nand U1855 (N_1855,In_201,In_304);
nor U1856 (N_1856,In_14,In_705);
or U1857 (N_1857,In_814,In_1268);
nand U1858 (N_1858,In_2,In_291);
nand U1859 (N_1859,In_1410,In_911);
nand U1860 (N_1860,In_865,In_552);
nor U1861 (N_1861,In_476,In_811);
and U1862 (N_1862,In_968,In_1082);
nor U1863 (N_1863,In_1031,In_285);
nand U1864 (N_1864,In_1037,In_1196);
or U1865 (N_1865,In_338,In_1405);
nand U1866 (N_1866,In_596,In_658);
nand U1867 (N_1867,In_776,In_463);
or U1868 (N_1868,In_330,In_1028);
nand U1869 (N_1869,In_55,In_1092);
nor U1870 (N_1870,In_1256,In_916);
and U1871 (N_1871,In_798,In_217);
nor U1872 (N_1872,In_1032,In_593);
or U1873 (N_1873,In_609,In_917);
and U1874 (N_1874,In_1212,In_526);
nand U1875 (N_1875,In_306,In_78);
nand U1876 (N_1876,In_518,In_1);
and U1877 (N_1877,In_1382,In_160);
and U1878 (N_1878,In_1042,In_566);
nor U1879 (N_1879,In_256,In_483);
or U1880 (N_1880,In_971,In_1355);
or U1881 (N_1881,In_1245,In_1143);
and U1882 (N_1882,In_1430,In_1452);
nor U1883 (N_1883,In_110,In_1278);
nor U1884 (N_1884,In_1056,In_769);
or U1885 (N_1885,In_974,In_772);
nor U1886 (N_1886,In_558,In_1138);
and U1887 (N_1887,In_303,In_478);
nor U1888 (N_1888,In_1285,In_632);
and U1889 (N_1889,In_771,In_1454);
and U1890 (N_1890,In_396,In_374);
and U1891 (N_1891,In_955,In_947);
nor U1892 (N_1892,In_1419,In_195);
and U1893 (N_1893,In_1158,In_398);
or U1894 (N_1894,In_594,In_161);
and U1895 (N_1895,In_326,In_918);
nor U1896 (N_1896,In_1046,In_1236);
and U1897 (N_1897,In_451,In_1132);
nor U1898 (N_1898,In_897,In_909);
nand U1899 (N_1899,In_538,In_1001);
or U1900 (N_1900,In_1322,In_511);
nand U1901 (N_1901,In_410,In_1381);
and U1902 (N_1902,In_378,In_1107);
nand U1903 (N_1903,In_924,In_679);
nor U1904 (N_1904,In_785,In_491);
and U1905 (N_1905,In_1212,In_1219);
or U1906 (N_1906,In_1302,In_355);
nand U1907 (N_1907,In_253,In_1387);
and U1908 (N_1908,In_1236,In_342);
nand U1909 (N_1909,In_1235,In_1213);
nor U1910 (N_1910,In_1143,In_1161);
and U1911 (N_1911,In_1387,In_694);
nand U1912 (N_1912,In_456,In_952);
nand U1913 (N_1913,In_574,In_1238);
nor U1914 (N_1914,In_1033,In_1031);
nand U1915 (N_1915,In_922,In_898);
nor U1916 (N_1916,In_1375,In_1472);
nand U1917 (N_1917,In_1156,In_847);
or U1918 (N_1918,In_259,In_50);
nor U1919 (N_1919,In_708,In_984);
nand U1920 (N_1920,In_1067,In_765);
and U1921 (N_1921,In_881,In_1454);
nand U1922 (N_1922,In_657,In_1282);
nor U1923 (N_1923,In_226,In_1190);
nor U1924 (N_1924,In_634,In_402);
nor U1925 (N_1925,In_1369,In_1189);
nor U1926 (N_1926,In_505,In_18);
and U1927 (N_1927,In_1411,In_1227);
nor U1928 (N_1928,In_80,In_645);
nor U1929 (N_1929,In_1480,In_1065);
nor U1930 (N_1930,In_641,In_183);
xor U1931 (N_1931,In_1498,In_1008);
or U1932 (N_1932,In_629,In_163);
nor U1933 (N_1933,In_104,In_1030);
nor U1934 (N_1934,In_1208,In_836);
nor U1935 (N_1935,In_282,In_24);
or U1936 (N_1936,In_462,In_61);
and U1937 (N_1937,In_843,In_122);
nand U1938 (N_1938,In_1087,In_495);
and U1939 (N_1939,In_44,In_1178);
nand U1940 (N_1940,In_846,In_111);
and U1941 (N_1941,In_7,In_511);
and U1942 (N_1942,In_665,In_430);
or U1943 (N_1943,In_1390,In_705);
or U1944 (N_1944,In_982,In_7);
nor U1945 (N_1945,In_1273,In_579);
or U1946 (N_1946,In_1430,In_1432);
nand U1947 (N_1947,In_1221,In_1400);
and U1948 (N_1948,In_472,In_781);
nor U1949 (N_1949,In_960,In_917);
and U1950 (N_1950,In_675,In_998);
nor U1951 (N_1951,In_1490,In_84);
nor U1952 (N_1952,In_22,In_567);
nand U1953 (N_1953,In_55,In_533);
nor U1954 (N_1954,In_422,In_600);
nor U1955 (N_1955,In_1271,In_1431);
or U1956 (N_1956,In_440,In_931);
and U1957 (N_1957,In_1382,In_746);
nor U1958 (N_1958,In_545,In_652);
nor U1959 (N_1959,In_1084,In_749);
xnor U1960 (N_1960,In_983,In_529);
xnor U1961 (N_1961,In_392,In_1125);
nor U1962 (N_1962,In_928,In_695);
and U1963 (N_1963,In_251,In_469);
nand U1964 (N_1964,In_1143,In_582);
nor U1965 (N_1965,In_1489,In_913);
nand U1966 (N_1966,In_268,In_1077);
or U1967 (N_1967,In_1285,In_253);
nor U1968 (N_1968,In_1396,In_127);
and U1969 (N_1969,In_21,In_1096);
or U1970 (N_1970,In_680,In_874);
or U1971 (N_1971,In_1164,In_1022);
nand U1972 (N_1972,In_498,In_1368);
nand U1973 (N_1973,In_627,In_413);
nor U1974 (N_1974,In_1350,In_629);
or U1975 (N_1975,In_949,In_56);
and U1976 (N_1976,In_488,In_707);
nor U1977 (N_1977,In_253,In_1421);
and U1978 (N_1978,In_458,In_691);
nand U1979 (N_1979,In_86,In_474);
xnor U1980 (N_1980,In_377,In_441);
and U1981 (N_1981,In_1494,In_914);
nor U1982 (N_1982,In_76,In_391);
nand U1983 (N_1983,In_1456,In_616);
and U1984 (N_1984,In_1263,In_82);
nor U1985 (N_1985,In_11,In_39);
or U1986 (N_1986,In_730,In_1175);
nor U1987 (N_1987,In_1003,In_1004);
and U1988 (N_1988,In_539,In_166);
nand U1989 (N_1989,In_1253,In_61);
and U1990 (N_1990,In_1115,In_916);
and U1991 (N_1991,In_1373,In_1470);
nand U1992 (N_1992,In_11,In_1333);
and U1993 (N_1993,In_1150,In_1333);
or U1994 (N_1994,In_621,In_1254);
nor U1995 (N_1995,In_401,In_361);
or U1996 (N_1996,In_1317,In_1068);
nand U1997 (N_1997,In_1120,In_1008);
nand U1998 (N_1998,In_603,In_685);
nor U1999 (N_1999,In_1195,In_321);
nand U2000 (N_2000,In_263,In_793);
or U2001 (N_2001,In_1259,In_385);
or U2002 (N_2002,In_160,In_1466);
or U2003 (N_2003,In_1249,In_1221);
nor U2004 (N_2004,In_1190,In_746);
nand U2005 (N_2005,In_724,In_121);
or U2006 (N_2006,In_585,In_874);
nand U2007 (N_2007,In_998,In_1051);
nor U2008 (N_2008,In_180,In_288);
nand U2009 (N_2009,In_140,In_531);
or U2010 (N_2010,In_1381,In_788);
or U2011 (N_2011,In_685,In_212);
nand U2012 (N_2012,In_155,In_147);
and U2013 (N_2013,In_863,In_1374);
or U2014 (N_2014,In_278,In_412);
or U2015 (N_2015,In_51,In_967);
nand U2016 (N_2016,In_268,In_1208);
nand U2017 (N_2017,In_830,In_723);
nand U2018 (N_2018,In_1391,In_1384);
and U2019 (N_2019,In_404,In_1426);
nor U2020 (N_2020,In_888,In_29);
nor U2021 (N_2021,In_207,In_585);
and U2022 (N_2022,In_879,In_490);
xor U2023 (N_2023,In_412,In_1200);
nor U2024 (N_2024,In_1430,In_782);
nor U2025 (N_2025,In_811,In_202);
or U2026 (N_2026,In_1226,In_1352);
nand U2027 (N_2027,In_651,In_1332);
nor U2028 (N_2028,In_1298,In_802);
and U2029 (N_2029,In_1121,In_56);
or U2030 (N_2030,In_1339,In_399);
and U2031 (N_2031,In_910,In_116);
nor U2032 (N_2032,In_163,In_1273);
nor U2033 (N_2033,In_1037,In_1478);
nor U2034 (N_2034,In_1386,In_1464);
nand U2035 (N_2035,In_901,In_153);
and U2036 (N_2036,In_117,In_629);
nand U2037 (N_2037,In_1278,In_438);
and U2038 (N_2038,In_98,In_1157);
and U2039 (N_2039,In_300,In_598);
and U2040 (N_2040,In_755,In_46);
nor U2041 (N_2041,In_967,In_624);
nor U2042 (N_2042,In_1449,In_754);
nor U2043 (N_2043,In_282,In_389);
and U2044 (N_2044,In_1449,In_1477);
nor U2045 (N_2045,In_89,In_232);
nor U2046 (N_2046,In_431,In_981);
nor U2047 (N_2047,In_1421,In_427);
and U2048 (N_2048,In_582,In_673);
nor U2049 (N_2049,In_539,In_754);
or U2050 (N_2050,In_667,In_1393);
or U2051 (N_2051,In_1336,In_943);
xor U2052 (N_2052,In_1027,In_1033);
and U2053 (N_2053,In_845,In_1406);
or U2054 (N_2054,In_1336,In_1181);
nand U2055 (N_2055,In_1407,In_453);
or U2056 (N_2056,In_9,In_506);
nor U2057 (N_2057,In_447,In_236);
and U2058 (N_2058,In_574,In_129);
nand U2059 (N_2059,In_160,In_486);
or U2060 (N_2060,In_850,In_876);
or U2061 (N_2061,In_71,In_467);
or U2062 (N_2062,In_956,In_1261);
or U2063 (N_2063,In_1263,In_375);
or U2064 (N_2064,In_497,In_924);
or U2065 (N_2065,In_855,In_858);
and U2066 (N_2066,In_784,In_1379);
nor U2067 (N_2067,In_1402,In_1459);
nor U2068 (N_2068,In_1273,In_136);
nand U2069 (N_2069,In_567,In_1127);
or U2070 (N_2070,In_49,In_557);
or U2071 (N_2071,In_1416,In_1107);
nand U2072 (N_2072,In_651,In_1319);
or U2073 (N_2073,In_1389,In_61);
nor U2074 (N_2074,In_957,In_1269);
or U2075 (N_2075,In_1001,In_498);
nand U2076 (N_2076,In_1235,In_132);
nor U2077 (N_2077,In_124,In_1133);
xnor U2078 (N_2078,In_1181,In_661);
nor U2079 (N_2079,In_732,In_1114);
nor U2080 (N_2080,In_9,In_274);
or U2081 (N_2081,In_1137,In_1031);
nor U2082 (N_2082,In_665,In_783);
or U2083 (N_2083,In_96,In_968);
or U2084 (N_2084,In_587,In_594);
nand U2085 (N_2085,In_821,In_928);
or U2086 (N_2086,In_1350,In_1177);
nand U2087 (N_2087,In_572,In_1424);
or U2088 (N_2088,In_1478,In_1196);
or U2089 (N_2089,In_1170,In_1400);
or U2090 (N_2090,In_1193,In_1119);
or U2091 (N_2091,In_1017,In_1469);
nand U2092 (N_2092,In_937,In_1321);
nor U2093 (N_2093,In_952,In_1384);
or U2094 (N_2094,In_1070,In_1133);
and U2095 (N_2095,In_738,In_22);
or U2096 (N_2096,In_564,In_67);
or U2097 (N_2097,In_1354,In_732);
nor U2098 (N_2098,In_1233,In_929);
nand U2099 (N_2099,In_140,In_352);
nor U2100 (N_2100,In_1361,In_1332);
or U2101 (N_2101,In_981,In_1411);
and U2102 (N_2102,In_973,In_904);
and U2103 (N_2103,In_471,In_1129);
nor U2104 (N_2104,In_348,In_90);
or U2105 (N_2105,In_225,In_922);
or U2106 (N_2106,In_1,In_1064);
nand U2107 (N_2107,In_613,In_950);
nor U2108 (N_2108,In_885,In_150);
or U2109 (N_2109,In_1327,In_842);
or U2110 (N_2110,In_130,In_800);
and U2111 (N_2111,In_551,In_69);
and U2112 (N_2112,In_1419,In_288);
and U2113 (N_2113,In_341,In_1438);
and U2114 (N_2114,In_550,In_1340);
and U2115 (N_2115,In_1339,In_525);
or U2116 (N_2116,In_601,In_413);
nand U2117 (N_2117,In_882,In_58);
and U2118 (N_2118,In_608,In_670);
or U2119 (N_2119,In_653,In_1232);
or U2120 (N_2120,In_1070,In_924);
nor U2121 (N_2121,In_1355,In_1354);
nor U2122 (N_2122,In_828,In_824);
or U2123 (N_2123,In_1010,In_123);
nor U2124 (N_2124,In_285,In_1047);
and U2125 (N_2125,In_811,In_973);
nand U2126 (N_2126,In_1165,In_699);
nor U2127 (N_2127,In_441,In_760);
or U2128 (N_2128,In_1028,In_1248);
or U2129 (N_2129,In_0,In_154);
or U2130 (N_2130,In_1363,In_1193);
xor U2131 (N_2131,In_87,In_1122);
nand U2132 (N_2132,In_724,In_444);
or U2133 (N_2133,In_4,In_98);
nand U2134 (N_2134,In_808,In_323);
or U2135 (N_2135,In_84,In_1351);
or U2136 (N_2136,In_1433,In_1111);
nor U2137 (N_2137,In_1097,In_36);
or U2138 (N_2138,In_456,In_1442);
or U2139 (N_2139,In_186,In_838);
or U2140 (N_2140,In_836,In_1377);
nor U2141 (N_2141,In_797,In_45);
or U2142 (N_2142,In_964,In_626);
nor U2143 (N_2143,In_1339,In_453);
and U2144 (N_2144,In_414,In_664);
nor U2145 (N_2145,In_740,In_1223);
nor U2146 (N_2146,In_1078,In_588);
or U2147 (N_2147,In_493,In_1451);
and U2148 (N_2148,In_745,In_907);
or U2149 (N_2149,In_49,In_50);
and U2150 (N_2150,In_965,In_691);
nand U2151 (N_2151,In_249,In_250);
nor U2152 (N_2152,In_1240,In_1326);
nand U2153 (N_2153,In_1033,In_991);
and U2154 (N_2154,In_1307,In_1046);
and U2155 (N_2155,In_1330,In_424);
nor U2156 (N_2156,In_589,In_688);
and U2157 (N_2157,In_67,In_908);
nor U2158 (N_2158,In_85,In_1313);
nand U2159 (N_2159,In_0,In_1121);
nand U2160 (N_2160,In_146,In_317);
nand U2161 (N_2161,In_1012,In_755);
nand U2162 (N_2162,In_17,In_505);
or U2163 (N_2163,In_1342,In_230);
or U2164 (N_2164,In_1437,In_1122);
nor U2165 (N_2165,In_200,In_890);
and U2166 (N_2166,In_1073,In_987);
or U2167 (N_2167,In_1273,In_424);
or U2168 (N_2168,In_166,In_512);
nor U2169 (N_2169,In_799,In_516);
nor U2170 (N_2170,In_1084,In_321);
nand U2171 (N_2171,In_486,In_589);
or U2172 (N_2172,In_134,In_966);
and U2173 (N_2173,In_311,In_1022);
nor U2174 (N_2174,In_35,In_145);
nor U2175 (N_2175,In_1319,In_330);
and U2176 (N_2176,In_456,In_689);
xnor U2177 (N_2177,In_1449,In_1033);
and U2178 (N_2178,In_430,In_974);
and U2179 (N_2179,In_975,In_795);
nor U2180 (N_2180,In_902,In_694);
and U2181 (N_2181,In_599,In_349);
and U2182 (N_2182,In_277,In_1082);
and U2183 (N_2183,In_1363,In_920);
nand U2184 (N_2184,In_941,In_1046);
or U2185 (N_2185,In_1447,In_514);
nand U2186 (N_2186,In_259,In_765);
nor U2187 (N_2187,In_949,In_398);
nand U2188 (N_2188,In_1364,In_154);
nand U2189 (N_2189,In_960,In_194);
nor U2190 (N_2190,In_881,In_765);
or U2191 (N_2191,In_1001,In_830);
xor U2192 (N_2192,In_1168,In_556);
or U2193 (N_2193,In_284,In_1382);
nand U2194 (N_2194,In_1484,In_917);
nor U2195 (N_2195,In_865,In_495);
or U2196 (N_2196,In_1089,In_1338);
or U2197 (N_2197,In_855,In_1427);
and U2198 (N_2198,In_1478,In_305);
nor U2199 (N_2199,In_166,In_190);
nor U2200 (N_2200,In_868,In_636);
and U2201 (N_2201,In_1339,In_890);
nand U2202 (N_2202,In_1334,In_1051);
nor U2203 (N_2203,In_1378,In_584);
nand U2204 (N_2204,In_1238,In_1290);
and U2205 (N_2205,In_801,In_1381);
nor U2206 (N_2206,In_1498,In_1442);
nand U2207 (N_2207,In_168,In_950);
and U2208 (N_2208,In_1070,In_407);
or U2209 (N_2209,In_852,In_591);
and U2210 (N_2210,In_1006,In_961);
nor U2211 (N_2211,In_1190,In_722);
and U2212 (N_2212,In_789,In_438);
nand U2213 (N_2213,In_521,In_1243);
nand U2214 (N_2214,In_1360,In_1121);
nand U2215 (N_2215,In_202,In_1463);
nand U2216 (N_2216,In_1195,In_521);
nor U2217 (N_2217,In_687,In_135);
nor U2218 (N_2218,In_1175,In_995);
or U2219 (N_2219,In_887,In_1108);
or U2220 (N_2220,In_1061,In_486);
nor U2221 (N_2221,In_35,In_648);
or U2222 (N_2222,In_1322,In_896);
and U2223 (N_2223,In_1315,In_1080);
or U2224 (N_2224,In_354,In_1184);
or U2225 (N_2225,In_1387,In_834);
nor U2226 (N_2226,In_382,In_632);
nand U2227 (N_2227,In_711,In_224);
nor U2228 (N_2228,In_1118,In_905);
or U2229 (N_2229,In_1301,In_1245);
or U2230 (N_2230,In_826,In_339);
xnor U2231 (N_2231,In_638,In_1423);
nor U2232 (N_2232,In_1020,In_420);
and U2233 (N_2233,In_828,In_1063);
or U2234 (N_2234,In_1024,In_600);
nand U2235 (N_2235,In_1422,In_874);
nand U2236 (N_2236,In_582,In_31);
nor U2237 (N_2237,In_243,In_1008);
nor U2238 (N_2238,In_1173,In_872);
nor U2239 (N_2239,In_590,In_1103);
and U2240 (N_2240,In_564,In_93);
and U2241 (N_2241,In_1194,In_1286);
nor U2242 (N_2242,In_582,In_931);
nor U2243 (N_2243,In_725,In_1084);
or U2244 (N_2244,In_1222,In_1191);
nor U2245 (N_2245,In_1392,In_171);
or U2246 (N_2246,In_616,In_87);
nor U2247 (N_2247,In_216,In_438);
nand U2248 (N_2248,In_533,In_270);
nor U2249 (N_2249,In_1007,In_240);
and U2250 (N_2250,In_1009,In_517);
and U2251 (N_2251,In_498,In_1453);
nor U2252 (N_2252,In_397,In_250);
and U2253 (N_2253,In_188,In_164);
nand U2254 (N_2254,In_622,In_424);
nor U2255 (N_2255,In_1361,In_886);
nor U2256 (N_2256,In_925,In_921);
nor U2257 (N_2257,In_989,In_829);
and U2258 (N_2258,In_1280,In_109);
or U2259 (N_2259,In_260,In_346);
and U2260 (N_2260,In_62,In_971);
nand U2261 (N_2261,In_1287,In_730);
nor U2262 (N_2262,In_318,In_1301);
or U2263 (N_2263,In_1,In_981);
nor U2264 (N_2264,In_705,In_721);
or U2265 (N_2265,In_1084,In_1255);
or U2266 (N_2266,In_1160,In_272);
or U2267 (N_2267,In_506,In_1137);
nand U2268 (N_2268,In_720,In_629);
nor U2269 (N_2269,In_1121,In_17);
and U2270 (N_2270,In_471,In_1433);
nor U2271 (N_2271,In_760,In_474);
nor U2272 (N_2272,In_51,In_74);
or U2273 (N_2273,In_924,In_290);
nor U2274 (N_2274,In_1405,In_555);
nor U2275 (N_2275,In_899,In_1295);
nor U2276 (N_2276,In_641,In_892);
nand U2277 (N_2277,In_810,In_525);
nor U2278 (N_2278,In_675,In_1434);
nor U2279 (N_2279,In_760,In_172);
and U2280 (N_2280,In_1087,In_351);
and U2281 (N_2281,In_658,In_464);
nor U2282 (N_2282,In_1214,In_744);
nor U2283 (N_2283,In_1280,In_900);
or U2284 (N_2284,In_1345,In_997);
nor U2285 (N_2285,In_667,In_1387);
or U2286 (N_2286,In_113,In_869);
and U2287 (N_2287,In_163,In_990);
nand U2288 (N_2288,In_1377,In_1343);
nand U2289 (N_2289,In_106,In_1086);
nor U2290 (N_2290,In_317,In_800);
nand U2291 (N_2291,In_176,In_397);
nand U2292 (N_2292,In_1123,In_621);
or U2293 (N_2293,In_1108,In_1084);
nand U2294 (N_2294,In_898,In_168);
or U2295 (N_2295,In_780,In_973);
or U2296 (N_2296,In_65,In_1055);
or U2297 (N_2297,In_598,In_835);
or U2298 (N_2298,In_343,In_329);
and U2299 (N_2299,In_485,In_1338);
and U2300 (N_2300,In_1232,In_458);
nand U2301 (N_2301,In_830,In_31);
nor U2302 (N_2302,In_914,In_24);
xor U2303 (N_2303,In_44,In_976);
nor U2304 (N_2304,In_90,In_639);
nor U2305 (N_2305,In_1106,In_912);
and U2306 (N_2306,In_1030,In_696);
nand U2307 (N_2307,In_708,In_627);
nand U2308 (N_2308,In_669,In_812);
and U2309 (N_2309,In_52,In_857);
and U2310 (N_2310,In_969,In_1459);
or U2311 (N_2311,In_477,In_250);
nand U2312 (N_2312,In_1083,In_832);
nor U2313 (N_2313,In_321,In_762);
nand U2314 (N_2314,In_1004,In_223);
nor U2315 (N_2315,In_917,In_426);
and U2316 (N_2316,In_567,In_251);
or U2317 (N_2317,In_1412,In_90);
nor U2318 (N_2318,In_148,In_145);
or U2319 (N_2319,In_38,In_147);
or U2320 (N_2320,In_1391,In_169);
nor U2321 (N_2321,In_1371,In_1122);
nor U2322 (N_2322,In_920,In_1037);
nor U2323 (N_2323,In_886,In_15);
nor U2324 (N_2324,In_1294,In_48);
nand U2325 (N_2325,In_268,In_1305);
and U2326 (N_2326,In_559,In_869);
nand U2327 (N_2327,In_681,In_1096);
or U2328 (N_2328,In_245,In_168);
and U2329 (N_2329,In_526,In_171);
and U2330 (N_2330,In_142,In_1055);
nand U2331 (N_2331,In_877,In_17);
nor U2332 (N_2332,In_1437,In_868);
nand U2333 (N_2333,In_1018,In_130);
and U2334 (N_2334,In_277,In_330);
and U2335 (N_2335,In_1176,In_1188);
nand U2336 (N_2336,In_448,In_308);
nor U2337 (N_2337,In_700,In_280);
and U2338 (N_2338,In_594,In_835);
nor U2339 (N_2339,In_767,In_457);
or U2340 (N_2340,In_1413,In_749);
nand U2341 (N_2341,In_867,In_1282);
or U2342 (N_2342,In_988,In_187);
or U2343 (N_2343,In_405,In_1390);
nor U2344 (N_2344,In_560,In_1121);
nor U2345 (N_2345,In_742,In_752);
nand U2346 (N_2346,In_361,In_1272);
or U2347 (N_2347,In_1194,In_523);
nor U2348 (N_2348,In_1251,In_478);
nand U2349 (N_2349,In_560,In_178);
or U2350 (N_2350,In_666,In_209);
nand U2351 (N_2351,In_722,In_459);
nor U2352 (N_2352,In_621,In_357);
or U2353 (N_2353,In_59,In_1475);
and U2354 (N_2354,In_69,In_202);
nand U2355 (N_2355,In_331,In_930);
or U2356 (N_2356,In_1379,In_18);
xor U2357 (N_2357,In_1229,In_437);
and U2358 (N_2358,In_833,In_716);
nor U2359 (N_2359,In_71,In_201);
or U2360 (N_2360,In_348,In_1447);
and U2361 (N_2361,In_742,In_43);
or U2362 (N_2362,In_1178,In_817);
xor U2363 (N_2363,In_1030,In_122);
nand U2364 (N_2364,In_226,In_1239);
nand U2365 (N_2365,In_204,In_461);
xor U2366 (N_2366,In_54,In_1377);
nand U2367 (N_2367,In_182,In_919);
or U2368 (N_2368,In_1054,In_250);
and U2369 (N_2369,In_170,In_311);
and U2370 (N_2370,In_1360,In_321);
and U2371 (N_2371,In_701,In_1346);
nor U2372 (N_2372,In_622,In_233);
nor U2373 (N_2373,In_325,In_80);
and U2374 (N_2374,In_1193,In_909);
nor U2375 (N_2375,In_1354,In_1174);
nor U2376 (N_2376,In_821,In_1095);
nor U2377 (N_2377,In_733,In_856);
and U2378 (N_2378,In_676,In_1191);
or U2379 (N_2379,In_188,In_1485);
or U2380 (N_2380,In_898,In_340);
nand U2381 (N_2381,In_995,In_1410);
nor U2382 (N_2382,In_357,In_820);
or U2383 (N_2383,In_403,In_737);
or U2384 (N_2384,In_553,In_734);
nand U2385 (N_2385,In_1009,In_885);
and U2386 (N_2386,In_901,In_1402);
and U2387 (N_2387,In_1212,In_1096);
or U2388 (N_2388,In_1193,In_775);
nand U2389 (N_2389,In_264,In_600);
nor U2390 (N_2390,In_1388,In_888);
and U2391 (N_2391,In_505,In_1256);
and U2392 (N_2392,In_1408,In_160);
or U2393 (N_2393,In_239,In_51);
or U2394 (N_2394,In_197,In_3);
nand U2395 (N_2395,In_994,In_832);
nand U2396 (N_2396,In_542,In_372);
xnor U2397 (N_2397,In_1061,In_72);
or U2398 (N_2398,In_1278,In_172);
or U2399 (N_2399,In_528,In_1040);
and U2400 (N_2400,In_276,In_58);
and U2401 (N_2401,In_423,In_1450);
and U2402 (N_2402,In_633,In_48);
or U2403 (N_2403,In_399,In_23);
nand U2404 (N_2404,In_58,In_498);
nand U2405 (N_2405,In_1203,In_173);
and U2406 (N_2406,In_1423,In_328);
or U2407 (N_2407,In_1069,In_155);
nand U2408 (N_2408,In_99,In_468);
nor U2409 (N_2409,In_641,In_635);
or U2410 (N_2410,In_1124,In_1083);
nand U2411 (N_2411,In_1328,In_840);
nor U2412 (N_2412,In_1363,In_334);
nor U2413 (N_2413,In_1151,In_1424);
and U2414 (N_2414,In_196,In_691);
nand U2415 (N_2415,In_520,In_439);
and U2416 (N_2416,In_289,In_947);
nor U2417 (N_2417,In_1123,In_633);
or U2418 (N_2418,In_516,In_1333);
and U2419 (N_2419,In_1273,In_94);
or U2420 (N_2420,In_370,In_573);
nor U2421 (N_2421,In_622,In_846);
nor U2422 (N_2422,In_624,In_1424);
nand U2423 (N_2423,In_1093,In_1277);
nand U2424 (N_2424,In_1081,In_1149);
and U2425 (N_2425,In_1000,In_861);
and U2426 (N_2426,In_1124,In_99);
nand U2427 (N_2427,In_1312,In_633);
nor U2428 (N_2428,In_331,In_588);
and U2429 (N_2429,In_1177,In_1388);
nor U2430 (N_2430,In_741,In_1163);
nor U2431 (N_2431,In_1318,In_1160);
nor U2432 (N_2432,In_1070,In_443);
nand U2433 (N_2433,In_1083,In_717);
nand U2434 (N_2434,In_566,In_1065);
and U2435 (N_2435,In_1168,In_848);
and U2436 (N_2436,In_1197,In_1105);
nand U2437 (N_2437,In_669,In_1281);
nand U2438 (N_2438,In_652,In_53);
nor U2439 (N_2439,In_382,In_332);
nor U2440 (N_2440,In_1322,In_1054);
and U2441 (N_2441,In_1196,In_801);
nand U2442 (N_2442,In_1215,In_856);
nand U2443 (N_2443,In_1459,In_1290);
and U2444 (N_2444,In_764,In_1182);
or U2445 (N_2445,In_518,In_1405);
and U2446 (N_2446,In_843,In_676);
nor U2447 (N_2447,In_256,In_1239);
nand U2448 (N_2448,In_279,In_1479);
nor U2449 (N_2449,In_767,In_1052);
and U2450 (N_2450,In_1337,In_1394);
nand U2451 (N_2451,In_1435,In_594);
or U2452 (N_2452,In_345,In_693);
nand U2453 (N_2453,In_1061,In_692);
nand U2454 (N_2454,In_1237,In_1362);
and U2455 (N_2455,In_772,In_868);
and U2456 (N_2456,In_6,In_717);
nor U2457 (N_2457,In_1207,In_455);
nor U2458 (N_2458,In_389,In_270);
nand U2459 (N_2459,In_590,In_1160);
xnor U2460 (N_2460,In_18,In_150);
and U2461 (N_2461,In_871,In_832);
nor U2462 (N_2462,In_1353,In_967);
and U2463 (N_2463,In_1315,In_1343);
nand U2464 (N_2464,In_804,In_947);
and U2465 (N_2465,In_204,In_1043);
and U2466 (N_2466,In_896,In_563);
xnor U2467 (N_2467,In_802,In_1304);
nor U2468 (N_2468,In_599,In_893);
and U2469 (N_2469,In_207,In_1293);
nand U2470 (N_2470,In_1274,In_76);
or U2471 (N_2471,In_149,In_596);
or U2472 (N_2472,In_1196,In_731);
and U2473 (N_2473,In_982,In_285);
or U2474 (N_2474,In_1425,In_1024);
or U2475 (N_2475,In_677,In_176);
nand U2476 (N_2476,In_1308,In_159);
nand U2477 (N_2477,In_1074,In_1159);
or U2478 (N_2478,In_737,In_745);
and U2479 (N_2479,In_1100,In_104);
nor U2480 (N_2480,In_1109,In_329);
nor U2481 (N_2481,In_197,In_323);
and U2482 (N_2482,In_1468,In_219);
or U2483 (N_2483,In_1394,In_1078);
nor U2484 (N_2484,In_766,In_633);
and U2485 (N_2485,In_581,In_1003);
nand U2486 (N_2486,In_1274,In_670);
nor U2487 (N_2487,In_844,In_20);
or U2488 (N_2488,In_1360,In_1290);
nor U2489 (N_2489,In_1322,In_861);
or U2490 (N_2490,In_179,In_631);
nand U2491 (N_2491,In_65,In_1110);
nor U2492 (N_2492,In_405,In_61);
nand U2493 (N_2493,In_1055,In_657);
or U2494 (N_2494,In_1097,In_1275);
and U2495 (N_2495,In_1054,In_979);
and U2496 (N_2496,In_1442,In_1414);
nor U2497 (N_2497,In_320,In_26);
nor U2498 (N_2498,In_1335,In_1258);
nor U2499 (N_2499,In_1198,In_166);
or U2500 (N_2500,In_1235,In_1039);
nand U2501 (N_2501,In_834,In_669);
and U2502 (N_2502,In_782,In_1237);
nor U2503 (N_2503,In_1393,In_1387);
or U2504 (N_2504,In_795,In_888);
nand U2505 (N_2505,In_606,In_300);
or U2506 (N_2506,In_1365,In_242);
or U2507 (N_2507,In_1137,In_1108);
or U2508 (N_2508,In_545,In_279);
and U2509 (N_2509,In_876,In_458);
nor U2510 (N_2510,In_35,In_706);
nand U2511 (N_2511,In_185,In_1454);
nand U2512 (N_2512,In_828,In_1499);
nand U2513 (N_2513,In_853,In_328);
nor U2514 (N_2514,In_1444,In_32);
or U2515 (N_2515,In_379,In_465);
and U2516 (N_2516,In_88,In_1360);
or U2517 (N_2517,In_1320,In_744);
nand U2518 (N_2518,In_1026,In_72);
or U2519 (N_2519,In_1353,In_201);
nor U2520 (N_2520,In_333,In_814);
nand U2521 (N_2521,In_409,In_488);
and U2522 (N_2522,In_1284,In_80);
nor U2523 (N_2523,In_657,In_846);
nand U2524 (N_2524,In_601,In_768);
and U2525 (N_2525,In_1352,In_256);
nor U2526 (N_2526,In_163,In_1419);
nor U2527 (N_2527,In_1130,In_423);
and U2528 (N_2528,In_1260,In_726);
and U2529 (N_2529,In_1417,In_95);
or U2530 (N_2530,In_926,In_371);
and U2531 (N_2531,In_239,In_248);
and U2532 (N_2532,In_456,In_206);
nor U2533 (N_2533,In_1196,In_1428);
and U2534 (N_2534,In_1354,In_383);
or U2535 (N_2535,In_1053,In_1080);
or U2536 (N_2536,In_336,In_366);
and U2537 (N_2537,In_152,In_501);
nand U2538 (N_2538,In_286,In_189);
or U2539 (N_2539,In_595,In_179);
or U2540 (N_2540,In_819,In_716);
and U2541 (N_2541,In_767,In_577);
or U2542 (N_2542,In_1399,In_1427);
or U2543 (N_2543,In_759,In_1258);
and U2544 (N_2544,In_1488,In_599);
and U2545 (N_2545,In_1492,In_1250);
or U2546 (N_2546,In_265,In_588);
nor U2547 (N_2547,In_701,In_46);
nand U2548 (N_2548,In_1346,In_431);
or U2549 (N_2549,In_679,In_124);
and U2550 (N_2550,In_343,In_334);
or U2551 (N_2551,In_204,In_1331);
or U2552 (N_2552,In_1274,In_724);
nand U2553 (N_2553,In_157,In_213);
nand U2554 (N_2554,In_995,In_1099);
and U2555 (N_2555,In_423,In_736);
and U2556 (N_2556,In_1334,In_167);
nor U2557 (N_2557,In_92,In_27);
and U2558 (N_2558,In_163,In_1483);
or U2559 (N_2559,In_1221,In_606);
or U2560 (N_2560,In_155,In_142);
nor U2561 (N_2561,In_308,In_1157);
nand U2562 (N_2562,In_255,In_781);
and U2563 (N_2563,In_597,In_1480);
nor U2564 (N_2564,In_912,In_826);
or U2565 (N_2565,In_535,In_1456);
and U2566 (N_2566,In_524,In_1030);
or U2567 (N_2567,In_320,In_515);
and U2568 (N_2568,In_1020,In_97);
nor U2569 (N_2569,In_100,In_1042);
nor U2570 (N_2570,In_669,In_758);
nor U2571 (N_2571,In_173,In_1424);
nand U2572 (N_2572,In_868,In_930);
nand U2573 (N_2573,In_1441,In_848);
or U2574 (N_2574,In_250,In_1479);
and U2575 (N_2575,In_1420,In_971);
nand U2576 (N_2576,In_264,In_939);
nand U2577 (N_2577,In_1443,In_637);
nor U2578 (N_2578,In_574,In_800);
and U2579 (N_2579,In_283,In_51);
or U2580 (N_2580,In_1172,In_994);
and U2581 (N_2581,In_1449,In_44);
or U2582 (N_2582,In_161,In_434);
nor U2583 (N_2583,In_1125,In_253);
nand U2584 (N_2584,In_186,In_612);
and U2585 (N_2585,In_869,In_687);
or U2586 (N_2586,In_923,In_689);
nor U2587 (N_2587,In_1046,In_821);
or U2588 (N_2588,In_206,In_29);
and U2589 (N_2589,In_263,In_69);
nand U2590 (N_2590,In_20,In_318);
and U2591 (N_2591,In_1471,In_1418);
nor U2592 (N_2592,In_446,In_833);
or U2593 (N_2593,In_1102,In_82);
nand U2594 (N_2594,In_43,In_479);
or U2595 (N_2595,In_967,In_1130);
and U2596 (N_2596,In_1393,In_43);
nand U2597 (N_2597,In_240,In_650);
nor U2598 (N_2598,In_14,In_807);
and U2599 (N_2599,In_676,In_1145);
nor U2600 (N_2600,In_1200,In_561);
nor U2601 (N_2601,In_717,In_1066);
nor U2602 (N_2602,In_136,In_986);
nand U2603 (N_2603,In_452,In_77);
nand U2604 (N_2604,In_341,In_793);
nor U2605 (N_2605,In_18,In_701);
nor U2606 (N_2606,In_280,In_683);
and U2607 (N_2607,In_638,In_384);
and U2608 (N_2608,In_650,In_333);
nor U2609 (N_2609,In_862,In_884);
or U2610 (N_2610,In_1407,In_439);
or U2611 (N_2611,In_853,In_1448);
and U2612 (N_2612,In_1458,In_316);
and U2613 (N_2613,In_357,In_761);
nand U2614 (N_2614,In_855,In_1038);
and U2615 (N_2615,In_1064,In_1019);
or U2616 (N_2616,In_381,In_911);
and U2617 (N_2617,In_283,In_562);
or U2618 (N_2618,In_445,In_1192);
and U2619 (N_2619,In_75,In_940);
and U2620 (N_2620,In_305,In_299);
or U2621 (N_2621,In_241,In_494);
nor U2622 (N_2622,In_394,In_169);
and U2623 (N_2623,In_1176,In_778);
and U2624 (N_2624,In_1022,In_1448);
and U2625 (N_2625,In_857,In_1314);
nor U2626 (N_2626,In_626,In_923);
nor U2627 (N_2627,In_461,In_1218);
or U2628 (N_2628,In_593,In_355);
or U2629 (N_2629,In_500,In_39);
nor U2630 (N_2630,In_913,In_288);
nor U2631 (N_2631,In_1136,In_362);
nor U2632 (N_2632,In_97,In_1101);
and U2633 (N_2633,In_155,In_1318);
xor U2634 (N_2634,In_961,In_891);
xor U2635 (N_2635,In_409,In_1191);
nor U2636 (N_2636,In_847,In_655);
nor U2637 (N_2637,In_990,In_761);
nand U2638 (N_2638,In_1017,In_1055);
and U2639 (N_2639,In_1291,In_426);
or U2640 (N_2640,In_1128,In_366);
or U2641 (N_2641,In_928,In_1440);
and U2642 (N_2642,In_448,In_1143);
nor U2643 (N_2643,In_881,In_1263);
nor U2644 (N_2644,In_1447,In_1375);
and U2645 (N_2645,In_287,In_1438);
nor U2646 (N_2646,In_1355,In_1064);
and U2647 (N_2647,In_525,In_1027);
or U2648 (N_2648,In_1357,In_593);
and U2649 (N_2649,In_825,In_1156);
nand U2650 (N_2650,In_1192,In_1072);
nand U2651 (N_2651,In_111,In_677);
and U2652 (N_2652,In_1291,In_281);
nor U2653 (N_2653,In_388,In_409);
or U2654 (N_2654,In_1456,In_1199);
or U2655 (N_2655,In_855,In_565);
and U2656 (N_2656,In_415,In_664);
nor U2657 (N_2657,In_221,In_744);
nor U2658 (N_2658,In_429,In_638);
or U2659 (N_2659,In_1469,In_1454);
or U2660 (N_2660,In_111,In_594);
and U2661 (N_2661,In_1333,In_470);
xor U2662 (N_2662,In_138,In_1064);
nor U2663 (N_2663,In_31,In_898);
nor U2664 (N_2664,In_40,In_1464);
nor U2665 (N_2665,In_644,In_1018);
nand U2666 (N_2666,In_916,In_718);
or U2667 (N_2667,In_544,In_1044);
and U2668 (N_2668,In_17,In_985);
nand U2669 (N_2669,In_981,In_634);
nor U2670 (N_2670,In_1188,In_1395);
and U2671 (N_2671,In_1118,In_124);
nor U2672 (N_2672,In_1170,In_306);
nand U2673 (N_2673,In_1421,In_359);
or U2674 (N_2674,In_1088,In_396);
nand U2675 (N_2675,In_147,In_940);
and U2676 (N_2676,In_1130,In_1028);
or U2677 (N_2677,In_856,In_240);
or U2678 (N_2678,In_266,In_280);
nor U2679 (N_2679,In_737,In_443);
nand U2680 (N_2680,In_453,In_411);
nor U2681 (N_2681,In_38,In_881);
nand U2682 (N_2682,In_793,In_1417);
and U2683 (N_2683,In_900,In_469);
nand U2684 (N_2684,In_135,In_322);
nor U2685 (N_2685,In_257,In_1349);
nand U2686 (N_2686,In_302,In_713);
nand U2687 (N_2687,In_947,In_758);
and U2688 (N_2688,In_1195,In_342);
and U2689 (N_2689,In_316,In_972);
nor U2690 (N_2690,In_37,In_527);
or U2691 (N_2691,In_401,In_1181);
xnor U2692 (N_2692,In_975,In_1025);
nor U2693 (N_2693,In_821,In_332);
and U2694 (N_2694,In_554,In_1252);
nand U2695 (N_2695,In_1230,In_566);
and U2696 (N_2696,In_1249,In_408);
xnor U2697 (N_2697,In_1346,In_242);
nor U2698 (N_2698,In_889,In_130);
or U2699 (N_2699,In_835,In_108);
nand U2700 (N_2700,In_50,In_303);
and U2701 (N_2701,In_872,In_838);
nand U2702 (N_2702,In_1497,In_930);
nor U2703 (N_2703,In_582,In_1177);
or U2704 (N_2704,In_106,In_1155);
nor U2705 (N_2705,In_1402,In_240);
and U2706 (N_2706,In_894,In_1101);
and U2707 (N_2707,In_961,In_16);
and U2708 (N_2708,In_41,In_146);
nor U2709 (N_2709,In_561,In_994);
or U2710 (N_2710,In_59,In_752);
and U2711 (N_2711,In_875,In_540);
nand U2712 (N_2712,In_962,In_226);
nor U2713 (N_2713,In_437,In_20);
and U2714 (N_2714,In_133,In_1235);
xnor U2715 (N_2715,In_112,In_929);
and U2716 (N_2716,In_1241,In_93);
or U2717 (N_2717,In_170,In_273);
or U2718 (N_2718,In_1012,In_844);
and U2719 (N_2719,In_1041,In_510);
or U2720 (N_2720,In_420,In_721);
nor U2721 (N_2721,In_75,In_870);
or U2722 (N_2722,In_91,In_614);
and U2723 (N_2723,In_792,In_1395);
nor U2724 (N_2724,In_160,In_78);
or U2725 (N_2725,In_748,In_674);
nor U2726 (N_2726,In_477,In_925);
nor U2727 (N_2727,In_510,In_419);
nand U2728 (N_2728,In_1398,In_700);
nor U2729 (N_2729,In_643,In_943);
nand U2730 (N_2730,In_834,In_731);
nor U2731 (N_2731,In_117,In_501);
or U2732 (N_2732,In_1472,In_385);
or U2733 (N_2733,In_1314,In_626);
or U2734 (N_2734,In_747,In_502);
and U2735 (N_2735,In_730,In_1186);
or U2736 (N_2736,In_627,In_1391);
nand U2737 (N_2737,In_624,In_530);
nor U2738 (N_2738,In_813,In_309);
nand U2739 (N_2739,In_702,In_1242);
or U2740 (N_2740,In_1189,In_23);
and U2741 (N_2741,In_451,In_311);
and U2742 (N_2742,In_1315,In_231);
xor U2743 (N_2743,In_204,In_313);
or U2744 (N_2744,In_1370,In_939);
nand U2745 (N_2745,In_110,In_911);
nand U2746 (N_2746,In_812,In_885);
nand U2747 (N_2747,In_433,In_1497);
nor U2748 (N_2748,In_1050,In_982);
nand U2749 (N_2749,In_1350,In_1414);
and U2750 (N_2750,In_47,In_799);
nor U2751 (N_2751,In_587,In_889);
and U2752 (N_2752,In_2,In_574);
nor U2753 (N_2753,In_477,In_1322);
nand U2754 (N_2754,In_1193,In_467);
and U2755 (N_2755,In_1233,In_49);
nor U2756 (N_2756,In_700,In_808);
nor U2757 (N_2757,In_674,In_220);
nand U2758 (N_2758,In_658,In_1390);
and U2759 (N_2759,In_390,In_630);
nand U2760 (N_2760,In_225,In_665);
nor U2761 (N_2761,In_599,In_12);
and U2762 (N_2762,In_386,In_656);
and U2763 (N_2763,In_1047,In_1238);
and U2764 (N_2764,In_666,In_79);
or U2765 (N_2765,In_694,In_279);
nand U2766 (N_2766,In_919,In_374);
or U2767 (N_2767,In_1066,In_728);
or U2768 (N_2768,In_50,In_44);
nand U2769 (N_2769,In_204,In_1437);
and U2770 (N_2770,In_398,In_1347);
or U2771 (N_2771,In_217,In_590);
and U2772 (N_2772,In_1465,In_58);
or U2773 (N_2773,In_1061,In_920);
or U2774 (N_2774,In_1392,In_528);
nand U2775 (N_2775,In_1116,In_58);
or U2776 (N_2776,In_398,In_291);
nand U2777 (N_2777,In_120,In_1396);
and U2778 (N_2778,In_127,In_286);
nor U2779 (N_2779,In_180,In_1130);
nor U2780 (N_2780,In_1394,In_599);
and U2781 (N_2781,In_786,In_1027);
and U2782 (N_2782,In_533,In_1309);
and U2783 (N_2783,In_1015,In_71);
nor U2784 (N_2784,In_738,In_56);
nand U2785 (N_2785,In_793,In_1420);
nor U2786 (N_2786,In_1245,In_1079);
and U2787 (N_2787,In_1020,In_503);
or U2788 (N_2788,In_1439,In_1125);
and U2789 (N_2789,In_558,In_77);
or U2790 (N_2790,In_1310,In_1009);
or U2791 (N_2791,In_940,In_915);
and U2792 (N_2792,In_1490,In_819);
nand U2793 (N_2793,In_950,In_1169);
and U2794 (N_2794,In_831,In_1241);
and U2795 (N_2795,In_407,In_415);
nor U2796 (N_2796,In_1213,In_560);
nand U2797 (N_2797,In_801,In_670);
or U2798 (N_2798,In_527,In_1220);
nand U2799 (N_2799,In_447,In_525);
nand U2800 (N_2800,In_470,In_1038);
nor U2801 (N_2801,In_584,In_1339);
and U2802 (N_2802,In_725,In_325);
nand U2803 (N_2803,In_869,In_838);
and U2804 (N_2804,In_1269,In_1158);
nand U2805 (N_2805,In_851,In_670);
nand U2806 (N_2806,In_282,In_456);
and U2807 (N_2807,In_823,In_1393);
and U2808 (N_2808,In_988,In_181);
and U2809 (N_2809,In_370,In_968);
nand U2810 (N_2810,In_1327,In_1147);
nor U2811 (N_2811,In_1228,In_636);
or U2812 (N_2812,In_437,In_400);
nor U2813 (N_2813,In_28,In_495);
or U2814 (N_2814,In_290,In_785);
and U2815 (N_2815,In_1152,In_497);
nand U2816 (N_2816,In_911,In_421);
and U2817 (N_2817,In_143,In_1400);
and U2818 (N_2818,In_330,In_939);
nor U2819 (N_2819,In_1272,In_679);
or U2820 (N_2820,In_1281,In_494);
or U2821 (N_2821,In_705,In_950);
and U2822 (N_2822,In_411,In_256);
or U2823 (N_2823,In_312,In_674);
nand U2824 (N_2824,In_261,In_1255);
nor U2825 (N_2825,In_183,In_824);
and U2826 (N_2826,In_323,In_140);
nand U2827 (N_2827,In_417,In_493);
nand U2828 (N_2828,In_379,In_865);
nand U2829 (N_2829,In_925,In_450);
nor U2830 (N_2830,In_409,In_1053);
and U2831 (N_2831,In_907,In_1127);
nand U2832 (N_2832,In_1350,In_901);
or U2833 (N_2833,In_1334,In_765);
or U2834 (N_2834,In_1365,In_247);
or U2835 (N_2835,In_1449,In_1175);
and U2836 (N_2836,In_163,In_1359);
nand U2837 (N_2837,In_1265,In_626);
or U2838 (N_2838,In_1057,In_1164);
nand U2839 (N_2839,In_551,In_1413);
and U2840 (N_2840,In_1484,In_678);
nor U2841 (N_2841,In_1446,In_1242);
or U2842 (N_2842,In_594,In_574);
nand U2843 (N_2843,In_1102,In_219);
and U2844 (N_2844,In_535,In_524);
or U2845 (N_2845,In_1395,In_8);
nor U2846 (N_2846,In_166,In_371);
and U2847 (N_2847,In_506,In_753);
nor U2848 (N_2848,In_1170,In_301);
nor U2849 (N_2849,In_448,In_279);
nor U2850 (N_2850,In_648,In_920);
or U2851 (N_2851,In_884,In_384);
nor U2852 (N_2852,In_931,In_603);
nor U2853 (N_2853,In_1431,In_532);
nand U2854 (N_2854,In_828,In_918);
or U2855 (N_2855,In_912,In_56);
nor U2856 (N_2856,In_505,In_219);
nand U2857 (N_2857,In_760,In_610);
or U2858 (N_2858,In_1137,In_862);
or U2859 (N_2859,In_577,In_497);
and U2860 (N_2860,In_562,In_631);
nand U2861 (N_2861,In_559,In_98);
nor U2862 (N_2862,In_1444,In_1309);
nand U2863 (N_2863,In_1180,In_414);
nor U2864 (N_2864,In_612,In_301);
or U2865 (N_2865,In_483,In_1098);
nor U2866 (N_2866,In_1274,In_846);
or U2867 (N_2867,In_378,In_1293);
nor U2868 (N_2868,In_720,In_673);
and U2869 (N_2869,In_1096,In_1210);
or U2870 (N_2870,In_795,In_1278);
or U2871 (N_2871,In_677,In_1343);
nor U2872 (N_2872,In_255,In_679);
and U2873 (N_2873,In_748,In_47);
and U2874 (N_2874,In_1043,In_1362);
nand U2875 (N_2875,In_11,In_1158);
or U2876 (N_2876,In_1318,In_1174);
nor U2877 (N_2877,In_933,In_151);
nand U2878 (N_2878,In_716,In_623);
or U2879 (N_2879,In_889,In_645);
nand U2880 (N_2880,In_466,In_100);
nand U2881 (N_2881,In_381,In_186);
or U2882 (N_2882,In_1496,In_569);
nand U2883 (N_2883,In_1414,In_1384);
and U2884 (N_2884,In_1423,In_737);
and U2885 (N_2885,In_1187,In_207);
nand U2886 (N_2886,In_389,In_36);
nor U2887 (N_2887,In_1460,In_608);
nor U2888 (N_2888,In_267,In_570);
nand U2889 (N_2889,In_666,In_1281);
and U2890 (N_2890,In_14,In_98);
nor U2891 (N_2891,In_553,In_608);
and U2892 (N_2892,In_668,In_806);
nand U2893 (N_2893,In_474,In_1463);
or U2894 (N_2894,In_447,In_1052);
and U2895 (N_2895,In_833,In_1308);
nand U2896 (N_2896,In_663,In_1054);
and U2897 (N_2897,In_76,In_584);
nand U2898 (N_2898,In_459,In_587);
nor U2899 (N_2899,In_265,In_1418);
nor U2900 (N_2900,In_1213,In_254);
and U2901 (N_2901,In_699,In_1301);
and U2902 (N_2902,In_1200,In_999);
nor U2903 (N_2903,In_1265,In_1285);
nor U2904 (N_2904,In_1113,In_393);
and U2905 (N_2905,In_1030,In_503);
nand U2906 (N_2906,In_265,In_474);
nand U2907 (N_2907,In_1231,In_63);
and U2908 (N_2908,In_968,In_619);
nand U2909 (N_2909,In_204,In_1275);
nand U2910 (N_2910,In_1327,In_334);
and U2911 (N_2911,In_533,In_1152);
or U2912 (N_2912,In_296,In_748);
nor U2913 (N_2913,In_760,In_175);
nor U2914 (N_2914,In_956,In_1086);
or U2915 (N_2915,In_182,In_1265);
nand U2916 (N_2916,In_1348,In_1472);
or U2917 (N_2917,In_102,In_107);
nand U2918 (N_2918,In_552,In_179);
nor U2919 (N_2919,In_1049,In_596);
or U2920 (N_2920,In_1490,In_1173);
or U2921 (N_2921,In_944,In_968);
nand U2922 (N_2922,In_276,In_465);
or U2923 (N_2923,In_363,In_1334);
and U2924 (N_2924,In_105,In_563);
or U2925 (N_2925,In_340,In_1475);
and U2926 (N_2926,In_414,In_336);
nor U2927 (N_2927,In_1,In_396);
nor U2928 (N_2928,In_1122,In_737);
nor U2929 (N_2929,In_362,In_273);
nand U2930 (N_2930,In_406,In_273);
nor U2931 (N_2931,In_966,In_1281);
and U2932 (N_2932,In_17,In_1442);
nor U2933 (N_2933,In_688,In_320);
nand U2934 (N_2934,In_488,In_1451);
nand U2935 (N_2935,In_986,In_1180);
nor U2936 (N_2936,In_932,In_504);
nor U2937 (N_2937,In_20,In_381);
or U2938 (N_2938,In_995,In_510);
nor U2939 (N_2939,In_756,In_328);
nor U2940 (N_2940,In_551,In_674);
nand U2941 (N_2941,In_278,In_1141);
and U2942 (N_2942,In_1345,In_1300);
nor U2943 (N_2943,In_823,In_876);
and U2944 (N_2944,In_1199,In_414);
and U2945 (N_2945,In_865,In_1271);
nor U2946 (N_2946,In_844,In_647);
nor U2947 (N_2947,In_1497,In_215);
nor U2948 (N_2948,In_1225,In_1490);
nand U2949 (N_2949,In_952,In_412);
nor U2950 (N_2950,In_834,In_158);
or U2951 (N_2951,In_281,In_874);
nor U2952 (N_2952,In_582,In_842);
nand U2953 (N_2953,In_327,In_1252);
nor U2954 (N_2954,In_316,In_899);
and U2955 (N_2955,In_1436,In_647);
nor U2956 (N_2956,In_181,In_1354);
or U2957 (N_2957,In_277,In_207);
nor U2958 (N_2958,In_96,In_974);
and U2959 (N_2959,In_1483,In_1104);
and U2960 (N_2960,In_180,In_1219);
or U2961 (N_2961,In_653,In_795);
nor U2962 (N_2962,In_1082,In_964);
or U2963 (N_2963,In_269,In_1482);
or U2964 (N_2964,In_348,In_1347);
nand U2965 (N_2965,In_871,In_386);
and U2966 (N_2966,In_1208,In_371);
or U2967 (N_2967,In_535,In_514);
and U2968 (N_2968,In_672,In_1443);
or U2969 (N_2969,In_1074,In_656);
or U2970 (N_2970,In_705,In_1430);
nor U2971 (N_2971,In_462,In_1358);
or U2972 (N_2972,In_1253,In_405);
or U2973 (N_2973,In_1140,In_1354);
nor U2974 (N_2974,In_591,In_958);
nand U2975 (N_2975,In_1330,In_1006);
and U2976 (N_2976,In_1279,In_738);
and U2977 (N_2977,In_1248,In_1115);
nand U2978 (N_2978,In_1411,In_1282);
or U2979 (N_2979,In_1294,In_838);
and U2980 (N_2980,In_1199,In_54);
or U2981 (N_2981,In_165,In_1034);
nand U2982 (N_2982,In_170,In_562);
and U2983 (N_2983,In_521,In_12);
or U2984 (N_2984,In_181,In_159);
nor U2985 (N_2985,In_1205,In_670);
or U2986 (N_2986,In_533,In_1383);
or U2987 (N_2987,In_1448,In_1258);
and U2988 (N_2988,In_114,In_557);
nor U2989 (N_2989,In_740,In_809);
or U2990 (N_2990,In_934,In_574);
xor U2991 (N_2991,In_1267,In_1167);
or U2992 (N_2992,In_52,In_254);
and U2993 (N_2993,In_1487,In_1195);
nand U2994 (N_2994,In_1053,In_800);
and U2995 (N_2995,In_846,In_183);
or U2996 (N_2996,In_883,In_849);
or U2997 (N_2997,In_336,In_425);
nor U2998 (N_2998,In_1422,In_408);
nor U2999 (N_2999,In_874,In_459);
and U3000 (N_3000,N_1949,N_31);
or U3001 (N_3001,N_902,N_1860);
or U3002 (N_3002,N_2225,N_1716);
and U3003 (N_3003,N_2267,N_2117);
or U3004 (N_3004,N_378,N_2410);
and U3005 (N_3005,N_1131,N_2269);
nor U3006 (N_3006,N_1407,N_543);
or U3007 (N_3007,N_2286,N_2726);
and U3008 (N_3008,N_1675,N_1891);
or U3009 (N_3009,N_1300,N_2378);
and U3010 (N_3010,N_395,N_1390);
nor U3011 (N_3011,N_2630,N_1046);
and U3012 (N_3012,N_821,N_908);
and U3013 (N_3013,N_1906,N_2150);
or U3014 (N_3014,N_1665,N_504);
nor U3015 (N_3015,N_878,N_1862);
nand U3016 (N_3016,N_398,N_219);
or U3017 (N_3017,N_611,N_1491);
nor U3018 (N_3018,N_1613,N_1393);
nor U3019 (N_3019,N_1766,N_1041);
and U3020 (N_3020,N_2454,N_781);
or U3021 (N_3021,N_2189,N_1098);
and U3022 (N_3022,N_2990,N_1115);
nand U3023 (N_3023,N_1615,N_602);
nor U3024 (N_3024,N_1264,N_2355);
nor U3025 (N_3025,N_1371,N_337);
and U3026 (N_3026,N_1343,N_664);
or U3027 (N_3027,N_468,N_605);
nor U3028 (N_3028,N_2908,N_2473);
or U3029 (N_3029,N_894,N_1494);
nor U3030 (N_3030,N_172,N_1480);
nand U3031 (N_3031,N_2377,N_32);
nand U3032 (N_3032,N_2558,N_2541);
or U3033 (N_3033,N_356,N_1247);
nor U3034 (N_3034,N_1322,N_2614);
and U3035 (N_3035,N_60,N_2825);
or U3036 (N_3036,N_2211,N_343);
and U3037 (N_3037,N_2492,N_2027);
and U3038 (N_3038,N_2668,N_485);
or U3039 (N_3039,N_1798,N_2539);
and U3040 (N_3040,N_1336,N_2300);
nand U3041 (N_3041,N_2640,N_647);
nor U3042 (N_3042,N_364,N_1749);
nor U3043 (N_3043,N_251,N_1717);
or U3044 (N_3044,N_2065,N_693);
or U3045 (N_3045,N_2464,N_1738);
or U3046 (N_3046,N_2689,N_1169);
or U3047 (N_3047,N_2238,N_1516);
nor U3048 (N_3048,N_1005,N_606);
and U3049 (N_3049,N_1700,N_2548);
and U3050 (N_3050,N_133,N_899);
and U3051 (N_3051,N_1340,N_2822);
and U3052 (N_3052,N_2025,N_216);
and U3053 (N_3053,N_1268,N_1959);
and U3054 (N_3054,N_1114,N_199);
and U3055 (N_3055,N_2873,N_1844);
and U3056 (N_3056,N_1653,N_2383);
nand U3057 (N_3057,N_182,N_1708);
nand U3058 (N_3058,N_1043,N_2111);
nor U3059 (N_3059,N_1463,N_951);
nor U3060 (N_3060,N_2859,N_2216);
and U3061 (N_3061,N_2317,N_234);
nor U3062 (N_3062,N_1807,N_249);
and U3063 (N_3063,N_1448,N_2368);
and U3064 (N_3064,N_2394,N_1026);
or U3065 (N_3065,N_660,N_152);
or U3066 (N_3066,N_1078,N_1012);
or U3067 (N_3067,N_1585,N_1377);
nor U3068 (N_3068,N_2890,N_2250);
and U3069 (N_3069,N_2666,N_203);
nor U3070 (N_3070,N_840,N_1584);
nor U3071 (N_3071,N_1559,N_2574);
nor U3072 (N_3072,N_1238,N_2680);
or U3073 (N_3073,N_547,N_2973);
or U3074 (N_3074,N_2006,N_1861);
nand U3075 (N_3075,N_1299,N_1755);
nand U3076 (N_3076,N_1873,N_589);
nor U3077 (N_3077,N_1878,N_1187);
xor U3078 (N_3078,N_515,N_920);
nor U3079 (N_3079,N_1089,N_1375);
or U3080 (N_3080,N_1313,N_2572);
and U3081 (N_3081,N_437,N_1261);
or U3082 (N_3082,N_2308,N_1353);
nor U3083 (N_3083,N_1705,N_1519);
and U3084 (N_3084,N_1142,N_639);
nand U3085 (N_3085,N_2984,N_2443);
nor U3086 (N_3086,N_1792,N_2352);
or U3087 (N_3087,N_2917,N_1603);
nand U3088 (N_3088,N_2370,N_2149);
nor U3089 (N_3089,N_2869,N_2838);
nor U3090 (N_3090,N_1571,N_1869);
and U3091 (N_3091,N_52,N_1751);
and U3092 (N_3092,N_2024,N_910);
or U3093 (N_3093,N_1863,N_1294);
or U3094 (N_3094,N_1944,N_2381);
nor U3095 (N_3095,N_2886,N_2369);
or U3096 (N_3096,N_671,N_381);
nor U3097 (N_3097,N_2993,N_2661);
nand U3098 (N_3098,N_2324,N_788);
or U3099 (N_3099,N_2561,N_191);
nand U3100 (N_3100,N_301,N_2339);
or U3101 (N_3101,N_108,N_520);
and U3102 (N_3102,N_223,N_2232);
nand U3103 (N_3103,N_2647,N_706);
nor U3104 (N_3104,N_2123,N_1984);
and U3105 (N_3105,N_1193,N_2891);
and U3106 (N_3106,N_526,N_2379);
and U3107 (N_3107,N_407,N_1765);
and U3108 (N_3108,N_101,N_569);
or U3109 (N_3109,N_1919,N_1179);
or U3110 (N_3110,N_1720,N_918);
nor U3111 (N_3111,N_2280,N_2625);
nand U3112 (N_3112,N_134,N_1172);
nor U3113 (N_3113,N_1376,N_1610);
and U3114 (N_3114,N_1667,N_1059);
nand U3115 (N_3115,N_846,N_698);
nor U3116 (N_3116,N_1021,N_1488);
nand U3117 (N_3117,N_287,N_651);
and U3118 (N_3118,N_474,N_1339);
and U3119 (N_3119,N_1835,N_2129);
or U3120 (N_3120,N_1245,N_74);
xor U3121 (N_3121,N_1432,N_1152);
nand U3122 (N_3122,N_1857,N_766);
or U3123 (N_3123,N_75,N_2184);
or U3124 (N_3124,N_2900,N_1562);
or U3125 (N_3125,N_2427,N_1147);
nor U3126 (N_3126,N_2944,N_132);
nor U3127 (N_3127,N_2444,N_2739);
and U3128 (N_3128,N_1301,N_1058);
nand U3129 (N_3129,N_2309,N_2063);
nor U3130 (N_3130,N_893,N_231);
and U3131 (N_3131,N_2981,N_741);
nor U3132 (N_3132,N_392,N_36);
and U3133 (N_3133,N_1129,N_2023);
nand U3134 (N_3134,N_571,N_2802);
xnor U3135 (N_3135,N_747,N_2135);
nand U3136 (N_3136,N_2830,N_2619);
nand U3137 (N_3137,N_2770,N_1706);
nor U3138 (N_3138,N_169,N_1797);
nand U3139 (N_3139,N_1223,N_1543);
nand U3140 (N_3140,N_154,N_2179);
or U3141 (N_3141,N_2380,N_1606);
and U3142 (N_3142,N_2503,N_1827);
nand U3143 (N_3143,N_1537,N_367);
and U3144 (N_3144,N_968,N_1345);
nand U3145 (N_3145,N_1305,N_2477);
or U3146 (N_3146,N_1400,N_986);
or U3147 (N_3147,N_1618,N_1221);
nand U3148 (N_3148,N_88,N_1699);
and U3149 (N_3149,N_1501,N_1985);
or U3150 (N_3150,N_947,N_66);
or U3151 (N_3151,N_2496,N_2060);
nor U3152 (N_3152,N_278,N_1594);
and U3153 (N_3153,N_604,N_1824);
nor U3154 (N_3154,N_214,N_2089);
nor U3155 (N_3155,N_2602,N_1538);
nand U3156 (N_3156,N_1572,N_2601);
nor U3157 (N_3157,N_1381,N_2453);
nand U3158 (N_3158,N_768,N_2092);
nand U3159 (N_3159,N_2698,N_1282);
or U3160 (N_3160,N_848,N_945);
nand U3161 (N_3161,N_1033,N_2846);
nand U3162 (N_3162,N_646,N_361);
nor U3163 (N_3163,N_552,N_276);
nand U3164 (N_3164,N_2745,N_1638);
nand U3165 (N_3165,N_1512,N_389);
or U3166 (N_3166,N_1583,N_1287);
or U3167 (N_3167,N_2794,N_2479);
nor U3168 (N_3168,N_833,N_815);
nor U3169 (N_3169,N_1391,N_141);
nor U3170 (N_3170,N_1595,N_415);
and U3171 (N_3171,N_2605,N_2667);
nand U3172 (N_3172,N_2285,N_2079);
nand U3173 (N_3173,N_2249,N_26);
nand U3174 (N_3174,N_673,N_1405);
and U3175 (N_3175,N_1894,N_898);
and U3176 (N_3176,N_1304,N_142);
nor U3177 (N_3177,N_1982,N_2939);
nand U3178 (N_3178,N_2449,N_2411);
and U3179 (N_3179,N_1229,N_517);
nand U3180 (N_3180,N_652,N_872);
or U3181 (N_3181,N_827,N_1761);
nor U3182 (N_3182,N_1234,N_1580);
or U3183 (N_3183,N_2969,N_923);
nor U3184 (N_3184,N_518,N_1714);
nand U3185 (N_3185,N_2279,N_644);
or U3186 (N_3186,N_1219,N_2559);
nor U3187 (N_3187,N_2043,N_252);
and U3188 (N_3188,N_1577,N_603);
and U3189 (N_3189,N_1703,N_2550);
or U3190 (N_3190,N_432,N_718);
nor U3191 (N_3191,N_2108,N_1009);
nand U3192 (N_3192,N_995,N_2041);
nand U3193 (N_3193,N_353,N_2775);
nor U3194 (N_3194,N_936,N_2);
nand U3195 (N_3195,N_1996,N_2224);
and U3196 (N_3196,N_1986,N_1323);
nor U3197 (N_3197,N_1847,N_812);
or U3198 (N_3198,N_2867,N_2163);
or U3199 (N_3199,N_2174,N_714);
nor U3200 (N_3200,N_2346,N_2544);
or U3201 (N_3201,N_2874,N_115);
nand U3202 (N_3202,N_805,N_2407);
nand U3203 (N_3203,N_2021,N_2519);
and U3204 (N_3204,N_709,N_1484);
nor U3205 (N_3205,N_244,N_1240);
and U3206 (N_3206,N_2725,N_1542);
xnor U3207 (N_3207,N_829,N_1564);
nand U3208 (N_3208,N_1877,N_613);
nand U3209 (N_3209,N_509,N_869);
and U3210 (N_3210,N_1655,N_1777);
nand U3211 (N_3211,N_1396,N_484);
nor U3212 (N_3212,N_2813,N_2916);
nand U3213 (N_3213,N_2796,N_769);
and U3214 (N_3214,N_1681,N_109);
or U3215 (N_3215,N_914,N_1898);
nand U3216 (N_3216,N_2056,N_1458);
or U3217 (N_3217,N_35,N_2430);
or U3218 (N_3218,N_2766,N_1470);
nor U3219 (N_3219,N_2798,N_2138);
nand U3220 (N_3220,N_2809,N_572);
or U3221 (N_3221,N_1023,N_790);
and U3222 (N_3222,N_1102,N_2552);
xor U3223 (N_3223,N_1269,N_1097);
or U3224 (N_3224,N_2084,N_524);
and U3225 (N_3225,N_1162,N_896);
nor U3226 (N_3226,N_1666,N_2997);
and U3227 (N_3227,N_1459,N_1940);
nor U3228 (N_3228,N_1293,N_1927);
nand U3229 (N_3229,N_1203,N_1151);
nand U3230 (N_3230,N_955,N_2435);
and U3231 (N_3231,N_1232,N_2599);
nor U3232 (N_3232,N_2696,N_2953);
nor U3233 (N_3233,N_1808,N_464);
nand U3234 (N_3234,N_167,N_1557);
nor U3235 (N_3235,N_2855,N_1013);
nand U3236 (N_3236,N_1546,N_2153);
or U3237 (N_3237,N_1382,N_2852);
and U3238 (N_3238,N_1465,N_973);
nand U3239 (N_3239,N_25,N_1796);
and U3240 (N_3240,N_1274,N_919);
nor U3241 (N_3241,N_2146,N_1036);
nand U3242 (N_3242,N_2710,N_332);
nand U3243 (N_3243,N_113,N_691);
and U3244 (N_3244,N_310,N_1983);
nor U3245 (N_3245,N_1998,N_1329);
nand U3246 (N_3246,N_784,N_2393);
and U3247 (N_3247,N_527,N_927);
nor U3248 (N_3248,N_2604,N_1579);
nor U3249 (N_3249,N_1200,N_2651);
or U3250 (N_3250,N_2497,N_1846);
nor U3251 (N_3251,N_740,N_186);
or U3252 (N_3252,N_2929,N_2199);
nor U3253 (N_3253,N_1660,N_787);
nor U3254 (N_3254,N_467,N_2649);
and U3255 (N_3255,N_2957,N_870);
or U3256 (N_3256,N_2942,N_1489);
nand U3257 (N_3257,N_334,N_1668);
nor U3258 (N_3258,N_2644,N_578);
nand U3259 (N_3259,N_1888,N_600);
nor U3260 (N_3260,N_2716,N_795);
nor U3261 (N_3261,N_2256,N_1601);
and U3262 (N_3262,N_2203,N_2312);
nor U3263 (N_3263,N_2597,N_705);
and U3264 (N_3264,N_724,N_2951);
nand U3265 (N_3265,N_716,N_617);
nor U3266 (N_3266,N_697,N_204);
or U3267 (N_3267,N_916,N_2046);
and U3268 (N_3268,N_2923,N_2052);
nand U3269 (N_3269,N_2881,N_1772);
xor U3270 (N_3270,N_847,N_471);
and U3271 (N_3271,N_1257,N_749);
and U3272 (N_3272,N_2687,N_2587);
or U3273 (N_3273,N_240,N_2821);
or U3274 (N_3274,N_490,N_2158);
nand U3275 (N_3275,N_2156,N_2704);
nand U3276 (N_3276,N_350,N_292);
nor U3277 (N_3277,N_535,N_2069);
nand U3278 (N_3278,N_2563,N_1556);
nand U3279 (N_3279,N_690,N_591);
nor U3280 (N_3280,N_50,N_262);
and U3281 (N_3281,N_2094,N_2814);
and U3282 (N_3282,N_917,N_1812);
nand U3283 (N_3283,N_2062,N_862);
and U3284 (N_3284,N_2621,N_321);
or U3285 (N_3285,N_772,N_1547);
and U3286 (N_3286,N_1143,N_565);
and U3287 (N_3287,N_750,N_1900);
or U3288 (N_3288,N_1803,N_2523);
and U3289 (N_3289,N_1587,N_102);
and U3290 (N_3290,N_2076,N_460);
nor U3291 (N_3291,N_2641,N_1817);
or U3292 (N_3292,N_620,N_506);
nand U3293 (N_3293,N_1995,N_842);
xnor U3294 (N_3294,N_440,N_519);
and U3295 (N_3295,N_2104,N_1416);
or U3296 (N_3296,N_256,N_2648);
and U3297 (N_3297,N_1380,N_129);
nor U3298 (N_3298,N_1292,N_584);
or U3299 (N_3299,N_2529,N_1575);
and U3300 (N_3300,N_217,N_1897);
and U3301 (N_3301,N_681,N_465);
nand U3302 (N_3302,N_1848,N_655);
nand U3303 (N_3303,N_2734,N_47);
nor U3304 (N_3304,N_2762,N_238);
or U3305 (N_3305,N_2728,N_2463);
and U3306 (N_3306,N_2899,N_554);
and U3307 (N_3307,N_156,N_1937);
nor U3308 (N_3308,N_2534,N_1704);
and U3309 (N_3309,N_643,N_1756);
nand U3310 (N_3310,N_2843,N_2996);
nor U3311 (N_3311,N_966,N_1492);
nor U3312 (N_3312,N_1016,N_2538);
and U3313 (N_3313,N_2134,N_2787);
or U3314 (N_3314,N_379,N_890);
and U3315 (N_3315,N_2290,N_2526);
and U3316 (N_3316,N_1933,N_505);
nand U3317 (N_3317,N_789,N_296);
and U3318 (N_3318,N_69,N_54);
nand U3319 (N_3319,N_640,N_811);
or U3320 (N_3320,N_674,N_68);
and U3321 (N_3321,N_2294,N_2659);
and U3322 (N_3322,N_1829,N_1389);
nor U3323 (N_3323,N_830,N_171);
and U3324 (N_3324,N_2888,N_213);
or U3325 (N_3325,N_1990,N_73);
or U3326 (N_3326,N_1527,N_1550);
and U3327 (N_3327,N_308,N_92);
nor U3328 (N_3328,N_579,N_1502);
and U3329 (N_3329,N_1225,N_2103);
xor U3330 (N_3330,N_1048,N_1789);
nor U3331 (N_3331,N_2161,N_2536);
and U3332 (N_3332,N_2272,N_885);
or U3333 (N_3333,N_1137,N_1816);
nand U3334 (N_3334,N_2259,N_160);
nand U3335 (N_3335,N_1923,N_1038);
nand U3336 (N_3336,N_2253,N_64);
and U3337 (N_3337,N_2498,N_2187);
or U3338 (N_3338,N_998,N_212);
nand U3339 (N_3339,N_1745,N_2044);
nand U3340 (N_3340,N_1241,N_1321);
nor U3341 (N_3341,N_2003,N_77);
nand U3342 (N_3342,N_866,N_2959);
nor U3343 (N_3343,N_1173,N_1442);
nand U3344 (N_3344,N_2201,N_2113);
and U3345 (N_3345,N_2302,N_96);
and U3346 (N_3346,N_2987,N_887);
nor U3347 (N_3347,N_2193,N_2703);
or U3348 (N_3348,N_889,N_779);
nand U3349 (N_3349,N_1002,N_734);
nand U3350 (N_3350,N_245,N_577);
nor U3351 (N_3351,N_2375,N_1124);
nor U3352 (N_3352,N_195,N_2940);
nand U3353 (N_3353,N_1077,N_1065);
or U3354 (N_3354,N_1387,N_2243);
or U3355 (N_3355,N_342,N_2826);
nor U3356 (N_3356,N_1368,N_2212);
nor U3357 (N_3357,N_257,N_863);
or U3358 (N_3358,N_683,N_2578);
nand U3359 (N_3359,N_637,N_2781);
nand U3360 (N_3360,N_798,N_972);
nand U3361 (N_3361,N_1874,N_399);
nand U3362 (N_3362,N_2247,N_2706);
nand U3363 (N_3363,N_1593,N_2580);
or U3364 (N_3364,N_1117,N_2854);
nand U3365 (N_3365,N_2226,N_2918);
and U3366 (N_3366,N_832,N_272);
or U3367 (N_3367,N_1483,N_1346);
nand U3368 (N_3368,N_1490,N_2709);
nand U3369 (N_3369,N_114,N_2754);
nor U3370 (N_3370,N_733,N_2635);
nor U3371 (N_3371,N_477,N_1555);
or U3372 (N_3372,N_421,N_149);
nor U3373 (N_3373,N_201,N_1678);
nor U3374 (N_3374,N_2196,N_63);
or U3375 (N_3375,N_2624,N_260);
nor U3376 (N_3376,N_7,N_1069);
nand U3377 (N_3377,N_1186,N_1473);
nand U3378 (N_3378,N_2974,N_2305);
or U3379 (N_3379,N_1724,N_689);
and U3380 (N_3380,N_2688,N_1076);
or U3381 (N_3381,N_2325,N_335);
and U3382 (N_3382,N_1980,N_2147);
nand U3383 (N_3383,N_561,N_166);
and U3384 (N_3384,N_1576,N_943);
and U3385 (N_3385,N_1295,N_1733);
or U3386 (N_3386,N_1320,N_548);
nor U3387 (N_3387,N_207,N_1973);
nor U3388 (N_3388,N_2815,N_2336);
or U3389 (N_3389,N_2832,N_1319);
nand U3390 (N_3390,N_1429,N_1842);
and U3391 (N_3391,N_402,N_1385);
nand U3392 (N_3392,N_1170,N_2522);
or U3393 (N_3393,N_1000,N_1464);
or U3394 (N_3394,N_553,N_2573);
or U3395 (N_3395,N_1534,N_2303);
or U3396 (N_3396,N_162,N_1227);
nand U3397 (N_3397,N_1341,N_1469);
nand U3398 (N_3398,N_347,N_2810);
xor U3399 (N_3399,N_1280,N_2295);
nor U3400 (N_3400,N_1083,N_1155);
or U3401 (N_3401,N_746,N_1330);
and U3402 (N_3402,N_76,N_976);
or U3403 (N_3403,N_275,N_2489);
nor U3404 (N_3404,N_155,N_949);
or U3405 (N_3405,N_1093,N_3);
and U3406 (N_3406,N_2876,N_290);
nand U3407 (N_3407,N_954,N_1437);
and U3408 (N_3408,N_237,N_39);
nor U3409 (N_3409,N_2773,N_462);
or U3410 (N_3410,N_1188,N_121);
nor U3411 (N_3411,N_2958,N_2844);
nor U3412 (N_3412,N_533,N_297);
and U3413 (N_3413,N_956,N_1974);
nor U3414 (N_3414,N_2960,N_1235);
or U3415 (N_3415,N_2565,N_1946);
or U3416 (N_3416,N_682,N_2611);
nor U3417 (N_3417,N_2977,N_1163);
or U3418 (N_3418,N_942,N_1876);
or U3419 (N_3419,N_2457,N_81);
or U3420 (N_3420,N_2307,N_2209);
or U3421 (N_3421,N_1426,N_2771);
or U3422 (N_3422,N_2717,N_806);
or U3423 (N_3423,N_2338,N_2350);
nand U3424 (N_3424,N_403,N_411);
or U3425 (N_3425,N_2206,N_568);
or U3426 (N_3426,N_315,N_2639);
nand U3427 (N_3427,N_2053,N_2758);
nor U3428 (N_3428,N_1003,N_580);
nand U3429 (N_3429,N_576,N_46);
nor U3430 (N_3430,N_765,N_939);
nand U3431 (N_3431,N_2109,N_2556);
or U3432 (N_3432,N_1500,N_1818);
nor U3433 (N_3433,N_2462,N_1410);
or U3434 (N_3434,N_657,N_2366);
and U3435 (N_3435,N_1809,N_796);
nor U3436 (N_3436,N_2445,N_1922);
nor U3437 (N_3437,N_1971,N_2595);
and U3438 (N_3438,N_215,N_1011);
xor U3439 (N_3439,N_1977,N_744);
nand U3440 (N_3440,N_1433,N_780);
nand U3441 (N_3441,N_313,N_473);
or U3442 (N_3442,N_2746,N_2011);
and U3443 (N_3443,N_1709,N_822);
or U3444 (N_3444,N_2208,N_1746);
or U3445 (N_3445,N_1684,N_67);
and U3446 (N_3446,N_306,N_2506);
nand U3447 (N_3447,N_1273,N_48);
and U3448 (N_3448,N_1635,N_928);
or U3449 (N_3449,N_446,N_2005);
and U3450 (N_3450,N_1112,N_592);
nor U3451 (N_3451,N_978,N_1830);
nand U3452 (N_3452,N_2875,N_458);
nand U3453 (N_3453,N_901,N_2330);
and U3454 (N_3454,N_2081,N_264);
nand U3455 (N_3455,N_2562,N_2926);
nand U3456 (N_3456,N_921,N_2829);
and U3457 (N_3457,N_2019,N_1248);
nand U3458 (N_3458,N_317,N_2950);
or U3459 (N_3459,N_2789,N_309);
nand U3460 (N_3460,N_376,N_585);
or U3461 (N_3461,N_501,N_853);
nor U3462 (N_3462,N_2753,N_428);
or U3463 (N_3463,N_1272,N_2141);
or U3464 (N_3464,N_70,N_1);
or U3465 (N_3465,N_1454,N_940);
or U3466 (N_3466,N_931,N_176);
nand U3467 (N_3467,N_630,N_1044);
nor U3468 (N_3468,N_2219,N_1401);
or U3469 (N_3469,N_1641,N_930);
and U3470 (N_3470,N_1916,N_963);
and U3471 (N_3471,N_1960,N_867);
nor U3472 (N_3472,N_849,N_418);
nor U3473 (N_3473,N_1440,N_302);
or U3474 (N_3474,N_1386,N_2397);
and U3475 (N_3475,N_1836,N_1398);
and U3476 (N_3476,N_607,N_2994);
nor U3477 (N_3477,N_105,N_582);
nand U3478 (N_3478,N_1311,N_2833);
nand U3479 (N_3479,N_1999,N_2862);
and U3480 (N_3480,N_2010,N_140);
and U3481 (N_3481,N_1056,N_329);
nand U3482 (N_3482,N_864,N_1725);
or U3483 (N_3483,N_144,N_2811);
and U3484 (N_3484,N_615,N_1338);
nor U3485 (N_3485,N_2136,N_502);
or U3486 (N_3486,N_2945,N_2507);
or U3487 (N_3487,N_346,N_336);
nor U3488 (N_3488,N_771,N_2588);
and U3489 (N_3489,N_2827,N_1471);
and U3490 (N_3490,N_824,N_2438);
and U3491 (N_3491,N_2433,N_563);
nand U3492 (N_3492,N_1518,N_1680);
nand U3493 (N_3493,N_2776,N_2200);
and U3494 (N_3494,N_1135,N_137);
nand U3495 (N_3495,N_2975,N_2218);
nand U3496 (N_3496,N_1318,N_1853);
nand U3497 (N_3497,N_1087,N_1524);
nand U3498 (N_3498,N_1530,N_1236);
nand U3499 (N_3499,N_1246,N_510);
nand U3500 (N_3500,N_2252,N_2695);
or U3501 (N_3501,N_1275,N_1820);
or U3502 (N_3502,N_2143,N_1478);
or U3503 (N_3503,N_2782,N_1160);
nor U3504 (N_3504,N_1648,N_470);
nand U3505 (N_3505,N_2245,N_1242);
or U3506 (N_3506,N_1769,N_178);
and U3507 (N_3507,N_1128,N_2995);
or U3508 (N_3508,N_439,N_277);
nand U3509 (N_3509,N_53,N_1030);
and U3510 (N_3510,N_226,N_2391);
or U3511 (N_3511,N_2665,N_952);
nor U3512 (N_3512,N_2490,N_1111);
nor U3513 (N_3513,N_28,N_661);
and U3514 (N_3514,N_1972,N_2516);
and U3515 (N_3515,N_1515,N_1722);
nor U3516 (N_3516,N_291,N_962);
or U3517 (N_3517,N_2097,N_650);
xnor U3518 (N_3518,N_1926,N_2265);
and U3519 (N_3519,N_594,N_2904);
nand U3520 (N_3520,N_181,N_202);
nand U3521 (N_3521,N_2828,N_2616);
nand U3522 (N_3522,N_2287,N_737);
nand U3523 (N_3523,N_269,N_1351);
nor U3524 (N_3524,N_1802,N_722);
nand U3525 (N_3525,N_816,N_1969);
or U3526 (N_3526,N_2261,N_2878);
nand U3527 (N_3527,N_120,N_933);
nor U3528 (N_3528,N_1425,N_1707);
and U3529 (N_3529,N_1510,N_487);
nor U3530 (N_3530,N_2927,N_2049);
and U3531 (N_3531,N_22,N_1460);
and U3532 (N_3532,N_2877,N_193);
or U3533 (N_3533,N_360,N_2576);
and U3534 (N_3534,N_649,N_396);
nor U3535 (N_3535,N_926,N_2839);
nor U3536 (N_3536,N_414,N_243);
nor U3537 (N_3537,N_354,N_626);
nand U3538 (N_3538,N_2448,N_1233);
or U3539 (N_3539,N_2152,N_1651);
and U3540 (N_3540,N_2871,N_1728);
nand U3541 (N_3541,N_900,N_522);
nor U3542 (N_3542,N_200,N_1921);
nand U3543 (N_3543,N_1090,N_2311);
or U3544 (N_3544,N_1834,N_1216);
and U3545 (N_3545,N_1183,N_247);
and U3546 (N_3546,N_1697,N_2425);
nor U3547 (N_3547,N_755,N_2155);
nor U3548 (N_3548,N_14,N_93);
or U3549 (N_3549,N_2629,N_1497);
and U3550 (N_3550,N_1190,N_1698);
nor U3551 (N_3551,N_280,N_33);
or U3552 (N_3552,N_2484,N_1545);
nand U3553 (N_3553,N_2807,N_450);
and U3554 (N_3554,N_2202,N_667);
nor U3555 (N_3555,N_1907,N_136);
nor U3556 (N_3556,N_979,N_837);
nor U3557 (N_3557,N_2535,N_1823);
nand U3558 (N_3558,N_1182,N_2007);
nor U3559 (N_3559,N_1526,N_873);
nand U3560 (N_3560,N_793,N_588);
or U3561 (N_3561,N_528,N_1549);
nor U3562 (N_3562,N_2986,N_761);
and U3563 (N_3563,N_1522,N_1932);
nand U3564 (N_3564,N_1711,N_323);
and U3565 (N_3565,N_1644,N_1408);
or U3566 (N_3566,N_622,N_2418);
nor U3567 (N_3567,N_748,N_2965);
or U3568 (N_3568,N_612,N_967);
nor U3569 (N_3569,N_2784,N_224);
nand U3570 (N_3570,N_365,N_1778);
nand U3571 (N_3571,N_2115,N_2157);
and U3572 (N_3572,N_1732,N_1206);
and U3573 (N_3573,N_1250,N_1328);
nand U3574 (N_3574,N_2868,N_1133);
nand U3575 (N_3575,N_1645,N_2568);
nand U3576 (N_3576,N_1418,N_1255);
and U3577 (N_3577,N_2315,N_2437);
and U3578 (N_3578,N_507,N_1787);
and U3579 (N_3579,N_2415,N_2172);
or U3580 (N_3580,N_1159,N_2557);
and U3581 (N_3581,N_1075,N_123);
nand U3582 (N_3582,N_2125,N_633);
and U3583 (N_3583,N_1348,N_1024);
nand U3584 (N_3584,N_729,N_2456);
nand U3585 (N_3585,N_124,N_1525);
nand U3586 (N_3586,N_503,N_2779);
nor U3587 (N_3587,N_875,N_409);
nand U3588 (N_3588,N_1161,N_1239);
and U3589 (N_3589,N_2610,N_1175);
or U3590 (N_3590,N_2306,N_720);
or U3591 (N_3591,N_1064,N_2185);
nand U3592 (N_3592,N_2471,N_2799);
nand U3593 (N_3593,N_2902,N_1867);
or U3594 (N_3594,N_2451,N_886);
nand U3595 (N_3595,N_2235,N_38);
or U3596 (N_3596,N_1503,N_2137);
and U3597 (N_3597,N_2173,N_2220);
nand U3598 (N_3598,N_2653,N_1551);
nand U3599 (N_3599,N_2847,N_372);
and U3600 (N_3600,N_669,N_702);
nor U3601 (N_3601,N_2909,N_1450);
and U3602 (N_3602,N_419,N_2275);
or U3603 (N_3603,N_2964,N_2797);
or U3604 (N_3604,N_2486,N_482);
nor U3605 (N_3605,N_197,N_1866);
nor U3606 (N_3606,N_2192,N_624);
and U3607 (N_3607,N_2546,N_1887);
nand U3608 (N_3608,N_2750,N_2702);
nor U3609 (N_3609,N_1811,N_1055);
and U3610 (N_3610,N_1068,N_562);
or U3611 (N_3611,N_2656,N_1879);
and U3612 (N_3612,N_422,N_1174);
and U3613 (N_3613,N_988,N_1285);
nand U3614 (N_3614,N_2778,N_1270);
nand U3615 (N_3615,N_2110,N_2882);
nand U3616 (N_3616,N_369,N_2459);
nor U3617 (N_3617,N_2505,N_656);
or U3618 (N_3618,N_320,N_1560);
or U3619 (N_3619,N_2991,N_2009);
nand U3620 (N_3620,N_2367,N_386);
nand U3621 (N_3621,N_2033,N_267);
nand U3622 (N_3622,N_2441,N_2405);
nand U3623 (N_3623,N_2057,N_1360);
nor U3624 (N_3624,N_233,N_2064);
or U3625 (N_3625,N_72,N_2026);
or U3626 (N_3626,N_721,N_1189);
nand U3627 (N_3627,N_2714,N_2061);
nor U3628 (N_3628,N_2731,N_623);
nand U3629 (N_3629,N_1687,N_286);
and U3630 (N_3630,N_2620,N_49);
nor U3631 (N_3631,N_2609,N_1832);
and U3632 (N_3632,N_1505,N_974);
nand U3633 (N_3633,N_29,N_903);
nand U3634 (N_3634,N_2030,N_2712);
nor U3635 (N_3635,N_2318,N_94);
nor U3636 (N_3636,N_831,N_1451);
nor U3637 (N_3637,N_2402,N_281);
or U3638 (N_3638,N_2893,N_838);
and U3639 (N_3639,N_1297,N_1992);
nand U3640 (N_3640,N_1122,N_1509);
or U3641 (N_3641,N_1799,N_438);
nand U3642 (N_3642,N_1513,N_2210);
nand U3643 (N_3643,N_410,N_2642);
nand U3644 (N_3644,N_1903,N_841);
or U3645 (N_3645,N_1198,N_2020);
nor U3646 (N_3646,N_4,N_2723);
and U3647 (N_3647,N_808,N_1917);
and U3648 (N_3648,N_937,N_2678);
and U3649 (N_3649,N_540,N_457);
or U3650 (N_3650,N_2607,N_59);
nor U3651 (N_3651,N_1506,N_2673);
and U3652 (N_3652,N_1804,N_2014);
nand U3653 (N_3653,N_1181,N_687);
and U3654 (N_3654,N_1207,N_393);
nor U3655 (N_3655,N_2655,N_1424);
and U3656 (N_3656,N_1156,N_128);
nor U3657 (N_3657,N_2040,N_1588);
nand U3658 (N_3658,N_2099,N_434);
or U3659 (N_3659,N_1028,N_1362);
and U3660 (N_3660,N_2263,N_1826);
nor U3661 (N_3661,N_1642,N_444);
nor U3662 (N_3662,N_2075,N_241);
nand U3663 (N_3663,N_1739,N_441);
nand U3664 (N_3664,N_2972,N_2623);
and U3665 (N_3665,N_508,N_2671);
nor U3666 (N_3666,N_1649,N_523);
and U3667 (N_3667,N_1378,N_1256);
nand U3668 (N_3668,N_935,N_1158);
and U3669 (N_3669,N_760,N_2424);
nand U3670 (N_3670,N_2145,N_139);
nand U3671 (N_3671,N_2528,N_2399);
nand U3672 (N_3672,N_431,N_89);
nor U3673 (N_3673,N_424,N_785);
and U3674 (N_3674,N_2683,N_420);
or U3675 (N_3675,N_814,N_1858);
and U3676 (N_3676,N_225,N_1130);
or U3677 (N_3677,N_1614,N_1040);
nor U3678 (N_3678,N_1701,N_2344);
and U3679 (N_3679,N_1763,N_823);
or U3680 (N_3680,N_2675,N_2419);
nand U3681 (N_3681,N_2654,N_2432);
and U3682 (N_3682,N_235,N_1785);
nand U3683 (N_3683,N_362,N_98);
or U3684 (N_3684,N_587,N_2035);
nand U3685 (N_3685,N_994,N_2022);
and U3686 (N_3686,N_150,N_1833);
nor U3687 (N_3687,N_888,N_1540);
nor U3688 (N_3688,N_1363,N_1327);
nor U3689 (N_3689,N_1199,N_839);
or U3690 (N_3690,N_969,N_1636);
and U3691 (N_3691,N_636,N_2329);
and U3692 (N_3692,N_2183,N_1611);
and U3693 (N_3693,N_1402,N_704);
or U3694 (N_3694,N_570,N_1734);
and U3695 (N_3695,N_65,N_688);
nand U3696 (N_3696,N_1394,N_2707);
nand U3697 (N_3697,N_2949,N_1523);
or U3698 (N_3698,N_1204,N_1567);
or U3699 (N_3699,N_1548,N_1107);
nor U3700 (N_3700,N_1904,N_2077);
and U3701 (N_3701,N_2761,N_2510);
and U3702 (N_3702,N_239,N_2442);
or U3703 (N_3703,N_2980,N_1596);
and U3704 (N_3704,N_1307,N_2051);
nor U3705 (N_3705,N_104,N_879);
nor U3706 (N_3706,N_1741,N_1214);
and U3707 (N_3707,N_2426,N_2645);
nand U3708 (N_3708,N_586,N_1885);
and U3709 (N_3709,N_2039,N_2313);
nor U3710 (N_3710,N_2319,N_1566);
nand U3711 (N_3711,N_1531,N_1754);
and U3712 (N_3712,N_675,N_2617);
nor U3713 (N_3713,N_2713,N_2343);
nor U3714 (N_3714,N_355,N_1053);
nor U3715 (N_3715,N_2735,N_1788);
nand U3716 (N_3716,N_2768,N_2806);
and U3717 (N_3717,N_957,N_2664);
nor U3718 (N_3718,N_2301,N_206);
and U3719 (N_3719,N_1951,N_1060);
or U3720 (N_3720,N_1476,N_1831);
nor U3721 (N_3721,N_665,N_2755);
nand U3722 (N_3722,N_631,N_11);
nand U3723 (N_3723,N_2637,N_857);
nor U3724 (N_3724,N_1767,N_2258);
and U3725 (N_3725,N_2361,N_2162);
nor U3726 (N_3726,N_2002,N_614);
nor U3727 (N_3727,N_2297,N_1621);
and U3728 (N_3728,N_2140,N_390);
nor U3729 (N_3729,N_2860,N_97);
and U3730 (N_3730,N_1956,N_2170);
nor U3731 (N_3731,N_529,N_1141);
and U3732 (N_3732,N_2205,N_1101);
nand U3733 (N_3733,N_1828,N_1496);
nor U3734 (N_3734,N_2582,N_601);
nor U3735 (N_3735,N_2674,N_1100);
or U3736 (N_3736,N_1084,N_1349);
nand U3737 (N_3737,N_2701,N_759);
and U3738 (N_3738,N_2889,N_1054);
or U3739 (N_3739,N_2594,N_1646);
nand U3740 (N_3740,N_159,N_250);
nor U3741 (N_3741,N_2816,N_1017);
nand U3742 (N_3742,N_2747,N_2310);
or U3743 (N_3743,N_1825,N_2298);
nand U3744 (N_3744,N_40,N_756);
nand U3745 (N_3745,N_1364,N_2906);
nand U3746 (N_3746,N_1372,N_608);
or U3747 (N_3747,N_2988,N_556);
nand U3748 (N_3748,N_1220,N_1337);
nand U3749 (N_3749,N_2142,N_2705);
or U3750 (N_3750,N_1192,N_363);
and U3751 (N_3751,N_2791,N_1196);
and U3752 (N_3752,N_2197,N_1582);
nand U3753 (N_3753,N_248,N_2898);
and U3754 (N_3754,N_1029,N_2818);
nand U3755 (N_3755,N_904,N_2941);
or U3756 (N_3756,N_751,N_1689);
nor U3757 (N_3757,N_2931,N_2513);
nor U3758 (N_3758,N_1813,N_2938);
nand U3759 (N_3759,N_316,N_51);
nor U3760 (N_3760,N_991,N_1067);
nand U3761 (N_3761,N_534,N_2121);
or U3762 (N_3762,N_1006,N_348);
nand U3763 (N_3763,N_2933,N_2333);
and U3764 (N_3764,N_752,N_1726);
nand U3765 (N_3765,N_638,N_1947);
and U3766 (N_3766,N_2055,N_163);
or U3767 (N_3767,N_2299,N_103);
nor U3768 (N_3768,N_742,N_1357);
or U3769 (N_3769,N_632,N_2222);
and U3770 (N_3770,N_2679,N_2947);
nor U3771 (N_3771,N_2542,N_2169);
nand U3772 (N_3772,N_2700,N_1176);
nand U3773 (N_3773,N_1520,N_495);
nand U3774 (N_3774,N_2892,N_1194);
and U3775 (N_3775,N_469,N_1118);
nand U3776 (N_3776,N_454,N_106);
or U3777 (N_3777,N_1178,N_2511);
or U3778 (N_3778,N_383,N_388);
nand U3779 (N_3779,N_227,N_668);
and U3780 (N_3780,N_2470,N_906);
nand U3781 (N_3781,N_1961,N_850);
nor U3782 (N_3782,N_408,N_1462);
nor U3783 (N_3783,N_95,N_151);
nand U3784 (N_3784,N_2567,N_2928);
nor U3785 (N_3785,N_514,N_1935);
nand U3786 (N_3786,N_1370,N_188);
and U3787 (N_3787,N_1875,N_2335);
nand U3788 (N_3788,N_2429,N_2122);
and U3789 (N_3789,N_609,N_2912);
nand U3790 (N_3790,N_999,N_2070);
nand U3791 (N_3791,N_1737,N_2634);
or U3792 (N_3792,N_1290,N_2591);
or U3793 (N_3793,N_711,N_2188);
nor U3794 (N_3794,N_1092,N_2527);
and U3795 (N_3795,N_1359,N_521);
nand U3796 (N_3796,N_2584,N_757);
or U3797 (N_3797,N_1790,N_2549);
or U3798 (N_3798,N_810,N_971);
nor U3799 (N_3799,N_1750,N_1852);
nand U3800 (N_3800,N_20,N_118);
or U3801 (N_3801,N_1631,N_461);
and U3802 (N_3802,N_2543,N_180);
nor U3803 (N_3803,N_2180,N_2545);
nor U3804 (N_3804,N_2413,N_1784);
xor U3805 (N_3805,N_1884,N_1712);
nand U3806 (N_3806,N_530,N_476);
nor U3807 (N_3807,N_1208,N_259);
nand U3808 (N_3808,N_1217,N_2764);
or U3809 (N_3809,N_80,N_1623);
nand U3810 (N_3810,N_2171,N_2968);
or U3811 (N_3811,N_2920,N_491);
nor U3812 (N_3812,N_2373,N_791);
and U3813 (N_3813,N_1664,N_1730);
nand U3814 (N_3814,N_1517,N_686);
nor U3815 (N_3815,N_2392,N_1383);
nor U3816 (N_3816,N_593,N_1915);
and U3817 (N_3817,N_2636,N_2460);
nand U3818 (N_3818,N_2291,N_1249);
and U3819 (N_3819,N_725,N_2772);
or U3820 (N_3820,N_513,N_1855);
and U3821 (N_3821,N_2452,N_125);
and U3822 (N_3822,N_2808,N_455);
or U3823 (N_3823,N_1654,N_135);
nand U3824 (N_3824,N_1431,N_1276);
nand U3825 (N_3825,N_2365,N_325);
and U3826 (N_3826,N_2744,N_1335);
xnor U3827 (N_3827,N_2504,N_2233);
or U3828 (N_3828,N_531,N_654);
xnor U3829 (N_3829,N_2101,N_1284);
and U3830 (N_3830,N_977,N_1632);
nand U3831 (N_3831,N_1252,N_2048);
nor U3832 (N_3832,N_738,N_953);
nand U3833 (N_3833,N_1231,N_2618);
nand U3834 (N_3834,N_1819,N_1747);
and U3835 (N_3835,N_876,N_87);
and U3836 (N_3836,N_2627,N_2450);
nor U3837 (N_3837,N_2347,N_2478);
nor U3838 (N_3838,N_1768,N_732);
or U3839 (N_3839,N_1081,N_2284);
or U3840 (N_3840,N_1742,N_1032);
and U3841 (N_3841,N_1775,N_2351);
and U3842 (N_3842,N_2722,N_2592);
or U3843 (N_3843,N_1355,N_1430);
nand U3844 (N_3844,N_255,N_980);
or U3845 (N_3845,N_2001,N_1347);
and U3846 (N_3846,N_1882,N_1309);
nor U3847 (N_3847,N_610,N_2168);
nor U3848 (N_3848,N_1521,N_1753);
or U3849 (N_3849,N_79,N_130);
and U3850 (N_3850,N_1105,N_1258);
nand U3851 (N_3851,N_2322,N_1210);
nand U3852 (N_3852,N_2708,N_417);
nand U3853 (N_3853,N_1931,N_2254);
nand U3854 (N_3854,N_1950,N_881);
nand U3855 (N_3855,N_1373,N_1640);
and U3856 (N_3856,N_2130,N_2488);
or U3857 (N_3857,N_2204,N_1920);
nor U3858 (N_3858,N_246,N_1539);
nor U3859 (N_3859,N_2699,N_2483);
and U3860 (N_3860,N_1670,N_90);
nand U3861 (N_3861,N_2371,N_147);
and U3862 (N_3862,N_710,N_2268);
nand U3863 (N_3863,N_1254,N_2388);
nor U3864 (N_3864,N_489,N_692);
nand U3865 (N_3865,N_2358,N_1066);
or U3866 (N_3866,N_2385,N_2566);
nand U3867 (N_3867,N_2160,N_1943);
and U3868 (N_3868,N_595,N_2553);
or U3869 (N_3869,N_1771,N_289);
nand U3870 (N_3870,N_349,N_2756);
nand U3871 (N_3871,N_1688,N_1108);
or U3872 (N_3872,N_494,N_1008);
or U3873 (N_3873,N_2176,N_1063);
nor U3874 (N_3874,N_2234,N_1125);
or U3875 (N_3875,N_303,N_2107);
nand U3876 (N_3876,N_703,N_34);
nor U3877 (N_3877,N_1629,N_1783);
nor U3878 (N_3878,N_83,N_1251);
and U3879 (N_3879,N_1815,N_1486);
and U3880 (N_3880,N_1317,N_634);
nor U3881 (N_3881,N_2669,N_1201);
and U3882 (N_3882,N_2191,N_877);
nor U3883 (N_3883,N_1202,N_987);
nor U3884 (N_3884,N_715,N_307);
or U3885 (N_3885,N_148,N_2686);
or U3886 (N_3886,N_685,N_1120);
and U3887 (N_3887,N_525,N_0);
nor U3888 (N_3888,N_2428,N_924);
or U3889 (N_3889,N_1864,N_512);
or U3890 (N_3890,N_2532,N_2583);
nor U3891 (N_3891,N_165,N_2148);
nor U3892 (N_3892,N_1149,N_2663);
and U3893 (N_3893,N_2164,N_2792);
nand U3894 (N_3894,N_2461,N_1511);
nor U3895 (N_3895,N_2114,N_1070);
nor U3896 (N_3896,N_330,N_2841);
and U3897 (N_3897,N_2045,N_168);
or U3898 (N_3898,N_913,N_1598);
nand U3899 (N_3899,N_1443,N_852);
nand U3900 (N_3900,N_1228,N_1306);
or U3901 (N_3901,N_1397,N_2439);
nand U3902 (N_3902,N_1116,N_1421);
and U3903 (N_3903,N_283,N_1461);
nand U3904 (N_3904,N_992,N_1119);
or U3905 (N_3905,N_1868,N_300);
nand U3906 (N_3906,N_1034,N_2364);
and U3907 (N_3907,N_274,N_1650);
nand U3908 (N_3908,N_268,N_1607);
and U3909 (N_3909,N_859,N_116);
nor U3910 (N_3910,N_1592,N_1657);
nand U3911 (N_3911,N_800,N_1086);
and U3912 (N_3912,N_1736,N_1358);
nand U3913 (N_3913,N_481,N_2221);
nand U3914 (N_3914,N_2288,N_912);
and U3915 (N_3915,N_2502,N_1166);
nand U3916 (N_3916,N_2100,N_1109);
and U3917 (N_3917,N_2853,N_1896);
and U3918 (N_3918,N_288,N_497);
and U3919 (N_3919,N_1696,N_2998);
or U3920 (N_3920,N_1487,N_1479);
or U3921 (N_3921,N_1865,N_2217);
and U3922 (N_3922,N_1843,N_1978);
nor U3923 (N_3923,N_2085,N_1455);
nand U3924 (N_3924,N_2600,N_146);
or U3925 (N_3925,N_312,N_1994);
or U3926 (N_3926,N_2091,N_2348);
nand U3927 (N_3927,N_874,N_157);
nor U3928 (N_3928,N_1457,N_1403);
and U3929 (N_3929,N_62,N_1740);
and U3930 (N_3930,N_2670,N_775);
nand U3931 (N_3931,N_339,N_2434);
xor U3932 (N_3932,N_2693,N_1814);
or U3933 (N_3933,N_958,N_1435);
nor U3934 (N_3934,N_1690,N_583);
and U3935 (N_3935,N_1637,N_1934);
and U3936 (N_3936,N_2691,N_2018);
or U3937 (N_3937,N_1001,N_2760);
nand U3938 (N_3938,N_2499,N_1303);
or U3939 (N_3939,N_2440,N_2078);
nand U3940 (N_3940,N_2836,N_1719);
or U3941 (N_3941,N_143,N_208);
and U3942 (N_3942,N_1964,N_2096);
nor U3943 (N_3943,N_2248,N_1552);
nand U3944 (N_3944,N_2017,N_2029);
nand U3945 (N_3945,N_2943,N_366);
and U3946 (N_3946,N_960,N_2447);
xor U3947 (N_3947,N_541,N_2660);
or U3948 (N_3948,N_2831,N_327);
or U3949 (N_3949,N_1929,N_322);
or U3950 (N_3950,N_2124,N_2922);
nand U3951 (N_3951,N_783,N_797);
and U3952 (N_3952,N_743,N_2495);
nor U3953 (N_3953,N_406,N_1103);
and U3954 (N_3954,N_1890,N_1332);
nor U3955 (N_3955,N_107,N_2865);
and U3956 (N_3956,N_258,N_2551);
nor U3957 (N_3957,N_560,N_2907);
nor U3958 (N_3958,N_2963,N_1296);
nand U3959 (N_3959,N_459,N_357);
and U3960 (N_3960,N_2334,N_2586);
or U3961 (N_3961,N_1849,N_1267);
nor U3962 (N_3962,N_442,N_559);
and U3963 (N_3963,N_498,N_58);
nor U3964 (N_3964,N_1770,N_1447);
and U3965 (N_3965,N_2682,N_1762);
nor U3966 (N_3966,N_1639,N_700);
and U3967 (N_3967,N_2903,N_333);
and U3968 (N_3968,N_1104,N_1909);
or U3969 (N_3969,N_205,N_2840);
and U3970 (N_3970,N_2257,N_2743);
and U3971 (N_3971,N_2281,N_2274);
xnor U3972 (N_3972,N_145,N_997);
or U3973 (N_3973,N_375,N_574);
and U3974 (N_3974,N_1695,N_1633);
or U3975 (N_3975,N_1672,N_723);
or U3976 (N_3976,N_844,N_1395);
nor U3977 (N_3977,N_295,N_642);
nor U3978 (N_3978,N_2105,N_61);
or U3979 (N_3979,N_736,N_2127);
and U3980 (N_3980,N_2540,N_735);
nor U3981 (N_3981,N_2032,N_1288);
and U3982 (N_3982,N_825,N_1079);
nor U3983 (N_3983,N_2672,N_1493);
or U3984 (N_3984,N_1422,N_86);
nor U3985 (N_3985,N_2345,N_2167);
or U3986 (N_3986,N_1743,N_2068);
and U3987 (N_3987,N_2042,N_1088);
or U3988 (N_3988,N_2304,N_1599);
or U3989 (N_3989,N_1507,N_659);
nor U3990 (N_3990,N_305,N_950);
nor U3991 (N_3991,N_2266,N_2622);
nand U3992 (N_3992,N_922,N_1168);
nor U3993 (N_3993,N_1110,N_1794);
or U3994 (N_3994,N_2978,N_834);
or U3995 (N_3995,N_1191,N_684);
nand U3996 (N_3996,N_2823,N_2067);
nor U3997 (N_3997,N_2790,N_1218);
nor U3998 (N_3998,N_1871,N_2646);
and U3999 (N_3999,N_1609,N_2866);
nor U4000 (N_4000,N_828,N_2036);
nand U4001 (N_4001,N_1872,N_1989);
or U4002 (N_4002,N_1039,N_2332);
and U4003 (N_4003,N_1643,N_2106);
and U4004 (N_4004,N_1018,N_1144);
or U4005 (N_4005,N_1841,N_2126);
or U4006 (N_4006,N_299,N_2752);
nand U4007 (N_4007,N_717,N_345);
nor U4008 (N_4008,N_2684,N_1744);
and U4009 (N_4009,N_331,N_483);
and U4010 (N_4010,N_2251,N_2031);
or U4011 (N_4011,N_1420,N_184);
nor U4012 (N_4012,N_1262,N_1308);
or U4013 (N_4013,N_2154,N_1968);
and U4014 (N_4014,N_273,N_663);
or U4015 (N_4015,N_2037,N_2612);
or U4016 (N_4016,N_2177,N_1485);
nor U4017 (N_4017,N_1057,N_2948);
and U4018 (N_4018,N_2895,N_1446);
or U4019 (N_4019,N_2554,N_285);
or U4020 (N_4020,N_2736,N_1139);
nand U4021 (N_4021,N_100,N_2494);
nor U4022 (N_4022,N_1616,N_1676);
nor U4023 (N_4023,N_845,N_1718);
nor U4024 (N_4024,N_1910,N_2512);
and U4025 (N_4025,N_695,N_1271);
nor U4026 (N_4026,N_2626,N_511);
nand U4027 (N_4027,N_222,N_2314);
or U4028 (N_4028,N_762,N_41);
and U4029 (N_4029,N_253,N_1154);
or U4030 (N_4030,N_2932,N_2093);
nor U4031 (N_4031,N_1356,N_1312);
and U4032 (N_4032,N_56,N_2491);
and U4033 (N_4033,N_1388,N_463);
or U4034 (N_4034,N_119,N_2276);
xnor U4035 (N_4035,N_2979,N_2227);
nor U4036 (N_4036,N_492,N_2737);
nand U4037 (N_4037,N_1062,N_802);
and U4038 (N_4038,N_230,N_1140);
nor U4039 (N_4039,N_499,N_279);
nor U4040 (N_4040,N_1266,N_1691);
or U4041 (N_4041,N_1180,N_635);
or U4042 (N_4042,N_1997,N_2468);
and U4043 (N_4043,N_2008,N_298);
nand U4044 (N_4044,N_2872,N_2521);
nand U4045 (N_4045,N_1211,N_1938);
nand U4046 (N_4046,N_447,N_2520);
nand U4047 (N_4047,N_404,N_2230);
or U4048 (N_4048,N_382,N_1991);
nand U4049 (N_4049,N_1682,N_516);
nand U4050 (N_4050,N_1047,N_573);
and U4051 (N_4051,N_2803,N_2905);
and U4052 (N_4052,N_2228,N_2555);
nor U4053 (N_4053,N_1757,N_1573);
or U4054 (N_4054,N_2738,N_194);
and U4055 (N_4055,N_621,N_1342);
and U4056 (N_4056,N_2718,N_2059);
nor U4057 (N_4057,N_1602,N_1955);
nor U4058 (N_4058,N_385,N_984);
nor U4059 (N_4059,N_2515,N_2751);
nor U4060 (N_4060,N_1445,N_284);
nor U4061 (N_4061,N_713,N_1886);
nand U4062 (N_4062,N_2412,N_1014);
or U4063 (N_4063,N_1565,N_1970);
nand U4064 (N_4064,N_1911,N_294);
and U4065 (N_4065,N_2255,N_1979);
nand U4066 (N_4066,N_2603,N_596);
and U4067 (N_4067,N_856,N_373);
or U4068 (N_4068,N_175,N_1630);
or U4069 (N_4069,N_719,N_293);
or U4070 (N_4070,N_2985,N_1310);
nor U4071 (N_4071,N_2400,N_701);
and U4072 (N_4072,N_2879,N_1279);
nor U4073 (N_4073,N_2894,N_228);
nor U4074 (N_4074,N_566,N_2631);
nor U4075 (N_4075,N_2119,N_91);
nand U4076 (N_4076,N_1051,N_1417);
or U4077 (N_4077,N_564,N_1415);
nor U4078 (N_4078,N_2729,N_1710);
or U4079 (N_4079,N_2034,N_2850);
or U4080 (N_4080,N_1893,N_2730);
xnor U4081 (N_4081,N_2416,N_221);
nor U4082 (N_4082,N_1071,N_764);
and U4083 (N_4083,N_1184,N_456);
xor U4084 (N_4084,N_1384,N_1619);
and U4085 (N_4085,N_1148,N_820);
nand U4086 (N_4086,N_1153,N_699);
or U4087 (N_4087,N_2765,N_2935);
xor U4088 (N_4088,N_2485,N_2817);
nand U4089 (N_4089,N_2780,N_1411);
or U4090 (N_4090,N_189,N_2514);
nand U4091 (N_4091,N_694,N_453);
nor U4092 (N_4092,N_311,N_413);
or U4093 (N_4093,N_2395,N_961);
or U4094 (N_4094,N_452,N_1597);
and U4095 (N_4095,N_198,N_30);
and U4096 (N_4096,N_2073,N_2732);
nand U4097 (N_4097,N_763,N_19);
nand U4098 (N_4098,N_2186,N_2525);
nand U4099 (N_4099,N_1895,N_1608);
and U4100 (N_4100,N_1366,N_2466);
and U4101 (N_4101,N_45,N_466);
or U4102 (N_4102,N_745,N_2401);
nand U4103 (N_4103,N_677,N_2652);
and U4104 (N_4104,N_2058,N_2223);
nand U4105 (N_4105,N_2404,N_27);
nand U4106 (N_4106,N_1764,N_809);
and U4107 (N_4107,N_1352,N_1177);
or U4108 (N_4108,N_401,N_1325);
and U4109 (N_4109,N_10,N_351);
nor U4110 (N_4110,N_1791,N_1851);
and U4111 (N_4111,N_2054,N_1881);
or U4112 (N_4112,N_2283,N_1966);
or U4113 (N_4113,N_2861,N_2740);
nand U4114 (N_4114,N_1715,N_1581);
nand U4115 (N_4115,N_37,N_2870);
nor U4116 (N_4116,N_1020,N_2356);
or U4117 (N_4117,N_2845,N_1035);
nor U4118 (N_4118,N_1693,N_486);
or U4119 (N_4119,N_1412,N_2074);
and U4120 (N_4120,N_1674,N_1409);
and U4121 (N_4121,N_728,N_2246);
or U4122 (N_4122,N_884,N_2354);
and U4123 (N_4123,N_44,N_860);
nand U4124 (N_4124,N_158,N_2363);
or U4125 (N_4125,N_1259,N_2396);
or U4126 (N_4126,N_1625,N_1612);
and U4127 (N_4127,N_2386,N_2864);
and U4128 (N_4128,N_532,N_2133);
nand U4129 (N_4129,N_1171,N_2072);
or U4130 (N_4130,N_627,N_1822);
nand U4131 (N_4131,N_1958,N_435);
nand U4132 (N_4132,N_211,N_21);
or U4133 (N_4133,N_2467,N_2733);
and U4134 (N_4134,N_2349,N_2095);
and U4135 (N_4135,N_941,N_2966);
nor U4136 (N_4136,N_1953,N_1948);
or U4137 (N_4137,N_99,N_2842);
and U4138 (N_4138,N_2328,N_17);
nand U4139 (N_4139,N_2721,N_1082);
nor U4140 (N_4140,N_1589,N_220);
nand U4141 (N_4141,N_558,N_488);
nand U4142 (N_4142,N_2786,N_2131);
or U4143 (N_4143,N_1671,N_907);
and U4144 (N_4144,N_84,N_1908);
or U4145 (N_4145,N_493,N_1782);
nand U4146 (N_4146,N_2819,N_2244);
and U4147 (N_4147,N_318,N_1106);
and U4148 (N_4148,N_1913,N_2741);
nand U4149 (N_4149,N_71,N_229);
nand U4150 (N_4150,N_1419,N_1495);
nor U4151 (N_4151,N_1015,N_567);
or U4152 (N_4152,N_1289,N_1806);
nand U4153 (N_4153,N_2593,N_1981);
and U4154 (N_4154,N_2983,N_2598);
nand U4155 (N_4155,N_1472,N_110);
and U4156 (N_4156,N_2374,N_1134);
nand U4157 (N_4157,N_1481,N_319);
nand U4158 (N_4158,N_1570,N_1467);
and U4159 (N_4159,N_599,N_126);
or U4160 (N_4160,N_1010,N_1475);
nor U4161 (N_4161,N_1423,N_1624);
xnor U4162 (N_4162,N_2004,N_1661);
or U4163 (N_4163,N_1685,N_2417);
or U4164 (N_4164,N_985,N_1988);
nand U4165 (N_4165,N_2015,N_1334);
nand U4166 (N_4166,N_2151,N_1072);
or U4167 (N_4167,N_619,N_1452);
or U4168 (N_4168,N_1541,N_2956);
nor U4169 (N_4169,N_1399,N_2331);
and U4170 (N_4170,N_803,N_2952);
or U4171 (N_4171,N_271,N_2524);
nor U4172 (N_4172,N_2262,N_2213);
and U4173 (N_4173,N_835,N_883);
and U4174 (N_4174,N_1662,N_792);
and U4175 (N_4175,N_1132,N_2264);
nand U4176 (N_4176,N_557,N_1253);
nor U4177 (N_4177,N_138,N_1936);
nor U4178 (N_4178,N_2501,N_1508);
and U4179 (N_4179,N_1529,N_1925);
and U4180 (N_4180,N_1620,N_2362);
and U4181 (N_4181,N_1226,N_2098);
and U4182 (N_4182,N_1627,N_2012);
nor U4183 (N_4183,N_2921,N_861);
and U4184 (N_4184,N_905,N_670);
nor U4185 (N_4185,N_993,N_1779);
nand U4186 (N_4186,N_2277,N_242);
nor U4187 (N_4187,N_2088,N_344);
nor U4188 (N_4188,N_1504,N_153);
nand U4189 (N_4189,N_2481,N_122);
nand U4190 (N_4190,N_1237,N_2856);
nor U4191 (N_4191,N_2812,N_2608);
or U4192 (N_4192,N_2681,N_254);
nand U4193 (N_4193,N_1535,N_731);
or U4194 (N_4194,N_2382,N_2804);
xnor U4195 (N_4195,N_2480,N_2589);
or U4196 (N_4196,N_1677,N_314);
and U4197 (N_4197,N_1215,N_2946);
nand U4198 (N_4198,N_996,N_2961);
or U4199 (N_4199,N_209,N_1025);
and U4200 (N_4200,N_1456,N_185);
nor U4201 (N_4201,N_2083,N_263);
and U4202 (N_4202,N_1324,N_712);
and U4203 (N_4203,N_2571,N_1007);
nor U4204 (N_4204,N_6,N_2585);
nor U4205 (N_4205,N_2913,N_753);
nor U4206 (N_4206,N_770,N_2769);
or U4207 (N_4207,N_2517,N_648);
or U4208 (N_4208,N_2848,N_1558);
nor U4209 (N_4209,N_1427,N_2824);
nor U4210 (N_4210,N_425,N_2518);
or U4211 (N_4211,N_1482,N_2372);
nor U4212 (N_4212,N_394,N_2785);
nand U4213 (N_4213,N_871,N_1533);
or U4214 (N_4214,N_1302,N_2884);
and U4215 (N_4215,N_2207,N_1019);
or U4216 (N_4216,N_2537,N_338);
nand U4217 (N_4217,N_542,N_2509);
nor U4218 (N_4218,N_1031,N_858);
nand U4219 (N_4219,N_57,N_1554);
nor U4220 (N_4220,N_1138,N_2967);
and U4221 (N_4221,N_676,N_1679);
nor U4222 (N_4222,N_758,N_1800);
and U4223 (N_4223,N_897,N_1127);
nand U4224 (N_4224,N_1095,N_575);
nor U4225 (N_4225,N_932,N_1453);
nand U4226 (N_4226,N_1436,N_1037);
or U4227 (N_4227,N_423,N_265);
xnor U4228 (N_4228,N_2883,N_1723);
nor U4229 (N_4229,N_2575,N_1622);
nand U4230 (N_4230,N_739,N_1962);
and U4231 (N_4231,N_2260,N_1049);
or U4232 (N_4232,N_2837,N_2320);
nor U4233 (N_4233,N_938,N_1773);
nor U4234 (N_4234,N_23,N_1121);
and U4235 (N_4235,N_2182,N_2090);
or U4236 (N_4236,N_1928,N_2783);
xor U4237 (N_4237,N_1365,N_2858);
nor U4238 (N_4238,N_1854,N_1369);
and U4239 (N_4239,N_12,N_2834);
or U4240 (N_4240,N_1930,N_946);
or U4241 (N_4241,N_1096,N_480);
nor U4242 (N_4242,N_1449,N_1126);
nand U4243 (N_4243,N_2240,N_2327);
and U4244 (N_4244,N_2615,N_819);
nor U4245 (N_4245,N_1514,N_1591);
nand U4246 (N_4246,N_2278,N_2237);
xnor U4247 (N_4247,N_590,N_2658);
nand U4248 (N_4248,N_786,N_2406);
nor U4249 (N_4249,N_1167,N_359);
and U4250 (N_4250,N_2178,N_625);
nand U4251 (N_4251,N_2936,N_2476);
nor U4252 (N_4252,N_2376,N_892);
or U4253 (N_4253,N_2694,N_2851);
and U4254 (N_4254,N_1795,N_368);
or U4255 (N_4255,N_550,N_2144);
nand U4256 (N_4256,N_2273,N_5);
and U4257 (N_4257,N_696,N_1438);
nand U4258 (N_4258,N_826,N_2547);
and U4259 (N_4259,N_2748,N_1392);
and U4260 (N_4260,N_794,N_2446);
or U4261 (N_4261,N_2066,N_436);
or U4262 (N_4262,N_2271,N_387);
nor U4263 (N_4263,N_1265,N_1850);
and U4264 (N_4264,N_855,N_2337);
nand U4265 (N_4265,N_2560,N_1604);
and U4266 (N_4266,N_2999,N_161);
nand U4267 (N_4267,N_131,N_475);
nand U4268 (N_4268,N_1941,N_24);
nand U4269 (N_4269,N_836,N_909);
or U4270 (N_4270,N_730,N_173);
and U4271 (N_4271,N_1165,N_370);
nor U4272 (N_4272,N_726,N_2777);
nor U4273 (N_4273,N_2914,N_1350);
nor U4274 (N_4274,N_2465,N_767);
or U4275 (N_4275,N_1837,N_2759);
and U4276 (N_4276,N_371,N_1686);
or U4277 (N_4277,N_1042,N_210);
nor U4278 (N_4278,N_433,N_400);
nand U4279 (N_4279,N_2643,N_2887);
nor U4280 (N_4280,N_2181,N_1892);
nor U4281 (N_4281,N_2241,N_1331);
nor U4282 (N_4282,N_1073,N_164);
nand U4283 (N_4283,N_818,N_2579);
nor U4284 (N_4284,N_1145,N_1856);
or U4285 (N_4285,N_679,N_2316);
or U4286 (N_4286,N_2409,N_1952);
and U4287 (N_4287,N_449,N_2132);
nand U4288 (N_4288,N_1136,N_658);
nand U4289 (N_4289,N_2357,N_2159);
nor U4290 (N_4290,N_2431,N_2774);
or U4291 (N_4291,N_1146,N_2458);
or U4292 (N_4292,N_1880,N_2590);
nand U4293 (N_4293,N_85,N_111);
or U4294 (N_4294,N_15,N_2757);
nor U4295 (N_4295,N_1291,N_1805);
and U4296 (N_4296,N_1683,N_778);
or U4297 (N_4297,N_2970,N_2650);
nor U4298 (N_4298,N_1954,N_2989);
or U4299 (N_4299,N_1702,N_2569);
or U4300 (N_4300,N_944,N_2229);
and U4301 (N_4301,N_112,N_549);
nand U4302 (N_4302,N_1840,N_2954);
nand U4303 (N_4303,N_1924,N_2628);
nand U4304 (N_4304,N_2632,N_55);
or U4305 (N_4305,N_1586,N_707);
nand U4306 (N_4306,N_598,N_426);
nand U4307 (N_4307,N_2606,N_429);
and U4308 (N_4308,N_1899,N_641);
and U4309 (N_4309,N_2711,N_500);
and U4310 (N_4310,N_1052,N_1213);
nand U4311 (N_4311,N_2166,N_2214);
or U4312 (N_4312,N_868,N_190);
nand U4313 (N_4313,N_2570,N_8);
nor U4314 (N_4314,N_1027,N_2805);
or U4315 (N_4315,N_555,N_1647);
or U4316 (N_4316,N_384,N_2487);
nor U4317 (N_4317,N_1939,N_774);
nand U4318 (N_4318,N_2896,N_2112);
or U4319 (N_4319,N_174,N_915);
and U4320 (N_4320,N_2086,N_680);
nand U4321 (N_4321,N_2390,N_1326);
or U4322 (N_4322,N_2982,N_2475);
nand U4323 (N_4323,N_1379,N_326);
or U4324 (N_4324,N_1801,N_1568);
nand U4325 (N_4325,N_324,N_1987);
or U4326 (N_4326,N_1839,N_2116);
and U4327 (N_4327,N_2676,N_1721);
or U4328 (N_4328,N_1870,N_538);
nor U4329 (N_4329,N_1344,N_1224);
nand U4330 (N_4330,N_882,N_1656);
or U4331 (N_4331,N_2795,N_982);
or U4332 (N_4332,N_2915,N_412);
nand U4333 (N_4333,N_380,N_328);
nor U4334 (N_4334,N_261,N_1185);
nand U4335 (N_4335,N_865,N_2530);
nor U4336 (N_4336,N_983,N_1793);
and U4337 (N_4337,N_1810,N_1760);
nor U4338 (N_4338,N_981,N_1441);
or U4339 (N_4339,N_18,N_1263);
and U4340 (N_4340,N_1967,N_2788);
nor U4341 (N_4341,N_1713,N_391);
and U4342 (N_4342,N_9,N_1976);
nand U4343 (N_4343,N_2910,N_1157);
nand U4344 (N_4344,N_1414,N_2071);
or U4345 (N_4345,N_727,N_2930);
and U4346 (N_4346,N_1957,N_2613);
or U4347 (N_4347,N_1094,N_1315);
nand U4348 (N_4348,N_1045,N_2293);
nand U4349 (N_4349,N_2937,N_964);
nor U4350 (N_4350,N_801,N_1314);
and U4351 (N_4351,N_2800,N_2139);
and U4352 (N_4352,N_1963,N_1694);
nor U4353 (N_4353,N_1912,N_1729);
or U4354 (N_4354,N_662,N_2715);
or U4355 (N_4355,N_1918,N_2102);
or U4356 (N_4356,N_1281,N_1945);
nand U4357 (N_4357,N_1727,N_597);
nand U4358 (N_4358,N_1298,N_266);
xnor U4359 (N_4359,N_1243,N_1786);
nor U4360 (N_4360,N_948,N_2436);
nor U4361 (N_4361,N_1477,N_2414);
nand U4362 (N_4362,N_2420,N_427);
nand U4363 (N_4363,N_1748,N_2087);
nand U4364 (N_4364,N_1468,N_2190);
and U4365 (N_4365,N_2028,N_416);
and U4366 (N_4366,N_1942,N_2849);
nor U4367 (N_4367,N_397,N_975);
and U4368 (N_4368,N_1905,N_1838);
nand U4369 (N_4369,N_2533,N_1466);
nand U4370 (N_4370,N_1354,N_817);
nor U4371 (N_4371,N_2321,N_496);
or U4372 (N_4372,N_2231,N_1536);
nand U4373 (N_4373,N_880,N_2934);
nand U4374 (N_4374,N_1845,N_2198);
or U4375 (N_4375,N_539,N_1113);
or U4376 (N_4376,N_2469,N_672);
or U4377 (N_4377,N_448,N_187);
and U4378 (N_4378,N_546,N_2474);
or U4379 (N_4379,N_1222,N_1499);
or U4380 (N_4380,N_1902,N_1244);
nor U4381 (N_4381,N_1406,N_1085);
nor U4382 (N_4382,N_2508,N_2564);
nor U4383 (N_4383,N_807,N_1883);
and U4384 (N_4384,N_1050,N_2793);
or U4385 (N_4385,N_2662,N_2962);
nand U4386 (N_4386,N_708,N_1563);
nand U4387 (N_4387,N_1230,N_2359);
nand U4388 (N_4388,N_1553,N_2924);
nand U4389 (N_4389,N_183,N_2398);
and U4390 (N_4390,N_236,N_965);
and U4391 (N_4391,N_2000,N_895);
or U4392 (N_4392,N_2165,N_2992);
xor U4393 (N_4393,N_358,N_2047);
and U4394 (N_4394,N_1164,N_374);
nand U4395 (N_4395,N_1669,N_127);
or U4396 (N_4396,N_478,N_813);
and U4397 (N_4397,N_544,N_2342);
nand U4398 (N_4398,N_678,N_1544);
and U4399 (N_4399,N_2050,N_2080);
nor U4400 (N_4400,N_990,N_782);
and U4401 (N_4401,N_2215,N_754);
nand U4402 (N_4402,N_1561,N_2897);
and U4403 (N_4403,N_777,N_1574);
and U4404 (N_4404,N_2801,N_2955);
and U4405 (N_4405,N_618,N_629);
nand U4406 (N_4406,N_1404,N_2971);
or U4407 (N_4407,N_666,N_616);
or U4408 (N_4408,N_1758,N_537);
or U4409 (N_4409,N_1022,N_304);
or U4410 (N_4410,N_2500,N_1099);
nor U4411 (N_4411,N_1600,N_925);
or U4412 (N_4412,N_2581,N_2353);
nand U4413 (N_4413,N_2911,N_551);
nor U4414 (N_4414,N_78,N_1752);
nor U4415 (N_4415,N_911,N_1212);
nand U4416 (N_4416,N_1061,N_1634);
nand U4417 (N_4417,N_776,N_377);
or U4418 (N_4418,N_1195,N_1091);
or U4419 (N_4419,N_445,N_179);
or U4420 (N_4420,N_628,N_2455);
or U4421 (N_4421,N_1209,N_970);
or U4422 (N_4422,N_2727,N_2016);
or U4423 (N_4423,N_799,N_2692);
nor U4424 (N_4424,N_1569,N_43);
nor U4425 (N_4425,N_2194,N_405);
or U4426 (N_4426,N_2925,N_1474);
and U4427 (N_4427,N_1731,N_2880);
nand U4428 (N_4428,N_1498,N_1150);
nand U4429 (N_4429,N_2690,N_1316);
or U4430 (N_4430,N_2835,N_1626);
or U4431 (N_4431,N_1528,N_2493);
nor U4432 (N_4432,N_2118,N_2633);
nand U4433 (N_4433,N_1652,N_804);
and U4434 (N_4434,N_2657,N_2038);
nand U4435 (N_4435,N_2638,N_2820);
nand U4436 (N_4436,N_451,N_170);
and U4437 (N_4437,N_2885,N_2677);
nand U4438 (N_4438,N_1965,N_1776);
or U4439 (N_4439,N_2270,N_2387);
and U4440 (N_4440,N_1277,N_2531);
nand U4441 (N_4441,N_479,N_2685);
nand U4442 (N_4442,N_282,N_1914);
or U4443 (N_4443,N_1361,N_2384);
or U4444 (N_4444,N_177,N_1659);
or U4445 (N_4445,N_2724,N_2767);
nor U4446 (N_4446,N_1617,N_2175);
and U4447 (N_4447,N_2901,N_1367);
and U4448 (N_4448,N_1434,N_1197);
nand U4449 (N_4449,N_1663,N_1692);
nand U4450 (N_4450,N_2720,N_1821);
nor U4451 (N_4451,N_536,N_959);
and U4452 (N_4452,N_1780,N_1444);
and U4453 (N_4453,N_1374,N_989);
or U4454 (N_4454,N_352,N_1975);
nor U4455 (N_4455,N_653,N_340);
nor U4456 (N_4456,N_1439,N_1774);
nor U4457 (N_4457,N_1889,N_192);
or U4458 (N_4458,N_2239,N_2749);
and U4459 (N_4459,N_1428,N_843);
nor U4460 (N_4460,N_2577,N_1074);
nand U4461 (N_4461,N_2421,N_1759);
nor U4462 (N_4462,N_2360,N_1004);
and U4463 (N_4463,N_1673,N_1658);
xnor U4464 (N_4464,N_1278,N_1859);
nor U4465 (N_4465,N_1628,N_232);
nand U4466 (N_4466,N_2128,N_2341);
nor U4467 (N_4467,N_2742,N_2919);
nand U4468 (N_4468,N_2596,N_545);
nand U4469 (N_4469,N_117,N_1413);
nand U4470 (N_4470,N_2389,N_2340);
nor U4471 (N_4471,N_1286,N_218);
and U4472 (N_4472,N_2423,N_2408);
and U4473 (N_4473,N_1532,N_2013);
nor U4474 (N_4474,N_2976,N_2292);
nor U4475 (N_4475,N_773,N_934);
xnor U4476 (N_4476,N_1993,N_2482);
and U4477 (N_4477,N_854,N_2422);
and U4478 (N_4478,N_851,N_1901);
or U4479 (N_4479,N_929,N_341);
and U4480 (N_4480,N_2323,N_472);
nor U4481 (N_4481,N_1333,N_891);
nand U4482 (N_4482,N_13,N_16);
or U4483 (N_4483,N_1735,N_2195);
and U4484 (N_4484,N_2326,N_1781);
nor U4485 (N_4485,N_1080,N_2082);
nor U4486 (N_4486,N_2472,N_2857);
and U4487 (N_4487,N_2863,N_270);
nor U4488 (N_4488,N_2719,N_2403);
nand U4489 (N_4489,N_1605,N_1205);
and U4490 (N_4490,N_1578,N_2697);
and U4491 (N_4491,N_42,N_1283);
nor U4492 (N_4492,N_2763,N_1590);
or U4493 (N_4493,N_1123,N_82);
nor U4494 (N_4494,N_581,N_2236);
nor U4495 (N_4495,N_2120,N_645);
or U4496 (N_4496,N_430,N_2289);
nand U4497 (N_4497,N_443,N_2282);
and U4498 (N_4498,N_2242,N_1260);
or U4499 (N_4499,N_2296,N_196);
or U4500 (N_4500,N_223,N_1962);
or U4501 (N_4501,N_1362,N_2381);
and U4502 (N_4502,N_2193,N_2540);
nand U4503 (N_4503,N_2263,N_993);
and U4504 (N_4504,N_1123,N_2572);
nor U4505 (N_4505,N_1486,N_2708);
nand U4506 (N_4506,N_1185,N_1422);
or U4507 (N_4507,N_2764,N_2744);
and U4508 (N_4508,N_2567,N_601);
nand U4509 (N_4509,N_751,N_436);
nor U4510 (N_4510,N_1132,N_81);
or U4511 (N_4511,N_450,N_1672);
nand U4512 (N_4512,N_2973,N_1030);
nand U4513 (N_4513,N_2062,N_1837);
nand U4514 (N_4514,N_1961,N_1507);
nand U4515 (N_4515,N_255,N_687);
and U4516 (N_4516,N_2157,N_1186);
nor U4517 (N_4517,N_681,N_2174);
and U4518 (N_4518,N_863,N_2316);
and U4519 (N_4519,N_413,N_864);
nand U4520 (N_4520,N_2861,N_1133);
and U4521 (N_4521,N_1689,N_623);
nor U4522 (N_4522,N_2820,N_87);
nand U4523 (N_4523,N_1766,N_124);
xor U4524 (N_4524,N_1520,N_12);
and U4525 (N_4525,N_1893,N_2528);
and U4526 (N_4526,N_165,N_1101);
and U4527 (N_4527,N_2874,N_2809);
and U4528 (N_4528,N_2244,N_829);
or U4529 (N_4529,N_1929,N_2369);
or U4530 (N_4530,N_8,N_423);
nand U4531 (N_4531,N_2772,N_2373);
nand U4532 (N_4532,N_839,N_2539);
nor U4533 (N_4533,N_2965,N_2859);
or U4534 (N_4534,N_733,N_1228);
or U4535 (N_4535,N_1474,N_2196);
and U4536 (N_4536,N_1739,N_1383);
or U4537 (N_4537,N_701,N_776);
and U4538 (N_4538,N_1906,N_74);
nor U4539 (N_4539,N_2501,N_2563);
and U4540 (N_4540,N_150,N_2100);
nand U4541 (N_4541,N_212,N_385);
and U4542 (N_4542,N_1422,N_2635);
or U4543 (N_4543,N_1588,N_1565);
or U4544 (N_4544,N_1045,N_1707);
and U4545 (N_4545,N_1668,N_2220);
nand U4546 (N_4546,N_2900,N_1991);
and U4547 (N_4547,N_2107,N_1872);
and U4548 (N_4548,N_547,N_1748);
and U4549 (N_4549,N_1931,N_2032);
and U4550 (N_4550,N_2747,N_1961);
or U4551 (N_4551,N_712,N_1090);
and U4552 (N_4552,N_1758,N_40);
and U4553 (N_4553,N_1548,N_574);
and U4554 (N_4554,N_1275,N_1221);
nor U4555 (N_4555,N_124,N_1123);
and U4556 (N_4556,N_1769,N_1331);
nand U4557 (N_4557,N_265,N_2217);
nor U4558 (N_4558,N_447,N_58);
nor U4559 (N_4559,N_2367,N_37);
or U4560 (N_4560,N_2079,N_41);
nor U4561 (N_4561,N_2625,N_275);
nor U4562 (N_4562,N_2996,N_2577);
nor U4563 (N_4563,N_156,N_1815);
or U4564 (N_4564,N_1741,N_774);
or U4565 (N_4565,N_2098,N_1435);
and U4566 (N_4566,N_2915,N_301);
nand U4567 (N_4567,N_1571,N_2632);
and U4568 (N_4568,N_2701,N_1683);
or U4569 (N_4569,N_2294,N_703);
nor U4570 (N_4570,N_2381,N_930);
and U4571 (N_4571,N_1677,N_671);
or U4572 (N_4572,N_1501,N_1406);
nor U4573 (N_4573,N_1212,N_1059);
and U4574 (N_4574,N_2998,N_1267);
nand U4575 (N_4575,N_2834,N_2382);
or U4576 (N_4576,N_402,N_238);
or U4577 (N_4577,N_1425,N_1603);
nand U4578 (N_4578,N_899,N_1053);
and U4579 (N_4579,N_36,N_2361);
nor U4580 (N_4580,N_1039,N_712);
or U4581 (N_4581,N_2377,N_1879);
and U4582 (N_4582,N_1985,N_2266);
and U4583 (N_4583,N_1262,N_1038);
or U4584 (N_4584,N_137,N_2675);
and U4585 (N_4585,N_518,N_1649);
and U4586 (N_4586,N_1794,N_1480);
and U4587 (N_4587,N_2812,N_1028);
xnor U4588 (N_4588,N_2647,N_2547);
and U4589 (N_4589,N_586,N_1309);
nand U4590 (N_4590,N_1871,N_424);
nand U4591 (N_4591,N_1597,N_2601);
nand U4592 (N_4592,N_299,N_1502);
nor U4593 (N_4593,N_1772,N_2092);
and U4594 (N_4594,N_43,N_360);
nand U4595 (N_4595,N_798,N_953);
nand U4596 (N_4596,N_1534,N_2829);
nand U4597 (N_4597,N_1046,N_1379);
nand U4598 (N_4598,N_2646,N_1793);
nand U4599 (N_4599,N_2427,N_287);
and U4600 (N_4600,N_2335,N_2924);
or U4601 (N_4601,N_2644,N_1156);
nor U4602 (N_4602,N_402,N_1986);
or U4603 (N_4603,N_926,N_52);
nand U4604 (N_4604,N_378,N_2067);
and U4605 (N_4605,N_666,N_1889);
nand U4606 (N_4606,N_208,N_1107);
or U4607 (N_4607,N_324,N_983);
and U4608 (N_4608,N_1320,N_1968);
or U4609 (N_4609,N_559,N_2497);
nand U4610 (N_4610,N_47,N_2924);
and U4611 (N_4611,N_2532,N_283);
nand U4612 (N_4612,N_817,N_1650);
or U4613 (N_4613,N_2952,N_443);
and U4614 (N_4614,N_665,N_2141);
nor U4615 (N_4615,N_1683,N_2360);
or U4616 (N_4616,N_380,N_1541);
or U4617 (N_4617,N_699,N_2239);
nand U4618 (N_4618,N_1164,N_2184);
or U4619 (N_4619,N_1963,N_312);
nand U4620 (N_4620,N_1884,N_2103);
and U4621 (N_4621,N_385,N_566);
and U4622 (N_4622,N_2905,N_2302);
nand U4623 (N_4623,N_273,N_976);
and U4624 (N_4624,N_1271,N_2375);
nor U4625 (N_4625,N_698,N_1063);
nand U4626 (N_4626,N_1174,N_1665);
or U4627 (N_4627,N_498,N_2034);
or U4628 (N_4628,N_1769,N_2353);
nand U4629 (N_4629,N_1246,N_1616);
nand U4630 (N_4630,N_439,N_1991);
or U4631 (N_4631,N_1476,N_1008);
nor U4632 (N_4632,N_1533,N_317);
or U4633 (N_4633,N_554,N_387);
and U4634 (N_4634,N_661,N_1006);
or U4635 (N_4635,N_348,N_2480);
or U4636 (N_4636,N_1610,N_1514);
or U4637 (N_4637,N_2199,N_2459);
or U4638 (N_4638,N_1738,N_1518);
or U4639 (N_4639,N_2004,N_307);
nor U4640 (N_4640,N_1256,N_2450);
nand U4641 (N_4641,N_14,N_1488);
nand U4642 (N_4642,N_2164,N_1620);
or U4643 (N_4643,N_1218,N_1930);
or U4644 (N_4644,N_167,N_2690);
and U4645 (N_4645,N_33,N_1020);
and U4646 (N_4646,N_2212,N_2979);
or U4647 (N_4647,N_840,N_1070);
or U4648 (N_4648,N_891,N_1115);
or U4649 (N_4649,N_2687,N_2994);
nor U4650 (N_4650,N_303,N_2661);
nand U4651 (N_4651,N_2339,N_90);
or U4652 (N_4652,N_2071,N_59);
and U4653 (N_4653,N_2098,N_1637);
or U4654 (N_4654,N_2349,N_908);
or U4655 (N_4655,N_1589,N_1141);
and U4656 (N_4656,N_1923,N_470);
or U4657 (N_4657,N_1780,N_175);
nand U4658 (N_4658,N_2259,N_2554);
or U4659 (N_4659,N_1483,N_2952);
or U4660 (N_4660,N_772,N_508);
nor U4661 (N_4661,N_545,N_1298);
nand U4662 (N_4662,N_2554,N_2753);
or U4663 (N_4663,N_1402,N_1346);
nand U4664 (N_4664,N_591,N_1268);
and U4665 (N_4665,N_2568,N_1592);
and U4666 (N_4666,N_2502,N_569);
and U4667 (N_4667,N_1851,N_2454);
or U4668 (N_4668,N_2378,N_552);
nand U4669 (N_4669,N_692,N_2179);
nand U4670 (N_4670,N_266,N_2433);
and U4671 (N_4671,N_2175,N_1598);
and U4672 (N_4672,N_655,N_940);
xnor U4673 (N_4673,N_2289,N_2378);
nor U4674 (N_4674,N_2412,N_2903);
nand U4675 (N_4675,N_2198,N_2440);
nand U4676 (N_4676,N_606,N_1924);
nor U4677 (N_4677,N_2254,N_1669);
nor U4678 (N_4678,N_2510,N_1852);
or U4679 (N_4679,N_1394,N_396);
nand U4680 (N_4680,N_274,N_2890);
and U4681 (N_4681,N_2495,N_2);
nor U4682 (N_4682,N_1228,N_1409);
and U4683 (N_4683,N_1794,N_2404);
nand U4684 (N_4684,N_2062,N_569);
nand U4685 (N_4685,N_2223,N_2247);
or U4686 (N_4686,N_2428,N_1068);
and U4687 (N_4687,N_509,N_1304);
nand U4688 (N_4688,N_1119,N_1537);
nor U4689 (N_4689,N_243,N_2812);
nand U4690 (N_4690,N_709,N_1411);
nand U4691 (N_4691,N_386,N_2116);
nand U4692 (N_4692,N_698,N_281);
and U4693 (N_4693,N_1619,N_1961);
or U4694 (N_4694,N_1779,N_2222);
nor U4695 (N_4695,N_2037,N_2671);
or U4696 (N_4696,N_2876,N_1721);
and U4697 (N_4697,N_1240,N_2588);
and U4698 (N_4698,N_416,N_2937);
nand U4699 (N_4699,N_1734,N_1026);
and U4700 (N_4700,N_2621,N_2643);
or U4701 (N_4701,N_2265,N_1435);
nand U4702 (N_4702,N_1203,N_1460);
or U4703 (N_4703,N_2324,N_914);
or U4704 (N_4704,N_808,N_1431);
nand U4705 (N_4705,N_2113,N_873);
nor U4706 (N_4706,N_2115,N_1461);
or U4707 (N_4707,N_1447,N_1796);
and U4708 (N_4708,N_1627,N_2296);
and U4709 (N_4709,N_1106,N_2524);
or U4710 (N_4710,N_808,N_2713);
nand U4711 (N_4711,N_2827,N_1304);
or U4712 (N_4712,N_1006,N_1086);
or U4713 (N_4713,N_712,N_151);
nor U4714 (N_4714,N_1064,N_1351);
nand U4715 (N_4715,N_740,N_1751);
or U4716 (N_4716,N_1442,N_653);
and U4717 (N_4717,N_1323,N_1538);
or U4718 (N_4718,N_349,N_1384);
nor U4719 (N_4719,N_1208,N_759);
or U4720 (N_4720,N_2564,N_2324);
or U4721 (N_4721,N_373,N_1951);
nand U4722 (N_4722,N_2775,N_893);
nand U4723 (N_4723,N_228,N_2529);
nand U4724 (N_4724,N_2847,N_1641);
or U4725 (N_4725,N_2520,N_2825);
and U4726 (N_4726,N_1311,N_1790);
nand U4727 (N_4727,N_60,N_659);
or U4728 (N_4728,N_1765,N_2052);
or U4729 (N_4729,N_1196,N_1286);
and U4730 (N_4730,N_2548,N_2499);
nand U4731 (N_4731,N_2228,N_2199);
nand U4732 (N_4732,N_613,N_2927);
nor U4733 (N_4733,N_2203,N_329);
and U4734 (N_4734,N_2758,N_2941);
xor U4735 (N_4735,N_2493,N_2095);
nand U4736 (N_4736,N_451,N_929);
xor U4737 (N_4737,N_2548,N_245);
and U4738 (N_4738,N_2204,N_2987);
nand U4739 (N_4739,N_2982,N_1034);
or U4740 (N_4740,N_82,N_186);
or U4741 (N_4741,N_1565,N_1638);
or U4742 (N_4742,N_1990,N_2138);
or U4743 (N_4743,N_2748,N_538);
and U4744 (N_4744,N_1250,N_1192);
and U4745 (N_4745,N_2506,N_565);
nor U4746 (N_4746,N_289,N_2275);
xnor U4747 (N_4747,N_1629,N_44);
and U4748 (N_4748,N_994,N_885);
and U4749 (N_4749,N_880,N_1354);
or U4750 (N_4750,N_1073,N_2415);
or U4751 (N_4751,N_2384,N_1899);
nand U4752 (N_4752,N_357,N_2327);
and U4753 (N_4753,N_873,N_2724);
or U4754 (N_4754,N_2931,N_669);
or U4755 (N_4755,N_1974,N_36);
nor U4756 (N_4756,N_2694,N_655);
and U4757 (N_4757,N_2023,N_366);
and U4758 (N_4758,N_646,N_2560);
and U4759 (N_4759,N_845,N_527);
nor U4760 (N_4760,N_765,N_171);
or U4761 (N_4761,N_1869,N_908);
or U4762 (N_4762,N_669,N_2113);
and U4763 (N_4763,N_126,N_2075);
nand U4764 (N_4764,N_731,N_2639);
or U4765 (N_4765,N_2574,N_248);
or U4766 (N_4766,N_310,N_1515);
and U4767 (N_4767,N_762,N_1694);
or U4768 (N_4768,N_1199,N_1742);
nor U4769 (N_4769,N_2030,N_2691);
and U4770 (N_4770,N_1092,N_282);
and U4771 (N_4771,N_2158,N_2370);
and U4772 (N_4772,N_1996,N_616);
nand U4773 (N_4773,N_2213,N_2370);
nor U4774 (N_4774,N_2850,N_429);
nor U4775 (N_4775,N_2418,N_537);
nor U4776 (N_4776,N_2855,N_2233);
or U4777 (N_4777,N_1918,N_988);
nand U4778 (N_4778,N_1967,N_1347);
or U4779 (N_4779,N_2130,N_2828);
nor U4780 (N_4780,N_1132,N_708);
and U4781 (N_4781,N_1534,N_1500);
or U4782 (N_4782,N_983,N_128);
nand U4783 (N_4783,N_992,N_2365);
and U4784 (N_4784,N_2938,N_2381);
nand U4785 (N_4785,N_2093,N_1685);
or U4786 (N_4786,N_2032,N_1771);
nor U4787 (N_4787,N_1901,N_2709);
nand U4788 (N_4788,N_1018,N_1015);
nand U4789 (N_4789,N_1367,N_2583);
nand U4790 (N_4790,N_1003,N_1818);
and U4791 (N_4791,N_1423,N_1225);
and U4792 (N_4792,N_1671,N_2129);
nor U4793 (N_4793,N_2528,N_335);
or U4794 (N_4794,N_345,N_2578);
or U4795 (N_4795,N_900,N_363);
nor U4796 (N_4796,N_1490,N_2146);
nand U4797 (N_4797,N_150,N_2521);
nor U4798 (N_4798,N_191,N_2084);
nor U4799 (N_4799,N_2842,N_2396);
and U4800 (N_4800,N_1067,N_1179);
nand U4801 (N_4801,N_744,N_969);
or U4802 (N_4802,N_796,N_2584);
and U4803 (N_4803,N_2125,N_35);
nor U4804 (N_4804,N_2428,N_2620);
and U4805 (N_4805,N_220,N_565);
and U4806 (N_4806,N_2223,N_2125);
and U4807 (N_4807,N_1241,N_2939);
nor U4808 (N_4808,N_468,N_344);
nand U4809 (N_4809,N_2698,N_502);
nor U4810 (N_4810,N_2899,N_1101);
nand U4811 (N_4811,N_74,N_2299);
and U4812 (N_4812,N_1637,N_1765);
nor U4813 (N_4813,N_628,N_2500);
nor U4814 (N_4814,N_2421,N_1453);
nor U4815 (N_4815,N_2488,N_640);
nand U4816 (N_4816,N_637,N_772);
or U4817 (N_4817,N_1718,N_2242);
and U4818 (N_4818,N_1448,N_1973);
nand U4819 (N_4819,N_1249,N_1236);
and U4820 (N_4820,N_1131,N_2109);
nor U4821 (N_4821,N_1448,N_8);
or U4822 (N_4822,N_501,N_291);
nor U4823 (N_4823,N_754,N_1519);
or U4824 (N_4824,N_2361,N_623);
or U4825 (N_4825,N_868,N_2282);
or U4826 (N_4826,N_441,N_1295);
nand U4827 (N_4827,N_2621,N_935);
and U4828 (N_4828,N_772,N_517);
nand U4829 (N_4829,N_2725,N_1091);
or U4830 (N_4830,N_36,N_1346);
nand U4831 (N_4831,N_392,N_2362);
and U4832 (N_4832,N_2791,N_2023);
or U4833 (N_4833,N_312,N_632);
nor U4834 (N_4834,N_600,N_145);
nand U4835 (N_4835,N_1195,N_165);
and U4836 (N_4836,N_1060,N_156);
or U4837 (N_4837,N_2011,N_1323);
nand U4838 (N_4838,N_2751,N_2041);
or U4839 (N_4839,N_2010,N_141);
or U4840 (N_4840,N_1239,N_2243);
nor U4841 (N_4841,N_600,N_224);
nand U4842 (N_4842,N_1663,N_778);
or U4843 (N_4843,N_1234,N_762);
nor U4844 (N_4844,N_437,N_1414);
nor U4845 (N_4845,N_1087,N_65);
or U4846 (N_4846,N_1826,N_1715);
or U4847 (N_4847,N_518,N_2217);
nor U4848 (N_4848,N_1304,N_1013);
nor U4849 (N_4849,N_2049,N_2729);
nand U4850 (N_4850,N_1891,N_2981);
nand U4851 (N_4851,N_1296,N_2637);
nand U4852 (N_4852,N_134,N_479);
or U4853 (N_4853,N_521,N_2820);
or U4854 (N_4854,N_262,N_1189);
and U4855 (N_4855,N_412,N_1774);
nor U4856 (N_4856,N_2522,N_2121);
or U4857 (N_4857,N_1697,N_1813);
and U4858 (N_4858,N_2065,N_2848);
nor U4859 (N_4859,N_822,N_2152);
and U4860 (N_4860,N_2147,N_899);
and U4861 (N_4861,N_1323,N_1203);
nor U4862 (N_4862,N_33,N_2059);
nand U4863 (N_4863,N_478,N_2831);
nand U4864 (N_4864,N_1242,N_2124);
nand U4865 (N_4865,N_846,N_1868);
or U4866 (N_4866,N_547,N_112);
nor U4867 (N_4867,N_2944,N_1179);
nand U4868 (N_4868,N_2321,N_2860);
and U4869 (N_4869,N_1246,N_714);
and U4870 (N_4870,N_1931,N_2612);
and U4871 (N_4871,N_650,N_1444);
nand U4872 (N_4872,N_2915,N_1907);
and U4873 (N_4873,N_2037,N_1470);
or U4874 (N_4874,N_1117,N_2098);
or U4875 (N_4875,N_2373,N_1905);
nand U4876 (N_4876,N_2218,N_1776);
and U4877 (N_4877,N_242,N_1425);
nor U4878 (N_4878,N_2109,N_2233);
nor U4879 (N_4879,N_2429,N_2209);
nand U4880 (N_4880,N_828,N_1778);
nand U4881 (N_4881,N_661,N_2794);
nand U4882 (N_4882,N_2529,N_2651);
or U4883 (N_4883,N_1462,N_1460);
nor U4884 (N_4884,N_2801,N_1697);
nor U4885 (N_4885,N_2786,N_2645);
nand U4886 (N_4886,N_986,N_436);
or U4887 (N_4887,N_2807,N_28);
and U4888 (N_4888,N_1873,N_198);
nand U4889 (N_4889,N_2834,N_1627);
nand U4890 (N_4890,N_1955,N_1205);
nand U4891 (N_4891,N_1102,N_2940);
nand U4892 (N_4892,N_2657,N_2943);
nor U4893 (N_4893,N_1694,N_2809);
and U4894 (N_4894,N_2628,N_1360);
nor U4895 (N_4895,N_1975,N_2781);
nor U4896 (N_4896,N_1351,N_2414);
and U4897 (N_4897,N_2801,N_964);
nand U4898 (N_4898,N_388,N_1257);
or U4899 (N_4899,N_1037,N_29);
or U4900 (N_4900,N_912,N_2360);
nand U4901 (N_4901,N_157,N_1587);
and U4902 (N_4902,N_1127,N_206);
nor U4903 (N_4903,N_2028,N_1258);
nand U4904 (N_4904,N_1811,N_2878);
nor U4905 (N_4905,N_427,N_1274);
nor U4906 (N_4906,N_1146,N_2787);
or U4907 (N_4907,N_1089,N_1834);
and U4908 (N_4908,N_2596,N_219);
and U4909 (N_4909,N_1241,N_1074);
nor U4910 (N_4910,N_1904,N_2826);
nor U4911 (N_4911,N_2157,N_672);
and U4912 (N_4912,N_2137,N_1836);
nand U4913 (N_4913,N_1592,N_2761);
or U4914 (N_4914,N_2302,N_2539);
nand U4915 (N_4915,N_2791,N_1238);
xor U4916 (N_4916,N_1271,N_78);
or U4917 (N_4917,N_930,N_2774);
or U4918 (N_4918,N_353,N_2636);
and U4919 (N_4919,N_202,N_1249);
or U4920 (N_4920,N_783,N_1266);
nand U4921 (N_4921,N_2662,N_700);
and U4922 (N_4922,N_1620,N_1006);
nor U4923 (N_4923,N_2025,N_2554);
and U4924 (N_4924,N_2983,N_114);
and U4925 (N_4925,N_957,N_1977);
and U4926 (N_4926,N_872,N_1199);
or U4927 (N_4927,N_2777,N_2395);
and U4928 (N_4928,N_2216,N_2647);
and U4929 (N_4929,N_2354,N_1143);
and U4930 (N_4930,N_1803,N_2149);
or U4931 (N_4931,N_650,N_1719);
and U4932 (N_4932,N_320,N_2746);
and U4933 (N_4933,N_2602,N_1988);
nor U4934 (N_4934,N_1026,N_1161);
or U4935 (N_4935,N_1439,N_417);
or U4936 (N_4936,N_324,N_56);
or U4937 (N_4937,N_1855,N_1094);
and U4938 (N_4938,N_2445,N_240);
nor U4939 (N_4939,N_2015,N_1432);
nand U4940 (N_4940,N_2155,N_2318);
nand U4941 (N_4941,N_300,N_682);
or U4942 (N_4942,N_1920,N_1517);
and U4943 (N_4943,N_1166,N_565);
or U4944 (N_4944,N_1891,N_1008);
or U4945 (N_4945,N_2018,N_971);
or U4946 (N_4946,N_1332,N_293);
nand U4947 (N_4947,N_1173,N_1775);
nand U4948 (N_4948,N_72,N_2420);
or U4949 (N_4949,N_1276,N_1879);
nor U4950 (N_4950,N_314,N_1026);
or U4951 (N_4951,N_483,N_1238);
or U4952 (N_4952,N_1069,N_1186);
nor U4953 (N_4953,N_847,N_2462);
or U4954 (N_4954,N_517,N_2459);
and U4955 (N_4955,N_1909,N_1384);
nor U4956 (N_4956,N_375,N_514);
or U4957 (N_4957,N_1386,N_1606);
nand U4958 (N_4958,N_1239,N_473);
and U4959 (N_4959,N_788,N_1438);
and U4960 (N_4960,N_2120,N_1050);
nor U4961 (N_4961,N_2478,N_1614);
or U4962 (N_4962,N_1976,N_989);
and U4963 (N_4963,N_2893,N_782);
and U4964 (N_4964,N_1314,N_1739);
or U4965 (N_4965,N_104,N_2310);
nand U4966 (N_4966,N_712,N_2502);
and U4967 (N_4967,N_2114,N_2385);
nor U4968 (N_4968,N_2347,N_1614);
and U4969 (N_4969,N_1627,N_525);
or U4970 (N_4970,N_1796,N_2352);
nor U4971 (N_4971,N_1084,N_2749);
nand U4972 (N_4972,N_878,N_1880);
or U4973 (N_4973,N_2936,N_2386);
and U4974 (N_4974,N_2051,N_2973);
and U4975 (N_4975,N_2853,N_1393);
nand U4976 (N_4976,N_150,N_1610);
nor U4977 (N_4977,N_2075,N_1327);
and U4978 (N_4978,N_2758,N_2012);
and U4979 (N_4979,N_45,N_1873);
and U4980 (N_4980,N_8,N_2907);
nand U4981 (N_4981,N_1853,N_216);
and U4982 (N_4982,N_2080,N_735);
or U4983 (N_4983,N_1141,N_2507);
nor U4984 (N_4984,N_368,N_585);
or U4985 (N_4985,N_957,N_2121);
or U4986 (N_4986,N_2454,N_2376);
and U4987 (N_4987,N_1670,N_2534);
and U4988 (N_4988,N_439,N_164);
and U4989 (N_4989,N_2845,N_2635);
or U4990 (N_4990,N_1997,N_77);
and U4991 (N_4991,N_2110,N_2271);
or U4992 (N_4992,N_2450,N_1013);
nor U4993 (N_4993,N_1764,N_35);
nand U4994 (N_4994,N_1158,N_840);
or U4995 (N_4995,N_804,N_2731);
and U4996 (N_4996,N_581,N_1011);
and U4997 (N_4997,N_2458,N_2761);
and U4998 (N_4998,N_120,N_1385);
and U4999 (N_4999,N_1724,N_1237);
or U5000 (N_5000,N_2036,N_1527);
nor U5001 (N_5001,N_1531,N_751);
and U5002 (N_5002,N_687,N_2616);
or U5003 (N_5003,N_6,N_1017);
or U5004 (N_5004,N_2580,N_2175);
nand U5005 (N_5005,N_1048,N_1436);
or U5006 (N_5006,N_2462,N_2263);
or U5007 (N_5007,N_2518,N_1530);
or U5008 (N_5008,N_1335,N_2286);
nand U5009 (N_5009,N_714,N_2140);
nor U5010 (N_5010,N_2036,N_1351);
nand U5011 (N_5011,N_314,N_2119);
nor U5012 (N_5012,N_769,N_2817);
nand U5013 (N_5013,N_2482,N_2988);
and U5014 (N_5014,N_1134,N_2274);
nand U5015 (N_5015,N_534,N_2469);
nor U5016 (N_5016,N_838,N_969);
nand U5017 (N_5017,N_2799,N_1568);
and U5018 (N_5018,N_1937,N_949);
or U5019 (N_5019,N_1772,N_256);
or U5020 (N_5020,N_1578,N_867);
nand U5021 (N_5021,N_2603,N_2554);
and U5022 (N_5022,N_288,N_29);
and U5023 (N_5023,N_2234,N_1521);
and U5024 (N_5024,N_1324,N_2265);
and U5025 (N_5025,N_1836,N_2728);
and U5026 (N_5026,N_1484,N_1191);
or U5027 (N_5027,N_2104,N_2986);
nand U5028 (N_5028,N_1445,N_1529);
nand U5029 (N_5029,N_987,N_1356);
nand U5030 (N_5030,N_187,N_2168);
nand U5031 (N_5031,N_1829,N_2776);
nand U5032 (N_5032,N_2460,N_570);
or U5033 (N_5033,N_1846,N_1169);
or U5034 (N_5034,N_681,N_556);
nand U5035 (N_5035,N_207,N_1551);
or U5036 (N_5036,N_1516,N_774);
nand U5037 (N_5037,N_2301,N_1793);
xnor U5038 (N_5038,N_2033,N_604);
and U5039 (N_5039,N_667,N_1360);
or U5040 (N_5040,N_601,N_155);
nor U5041 (N_5041,N_775,N_720);
nor U5042 (N_5042,N_1522,N_543);
and U5043 (N_5043,N_1189,N_1310);
or U5044 (N_5044,N_2291,N_1394);
nand U5045 (N_5045,N_729,N_935);
or U5046 (N_5046,N_1984,N_979);
nor U5047 (N_5047,N_2781,N_2498);
nor U5048 (N_5048,N_2461,N_2829);
xor U5049 (N_5049,N_2770,N_136);
or U5050 (N_5050,N_260,N_2774);
or U5051 (N_5051,N_622,N_2675);
and U5052 (N_5052,N_1037,N_183);
nor U5053 (N_5053,N_937,N_2293);
and U5054 (N_5054,N_361,N_1473);
nand U5055 (N_5055,N_992,N_211);
and U5056 (N_5056,N_1151,N_88);
nand U5057 (N_5057,N_2520,N_2477);
nor U5058 (N_5058,N_648,N_2898);
and U5059 (N_5059,N_365,N_2924);
nand U5060 (N_5060,N_2382,N_1578);
or U5061 (N_5061,N_162,N_1390);
or U5062 (N_5062,N_787,N_1397);
nor U5063 (N_5063,N_638,N_2309);
or U5064 (N_5064,N_41,N_1728);
nand U5065 (N_5065,N_195,N_2343);
and U5066 (N_5066,N_1438,N_2926);
nand U5067 (N_5067,N_2170,N_730);
and U5068 (N_5068,N_1678,N_2977);
or U5069 (N_5069,N_275,N_2515);
nor U5070 (N_5070,N_2211,N_118);
nor U5071 (N_5071,N_2631,N_806);
nand U5072 (N_5072,N_1378,N_1411);
nor U5073 (N_5073,N_2630,N_289);
nand U5074 (N_5074,N_1967,N_1571);
nand U5075 (N_5075,N_61,N_2);
nor U5076 (N_5076,N_2815,N_131);
and U5077 (N_5077,N_1054,N_2649);
and U5078 (N_5078,N_82,N_227);
or U5079 (N_5079,N_1717,N_2);
nand U5080 (N_5080,N_138,N_1533);
nand U5081 (N_5081,N_488,N_430);
nand U5082 (N_5082,N_1237,N_1504);
nand U5083 (N_5083,N_197,N_373);
or U5084 (N_5084,N_277,N_1821);
or U5085 (N_5085,N_91,N_2487);
nand U5086 (N_5086,N_127,N_2746);
or U5087 (N_5087,N_1459,N_2913);
or U5088 (N_5088,N_2653,N_820);
nand U5089 (N_5089,N_2089,N_1344);
and U5090 (N_5090,N_2519,N_69);
nor U5091 (N_5091,N_626,N_224);
and U5092 (N_5092,N_2145,N_1841);
nand U5093 (N_5093,N_1692,N_2954);
nand U5094 (N_5094,N_192,N_2469);
or U5095 (N_5095,N_2153,N_728);
and U5096 (N_5096,N_2581,N_941);
or U5097 (N_5097,N_49,N_2899);
nor U5098 (N_5098,N_1207,N_2740);
nor U5099 (N_5099,N_644,N_1542);
or U5100 (N_5100,N_1334,N_1299);
and U5101 (N_5101,N_2398,N_172);
or U5102 (N_5102,N_1307,N_929);
nor U5103 (N_5103,N_2243,N_1822);
or U5104 (N_5104,N_294,N_2399);
nor U5105 (N_5105,N_2085,N_2914);
nand U5106 (N_5106,N_1924,N_2213);
nand U5107 (N_5107,N_1749,N_189);
nand U5108 (N_5108,N_463,N_2681);
or U5109 (N_5109,N_2334,N_1875);
or U5110 (N_5110,N_1473,N_688);
or U5111 (N_5111,N_888,N_2782);
nor U5112 (N_5112,N_2539,N_134);
nand U5113 (N_5113,N_2126,N_227);
nor U5114 (N_5114,N_479,N_80);
nor U5115 (N_5115,N_1393,N_80);
and U5116 (N_5116,N_790,N_2151);
and U5117 (N_5117,N_2717,N_112);
and U5118 (N_5118,N_144,N_2413);
and U5119 (N_5119,N_1614,N_937);
and U5120 (N_5120,N_909,N_386);
nor U5121 (N_5121,N_212,N_1721);
and U5122 (N_5122,N_761,N_1292);
nand U5123 (N_5123,N_2088,N_1542);
or U5124 (N_5124,N_1770,N_1328);
nor U5125 (N_5125,N_588,N_2028);
nand U5126 (N_5126,N_574,N_474);
nor U5127 (N_5127,N_1170,N_1325);
nand U5128 (N_5128,N_774,N_388);
and U5129 (N_5129,N_2338,N_1344);
and U5130 (N_5130,N_2023,N_544);
nand U5131 (N_5131,N_2003,N_1125);
or U5132 (N_5132,N_1952,N_945);
and U5133 (N_5133,N_361,N_15);
and U5134 (N_5134,N_613,N_2702);
nand U5135 (N_5135,N_1583,N_867);
nor U5136 (N_5136,N_1972,N_1289);
or U5137 (N_5137,N_1977,N_194);
and U5138 (N_5138,N_881,N_306);
nor U5139 (N_5139,N_1183,N_1019);
and U5140 (N_5140,N_680,N_2605);
nand U5141 (N_5141,N_1942,N_1271);
nand U5142 (N_5142,N_2744,N_499);
and U5143 (N_5143,N_1018,N_2723);
nor U5144 (N_5144,N_1258,N_2810);
and U5145 (N_5145,N_1448,N_1908);
nand U5146 (N_5146,N_944,N_928);
nor U5147 (N_5147,N_689,N_2612);
nand U5148 (N_5148,N_329,N_2385);
or U5149 (N_5149,N_422,N_2017);
nor U5150 (N_5150,N_2744,N_2389);
nand U5151 (N_5151,N_2200,N_882);
or U5152 (N_5152,N_1796,N_132);
or U5153 (N_5153,N_1202,N_2056);
and U5154 (N_5154,N_1774,N_553);
nand U5155 (N_5155,N_966,N_1271);
and U5156 (N_5156,N_1738,N_315);
or U5157 (N_5157,N_790,N_566);
nor U5158 (N_5158,N_334,N_29);
and U5159 (N_5159,N_865,N_89);
or U5160 (N_5160,N_1574,N_707);
or U5161 (N_5161,N_1609,N_1070);
nand U5162 (N_5162,N_2536,N_2779);
or U5163 (N_5163,N_1998,N_2824);
nand U5164 (N_5164,N_2807,N_1890);
or U5165 (N_5165,N_1546,N_476);
and U5166 (N_5166,N_141,N_2275);
nor U5167 (N_5167,N_810,N_2673);
nand U5168 (N_5168,N_2402,N_1054);
or U5169 (N_5169,N_454,N_840);
nand U5170 (N_5170,N_2767,N_618);
nand U5171 (N_5171,N_250,N_2964);
nand U5172 (N_5172,N_1726,N_412);
or U5173 (N_5173,N_2933,N_2059);
or U5174 (N_5174,N_1041,N_1311);
nor U5175 (N_5175,N_459,N_790);
nand U5176 (N_5176,N_2905,N_589);
or U5177 (N_5177,N_213,N_2295);
nor U5178 (N_5178,N_50,N_2960);
nand U5179 (N_5179,N_2401,N_182);
or U5180 (N_5180,N_158,N_2617);
nand U5181 (N_5181,N_1397,N_1364);
nor U5182 (N_5182,N_1077,N_2132);
nor U5183 (N_5183,N_467,N_2524);
and U5184 (N_5184,N_1049,N_1970);
or U5185 (N_5185,N_1231,N_1369);
and U5186 (N_5186,N_2089,N_2907);
nor U5187 (N_5187,N_2925,N_453);
and U5188 (N_5188,N_1603,N_2192);
xor U5189 (N_5189,N_1665,N_298);
nor U5190 (N_5190,N_1312,N_219);
nand U5191 (N_5191,N_2794,N_99);
and U5192 (N_5192,N_798,N_2944);
and U5193 (N_5193,N_2024,N_2200);
nor U5194 (N_5194,N_1181,N_430);
or U5195 (N_5195,N_793,N_1783);
or U5196 (N_5196,N_18,N_1814);
or U5197 (N_5197,N_1936,N_2098);
nor U5198 (N_5198,N_2605,N_2845);
nor U5199 (N_5199,N_2230,N_2589);
nor U5200 (N_5200,N_2999,N_702);
nor U5201 (N_5201,N_1114,N_1595);
or U5202 (N_5202,N_508,N_2728);
or U5203 (N_5203,N_1304,N_1842);
and U5204 (N_5204,N_89,N_2194);
and U5205 (N_5205,N_2791,N_1267);
or U5206 (N_5206,N_2502,N_572);
and U5207 (N_5207,N_2437,N_1765);
nor U5208 (N_5208,N_505,N_2447);
nor U5209 (N_5209,N_1657,N_2021);
xor U5210 (N_5210,N_1938,N_1177);
nor U5211 (N_5211,N_1639,N_2749);
and U5212 (N_5212,N_2468,N_238);
and U5213 (N_5213,N_2548,N_2298);
and U5214 (N_5214,N_803,N_1806);
nand U5215 (N_5215,N_2581,N_53);
or U5216 (N_5216,N_2232,N_1971);
nand U5217 (N_5217,N_493,N_1278);
nand U5218 (N_5218,N_2958,N_1128);
and U5219 (N_5219,N_1783,N_2502);
or U5220 (N_5220,N_1251,N_778);
or U5221 (N_5221,N_2941,N_2929);
xnor U5222 (N_5222,N_1037,N_87);
nor U5223 (N_5223,N_723,N_1756);
nand U5224 (N_5224,N_2385,N_2586);
and U5225 (N_5225,N_2064,N_1166);
nand U5226 (N_5226,N_1269,N_956);
nand U5227 (N_5227,N_1829,N_85);
and U5228 (N_5228,N_2733,N_584);
and U5229 (N_5229,N_2503,N_2807);
nand U5230 (N_5230,N_1499,N_1448);
nand U5231 (N_5231,N_736,N_1635);
nand U5232 (N_5232,N_1982,N_1877);
and U5233 (N_5233,N_2233,N_939);
or U5234 (N_5234,N_2526,N_849);
nand U5235 (N_5235,N_2409,N_1613);
or U5236 (N_5236,N_1403,N_2731);
and U5237 (N_5237,N_422,N_834);
nand U5238 (N_5238,N_2903,N_373);
nor U5239 (N_5239,N_2703,N_2057);
nor U5240 (N_5240,N_418,N_857);
nor U5241 (N_5241,N_558,N_2906);
nand U5242 (N_5242,N_2641,N_2773);
nand U5243 (N_5243,N_1340,N_989);
or U5244 (N_5244,N_919,N_2127);
nor U5245 (N_5245,N_2523,N_2556);
nor U5246 (N_5246,N_530,N_203);
and U5247 (N_5247,N_1906,N_760);
nor U5248 (N_5248,N_2083,N_1612);
nor U5249 (N_5249,N_2230,N_1654);
nand U5250 (N_5250,N_2012,N_2081);
or U5251 (N_5251,N_1448,N_1301);
and U5252 (N_5252,N_666,N_2128);
or U5253 (N_5253,N_654,N_1193);
or U5254 (N_5254,N_1939,N_2138);
nor U5255 (N_5255,N_1744,N_93);
nor U5256 (N_5256,N_1285,N_698);
or U5257 (N_5257,N_183,N_963);
or U5258 (N_5258,N_260,N_376);
and U5259 (N_5259,N_900,N_248);
and U5260 (N_5260,N_1601,N_1846);
xor U5261 (N_5261,N_869,N_2430);
and U5262 (N_5262,N_1926,N_1550);
and U5263 (N_5263,N_1153,N_1609);
nand U5264 (N_5264,N_1990,N_1925);
nor U5265 (N_5265,N_237,N_18);
or U5266 (N_5266,N_1189,N_1842);
nor U5267 (N_5267,N_2104,N_2924);
and U5268 (N_5268,N_2118,N_57);
nand U5269 (N_5269,N_1918,N_1248);
xnor U5270 (N_5270,N_917,N_1786);
nand U5271 (N_5271,N_1780,N_1418);
or U5272 (N_5272,N_1806,N_2228);
nand U5273 (N_5273,N_2170,N_287);
nand U5274 (N_5274,N_2253,N_942);
or U5275 (N_5275,N_29,N_1750);
nand U5276 (N_5276,N_1450,N_1688);
nand U5277 (N_5277,N_872,N_84);
and U5278 (N_5278,N_1112,N_1130);
nor U5279 (N_5279,N_2827,N_2932);
and U5280 (N_5280,N_12,N_2339);
nand U5281 (N_5281,N_604,N_1833);
and U5282 (N_5282,N_1938,N_2163);
nor U5283 (N_5283,N_220,N_1438);
nand U5284 (N_5284,N_1824,N_1092);
and U5285 (N_5285,N_2186,N_2913);
and U5286 (N_5286,N_1810,N_2241);
nor U5287 (N_5287,N_29,N_1423);
or U5288 (N_5288,N_2747,N_273);
or U5289 (N_5289,N_696,N_148);
and U5290 (N_5290,N_2035,N_2873);
nand U5291 (N_5291,N_2616,N_1436);
and U5292 (N_5292,N_2497,N_493);
or U5293 (N_5293,N_1599,N_467);
nand U5294 (N_5294,N_901,N_2667);
nor U5295 (N_5295,N_29,N_2402);
nand U5296 (N_5296,N_1955,N_2809);
and U5297 (N_5297,N_2437,N_2951);
and U5298 (N_5298,N_1865,N_974);
and U5299 (N_5299,N_1843,N_2870);
nand U5300 (N_5300,N_885,N_1289);
or U5301 (N_5301,N_868,N_2868);
or U5302 (N_5302,N_2717,N_1101);
nor U5303 (N_5303,N_2495,N_2871);
or U5304 (N_5304,N_675,N_2447);
and U5305 (N_5305,N_262,N_31);
and U5306 (N_5306,N_2299,N_579);
or U5307 (N_5307,N_29,N_350);
and U5308 (N_5308,N_2296,N_2660);
and U5309 (N_5309,N_201,N_1091);
nand U5310 (N_5310,N_2357,N_2778);
and U5311 (N_5311,N_68,N_759);
nor U5312 (N_5312,N_1891,N_546);
or U5313 (N_5313,N_1459,N_1282);
nor U5314 (N_5314,N_1285,N_2807);
and U5315 (N_5315,N_1177,N_2273);
or U5316 (N_5316,N_2894,N_717);
and U5317 (N_5317,N_1882,N_1363);
nand U5318 (N_5318,N_73,N_2631);
nor U5319 (N_5319,N_1891,N_2262);
nor U5320 (N_5320,N_1524,N_752);
nand U5321 (N_5321,N_380,N_988);
nor U5322 (N_5322,N_2471,N_1561);
nor U5323 (N_5323,N_1597,N_1489);
nor U5324 (N_5324,N_2762,N_2837);
nor U5325 (N_5325,N_2353,N_1756);
and U5326 (N_5326,N_200,N_2382);
nor U5327 (N_5327,N_1808,N_1721);
or U5328 (N_5328,N_1278,N_2827);
or U5329 (N_5329,N_2451,N_2833);
and U5330 (N_5330,N_1000,N_1368);
nand U5331 (N_5331,N_453,N_1458);
or U5332 (N_5332,N_2595,N_1469);
and U5333 (N_5333,N_2132,N_1617);
nor U5334 (N_5334,N_2953,N_694);
and U5335 (N_5335,N_1853,N_451);
and U5336 (N_5336,N_2506,N_2269);
nand U5337 (N_5337,N_128,N_414);
nand U5338 (N_5338,N_772,N_297);
nand U5339 (N_5339,N_1391,N_1577);
or U5340 (N_5340,N_2842,N_2507);
or U5341 (N_5341,N_2096,N_1743);
or U5342 (N_5342,N_456,N_2253);
or U5343 (N_5343,N_194,N_2407);
or U5344 (N_5344,N_1934,N_339);
nand U5345 (N_5345,N_1993,N_2904);
nand U5346 (N_5346,N_984,N_1348);
or U5347 (N_5347,N_1618,N_281);
nand U5348 (N_5348,N_1292,N_2062);
and U5349 (N_5349,N_1455,N_1196);
or U5350 (N_5350,N_704,N_1113);
and U5351 (N_5351,N_309,N_606);
nor U5352 (N_5352,N_1149,N_2626);
nand U5353 (N_5353,N_1977,N_2166);
nand U5354 (N_5354,N_2545,N_1210);
and U5355 (N_5355,N_2554,N_2079);
and U5356 (N_5356,N_392,N_1579);
xnor U5357 (N_5357,N_1917,N_1650);
or U5358 (N_5358,N_1919,N_790);
or U5359 (N_5359,N_1968,N_829);
nand U5360 (N_5360,N_1171,N_1302);
or U5361 (N_5361,N_437,N_2056);
nand U5362 (N_5362,N_1765,N_1745);
nor U5363 (N_5363,N_2018,N_290);
nor U5364 (N_5364,N_519,N_1839);
nor U5365 (N_5365,N_576,N_660);
nor U5366 (N_5366,N_1054,N_2049);
and U5367 (N_5367,N_1540,N_346);
nor U5368 (N_5368,N_2502,N_1447);
nor U5369 (N_5369,N_1522,N_230);
or U5370 (N_5370,N_2958,N_1579);
or U5371 (N_5371,N_667,N_1476);
nor U5372 (N_5372,N_2049,N_2481);
nor U5373 (N_5373,N_1343,N_1327);
nand U5374 (N_5374,N_2065,N_2551);
nor U5375 (N_5375,N_2329,N_18);
or U5376 (N_5376,N_1632,N_1950);
or U5377 (N_5377,N_1523,N_2875);
nor U5378 (N_5378,N_2847,N_565);
or U5379 (N_5379,N_1139,N_2968);
nor U5380 (N_5380,N_1110,N_547);
or U5381 (N_5381,N_1954,N_2055);
or U5382 (N_5382,N_1267,N_877);
nand U5383 (N_5383,N_1347,N_2945);
or U5384 (N_5384,N_2607,N_141);
nand U5385 (N_5385,N_2678,N_199);
or U5386 (N_5386,N_1916,N_1354);
nor U5387 (N_5387,N_2547,N_2206);
nand U5388 (N_5388,N_2541,N_2016);
and U5389 (N_5389,N_2463,N_1739);
or U5390 (N_5390,N_151,N_600);
or U5391 (N_5391,N_2474,N_1696);
nand U5392 (N_5392,N_1348,N_2004);
or U5393 (N_5393,N_321,N_1445);
nor U5394 (N_5394,N_1489,N_562);
or U5395 (N_5395,N_1620,N_1687);
nand U5396 (N_5396,N_1756,N_176);
or U5397 (N_5397,N_1703,N_685);
nand U5398 (N_5398,N_666,N_1602);
nor U5399 (N_5399,N_1903,N_383);
and U5400 (N_5400,N_941,N_749);
nand U5401 (N_5401,N_592,N_1973);
nor U5402 (N_5402,N_2388,N_446);
and U5403 (N_5403,N_979,N_1453);
nand U5404 (N_5404,N_2879,N_1710);
or U5405 (N_5405,N_614,N_1994);
nand U5406 (N_5406,N_1048,N_1837);
nand U5407 (N_5407,N_269,N_1681);
nand U5408 (N_5408,N_775,N_2868);
nor U5409 (N_5409,N_2864,N_2521);
and U5410 (N_5410,N_167,N_579);
and U5411 (N_5411,N_1700,N_816);
nand U5412 (N_5412,N_564,N_553);
nand U5413 (N_5413,N_1192,N_357);
and U5414 (N_5414,N_1664,N_795);
and U5415 (N_5415,N_2036,N_1749);
nand U5416 (N_5416,N_1545,N_2291);
nor U5417 (N_5417,N_583,N_1682);
nand U5418 (N_5418,N_439,N_1195);
xor U5419 (N_5419,N_361,N_2664);
and U5420 (N_5420,N_1339,N_2819);
nand U5421 (N_5421,N_1346,N_1730);
or U5422 (N_5422,N_786,N_331);
nand U5423 (N_5423,N_2523,N_830);
or U5424 (N_5424,N_2139,N_1559);
nor U5425 (N_5425,N_2027,N_115);
and U5426 (N_5426,N_11,N_1927);
nand U5427 (N_5427,N_2913,N_2383);
nand U5428 (N_5428,N_1308,N_151);
and U5429 (N_5429,N_544,N_26);
and U5430 (N_5430,N_620,N_2516);
and U5431 (N_5431,N_2494,N_1136);
nand U5432 (N_5432,N_2970,N_1176);
nor U5433 (N_5433,N_2550,N_575);
nand U5434 (N_5434,N_466,N_1571);
or U5435 (N_5435,N_136,N_2075);
and U5436 (N_5436,N_1152,N_898);
nor U5437 (N_5437,N_874,N_519);
nor U5438 (N_5438,N_519,N_2572);
and U5439 (N_5439,N_2198,N_2695);
nand U5440 (N_5440,N_1913,N_321);
nor U5441 (N_5441,N_2202,N_61);
nor U5442 (N_5442,N_141,N_1050);
or U5443 (N_5443,N_2823,N_931);
and U5444 (N_5444,N_1041,N_153);
or U5445 (N_5445,N_870,N_1994);
nor U5446 (N_5446,N_589,N_2224);
or U5447 (N_5447,N_2223,N_75);
nor U5448 (N_5448,N_1138,N_152);
nor U5449 (N_5449,N_2276,N_1214);
nand U5450 (N_5450,N_291,N_3);
or U5451 (N_5451,N_805,N_257);
or U5452 (N_5452,N_910,N_1543);
nor U5453 (N_5453,N_2246,N_244);
and U5454 (N_5454,N_2141,N_712);
and U5455 (N_5455,N_2343,N_853);
or U5456 (N_5456,N_2715,N_1266);
nor U5457 (N_5457,N_2140,N_2733);
or U5458 (N_5458,N_2497,N_1767);
nor U5459 (N_5459,N_2363,N_259);
or U5460 (N_5460,N_2777,N_1171);
nor U5461 (N_5461,N_181,N_354);
and U5462 (N_5462,N_2983,N_1222);
nor U5463 (N_5463,N_2459,N_2220);
or U5464 (N_5464,N_276,N_2213);
or U5465 (N_5465,N_895,N_533);
and U5466 (N_5466,N_138,N_150);
nor U5467 (N_5467,N_385,N_557);
or U5468 (N_5468,N_1273,N_360);
and U5469 (N_5469,N_386,N_1970);
nor U5470 (N_5470,N_2587,N_2546);
nand U5471 (N_5471,N_201,N_343);
nand U5472 (N_5472,N_987,N_316);
nor U5473 (N_5473,N_1026,N_2378);
or U5474 (N_5474,N_2717,N_2890);
nor U5475 (N_5475,N_352,N_2289);
xor U5476 (N_5476,N_1817,N_495);
or U5477 (N_5477,N_2635,N_530);
nor U5478 (N_5478,N_1637,N_449);
or U5479 (N_5479,N_1081,N_354);
and U5480 (N_5480,N_2287,N_436);
nand U5481 (N_5481,N_1277,N_1996);
nor U5482 (N_5482,N_2183,N_2552);
or U5483 (N_5483,N_1508,N_1790);
nand U5484 (N_5484,N_1605,N_1618);
nand U5485 (N_5485,N_2456,N_653);
nand U5486 (N_5486,N_2740,N_1423);
nand U5487 (N_5487,N_1861,N_1170);
nor U5488 (N_5488,N_1326,N_646);
nor U5489 (N_5489,N_149,N_2440);
or U5490 (N_5490,N_1102,N_1494);
nor U5491 (N_5491,N_604,N_2847);
and U5492 (N_5492,N_332,N_119);
and U5493 (N_5493,N_2350,N_2130);
and U5494 (N_5494,N_2946,N_1917);
and U5495 (N_5495,N_309,N_701);
or U5496 (N_5496,N_1479,N_1729);
nand U5497 (N_5497,N_1250,N_1481);
nand U5498 (N_5498,N_1081,N_1768);
nand U5499 (N_5499,N_1691,N_1119);
nand U5500 (N_5500,N_1188,N_1845);
nor U5501 (N_5501,N_622,N_1930);
or U5502 (N_5502,N_2844,N_1699);
nor U5503 (N_5503,N_67,N_2865);
and U5504 (N_5504,N_126,N_1198);
nand U5505 (N_5505,N_19,N_2188);
and U5506 (N_5506,N_597,N_577);
or U5507 (N_5507,N_1647,N_1972);
and U5508 (N_5508,N_1459,N_1041);
and U5509 (N_5509,N_1753,N_1506);
and U5510 (N_5510,N_429,N_693);
nand U5511 (N_5511,N_2660,N_147);
nor U5512 (N_5512,N_597,N_332);
or U5513 (N_5513,N_1915,N_1974);
and U5514 (N_5514,N_2520,N_2436);
nand U5515 (N_5515,N_490,N_1202);
and U5516 (N_5516,N_255,N_985);
nor U5517 (N_5517,N_470,N_1195);
nand U5518 (N_5518,N_1214,N_533);
and U5519 (N_5519,N_2252,N_632);
or U5520 (N_5520,N_360,N_1790);
or U5521 (N_5521,N_397,N_2715);
or U5522 (N_5522,N_2010,N_897);
nand U5523 (N_5523,N_1207,N_2225);
xnor U5524 (N_5524,N_2092,N_2227);
or U5525 (N_5525,N_1648,N_1120);
xor U5526 (N_5526,N_1851,N_1559);
and U5527 (N_5527,N_2433,N_2279);
nand U5528 (N_5528,N_2590,N_2953);
nand U5529 (N_5529,N_1589,N_201);
nand U5530 (N_5530,N_1312,N_1283);
nand U5531 (N_5531,N_783,N_1753);
nand U5532 (N_5532,N_648,N_2938);
nor U5533 (N_5533,N_504,N_1838);
or U5534 (N_5534,N_651,N_1853);
nand U5535 (N_5535,N_2518,N_749);
nand U5536 (N_5536,N_2103,N_2789);
nor U5537 (N_5537,N_1623,N_29);
nand U5538 (N_5538,N_384,N_2389);
nor U5539 (N_5539,N_2928,N_82);
or U5540 (N_5540,N_386,N_2351);
nor U5541 (N_5541,N_309,N_1447);
nor U5542 (N_5542,N_1094,N_262);
and U5543 (N_5543,N_1377,N_2980);
or U5544 (N_5544,N_2365,N_2114);
or U5545 (N_5545,N_703,N_2546);
or U5546 (N_5546,N_1286,N_1744);
nand U5547 (N_5547,N_1311,N_1345);
and U5548 (N_5548,N_1538,N_1807);
nor U5549 (N_5549,N_239,N_1777);
nand U5550 (N_5550,N_1901,N_2224);
nand U5551 (N_5551,N_173,N_2396);
nor U5552 (N_5552,N_746,N_2377);
or U5553 (N_5553,N_2962,N_1014);
nor U5554 (N_5554,N_2985,N_185);
and U5555 (N_5555,N_2889,N_2916);
or U5556 (N_5556,N_1351,N_2338);
or U5557 (N_5557,N_1225,N_779);
xor U5558 (N_5558,N_2573,N_1216);
nand U5559 (N_5559,N_2660,N_1750);
xor U5560 (N_5560,N_2075,N_2707);
nand U5561 (N_5561,N_387,N_49);
nand U5562 (N_5562,N_1802,N_90);
and U5563 (N_5563,N_180,N_1426);
nand U5564 (N_5564,N_153,N_2922);
nand U5565 (N_5565,N_444,N_2401);
nand U5566 (N_5566,N_2902,N_1924);
nand U5567 (N_5567,N_1761,N_2110);
nand U5568 (N_5568,N_1790,N_1522);
nand U5569 (N_5569,N_492,N_463);
nand U5570 (N_5570,N_1164,N_1869);
and U5571 (N_5571,N_2386,N_617);
and U5572 (N_5572,N_1657,N_1273);
nor U5573 (N_5573,N_770,N_1879);
or U5574 (N_5574,N_2617,N_2523);
and U5575 (N_5575,N_859,N_734);
nand U5576 (N_5576,N_1037,N_2901);
and U5577 (N_5577,N_2475,N_2625);
or U5578 (N_5578,N_1473,N_1868);
or U5579 (N_5579,N_2400,N_618);
or U5580 (N_5580,N_1512,N_1173);
nor U5581 (N_5581,N_2029,N_1545);
nand U5582 (N_5582,N_2788,N_56);
and U5583 (N_5583,N_672,N_1558);
nand U5584 (N_5584,N_958,N_1372);
nor U5585 (N_5585,N_1748,N_73);
and U5586 (N_5586,N_1473,N_1045);
nor U5587 (N_5587,N_1282,N_1557);
nor U5588 (N_5588,N_875,N_2925);
or U5589 (N_5589,N_2982,N_1912);
nand U5590 (N_5590,N_546,N_1873);
or U5591 (N_5591,N_1607,N_635);
nand U5592 (N_5592,N_1892,N_625);
nor U5593 (N_5593,N_130,N_2571);
nor U5594 (N_5594,N_1199,N_454);
nor U5595 (N_5595,N_115,N_243);
nand U5596 (N_5596,N_162,N_2346);
nor U5597 (N_5597,N_1398,N_1549);
nor U5598 (N_5598,N_2764,N_1444);
or U5599 (N_5599,N_2059,N_1221);
or U5600 (N_5600,N_737,N_2248);
or U5601 (N_5601,N_697,N_1584);
and U5602 (N_5602,N_1261,N_1242);
and U5603 (N_5603,N_2256,N_599);
nand U5604 (N_5604,N_533,N_475);
and U5605 (N_5605,N_2305,N_696);
nand U5606 (N_5606,N_2217,N_2967);
or U5607 (N_5607,N_520,N_1640);
or U5608 (N_5608,N_1601,N_175);
nand U5609 (N_5609,N_1794,N_449);
nor U5610 (N_5610,N_996,N_442);
or U5611 (N_5611,N_811,N_181);
nand U5612 (N_5612,N_1453,N_2256);
nor U5613 (N_5613,N_1567,N_61);
or U5614 (N_5614,N_2943,N_2949);
nor U5615 (N_5615,N_324,N_1366);
nand U5616 (N_5616,N_1946,N_1310);
or U5617 (N_5617,N_1441,N_1069);
or U5618 (N_5618,N_1915,N_2240);
nor U5619 (N_5619,N_970,N_879);
or U5620 (N_5620,N_1505,N_249);
nand U5621 (N_5621,N_2340,N_175);
xnor U5622 (N_5622,N_2557,N_2407);
and U5623 (N_5623,N_439,N_1778);
nand U5624 (N_5624,N_1420,N_1851);
nor U5625 (N_5625,N_1097,N_1963);
nand U5626 (N_5626,N_1255,N_1487);
nor U5627 (N_5627,N_2743,N_1841);
nand U5628 (N_5628,N_621,N_77);
nor U5629 (N_5629,N_2518,N_2156);
and U5630 (N_5630,N_967,N_639);
or U5631 (N_5631,N_2392,N_2467);
nor U5632 (N_5632,N_683,N_2983);
nor U5633 (N_5633,N_799,N_1216);
and U5634 (N_5634,N_1451,N_1970);
or U5635 (N_5635,N_2583,N_1887);
and U5636 (N_5636,N_1685,N_1616);
and U5637 (N_5637,N_1524,N_589);
nand U5638 (N_5638,N_1543,N_770);
nand U5639 (N_5639,N_1359,N_2802);
xor U5640 (N_5640,N_1891,N_1092);
nor U5641 (N_5641,N_1616,N_1658);
and U5642 (N_5642,N_581,N_39);
nand U5643 (N_5643,N_744,N_2358);
nor U5644 (N_5644,N_1406,N_1539);
nand U5645 (N_5645,N_1015,N_2935);
nor U5646 (N_5646,N_2548,N_1671);
or U5647 (N_5647,N_844,N_175);
nor U5648 (N_5648,N_2688,N_1296);
and U5649 (N_5649,N_1244,N_2514);
nand U5650 (N_5650,N_141,N_2823);
nor U5651 (N_5651,N_2857,N_2327);
or U5652 (N_5652,N_2811,N_1467);
nor U5653 (N_5653,N_1727,N_2844);
nor U5654 (N_5654,N_1907,N_1993);
nor U5655 (N_5655,N_290,N_1723);
and U5656 (N_5656,N_2708,N_731);
or U5657 (N_5657,N_1697,N_1399);
nor U5658 (N_5658,N_118,N_2876);
and U5659 (N_5659,N_693,N_2724);
nand U5660 (N_5660,N_1476,N_2437);
or U5661 (N_5661,N_660,N_815);
or U5662 (N_5662,N_2726,N_1465);
nand U5663 (N_5663,N_2426,N_339);
or U5664 (N_5664,N_1300,N_2751);
and U5665 (N_5665,N_2419,N_1191);
and U5666 (N_5666,N_400,N_2054);
nand U5667 (N_5667,N_2256,N_2762);
nor U5668 (N_5668,N_2187,N_2446);
and U5669 (N_5669,N_483,N_202);
nand U5670 (N_5670,N_2197,N_1812);
nor U5671 (N_5671,N_1694,N_338);
or U5672 (N_5672,N_1836,N_972);
or U5673 (N_5673,N_515,N_2950);
nor U5674 (N_5674,N_594,N_1655);
nand U5675 (N_5675,N_2833,N_776);
nand U5676 (N_5676,N_1456,N_1050);
nor U5677 (N_5677,N_83,N_31);
and U5678 (N_5678,N_419,N_2917);
nand U5679 (N_5679,N_1031,N_2317);
nor U5680 (N_5680,N_2124,N_2004);
nand U5681 (N_5681,N_1955,N_1864);
nor U5682 (N_5682,N_1662,N_1701);
nand U5683 (N_5683,N_2874,N_507);
nand U5684 (N_5684,N_2513,N_2133);
nor U5685 (N_5685,N_662,N_2935);
nor U5686 (N_5686,N_1588,N_955);
nand U5687 (N_5687,N_2975,N_717);
nand U5688 (N_5688,N_1944,N_1348);
and U5689 (N_5689,N_1855,N_2677);
nand U5690 (N_5690,N_2854,N_1326);
and U5691 (N_5691,N_1460,N_1579);
nand U5692 (N_5692,N_2162,N_2004);
and U5693 (N_5693,N_2905,N_194);
nor U5694 (N_5694,N_1492,N_1458);
nand U5695 (N_5695,N_1927,N_523);
and U5696 (N_5696,N_2713,N_638);
or U5697 (N_5697,N_799,N_1680);
or U5698 (N_5698,N_2092,N_2154);
nor U5699 (N_5699,N_387,N_1247);
nor U5700 (N_5700,N_2204,N_2608);
nor U5701 (N_5701,N_1234,N_278);
nor U5702 (N_5702,N_791,N_2028);
or U5703 (N_5703,N_1656,N_2272);
nand U5704 (N_5704,N_2666,N_2779);
nor U5705 (N_5705,N_2115,N_49);
nor U5706 (N_5706,N_1454,N_1251);
nor U5707 (N_5707,N_470,N_857);
and U5708 (N_5708,N_289,N_1411);
and U5709 (N_5709,N_793,N_2703);
and U5710 (N_5710,N_1844,N_2877);
or U5711 (N_5711,N_1815,N_1261);
and U5712 (N_5712,N_2282,N_1965);
and U5713 (N_5713,N_1813,N_1184);
and U5714 (N_5714,N_2895,N_2030);
or U5715 (N_5715,N_1917,N_2380);
and U5716 (N_5716,N_1103,N_2213);
or U5717 (N_5717,N_1860,N_2102);
nand U5718 (N_5718,N_649,N_2473);
and U5719 (N_5719,N_29,N_1993);
nor U5720 (N_5720,N_259,N_2998);
nand U5721 (N_5721,N_2445,N_1698);
nand U5722 (N_5722,N_1435,N_1238);
nor U5723 (N_5723,N_1650,N_1547);
and U5724 (N_5724,N_46,N_2930);
nor U5725 (N_5725,N_1400,N_2890);
and U5726 (N_5726,N_1577,N_2414);
nor U5727 (N_5727,N_935,N_1656);
and U5728 (N_5728,N_2963,N_484);
and U5729 (N_5729,N_2761,N_2442);
nor U5730 (N_5730,N_1601,N_2821);
nand U5731 (N_5731,N_1936,N_1304);
nor U5732 (N_5732,N_69,N_2242);
and U5733 (N_5733,N_114,N_1386);
or U5734 (N_5734,N_1764,N_2330);
or U5735 (N_5735,N_2551,N_419);
or U5736 (N_5736,N_1857,N_2065);
nor U5737 (N_5737,N_45,N_185);
nor U5738 (N_5738,N_1463,N_1926);
nor U5739 (N_5739,N_38,N_1074);
or U5740 (N_5740,N_2810,N_1068);
nor U5741 (N_5741,N_2074,N_1472);
nor U5742 (N_5742,N_2715,N_302);
nand U5743 (N_5743,N_88,N_2942);
nand U5744 (N_5744,N_1163,N_1057);
nand U5745 (N_5745,N_2932,N_2964);
nand U5746 (N_5746,N_2413,N_887);
nand U5747 (N_5747,N_2217,N_792);
nor U5748 (N_5748,N_529,N_996);
nand U5749 (N_5749,N_840,N_535);
and U5750 (N_5750,N_1843,N_1318);
or U5751 (N_5751,N_1724,N_623);
and U5752 (N_5752,N_1261,N_5);
nor U5753 (N_5753,N_934,N_2059);
xor U5754 (N_5754,N_2663,N_1102);
nand U5755 (N_5755,N_2109,N_1737);
nor U5756 (N_5756,N_56,N_2780);
nor U5757 (N_5757,N_1973,N_903);
or U5758 (N_5758,N_2642,N_628);
nor U5759 (N_5759,N_2894,N_2581);
and U5760 (N_5760,N_437,N_2621);
and U5761 (N_5761,N_1383,N_553);
or U5762 (N_5762,N_2076,N_2950);
nand U5763 (N_5763,N_492,N_2462);
nor U5764 (N_5764,N_1278,N_967);
nand U5765 (N_5765,N_1838,N_1352);
or U5766 (N_5766,N_2335,N_1641);
nor U5767 (N_5767,N_1351,N_2954);
nor U5768 (N_5768,N_369,N_2845);
and U5769 (N_5769,N_2744,N_1917);
and U5770 (N_5770,N_1122,N_1880);
and U5771 (N_5771,N_2217,N_1882);
and U5772 (N_5772,N_2201,N_1515);
and U5773 (N_5773,N_1770,N_530);
and U5774 (N_5774,N_1977,N_2440);
and U5775 (N_5775,N_702,N_2731);
nor U5776 (N_5776,N_2447,N_1421);
nand U5777 (N_5777,N_772,N_1731);
and U5778 (N_5778,N_274,N_479);
nor U5779 (N_5779,N_1180,N_476);
nand U5780 (N_5780,N_761,N_1710);
or U5781 (N_5781,N_787,N_2862);
and U5782 (N_5782,N_1297,N_204);
nor U5783 (N_5783,N_733,N_2567);
nor U5784 (N_5784,N_609,N_2900);
nand U5785 (N_5785,N_1771,N_1291);
nor U5786 (N_5786,N_705,N_1053);
and U5787 (N_5787,N_570,N_736);
or U5788 (N_5788,N_1283,N_163);
or U5789 (N_5789,N_1444,N_856);
and U5790 (N_5790,N_2509,N_1892);
and U5791 (N_5791,N_1065,N_1388);
and U5792 (N_5792,N_2706,N_2198);
or U5793 (N_5793,N_2625,N_1637);
nor U5794 (N_5794,N_1336,N_281);
nor U5795 (N_5795,N_2565,N_156);
nand U5796 (N_5796,N_2161,N_2392);
nor U5797 (N_5797,N_326,N_1401);
nor U5798 (N_5798,N_1090,N_402);
nor U5799 (N_5799,N_2889,N_5);
or U5800 (N_5800,N_713,N_699);
or U5801 (N_5801,N_1039,N_985);
nor U5802 (N_5802,N_2599,N_1187);
nor U5803 (N_5803,N_1048,N_326);
and U5804 (N_5804,N_1413,N_1498);
and U5805 (N_5805,N_1063,N_175);
nand U5806 (N_5806,N_757,N_1940);
nand U5807 (N_5807,N_884,N_2159);
and U5808 (N_5808,N_125,N_1297);
and U5809 (N_5809,N_413,N_489);
and U5810 (N_5810,N_228,N_152);
and U5811 (N_5811,N_1695,N_2816);
and U5812 (N_5812,N_1764,N_1539);
nand U5813 (N_5813,N_1610,N_1742);
nor U5814 (N_5814,N_2440,N_952);
nor U5815 (N_5815,N_2091,N_2564);
or U5816 (N_5816,N_1312,N_2137);
nor U5817 (N_5817,N_2377,N_1736);
nor U5818 (N_5818,N_1583,N_383);
or U5819 (N_5819,N_1224,N_689);
nand U5820 (N_5820,N_260,N_2386);
or U5821 (N_5821,N_1044,N_1979);
or U5822 (N_5822,N_2789,N_1727);
and U5823 (N_5823,N_1297,N_2295);
or U5824 (N_5824,N_2623,N_299);
nor U5825 (N_5825,N_910,N_762);
and U5826 (N_5826,N_2856,N_102);
or U5827 (N_5827,N_1793,N_2674);
or U5828 (N_5828,N_2987,N_2872);
and U5829 (N_5829,N_651,N_512);
nor U5830 (N_5830,N_2365,N_1619);
nand U5831 (N_5831,N_585,N_1154);
nand U5832 (N_5832,N_1595,N_657);
and U5833 (N_5833,N_2375,N_2170);
nor U5834 (N_5834,N_2859,N_2313);
and U5835 (N_5835,N_1030,N_596);
nand U5836 (N_5836,N_2366,N_1437);
nor U5837 (N_5837,N_158,N_1709);
nand U5838 (N_5838,N_993,N_2358);
or U5839 (N_5839,N_2857,N_483);
and U5840 (N_5840,N_2315,N_2598);
nor U5841 (N_5841,N_1354,N_66);
and U5842 (N_5842,N_2851,N_1327);
or U5843 (N_5843,N_2202,N_1932);
and U5844 (N_5844,N_1458,N_139);
nand U5845 (N_5845,N_1480,N_623);
nor U5846 (N_5846,N_1387,N_1609);
nand U5847 (N_5847,N_2493,N_388);
nand U5848 (N_5848,N_948,N_1964);
and U5849 (N_5849,N_634,N_2445);
and U5850 (N_5850,N_785,N_130);
or U5851 (N_5851,N_1603,N_2884);
and U5852 (N_5852,N_130,N_640);
and U5853 (N_5853,N_636,N_1711);
or U5854 (N_5854,N_1273,N_1373);
nor U5855 (N_5855,N_2203,N_2941);
or U5856 (N_5856,N_883,N_215);
nor U5857 (N_5857,N_224,N_2386);
and U5858 (N_5858,N_2790,N_2579);
nor U5859 (N_5859,N_1703,N_1448);
or U5860 (N_5860,N_1617,N_2198);
nand U5861 (N_5861,N_860,N_1591);
nand U5862 (N_5862,N_2906,N_1440);
and U5863 (N_5863,N_1672,N_1270);
nor U5864 (N_5864,N_448,N_1826);
and U5865 (N_5865,N_629,N_2975);
nor U5866 (N_5866,N_90,N_1393);
and U5867 (N_5867,N_1933,N_2134);
or U5868 (N_5868,N_1370,N_576);
and U5869 (N_5869,N_798,N_2053);
or U5870 (N_5870,N_1320,N_253);
or U5871 (N_5871,N_2285,N_2996);
and U5872 (N_5872,N_374,N_1864);
and U5873 (N_5873,N_1902,N_1407);
nor U5874 (N_5874,N_1447,N_2280);
nor U5875 (N_5875,N_405,N_2863);
nor U5876 (N_5876,N_309,N_1572);
nand U5877 (N_5877,N_650,N_2699);
or U5878 (N_5878,N_2447,N_1033);
or U5879 (N_5879,N_2046,N_2142);
nor U5880 (N_5880,N_2522,N_2249);
or U5881 (N_5881,N_1201,N_15);
nor U5882 (N_5882,N_1697,N_903);
and U5883 (N_5883,N_1845,N_501);
nor U5884 (N_5884,N_1252,N_1262);
nor U5885 (N_5885,N_522,N_1259);
nor U5886 (N_5886,N_127,N_63);
nor U5887 (N_5887,N_1889,N_1249);
or U5888 (N_5888,N_1712,N_1407);
and U5889 (N_5889,N_863,N_286);
nand U5890 (N_5890,N_2414,N_1547);
nand U5891 (N_5891,N_1945,N_1764);
and U5892 (N_5892,N_23,N_679);
nor U5893 (N_5893,N_2690,N_375);
or U5894 (N_5894,N_1406,N_1033);
nor U5895 (N_5895,N_2104,N_1737);
or U5896 (N_5896,N_1545,N_1843);
and U5897 (N_5897,N_638,N_2668);
nor U5898 (N_5898,N_904,N_1075);
nor U5899 (N_5899,N_1838,N_85);
or U5900 (N_5900,N_1580,N_2175);
and U5901 (N_5901,N_2362,N_2576);
and U5902 (N_5902,N_2457,N_2117);
and U5903 (N_5903,N_1622,N_52);
or U5904 (N_5904,N_2332,N_1993);
or U5905 (N_5905,N_1897,N_76);
nand U5906 (N_5906,N_2435,N_2194);
or U5907 (N_5907,N_39,N_1137);
or U5908 (N_5908,N_2553,N_1048);
nand U5909 (N_5909,N_731,N_210);
or U5910 (N_5910,N_1161,N_1269);
nand U5911 (N_5911,N_2015,N_2375);
or U5912 (N_5912,N_1840,N_1739);
and U5913 (N_5913,N_2520,N_1117);
or U5914 (N_5914,N_1118,N_1180);
and U5915 (N_5915,N_1705,N_2994);
nand U5916 (N_5916,N_686,N_364);
or U5917 (N_5917,N_1641,N_108);
or U5918 (N_5918,N_1221,N_1555);
nand U5919 (N_5919,N_292,N_2286);
and U5920 (N_5920,N_2463,N_2032);
or U5921 (N_5921,N_808,N_2259);
and U5922 (N_5922,N_2802,N_2653);
nor U5923 (N_5923,N_2114,N_1135);
or U5924 (N_5924,N_1916,N_1986);
nor U5925 (N_5925,N_631,N_2460);
and U5926 (N_5926,N_1840,N_1417);
nand U5927 (N_5927,N_2352,N_1418);
nor U5928 (N_5928,N_14,N_1474);
and U5929 (N_5929,N_2821,N_2395);
or U5930 (N_5930,N_1646,N_1898);
and U5931 (N_5931,N_2442,N_2620);
or U5932 (N_5932,N_2454,N_545);
nor U5933 (N_5933,N_2541,N_1924);
nand U5934 (N_5934,N_2842,N_1130);
or U5935 (N_5935,N_122,N_111);
nand U5936 (N_5936,N_2436,N_2654);
or U5937 (N_5937,N_2946,N_2695);
or U5938 (N_5938,N_1162,N_2479);
nor U5939 (N_5939,N_2940,N_426);
or U5940 (N_5940,N_575,N_2559);
nor U5941 (N_5941,N_911,N_949);
or U5942 (N_5942,N_423,N_2875);
nand U5943 (N_5943,N_1909,N_1220);
nor U5944 (N_5944,N_2775,N_223);
or U5945 (N_5945,N_437,N_1564);
nand U5946 (N_5946,N_1478,N_836);
nand U5947 (N_5947,N_2468,N_1400);
nor U5948 (N_5948,N_2173,N_1156);
and U5949 (N_5949,N_82,N_510);
or U5950 (N_5950,N_1683,N_2408);
and U5951 (N_5951,N_1974,N_2404);
nand U5952 (N_5952,N_1124,N_2003);
or U5953 (N_5953,N_2816,N_775);
nor U5954 (N_5954,N_934,N_1141);
nor U5955 (N_5955,N_1386,N_2301);
nor U5956 (N_5956,N_1431,N_1789);
and U5957 (N_5957,N_1586,N_1172);
and U5958 (N_5958,N_2577,N_1937);
nand U5959 (N_5959,N_706,N_2947);
nand U5960 (N_5960,N_874,N_2720);
or U5961 (N_5961,N_28,N_1320);
and U5962 (N_5962,N_1946,N_964);
or U5963 (N_5963,N_1358,N_2016);
or U5964 (N_5964,N_1604,N_371);
nor U5965 (N_5965,N_2392,N_2840);
nand U5966 (N_5966,N_1466,N_1372);
and U5967 (N_5967,N_2325,N_538);
and U5968 (N_5968,N_1128,N_1610);
nand U5969 (N_5969,N_1713,N_2599);
or U5970 (N_5970,N_1693,N_397);
and U5971 (N_5971,N_1471,N_990);
or U5972 (N_5972,N_397,N_2368);
nor U5973 (N_5973,N_1335,N_193);
and U5974 (N_5974,N_2308,N_2709);
nor U5975 (N_5975,N_2435,N_1236);
nand U5976 (N_5976,N_1180,N_2082);
nor U5977 (N_5977,N_1021,N_2715);
and U5978 (N_5978,N_1091,N_539);
or U5979 (N_5979,N_486,N_2605);
nand U5980 (N_5980,N_1843,N_2715);
nor U5981 (N_5981,N_1231,N_2685);
or U5982 (N_5982,N_1975,N_1166);
nor U5983 (N_5983,N_1897,N_137);
and U5984 (N_5984,N_424,N_1003);
nand U5985 (N_5985,N_108,N_2834);
and U5986 (N_5986,N_1569,N_215);
nor U5987 (N_5987,N_2315,N_1660);
nor U5988 (N_5988,N_1631,N_1559);
nor U5989 (N_5989,N_568,N_2276);
nand U5990 (N_5990,N_2307,N_625);
nand U5991 (N_5991,N_1339,N_2064);
nor U5992 (N_5992,N_224,N_301);
nand U5993 (N_5993,N_2261,N_2648);
and U5994 (N_5994,N_608,N_514);
nand U5995 (N_5995,N_2787,N_545);
or U5996 (N_5996,N_469,N_742);
or U5997 (N_5997,N_683,N_2506);
or U5998 (N_5998,N_543,N_2050);
nor U5999 (N_5999,N_1449,N_1545);
or U6000 (N_6000,N_4796,N_5076);
or U6001 (N_6001,N_3456,N_4326);
and U6002 (N_6002,N_4173,N_3061);
and U6003 (N_6003,N_4163,N_3928);
and U6004 (N_6004,N_5832,N_5389);
nand U6005 (N_6005,N_5689,N_5823);
and U6006 (N_6006,N_4878,N_5403);
and U6007 (N_6007,N_4423,N_5635);
nor U6008 (N_6008,N_5856,N_4763);
nand U6009 (N_6009,N_5359,N_4881);
nand U6010 (N_6010,N_3007,N_4202);
and U6011 (N_6011,N_5758,N_4673);
and U6012 (N_6012,N_3398,N_4575);
and U6013 (N_6013,N_5464,N_3245);
nor U6014 (N_6014,N_5813,N_5842);
or U6015 (N_6015,N_4043,N_5791);
nor U6016 (N_6016,N_5433,N_3380);
or U6017 (N_6017,N_3560,N_3680);
or U6018 (N_6018,N_5866,N_4671);
nand U6019 (N_6019,N_3949,N_4375);
and U6020 (N_6020,N_5744,N_4468);
or U6021 (N_6021,N_3073,N_4503);
nor U6022 (N_6022,N_4051,N_3828);
nand U6023 (N_6023,N_5330,N_3113);
nor U6024 (N_6024,N_5849,N_5937);
xor U6025 (N_6025,N_4623,N_3466);
nand U6026 (N_6026,N_5201,N_4061);
nand U6027 (N_6027,N_4121,N_4015);
or U6028 (N_6028,N_5156,N_4209);
or U6029 (N_6029,N_3405,N_4104);
nor U6030 (N_6030,N_5254,N_3299);
nand U6031 (N_6031,N_3208,N_4258);
nand U6032 (N_6032,N_4280,N_5294);
nor U6033 (N_6033,N_4985,N_4789);
nor U6034 (N_6034,N_3328,N_4667);
and U6035 (N_6035,N_4569,N_4198);
nand U6036 (N_6036,N_3078,N_5537);
nor U6037 (N_6037,N_5003,N_4871);
nor U6038 (N_6038,N_4780,N_3538);
nor U6039 (N_6039,N_5134,N_3683);
or U6040 (N_6040,N_4620,N_3576);
nor U6041 (N_6041,N_4894,N_5692);
nor U6042 (N_6042,N_4825,N_4875);
and U6043 (N_6043,N_3451,N_3378);
nand U6044 (N_6044,N_4839,N_3394);
nand U6045 (N_6045,N_3704,N_5239);
nor U6046 (N_6046,N_4688,N_5089);
or U6047 (N_6047,N_3333,N_5595);
nand U6048 (N_6048,N_3728,N_5043);
or U6049 (N_6049,N_3020,N_5863);
and U6050 (N_6050,N_5638,N_3510);
nor U6051 (N_6051,N_3251,N_4382);
nor U6052 (N_6052,N_5442,N_5504);
and U6053 (N_6053,N_3454,N_5923);
or U6054 (N_6054,N_4835,N_4803);
and U6055 (N_6055,N_3998,N_4031);
nor U6056 (N_6056,N_3238,N_5084);
and U6057 (N_6057,N_5615,N_3102);
and U6058 (N_6058,N_4272,N_4800);
nand U6059 (N_6059,N_4231,N_4453);
nand U6060 (N_6060,N_3037,N_5910);
or U6061 (N_6061,N_5404,N_5878);
nand U6062 (N_6062,N_4293,N_5009);
or U6063 (N_6063,N_3977,N_4896);
nor U6064 (N_6064,N_4139,N_5745);
and U6065 (N_6065,N_4256,N_3313);
or U6066 (N_6066,N_3422,N_4903);
nand U6067 (N_6067,N_5341,N_4073);
nor U6068 (N_6068,N_4097,N_4033);
nor U6069 (N_6069,N_5691,N_5492);
nand U6070 (N_6070,N_5713,N_4702);
or U6071 (N_6071,N_5748,N_4837);
and U6072 (N_6072,N_3866,N_4744);
nand U6073 (N_6073,N_5232,N_4479);
and U6074 (N_6074,N_3534,N_5115);
or U6075 (N_6075,N_4373,N_3602);
nor U6076 (N_6076,N_5574,N_5315);
nand U6077 (N_6077,N_5822,N_3529);
and U6078 (N_6078,N_4314,N_4311);
or U6079 (N_6079,N_5209,N_4296);
or U6080 (N_6080,N_5766,N_4217);
or U6081 (N_6081,N_4684,N_3541);
nand U6082 (N_6082,N_4169,N_5977);
or U6083 (N_6083,N_5013,N_3899);
and U6084 (N_6084,N_3823,N_3209);
nand U6085 (N_6085,N_3901,N_5704);
and U6086 (N_6086,N_5533,N_5361);
nand U6087 (N_6087,N_4644,N_4427);
nor U6088 (N_6088,N_4906,N_5186);
or U6089 (N_6089,N_5656,N_4931);
nand U6090 (N_6090,N_4568,N_4670);
and U6091 (N_6091,N_4002,N_5888);
nand U6092 (N_6092,N_5367,N_5346);
xnor U6093 (N_6093,N_4064,N_3980);
and U6094 (N_6094,N_5234,N_5978);
and U6095 (N_6095,N_4579,N_3801);
nor U6096 (N_6096,N_5279,N_3483);
nand U6097 (N_6097,N_3679,N_4443);
and U6098 (N_6098,N_4384,N_3045);
nand U6099 (N_6099,N_5406,N_3648);
nand U6100 (N_6100,N_4257,N_5340);
and U6101 (N_6101,N_5995,N_3411);
and U6102 (N_6102,N_3882,N_4787);
nand U6103 (N_6103,N_5733,N_4666);
or U6104 (N_6104,N_4542,N_3206);
and U6105 (N_6105,N_3614,N_5071);
nand U6106 (N_6106,N_5943,N_3152);
nand U6107 (N_6107,N_5618,N_4084);
nand U6108 (N_6108,N_5235,N_4957);
or U6109 (N_6109,N_5628,N_3668);
nor U6110 (N_6110,N_5883,N_3049);
or U6111 (N_6111,N_4070,N_5461);
or U6112 (N_6112,N_5073,N_4027);
and U6113 (N_6113,N_4678,N_4926);
or U6114 (N_6114,N_3484,N_4607);
nor U6115 (N_6115,N_5962,N_3481);
nor U6116 (N_6116,N_5747,N_4372);
and U6117 (N_6117,N_5990,N_5308);
nor U6118 (N_6118,N_4327,N_4157);
nand U6119 (N_6119,N_5875,N_5731);
and U6120 (N_6120,N_5440,N_4940);
nor U6121 (N_6121,N_3724,N_4393);
nor U6122 (N_6122,N_3262,N_4037);
and U6123 (N_6123,N_3189,N_5019);
nand U6124 (N_6124,N_5070,N_3829);
nand U6125 (N_6125,N_5117,N_3846);
or U6126 (N_6126,N_5011,N_4411);
nor U6127 (N_6127,N_4923,N_3205);
or U6128 (N_6128,N_5954,N_3742);
nand U6129 (N_6129,N_3867,N_4433);
and U6130 (N_6130,N_4227,N_5262);
nand U6131 (N_6131,N_4273,N_5260);
xnor U6132 (N_6132,N_4584,N_5365);
or U6133 (N_6133,N_4741,N_5735);
and U6134 (N_6134,N_5229,N_5032);
xnor U6135 (N_6135,N_3825,N_3270);
nand U6136 (N_6136,N_5217,N_3107);
and U6137 (N_6137,N_4442,N_3835);
and U6138 (N_6138,N_3219,N_5306);
nor U6139 (N_6139,N_3459,N_4737);
or U6140 (N_6140,N_3369,N_5782);
or U6141 (N_6141,N_3229,N_4193);
nor U6142 (N_6142,N_4981,N_5455);
nand U6143 (N_6143,N_4880,N_5933);
and U6144 (N_6144,N_5049,N_4485);
nor U6145 (N_6145,N_5899,N_4040);
nand U6146 (N_6146,N_4358,N_3243);
nor U6147 (N_6147,N_4378,N_3851);
or U6148 (N_6148,N_4762,N_5776);
and U6149 (N_6149,N_3293,N_3282);
nor U6150 (N_6150,N_5012,N_5028);
nand U6151 (N_6151,N_5203,N_4580);
and U6152 (N_6152,N_4392,N_4545);
and U6153 (N_6153,N_3730,N_3936);
nor U6154 (N_6154,N_4840,N_4802);
nand U6155 (N_6155,N_5793,N_4638);
and U6156 (N_6156,N_5489,N_3120);
and U6157 (N_6157,N_3160,N_4298);
and U6158 (N_6158,N_5318,N_4813);
nand U6159 (N_6159,N_3403,N_5624);
nand U6160 (N_6160,N_3666,N_3550);
or U6161 (N_6161,N_5123,N_3464);
and U6162 (N_6162,N_3275,N_5792);
nand U6163 (N_6163,N_4264,N_5021);
nor U6164 (N_6164,N_3496,N_4980);
and U6165 (N_6165,N_5268,N_3091);
nor U6166 (N_6166,N_4548,N_3859);
or U6167 (N_6167,N_3144,N_3253);
nand U6168 (N_6168,N_5802,N_3324);
or U6169 (N_6169,N_4654,N_4941);
and U6170 (N_6170,N_4549,N_5577);
and U6171 (N_6171,N_3658,N_3857);
nor U6172 (N_6172,N_3645,N_4420);
and U6173 (N_6173,N_5042,N_3840);
nor U6174 (N_6174,N_3134,N_3771);
nand U6175 (N_6175,N_5351,N_5121);
nand U6176 (N_6176,N_5760,N_4480);
or U6177 (N_6177,N_4275,N_3927);
nand U6178 (N_6178,N_5771,N_4228);
or U6179 (N_6179,N_5145,N_3590);
nand U6180 (N_6180,N_3697,N_4005);
nor U6181 (N_6181,N_4446,N_3312);
nand U6182 (N_6182,N_4165,N_5007);
nand U6183 (N_6183,N_4464,N_4860);
nand U6184 (N_6184,N_3086,N_3636);
and U6185 (N_6185,N_4074,N_5027);
and U6186 (N_6186,N_4016,N_3438);
nand U6187 (N_6187,N_4619,N_4270);
nand U6188 (N_6188,N_4652,N_4947);
nand U6189 (N_6189,N_5512,N_3946);
nor U6190 (N_6190,N_3997,N_4733);
nand U6191 (N_6191,N_4476,N_3470);
or U6192 (N_6192,N_3213,N_4588);
nor U6193 (N_6193,N_5085,N_3446);
or U6194 (N_6194,N_3995,N_4754);
and U6195 (N_6195,N_4412,N_5321);
nand U6196 (N_6196,N_3480,N_4036);
and U6197 (N_6197,N_5449,N_4204);
and U6198 (N_6198,N_5467,N_3616);
nor U6199 (N_6199,N_4137,N_4492);
nor U6200 (N_6200,N_3729,N_4861);
nor U6201 (N_6201,N_3501,N_5852);
nand U6202 (N_6202,N_5197,N_5329);
or U6203 (N_6203,N_4429,N_4328);
or U6204 (N_6204,N_3316,N_3231);
nor U6205 (N_6205,N_3630,N_4434);
nor U6206 (N_6206,N_3407,N_4351);
and U6207 (N_6207,N_3522,N_3844);
xnor U6208 (N_6208,N_3286,N_3611);
nand U6209 (N_6209,N_3563,N_5907);
and U6210 (N_6210,N_3987,N_5999);
nor U6211 (N_6211,N_5081,N_3039);
or U6212 (N_6212,N_4366,N_5569);
xnor U6213 (N_6213,N_5687,N_4971);
and U6214 (N_6214,N_4630,N_4919);
nor U6215 (N_6215,N_4783,N_5526);
and U6216 (N_6216,N_3311,N_3461);
and U6217 (N_6217,N_5958,N_3352);
and U6218 (N_6218,N_5447,N_3399);
nand U6219 (N_6219,N_5041,N_5746);
nor U6220 (N_6220,N_4007,N_5607);
nor U6221 (N_6221,N_4844,N_3767);
and U6222 (N_6222,N_4451,N_5617);
nand U6223 (N_6223,N_3338,N_3922);
nor U6224 (N_6224,N_5546,N_3148);
and U6225 (N_6225,N_5106,N_3214);
nor U6226 (N_6226,N_5700,N_5036);
or U6227 (N_6227,N_5398,N_3706);
or U6228 (N_6228,N_3237,N_4624);
nand U6229 (N_6229,N_4409,N_5188);
nor U6230 (N_6230,N_4085,N_3890);
or U6231 (N_6231,N_3332,N_3824);
nor U6232 (N_6232,N_4959,N_4723);
and U6233 (N_6233,N_4238,N_5720);
nand U6234 (N_6234,N_3942,N_3548);
and U6235 (N_6235,N_3633,N_4938);
and U6236 (N_6236,N_3334,N_5238);
or U6237 (N_6237,N_3693,N_4457);
and U6238 (N_6238,N_5065,N_5418);
and U6239 (N_6239,N_3048,N_5103);
or U6240 (N_6240,N_4136,N_3717);
nor U6241 (N_6241,N_3800,N_5989);
nand U6242 (N_6242,N_4533,N_3878);
nor U6243 (N_6243,N_5290,N_5901);
nor U6244 (N_6244,N_4658,N_3121);
or U6245 (N_6245,N_3701,N_3958);
or U6246 (N_6246,N_4912,N_5307);
nand U6247 (N_6247,N_5947,N_5696);
nor U6248 (N_6248,N_3079,N_5383);
or U6249 (N_6249,N_3832,N_5069);
nor U6250 (N_6250,N_4415,N_4738);
nand U6251 (N_6251,N_3123,N_4215);
or U6252 (N_6252,N_5592,N_3010);
and U6253 (N_6253,N_5818,N_3343);
nor U6254 (N_6254,N_3386,N_5803);
and U6255 (N_6255,N_3181,N_4025);
and U6256 (N_6256,N_5267,N_3695);
nand U6257 (N_6257,N_3241,N_5566);
nand U6258 (N_6258,N_3687,N_4312);
or U6259 (N_6259,N_4368,N_5718);
or U6260 (N_6260,N_3468,N_4347);
nor U6261 (N_6261,N_5285,N_3193);
or U6262 (N_6262,N_4076,N_5814);
nor U6263 (N_6263,N_5547,N_5474);
or U6264 (N_6264,N_3607,N_4720);
and U6265 (N_6265,N_4179,N_3439);
and U6266 (N_6266,N_3774,N_5044);
or U6267 (N_6267,N_3690,N_5006);
nand U6268 (N_6268,N_4172,N_4018);
or U6269 (N_6269,N_3793,N_4521);
nand U6270 (N_6270,N_3361,N_4657);
nor U6271 (N_6271,N_5396,N_4963);
nor U6272 (N_6272,N_5596,N_3240);
and U6273 (N_6273,N_4161,N_5709);
nor U6274 (N_6274,N_3856,N_5850);
and U6275 (N_6275,N_4029,N_3082);
and U6276 (N_6276,N_4817,N_3650);
and U6277 (N_6277,N_5819,N_5921);
nand U6278 (N_6278,N_4124,N_4331);
and U6279 (N_6279,N_4700,N_4340);
nor U6280 (N_6280,N_3902,N_4487);
and U6281 (N_6281,N_4413,N_3167);
nand U6282 (N_6282,N_5353,N_4822);
nor U6283 (N_6283,N_4252,N_4973);
or U6284 (N_6284,N_5038,N_5453);
or U6285 (N_6285,N_3390,N_3106);
or U6286 (N_6286,N_3430,N_4180);
nand U6287 (N_6287,N_4035,N_4364);
and U6288 (N_6288,N_5171,N_5892);
nand U6289 (N_6289,N_3178,N_3002);
nand U6290 (N_6290,N_3285,N_4782);
nand U6291 (N_6291,N_3132,N_3659);
and U6292 (N_6292,N_4633,N_4911);
or U6293 (N_6293,N_5797,N_3551);
nor U6294 (N_6294,N_5862,N_5130);
nand U6295 (N_6295,N_3268,N_3447);
and U6296 (N_6296,N_3626,N_4815);
and U6297 (N_6297,N_3104,N_4463);
and U6298 (N_6298,N_4742,N_3649);
or U6299 (N_6299,N_4461,N_4904);
nor U6300 (N_6300,N_4523,N_5451);
and U6301 (N_6301,N_5193,N_3184);
or U6302 (N_6302,N_3696,N_4602);
nand U6303 (N_6303,N_5488,N_5435);
and U6304 (N_6304,N_5939,N_4297);
or U6305 (N_6305,N_4722,N_3008);
nand U6306 (N_6306,N_5487,N_3580);
or U6307 (N_6307,N_3096,N_4982);
or U6308 (N_6308,N_3939,N_3067);
or U6309 (N_6309,N_5362,N_3723);
nor U6310 (N_6310,N_3026,N_4019);
nand U6311 (N_6311,N_3495,N_4539);
or U6312 (N_6312,N_4555,N_4646);
nand U6313 (N_6313,N_3564,N_4788);
or U6314 (N_6314,N_5559,N_5909);
nand U6315 (N_6315,N_5919,N_3678);
or U6316 (N_6316,N_3689,N_3246);
nor U6317 (N_6317,N_5491,N_4887);
or U6318 (N_6318,N_4761,N_5142);
and U6319 (N_6319,N_4240,N_3596);
or U6320 (N_6320,N_5183,N_4529);
and U6321 (N_6321,N_5839,N_5018);
nand U6322 (N_6322,N_5111,N_3609);
and U6323 (N_6323,N_5774,N_5015);
or U6324 (N_6324,N_5247,N_3926);
nor U6325 (N_6325,N_3013,N_3040);
or U6326 (N_6326,N_4997,N_4417);
nand U6327 (N_6327,N_5622,N_4099);
or U6328 (N_6328,N_4160,N_3852);
and U6329 (N_6329,N_3457,N_5975);
nor U6330 (N_6330,N_3671,N_5683);
nor U6331 (N_6331,N_5258,N_5244);
nor U6332 (N_6332,N_5931,N_5213);
nor U6333 (N_6333,N_4512,N_3103);
and U6334 (N_6334,N_3250,N_5326);
or U6335 (N_6335,N_5784,N_3440);
and U6336 (N_6336,N_5506,N_4914);
and U6337 (N_6337,N_3960,N_4632);
nand U6338 (N_6338,N_4901,N_5058);
nor U6339 (N_6339,N_4816,N_5332);
nand U6340 (N_6340,N_5633,N_5997);
nand U6341 (N_6341,N_3727,N_3874);
nand U6342 (N_6342,N_5529,N_3076);
nand U6343 (N_6343,N_3778,N_4484);
and U6344 (N_6344,N_4544,N_3733);
or U6345 (N_6345,N_3119,N_3546);
nand U6346 (N_6346,N_3883,N_3570);
and U6347 (N_6347,N_4534,N_4301);
and U6348 (N_6348,N_4677,N_4642);
or U6349 (N_6349,N_4462,N_5681);
nand U6350 (N_6350,N_4026,N_5705);
or U6351 (N_6351,N_4060,N_3218);
nand U6352 (N_6352,N_3383,N_5988);
nor U6353 (N_6353,N_3269,N_3164);
or U6354 (N_6354,N_5490,N_4474);
nor U6355 (N_6355,N_3544,N_5684);
or U6356 (N_6356,N_5973,N_3223);
or U6357 (N_6357,N_3631,N_4907);
nor U6358 (N_6358,N_3613,N_5528);
nor U6359 (N_6359,N_5558,N_5916);
xor U6360 (N_6360,N_3937,N_5462);
xnor U6361 (N_6361,N_4426,N_5377);
and U6362 (N_6362,N_5154,N_4984);
nor U6363 (N_6363,N_5889,N_3819);
and U6364 (N_6364,N_5310,N_4224);
nand U6365 (N_6365,N_3101,N_4406);
nor U6366 (N_6366,N_3996,N_3493);
or U6367 (N_6367,N_3153,N_4247);
or U6368 (N_6368,N_3034,N_4158);
nand U6369 (N_6369,N_4481,N_5945);
nor U6370 (N_6370,N_5532,N_5804);
nand U6371 (N_6371,N_4653,N_4396);
or U6372 (N_6372,N_4318,N_4955);
and U6373 (N_6373,N_4236,N_3620);
and U6374 (N_6374,N_3978,N_5345);
nor U6375 (N_6375,N_4701,N_3331);
or U6376 (N_6376,N_3281,N_3228);
or U6377 (N_6377,N_4313,N_3809);
or U6378 (N_6378,N_5296,N_5620);
and U6379 (N_6379,N_4853,N_5328);
and U6380 (N_6380,N_3089,N_5877);
nor U6381 (N_6381,N_5903,N_3940);
nand U6382 (N_6382,N_4905,N_5074);
and U6383 (N_6383,N_5757,N_3477);
nor U6384 (N_6384,N_3449,N_4974);
nand U6385 (N_6385,N_4552,N_4553);
nand U6386 (N_6386,N_3363,N_4316);
or U6387 (N_6387,N_5717,N_3950);
nor U6388 (N_6388,N_5360,N_4972);
and U6389 (N_6389,N_4942,N_5458);
and U6390 (N_6390,N_3804,N_3612);
or U6391 (N_6391,N_5116,N_3431);
nand U6392 (N_6392,N_4759,N_3655);
nor U6393 (N_6393,N_3872,N_5680);
nand U6394 (N_6394,N_5348,N_3325);
and U6395 (N_6395,N_3017,N_5048);
nor U6396 (N_6396,N_4626,N_5544);
nand U6397 (N_6397,N_4801,N_5865);
and U6398 (N_6398,N_5140,N_3349);
nor U6399 (N_6399,N_4819,N_5192);
nor U6400 (N_6400,N_4609,N_4363);
nand U6401 (N_6401,N_3179,N_3058);
nand U6402 (N_6402,N_3256,N_4181);
and U6403 (N_6403,N_4572,N_4081);
or U6404 (N_6404,N_5579,N_4961);
and U6405 (N_6405,N_5429,N_3276);
nor U6406 (N_6406,N_5194,N_4122);
nand U6407 (N_6407,N_5535,N_3307);
nor U6408 (N_6408,N_3122,N_4842);
or U6409 (N_6409,N_5198,N_4836);
or U6410 (N_6410,N_5205,N_4034);
nand U6411 (N_6411,N_3216,N_5690);
or U6412 (N_6412,N_3662,N_5493);
nor U6413 (N_6413,N_3267,N_4459);
nor U6414 (N_6414,N_5721,N_5059);
and U6415 (N_6415,N_4159,N_5957);
nand U6416 (N_6416,N_5556,N_4556);
nor U6417 (N_6417,N_3956,N_5052);
nand U6418 (N_6418,N_4593,N_5664);
nand U6419 (N_6419,N_4192,N_3083);
and U6420 (N_6420,N_4115,N_4937);
nor U6421 (N_6421,N_5466,N_5930);
nand U6422 (N_6422,N_5867,N_5327);
and U6423 (N_6423,N_4987,N_3948);
and U6424 (N_6424,N_3195,N_4715);
or U6425 (N_6425,N_5510,N_4319);
nor U6426 (N_6426,N_5502,N_3173);
and U6427 (N_6427,N_5926,N_4407);
nor U6428 (N_6428,N_4200,N_3854);
and U6429 (N_6429,N_5716,N_5181);
nand U6430 (N_6430,N_5151,N_3156);
nand U6431 (N_6431,N_3552,N_3302);
nand U6432 (N_6432,N_4932,N_5093);
and U6433 (N_6433,N_4248,N_3317);
nor U6434 (N_6434,N_4149,N_4517);
and U6435 (N_6435,N_4403,N_5825);
nand U6436 (N_6436,N_3041,N_3663);
or U6437 (N_6437,N_5165,N_4354);
nand U6438 (N_6438,N_5851,N_3578);
nand U6439 (N_6439,N_5987,N_5104);
nand U6440 (N_6440,N_3395,N_4329);
nand U6441 (N_6441,N_3808,N_4691);
and U6442 (N_6442,N_5414,N_4105);
and U6443 (N_6443,N_5379,N_5139);
nand U6444 (N_6444,N_5563,N_5114);
or U6445 (N_6445,N_4511,N_4376);
nor U6446 (N_6446,N_4551,N_4869);
nand U6447 (N_6447,N_3756,N_5612);
nand U6448 (N_6448,N_4683,N_5484);
nor U6449 (N_6449,N_3441,N_3681);
nor U6450 (N_6450,N_3192,N_3722);
nor U6451 (N_6451,N_5756,N_5739);
nand U6452 (N_6452,N_3358,N_3657);
nor U6453 (N_6453,N_5788,N_3515);
nor U6454 (N_6454,N_3374,N_3935);
nor U6455 (N_6455,N_5179,N_3029);
nor U6456 (N_6456,N_4879,N_4205);
nand U6457 (N_6457,N_3537,N_3549);
or U6458 (N_6458,N_5463,N_5266);
nand U6459 (N_6459,N_4402,N_3907);
and U6460 (N_6460,N_5800,N_4970);
and U6461 (N_6461,N_5854,N_3095);
or U6462 (N_6462,N_5241,N_3341);
xor U6463 (N_6463,N_3056,N_5356);
or U6464 (N_6464,N_4466,N_5108);
and U6465 (N_6465,N_5831,N_5645);
xor U6466 (N_6466,N_3992,N_4108);
nor U6467 (N_6467,N_4703,N_5913);
nor U6468 (N_6468,N_3309,N_3221);
xor U6469 (N_6469,N_4739,N_3779);
and U6470 (N_6470,N_4611,N_5347);
and U6471 (N_6471,N_5523,N_5388);
or U6472 (N_6472,N_3188,N_5162);
and U6473 (N_6473,N_5411,N_5163);
and U6474 (N_6474,N_3210,N_5561);
and U6475 (N_6475,N_4855,N_5001);
and U6476 (N_6476,N_5698,N_4438);
and U6477 (N_6477,N_4381,N_5643);
or U6478 (N_6478,N_5815,N_5299);
and U6479 (N_6479,N_5441,N_5672);
or U6480 (N_6480,N_3572,N_3985);
nor U6481 (N_6481,N_3865,N_4645);
nand U6482 (N_6482,N_5855,N_5940);
nor U6483 (N_6483,N_4501,N_5068);
and U6484 (N_6484,N_3777,N_4212);
nand U6485 (N_6485,N_5562,N_4877);
or U6486 (N_6486,N_5657,N_3085);
or U6487 (N_6487,N_4705,N_3743);
or U6488 (N_6488,N_5964,N_5702);
nor U6489 (N_6489,N_3861,N_5251);
and U6490 (N_6490,N_4008,N_4864);
nor U6491 (N_6491,N_3402,N_4920);
and U6492 (N_6492,N_4057,N_3226);
and U6493 (N_6493,N_5083,N_3090);
nand U6494 (N_6494,N_5090,N_5991);
nor U6495 (N_6495,N_3488,N_5986);
nand U6496 (N_6496,N_3732,N_3360);
and U6497 (N_6497,N_5184,N_3877);
and U6498 (N_6498,N_3478,N_4820);
nor U6499 (N_6499,N_3962,N_3752);
nor U6500 (N_6500,N_3025,N_4194);
and U6501 (N_6501,N_3543,N_3860);
or U6502 (N_6502,N_5334,N_5298);
nand U6503 (N_6503,N_3437,N_3532);
and U6504 (N_6504,N_4253,N_5591);
nor U6505 (N_6505,N_3344,N_3052);
nor U6506 (N_6506,N_3465,N_5868);
and U6507 (N_6507,N_4708,N_4475);
nor U6508 (N_6508,N_5611,N_4740);
nand U6509 (N_6509,N_4473,N_4509);
or U6510 (N_6510,N_4718,N_4103);
nand U6511 (N_6511,N_4142,N_3869);
nor U6512 (N_6512,N_4148,N_3897);
nor U6513 (N_6513,N_4053,N_3589);
and U6514 (N_6514,N_4478,N_4989);
nor U6515 (N_6515,N_5175,N_5799);
nand U6516 (N_6516,N_5876,N_4766);
nor U6517 (N_6517,N_4325,N_3975);
nand U6518 (N_6518,N_3610,N_5589);
or U6519 (N_6519,N_5270,N_4261);
nor U6520 (N_6520,N_5764,N_3426);
nor U6521 (N_6521,N_4141,N_4929);
nand U6522 (N_6522,N_3896,N_4858);
and U6523 (N_6523,N_3716,N_4006);
nor U6524 (N_6524,N_4041,N_3116);
nor U6525 (N_6525,N_3366,N_4092);
and U6526 (N_6526,N_5509,N_4456);
and U6527 (N_6527,N_5801,N_3763);
nor U6528 (N_6528,N_3919,N_4799);
or U6529 (N_6529,N_4730,N_5312);
nand U6530 (N_6530,N_5037,N_3517);
and U6531 (N_6531,N_5917,N_5159);
nand U6532 (N_6532,N_3619,N_3700);
nand U6533 (N_6533,N_4388,N_3904);
nand U6534 (N_6534,N_5723,N_5654);
nor U6535 (N_6535,N_5166,N_5333);
and U6536 (N_6536,N_5372,N_4093);
nand U6537 (N_6537,N_4591,N_5750);
nor U6538 (N_6538,N_5167,N_5873);
nand U6539 (N_6539,N_5086,N_5264);
nand U6540 (N_6540,N_5751,N_5160);
or U6541 (N_6541,N_4221,N_3617);
nor U6542 (N_6542,N_4682,N_4687);
nand U6543 (N_6543,N_4095,N_5082);
or U6544 (N_6544,N_3345,N_4967);
and U6545 (N_6545,N_3947,N_5824);
and U6546 (N_6546,N_5407,N_5176);
nor U6547 (N_6547,N_4174,N_4828);
and U6548 (N_6548,N_5539,N_3014);
and U6549 (N_6549,N_4599,N_5550);
or U6550 (N_6550,N_5230,N_5056);
nand U6551 (N_6551,N_5714,N_4606);
or U6552 (N_6552,N_5830,N_4774);
and U6553 (N_6553,N_4757,N_5099);
nand U6554 (N_6554,N_3232,N_4806);
nor U6555 (N_6555,N_3044,N_3559);
or U6556 (N_6556,N_5548,N_4353);
or U6557 (N_6557,N_5412,N_4399);
nor U6558 (N_6558,N_5033,N_5152);
nor U6559 (N_6559,N_5382,N_3295);
or U6560 (N_6560,N_3858,N_4047);
and U6561 (N_6561,N_4953,N_3442);
or U6562 (N_6562,N_5786,N_3539);
nand U6563 (N_6563,N_3755,N_3908);
nand U6564 (N_6564,N_5051,N_4385);
nor U6565 (N_6565,N_3817,N_3423);
or U6566 (N_6566,N_4899,N_3051);
and U6567 (N_6567,N_5514,N_4917);
and U6568 (N_6568,N_3761,N_3301);
or U6569 (N_6569,N_3964,N_5811);
or U6570 (N_6570,N_3400,N_5105);
or U6571 (N_6571,N_3359,N_4362);
nand U6572 (N_6572,N_3200,N_5726);
or U6573 (N_6573,N_4419,N_4335);
and U6574 (N_6574,N_5588,N_3419);
and U6575 (N_6575,N_4023,N_4884);
or U6576 (N_6576,N_5400,N_3837);
or U6577 (N_6577,N_5606,N_4531);
or U6578 (N_6578,N_5295,N_4935);
nor U6579 (N_6579,N_4400,N_5661);
nor U6580 (N_6580,N_3601,N_4255);
or U6581 (N_6581,N_5906,N_4731);
and U6582 (N_6582,N_3350,N_4144);
nor U6583 (N_6583,N_4190,N_3989);
or U6584 (N_6584,N_3435,N_4751);
or U6585 (N_6585,N_4681,N_4470);
or U6586 (N_6586,N_3768,N_4243);
nand U6587 (N_6587,N_3796,N_4250);
nand U6588 (N_6588,N_4927,N_3081);
or U6589 (N_6589,N_5951,N_4440);
nand U6590 (N_6590,N_4483,N_4567);
nor U6591 (N_6591,N_4488,N_3003);
nor U6592 (N_6592,N_5730,N_5675);
or U6593 (N_6593,N_3236,N_5828);
and U6594 (N_6594,N_5250,N_5237);
nor U6595 (N_6595,N_3158,N_5971);
nor U6596 (N_6596,N_5337,N_3445);
nand U6597 (N_6597,N_4303,N_5838);
nand U6598 (N_6598,N_3664,N_5132);
nand U6599 (N_6599,N_4746,N_4793);
and U6600 (N_6600,N_4686,N_3892);
and U6601 (N_6601,N_3023,N_3673);
nor U6602 (N_6602,N_5158,N_5670);
or U6603 (N_6603,N_3795,N_5317);
and U6604 (N_6604,N_3586,N_3077);
nor U6605 (N_6605,N_5642,N_4797);
xnor U6606 (N_6606,N_5604,N_4398);
or U6607 (N_6607,N_3565,N_3581);
or U6608 (N_6608,N_5541,N_4647);
or U6609 (N_6609,N_5438,N_4379);
nand U6610 (N_6610,N_3384,N_4581);
nand U6611 (N_6611,N_3963,N_3409);
nor U6612 (N_6612,N_4009,N_4753);
or U6613 (N_6613,N_4656,N_5941);
nand U6614 (N_6614,N_3688,N_4226);
nor U6615 (N_6615,N_4486,N_5527);
and U6616 (N_6616,N_5820,N_4156);
nand U6617 (N_6617,N_4333,N_5202);
or U6618 (N_6618,N_5715,N_5240);
or U6619 (N_6619,N_4535,N_5685);
nand U6620 (N_6620,N_4222,N_4305);
nand U6621 (N_6621,N_3207,N_3233);
and U6622 (N_6622,N_5665,N_4775);
or U6623 (N_6623,N_4153,N_3595);
nand U6624 (N_6624,N_3830,N_3059);
nand U6625 (N_6625,N_4482,N_5062);
and U6626 (N_6626,N_4850,N_5511);
and U6627 (N_6627,N_5603,N_4214);
nor U6628 (N_6628,N_3932,N_4514);
nand U6629 (N_6629,N_5350,N_5014);
and U6630 (N_6630,N_3615,N_4900);
and U6631 (N_6631,N_4622,N_4617);
nand U6632 (N_6632,N_3053,N_5630);
nor U6633 (N_6633,N_3455,N_3863);
and U6634 (N_6634,N_3162,N_5335);
nor U6635 (N_6635,N_3976,N_5965);
or U6636 (N_6636,N_3929,N_4713);
nand U6637 (N_6637,N_4726,N_5272);
or U6638 (N_6638,N_3355,N_3163);
nand U6639 (N_6639,N_4283,N_4206);
nor U6640 (N_6640,N_5276,N_5182);
or U6641 (N_6641,N_4563,N_4045);
or U6642 (N_6642,N_3781,N_3462);
or U6643 (N_6643,N_4504,N_3117);
nor U6644 (N_6644,N_5884,N_3127);
nor U6645 (N_6645,N_3748,N_3306);
and U6646 (N_6646,N_5273,N_5749);
and U6647 (N_6647,N_4675,N_4120);
nor U6648 (N_6648,N_3911,N_3672);
nand U6649 (N_6649,N_4066,N_5196);
nand U6650 (N_6650,N_4958,N_4665);
nor U6651 (N_6651,N_3087,N_4263);
nor U6652 (N_6652,N_3850,N_5499);
nand U6653 (N_6653,N_4489,N_5844);
or U6654 (N_6654,N_4830,N_5495);
or U6655 (N_6655,N_4674,N_3110);
or U6656 (N_6656,N_5707,N_4125);
and U6657 (N_6657,N_5513,N_4999);
nor U6658 (N_6658,N_5742,N_5439);
nor U6659 (N_6659,N_3272,N_5732);
nand U6660 (N_6660,N_4201,N_5778);
xnor U6661 (N_6661,N_3050,N_3146);
nor U6662 (N_6662,N_3821,N_3953);
nand U6663 (N_6663,N_5236,N_5399);
nor U6664 (N_6664,N_3006,N_3257);
or U6665 (N_6665,N_3217,N_5682);
or U6666 (N_6666,N_4164,N_3557);
or U6667 (N_6667,N_5172,N_3469);
nor U6668 (N_6668,N_4930,N_4507);
or U6669 (N_6669,N_4621,N_4211);
or U6670 (N_6670,N_3739,N_5845);
nor U6671 (N_6671,N_5384,N_3784);
and U6672 (N_6672,N_5605,N_5039);
or U6673 (N_6673,N_3691,N_5391);
or U6674 (N_6674,N_4177,N_3737);
nor U6675 (N_6675,N_4265,N_5826);
nor U6676 (N_6676,N_3443,N_4976);
xnor U6677 (N_6677,N_5816,N_4435);
nor U6678 (N_6678,N_5996,N_4251);
nand U6679 (N_6679,N_4138,N_4990);
or U6680 (N_6680,N_4873,N_5998);
or U6681 (N_6681,N_4515,N_4809);
nor U6682 (N_6682,N_5770,N_3347);
nor U6683 (N_6683,N_4516,N_4676);
or U6684 (N_6684,N_3849,N_4166);
and U6685 (N_6685,N_3972,N_3244);
and U6686 (N_6686,N_5064,N_5521);
and U6687 (N_6687,N_5787,N_3027);
and U6688 (N_6688,N_3864,N_3647);
nand U6689 (N_6689,N_4395,N_4867);
nor U6690 (N_6690,N_3898,N_3838);
nor U6691 (N_6691,N_3322,N_5741);
or U6692 (N_6692,N_4784,N_5835);
nand U6693 (N_6693,N_4791,N_5078);
nor U6694 (N_6694,N_3624,N_3893);
and U6695 (N_6695,N_4497,N_4964);
or U6696 (N_6696,N_5695,N_3487);
or U6697 (N_6697,N_5402,N_3393);
nor U6698 (N_6698,N_3004,N_5436);
and U6699 (N_6699,N_5291,N_5821);
or U6700 (N_6700,N_5555,N_4826);
and U6701 (N_6701,N_3062,N_4949);
nand U6702 (N_6702,N_3661,N_3310);
nand U6703 (N_6703,N_3562,N_3174);
or U6704 (N_6704,N_4596,N_3249);
or U6705 (N_6705,N_3915,N_3785);
and U6706 (N_6706,N_5583,N_3147);
nand U6707 (N_6707,N_3554,N_3124);
nor U6708 (N_6708,N_3891,N_5316);
and U6709 (N_6709,N_4203,N_3097);
or U6710 (N_6710,N_4133,N_3749);
or U6711 (N_6711,N_5869,N_3711);
and U6712 (N_6712,N_4721,N_3802);
nand U6713 (N_6713,N_5572,N_4010);
or U6714 (N_6714,N_4336,N_5128);
nand U6715 (N_6715,N_5754,N_5452);
nor U6716 (N_6716,N_3263,N_5497);
nor U6717 (N_6717,N_3497,N_3308);
nor U6718 (N_6718,N_3064,N_3396);
and U6719 (N_6719,N_3660,N_3379);
and U6720 (N_6720,N_3186,N_5891);
and U6721 (N_6721,N_4425,N_4234);
nor U6722 (N_6722,N_5180,N_3284);
nand U6723 (N_6723,N_3641,N_4281);
nor U6724 (N_6724,N_5627,N_5631);
nand U6725 (N_6725,N_4641,N_3018);
nor U6726 (N_6726,N_4979,N_4557);
nor U6727 (N_6727,N_5199,N_3587);
or U6728 (N_6728,N_4526,N_5538);
xor U6729 (N_6729,N_4056,N_3265);
xor U6730 (N_6730,N_3212,N_4380);
or U6731 (N_6731,N_5531,N_3786);
nor U6732 (N_6732,N_3621,N_4892);
nand U6733 (N_6733,N_5177,N_5421);
or U6734 (N_6734,N_3508,N_4028);
or U6735 (N_6735,N_4547,N_3458);
or U6736 (N_6736,N_3412,N_3471);
nand U6737 (N_6737,N_4893,N_3862);
or U6738 (N_6738,N_5543,N_4594);
nor U6739 (N_6739,N_5623,N_3415);
and U6740 (N_6740,N_5161,N_5055);
or U6741 (N_6741,N_4274,N_4260);
and U6742 (N_6742,N_3606,N_4151);
or U6743 (N_6743,N_5843,N_4096);
or U6744 (N_6744,N_5560,N_3764);
or U6745 (N_6745,N_5805,N_4859);
and U6746 (N_6746,N_5434,N_5375);
nor U6747 (N_6747,N_4285,N_5922);
or U6748 (N_6748,N_5753,N_4934);
nand U6749 (N_6749,N_3075,N_4162);
and U6750 (N_6750,N_4945,N_4129);
and U6751 (N_6751,N_3420,N_4242);
and U6752 (N_6752,N_5323,N_3151);
nor U6753 (N_6753,N_4760,N_5113);
or U6754 (N_6754,N_5966,N_4614);
or U6755 (N_6755,N_3599,N_3414);
nand U6756 (N_6756,N_4321,N_4356);
nor U6757 (N_6757,N_5381,N_5143);
nor U6758 (N_6758,N_5545,N_4128);
nor U6759 (N_6759,N_5405,N_4528);
nand U6760 (N_6760,N_3329,N_3182);
and U6761 (N_6761,N_5676,N_4833);
nor U6762 (N_6762,N_5061,N_5067);
nor U6763 (N_6763,N_5515,N_5077);
nand U6764 (N_6764,N_4794,N_5080);
nor U6765 (N_6765,N_5257,N_4237);
nand U6766 (N_6766,N_3637,N_5568);
nand U6767 (N_6767,N_5729,N_3099);
or U6768 (N_6768,N_5500,N_3714);
or U6769 (N_6769,N_4432,N_4155);
nor U6770 (N_6770,N_3137,N_4882);
or U6771 (N_6771,N_3813,N_4745);
or U6772 (N_6772,N_3521,N_3071);
and U6773 (N_6773,N_4662,N_3734);
nor U6774 (N_6774,N_3568,N_5578);
nor U6775 (N_6775,N_5302,N_3503);
and U6776 (N_6776,N_3642,N_5893);
and U6777 (N_6777,N_4452,N_3993);
and U6778 (N_6778,N_3881,N_5185);
nand U6779 (N_6779,N_5666,N_3833);
nand U6780 (N_6780,N_5710,N_3981);
and U6781 (N_6781,N_3142,N_5669);
and U6782 (N_6782,N_4928,N_5355);
and U6783 (N_6783,N_5319,N_4712);
or U6784 (N_6784,N_4350,N_3588);
nor U6785 (N_6785,N_5428,N_5417);
nand U6786 (N_6786,N_3305,N_5075);
or U6787 (N_6787,N_4170,N_4779);
nor U6788 (N_6788,N_4527,N_5129);
nor U6789 (N_6789,N_4262,N_5373);
and U6790 (N_6790,N_4001,N_5779);
and U6791 (N_6791,N_3959,N_4991);
nor U6792 (N_6792,N_3154,N_3166);
and U6793 (N_6793,N_5894,N_5023);
and U6794 (N_6794,N_5107,N_5525);
nand U6795 (N_6795,N_3703,N_4123);
or U6796 (N_6796,N_5005,N_5840);
and U6797 (N_6797,N_5518,N_5390);
nor U6798 (N_6798,N_3482,N_5227);
or U6799 (N_6799,N_4088,N_4213);
and U6800 (N_6800,N_5678,N_5206);
or U6801 (N_6801,N_3747,N_3060);
nand U6802 (N_6802,N_4334,N_3632);
or U6803 (N_6803,N_3791,N_4054);
and U6804 (N_6804,N_3628,N_3841);
and U6805 (N_6805,N_3925,N_5047);
and U6806 (N_6806,N_5287,N_5226);
xnor U6807 (N_6807,N_5246,N_3479);
nor U6808 (N_6808,N_5915,N_5609);
and U6809 (N_6809,N_4918,N_4966);
and U6810 (N_6810,N_3931,N_3171);
nor U6811 (N_6811,N_4289,N_3001);
nor U6812 (N_6812,N_3063,N_3968);
or U6813 (N_6813,N_3012,N_4277);
nand U6814 (N_6814,N_5616,N_5008);
nor U6815 (N_6815,N_3165,N_5289);
and U6816 (N_6816,N_4246,N_3201);
or U6817 (N_6817,N_3485,N_5137);
or U6818 (N_6818,N_3070,N_5660);
nor U6819 (N_6819,N_4808,N_4598);
or U6820 (N_6820,N_4304,N_5444);
or U6821 (N_6821,N_3842,N_4369);
nand U6822 (N_6822,N_5636,N_4939);
nand U6823 (N_6823,N_4562,N_4341);
nand U6824 (N_6824,N_3354,N_4448);
and U6825 (N_6825,N_4307,N_5415);
nor U6826 (N_6826,N_4807,N_5035);
or U6827 (N_6827,N_3561,N_4943);
nand U6828 (N_6828,N_3365,N_4902);
and U6829 (N_6829,N_4725,N_3128);
and U6830 (N_6830,N_4592,N_4225);
nor U6831 (N_6831,N_3816,N_4437);
and U6832 (N_6832,N_4778,N_3024);
nor U6833 (N_6833,N_4408,N_4495);
and U6834 (N_6834,N_4854,N_4576);
nor U6835 (N_6835,N_3136,N_4292);
or U6836 (N_6836,N_4345,N_3684);
nand U6837 (N_6837,N_4387,N_4117);
and U6838 (N_6838,N_3787,N_4079);
or U6839 (N_6839,N_4140,N_3514);
or U6840 (N_6840,N_5542,N_3413);
nand U6841 (N_6841,N_3092,N_4284);
or U6842 (N_6842,N_4874,N_3291);
and U6843 (N_6843,N_4672,N_5781);
or U6844 (N_6844,N_5775,N_3772);
or U6845 (N_6845,N_5655,N_5908);
or U6846 (N_6846,N_5736,N_3556);
nor U6847 (N_6847,N_3686,N_5413);
and U6848 (N_6848,N_5520,N_3065);
nor U6849 (N_6849,N_5000,N_5581);
nor U6850 (N_6850,N_3839,N_4897);
or U6851 (N_6851,N_5837,N_3519);
or U6852 (N_6852,N_3094,N_4578);
nand U6853 (N_6853,N_4520,N_4175);
nor U6854 (N_6854,N_3187,N_4643);
or U6855 (N_6855,N_5674,N_5010);
nand U6856 (N_6856,N_3215,N_5094);
and U6857 (N_6857,N_5218,N_4477);
and U6858 (N_6858,N_5102,N_4267);
nand U6859 (N_6859,N_4639,N_5265);
nand U6860 (N_6860,N_4995,N_5719);
or U6861 (N_6861,N_3741,N_3744);
nor U6862 (N_6862,N_4447,N_5366);
and U6863 (N_6863,N_4290,N_5164);
nor U6864 (N_6864,N_4024,N_3811);
and U6865 (N_6865,N_5282,N_4689);
and U6866 (N_6866,N_3870,N_5066);
and U6867 (N_6867,N_3692,N_3634);
or U6868 (N_6868,N_3982,N_5283);
or U6869 (N_6869,N_5419,N_3375);
nand U6870 (N_6870,N_5425,N_4913);
and U6871 (N_6871,N_3675,N_3069);
nor U6872 (N_6872,N_3377,N_5040);
or U6873 (N_6873,N_5187,N_5712);
and U6874 (N_6874,N_4768,N_4608);
nor U6875 (N_6875,N_4431,N_3783);
and U6876 (N_6876,N_3594,N_5168);
or U6877 (N_6877,N_4685,N_3712);
nor U6878 (N_6878,N_4765,N_3951);
nand U6879 (N_6879,N_5170,N_3452);
nor U6880 (N_6880,N_3608,N_5223);
nand U6881 (N_6881,N_3258,N_3654);
nor U6882 (N_6882,N_3191,N_3873);
or U6883 (N_6883,N_5479,N_4218);
nand U6884 (N_6884,N_4560,N_5598);
nand U6885 (N_6885,N_4320,N_3080);
and U6886 (N_6886,N_3108,N_5608);
and U6887 (N_6887,N_3492,N_5004);
nand U6888 (N_6888,N_3803,N_5519);
nand U6889 (N_6889,N_3247,N_4230);
or U6890 (N_6890,N_5944,N_4143);
nor U6891 (N_6891,N_4185,N_4538);
or U6892 (N_6892,N_5496,N_5505);
and U6893 (N_6893,N_4352,N_4695);
nor U6894 (N_6894,N_3986,N_4330);
or U6895 (N_6895,N_5220,N_4229);
nand U6896 (N_6896,N_5410,N_4993);
nand U6897 (N_6897,N_3381,N_4536);
nor U6898 (N_6898,N_3794,N_4113);
and U6899 (N_6899,N_5703,N_5651);
or U6900 (N_6900,N_5380,N_3920);
and U6901 (N_6901,N_5342,N_4410);
nand U6902 (N_6902,N_3252,N_3600);
and U6903 (N_6903,N_5087,N_4068);
nand U6904 (N_6904,N_5271,N_5738);
or U6905 (N_6905,N_4648,N_3125);
nor U6906 (N_6906,N_3725,N_3498);
and U6907 (N_6907,N_3751,N_5476);
nand U6908 (N_6908,N_3406,N_3368);
nor U6909 (N_6909,N_4032,N_4640);
and U6910 (N_6910,N_4196,N_5980);
nand U6911 (N_6911,N_4600,N_4197);
nand U6912 (N_6912,N_5478,N_5498);
nor U6913 (N_6913,N_3973,N_5693);
or U6914 (N_6914,N_3336,N_4921);
and U6915 (N_6915,N_5280,N_5983);
or U6916 (N_6916,N_4767,N_5325);
or U6917 (N_6917,N_3705,N_4276);
nand U6918 (N_6918,N_4570,N_5460);
or U6919 (N_6919,N_4498,N_5858);
or U6920 (N_6920,N_3888,N_3868);
nor U6921 (N_6921,N_3150,N_5485);
or U6922 (N_6922,N_4469,N_4323);
nand U6923 (N_6923,N_5798,N_4439);
and U6924 (N_6924,N_5016,N_4506);
nand U6925 (N_6925,N_4332,N_3567);
and U6926 (N_6926,N_3131,N_5357);
and U6927 (N_6927,N_3155,N_3175);
or U6928 (N_6928,N_3524,N_4390);
and U6929 (N_6929,N_3264,N_3558);
and U6930 (N_6930,N_3527,N_5110);
nor U6931 (N_6931,N_3190,N_4559);
or U6932 (N_6932,N_4004,N_5982);
and U6933 (N_6933,N_5571,N_3370);
and U6934 (N_6934,N_3836,N_4003);
and U6935 (N_6935,N_5881,N_3093);
nand U6936 (N_6936,N_4383,N_5395);
nor U6937 (N_6937,N_3475,N_4752);
nand U6938 (N_6938,N_3339,N_4969);
and U6939 (N_6939,N_4554,N_5841);
and U6940 (N_6940,N_3715,N_5586);
nor U6941 (N_6941,N_3957,N_3130);
and U6942 (N_6942,N_5331,N_3629);
or U6943 (N_6943,N_4134,N_5653);
nand U6944 (N_6944,N_5848,N_3211);
or U6945 (N_6945,N_5584,N_3670);
nand U6946 (N_6946,N_5701,N_5763);
and U6947 (N_6947,N_3644,N_5817);
nor U6948 (N_6948,N_5426,N_3635);
nand U6949 (N_6949,N_3224,N_5138);
and U6950 (N_6950,N_3157,N_4834);
and U6951 (N_6951,N_4707,N_4176);
nand U6952 (N_6952,N_5874,N_3945);
and U6953 (N_6953,N_5904,N_4235);
or U6954 (N_6954,N_5133,N_4604);
or U6955 (N_6955,N_5765,N_5149);
or U6956 (N_6956,N_4649,N_4111);
nand U6957 (N_6957,N_3766,N_3884);
nor U6958 (N_6958,N_3740,N_5189);
nor U6959 (N_6959,N_4116,N_4048);
nand U6960 (N_6960,N_4278,N_3640);
nand U6961 (N_6961,N_5017,N_4613);
nand U6962 (N_6962,N_5573,N_4543);
or U6963 (N_6963,N_4631,N_4186);
and U6964 (N_6964,N_5898,N_4664);
nor U6965 (N_6965,N_3685,N_4824);
nand U6966 (N_6966,N_3895,N_3905);
nand U6967 (N_6967,N_3463,N_4349);
xnor U6968 (N_6968,N_4848,N_4916);
and U6969 (N_6969,N_5686,N_4863);
nor U6970 (N_6970,N_4951,N_5026);
xor U6971 (N_6971,N_3909,N_5697);
and U6972 (N_6972,N_5885,N_3708);
nand U6973 (N_6973,N_3583,N_4416);
or U6974 (N_6974,N_5045,N_4428);
and U6975 (N_6975,N_5482,N_5905);
nand U6976 (N_6976,N_4843,N_3638);
and U6977 (N_6977,N_5212,N_4467);
nand U6978 (N_6978,N_4337,N_3798);
and U6979 (N_6979,N_4131,N_3100);
nand U6980 (N_6980,N_5920,N_5471);
nand U6981 (N_6981,N_5708,N_4346);
nand U6982 (N_6982,N_4490,N_3432);
and U6983 (N_6983,N_3773,N_3397);
or U6984 (N_6984,N_5981,N_4233);
nor U6985 (N_6985,N_5457,N_4317);
and U6986 (N_6986,N_4450,N_4184);
nand U6987 (N_6987,N_5256,N_3651);
nor U6988 (N_6988,N_3894,N_4063);
nor U6989 (N_6989,N_4770,N_5454);
nor U6990 (N_6990,N_3750,N_5269);
and U6991 (N_6991,N_3542,N_4749);
nand U6992 (N_6992,N_3453,N_3138);
and U6993 (N_6993,N_3707,N_4127);
nor U6994 (N_6994,N_4812,N_3887);
or U6995 (N_6995,N_4430,N_3057);
nand U6996 (N_6996,N_3294,N_3319);
or U6997 (N_6997,N_4663,N_4697);
and U6998 (N_6998,N_5641,N_5124);
or U6999 (N_6999,N_3030,N_5948);
nor U7000 (N_7000,N_4540,N_3424);
and U7001 (N_7001,N_3520,N_4168);
nand U7002 (N_7002,N_5864,N_5371);
nor U7003 (N_7003,N_5658,N_4182);
nor U7004 (N_7004,N_3843,N_5304);
nor U7005 (N_7005,N_4132,N_3579);
and U7006 (N_7006,N_4342,N_5659);
nor U7007 (N_7007,N_5473,N_5599);
nand U7008 (N_7008,N_5224,N_4706);
and U7009 (N_7009,N_3323,N_5861);
nand U7010 (N_7010,N_3196,N_5135);
nor U7011 (N_7011,N_3758,N_5300);
nor U7012 (N_7012,N_4998,N_4055);
nand U7013 (N_7013,N_3990,N_3404);
or U7014 (N_7014,N_5125,N_4655);
nand U7015 (N_7015,N_5650,N_4693);
and U7016 (N_7016,N_5153,N_4769);
and U7017 (N_7017,N_4147,N_4360);
and U7018 (N_7018,N_3185,N_4282);
nor U7019 (N_7019,N_4736,N_5974);
or U7020 (N_7020,N_5369,N_4698);
nor U7021 (N_7021,N_5992,N_3933);
and U7022 (N_7022,N_3797,N_3699);
and U7023 (N_7023,N_4915,N_5141);
and U7024 (N_7024,N_5959,N_5096);
and U7025 (N_7025,N_3260,N_4210);
nand U7026 (N_7026,N_5644,N_5946);
or U7027 (N_7027,N_5935,N_3653);
and U7028 (N_7028,N_3373,N_5480);
nand U7029 (N_7029,N_5088,N_3597);
and U7030 (N_7030,N_4391,N_4306);
nor U7031 (N_7031,N_5157,N_3417);
or U7032 (N_7032,N_3506,N_3924);
or U7033 (N_7033,N_3525,N_5646);
nand U7034 (N_7034,N_4072,N_4865);
and U7035 (N_7035,N_3019,N_3598);
and U7036 (N_7036,N_5098,N_4615);
or U7037 (N_7037,N_5929,N_4012);
nand U7038 (N_7038,N_3072,N_3812);
nor U7039 (N_7039,N_3569,N_3623);
nand U7040 (N_7040,N_5953,N_4098);
nand U7041 (N_7041,N_4367,N_3643);
nor U7042 (N_7042,N_3938,N_3709);
and U7043 (N_7043,N_5336,N_4444);
and U7044 (N_7044,N_5274,N_4150);
and U7045 (N_7045,N_5155,N_4750);
and U7046 (N_7046,N_4039,N_5600);
and U7047 (N_7047,N_3304,N_3169);
or U7048 (N_7048,N_3011,N_3918);
and U7049 (N_7049,N_3183,N_3776);
nand U7050 (N_7050,N_5432,N_3170);
nor U7051 (N_7051,N_4189,N_4223);
or U7052 (N_7052,N_4595,N_4888);
nand U7053 (N_7053,N_5647,N_3738);
and U7054 (N_7054,N_5972,N_3074);
nor U7055 (N_7055,N_4154,N_5743);
nor U7056 (N_7056,N_5530,N_5711);
or U7057 (N_7057,N_3230,N_4000);
or U7058 (N_7058,N_5810,N_3694);
nor U7059 (N_7059,N_4944,N_3112);
and U7060 (N_7060,N_5724,N_5219);
nand U7061 (N_7061,N_3677,N_3287);
nor U7062 (N_7062,N_3318,N_3042);
nor U7063 (N_7063,N_3371,N_4846);
and U7064 (N_7064,N_5570,N_5769);
nand U7065 (N_7065,N_3745,N_5101);
or U7066 (N_7066,N_5790,N_4254);
nand U7067 (N_7067,N_4933,N_5985);
and U7068 (N_7068,N_3141,N_4699);
or U7069 (N_7069,N_4359,N_4365);
nor U7070 (N_7070,N_4831,N_5794);
nand U7071 (N_7071,N_5886,N_4908);
nand U7072 (N_7072,N_5872,N_3910);
nand U7073 (N_7073,N_3489,N_5286);
and U7074 (N_7074,N_5613,N_4574);
nor U7075 (N_7075,N_3279,N_4716);
or U7076 (N_7076,N_5054,N_5364);
or U7077 (N_7077,N_5597,N_4471);
nand U7078 (N_7078,N_5918,N_4610);
nor U7079 (N_7079,N_4269,N_3818);
and U7080 (N_7080,N_4424,N_3702);
or U7081 (N_7081,N_4109,N_4502);
and U7082 (N_7082,N_5755,N_5846);
nor U7083 (N_7083,N_4786,N_4106);
nor U7084 (N_7084,N_3789,N_4130);
nand U7085 (N_7085,N_5662,N_5100);
and U7086 (N_7086,N_5148,N_4975);
nor U7087 (N_7087,N_4500,N_3448);
or U7088 (N_7088,N_4886,N_5976);
nand U7089 (N_7089,N_4852,N_5575);
nor U7090 (N_7090,N_3676,N_4790);
nand U7091 (N_7091,N_4421,N_4344);
nand U7092 (N_7092,N_5836,N_4338);
and U7093 (N_7093,N_3367,N_3476);
and U7094 (N_7094,N_3988,N_3421);
nand U7095 (N_7095,N_4792,N_3429);
or U7096 (N_7096,N_3831,N_3266);
and U7097 (N_7097,N_3274,N_5079);
nor U7098 (N_7098,N_3234,N_4795);
nand U7099 (N_7099,N_3114,N_4525);
and U7100 (N_7100,N_4719,N_4660);
nor U7101 (N_7101,N_3444,N_3871);
nand U7102 (N_7102,N_3356,N_3916);
nor U7103 (N_7103,N_5309,N_3526);
or U7104 (N_7104,N_5955,N_4898);
and U7105 (N_7105,N_4195,N_3277);
nand U7106 (N_7106,N_5979,N_5870);
or U7107 (N_7107,N_3273,N_3879);
and U7108 (N_7108,N_4711,N_3698);
nor U7109 (N_7109,N_3971,N_3161);
or U7110 (N_7110,N_4401,N_5210);
and U7111 (N_7111,N_3376,N_3536);
nand U7112 (N_7112,N_3047,N_4936);
nand U7113 (N_7113,N_4597,N_5109);
nand U7114 (N_7114,N_3327,N_3427);
and U7115 (N_7115,N_4992,N_3782);
or U7116 (N_7116,N_3889,N_5472);
xnor U7117 (N_7117,N_4178,N_4755);
nand U7118 (N_7118,N_3720,N_3806);
nor U7119 (N_7119,N_3848,N_5002);
nor U7120 (N_7120,N_3425,N_5773);
and U7121 (N_7121,N_5777,N_3792);
nand U7122 (N_7122,N_4295,N_5393);
nand U7123 (N_7123,N_4709,N_5486);
or U7124 (N_7124,N_5540,N_3408);
or U7125 (N_7125,N_4661,N_5303);
or U7126 (N_7126,N_4823,N_5967);
nor U7127 (N_7127,N_4418,N_5632);
nand U7128 (N_7128,N_3622,N_4508);
nor U7129 (N_7129,N_3912,N_4637);
or U7130 (N_7130,N_3261,N_4541);
or U7131 (N_7131,N_4049,N_5728);
nor U7132 (N_7132,N_3143,N_4013);
nand U7133 (N_7133,N_3473,N_4895);
nand U7134 (N_7134,N_3242,N_3351);
or U7135 (N_7135,N_5261,N_5445);
or U7136 (N_7136,N_4690,N_5120);
nor U7137 (N_7137,N_5169,N_4146);
or U7138 (N_7138,N_3999,N_3467);
nor U7139 (N_7139,N_3769,N_5278);
and U7140 (N_7140,N_4118,N_5204);
or U7141 (N_7141,N_4059,N_4862);
nand U7142 (N_7142,N_5430,N_4889);
or U7143 (N_7143,N_3126,N_5060);
nand U7144 (N_7144,N_4052,N_4355);
or U7145 (N_7145,N_4348,N_3921);
or U7146 (N_7146,N_5200,N_4505);
or U7147 (N_7147,N_4717,N_4119);
or U7148 (N_7148,N_3254,N_5385);
nor U7149 (N_7149,N_3388,N_5902);
or U7150 (N_7150,N_5637,N_3203);
nand U7151 (N_7151,N_5173,N_4612);
xor U7152 (N_7152,N_3474,N_5549);
or U7153 (N_7153,N_5812,N_4339);
nor U7154 (N_7154,N_4044,N_5761);
or U7155 (N_7155,N_4891,N_5890);
or U7156 (N_7156,N_4764,N_5629);
and U7157 (N_7157,N_3807,N_4499);
nand U7158 (N_7158,N_5242,N_4727);
nor U7159 (N_7159,N_3965,N_5796);
nor U7160 (N_7160,N_4590,N_4714);
or U7161 (N_7161,N_5150,N_4832);
nor U7162 (N_7162,N_3505,N_4827);
and U7163 (N_7163,N_5216,N_5896);
nor U7164 (N_7164,N_5503,N_4397);
nand U7165 (N_7165,N_3364,N_5834);
nand U7166 (N_7166,N_5394,N_4857);
nor U7167 (N_7167,N_5127,N_5648);
and U7168 (N_7168,N_4668,N_3625);
nor U7169 (N_7169,N_4582,N_4618);
or U7170 (N_7170,N_4020,N_4449);
and U7171 (N_7171,N_3168,N_3955);
and U7172 (N_7172,N_5263,N_4030);
nand U7173 (N_7173,N_4370,N_5475);
or U7174 (N_7174,N_5673,N_4493);
nor U7175 (N_7175,N_4872,N_3135);
nand U7176 (N_7176,N_5221,N_5806);
or U7177 (N_7177,N_4564,N_3906);
nor U7178 (N_7178,N_3084,N_3682);
and U7179 (N_7179,N_4219,N_4694);
or U7180 (N_7180,N_5416,N_3952);
nor U7181 (N_7181,N_5112,N_3288);
and U7182 (N_7182,N_3342,N_5737);
nand U7183 (N_7183,N_3941,N_4849);
or U7184 (N_7184,N_4628,N_3762);
nor U7185 (N_7185,N_3290,N_3416);
nor U7186 (N_7186,N_3810,N_3314);
or U7187 (N_7187,N_4946,N_5582);
or U7188 (N_7188,N_5352,N_5401);
xnor U7189 (N_7189,N_3746,N_5752);
nor U7190 (N_7190,N_5243,N_4460);
or U7191 (N_7191,N_5553,N_5772);
or U7192 (N_7192,N_5349,N_5619);
nand U7193 (N_7193,N_3055,N_4510);
and U7194 (N_7194,N_5233,N_5431);
nor U7195 (N_7195,N_3105,N_4566);
nor U7196 (N_7196,N_3239,N_4062);
and U7197 (N_7197,N_4868,N_4145);
nand U7198 (N_7198,N_3757,N_5882);
and U7199 (N_7199,N_5602,N_5785);
and U7200 (N_7200,N_5305,N_5228);
nor U7201 (N_7201,N_5408,N_3353);
or U7202 (N_7202,N_5634,N_3531);
and U7203 (N_7203,N_3490,N_4374);
and U7204 (N_7204,N_4310,N_5554);
nor U7205 (N_7205,N_4704,N_4361);
nor U7206 (N_7206,N_5477,N_3923);
xnor U7207 (N_7207,N_3046,N_4583);
and U7208 (N_7208,N_3315,N_5456);
or U7209 (N_7209,N_3499,N_3486);
nor U7210 (N_7210,N_3618,N_3726);
nor U7211 (N_7211,N_4986,N_5960);
nand U7212 (N_7212,N_5470,N_5507);
and U7213 (N_7213,N_4729,N_5231);
nor U7214 (N_7214,N_4732,N_4069);
nand U7215 (N_7215,N_5833,N_5927);
or U7216 (N_7216,N_4102,N_3194);
nand U7217 (N_7217,N_5245,N_3022);
nor U7218 (N_7218,N_5423,N_5030);
nor U7219 (N_7219,N_5706,N_5313);
or U7220 (N_7220,N_4710,N_3109);
nand U7221 (N_7221,N_4747,N_3855);
nor U7222 (N_7222,N_5050,N_3033);
and U7223 (N_7223,N_4960,N_4829);
nand U7224 (N_7224,N_3326,N_5370);
nor U7225 (N_7225,N_3436,N_4187);
nor U7226 (N_7226,N_4565,N_4017);
or U7227 (N_7227,N_5072,N_5952);
nand U7228 (N_7228,N_5789,N_3391);
nor U7229 (N_7229,N_3068,N_3298);
nand U7230 (N_7230,N_3227,N_4651);
and U7231 (N_7231,N_3472,N_3913);
or U7232 (N_7232,N_4573,N_5354);
or U7233 (N_7233,N_4294,N_3547);
nor U7234 (N_7234,N_5195,N_3271);
nor U7235 (N_7235,N_3346,N_4288);
nor U7236 (N_7236,N_4577,N_4748);
nor U7237 (N_7237,N_3387,N_5031);
nor U7238 (N_7238,N_3885,N_5567);
and U7239 (N_7239,N_5580,N_5034);
or U7240 (N_7240,N_5847,N_3098);
and U7241 (N_7241,N_3903,N_3199);
and U7242 (N_7242,N_4300,N_5338);
and U7243 (N_7243,N_4065,N_3853);
or U7244 (N_7244,N_3335,N_5136);
nor U7245 (N_7245,N_3021,N_5450);
nand U7246 (N_7246,N_5564,N_3790);
or U7247 (N_7247,N_5118,N_5667);
nor U7248 (N_7248,N_4414,N_4773);
nor U7249 (N_7249,N_4491,N_3337);
and U7250 (N_7250,N_5378,N_4216);
and U7251 (N_7251,N_4851,N_4126);
and U7252 (N_7252,N_5956,N_4011);
and U7253 (N_7253,N_4114,N_3512);
nor U7254 (N_7254,N_3000,N_3805);
nand U7255 (N_7255,N_3585,N_5934);
nor U7256 (N_7256,N_5255,N_3574);
nor U7257 (N_7257,N_5249,N_4389);
nand U7258 (N_7258,N_3235,N_3220);
and U7259 (N_7259,N_3591,N_4075);
nand U7260 (N_7260,N_5688,N_4950);
nand U7261 (N_7261,N_4046,N_4279);
nand U7262 (N_7262,N_3392,N_4472);
or U7263 (N_7263,N_3770,N_4239);
or U7264 (N_7264,N_5422,N_4309);
nor U7265 (N_7265,N_3385,N_4494);
or U7266 (N_7266,N_3043,N_3799);
nand U7267 (N_7267,N_4692,N_5501);
and U7268 (N_7268,N_4291,N_3248);
nand U7269 (N_7269,N_5740,N_3983);
or U7270 (N_7270,N_3292,N_5968);
nor U7271 (N_7271,N_5911,N_5783);
nand U7272 (N_7272,N_5938,N_3180);
nor U7273 (N_7273,N_5522,N_4286);
nor U7274 (N_7274,N_5095,N_3605);
nor U7275 (N_7275,N_4083,N_4798);
xor U7276 (N_7276,N_4605,N_3674);
or U7277 (N_7277,N_5594,N_5601);
nor U7278 (N_7278,N_4518,N_4546);
and U7279 (N_7279,N_5437,N_3540);
nand U7280 (N_7280,N_4994,N_3389);
nand U7281 (N_7281,N_3518,N_4734);
nor U7282 (N_7282,N_4781,N_4080);
or U7283 (N_7283,N_3718,N_5020);
nand U7284 (N_7284,N_4978,N_3297);
or U7285 (N_7285,N_5053,N_4357);
or U7286 (N_7286,N_3372,N_3428);
xor U7287 (N_7287,N_5668,N_5887);
and U7288 (N_7288,N_3204,N_5827);
and U7289 (N_7289,N_5795,N_3917);
xnor U7290 (N_7290,N_5925,N_4634);
or U7291 (N_7291,N_5248,N_4038);
and U7292 (N_7292,N_3820,N_5386);
nor U7293 (N_7293,N_4805,N_5994);
nand U7294 (N_7294,N_3780,N_5880);
nand U7295 (N_7295,N_4724,N_3765);
or U7296 (N_7296,N_5483,N_5277);
nand U7297 (N_7297,N_4245,N_4743);
nor U7298 (N_7298,N_3970,N_4050);
nand U7299 (N_7299,N_4241,N_4441);
and U7300 (N_7300,N_5551,N_3129);
and U7301 (N_7301,N_4244,N_3665);
or U7302 (N_7302,N_5626,N_3646);
nor U7303 (N_7303,N_5593,N_3340);
nand U7304 (N_7304,N_4207,N_4616);
and U7305 (N_7305,N_3603,N_5091);
nor U7306 (N_7306,N_5517,N_5022);
nand U7307 (N_7307,N_3760,N_4922);
or U7308 (N_7308,N_5576,N_5046);
nand U7309 (N_7309,N_5427,N_5879);
or U7310 (N_7310,N_4089,N_4811);
or U7311 (N_7311,N_5131,N_4601);
or U7312 (N_7312,N_4776,N_3280);
or U7313 (N_7313,N_5565,N_3914);
nor U7314 (N_7314,N_3418,N_5508);
nor U7315 (N_7315,N_3826,N_3502);
and U7316 (N_7316,N_3604,N_4804);
nor U7317 (N_7317,N_5557,N_3516);
or U7318 (N_7318,N_5984,N_4669);
and U7319 (N_7319,N_4094,N_5928);
or U7320 (N_7320,N_5225,N_5897);
and U7321 (N_7321,N_3088,N_3111);
and U7322 (N_7322,N_5092,N_3582);
and U7323 (N_7323,N_4890,N_3278);
nand U7324 (N_7324,N_5912,N_5808);
and U7325 (N_7325,N_5119,N_4519);
and U7326 (N_7326,N_3969,N_3593);
or U7327 (N_7327,N_3513,N_4183);
or U7328 (N_7328,N_5397,N_4818);
nand U7329 (N_7329,N_4537,N_5809);
nor U7330 (N_7330,N_4650,N_4042);
nand U7331 (N_7331,N_5640,N_5871);
and U7332 (N_7332,N_3822,N_5694);
and U7333 (N_7333,N_5146,N_4522);
nand U7334 (N_7334,N_5829,N_3500);
and U7335 (N_7335,N_4635,N_3202);
nor U7336 (N_7336,N_5621,N_3255);
and U7337 (N_7337,N_4268,N_5063);
and U7338 (N_7338,N_3149,N_5207);
and U7339 (N_7339,N_4627,N_3362);
nand U7340 (N_7340,N_4965,N_3523);
nor U7341 (N_7341,N_5253,N_5122);
nand U7342 (N_7342,N_3015,N_3979);
nand U7343 (N_7343,N_4058,N_3330);
or U7344 (N_7344,N_5585,N_4785);
nand U7345 (N_7345,N_5961,N_3876);
or U7346 (N_7346,N_4386,N_3259);
nor U7347 (N_7347,N_4821,N_4496);
nand U7348 (N_7348,N_3115,N_5387);
or U7349 (N_7349,N_4988,N_4220);
or U7350 (N_7350,N_4199,N_4287);
nand U7351 (N_7351,N_3943,N_4885);
nand U7352 (N_7352,N_3159,N_4636);
and U7353 (N_7353,N_4558,N_3991);
nor U7354 (N_7354,N_3197,N_5448);
nand U7355 (N_7355,N_4756,N_4550);
and U7356 (N_7356,N_3535,N_4925);
nor U7357 (N_7357,N_4302,N_4377);
nand U7358 (N_7358,N_3652,N_4454);
nand U7359 (N_7359,N_5297,N_5949);
nand U7360 (N_7360,N_3176,N_5552);
and U7361 (N_7361,N_4191,N_5292);
and U7362 (N_7362,N_3566,N_3944);
nand U7363 (N_7363,N_4188,N_4078);
or U7364 (N_7364,N_5481,N_4322);
nand U7365 (N_7365,N_3961,N_5469);
or U7366 (N_7366,N_3731,N_3321);
or U7367 (N_7367,N_5029,N_4112);
nand U7368 (N_7368,N_4343,N_5374);
nor U7369 (N_7369,N_3573,N_3118);
nor U7370 (N_7370,N_5025,N_3934);
or U7371 (N_7371,N_3553,N_5459);
nor U7372 (N_7372,N_3460,N_5301);
and U7373 (N_7373,N_3639,N_4561);
nand U7374 (N_7374,N_4371,N_3009);
nand U7375 (N_7375,N_5759,N_4883);
or U7376 (N_7376,N_5409,N_4404);
or U7377 (N_7377,N_5524,N_5494);
nor U7378 (N_7378,N_4394,N_5344);
or U7379 (N_7379,N_3504,N_3530);
xor U7380 (N_7380,N_3172,N_4022);
and U7381 (N_7381,N_5420,N_4077);
and U7382 (N_7382,N_3845,N_4100);
nand U7383 (N_7383,N_3198,N_3815);
nand U7384 (N_7384,N_4952,N_4315);
nor U7385 (N_7385,N_4082,N_4324);
nor U7386 (N_7386,N_3759,N_3054);
and U7387 (N_7387,N_5363,N_4107);
and U7388 (N_7388,N_4810,N_4101);
nor U7389 (N_7389,N_4856,N_4014);
nand U7390 (N_7390,N_4152,N_3954);
and U7391 (N_7391,N_4680,N_5324);
nand U7392 (N_7392,N_4735,N_3289);
nor U7393 (N_7393,N_5963,N_3303);
or U7394 (N_7394,N_3028,N_4167);
nor U7395 (N_7395,N_5376,N_3656);
nand U7396 (N_7396,N_3035,N_5857);
or U7397 (N_7397,N_5320,N_5288);
and U7398 (N_7398,N_5208,N_4845);
or U7399 (N_7399,N_3966,N_3788);
nor U7400 (N_7400,N_3571,N_4772);
nor U7401 (N_7401,N_4299,N_5699);
and U7402 (N_7402,N_5727,N_5126);
or U7403 (N_7403,N_3994,N_3967);
nor U7404 (N_7404,N_5275,N_3735);
and U7405 (N_7405,N_5625,N_5663);
or U7406 (N_7406,N_4587,N_4983);
or U7407 (N_7407,N_3713,N_4909);
nand U7408 (N_7408,N_3038,N_5339);
nand U7409 (N_7409,N_3834,N_5284);
nor U7410 (N_7410,N_4208,N_4679);
and U7411 (N_7411,N_5057,N_5259);
nand U7412 (N_7412,N_4847,N_4659);
and U7413 (N_7413,N_4458,N_3433);
nor U7414 (N_7414,N_3719,N_5144);
nor U7415 (N_7415,N_5859,N_4603);
nor U7416 (N_7416,N_5679,N_3592);
and U7417 (N_7417,N_5677,N_5652);
nand U7418 (N_7418,N_5649,N_5358);
and U7419 (N_7419,N_5252,N_3296);
and U7420 (N_7420,N_3753,N_5900);
xor U7421 (N_7421,N_4585,N_5610);
nand U7422 (N_7422,N_5768,N_4956);
nand U7423 (N_7423,N_4071,N_3005);
nand U7424 (N_7424,N_4968,N_4455);
and U7425 (N_7425,N_3577,N_3494);
nand U7426 (N_7426,N_4067,N_4249);
nand U7427 (N_7427,N_4696,N_3300);
nor U7428 (N_7428,N_5614,N_3382);
nor U7429 (N_7429,N_5936,N_3847);
nor U7430 (N_7430,N_3667,N_4110);
or U7431 (N_7431,N_4091,N_3880);
or U7432 (N_7432,N_5368,N_3225);
nand U7433 (N_7433,N_4910,N_3507);
and U7434 (N_7434,N_5671,N_4171);
nand U7435 (N_7435,N_4876,N_4838);
nor U7436 (N_7436,N_4021,N_4589);
nor U7437 (N_7437,N_5853,N_4266);
or U7438 (N_7438,N_3491,N_5780);
nand U7439 (N_7439,N_3036,N_5443);
and U7440 (N_7440,N_5807,N_4232);
nor U7441 (N_7441,N_5993,N_3140);
nand U7442 (N_7442,N_3584,N_4870);
or U7443 (N_7443,N_4524,N_4090);
nand U7444 (N_7444,N_3886,N_4977);
nor U7445 (N_7445,N_4777,N_5734);
nor U7446 (N_7446,N_4954,N_5281);
or U7447 (N_7447,N_5932,N_5914);
nand U7448 (N_7448,N_5536,N_5860);
or U7449 (N_7449,N_4841,N_3827);
and U7450 (N_7450,N_3401,N_4422);
nor U7451 (N_7451,N_4445,N_3900);
nand U7452 (N_7452,N_5024,N_3410);
and U7453 (N_7453,N_5970,N_3575);
nand U7454 (N_7454,N_5293,N_3133);
and U7455 (N_7455,N_5587,N_5392);
and U7456 (N_7456,N_3669,N_3736);
or U7457 (N_7457,N_3814,N_4086);
or U7458 (N_7458,N_3066,N_4271);
nand U7459 (N_7459,N_4758,N_5924);
nor U7460 (N_7460,N_5190,N_3320);
or U7461 (N_7461,N_5314,N_3222);
or U7462 (N_7462,N_4948,N_4513);
or U7463 (N_7463,N_3511,N_5147);
nor U7464 (N_7464,N_5322,N_3434);
nand U7465 (N_7465,N_3721,N_3627);
and U7466 (N_7466,N_5722,N_3032);
nand U7467 (N_7467,N_5191,N_3710);
or U7468 (N_7468,N_4405,N_3775);
xor U7469 (N_7469,N_5343,N_5942);
and U7470 (N_7470,N_5725,N_5762);
and U7471 (N_7471,N_3930,N_4814);
nand U7472 (N_7472,N_4924,N_5222);
nor U7473 (N_7473,N_3283,N_3145);
nand U7474 (N_7474,N_5214,N_4571);
nor U7475 (N_7475,N_3139,N_5097);
nand U7476 (N_7476,N_5174,N_3357);
and U7477 (N_7477,N_3348,N_5178);
nor U7478 (N_7478,N_3533,N_3528);
nor U7479 (N_7479,N_5950,N_5465);
and U7480 (N_7480,N_3974,N_5211);
nand U7481 (N_7481,N_5311,N_4962);
nor U7482 (N_7482,N_3754,N_4771);
and U7483 (N_7483,N_5534,N_5969);
and U7484 (N_7484,N_3016,N_4586);
nand U7485 (N_7485,N_4308,N_5424);
and U7486 (N_7486,N_5215,N_4087);
and U7487 (N_7487,N_4532,N_4135);
and U7488 (N_7488,N_4436,N_3509);
nand U7489 (N_7489,N_4530,N_3177);
nand U7490 (N_7490,N_3555,N_5516);
and U7491 (N_7491,N_4866,N_3031);
or U7492 (N_7492,N_5767,N_3875);
or U7493 (N_7493,N_3450,N_5468);
nor U7494 (N_7494,N_4728,N_5590);
nand U7495 (N_7495,N_4629,N_5639);
and U7496 (N_7496,N_4465,N_5446);
or U7497 (N_7497,N_4259,N_4625);
or U7498 (N_7498,N_5895,N_3545);
and U7499 (N_7499,N_3984,N_4996);
nor U7500 (N_7500,N_4659,N_3905);
nor U7501 (N_7501,N_4723,N_3640);
nand U7502 (N_7502,N_4119,N_3558);
nor U7503 (N_7503,N_5529,N_4251);
and U7504 (N_7504,N_3442,N_4610);
nor U7505 (N_7505,N_5504,N_3938);
and U7506 (N_7506,N_3925,N_4575);
xor U7507 (N_7507,N_3842,N_4755);
and U7508 (N_7508,N_4477,N_5390);
nand U7509 (N_7509,N_5862,N_4537);
or U7510 (N_7510,N_4795,N_5777);
xor U7511 (N_7511,N_3721,N_3086);
or U7512 (N_7512,N_3976,N_3638);
and U7513 (N_7513,N_4013,N_5447);
or U7514 (N_7514,N_4853,N_4653);
or U7515 (N_7515,N_3281,N_3937);
nor U7516 (N_7516,N_5000,N_4542);
nand U7517 (N_7517,N_5814,N_3130);
nand U7518 (N_7518,N_5736,N_3096);
nand U7519 (N_7519,N_3582,N_4372);
nor U7520 (N_7520,N_3135,N_4049);
nand U7521 (N_7521,N_5350,N_3333);
xor U7522 (N_7522,N_5602,N_3269);
and U7523 (N_7523,N_3928,N_4602);
and U7524 (N_7524,N_5212,N_3325);
nand U7525 (N_7525,N_5426,N_5906);
and U7526 (N_7526,N_3988,N_3666);
or U7527 (N_7527,N_5845,N_3084);
or U7528 (N_7528,N_5534,N_5210);
or U7529 (N_7529,N_3912,N_4769);
nor U7530 (N_7530,N_4945,N_4664);
and U7531 (N_7531,N_4786,N_3111);
nor U7532 (N_7532,N_3439,N_5283);
or U7533 (N_7533,N_3685,N_3111);
and U7534 (N_7534,N_3361,N_4990);
nand U7535 (N_7535,N_4104,N_5210);
or U7536 (N_7536,N_4591,N_4473);
nor U7537 (N_7537,N_4782,N_5995);
nor U7538 (N_7538,N_3130,N_5807);
or U7539 (N_7539,N_5395,N_3238);
nand U7540 (N_7540,N_4500,N_3723);
or U7541 (N_7541,N_3157,N_3580);
nand U7542 (N_7542,N_5370,N_4857);
nand U7543 (N_7543,N_4338,N_3592);
nand U7544 (N_7544,N_3603,N_5382);
and U7545 (N_7545,N_5441,N_3913);
nor U7546 (N_7546,N_5140,N_4107);
or U7547 (N_7547,N_5845,N_5774);
nor U7548 (N_7548,N_3836,N_4718);
nand U7549 (N_7549,N_4844,N_4663);
nor U7550 (N_7550,N_5418,N_5279);
and U7551 (N_7551,N_5199,N_4448);
nand U7552 (N_7552,N_4334,N_5874);
or U7553 (N_7553,N_4653,N_3685);
or U7554 (N_7554,N_4351,N_5889);
nor U7555 (N_7555,N_5642,N_4613);
xnor U7556 (N_7556,N_5939,N_4416);
and U7557 (N_7557,N_5419,N_4726);
and U7558 (N_7558,N_5013,N_3493);
or U7559 (N_7559,N_4110,N_3520);
nand U7560 (N_7560,N_3137,N_3798);
or U7561 (N_7561,N_5164,N_5109);
and U7562 (N_7562,N_5829,N_5375);
nand U7563 (N_7563,N_3711,N_3008);
nand U7564 (N_7564,N_4598,N_4471);
and U7565 (N_7565,N_5725,N_3456);
or U7566 (N_7566,N_5676,N_3742);
nor U7567 (N_7567,N_4997,N_4760);
nand U7568 (N_7568,N_5866,N_4166);
or U7569 (N_7569,N_3627,N_4666);
nor U7570 (N_7570,N_5933,N_5740);
and U7571 (N_7571,N_4464,N_3501);
or U7572 (N_7572,N_4083,N_5018);
xnor U7573 (N_7573,N_4240,N_3785);
nand U7574 (N_7574,N_5997,N_4450);
or U7575 (N_7575,N_3601,N_5148);
nor U7576 (N_7576,N_5771,N_5911);
xnor U7577 (N_7577,N_3021,N_4375);
nor U7578 (N_7578,N_4219,N_5433);
and U7579 (N_7579,N_5231,N_5077);
and U7580 (N_7580,N_3131,N_3264);
and U7581 (N_7581,N_5357,N_4865);
or U7582 (N_7582,N_4773,N_4813);
nor U7583 (N_7583,N_4602,N_5208);
nor U7584 (N_7584,N_4218,N_5993);
nand U7585 (N_7585,N_4164,N_4121);
or U7586 (N_7586,N_5869,N_5599);
nor U7587 (N_7587,N_5862,N_5952);
nand U7588 (N_7588,N_5052,N_3060);
and U7589 (N_7589,N_4649,N_5365);
nor U7590 (N_7590,N_5920,N_4822);
and U7591 (N_7591,N_3616,N_3927);
and U7592 (N_7592,N_3029,N_5787);
nand U7593 (N_7593,N_4498,N_5571);
nor U7594 (N_7594,N_4776,N_3341);
and U7595 (N_7595,N_4068,N_4357);
nor U7596 (N_7596,N_5591,N_4459);
or U7597 (N_7597,N_3061,N_5562);
and U7598 (N_7598,N_5356,N_5392);
or U7599 (N_7599,N_3792,N_5702);
nor U7600 (N_7600,N_5676,N_4643);
or U7601 (N_7601,N_4623,N_4932);
nand U7602 (N_7602,N_4632,N_4222);
nor U7603 (N_7603,N_4693,N_5376);
nor U7604 (N_7604,N_5342,N_3622);
and U7605 (N_7605,N_4295,N_4776);
or U7606 (N_7606,N_4270,N_5342);
nor U7607 (N_7607,N_4449,N_4226);
or U7608 (N_7608,N_4515,N_5879);
nand U7609 (N_7609,N_5354,N_4510);
nand U7610 (N_7610,N_4955,N_3502);
or U7611 (N_7611,N_5233,N_3523);
nor U7612 (N_7612,N_4435,N_3937);
and U7613 (N_7613,N_3887,N_4876);
nand U7614 (N_7614,N_3771,N_5235);
and U7615 (N_7615,N_3030,N_5460);
nor U7616 (N_7616,N_4207,N_4278);
nor U7617 (N_7617,N_4006,N_5959);
nor U7618 (N_7618,N_4405,N_5222);
nor U7619 (N_7619,N_3213,N_5188);
nor U7620 (N_7620,N_4407,N_3734);
nor U7621 (N_7621,N_3733,N_3644);
nor U7622 (N_7622,N_5542,N_4079);
or U7623 (N_7623,N_3513,N_4914);
nor U7624 (N_7624,N_5747,N_5322);
nand U7625 (N_7625,N_4010,N_3002);
nand U7626 (N_7626,N_5367,N_3854);
nor U7627 (N_7627,N_4071,N_5458);
and U7628 (N_7628,N_5331,N_4341);
nor U7629 (N_7629,N_3174,N_4367);
and U7630 (N_7630,N_5364,N_4371);
nand U7631 (N_7631,N_3037,N_4871);
nand U7632 (N_7632,N_4475,N_5130);
or U7633 (N_7633,N_3210,N_3774);
nor U7634 (N_7634,N_3354,N_5928);
and U7635 (N_7635,N_4779,N_4897);
or U7636 (N_7636,N_4135,N_3451);
or U7637 (N_7637,N_4801,N_4710);
nand U7638 (N_7638,N_5794,N_5095);
or U7639 (N_7639,N_3936,N_3149);
and U7640 (N_7640,N_4741,N_5265);
or U7641 (N_7641,N_3253,N_4007);
nor U7642 (N_7642,N_5396,N_3777);
and U7643 (N_7643,N_4742,N_3311);
and U7644 (N_7644,N_3573,N_3213);
nor U7645 (N_7645,N_5209,N_5483);
nand U7646 (N_7646,N_3779,N_4618);
nor U7647 (N_7647,N_4256,N_3899);
or U7648 (N_7648,N_3473,N_3058);
or U7649 (N_7649,N_5980,N_5535);
and U7650 (N_7650,N_3809,N_3735);
nand U7651 (N_7651,N_5592,N_3227);
and U7652 (N_7652,N_5078,N_4322);
nor U7653 (N_7653,N_4569,N_5221);
nor U7654 (N_7654,N_4497,N_4863);
nor U7655 (N_7655,N_4979,N_4190);
or U7656 (N_7656,N_3543,N_4976);
or U7657 (N_7657,N_4126,N_4269);
and U7658 (N_7658,N_5262,N_4930);
and U7659 (N_7659,N_3083,N_5366);
or U7660 (N_7660,N_4416,N_4955);
nor U7661 (N_7661,N_4259,N_5920);
or U7662 (N_7662,N_3730,N_3919);
and U7663 (N_7663,N_5529,N_3784);
nor U7664 (N_7664,N_5442,N_5687);
or U7665 (N_7665,N_3063,N_4936);
nand U7666 (N_7666,N_4164,N_5321);
or U7667 (N_7667,N_4254,N_3169);
nor U7668 (N_7668,N_5693,N_5994);
and U7669 (N_7669,N_4808,N_3550);
and U7670 (N_7670,N_3790,N_4789);
or U7671 (N_7671,N_5869,N_3486);
and U7672 (N_7672,N_4056,N_3678);
and U7673 (N_7673,N_3556,N_5961);
and U7674 (N_7674,N_4193,N_4775);
nand U7675 (N_7675,N_3666,N_4639);
or U7676 (N_7676,N_5959,N_4087);
nand U7677 (N_7677,N_5244,N_3083);
and U7678 (N_7678,N_3830,N_5821);
nor U7679 (N_7679,N_4690,N_5473);
or U7680 (N_7680,N_4804,N_4547);
and U7681 (N_7681,N_3528,N_4931);
nand U7682 (N_7682,N_3144,N_4809);
or U7683 (N_7683,N_4942,N_5517);
or U7684 (N_7684,N_5842,N_3410);
and U7685 (N_7685,N_4435,N_4869);
nand U7686 (N_7686,N_4033,N_4133);
and U7687 (N_7687,N_5480,N_5550);
and U7688 (N_7688,N_4305,N_5901);
or U7689 (N_7689,N_5420,N_3189);
or U7690 (N_7690,N_5483,N_4502);
nand U7691 (N_7691,N_3642,N_3159);
nor U7692 (N_7692,N_5574,N_5707);
nand U7693 (N_7693,N_3901,N_5556);
nand U7694 (N_7694,N_5800,N_5121);
nor U7695 (N_7695,N_4208,N_3533);
and U7696 (N_7696,N_3830,N_5717);
nor U7697 (N_7697,N_5526,N_3019);
or U7698 (N_7698,N_5196,N_3318);
or U7699 (N_7699,N_5632,N_5458);
nor U7700 (N_7700,N_5730,N_3815);
and U7701 (N_7701,N_5029,N_5981);
nand U7702 (N_7702,N_5084,N_4095);
nand U7703 (N_7703,N_5320,N_5744);
nor U7704 (N_7704,N_5884,N_3876);
or U7705 (N_7705,N_3091,N_4584);
xnor U7706 (N_7706,N_5202,N_4891);
or U7707 (N_7707,N_5596,N_3461);
or U7708 (N_7708,N_3731,N_3945);
nand U7709 (N_7709,N_5004,N_4203);
nand U7710 (N_7710,N_4348,N_4591);
nand U7711 (N_7711,N_3710,N_3082);
and U7712 (N_7712,N_3211,N_5414);
or U7713 (N_7713,N_5178,N_4307);
nand U7714 (N_7714,N_4928,N_3167);
nand U7715 (N_7715,N_5199,N_5735);
or U7716 (N_7716,N_5396,N_4331);
and U7717 (N_7717,N_5649,N_4061);
nor U7718 (N_7718,N_4893,N_3057);
and U7719 (N_7719,N_4754,N_4326);
xnor U7720 (N_7720,N_3877,N_5109);
or U7721 (N_7721,N_4413,N_4695);
or U7722 (N_7722,N_4316,N_4328);
or U7723 (N_7723,N_5170,N_3028);
or U7724 (N_7724,N_3257,N_5400);
and U7725 (N_7725,N_3356,N_5817);
and U7726 (N_7726,N_4821,N_4087);
or U7727 (N_7727,N_3371,N_3545);
xor U7728 (N_7728,N_5570,N_3019);
and U7729 (N_7729,N_4124,N_3739);
nand U7730 (N_7730,N_5199,N_3430);
and U7731 (N_7731,N_4516,N_5084);
or U7732 (N_7732,N_5822,N_5211);
or U7733 (N_7733,N_4933,N_3358);
or U7734 (N_7734,N_4284,N_3742);
nor U7735 (N_7735,N_4502,N_5755);
or U7736 (N_7736,N_4812,N_4455);
nor U7737 (N_7737,N_5311,N_4341);
nand U7738 (N_7738,N_4579,N_5298);
nand U7739 (N_7739,N_5703,N_5286);
nor U7740 (N_7740,N_3616,N_3606);
nor U7741 (N_7741,N_3952,N_3009);
or U7742 (N_7742,N_5549,N_3420);
nand U7743 (N_7743,N_3556,N_3448);
or U7744 (N_7744,N_5614,N_5378);
and U7745 (N_7745,N_4343,N_5901);
or U7746 (N_7746,N_3046,N_5278);
or U7747 (N_7747,N_3884,N_4319);
nand U7748 (N_7748,N_4619,N_3639);
nor U7749 (N_7749,N_3937,N_5750);
or U7750 (N_7750,N_4990,N_4625);
and U7751 (N_7751,N_3417,N_3445);
nor U7752 (N_7752,N_3725,N_5597);
and U7753 (N_7753,N_3797,N_3294);
nand U7754 (N_7754,N_5065,N_3156);
or U7755 (N_7755,N_4142,N_3040);
and U7756 (N_7756,N_4748,N_3631);
or U7757 (N_7757,N_4490,N_4361);
and U7758 (N_7758,N_4639,N_4968);
nand U7759 (N_7759,N_5535,N_5893);
nand U7760 (N_7760,N_3962,N_5812);
or U7761 (N_7761,N_4027,N_4210);
and U7762 (N_7762,N_4271,N_3475);
nor U7763 (N_7763,N_4887,N_3056);
nand U7764 (N_7764,N_3518,N_4651);
nor U7765 (N_7765,N_4111,N_4587);
nor U7766 (N_7766,N_4208,N_5935);
or U7767 (N_7767,N_5723,N_3201);
nor U7768 (N_7768,N_5511,N_5103);
or U7769 (N_7769,N_3437,N_4375);
nor U7770 (N_7770,N_4683,N_5069);
nor U7771 (N_7771,N_4230,N_4190);
nor U7772 (N_7772,N_4283,N_3767);
xnor U7773 (N_7773,N_4969,N_4054);
nand U7774 (N_7774,N_5517,N_5388);
nand U7775 (N_7775,N_3115,N_5937);
and U7776 (N_7776,N_3385,N_4921);
nand U7777 (N_7777,N_3053,N_3626);
or U7778 (N_7778,N_4544,N_5212);
nor U7779 (N_7779,N_5148,N_4939);
and U7780 (N_7780,N_5835,N_5686);
or U7781 (N_7781,N_4401,N_5202);
or U7782 (N_7782,N_4589,N_4102);
and U7783 (N_7783,N_5908,N_3649);
and U7784 (N_7784,N_5646,N_5868);
nor U7785 (N_7785,N_4556,N_3486);
or U7786 (N_7786,N_5512,N_5839);
nor U7787 (N_7787,N_5079,N_5158);
or U7788 (N_7788,N_3424,N_5818);
nor U7789 (N_7789,N_4458,N_3169);
or U7790 (N_7790,N_4179,N_3471);
or U7791 (N_7791,N_5025,N_3261);
nand U7792 (N_7792,N_4328,N_3285);
nand U7793 (N_7793,N_5637,N_5325);
and U7794 (N_7794,N_3660,N_3370);
or U7795 (N_7795,N_3896,N_4668);
nand U7796 (N_7796,N_4047,N_5895);
or U7797 (N_7797,N_5410,N_5642);
nor U7798 (N_7798,N_5224,N_3071);
and U7799 (N_7799,N_4365,N_5874);
or U7800 (N_7800,N_4058,N_4977);
nor U7801 (N_7801,N_3562,N_4673);
nor U7802 (N_7802,N_5675,N_3982);
nand U7803 (N_7803,N_3219,N_3432);
nand U7804 (N_7804,N_5846,N_4280);
or U7805 (N_7805,N_5401,N_3525);
nor U7806 (N_7806,N_3742,N_3942);
and U7807 (N_7807,N_5386,N_5142);
nor U7808 (N_7808,N_3788,N_3275);
nand U7809 (N_7809,N_5869,N_5337);
or U7810 (N_7810,N_5865,N_4794);
and U7811 (N_7811,N_5390,N_5140);
and U7812 (N_7812,N_4558,N_4923);
and U7813 (N_7813,N_5586,N_4311);
nor U7814 (N_7814,N_4383,N_3831);
and U7815 (N_7815,N_3888,N_5118);
xor U7816 (N_7816,N_5743,N_3361);
nor U7817 (N_7817,N_4119,N_5508);
nor U7818 (N_7818,N_3839,N_5302);
nor U7819 (N_7819,N_4570,N_3403);
or U7820 (N_7820,N_5164,N_4897);
nand U7821 (N_7821,N_5193,N_4327);
nand U7822 (N_7822,N_3982,N_3585);
or U7823 (N_7823,N_4915,N_5062);
and U7824 (N_7824,N_5534,N_3245);
or U7825 (N_7825,N_5380,N_3912);
nand U7826 (N_7826,N_3357,N_5089);
nor U7827 (N_7827,N_5018,N_4704);
nand U7828 (N_7828,N_3230,N_5842);
nand U7829 (N_7829,N_5895,N_5430);
nand U7830 (N_7830,N_5360,N_3195);
or U7831 (N_7831,N_4769,N_4122);
and U7832 (N_7832,N_4441,N_5695);
nand U7833 (N_7833,N_4581,N_4894);
and U7834 (N_7834,N_5842,N_4300);
nor U7835 (N_7835,N_4735,N_4284);
nor U7836 (N_7836,N_3312,N_3441);
and U7837 (N_7837,N_4910,N_4276);
nor U7838 (N_7838,N_5147,N_4227);
and U7839 (N_7839,N_3465,N_3038);
and U7840 (N_7840,N_4342,N_3375);
xnor U7841 (N_7841,N_4084,N_5187);
nand U7842 (N_7842,N_4429,N_3179);
nand U7843 (N_7843,N_5248,N_4040);
or U7844 (N_7844,N_4834,N_3459);
and U7845 (N_7845,N_3849,N_3947);
nor U7846 (N_7846,N_3021,N_5703);
or U7847 (N_7847,N_5007,N_4984);
or U7848 (N_7848,N_3719,N_4493);
or U7849 (N_7849,N_5966,N_3453);
nor U7850 (N_7850,N_3055,N_4076);
and U7851 (N_7851,N_4962,N_3627);
nand U7852 (N_7852,N_5711,N_4110);
or U7853 (N_7853,N_4256,N_4497);
or U7854 (N_7854,N_3512,N_5146);
and U7855 (N_7855,N_3964,N_5392);
nand U7856 (N_7856,N_4634,N_3016);
or U7857 (N_7857,N_4857,N_5835);
or U7858 (N_7858,N_3726,N_3546);
and U7859 (N_7859,N_3265,N_3758);
and U7860 (N_7860,N_4638,N_4781);
nor U7861 (N_7861,N_4886,N_3161);
nand U7862 (N_7862,N_5948,N_3381);
nor U7863 (N_7863,N_5020,N_3985);
or U7864 (N_7864,N_3492,N_5141);
and U7865 (N_7865,N_5370,N_3432);
and U7866 (N_7866,N_5049,N_4093);
nor U7867 (N_7867,N_3982,N_5773);
xnor U7868 (N_7868,N_5138,N_4284);
or U7869 (N_7869,N_3895,N_3896);
nor U7870 (N_7870,N_3735,N_3600);
and U7871 (N_7871,N_3093,N_5843);
xor U7872 (N_7872,N_3414,N_4342);
and U7873 (N_7873,N_5314,N_4043);
or U7874 (N_7874,N_5694,N_4781);
or U7875 (N_7875,N_3384,N_4070);
nor U7876 (N_7876,N_5568,N_3396);
nand U7877 (N_7877,N_5876,N_3996);
or U7878 (N_7878,N_3426,N_5567);
nor U7879 (N_7879,N_3664,N_5769);
and U7880 (N_7880,N_5649,N_3622);
and U7881 (N_7881,N_5719,N_4638);
nand U7882 (N_7882,N_4189,N_4480);
nand U7883 (N_7883,N_3038,N_3908);
and U7884 (N_7884,N_5296,N_5205);
and U7885 (N_7885,N_5967,N_5106);
nand U7886 (N_7886,N_5103,N_4460);
nor U7887 (N_7887,N_5599,N_4252);
and U7888 (N_7888,N_4506,N_3060);
nand U7889 (N_7889,N_3420,N_4661);
and U7890 (N_7890,N_3718,N_3272);
nor U7891 (N_7891,N_3474,N_5154);
xnor U7892 (N_7892,N_5883,N_5399);
nand U7893 (N_7893,N_4332,N_3607);
nand U7894 (N_7894,N_3309,N_3126);
nand U7895 (N_7895,N_5512,N_4796);
nor U7896 (N_7896,N_4414,N_5027);
or U7897 (N_7897,N_3240,N_5069);
and U7898 (N_7898,N_3398,N_4790);
nor U7899 (N_7899,N_4567,N_5694);
or U7900 (N_7900,N_5239,N_3383);
or U7901 (N_7901,N_5905,N_5853);
nor U7902 (N_7902,N_3688,N_3759);
nor U7903 (N_7903,N_4784,N_4801);
nand U7904 (N_7904,N_3554,N_4481);
nand U7905 (N_7905,N_4599,N_4942);
nand U7906 (N_7906,N_4779,N_5550);
nor U7907 (N_7907,N_3409,N_3885);
nand U7908 (N_7908,N_5962,N_5590);
or U7909 (N_7909,N_5693,N_5774);
or U7910 (N_7910,N_5391,N_3915);
and U7911 (N_7911,N_3448,N_3575);
nand U7912 (N_7912,N_4245,N_3345);
or U7913 (N_7913,N_5658,N_5416);
and U7914 (N_7914,N_5485,N_4510);
nand U7915 (N_7915,N_5351,N_3223);
nor U7916 (N_7916,N_3855,N_3871);
xnor U7917 (N_7917,N_5692,N_5072);
or U7918 (N_7918,N_4293,N_4385);
or U7919 (N_7919,N_3063,N_5021);
nor U7920 (N_7920,N_3563,N_4085);
and U7921 (N_7921,N_3569,N_5593);
nand U7922 (N_7922,N_3205,N_4778);
nor U7923 (N_7923,N_5995,N_3231);
or U7924 (N_7924,N_5686,N_5394);
or U7925 (N_7925,N_5274,N_3270);
and U7926 (N_7926,N_5313,N_5009);
nor U7927 (N_7927,N_3352,N_3933);
nand U7928 (N_7928,N_3780,N_3898);
and U7929 (N_7929,N_5301,N_5746);
nor U7930 (N_7930,N_3624,N_5030);
nand U7931 (N_7931,N_5232,N_4297);
nor U7932 (N_7932,N_5174,N_3245);
nor U7933 (N_7933,N_3906,N_3330);
and U7934 (N_7934,N_5918,N_3308);
nand U7935 (N_7935,N_5485,N_3308);
xor U7936 (N_7936,N_5798,N_3498);
nand U7937 (N_7937,N_4157,N_3483);
nor U7938 (N_7938,N_4586,N_3375);
and U7939 (N_7939,N_4897,N_3000);
nor U7940 (N_7940,N_5499,N_3185);
or U7941 (N_7941,N_4676,N_3807);
nand U7942 (N_7942,N_4999,N_4128);
nand U7943 (N_7943,N_3047,N_4144);
nand U7944 (N_7944,N_5729,N_3320);
nand U7945 (N_7945,N_4149,N_3620);
nor U7946 (N_7946,N_3297,N_5268);
nand U7947 (N_7947,N_4596,N_3679);
and U7948 (N_7948,N_5117,N_4856);
nor U7949 (N_7949,N_4687,N_4755);
nand U7950 (N_7950,N_4146,N_4654);
and U7951 (N_7951,N_5833,N_5600);
xor U7952 (N_7952,N_4961,N_5219);
and U7953 (N_7953,N_5561,N_5490);
nand U7954 (N_7954,N_4967,N_3050);
nor U7955 (N_7955,N_5775,N_5823);
and U7956 (N_7956,N_3410,N_3101);
nor U7957 (N_7957,N_4734,N_4191);
and U7958 (N_7958,N_3410,N_3197);
or U7959 (N_7959,N_4594,N_5100);
or U7960 (N_7960,N_3713,N_3234);
and U7961 (N_7961,N_4192,N_4929);
nor U7962 (N_7962,N_4194,N_3219);
and U7963 (N_7963,N_5344,N_5117);
nand U7964 (N_7964,N_4911,N_4649);
nand U7965 (N_7965,N_5259,N_5332);
nand U7966 (N_7966,N_3492,N_5388);
and U7967 (N_7967,N_3043,N_5014);
nor U7968 (N_7968,N_4146,N_4989);
nor U7969 (N_7969,N_3375,N_4570);
and U7970 (N_7970,N_5850,N_4600);
or U7971 (N_7971,N_4078,N_5620);
nor U7972 (N_7972,N_3791,N_5559);
or U7973 (N_7973,N_3266,N_5491);
and U7974 (N_7974,N_3527,N_4264);
nor U7975 (N_7975,N_5300,N_3444);
nand U7976 (N_7976,N_4586,N_4231);
nor U7977 (N_7977,N_3544,N_3048);
and U7978 (N_7978,N_3112,N_4685);
nor U7979 (N_7979,N_3209,N_4841);
nor U7980 (N_7980,N_4589,N_5012);
nand U7981 (N_7981,N_3126,N_5301);
and U7982 (N_7982,N_5170,N_4180);
nand U7983 (N_7983,N_3326,N_3019);
nand U7984 (N_7984,N_4418,N_3139);
nor U7985 (N_7985,N_5557,N_4201);
nor U7986 (N_7986,N_5722,N_5158);
or U7987 (N_7987,N_4869,N_5430);
and U7988 (N_7988,N_4382,N_5177);
nor U7989 (N_7989,N_4647,N_5034);
nand U7990 (N_7990,N_3985,N_3661);
and U7991 (N_7991,N_5456,N_5470);
nor U7992 (N_7992,N_5317,N_4641);
and U7993 (N_7993,N_3579,N_3094);
nor U7994 (N_7994,N_3431,N_4966);
nand U7995 (N_7995,N_3911,N_5255);
or U7996 (N_7996,N_4241,N_3256);
nor U7997 (N_7997,N_4805,N_3579);
nor U7998 (N_7998,N_4114,N_5910);
and U7999 (N_7999,N_3683,N_5618);
nor U8000 (N_8000,N_3561,N_5211);
nand U8001 (N_8001,N_3324,N_3034);
and U8002 (N_8002,N_3983,N_3565);
nand U8003 (N_8003,N_3365,N_5156);
or U8004 (N_8004,N_3384,N_4016);
nor U8005 (N_8005,N_4107,N_5216);
and U8006 (N_8006,N_3026,N_4991);
nand U8007 (N_8007,N_4285,N_4842);
nand U8008 (N_8008,N_3978,N_3154);
or U8009 (N_8009,N_3782,N_4490);
nand U8010 (N_8010,N_3575,N_3979);
nand U8011 (N_8011,N_3182,N_4502);
nor U8012 (N_8012,N_3698,N_3124);
xor U8013 (N_8013,N_3651,N_4906);
nand U8014 (N_8014,N_4891,N_3428);
nand U8015 (N_8015,N_3686,N_5585);
and U8016 (N_8016,N_5265,N_3404);
nor U8017 (N_8017,N_4898,N_5744);
nor U8018 (N_8018,N_3654,N_5230);
and U8019 (N_8019,N_3574,N_3251);
nor U8020 (N_8020,N_3622,N_5651);
and U8021 (N_8021,N_4405,N_4349);
or U8022 (N_8022,N_3064,N_5005);
or U8023 (N_8023,N_3184,N_3870);
or U8024 (N_8024,N_5615,N_4899);
nand U8025 (N_8025,N_3935,N_3377);
or U8026 (N_8026,N_5881,N_5777);
nand U8027 (N_8027,N_4372,N_4170);
nor U8028 (N_8028,N_3840,N_4161);
or U8029 (N_8029,N_4520,N_4476);
and U8030 (N_8030,N_5540,N_4231);
and U8031 (N_8031,N_4098,N_4373);
nand U8032 (N_8032,N_3183,N_4409);
nand U8033 (N_8033,N_3854,N_5188);
or U8034 (N_8034,N_3673,N_4359);
nand U8035 (N_8035,N_4819,N_3034);
or U8036 (N_8036,N_3870,N_4931);
or U8037 (N_8037,N_4566,N_3370);
nand U8038 (N_8038,N_5957,N_4651);
or U8039 (N_8039,N_5900,N_3035);
and U8040 (N_8040,N_4550,N_4486);
or U8041 (N_8041,N_4666,N_4652);
and U8042 (N_8042,N_4496,N_4905);
nand U8043 (N_8043,N_5503,N_3287);
nor U8044 (N_8044,N_4538,N_3693);
nor U8045 (N_8045,N_3862,N_4775);
and U8046 (N_8046,N_3907,N_5894);
nand U8047 (N_8047,N_3742,N_5433);
or U8048 (N_8048,N_4082,N_4989);
nor U8049 (N_8049,N_3171,N_4757);
nand U8050 (N_8050,N_3812,N_3223);
and U8051 (N_8051,N_5384,N_3162);
nor U8052 (N_8052,N_3191,N_5356);
and U8053 (N_8053,N_3211,N_3332);
nand U8054 (N_8054,N_3062,N_3239);
nand U8055 (N_8055,N_5044,N_4188);
and U8056 (N_8056,N_4260,N_4517);
nor U8057 (N_8057,N_3419,N_3059);
and U8058 (N_8058,N_4928,N_5273);
nor U8059 (N_8059,N_3404,N_5008);
nor U8060 (N_8060,N_3872,N_5369);
nor U8061 (N_8061,N_3811,N_5240);
and U8062 (N_8062,N_3856,N_4754);
and U8063 (N_8063,N_3892,N_4599);
and U8064 (N_8064,N_5350,N_3537);
nor U8065 (N_8065,N_3728,N_5016);
or U8066 (N_8066,N_5525,N_3086);
nor U8067 (N_8067,N_3058,N_3798);
and U8068 (N_8068,N_3267,N_5777);
nand U8069 (N_8069,N_5058,N_5830);
and U8070 (N_8070,N_3162,N_3205);
nor U8071 (N_8071,N_4608,N_4255);
nand U8072 (N_8072,N_4609,N_3719);
nor U8073 (N_8073,N_5845,N_3825);
nand U8074 (N_8074,N_5631,N_4738);
and U8075 (N_8075,N_5490,N_5387);
and U8076 (N_8076,N_5963,N_5836);
nand U8077 (N_8077,N_5083,N_3107);
and U8078 (N_8078,N_5291,N_3757);
or U8079 (N_8079,N_4383,N_4645);
nand U8080 (N_8080,N_5315,N_5569);
and U8081 (N_8081,N_3381,N_4514);
xor U8082 (N_8082,N_3861,N_3443);
nand U8083 (N_8083,N_5261,N_4627);
and U8084 (N_8084,N_5973,N_5845);
or U8085 (N_8085,N_3550,N_3255);
and U8086 (N_8086,N_4093,N_3782);
and U8087 (N_8087,N_3565,N_5260);
nor U8088 (N_8088,N_5299,N_4291);
nand U8089 (N_8089,N_3796,N_4838);
nand U8090 (N_8090,N_3897,N_3881);
and U8091 (N_8091,N_5396,N_5274);
and U8092 (N_8092,N_3927,N_3531);
nor U8093 (N_8093,N_3295,N_5987);
or U8094 (N_8094,N_5108,N_3757);
nor U8095 (N_8095,N_5336,N_5126);
nor U8096 (N_8096,N_4402,N_3314);
or U8097 (N_8097,N_3313,N_3788);
and U8098 (N_8098,N_3414,N_4069);
nor U8099 (N_8099,N_4369,N_5263);
and U8100 (N_8100,N_4451,N_3591);
and U8101 (N_8101,N_4431,N_4417);
and U8102 (N_8102,N_4760,N_3899);
nand U8103 (N_8103,N_3413,N_3041);
nor U8104 (N_8104,N_4379,N_5321);
nand U8105 (N_8105,N_3609,N_4880);
nand U8106 (N_8106,N_5902,N_4935);
or U8107 (N_8107,N_5800,N_5755);
and U8108 (N_8108,N_5063,N_3024);
or U8109 (N_8109,N_3121,N_3362);
and U8110 (N_8110,N_3106,N_3992);
nand U8111 (N_8111,N_5843,N_4674);
nand U8112 (N_8112,N_4776,N_5624);
or U8113 (N_8113,N_5140,N_4573);
or U8114 (N_8114,N_5484,N_4500);
nor U8115 (N_8115,N_5446,N_3196);
nor U8116 (N_8116,N_4166,N_4325);
and U8117 (N_8117,N_4742,N_3199);
or U8118 (N_8118,N_4309,N_5483);
nor U8119 (N_8119,N_5081,N_5999);
and U8120 (N_8120,N_3067,N_3561);
and U8121 (N_8121,N_5742,N_3854);
nand U8122 (N_8122,N_3832,N_4156);
nor U8123 (N_8123,N_4586,N_4577);
or U8124 (N_8124,N_4166,N_3105);
nor U8125 (N_8125,N_4587,N_3788);
nand U8126 (N_8126,N_3170,N_4646);
and U8127 (N_8127,N_4010,N_5242);
nor U8128 (N_8128,N_5381,N_3241);
and U8129 (N_8129,N_5275,N_3816);
and U8130 (N_8130,N_4163,N_4656);
nand U8131 (N_8131,N_4706,N_3656);
and U8132 (N_8132,N_3397,N_4120);
and U8133 (N_8133,N_5703,N_3640);
nor U8134 (N_8134,N_4607,N_4703);
or U8135 (N_8135,N_5603,N_4787);
and U8136 (N_8136,N_4008,N_3469);
nand U8137 (N_8137,N_3200,N_4319);
or U8138 (N_8138,N_3251,N_4473);
or U8139 (N_8139,N_4331,N_4968);
and U8140 (N_8140,N_4825,N_3419);
nand U8141 (N_8141,N_5811,N_5916);
nand U8142 (N_8142,N_3160,N_3012);
or U8143 (N_8143,N_5084,N_4834);
nand U8144 (N_8144,N_5020,N_3413);
or U8145 (N_8145,N_5555,N_4566);
or U8146 (N_8146,N_3837,N_4685);
or U8147 (N_8147,N_5863,N_4935);
or U8148 (N_8148,N_5931,N_5886);
or U8149 (N_8149,N_4591,N_3932);
and U8150 (N_8150,N_3153,N_3719);
nor U8151 (N_8151,N_4391,N_3140);
and U8152 (N_8152,N_4530,N_3785);
nand U8153 (N_8153,N_5537,N_5982);
nor U8154 (N_8154,N_5887,N_3941);
nand U8155 (N_8155,N_3561,N_3587);
and U8156 (N_8156,N_3492,N_4836);
nand U8157 (N_8157,N_4513,N_5895);
or U8158 (N_8158,N_5642,N_4880);
and U8159 (N_8159,N_3487,N_5375);
nand U8160 (N_8160,N_3410,N_3882);
nand U8161 (N_8161,N_3367,N_3139);
and U8162 (N_8162,N_4454,N_5708);
nor U8163 (N_8163,N_5350,N_4327);
or U8164 (N_8164,N_4644,N_4415);
nor U8165 (N_8165,N_5792,N_4253);
nand U8166 (N_8166,N_3815,N_4216);
nor U8167 (N_8167,N_5158,N_3216);
or U8168 (N_8168,N_4257,N_3807);
and U8169 (N_8169,N_5845,N_3929);
or U8170 (N_8170,N_4131,N_4004);
and U8171 (N_8171,N_3807,N_5013);
nor U8172 (N_8172,N_3986,N_3487);
nand U8173 (N_8173,N_4905,N_3093);
or U8174 (N_8174,N_4891,N_5200);
and U8175 (N_8175,N_4900,N_3195);
nor U8176 (N_8176,N_5595,N_4768);
nand U8177 (N_8177,N_4160,N_4091);
or U8178 (N_8178,N_4403,N_3212);
nor U8179 (N_8179,N_3211,N_5313);
and U8180 (N_8180,N_3751,N_5820);
and U8181 (N_8181,N_3392,N_5646);
nor U8182 (N_8182,N_3395,N_5480);
or U8183 (N_8183,N_3493,N_5364);
nand U8184 (N_8184,N_4031,N_4960);
and U8185 (N_8185,N_3952,N_3740);
nand U8186 (N_8186,N_3833,N_4865);
nor U8187 (N_8187,N_3139,N_5268);
xor U8188 (N_8188,N_4738,N_4574);
nand U8189 (N_8189,N_3439,N_4627);
nor U8190 (N_8190,N_3155,N_4629);
or U8191 (N_8191,N_4211,N_5870);
or U8192 (N_8192,N_3480,N_4031);
or U8193 (N_8193,N_3468,N_3815);
and U8194 (N_8194,N_4343,N_5153);
or U8195 (N_8195,N_5810,N_3537);
nand U8196 (N_8196,N_5417,N_5144);
nor U8197 (N_8197,N_5215,N_5653);
or U8198 (N_8198,N_5231,N_4690);
or U8199 (N_8199,N_4571,N_5760);
nor U8200 (N_8200,N_4501,N_4288);
nand U8201 (N_8201,N_3448,N_3665);
nand U8202 (N_8202,N_5229,N_4231);
and U8203 (N_8203,N_5551,N_4958);
or U8204 (N_8204,N_4972,N_5996);
and U8205 (N_8205,N_5585,N_3985);
and U8206 (N_8206,N_3670,N_3460);
and U8207 (N_8207,N_4600,N_5593);
nor U8208 (N_8208,N_4412,N_5464);
xor U8209 (N_8209,N_5404,N_5420);
nor U8210 (N_8210,N_3308,N_5256);
nor U8211 (N_8211,N_3308,N_3143);
and U8212 (N_8212,N_4005,N_5443);
nor U8213 (N_8213,N_5593,N_4939);
nand U8214 (N_8214,N_5865,N_4928);
or U8215 (N_8215,N_3608,N_4414);
nor U8216 (N_8216,N_3381,N_5459);
or U8217 (N_8217,N_3326,N_4659);
nand U8218 (N_8218,N_4993,N_3071);
nor U8219 (N_8219,N_5389,N_3837);
or U8220 (N_8220,N_5398,N_5368);
or U8221 (N_8221,N_5136,N_3578);
xnor U8222 (N_8222,N_3261,N_4070);
nand U8223 (N_8223,N_5662,N_4933);
or U8224 (N_8224,N_5796,N_5918);
nor U8225 (N_8225,N_3238,N_3656);
nor U8226 (N_8226,N_5761,N_3121);
nand U8227 (N_8227,N_3371,N_4213);
nand U8228 (N_8228,N_3463,N_5026);
nand U8229 (N_8229,N_3396,N_3569);
nand U8230 (N_8230,N_5747,N_5402);
and U8231 (N_8231,N_5472,N_3783);
or U8232 (N_8232,N_4711,N_4863);
and U8233 (N_8233,N_5109,N_3433);
nor U8234 (N_8234,N_3170,N_5352);
and U8235 (N_8235,N_5532,N_4541);
or U8236 (N_8236,N_5351,N_3024);
or U8237 (N_8237,N_5194,N_5252);
nor U8238 (N_8238,N_5823,N_3817);
nand U8239 (N_8239,N_3530,N_3519);
or U8240 (N_8240,N_3047,N_4759);
or U8241 (N_8241,N_5981,N_4998);
and U8242 (N_8242,N_5172,N_3217);
xnor U8243 (N_8243,N_4284,N_3195);
or U8244 (N_8244,N_4111,N_5592);
nor U8245 (N_8245,N_4710,N_3270);
and U8246 (N_8246,N_4240,N_3224);
or U8247 (N_8247,N_4441,N_5744);
and U8248 (N_8248,N_4972,N_5861);
and U8249 (N_8249,N_4952,N_5481);
nor U8250 (N_8250,N_5138,N_4101);
or U8251 (N_8251,N_4544,N_4811);
nor U8252 (N_8252,N_3558,N_3646);
and U8253 (N_8253,N_3473,N_4681);
and U8254 (N_8254,N_3277,N_4699);
nand U8255 (N_8255,N_3903,N_5996);
nand U8256 (N_8256,N_3118,N_4808);
or U8257 (N_8257,N_4697,N_5336);
and U8258 (N_8258,N_3015,N_3776);
and U8259 (N_8259,N_5871,N_5894);
and U8260 (N_8260,N_5737,N_5844);
nor U8261 (N_8261,N_3016,N_4170);
nor U8262 (N_8262,N_3490,N_5390);
and U8263 (N_8263,N_5412,N_5437);
nand U8264 (N_8264,N_5160,N_5081);
or U8265 (N_8265,N_3886,N_4087);
nor U8266 (N_8266,N_3727,N_3217);
nand U8267 (N_8267,N_5998,N_3009);
nor U8268 (N_8268,N_3649,N_5820);
and U8269 (N_8269,N_5870,N_4036);
nor U8270 (N_8270,N_4211,N_3986);
nand U8271 (N_8271,N_3525,N_5683);
nor U8272 (N_8272,N_4580,N_4990);
or U8273 (N_8273,N_5831,N_5215);
or U8274 (N_8274,N_5602,N_4432);
and U8275 (N_8275,N_4701,N_3093);
nor U8276 (N_8276,N_4594,N_4297);
and U8277 (N_8277,N_4539,N_4121);
nand U8278 (N_8278,N_3986,N_4536);
or U8279 (N_8279,N_5138,N_3487);
nand U8280 (N_8280,N_3991,N_5322);
and U8281 (N_8281,N_4895,N_4225);
nor U8282 (N_8282,N_5765,N_4151);
nor U8283 (N_8283,N_3287,N_4843);
nand U8284 (N_8284,N_3617,N_4568);
or U8285 (N_8285,N_5604,N_4539);
nor U8286 (N_8286,N_4035,N_3985);
nor U8287 (N_8287,N_5369,N_3997);
or U8288 (N_8288,N_4211,N_5536);
nor U8289 (N_8289,N_5407,N_5769);
nand U8290 (N_8290,N_5257,N_3810);
nand U8291 (N_8291,N_3225,N_5744);
or U8292 (N_8292,N_3159,N_4549);
nand U8293 (N_8293,N_3472,N_4829);
nand U8294 (N_8294,N_3227,N_5003);
and U8295 (N_8295,N_3372,N_3793);
and U8296 (N_8296,N_3153,N_5392);
or U8297 (N_8297,N_5775,N_3653);
and U8298 (N_8298,N_4389,N_4687);
nor U8299 (N_8299,N_4347,N_5681);
nand U8300 (N_8300,N_3649,N_4127);
or U8301 (N_8301,N_4415,N_3928);
nand U8302 (N_8302,N_5002,N_4375);
nor U8303 (N_8303,N_3896,N_3245);
and U8304 (N_8304,N_4420,N_4697);
or U8305 (N_8305,N_4508,N_4958);
and U8306 (N_8306,N_4919,N_4966);
nand U8307 (N_8307,N_4839,N_4345);
and U8308 (N_8308,N_3111,N_3259);
or U8309 (N_8309,N_5206,N_5385);
or U8310 (N_8310,N_4816,N_5385);
and U8311 (N_8311,N_3603,N_5068);
or U8312 (N_8312,N_4535,N_3498);
and U8313 (N_8313,N_5579,N_4732);
and U8314 (N_8314,N_5932,N_3291);
and U8315 (N_8315,N_4571,N_5775);
or U8316 (N_8316,N_4160,N_3443);
nand U8317 (N_8317,N_3278,N_3155);
nand U8318 (N_8318,N_3254,N_4511);
or U8319 (N_8319,N_5288,N_3122);
nand U8320 (N_8320,N_5785,N_4185);
nor U8321 (N_8321,N_3977,N_4495);
nor U8322 (N_8322,N_4516,N_3966);
nor U8323 (N_8323,N_3146,N_3465);
or U8324 (N_8324,N_4220,N_5994);
nor U8325 (N_8325,N_5751,N_3855);
nor U8326 (N_8326,N_3854,N_3087);
and U8327 (N_8327,N_3077,N_3822);
and U8328 (N_8328,N_5185,N_5464);
and U8329 (N_8329,N_4483,N_5697);
nor U8330 (N_8330,N_5320,N_5143);
nand U8331 (N_8331,N_5568,N_4906);
and U8332 (N_8332,N_5875,N_3195);
or U8333 (N_8333,N_4368,N_4513);
and U8334 (N_8334,N_4997,N_4811);
or U8335 (N_8335,N_5617,N_5243);
or U8336 (N_8336,N_3303,N_3243);
or U8337 (N_8337,N_4399,N_5484);
nand U8338 (N_8338,N_4390,N_4201);
nor U8339 (N_8339,N_3759,N_5201);
or U8340 (N_8340,N_5516,N_5857);
nor U8341 (N_8341,N_5527,N_4044);
and U8342 (N_8342,N_5364,N_3820);
and U8343 (N_8343,N_5214,N_4746);
or U8344 (N_8344,N_5598,N_3784);
xor U8345 (N_8345,N_3714,N_5422);
or U8346 (N_8346,N_5508,N_4573);
and U8347 (N_8347,N_5618,N_3983);
nor U8348 (N_8348,N_3527,N_4855);
and U8349 (N_8349,N_5406,N_4266);
nand U8350 (N_8350,N_3792,N_5117);
nor U8351 (N_8351,N_5954,N_3401);
or U8352 (N_8352,N_3650,N_4916);
and U8353 (N_8353,N_4295,N_3786);
nand U8354 (N_8354,N_4989,N_5953);
nor U8355 (N_8355,N_3645,N_4997);
or U8356 (N_8356,N_5935,N_4250);
nand U8357 (N_8357,N_3220,N_4622);
and U8358 (N_8358,N_3369,N_4894);
or U8359 (N_8359,N_4511,N_3424);
nor U8360 (N_8360,N_4389,N_4744);
nor U8361 (N_8361,N_5930,N_3597);
xnor U8362 (N_8362,N_3971,N_5430);
or U8363 (N_8363,N_3513,N_3350);
and U8364 (N_8364,N_5190,N_4694);
or U8365 (N_8365,N_3711,N_5575);
and U8366 (N_8366,N_3273,N_4594);
nor U8367 (N_8367,N_4889,N_3788);
and U8368 (N_8368,N_4667,N_4298);
and U8369 (N_8369,N_5145,N_4897);
or U8370 (N_8370,N_3972,N_3686);
nor U8371 (N_8371,N_3286,N_4577);
or U8372 (N_8372,N_4571,N_3340);
nand U8373 (N_8373,N_5863,N_4294);
and U8374 (N_8374,N_3626,N_5432);
or U8375 (N_8375,N_3025,N_5615);
nor U8376 (N_8376,N_4331,N_4261);
nand U8377 (N_8377,N_4071,N_4813);
or U8378 (N_8378,N_4897,N_3303);
or U8379 (N_8379,N_4945,N_5496);
xor U8380 (N_8380,N_3558,N_5905);
and U8381 (N_8381,N_4179,N_3892);
or U8382 (N_8382,N_5767,N_5315);
or U8383 (N_8383,N_5444,N_3101);
or U8384 (N_8384,N_5076,N_3083);
nor U8385 (N_8385,N_4352,N_5694);
or U8386 (N_8386,N_5930,N_4732);
or U8387 (N_8387,N_4620,N_5262);
nor U8388 (N_8388,N_5764,N_4239);
and U8389 (N_8389,N_4043,N_4694);
or U8390 (N_8390,N_3013,N_3137);
nand U8391 (N_8391,N_3051,N_3566);
nand U8392 (N_8392,N_3415,N_5233);
or U8393 (N_8393,N_5749,N_3733);
nor U8394 (N_8394,N_4777,N_3341);
nand U8395 (N_8395,N_3772,N_4551);
and U8396 (N_8396,N_4602,N_4015);
and U8397 (N_8397,N_4292,N_3171);
nand U8398 (N_8398,N_3309,N_5641);
nor U8399 (N_8399,N_5690,N_5956);
nor U8400 (N_8400,N_5041,N_3147);
nor U8401 (N_8401,N_3023,N_5565);
nand U8402 (N_8402,N_4622,N_4612);
nor U8403 (N_8403,N_4930,N_3481);
nand U8404 (N_8404,N_4883,N_5055);
or U8405 (N_8405,N_3322,N_3407);
xor U8406 (N_8406,N_5602,N_4792);
nor U8407 (N_8407,N_4463,N_5637);
nand U8408 (N_8408,N_5858,N_3495);
nand U8409 (N_8409,N_4385,N_5866);
or U8410 (N_8410,N_5161,N_3324);
nand U8411 (N_8411,N_3795,N_3341);
nor U8412 (N_8412,N_3143,N_5302);
and U8413 (N_8413,N_5386,N_3216);
or U8414 (N_8414,N_5055,N_5635);
or U8415 (N_8415,N_3782,N_5738);
nand U8416 (N_8416,N_3581,N_5280);
and U8417 (N_8417,N_5260,N_5974);
or U8418 (N_8418,N_4066,N_3717);
nand U8419 (N_8419,N_3501,N_3195);
nand U8420 (N_8420,N_5984,N_4177);
nor U8421 (N_8421,N_4151,N_5473);
nand U8422 (N_8422,N_5259,N_4330);
nand U8423 (N_8423,N_3130,N_4065);
and U8424 (N_8424,N_3550,N_3289);
nand U8425 (N_8425,N_3213,N_5108);
nor U8426 (N_8426,N_4480,N_3530);
nand U8427 (N_8427,N_3188,N_4334);
and U8428 (N_8428,N_3002,N_4055);
and U8429 (N_8429,N_5149,N_5950);
nor U8430 (N_8430,N_3136,N_5450);
or U8431 (N_8431,N_4860,N_3455);
or U8432 (N_8432,N_5179,N_5047);
nand U8433 (N_8433,N_5364,N_3276);
or U8434 (N_8434,N_4491,N_4059);
and U8435 (N_8435,N_4233,N_4431);
nor U8436 (N_8436,N_4997,N_4485);
or U8437 (N_8437,N_4119,N_3214);
nor U8438 (N_8438,N_5328,N_3159);
or U8439 (N_8439,N_3466,N_5646);
nor U8440 (N_8440,N_3261,N_5978);
and U8441 (N_8441,N_4660,N_4274);
or U8442 (N_8442,N_4779,N_4550);
nand U8443 (N_8443,N_3890,N_5392);
and U8444 (N_8444,N_4337,N_4715);
or U8445 (N_8445,N_4393,N_4320);
and U8446 (N_8446,N_5167,N_3837);
or U8447 (N_8447,N_4724,N_4876);
or U8448 (N_8448,N_4011,N_3825);
nand U8449 (N_8449,N_5093,N_5042);
and U8450 (N_8450,N_4204,N_3369);
nor U8451 (N_8451,N_4391,N_3735);
xor U8452 (N_8452,N_5033,N_4431);
or U8453 (N_8453,N_4320,N_3743);
or U8454 (N_8454,N_4485,N_3395);
or U8455 (N_8455,N_4845,N_3772);
nor U8456 (N_8456,N_5809,N_3865);
nor U8457 (N_8457,N_5746,N_4750);
nor U8458 (N_8458,N_4753,N_4347);
or U8459 (N_8459,N_4301,N_4903);
and U8460 (N_8460,N_3959,N_3956);
and U8461 (N_8461,N_4415,N_4848);
or U8462 (N_8462,N_4515,N_3278);
or U8463 (N_8463,N_3100,N_4677);
and U8464 (N_8464,N_5552,N_4237);
or U8465 (N_8465,N_4867,N_4839);
nand U8466 (N_8466,N_5898,N_4383);
nand U8467 (N_8467,N_5791,N_5964);
nand U8468 (N_8468,N_4170,N_4951);
or U8469 (N_8469,N_4999,N_4709);
or U8470 (N_8470,N_3059,N_4693);
xor U8471 (N_8471,N_4679,N_3017);
and U8472 (N_8472,N_4551,N_3563);
or U8473 (N_8473,N_3976,N_4898);
and U8474 (N_8474,N_3134,N_5087);
nor U8475 (N_8475,N_3354,N_3271);
nor U8476 (N_8476,N_3325,N_5047);
nand U8477 (N_8477,N_5875,N_4718);
or U8478 (N_8478,N_5947,N_4915);
or U8479 (N_8479,N_5314,N_5878);
or U8480 (N_8480,N_5927,N_4290);
nor U8481 (N_8481,N_4628,N_4999);
and U8482 (N_8482,N_3995,N_4853);
nand U8483 (N_8483,N_5177,N_5112);
or U8484 (N_8484,N_5542,N_5514);
nand U8485 (N_8485,N_5648,N_5877);
or U8486 (N_8486,N_3532,N_3477);
nand U8487 (N_8487,N_5388,N_4826);
nor U8488 (N_8488,N_4082,N_4391);
or U8489 (N_8489,N_3073,N_3010);
nor U8490 (N_8490,N_3145,N_5580);
nor U8491 (N_8491,N_5413,N_3654);
and U8492 (N_8492,N_5074,N_4724);
nor U8493 (N_8493,N_5118,N_5422);
nand U8494 (N_8494,N_3337,N_4459);
nor U8495 (N_8495,N_5343,N_3421);
nor U8496 (N_8496,N_5853,N_4691);
nand U8497 (N_8497,N_3554,N_4083);
nor U8498 (N_8498,N_3159,N_5693);
nor U8499 (N_8499,N_4870,N_3088);
or U8500 (N_8500,N_4215,N_4827);
nor U8501 (N_8501,N_5486,N_4220);
or U8502 (N_8502,N_5673,N_4668);
nor U8503 (N_8503,N_3938,N_5799);
nor U8504 (N_8504,N_3297,N_3997);
nand U8505 (N_8505,N_3489,N_5504);
or U8506 (N_8506,N_3228,N_3543);
nor U8507 (N_8507,N_4773,N_5365);
nor U8508 (N_8508,N_5285,N_5582);
and U8509 (N_8509,N_3586,N_3998);
and U8510 (N_8510,N_4839,N_3404);
nand U8511 (N_8511,N_5499,N_5871);
nor U8512 (N_8512,N_4231,N_4148);
or U8513 (N_8513,N_4828,N_5479);
nor U8514 (N_8514,N_4477,N_5703);
and U8515 (N_8515,N_4891,N_4804);
or U8516 (N_8516,N_4475,N_4048);
or U8517 (N_8517,N_3874,N_5302);
nor U8518 (N_8518,N_3203,N_4861);
nor U8519 (N_8519,N_4519,N_4886);
or U8520 (N_8520,N_4086,N_3315);
nor U8521 (N_8521,N_3443,N_5718);
xor U8522 (N_8522,N_5726,N_3212);
or U8523 (N_8523,N_5281,N_4117);
or U8524 (N_8524,N_4889,N_3490);
nand U8525 (N_8525,N_5298,N_4971);
nor U8526 (N_8526,N_3335,N_3283);
and U8527 (N_8527,N_3567,N_5701);
nand U8528 (N_8528,N_4853,N_5336);
nand U8529 (N_8529,N_5969,N_3669);
and U8530 (N_8530,N_4421,N_3489);
or U8531 (N_8531,N_4309,N_3175);
nor U8532 (N_8532,N_4423,N_5056);
nor U8533 (N_8533,N_5403,N_3462);
or U8534 (N_8534,N_5840,N_4744);
and U8535 (N_8535,N_5653,N_4033);
and U8536 (N_8536,N_4401,N_5903);
and U8537 (N_8537,N_3014,N_4412);
or U8538 (N_8538,N_5453,N_4943);
nor U8539 (N_8539,N_4446,N_4300);
nand U8540 (N_8540,N_4107,N_4004);
nor U8541 (N_8541,N_3477,N_4077);
or U8542 (N_8542,N_5195,N_5197);
nor U8543 (N_8543,N_3263,N_4694);
nand U8544 (N_8544,N_4668,N_3455);
nand U8545 (N_8545,N_5523,N_3992);
nor U8546 (N_8546,N_3337,N_4932);
or U8547 (N_8547,N_5970,N_5892);
nor U8548 (N_8548,N_5532,N_3290);
and U8549 (N_8549,N_5155,N_3728);
or U8550 (N_8550,N_4687,N_3653);
nand U8551 (N_8551,N_5843,N_5539);
nand U8552 (N_8552,N_3281,N_3729);
or U8553 (N_8553,N_5974,N_5177);
and U8554 (N_8554,N_5334,N_5813);
nand U8555 (N_8555,N_3415,N_3129);
and U8556 (N_8556,N_4588,N_4999);
and U8557 (N_8557,N_5243,N_3431);
nand U8558 (N_8558,N_4922,N_3408);
and U8559 (N_8559,N_5170,N_5510);
nor U8560 (N_8560,N_4921,N_5169);
nand U8561 (N_8561,N_4529,N_5587);
nor U8562 (N_8562,N_4075,N_3311);
or U8563 (N_8563,N_4436,N_3031);
or U8564 (N_8564,N_3509,N_4807);
nand U8565 (N_8565,N_4975,N_4208);
nor U8566 (N_8566,N_5148,N_5076);
nor U8567 (N_8567,N_4933,N_5913);
or U8568 (N_8568,N_5583,N_4421);
and U8569 (N_8569,N_3974,N_3644);
and U8570 (N_8570,N_5782,N_5450);
or U8571 (N_8571,N_5278,N_5083);
nor U8572 (N_8572,N_3417,N_4548);
and U8573 (N_8573,N_3930,N_3742);
nand U8574 (N_8574,N_4497,N_5360);
and U8575 (N_8575,N_5385,N_4854);
or U8576 (N_8576,N_3301,N_4586);
xnor U8577 (N_8577,N_5383,N_3804);
xor U8578 (N_8578,N_5888,N_3978);
nand U8579 (N_8579,N_4993,N_3079);
or U8580 (N_8580,N_5340,N_3968);
or U8581 (N_8581,N_4681,N_3487);
nor U8582 (N_8582,N_4485,N_3088);
and U8583 (N_8583,N_5143,N_4869);
nor U8584 (N_8584,N_4099,N_4987);
nand U8585 (N_8585,N_5037,N_5602);
nor U8586 (N_8586,N_5257,N_4462);
and U8587 (N_8587,N_3252,N_5573);
nor U8588 (N_8588,N_5404,N_3576);
and U8589 (N_8589,N_3948,N_3647);
nand U8590 (N_8590,N_4281,N_3852);
nand U8591 (N_8591,N_4151,N_4462);
nand U8592 (N_8592,N_4261,N_5470);
and U8593 (N_8593,N_4319,N_3408);
nand U8594 (N_8594,N_4059,N_4895);
nor U8595 (N_8595,N_5153,N_3657);
and U8596 (N_8596,N_5700,N_3802);
nand U8597 (N_8597,N_5211,N_5611);
and U8598 (N_8598,N_4890,N_3958);
or U8599 (N_8599,N_4469,N_5603);
or U8600 (N_8600,N_3533,N_5741);
and U8601 (N_8601,N_4963,N_4458);
or U8602 (N_8602,N_3023,N_3479);
nor U8603 (N_8603,N_5815,N_3818);
nor U8604 (N_8604,N_4566,N_5832);
or U8605 (N_8605,N_5581,N_3117);
nand U8606 (N_8606,N_3205,N_5832);
or U8607 (N_8607,N_3026,N_3818);
nor U8608 (N_8608,N_3272,N_3463);
and U8609 (N_8609,N_4179,N_4621);
nand U8610 (N_8610,N_5763,N_3051);
and U8611 (N_8611,N_3192,N_4338);
xnor U8612 (N_8612,N_3711,N_3580);
nand U8613 (N_8613,N_5065,N_4179);
and U8614 (N_8614,N_5686,N_4872);
or U8615 (N_8615,N_3338,N_5890);
or U8616 (N_8616,N_4749,N_4658);
or U8617 (N_8617,N_4637,N_5373);
and U8618 (N_8618,N_3228,N_3796);
and U8619 (N_8619,N_3133,N_4483);
and U8620 (N_8620,N_3280,N_3968);
nor U8621 (N_8621,N_3483,N_5304);
nor U8622 (N_8622,N_5142,N_4260);
nor U8623 (N_8623,N_4923,N_5931);
and U8624 (N_8624,N_5011,N_5721);
nand U8625 (N_8625,N_5386,N_4563);
and U8626 (N_8626,N_5552,N_5725);
nand U8627 (N_8627,N_4273,N_4278);
or U8628 (N_8628,N_5740,N_4436);
nor U8629 (N_8629,N_5832,N_5624);
and U8630 (N_8630,N_3568,N_3860);
or U8631 (N_8631,N_5474,N_3967);
nor U8632 (N_8632,N_4778,N_3402);
nand U8633 (N_8633,N_4050,N_5590);
or U8634 (N_8634,N_3191,N_5732);
nand U8635 (N_8635,N_3526,N_3573);
nor U8636 (N_8636,N_3017,N_5459);
and U8637 (N_8637,N_4813,N_5328);
nand U8638 (N_8638,N_4931,N_4661);
nor U8639 (N_8639,N_4861,N_4457);
or U8640 (N_8640,N_4753,N_5318);
nor U8641 (N_8641,N_3012,N_3427);
nand U8642 (N_8642,N_3607,N_4610);
and U8643 (N_8643,N_5217,N_4662);
nor U8644 (N_8644,N_4945,N_3581);
nor U8645 (N_8645,N_4360,N_4775);
nor U8646 (N_8646,N_5747,N_3798);
or U8647 (N_8647,N_5903,N_4676);
nor U8648 (N_8648,N_5682,N_3310);
nor U8649 (N_8649,N_4500,N_5853);
or U8650 (N_8650,N_3416,N_5182);
or U8651 (N_8651,N_3331,N_3397);
nor U8652 (N_8652,N_4125,N_5135);
nand U8653 (N_8653,N_4645,N_3541);
nand U8654 (N_8654,N_3764,N_4134);
nor U8655 (N_8655,N_4727,N_5353);
and U8656 (N_8656,N_3462,N_5444);
or U8657 (N_8657,N_4610,N_5294);
or U8658 (N_8658,N_4965,N_3236);
nor U8659 (N_8659,N_4656,N_4968);
or U8660 (N_8660,N_3187,N_4650);
nor U8661 (N_8661,N_4924,N_5219);
and U8662 (N_8662,N_4801,N_5670);
or U8663 (N_8663,N_5551,N_5706);
and U8664 (N_8664,N_3406,N_3908);
and U8665 (N_8665,N_3661,N_5864);
nand U8666 (N_8666,N_3993,N_3755);
nand U8667 (N_8667,N_5002,N_4134);
and U8668 (N_8668,N_5249,N_4763);
or U8669 (N_8669,N_3573,N_5218);
nand U8670 (N_8670,N_3213,N_3519);
nor U8671 (N_8671,N_5283,N_5130);
nor U8672 (N_8672,N_3723,N_3868);
nor U8673 (N_8673,N_3218,N_4890);
nand U8674 (N_8674,N_4380,N_4520);
nor U8675 (N_8675,N_3592,N_3499);
and U8676 (N_8676,N_3593,N_3821);
nor U8677 (N_8677,N_4879,N_4422);
and U8678 (N_8678,N_4424,N_3270);
and U8679 (N_8679,N_4913,N_3552);
or U8680 (N_8680,N_3726,N_4400);
nor U8681 (N_8681,N_4429,N_4916);
or U8682 (N_8682,N_5946,N_4175);
nand U8683 (N_8683,N_5680,N_4573);
nor U8684 (N_8684,N_5840,N_5700);
nor U8685 (N_8685,N_3260,N_3621);
or U8686 (N_8686,N_4569,N_3241);
and U8687 (N_8687,N_4736,N_5294);
nor U8688 (N_8688,N_3702,N_3195);
nor U8689 (N_8689,N_5765,N_5169);
and U8690 (N_8690,N_4163,N_4497);
nor U8691 (N_8691,N_5221,N_3675);
or U8692 (N_8692,N_3121,N_5049);
or U8693 (N_8693,N_5312,N_3597);
and U8694 (N_8694,N_3346,N_4809);
nor U8695 (N_8695,N_5653,N_3634);
nor U8696 (N_8696,N_5636,N_5341);
nand U8697 (N_8697,N_4842,N_4615);
and U8698 (N_8698,N_3695,N_5162);
nor U8699 (N_8699,N_5275,N_5238);
xnor U8700 (N_8700,N_4655,N_3472);
nor U8701 (N_8701,N_3316,N_3892);
or U8702 (N_8702,N_3923,N_4907);
nor U8703 (N_8703,N_4298,N_3088);
or U8704 (N_8704,N_4486,N_3980);
nand U8705 (N_8705,N_3668,N_4865);
nor U8706 (N_8706,N_3203,N_4429);
nand U8707 (N_8707,N_4943,N_3446);
nor U8708 (N_8708,N_4720,N_3541);
or U8709 (N_8709,N_5412,N_5395);
and U8710 (N_8710,N_5662,N_5786);
and U8711 (N_8711,N_5330,N_3153);
or U8712 (N_8712,N_3025,N_3448);
or U8713 (N_8713,N_3240,N_4808);
or U8714 (N_8714,N_5089,N_5887);
or U8715 (N_8715,N_4735,N_4027);
nor U8716 (N_8716,N_3608,N_3709);
or U8717 (N_8717,N_3266,N_4019);
or U8718 (N_8718,N_4739,N_5366);
and U8719 (N_8719,N_3075,N_4975);
or U8720 (N_8720,N_3340,N_4933);
nand U8721 (N_8721,N_5313,N_3472);
nor U8722 (N_8722,N_4666,N_3463);
nand U8723 (N_8723,N_3086,N_3799);
nor U8724 (N_8724,N_4964,N_5817);
nor U8725 (N_8725,N_4803,N_5724);
or U8726 (N_8726,N_3049,N_3386);
nor U8727 (N_8727,N_4908,N_3362);
and U8728 (N_8728,N_5400,N_3105);
and U8729 (N_8729,N_4614,N_4057);
nand U8730 (N_8730,N_4882,N_3683);
and U8731 (N_8731,N_5896,N_3034);
and U8732 (N_8732,N_3531,N_4948);
nand U8733 (N_8733,N_4401,N_4701);
nor U8734 (N_8734,N_5334,N_5468);
nand U8735 (N_8735,N_4409,N_3832);
or U8736 (N_8736,N_4482,N_4286);
nand U8737 (N_8737,N_3636,N_5393);
nor U8738 (N_8738,N_4989,N_4118);
or U8739 (N_8739,N_4721,N_4285);
nand U8740 (N_8740,N_4651,N_4871);
and U8741 (N_8741,N_4809,N_5229);
and U8742 (N_8742,N_4780,N_3347);
nor U8743 (N_8743,N_3289,N_5176);
nor U8744 (N_8744,N_5797,N_4128);
or U8745 (N_8745,N_5561,N_3961);
and U8746 (N_8746,N_4343,N_5883);
nand U8747 (N_8747,N_3229,N_3301);
nand U8748 (N_8748,N_4822,N_4481);
or U8749 (N_8749,N_5234,N_5913);
and U8750 (N_8750,N_3974,N_5077);
and U8751 (N_8751,N_5660,N_4200);
and U8752 (N_8752,N_4408,N_5362);
and U8753 (N_8753,N_5727,N_3897);
nand U8754 (N_8754,N_5331,N_5269);
or U8755 (N_8755,N_4729,N_5346);
nand U8756 (N_8756,N_4681,N_5513);
nor U8757 (N_8757,N_4848,N_3916);
nor U8758 (N_8758,N_5977,N_5273);
nand U8759 (N_8759,N_3431,N_4538);
nor U8760 (N_8760,N_4697,N_3232);
and U8761 (N_8761,N_3883,N_3702);
and U8762 (N_8762,N_3663,N_5101);
or U8763 (N_8763,N_4049,N_5724);
and U8764 (N_8764,N_4130,N_4354);
nor U8765 (N_8765,N_3565,N_4393);
and U8766 (N_8766,N_3451,N_4861);
and U8767 (N_8767,N_3459,N_5647);
and U8768 (N_8768,N_4515,N_3585);
nor U8769 (N_8769,N_4922,N_4736);
or U8770 (N_8770,N_3557,N_5466);
or U8771 (N_8771,N_4909,N_4673);
nor U8772 (N_8772,N_4620,N_3473);
and U8773 (N_8773,N_4239,N_3685);
nor U8774 (N_8774,N_5190,N_4422);
nand U8775 (N_8775,N_4316,N_4499);
nand U8776 (N_8776,N_4066,N_3727);
nand U8777 (N_8777,N_5482,N_3550);
nor U8778 (N_8778,N_3275,N_5356);
nand U8779 (N_8779,N_3665,N_5712);
and U8780 (N_8780,N_5592,N_4984);
or U8781 (N_8781,N_3355,N_4753);
or U8782 (N_8782,N_3611,N_3288);
nor U8783 (N_8783,N_4705,N_5575);
or U8784 (N_8784,N_5799,N_3914);
and U8785 (N_8785,N_3975,N_5930);
nor U8786 (N_8786,N_4491,N_4102);
nor U8787 (N_8787,N_5108,N_4730);
nand U8788 (N_8788,N_5137,N_3182);
nor U8789 (N_8789,N_4973,N_3959);
or U8790 (N_8790,N_5847,N_3117);
or U8791 (N_8791,N_5305,N_5773);
nor U8792 (N_8792,N_5328,N_3281);
and U8793 (N_8793,N_4747,N_4655);
nor U8794 (N_8794,N_5244,N_4760);
nor U8795 (N_8795,N_3456,N_3549);
nand U8796 (N_8796,N_5163,N_4094);
or U8797 (N_8797,N_4731,N_4798);
or U8798 (N_8798,N_5052,N_4594);
or U8799 (N_8799,N_5100,N_4644);
or U8800 (N_8800,N_5601,N_5224);
and U8801 (N_8801,N_4134,N_4000);
and U8802 (N_8802,N_4207,N_3270);
nor U8803 (N_8803,N_3669,N_4486);
nand U8804 (N_8804,N_5726,N_3676);
or U8805 (N_8805,N_4577,N_4954);
nor U8806 (N_8806,N_4690,N_5772);
nor U8807 (N_8807,N_4506,N_4756);
or U8808 (N_8808,N_3981,N_3951);
and U8809 (N_8809,N_4205,N_3335);
nand U8810 (N_8810,N_4962,N_4344);
and U8811 (N_8811,N_4563,N_5086);
and U8812 (N_8812,N_5602,N_4129);
and U8813 (N_8813,N_4078,N_3512);
nand U8814 (N_8814,N_3521,N_5333);
and U8815 (N_8815,N_5267,N_3285);
nand U8816 (N_8816,N_4576,N_5212);
nand U8817 (N_8817,N_4375,N_3022);
nor U8818 (N_8818,N_4115,N_5847);
nor U8819 (N_8819,N_3295,N_3862);
nand U8820 (N_8820,N_3908,N_4137);
or U8821 (N_8821,N_3255,N_5626);
and U8822 (N_8822,N_4436,N_4194);
nor U8823 (N_8823,N_5400,N_3630);
or U8824 (N_8824,N_4705,N_5234);
nand U8825 (N_8825,N_5422,N_3984);
nand U8826 (N_8826,N_3069,N_3166);
nor U8827 (N_8827,N_3822,N_5888);
and U8828 (N_8828,N_3406,N_4019);
or U8829 (N_8829,N_4084,N_3235);
and U8830 (N_8830,N_5322,N_3446);
nand U8831 (N_8831,N_5995,N_4408);
nand U8832 (N_8832,N_3487,N_5840);
nor U8833 (N_8833,N_5668,N_3487);
nand U8834 (N_8834,N_5718,N_5081);
nand U8835 (N_8835,N_3368,N_4385);
nor U8836 (N_8836,N_3170,N_4847);
nor U8837 (N_8837,N_4396,N_3643);
nor U8838 (N_8838,N_3164,N_4575);
nor U8839 (N_8839,N_5008,N_4194);
nor U8840 (N_8840,N_3245,N_5653);
or U8841 (N_8841,N_4836,N_5607);
and U8842 (N_8842,N_3126,N_5941);
or U8843 (N_8843,N_4717,N_4039);
nand U8844 (N_8844,N_4901,N_5558);
or U8845 (N_8845,N_5259,N_3320);
nor U8846 (N_8846,N_5445,N_3624);
nor U8847 (N_8847,N_3005,N_4212);
nand U8848 (N_8848,N_3540,N_3335);
nor U8849 (N_8849,N_4258,N_5963);
nor U8850 (N_8850,N_3407,N_4205);
nor U8851 (N_8851,N_5792,N_3552);
nand U8852 (N_8852,N_3332,N_4057);
nand U8853 (N_8853,N_4255,N_3442);
and U8854 (N_8854,N_5420,N_4652);
or U8855 (N_8855,N_5246,N_5655);
and U8856 (N_8856,N_5403,N_3910);
and U8857 (N_8857,N_4703,N_3219);
nor U8858 (N_8858,N_5916,N_3133);
nor U8859 (N_8859,N_3228,N_3126);
or U8860 (N_8860,N_5559,N_3016);
nand U8861 (N_8861,N_4282,N_3881);
and U8862 (N_8862,N_5428,N_5764);
nand U8863 (N_8863,N_5333,N_3868);
nor U8864 (N_8864,N_5197,N_3522);
nand U8865 (N_8865,N_5235,N_4793);
and U8866 (N_8866,N_4421,N_4666);
nand U8867 (N_8867,N_5954,N_3160);
nor U8868 (N_8868,N_4201,N_5070);
nand U8869 (N_8869,N_3070,N_4816);
nor U8870 (N_8870,N_4867,N_3085);
nand U8871 (N_8871,N_3393,N_5660);
nor U8872 (N_8872,N_5316,N_5121);
or U8873 (N_8873,N_3995,N_4896);
nand U8874 (N_8874,N_3674,N_3508);
nor U8875 (N_8875,N_3888,N_3225);
nand U8876 (N_8876,N_5557,N_4067);
and U8877 (N_8877,N_4947,N_4612);
nand U8878 (N_8878,N_4851,N_4858);
nor U8879 (N_8879,N_4905,N_4473);
nor U8880 (N_8880,N_4049,N_5399);
and U8881 (N_8881,N_4924,N_4128);
or U8882 (N_8882,N_3345,N_3773);
nor U8883 (N_8883,N_3872,N_3079);
nand U8884 (N_8884,N_3928,N_5329);
nor U8885 (N_8885,N_5731,N_4153);
nand U8886 (N_8886,N_3691,N_3034);
nor U8887 (N_8887,N_5003,N_4093);
and U8888 (N_8888,N_3144,N_3137);
and U8889 (N_8889,N_4163,N_3410);
and U8890 (N_8890,N_3409,N_5524);
nand U8891 (N_8891,N_3064,N_5461);
and U8892 (N_8892,N_3786,N_5888);
nand U8893 (N_8893,N_3054,N_4110);
nand U8894 (N_8894,N_5493,N_3930);
or U8895 (N_8895,N_5518,N_4189);
or U8896 (N_8896,N_3963,N_3660);
nor U8897 (N_8897,N_3002,N_4344);
nand U8898 (N_8898,N_4653,N_5488);
nand U8899 (N_8899,N_3874,N_5010);
nor U8900 (N_8900,N_5598,N_4508);
nand U8901 (N_8901,N_3564,N_3114);
or U8902 (N_8902,N_5290,N_5897);
nor U8903 (N_8903,N_5320,N_5882);
nand U8904 (N_8904,N_5763,N_5157);
and U8905 (N_8905,N_3921,N_4759);
and U8906 (N_8906,N_5122,N_5223);
or U8907 (N_8907,N_3147,N_3701);
and U8908 (N_8908,N_3425,N_3319);
and U8909 (N_8909,N_5195,N_4226);
and U8910 (N_8910,N_4324,N_3989);
nand U8911 (N_8911,N_5487,N_5959);
and U8912 (N_8912,N_3325,N_5236);
nor U8913 (N_8913,N_3436,N_4125);
nor U8914 (N_8914,N_5414,N_3223);
and U8915 (N_8915,N_4454,N_4151);
nand U8916 (N_8916,N_3571,N_3715);
and U8917 (N_8917,N_3383,N_3900);
nor U8918 (N_8918,N_5002,N_4274);
nand U8919 (N_8919,N_4042,N_5388);
nand U8920 (N_8920,N_5895,N_3055);
or U8921 (N_8921,N_5587,N_5816);
nand U8922 (N_8922,N_5747,N_3293);
nor U8923 (N_8923,N_5888,N_5020);
nand U8924 (N_8924,N_5257,N_4170);
nand U8925 (N_8925,N_3783,N_3743);
or U8926 (N_8926,N_4488,N_4627);
and U8927 (N_8927,N_4518,N_3353);
nand U8928 (N_8928,N_5574,N_5935);
and U8929 (N_8929,N_4496,N_4644);
or U8930 (N_8930,N_4472,N_4839);
and U8931 (N_8931,N_5658,N_5399);
nand U8932 (N_8932,N_5959,N_5582);
and U8933 (N_8933,N_5141,N_3061);
nand U8934 (N_8934,N_5972,N_4855);
and U8935 (N_8935,N_5872,N_3954);
nor U8936 (N_8936,N_5021,N_3187);
or U8937 (N_8937,N_5517,N_4036);
nand U8938 (N_8938,N_4432,N_4559);
nor U8939 (N_8939,N_5295,N_5695);
nor U8940 (N_8940,N_3570,N_5846);
or U8941 (N_8941,N_3126,N_3615);
nor U8942 (N_8942,N_5752,N_3884);
and U8943 (N_8943,N_3616,N_3628);
or U8944 (N_8944,N_3594,N_4657);
and U8945 (N_8945,N_4488,N_5762);
and U8946 (N_8946,N_3725,N_5280);
and U8947 (N_8947,N_4845,N_5792);
nor U8948 (N_8948,N_3657,N_5269);
nor U8949 (N_8949,N_4582,N_5368);
nor U8950 (N_8950,N_4989,N_3760);
nor U8951 (N_8951,N_5138,N_5987);
nand U8952 (N_8952,N_3670,N_5341);
and U8953 (N_8953,N_4339,N_4234);
or U8954 (N_8954,N_4114,N_5291);
nor U8955 (N_8955,N_5661,N_5034);
or U8956 (N_8956,N_5637,N_5165);
nor U8957 (N_8957,N_3773,N_4422);
nand U8958 (N_8958,N_3467,N_3677);
and U8959 (N_8959,N_5520,N_4676);
or U8960 (N_8960,N_4229,N_5527);
and U8961 (N_8961,N_5984,N_4942);
and U8962 (N_8962,N_5545,N_4215);
nor U8963 (N_8963,N_4036,N_4739);
and U8964 (N_8964,N_4773,N_4260);
or U8965 (N_8965,N_5537,N_5395);
and U8966 (N_8966,N_4648,N_3663);
nand U8967 (N_8967,N_5539,N_3712);
nand U8968 (N_8968,N_3331,N_4570);
nand U8969 (N_8969,N_5119,N_4788);
and U8970 (N_8970,N_4625,N_3764);
or U8971 (N_8971,N_3618,N_4378);
or U8972 (N_8972,N_3329,N_3210);
nand U8973 (N_8973,N_3034,N_3825);
or U8974 (N_8974,N_5565,N_3287);
nor U8975 (N_8975,N_4565,N_3104);
nand U8976 (N_8976,N_4450,N_3864);
and U8977 (N_8977,N_5541,N_4094);
and U8978 (N_8978,N_5530,N_3643);
and U8979 (N_8979,N_5533,N_5584);
and U8980 (N_8980,N_4753,N_4927);
nor U8981 (N_8981,N_5787,N_5056);
and U8982 (N_8982,N_3848,N_4367);
nor U8983 (N_8983,N_4032,N_4751);
nor U8984 (N_8984,N_3330,N_5206);
nand U8985 (N_8985,N_5618,N_5311);
nand U8986 (N_8986,N_5588,N_5420);
nand U8987 (N_8987,N_3080,N_4399);
nand U8988 (N_8988,N_4409,N_4243);
and U8989 (N_8989,N_5782,N_5762);
nand U8990 (N_8990,N_5094,N_4404);
nand U8991 (N_8991,N_3341,N_4131);
nand U8992 (N_8992,N_4674,N_5432);
nand U8993 (N_8993,N_4155,N_5868);
and U8994 (N_8994,N_3573,N_4206);
nand U8995 (N_8995,N_4436,N_5248);
or U8996 (N_8996,N_5829,N_4687);
nand U8997 (N_8997,N_5459,N_3038);
or U8998 (N_8998,N_4503,N_5067);
or U8999 (N_8999,N_4440,N_3651);
or U9000 (N_9000,N_7113,N_8297);
or U9001 (N_9001,N_6121,N_6308);
or U9002 (N_9002,N_8379,N_7766);
nor U9003 (N_9003,N_8210,N_6527);
nand U9004 (N_9004,N_7206,N_8591);
nor U9005 (N_9005,N_8540,N_6889);
or U9006 (N_9006,N_8994,N_8854);
nand U9007 (N_9007,N_6873,N_8174);
nand U9008 (N_9008,N_6325,N_8140);
or U9009 (N_9009,N_6459,N_8154);
nor U9010 (N_9010,N_8513,N_7239);
or U9011 (N_9011,N_8437,N_6736);
or U9012 (N_9012,N_6091,N_6200);
nor U9013 (N_9013,N_8902,N_8915);
nand U9014 (N_9014,N_8725,N_7467);
nand U9015 (N_9015,N_7472,N_6084);
nor U9016 (N_9016,N_6673,N_8380);
or U9017 (N_9017,N_7733,N_6102);
or U9018 (N_9018,N_6418,N_6001);
or U9019 (N_9019,N_6123,N_6570);
nor U9020 (N_9020,N_7145,N_7748);
or U9021 (N_9021,N_8441,N_6111);
and U9022 (N_9022,N_6843,N_7533);
nor U9023 (N_9023,N_6709,N_7009);
nor U9024 (N_9024,N_8081,N_6811);
or U9025 (N_9025,N_6161,N_7085);
or U9026 (N_9026,N_8518,N_7163);
and U9027 (N_9027,N_7875,N_8622);
nand U9028 (N_9028,N_7985,N_6810);
and U9029 (N_9029,N_8473,N_6993);
nand U9030 (N_9030,N_8044,N_8486);
or U9031 (N_9031,N_7799,N_8791);
nor U9032 (N_9032,N_8456,N_7922);
and U9033 (N_9033,N_6310,N_8980);
or U9034 (N_9034,N_6734,N_6557);
or U9035 (N_9035,N_7258,N_7696);
nand U9036 (N_9036,N_7908,N_8306);
nor U9037 (N_9037,N_7785,N_8179);
and U9038 (N_9038,N_8776,N_8218);
nand U9039 (N_9039,N_7606,N_6732);
or U9040 (N_9040,N_7599,N_6501);
nand U9041 (N_9041,N_8386,N_7381);
and U9042 (N_9042,N_6518,N_6417);
and U9043 (N_9043,N_6846,N_7192);
and U9044 (N_9044,N_7464,N_6405);
and U9045 (N_9045,N_8760,N_7168);
or U9046 (N_9046,N_8423,N_8021);
and U9047 (N_9047,N_7992,N_7105);
or U9048 (N_9048,N_7323,N_6723);
or U9049 (N_9049,N_6611,N_8624);
nor U9050 (N_9050,N_7614,N_6287);
nand U9051 (N_9051,N_7382,N_7889);
or U9052 (N_9052,N_6231,N_8975);
nor U9053 (N_9053,N_6593,N_8837);
nor U9054 (N_9054,N_6090,N_8178);
nand U9055 (N_9055,N_8199,N_7829);
nor U9056 (N_9056,N_7413,N_6982);
and U9057 (N_9057,N_6686,N_8057);
or U9058 (N_9058,N_6916,N_6027);
nand U9059 (N_9059,N_8598,N_8389);
or U9060 (N_9060,N_7132,N_6715);
and U9061 (N_9061,N_6936,N_6143);
and U9062 (N_9062,N_7135,N_7406);
nand U9063 (N_9063,N_7418,N_7705);
nor U9064 (N_9064,N_7964,N_7180);
or U9065 (N_9065,N_8069,N_7811);
and U9066 (N_9066,N_8692,N_7454);
or U9067 (N_9067,N_8283,N_8928);
and U9068 (N_9068,N_7111,N_8275);
nand U9069 (N_9069,N_6115,N_8601);
nand U9070 (N_9070,N_8876,N_7372);
nor U9071 (N_9071,N_8856,N_7230);
nor U9072 (N_9072,N_7063,N_8260);
or U9073 (N_9073,N_6549,N_7802);
and U9074 (N_9074,N_7336,N_6434);
nand U9075 (N_9075,N_6733,N_6623);
nor U9076 (N_9076,N_7858,N_7601);
nand U9077 (N_9077,N_7965,N_7888);
or U9078 (N_9078,N_7213,N_6770);
and U9079 (N_9079,N_7828,N_6573);
or U9080 (N_9080,N_7010,N_8807);
or U9081 (N_9081,N_6666,N_8961);
nor U9082 (N_9082,N_7668,N_7819);
nor U9083 (N_9083,N_6671,N_6995);
nand U9084 (N_9084,N_6924,N_8922);
and U9085 (N_9085,N_8214,N_8996);
or U9086 (N_9086,N_7879,N_8449);
and U9087 (N_9087,N_7319,N_8801);
nor U9088 (N_9088,N_6653,N_7591);
or U9089 (N_9089,N_7104,N_8477);
nor U9090 (N_9090,N_8372,N_7366);
nor U9091 (N_9091,N_8545,N_8819);
nor U9092 (N_9092,N_6324,N_6469);
and U9093 (N_9093,N_6941,N_6029);
nand U9094 (N_9094,N_7006,N_7184);
or U9095 (N_9095,N_7208,N_7298);
nand U9096 (N_9096,N_6712,N_6532);
and U9097 (N_9097,N_8217,N_8722);
nand U9098 (N_9098,N_8618,N_7855);
or U9099 (N_9099,N_7091,N_7868);
or U9100 (N_9100,N_7959,N_6250);
nor U9101 (N_9101,N_7337,N_6006);
nor U9102 (N_9102,N_6104,N_7334);
nand U9103 (N_9103,N_6689,N_7277);
nand U9104 (N_9104,N_7968,N_6510);
nand U9105 (N_9105,N_8172,N_7330);
and U9106 (N_9106,N_6122,N_7747);
nand U9107 (N_9107,N_8944,N_6453);
nor U9108 (N_9108,N_6462,N_6293);
or U9109 (N_9109,N_8409,N_8755);
nand U9110 (N_9110,N_6322,N_7867);
or U9111 (N_9111,N_8484,N_6050);
nand U9112 (N_9112,N_7436,N_7583);
nand U9113 (N_9113,N_8971,N_8194);
nor U9114 (N_9114,N_7942,N_8892);
nand U9115 (N_9115,N_6744,N_8553);
nand U9116 (N_9116,N_8352,N_8012);
nand U9117 (N_9117,N_7348,N_6270);
nand U9118 (N_9118,N_8036,N_8799);
or U9119 (N_9119,N_6368,N_6603);
nor U9120 (N_9120,N_6098,N_7592);
or U9121 (N_9121,N_6389,N_6222);
and U9122 (N_9122,N_7247,N_7934);
or U9123 (N_9123,N_6249,N_6407);
nor U9124 (N_9124,N_8170,N_7229);
and U9125 (N_9125,N_6705,N_6692);
nor U9126 (N_9126,N_8138,N_8815);
and U9127 (N_9127,N_6774,N_6632);
or U9128 (N_9128,N_6571,N_8030);
nor U9129 (N_9129,N_6391,N_7845);
or U9130 (N_9130,N_8060,N_7276);
nor U9131 (N_9131,N_7327,N_8497);
nand U9132 (N_9132,N_7417,N_8114);
or U9133 (N_9133,N_8511,N_6410);
nand U9134 (N_9134,N_8014,N_6708);
and U9135 (N_9135,N_7235,N_8623);
nor U9136 (N_9136,N_7448,N_7031);
nor U9137 (N_9137,N_7988,N_6254);
and U9138 (N_9138,N_8750,N_7181);
nand U9139 (N_9139,N_8318,N_8336);
nand U9140 (N_9140,N_7832,N_8781);
nor U9141 (N_9141,N_6536,N_6569);
nor U9142 (N_9142,N_7739,N_8538);
or U9143 (N_9143,N_6038,N_7000);
and U9144 (N_9144,N_8333,N_6721);
and U9145 (N_9145,N_7147,N_6826);
and U9146 (N_9146,N_6497,N_7118);
and U9147 (N_9147,N_7175,N_8914);
nand U9148 (N_9148,N_7201,N_7082);
and U9149 (N_9149,N_8888,N_6667);
nand U9150 (N_9150,N_7585,N_7919);
nor U9151 (N_9151,N_8300,N_7232);
nand U9152 (N_9152,N_6514,N_7289);
nand U9153 (N_9153,N_6042,N_7011);
nand U9154 (N_9154,N_6943,N_6897);
nor U9155 (N_9155,N_8316,N_6504);
nand U9156 (N_9156,N_6577,N_8146);
and U9157 (N_9157,N_6975,N_8433);
nand U9158 (N_9158,N_7822,N_6678);
or U9159 (N_9159,N_8880,N_7326);
and U9160 (N_9160,N_7291,N_8688);
or U9161 (N_9161,N_6302,N_7353);
nor U9162 (N_9162,N_7073,N_8071);
or U9163 (N_9163,N_7565,N_6074);
or U9164 (N_9164,N_8416,N_6500);
and U9165 (N_9165,N_8884,N_7633);
or U9166 (N_9166,N_6711,N_7935);
nor U9167 (N_9167,N_7646,N_8224);
and U9168 (N_9168,N_7831,N_7282);
or U9169 (N_9169,N_8662,N_8483);
nand U9170 (N_9170,N_6015,N_6145);
xnor U9171 (N_9171,N_8070,N_7301);
or U9172 (N_9172,N_7989,N_8939);
or U9173 (N_9173,N_7788,N_8699);
nor U9174 (N_9174,N_6512,N_6760);
xor U9175 (N_9175,N_7746,N_6220);
nor U9176 (N_9176,N_7316,N_8759);
and U9177 (N_9177,N_7424,N_6072);
and U9178 (N_9178,N_6358,N_8574);
nand U9179 (N_9179,N_7146,N_7459);
nand U9180 (N_9180,N_6830,N_8522);
and U9181 (N_9181,N_8577,N_6726);
and U9182 (N_9182,N_6820,N_7776);
nand U9183 (N_9183,N_6552,N_7440);
nand U9184 (N_9184,N_6968,N_8705);
nor U9185 (N_9185,N_7516,N_6725);
nand U9186 (N_9186,N_8698,N_6329);
or U9187 (N_9187,N_6352,N_8887);
nand U9188 (N_9188,N_7661,N_8842);
and U9189 (N_9189,N_7854,N_6173);
nor U9190 (N_9190,N_7245,N_8749);
and U9191 (N_9191,N_7153,N_8774);
nor U9192 (N_9192,N_6952,N_6039);
nand U9193 (N_9193,N_6581,N_7209);
nand U9194 (N_9194,N_6963,N_7364);
and U9195 (N_9195,N_6153,N_6258);
nand U9196 (N_9196,N_8637,N_7607);
nand U9197 (N_9197,N_8830,N_8615);
nor U9198 (N_9198,N_8335,N_6940);
and U9199 (N_9199,N_7223,N_8547);
and U9200 (N_9200,N_7665,N_8008);
or U9201 (N_9201,N_8960,N_8027);
nor U9202 (N_9202,N_8461,N_6208);
or U9203 (N_9203,N_7090,N_6735);
nand U9204 (N_9204,N_7021,N_6010);
nand U9205 (N_9205,N_8289,N_8765);
nor U9206 (N_9206,N_6845,N_7707);
nor U9207 (N_9207,N_8909,N_8422);
or U9208 (N_9208,N_6194,N_8225);
and U9209 (N_9209,N_6592,N_6065);
nor U9210 (N_9210,N_8671,N_8576);
nor U9211 (N_9211,N_7621,N_8459);
nand U9212 (N_9212,N_8093,N_7126);
nand U9213 (N_9213,N_8200,N_7331);
and U9214 (N_9214,N_7830,N_7904);
nand U9215 (N_9215,N_7625,N_8309);
or U9216 (N_9216,N_6199,N_6252);
or U9217 (N_9217,N_8764,N_8653);
or U9218 (N_9218,N_8703,N_6842);
nor U9219 (N_9219,N_7341,N_7624);
nand U9220 (N_9220,N_8083,N_8525);
and U9221 (N_9221,N_6400,N_7219);
nand U9222 (N_9222,N_8353,N_7664);
nand U9223 (N_9223,N_8492,N_8462);
or U9224 (N_9224,N_8312,N_6408);
nor U9225 (N_9225,N_7254,N_7900);
or U9226 (N_9226,N_8654,N_7752);
nand U9227 (N_9227,N_7347,N_7461);
nor U9228 (N_9228,N_8936,N_6881);
or U9229 (N_9229,N_6402,N_8908);
nor U9230 (N_9230,N_7984,N_6095);
or U9231 (N_9231,N_7619,N_8921);
nor U9232 (N_9232,N_7283,N_8519);
nand U9233 (N_9233,N_8120,N_6089);
or U9234 (N_9234,N_6991,N_7704);
and U9235 (N_9235,N_8421,N_6808);
nand U9236 (N_9236,N_7953,N_6851);
and U9237 (N_9237,N_6463,N_7342);
nand U9238 (N_9238,N_8916,N_8932);
nor U9239 (N_9239,N_8682,N_8208);
nor U9240 (N_9240,N_6766,N_8090);
or U9241 (N_9241,N_7026,N_8464);
and U9242 (N_9242,N_8374,N_7398);
nor U9243 (N_9243,N_6019,N_6583);
or U9244 (N_9244,N_6366,N_8162);
nor U9245 (N_9245,N_6687,N_7151);
nor U9246 (N_9246,N_7380,N_6786);
and U9247 (N_9247,N_6318,N_7610);
nor U9248 (N_9248,N_6765,N_8629);
nand U9249 (N_9249,N_7658,N_7916);
nor U9250 (N_9250,N_8667,N_7495);
or U9251 (N_9251,N_7269,N_8118);
nand U9252 (N_9252,N_7048,N_8206);
nand U9253 (N_9253,N_8106,N_8500);
and U9254 (N_9254,N_6460,N_7582);
nand U9255 (N_9255,N_6520,N_6567);
or U9256 (N_9256,N_7651,N_7886);
nor U9257 (N_9257,N_6507,N_7991);
nand U9258 (N_9258,N_7553,N_8579);
and U9259 (N_9259,N_8498,N_7540);
nor U9260 (N_9260,N_8376,N_6396);
nand U9261 (N_9261,N_7713,N_7098);
nor U9262 (N_9262,N_6763,N_6620);
nor U9263 (N_9263,N_6761,N_7487);
or U9264 (N_9264,N_8526,N_7532);
and U9265 (N_9265,N_6175,N_7825);
or U9266 (N_9266,N_7772,N_7051);
and U9267 (N_9267,N_6850,N_7689);
or U9268 (N_9268,N_8331,N_8544);
nand U9269 (N_9269,N_6238,N_8038);
or U9270 (N_9270,N_7499,N_6893);
nor U9271 (N_9271,N_8867,N_7352);
nand U9272 (N_9272,N_7268,N_8633);
or U9273 (N_9273,N_7370,N_8963);
or U9274 (N_9274,N_6132,N_6605);
nand U9275 (N_9275,N_8866,N_6861);
nor U9276 (N_9276,N_8864,N_7195);
nor U9277 (N_9277,N_7311,N_6730);
or U9278 (N_9278,N_8229,N_8677);
and U9279 (N_9279,N_6355,N_6246);
nand U9280 (N_9280,N_6664,N_6411);
nor U9281 (N_9281,N_6644,N_6607);
or U9282 (N_9282,N_8125,N_7906);
nor U9283 (N_9283,N_8542,N_7156);
and U9284 (N_9284,N_7310,N_6007);
nor U9285 (N_9285,N_7727,N_8643);
nor U9286 (N_9286,N_8778,N_7620);
nor U9287 (N_9287,N_7617,N_7067);
nor U9288 (N_9288,N_8142,N_6745);
nor U9289 (N_9289,N_7270,N_6415);
or U9290 (N_9290,N_8246,N_8109);
and U9291 (N_9291,N_7231,N_7481);
or U9292 (N_9292,N_8753,N_6904);
or U9293 (N_9293,N_8391,N_8238);
xor U9294 (N_9294,N_7027,N_6277);
or U9295 (N_9295,N_6638,N_7237);
and U9296 (N_9296,N_8895,N_7806);
nor U9297 (N_9297,N_7884,N_8950);
or U9298 (N_9298,N_6420,N_8382);
and U9299 (N_9299,N_8905,N_6909);
nand U9300 (N_9300,N_8097,N_7715);
nor U9301 (N_9301,N_6630,N_6868);
or U9302 (N_9302,N_6379,N_8323);
nand U9303 (N_9303,N_6409,N_6443);
nand U9304 (N_9304,N_6013,N_6890);
and U9305 (N_9305,N_8746,N_7567);
or U9306 (N_9306,N_6719,N_6061);
nor U9307 (N_9307,N_6346,N_8192);
nand U9308 (N_9308,N_6315,N_8346);
and U9309 (N_9309,N_8065,N_8619);
or U9310 (N_9310,N_8990,N_7912);
and U9311 (N_9311,N_7020,N_6369);
and U9312 (N_9312,N_8752,N_6838);
nand U9313 (N_9313,N_8509,N_8689);
or U9314 (N_9314,N_8797,N_6584);
and U9315 (N_9315,N_7386,N_6296);
nor U9316 (N_9316,N_6706,N_7182);
or U9317 (N_9317,N_6588,N_6377);
or U9318 (N_9318,N_7155,N_6471);
nand U9319 (N_9319,N_7936,N_7489);
and U9320 (N_9320,N_8475,N_6847);
nor U9321 (N_9321,N_7221,N_6187);
nor U9322 (N_9322,N_6781,N_7123);
nand U9323 (N_9323,N_6729,N_8239);
nand U9324 (N_9324,N_6449,N_8517);
and U9325 (N_9325,N_7076,N_6882);
nand U9326 (N_9326,N_7226,N_7969);
and U9327 (N_9327,N_8453,N_8670);
or U9328 (N_9328,N_7509,N_8103);
or U9329 (N_9329,N_8638,N_8358);
nor U9330 (N_9330,N_6236,N_8898);
nor U9331 (N_9331,N_6937,N_7400);
nor U9332 (N_9332,N_7143,N_7497);
or U9333 (N_9333,N_6951,N_8155);
and U9334 (N_9334,N_6643,N_8332);
or U9335 (N_9335,N_6886,N_6590);
or U9336 (N_9336,N_8078,N_6752);
nor U9337 (N_9337,N_8468,N_6836);
nand U9338 (N_9338,N_6134,N_8712);
nor U9339 (N_9339,N_8651,N_7631);
nor U9340 (N_9340,N_7477,N_8933);
or U9341 (N_9341,N_6235,N_6784);
or U9342 (N_9342,N_7305,N_8706);
or U9343 (N_9343,N_7526,N_8878);
nor U9344 (N_9344,N_6544,N_6896);
and U9345 (N_9345,N_6515,N_6964);
nand U9346 (N_9346,N_7358,N_6870);
nand U9347 (N_9347,N_6044,N_6362);
nand U9348 (N_9348,N_7641,N_6468);
or U9349 (N_9349,N_8285,N_7340);
nand U9350 (N_9350,N_8969,N_8405);
and U9351 (N_9351,N_6360,N_7602);
and U9352 (N_9352,N_6164,N_7684);
nand U9353 (N_9353,N_8885,N_7172);
or U9354 (N_9354,N_6912,N_8116);
and U9355 (N_9355,N_6867,N_8567);
nand U9356 (N_9356,N_6969,N_8427);
nand U9357 (N_9357,N_8344,N_8582);
nor U9358 (N_9358,N_7202,N_8485);
and U9359 (N_9359,N_6455,N_8701);
or U9360 (N_9360,N_8953,N_8274);
or U9361 (N_9361,N_6342,N_8167);
and U9362 (N_9362,N_6910,N_8041);
nor U9363 (N_9363,N_8853,N_7753);
nand U9364 (N_9364,N_8700,N_6048);
or U9365 (N_9365,N_7470,N_6679);
nand U9366 (N_9366,N_8621,N_8228);
and U9367 (N_9367,N_6777,N_8448);
nand U9368 (N_9368,N_7843,N_6124);
and U9369 (N_9369,N_8899,N_8434);
nand U9370 (N_9370,N_6269,N_6414);
nand U9371 (N_9371,N_8834,N_8438);
or U9372 (N_9372,N_6382,N_7608);
and U9373 (N_9373,N_8089,N_8010);
or U9374 (N_9374,N_7675,N_7257);
and U9375 (N_9375,N_8173,N_6917);
and U9376 (N_9376,N_8478,N_6509);
nand U9377 (N_9377,N_6107,N_6722);
and U9378 (N_9378,N_8197,N_8148);
or U9379 (N_9379,N_6742,N_8847);
or U9380 (N_9380,N_6802,N_8641);
nand U9381 (N_9381,N_7244,N_7913);
nand U9382 (N_9382,N_6884,N_6997);
and U9383 (N_9383,N_7449,N_6985);
and U9384 (N_9384,N_8958,N_8292);
nor U9385 (N_9385,N_6797,N_6171);
or U9386 (N_9386,N_8366,N_8691);
nand U9387 (N_9387,N_6697,N_8613);
or U9388 (N_9388,N_6189,N_7910);
nor U9389 (N_9389,N_6427,N_6621);
nor U9390 (N_9390,N_6096,N_7273);
nor U9391 (N_9391,N_8100,N_8020);
and U9392 (N_9392,N_6141,N_7948);
nor U9393 (N_9393,N_6147,N_8890);
or U9394 (N_9394,N_7199,N_8852);
and U9395 (N_9395,N_6755,N_8543);
nor U9396 (N_9396,N_8054,N_8989);
nor U9397 (N_9397,N_6388,N_7078);
nand U9398 (N_9398,N_8003,N_7018);
and U9399 (N_9399,N_7022,N_8767);
and U9400 (N_9400,N_7649,N_7432);
or U9401 (N_9401,N_7214,N_8270);
and U9402 (N_9402,N_8603,N_7850);
or U9403 (N_9403,N_6618,N_6680);
and U9404 (N_9404,N_6412,N_7049);
nand U9405 (N_9405,N_8411,N_8645);
nand U9406 (N_9406,N_7630,N_7429);
nand U9407 (N_9407,N_8957,N_8988);
and U9408 (N_9408,N_6986,N_6767);
nand U9409 (N_9409,N_7503,N_7399);
xor U9410 (N_9410,N_8308,N_7343);
nor U9411 (N_9411,N_8773,N_8810);
nor U9412 (N_9412,N_7929,N_6298);
or U9413 (N_9413,N_7137,N_7815);
and U9414 (N_9414,N_6057,N_6565);
and U9415 (N_9415,N_8049,N_6780);
nor U9416 (N_9416,N_6608,N_7584);
and U9417 (N_9417,N_7566,N_8304);
or U9418 (N_9418,N_8945,N_6987);
or U9419 (N_9419,N_8600,N_6645);
nor U9420 (N_9420,N_7166,N_7158);
nor U9421 (N_9421,N_8666,N_8663);
or U9422 (N_9422,N_6320,N_8278);
or U9423 (N_9423,N_6465,N_6676);
nand U9424 (N_9424,N_7212,N_6421);
and U9425 (N_9425,N_8973,N_8396);
nand U9426 (N_9426,N_7821,N_6399);
or U9427 (N_9427,N_8658,N_8233);
and U9428 (N_9428,N_7874,N_7657);
nand U9429 (N_9429,N_7263,N_7387);
or U9430 (N_9430,N_8570,N_8145);
or U9431 (N_9431,N_7652,N_7309);
and U9432 (N_9432,N_7426,N_6373);
or U9433 (N_9433,N_7852,N_7248);
nor U9434 (N_9434,N_7218,N_7545);
or U9435 (N_9435,N_7933,N_6540);
and U9436 (N_9436,N_8606,N_8368);
and U9437 (N_9437,N_6387,N_8037);
and U9438 (N_9438,N_8609,N_7148);
nor U9439 (N_9439,N_7278,N_6306);
nand U9440 (N_9440,N_7924,N_8839);
and U9441 (N_9441,N_6158,N_7307);
nor U9442 (N_9442,N_7150,N_7292);
nor U9443 (N_9443,N_7109,N_6472);
and U9444 (N_9444,N_8501,N_7890);
and U9445 (N_9445,N_7297,N_7012);
and U9446 (N_9446,N_6345,N_6785);
nor U9447 (N_9447,N_7447,N_7719);
or U9448 (N_9448,N_8320,N_8965);
or U9449 (N_9449,N_7701,N_6751);
nor U9450 (N_9450,N_8171,N_7046);
or U9451 (N_9451,N_6183,N_8436);
nor U9452 (N_9452,N_6718,N_6641);
or U9453 (N_9453,N_6610,N_8182);
or U9454 (N_9454,N_6159,N_7303);
nor U9455 (N_9455,N_7070,N_6028);
and U9456 (N_9456,N_6833,N_7967);
or U9457 (N_9457,N_7589,N_7878);
nand U9458 (N_9458,N_8067,N_8018);
or U9459 (N_9459,N_6753,N_6077);
nor U9460 (N_9460,N_7355,N_8105);
nand U9461 (N_9461,N_7198,N_6340);
nor U9462 (N_9462,N_8001,N_7590);
and U9463 (N_9463,N_6218,N_7412);
nand U9464 (N_9464,N_7655,N_8860);
and U9465 (N_9465,N_7228,N_8465);
nor U9466 (N_9466,N_7826,N_6155);
nand U9467 (N_9467,N_8910,N_6349);
nor U9468 (N_9468,N_7650,N_7981);
and U9469 (N_9469,N_8446,N_8400);
or U9470 (N_9470,N_7521,N_7669);
or U9471 (N_9471,N_7600,N_6927);
and U9472 (N_9472,N_7869,N_7127);
or U9473 (N_9473,N_8552,N_6140);
or U9474 (N_9474,N_8151,N_6871);
nand U9475 (N_9475,N_8452,N_6008);
nor U9476 (N_9476,N_6972,N_7133);
nor U9477 (N_9477,N_7511,N_6865);
nand U9478 (N_9478,N_7494,N_8707);
or U9479 (N_9479,N_7036,N_8045);
or U9480 (N_9480,N_8982,N_6572);
nand U9481 (N_9481,N_7549,N_7409);
nand U9482 (N_9482,N_7420,N_7042);
or U9483 (N_9483,N_7528,N_8467);
nor U9484 (N_9484,N_6051,N_6551);
nand U9485 (N_9485,N_6775,N_7667);
and U9486 (N_9486,N_7573,N_8076);
and U9487 (N_9487,N_8403,N_7741);
nor U9488 (N_9488,N_8310,N_7217);
nand U9489 (N_9489,N_6973,N_8798);
nand U9490 (N_9490,N_8868,N_7434);
or U9491 (N_9491,N_7207,N_7708);
or U9492 (N_9492,N_6849,N_7859);
xor U9493 (N_9493,N_6481,N_7853);
or U9494 (N_9494,N_7473,N_8087);
and U9495 (N_9495,N_6834,N_7140);
and U9496 (N_9496,N_6146,N_7029);
or U9497 (N_9497,N_7937,N_6696);
or U9498 (N_9498,N_7083,N_6280);
nor U9499 (N_9499,N_8882,N_6052);
or U9500 (N_9500,N_8803,N_6185);
nor U9501 (N_9501,N_7654,N_8630);
nand U9502 (N_9502,N_6063,N_6848);
nand U9503 (N_9503,N_7392,N_8241);
nand U9504 (N_9504,N_8978,N_6548);
or U9505 (N_9505,N_7881,N_6292);
nand U9506 (N_9506,N_7982,N_8286);
nor U9507 (N_9507,N_6274,N_8693);
nor U9508 (N_9508,N_8408,N_6169);
or U9509 (N_9509,N_7157,N_8548);
or U9510 (N_9510,N_6542,N_6702);
nand U9511 (N_9511,N_7446,N_6984);
nand U9512 (N_9512,N_6492,N_7222);
nor U9513 (N_9513,N_8930,N_6788);
and U9514 (N_9514,N_6365,N_8959);
nand U9515 (N_9515,N_8339,N_8367);
nor U9516 (N_9516,N_8967,N_7609);
nand U9517 (N_9517,N_6604,N_8748);
nor U9518 (N_9518,N_7290,N_7275);
or U9519 (N_9519,N_7108,N_6499);
nand U9520 (N_9520,N_7542,N_7883);
nor U9521 (N_9521,N_7349,N_6299);
nand U9522 (N_9522,N_7040,N_7866);
and U9523 (N_9523,N_7317,N_6474);
and U9524 (N_9524,N_8313,N_7714);
and U9525 (N_9525,N_6447,N_8407);
and U9526 (N_9526,N_6866,N_6945);
and U9527 (N_9527,N_6263,N_7486);
or U9528 (N_9528,N_7357,N_6976);
nand U9529 (N_9529,N_7069,N_6339);
nand U9530 (N_9530,N_7525,N_7068);
and U9531 (N_9531,N_8463,N_7014);
or U9532 (N_9532,N_7836,N_8432);
or U9533 (N_9533,N_7087,N_6477);
nand U9534 (N_9534,N_7575,N_7496);
nor U9535 (N_9535,N_8596,N_6559);
and U9536 (N_9536,N_7980,N_8190);
nor U9537 (N_9537,N_6311,N_6338);
and U9538 (N_9538,N_8032,N_8495);
nand U9539 (N_9539,N_6841,N_8028);
and U9540 (N_9540,N_7954,N_8679);
or U9541 (N_9541,N_8795,N_8169);
nand U9542 (N_9542,N_7117,N_7138);
nand U9543 (N_9543,N_7504,N_8551);
or U9544 (N_9544,N_7880,N_8835);
and U9545 (N_9545,N_8137,N_8938);
or U9546 (N_9546,N_8072,N_7756);
or U9547 (N_9547,N_8326,N_8595);
nand U9548 (N_9548,N_8625,N_7286);
and U9549 (N_9549,N_8636,N_6117);
nor U9550 (N_9550,N_6922,N_6869);
and U9551 (N_9551,N_8563,N_8825);
nor U9552 (N_9552,N_6546,N_8786);
nor U9553 (N_9553,N_7827,N_6022);
nand U9554 (N_9554,N_7813,N_6907);
nand U9555 (N_9555,N_6395,N_7488);
or U9556 (N_9556,N_7564,N_7227);
or U9557 (N_9557,N_6478,N_8796);
nor U9558 (N_9558,N_7103,N_6020);
nor U9559 (N_9559,N_7579,N_8766);
nand U9560 (N_9560,N_7623,N_8634);
or U9561 (N_9561,N_8572,N_6994);
or U9562 (N_9562,N_8974,N_8530);
nor U9563 (N_9563,N_8804,N_8288);
or U9564 (N_9564,N_6083,N_6799);
nand U9565 (N_9565,N_8077,N_8979);
and U9566 (N_9566,N_7512,N_8829);
or U9567 (N_9567,N_8115,N_6919);
nand U9568 (N_9568,N_6212,N_7837);
or U9569 (N_9569,N_6162,N_8136);
and U9570 (N_9570,N_6386,N_8482);
and U9571 (N_9571,N_6361,N_8535);
nor U9572 (N_9572,N_6467,N_8558);
or U9573 (N_9573,N_6764,N_8529);
nand U9574 (N_9574,N_8581,N_6404);
nor U9575 (N_9575,N_8052,N_8510);
or U9576 (N_9576,N_7302,N_7110);
nand U9577 (N_9577,N_7864,N_7946);
and U9578 (N_9578,N_7013,N_8481);
and U9579 (N_9579,N_7405,N_6815);
nand U9580 (N_9580,N_6275,N_7491);
nor U9581 (N_9581,N_7568,N_7056);
and U9582 (N_9582,N_6609,N_8232);
nor U9583 (N_9583,N_6589,N_6628);
or U9584 (N_9584,N_7122,N_8187);
nand U9585 (N_9585,N_7299,N_7401);
or U9586 (N_9586,N_7717,N_6495);
and U9587 (N_9587,N_6486,N_8296);
or U9588 (N_9588,N_7120,N_7834);
and U9589 (N_9589,N_8127,N_6773);
nor U9590 (N_9590,N_8234,N_6343);
and U9591 (N_9591,N_8413,N_8307);
nand U9592 (N_9592,N_7718,N_7431);
and U9593 (N_9593,N_8317,N_6880);
and U9594 (N_9594,N_8254,N_8681);
and U9595 (N_9595,N_8647,N_8425);
nor U9596 (N_9596,N_7692,N_6018);
or U9597 (N_9597,N_7478,N_7178);
or U9598 (N_9598,N_8337,N_8757);
nor U9599 (N_9599,N_7952,N_6452);
xnor U9600 (N_9600,N_8479,N_8727);
nor U9601 (N_9601,N_7377,N_6385);
nor U9602 (N_9602,N_6363,N_6071);
nor U9603 (N_9603,N_7736,N_6961);
nand U9604 (N_9604,N_8664,N_6717);
nand U9605 (N_9605,N_7320,N_7075);
nand U9606 (N_9606,N_8585,N_8782);
nor U9607 (N_9607,N_8435,N_7999);
or U9608 (N_9608,N_8818,N_7427);
nor U9609 (N_9609,N_6531,N_7750);
or U9610 (N_9610,N_7131,N_6506);
nor U9611 (N_9611,N_7743,N_7994);
nand U9612 (N_9612,N_6999,N_6313);
and U9613 (N_9613,N_7844,N_6290);
and U9614 (N_9614,N_6652,N_8019);
nand U9615 (N_9615,N_8954,N_8098);
nand U9616 (N_9616,N_6891,N_6446);
or U9617 (N_9617,N_7892,N_7215);
nor U9618 (N_9618,N_6075,N_7998);
nand U9619 (N_9619,N_8524,N_8783);
nor U9620 (N_9620,N_6436,N_6023);
and U9621 (N_9621,N_7637,N_7116);
nand U9622 (N_9622,N_6930,N_6367);
and U9623 (N_9623,N_7315,N_7928);
and U9624 (N_9624,N_8756,N_7345);
nor U9625 (N_9625,N_6088,N_8772);
or U9626 (N_9626,N_7089,N_6996);
and U9627 (N_9627,N_6305,N_6574);
nand U9628 (N_9628,N_6055,N_7445);
and U9629 (N_9629,N_8997,N_6243);
and U9630 (N_9630,N_6168,N_7045);
xnor U9631 (N_9631,N_7693,N_7955);
nand U9632 (N_9632,N_7930,N_7164);
nand U9633 (N_9633,N_6179,N_8875);
nor U9634 (N_9634,N_7957,N_7442);
and U9635 (N_9635,N_8935,N_8424);
and U9636 (N_9636,N_6012,N_6668);
nor U9637 (N_9637,N_7430,N_6646);
or U9638 (N_9638,N_8929,N_7862);
nand U9639 (N_9639,N_7923,N_7676);
nand U9640 (N_9640,N_6440,N_7578);
nor U9641 (N_9641,N_6648,N_8754);
nand U9642 (N_9642,N_8159,N_6204);
nand U9643 (N_9643,N_6461,N_8620);
nor U9644 (N_9644,N_7622,N_6598);
and U9645 (N_9645,N_6066,N_6174);
nor U9646 (N_9646,N_7513,N_8769);
nand U9647 (N_9647,N_8454,N_8363);
nand U9648 (N_9648,N_7546,N_7035);
and U9649 (N_9649,N_7917,N_6911);
and U9650 (N_9650,N_7997,N_8135);
or U9651 (N_9651,N_8840,N_8350);
nand U9652 (N_9652,N_6151,N_6196);
nor U9653 (N_9653,N_6526,N_7800);
and U9654 (N_9654,N_7775,N_6047);
and U9655 (N_9655,N_7462,N_7416);
nor U9656 (N_9656,N_7267,N_7190);
nor U9657 (N_9657,N_6827,N_7136);
or U9658 (N_9658,N_8271,N_8040);
and U9659 (N_9659,N_7898,N_7793);
nand U9660 (N_9660,N_7945,N_6939);
nor U9661 (N_9661,N_7313,N_6017);
nor U9662 (N_9662,N_8720,N_7950);
nor U9663 (N_9663,N_7096,N_6073);
nand U9664 (N_9664,N_6378,N_7807);
nor U9665 (N_9665,N_7414,N_7004);
nor U9666 (N_9666,N_7433,N_7662);
nor U9667 (N_9667,N_6156,N_6284);
nor U9668 (N_9668,N_8442,N_8573);
or U9669 (N_9669,N_7863,N_8132);
or U9670 (N_9670,N_7673,N_7160);
or U9671 (N_9671,N_6203,N_7037);
or U9672 (N_9672,N_6519,N_6631);
nand U9673 (N_9673,N_6247,N_6351);
and U9674 (N_9674,N_6606,N_8102);
nand U9675 (N_9675,N_7970,N_8005);
and U9676 (N_9676,N_6674,N_8053);
nor U9677 (N_9677,N_7961,N_6923);
and U9678 (N_9678,N_8447,N_6424);
and U9679 (N_9679,N_7086,N_7947);
nand U9680 (N_9680,N_6129,N_6135);
and U9681 (N_9681,N_8977,N_8360);
and U9682 (N_9682,N_8602,N_8470);
and U9683 (N_9683,N_7457,N_7949);
or U9684 (N_9684,N_8583,N_6069);
nand U9685 (N_9685,N_6683,N_6494);
and U9686 (N_9686,N_8133,N_6166);
or U9687 (N_9687,N_8833,N_8657);
or U9688 (N_9688,N_7066,N_8695);
nor U9689 (N_9689,N_8047,N_8665);
and U9690 (N_9690,N_6224,N_8257);
nor U9691 (N_9691,N_6707,N_8362);
or U9692 (N_9692,N_8160,N_7072);
or U9693 (N_9693,N_6457,N_8923);
nand U9694 (N_9694,N_8420,N_8016);
or U9695 (N_9695,N_8341,N_7724);
or U9696 (N_9696,N_8401,N_6078);
nand U9697 (N_9697,N_7877,N_6601);
nand U9698 (N_9698,N_6348,N_7993);
or U9699 (N_9699,N_8043,N_7407);
nor U9700 (N_9700,N_8302,N_7196);
nand U9701 (N_9701,N_6778,N_7365);
nor U9702 (N_9702,N_7849,N_8157);
nand U9703 (N_9703,N_6928,N_8702);
and U9704 (N_9704,N_7304,N_7015);
and U9705 (N_9705,N_8911,N_8377);
nor U9706 (N_9706,N_6304,N_8236);
nor U9707 (N_9707,N_6860,N_7119);
nand U9708 (N_9708,N_6690,N_7795);
nor U9709 (N_9709,N_7474,N_8277);
nor U9710 (N_9710,N_6675,N_6148);
and U9711 (N_9711,N_6108,N_8414);
and U9712 (N_9712,N_6594,N_7902);
and U9713 (N_9713,N_8281,N_7716);
nor U9714 (N_9714,N_8319,N_8451);
nand U9715 (N_9715,N_7710,N_7911);
nand U9716 (N_9716,N_8279,N_8298);
nor U9717 (N_9717,N_6965,N_7121);
xor U9718 (N_9718,N_7041,N_7514);
or U9719 (N_9719,N_7644,N_6257);
nand U9720 (N_9720,N_6303,N_6438);
and U9721 (N_9721,N_7539,N_6724);
nor U9722 (N_9722,N_8792,N_8042);
or U9723 (N_9723,N_7783,N_8177);
or U9724 (N_9724,N_6403,N_6265);
or U9725 (N_9725,N_6230,N_7475);
or U9726 (N_9726,N_7538,N_7958);
and U9727 (N_9727,N_8355,N_8684);
nand U9728 (N_9728,N_8846,N_6233);
and U9729 (N_9729,N_7114,N_6980);
nor U9730 (N_9730,N_8533,N_6289);
nor U9731 (N_9731,N_7019,N_7321);
and U9732 (N_9732,N_6079,N_8985);
nand U9733 (N_9733,N_6428,N_7165);
or U9734 (N_9734,N_6353,N_7216);
nand U9735 (N_9735,N_7897,N_7373);
and U9736 (N_9736,N_6337,N_8265);
or U9737 (N_9737,N_8881,N_8342);
and U9738 (N_9738,N_6336,N_6261);
or U9739 (N_9739,N_6334,N_8439);
or U9740 (N_9740,N_6872,N_6864);
nor U9741 (N_9741,N_7596,N_7860);
and U9742 (N_9742,N_7876,N_6710);
or U9743 (N_9743,N_6375,N_8430);
or U9744 (N_9744,N_6914,N_7141);
or U9745 (N_9745,N_8877,N_8836);
nand U9746 (N_9746,N_6037,N_7439);
nand U9747 (N_9747,N_7523,N_7547);
nand U9748 (N_9748,N_7926,N_6649);
and U9749 (N_9749,N_8649,N_8294);
nor U9750 (N_9750,N_7515,N_7253);
xnor U9751 (N_9751,N_6942,N_6295);
and U9752 (N_9752,N_7951,N_8023);
nor U9753 (N_9753,N_7328,N_8196);
or U9754 (N_9754,N_7351,N_6371);
nor U9755 (N_9755,N_6268,N_8527);
and U9756 (N_9756,N_7761,N_6054);
nand U9757 (N_9757,N_6561,N_6234);
nor U9758 (N_9758,N_8266,N_6271);
nor U9759 (N_9759,N_8085,N_8942);
nor U9760 (N_9760,N_7570,N_8491);
nor U9761 (N_9761,N_7960,N_6701);
and U9762 (N_9762,N_6556,N_8984);
nand U9763 (N_9763,N_6030,N_7893);
nand U9764 (N_9764,N_8571,N_6524);
nor U9765 (N_9765,N_7394,N_6464);
nor U9766 (N_9766,N_8295,N_6125);
nor U9767 (N_9767,N_6330,N_8869);
nor U9768 (N_9768,N_8176,N_7259);
nor U9769 (N_9769,N_7017,N_8369);
nor U9770 (N_9770,N_8301,N_6491);
or U9771 (N_9771,N_6684,N_7847);
nor U9772 (N_9772,N_8340,N_7306);
and U9773 (N_9773,N_7179,N_7099);
and U9774 (N_9774,N_7817,N_7780);
and U9775 (N_9775,N_7790,N_7551);
or U9776 (N_9776,N_7786,N_7312);
nand U9777 (N_9777,N_8843,N_6413);
nand U9778 (N_9778,N_7694,N_6482);
or U9779 (N_9779,N_8195,N_8450);
nand U9780 (N_9780,N_8956,N_8696);
nand U9781 (N_9781,N_8805,N_7233);
nor U9782 (N_9782,N_7576,N_7808);
or U9783 (N_9783,N_7774,N_7846);
nand U9784 (N_9784,N_7636,N_7534);
nand U9785 (N_9785,N_8784,N_6956);
nand U9786 (N_9786,N_8082,N_6458);
and U9787 (N_9787,N_8476,N_6824);
nand U9788 (N_9788,N_7396,N_6267);
and U9789 (N_9789,N_7789,N_7125);
nand U9790 (N_9790,N_8489,N_7674);
and U9791 (N_9791,N_7851,N_6131);
or U9792 (N_9792,N_8787,N_7870);
nor U9793 (N_9793,N_8612,N_7084);
and U9794 (N_9794,N_6728,N_8250);
nor U9795 (N_9795,N_7144,N_8894);
or U9796 (N_9796,N_8589,N_7560);
nand U9797 (N_9797,N_8024,N_7452);
nand U9798 (N_9798,N_8378,N_7618);
nand U9799 (N_9799,N_7225,N_8775);
and U9800 (N_9800,N_6035,N_7971);
nor U9801 (N_9801,N_8900,N_6319);
and U9802 (N_9802,N_8412,N_7450);
nand U9803 (N_9803,N_8007,N_8680);
or U9804 (N_9804,N_6207,N_8119);
or U9805 (N_9805,N_6307,N_6016);
or U9806 (N_9806,N_7279,N_6757);
and U9807 (N_9807,N_6118,N_7055);
or U9808 (N_9808,N_7905,N_6627);
nor U9809 (N_9809,N_7865,N_7562);
or U9810 (N_9810,N_7663,N_8096);
or U9811 (N_9811,N_6803,N_7966);
and U9812 (N_9812,N_6456,N_6754);
nor U9813 (N_9813,N_8927,N_8889);
or U9814 (N_9814,N_8381,N_8718);
nand U9815 (N_9815,N_7193,N_6092);
nand U9816 (N_9816,N_7986,N_8611);
nor U9817 (N_9817,N_6550,N_6064);
nor U9818 (N_9818,N_6772,N_7032);
or U9819 (N_9819,N_6401,N_7581);
nor U9820 (N_9820,N_7139,N_6192);
nor U9821 (N_9821,N_7359,N_6288);
or U9822 (N_9822,N_7074,N_6855);
or U9823 (N_9823,N_8731,N_7722);
nand U9824 (N_9824,N_8924,N_7483);
or U9825 (N_9825,N_7764,N_8981);
nand U9826 (N_9826,N_6647,N_7500);
nor U9827 (N_9827,N_6193,N_7687);
or U9828 (N_9828,N_8516,N_7757);
nand U9829 (N_9829,N_6576,N_6264);
or U9830 (N_9830,N_8995,N_7781);
and U9831 (N_9831,N_8419,N_7052);
nor U9832 (N_9832,N_7463,N_8264);
nor U9833 (N_9833,N_7973,N_8293);
nand U9834 (N_9834,N_7901,N_7887);
and U9835 (N_9835,N_7702,N_7064);
nand U9836 (N_9836,N_8406,N_7458);
and U9837 (N_9837,N_7773,N_7422);
nand U9838 (N_9838,N_7314,N_8813);
nand U9839 (N_9839,N_7726,N_8128);
nand U9840 (N_9840,N_6537,N_6935);
or U9841 (N_9841,N_8742,N_6045);
and U9842 (N_9842,N_7058,N_7839);
or U9843 (N_9843,N_8084,N_6558);
nor U9844 (N_9844,N_8687,N_7030);
nand U9845 (N_9845,N_6043,N_6955);
nand U9846 (N_9846,N_6149,N_7423);
nor U9847 (N_9847,N_6432,N_6892);
and U9848 (N_9848,N_7397,N_6285);
nor U9849 (N_9849,N_7002,N_6714);
and U9850 (N_9850,N_7681,N_6691);
nor U9851 (N_9851,N_7648,N_8418);
and U9852 (N_9852,N_8215,N_6144);
or U9853 (N_9853,N_8443,N_6202);
or U9854 (N_9854,N_6517,N_7081);
nand U9855 (N_9855,N_7682,N_7760);
or U9856 (N_9856,N_8268,N_6489);
and U9857 (N_9857,N_6783,N_7065);
or U9858 (N_9858,N_7034,N_6490);
nor U9859 (N_9859,N_8164,N_8113);
or U9860 (N_9860,N_8861,N_8086);
and U9861 (N_9861,N_7779,N_7057);
and U9862 (N_9862,N_7187,N_8690);
and U9863 (N_9863,N_6281,N_7490);
and U9864 (N_9864,N_8385,N_7251);
nor U9865 (N_9865,N_7335,N_6244);
xnor U9866 (N_9866,N_6768,N_8466);
nor U9867 (N_9867,N_7294,N_7411);
or U9868 (N_9868,N_7053,N_7107);
nor U9869 (N_9869,N_8557,N_7451);
or U9870 (N_9870,N_7043,N_8088);
nand U9871 (N_9871,N_7796,N_8213);
nor U9872 (N_9872,N_6727,N_8751);
nand U9873 (N_9873,N_6809,N_8987);
or U9874 (N_9874,N_8144,N_7468);
and U9875 (N_9875,N_6392,N_6839);
or U9876 (N_9876,N_6894,N_6239);
nand U9877 (N_9877,N_7522,N_7152);
nor U9878 (N_9878,N_8370,N_7255);
nor U9879 (N_9879,N_6128,N_7023);
and U9880 (N_9880,N_7185,N_7001);
and U9881 (N_9881,N_8821,N_6814);
nor U9882 (N_9882,N_7102,N_8913);
nand U9883 (N_9883,N_7480,N_8628);
or U9884 (N_9884,N_8844,N_8506);
and U9885 (N_9885,N_6014,N_8230);
nor U9886 (N_9886,N_7374,N_8678);
or U9887 (N_9887,N_6913,N_6223);
nand U9888 (N_9888,N_8831,N_6575);
or U9889 (N_9889,N_6454,N_6529);
nand U9890 (N_9890,N_7039,N_6364);
and U9891 (N_9891,N_6856,N_7519);
and U9892 (N_9892,N_7616,N_7769);
or U9893 (N_9893,N_8536,N_8322);
and U9894 (N_9894,N_7605,N_8458);
or U9895 (N_9895,N_6555,N_6226);
nand U9896 (N_9896,N_7325,N_6372);
nand U9897 (N_9897,N_6276,N_8039);
nand U9898 (N_9898,N_8112,N_6637);
or U9899 (N_9899,N_8659,N_8361);
or U9900 (N_9900,N_6700,N_8272);
nor U9901 (N_9901,N_6949,N_8445);
nand U9902 (N_9902,N_8111,N_7861);
nand U9903 (N_9903,N_7379,N_8101);
and U9904 (N_9904,N_7734,N_7322);
nand U9905 (N_9905,N_7730,N_6466);
or U9906 (N_9906,N_6835,N_8793);
and U9907 (N_9907,N_8387,N_8943);
or U9908 (N_9908,N_7943,N_6658);
xor U9909 (N_9909,N_7569,N_7848);
or U9910 (N_9910,N_6762,N_7720);
xnor U9911 (N_9911,N_7402,N_6779);
nand U9912 (N_9912,N_8616,N_8222);
or U9913 (N_9913,N_8568,N_8721);
nor U9914 (N_9914,N_7471,N_7666);
and U9915 (N_9915,N_7731,N_8488);
and U9916 (N_9916,N_8608,N_6000);
or U9917 (N_9917,N_8094,N_7530);
and U9918 (N_9918,N_6333,N_7389);
and U9919 (N_9919,N_8808,N_7410);
nand U9920 (N_9920,N_6034,N_7536);
nand U9921 (N_9921,N_7100,N_7700);
and U9922 (N_9922,N_8026,N_7577);
and U9923 (N_9923,N_7346,N_6227);
or U9924 (N_9924,N_7188,N_7638);
nand U9925 (N_9925,N_8940,N_8986);
nor U9926 (N_9926,N_7088,N_6789);
nor U9927 (N_9927,N_6817,N_8745);
nor U9928 (N_9928,N_7755,N_8207);
nand U9929 (N_9929,N_6944,N_8763);
and U9930 (N_9930,N_7794,N_6327);
and U9931 (N_9931,N_8870,N_7395);
nor U9932 (N_9932,N_8460,N_7203);
or U9933 (N_9933,N_6473,N_8092);
nor U9934 (N_9934,N_8402,N_6138);
and U9935 (N_9935,N_7517,N_6496);
or U9936 (N_9936,N_6642,N_6616);
and U9937 (N_9937,N_7918,N_8554);
nor U9938 (N_9938,N_6278,N_6229);
nor U9939 (N_9939,N_7518,N_6992);
or U9940 (N_9940,N_7563,N_6126);
or U9941 (N_9941,N_7261,N_6341);
nor U9942 (N_9942,N_7194,N_6812);
and U9943 (N_9943,N_6819,N_6331);
nand U9944 (N_9944,N_7944,N_8284);
and U9945 (N_9945,N_8931,N_6487);
nor U9946 (N_9946,N_8685,N_6533);
nor U9947 (N_9947,N_8580,N_7721);
nand U9948 (N_9948,N_7842,N_7338);
nand U9949 (N_9949,N_6470,N_6998);
and U9950 (N_9950,N_8129,N_6217);
and U9951 (N_9951,N_7762,N_8896);
nand U9952 (N_9952,N_6585,N_6294);
nor U9953 (N_9953,N_6011,N_7050);
or U9954 (N_9954,N_8639,N_7677);
nand U9955 (N_9955,N_8917,N_8108);
nand U9956 (N_9956,N_6769,N_7363);
nor U9957 (N_9957,N_7205,N_8604);
or U9958 (N_9958,N_8897,N_8710);
nor U9959 (N_9959,N_8099,N_7211);
nor U9960 (N_9960,N_7907,N_8672);
and U9961 (N_9961,N_7284,N_6316);
and U9962 (N_9962,N_7077,N_8848);
nor U9963 (N_9963,N_7176,N_6614);
or U9964 (N_9964,N_7243,N_6863);
and U9965 (N_9965,N_8841,N_7639);
nand U9966 (N_9966,N_8610,N_8972);
nand U9967 (N_9967,N_8723,N_8586);
nand U9968 (N_9968,N_8809,N_8919);
nand U9969 (N_9969,N_6523,N_6947);
or U9970 (N_9970,N_7170,N_6390);
or U9971 (N_9971,N_6350,N_6286);
nor U9972 (N_9972,N_8175,N_6493);
nor U9973 (N_9973,N_8523,N_6093);
and U9974 (N_9974,N_7645,N_6837);
or U9975 (N_9975,N_7552,N_6087);
nand U9976 (N_9976,N_7909,N_6381);
nor U9977 (N_9977,N_8062,N_8158);
and U9978 (N_9978,N_8771,N_6685);
nand U9979 (N_9979,N_6920,N_7856);
and U9980 (N_9980,N_7061,N_8575);
or U9981 (N_9981,N_6317,N_8189);
nor U9982 (N_9982,N_6256,N_6120);
or U9983 (N_9983,N_7558,N_6966);
nor U9984 (N_9984,N_6790,N_8141);
nand U9985 (N_9985,N_7695,N_6100);
and U9986 (N_9986,N_6967,N_6251);
nor U9987 (N_9987,N_6731,N_6036);
and U9988 (N_9988,N_8714,N_6357);
or U9989 (N_9989,N_8514,N_6356);
nand U9990 (N_9990,N_8656,N_6116);
nand U9991 (N_9991,N_6624,N_8163);
and U9992 (N_9992,N_7697,N_6521);
nor U9993 (N_9993,N_6938,N_7524);
nand U9994 (N_9994,N_6950,N_6600);
or U9995 (N_9995,N_7770,N_8004);
and U9996 (N_9996,N_8918,N_6596);
nor U9997 (N_9997,N_8569,N_7362);
or U9998 (N_9998,N_7903,N_8904);
or U9999 (N_9999,N_8104,N_8635);
nor U10000 (N_10000,N_7643,N_8859);
nor U10001 (N_10001,N_8537,N_8744);
and U10002 (N_10002,N_8287,N_8291);
and U10003 (N_10003,N_8814,N_6586);
or U10004 (N_10004,N_8117,N_8276);
and U10005 (N_10005,N_7456,N_7812);
and U10006 (N_10006,N_7873,N_6032);
and U10007 (N_10007,N_8180,N_6154);
nor U10008 (N_10008,N_7169,N_8273);
or U10009 (N_10009,N_6210,N_8126);
nor U10010 (N_10010,N_7520,N_8243);
nand U10011 (N_10011,N_6215,N_6314);
nand U10012 (N_10012,N_6669,N_6216);
or U10013 (N_10013,N_8011,N_7803);
nand U10014 (N_10014,N_8512,N_6335);
nor U10015 (N_10015,N_6921,N_8017);
nor U10016 (N_10016,N_6480,N_7332);
and U10017 (N_10017,N_6535,N_6445);
or U10018 (N_10018,N_7679,N_6142);
nor U10019 (N_10019,N_8280,N_8879);
nand U10020 (N_10020,N_7975,N_7240);
nand U10021 (N_10021,N_8033,N_6538);
nand U10022 (N_10022,N_6875,N_6347);
nor U10023 (N_10023,N_6615,N_6119);
nand U10024 (N_10024,N_8719,N_6908);
nand U10025 (N_10025,N_8717,N_6798);
nor U10026 (N_10026,N_7962,N_8393);
and U10027 (N_10027,N_7782,N_7559);
nor U10028 (N_10028,N_6853,N_6326);
nand U10029 (N_10029,N_6058,N_7749);
or U10030 (N_10030,N_6237,N_6475);
nand U10031 (N_10031,N_7557,N_7632);
nor U10032 (N_10032,N_8364,N_8966);
nand U10033 (N_10033,N_7095,N_8357);
nor U10034 (N_10034,N_6150,N_7465);
or U10035 (N_10035,N_7242,N_7891);
nor U10036 (N_10036,N_7972,N_8590);
nand U10037 (N_10037,N_6451,N_6167);
nand U10038 (N_10038,N_6716,N_7324);
and U10039 (N_10039,N_6958,N_8507);
or U10040 (N_10040,N_7186,N_8941);
or U10041 (N_10041,N_6682,N_8269);
nor U10042 (N_10042,N_8785,N_8874);
nand U10043 (N_10043,N_7894,N_6829);
nor U10044 (N_10044,N_7272,N_6959);
xnor U10045 (N_10045,N_7250,N_7008);
nand U10046 (N_10046,N_8139,N_6651);
nand U10047 (N_10047,N_6205,N_7550);
nand U10048 (N_10048,N_7384,N_8627);
or U10049 (N_10049,N_8417,N_7393);
nor U10050 (N_10050,N_6081,N_6918);
or U10051 (N_10051,N_6634,N_7371);
or U10052 (N_10052,N_8559,N_7595);
nor U10053 (N_10053,N_6857,N_8733);
or U10054 (N_10054,N_7476,N_6582);
or U10055 (N_10055,N_8354,N_6971);
nand U10056 (N_10056,N_7262,N_8499);
nand U10057 (N_10057,N_8327,N_6076);
nand U10058 (N_10058,N_7995,N_7189);
or U10059 (N_10059,N_6444,N_8726);
or U10060 (N_10060,N_6003,N_7979);
nand U10061 (N_10061,N_6240,N_7115);
or U10062 (N_10062,N_6749,N_7112);
nand U10063 (N_10063,N_7469,N_8147);
or U10064 (N_10064,N_6635,N_6541);
and U10065 (N_10065,N_6323,N_8343);
nor U10066 (N_10066,N_8976,N_6879);
or U10067 (N_10067,N_8075,N_7281);
or U10068 (N_10068,N_8348,N_8251);
or U10069 (N_10069,N_7963,N_7288);
nor U10070 (N_10070,N_8903,N_7818);
nand U10071 (N_10071,N_6059,N_7629);
nand U10072 (N_10072,N_8502,N_6260);
nand U10073 (N_10073,N_6688,N_7264);
or U10074 (N_10074,N_7735,N_8588);
nor U10075 (N_10075,N_8161,N_7360);
nor U10076 (N_10076,N_8907,N_6374);
or U10077 (N_10077,N_8812,N_7234);
or U10078 (N_10078,N_7271,N_7308);
nand U10079 (N_10079,N_8893,N_8048);
or U10080 (N_10080,N_7754,N_7732);
nor U10081 (N_10081,N_6698,N_7857);
nand U10082 (N_10082,N_7390,N_8735);
or U10083 (N_10083,N_8345,N_8762);
nand U10084 (N_10084,N_8951,N_8546);
nand U10085 (N_10085,N_6990,N_6954);
or U10086 (N_10086,N_7835,N_8683);
nand U10087 (N_10087,N_7940,N_7613);
nor U10088 (N_10088,N_7976,N_8259);
or U10089 (N_10089,N_7149,N_8730);
and U10090 (N_10090,N_6979,N_6282);
and U10091 (N_10091,N_8855,N_6114);
and U10092 (N_10092,N_7383,N_7285);
or U10093 (N_10093,N_7872,N_8541);
nor U10094 (N_10094,N_8789,N_6170);
and U10095 (N_10095,N_7354,N_7106);
or U10096 (N_10096,N_6888,N_6823);
nand U10097 (N_10097,N_8816,N_8383);
nand U10098 (N_10098,N_6321,N_6633);
and U10099 (N_10099,N_8152,N_7660);
or U10100 (N_10100,N_7159,N_7200);
and U10101 (N_10101,N_6067,N_7598);
nand U10102 (N_10102,N_8035,N_6053);
and U10103 (N_10103,N_8063,N_7742);
nand U10104 (N_10104,N_7505,N_8832);
or U10105 (N_10105,N_6878,N_8949);
nand U10106 (N_10106,N_7403,N_8124);
and U10107 (N_10107,N_7706,N_7531);
and U10108 (N_10108,N_7388,N_6359);
nor U10109 (N_10109,N_6112,N_7038);
nor U10110 (N_10110,N_6662,N_8508);
or U10111 (N_10111,N_6026,N_6152);
nor U10112 (N_10112,N_8652,N_8964);
or U10113 (N_10113,N_8328,N_6568);
or U10114 (N_10114,N_6219,N_6931);
and U10115 (N_10115,N_7274,N_6398);
nor U10116 (N_10116,N_6832,N_6182);
nand U10117 (N_10117,N_6748,N_8650);
and U10118 (N_10118,N_6062,N_6665);
nor U10119 (N_10119,N_7419,N_7266);
nand U10120 (N_10120,N_6564,N_6021);
nor U10121 (N_10121,N_7101,N_8962);
nor U10122 (N_10122,N_8648,N_7391);
nor U10123 (N_10123,N_7054,N_6883);
and U10124 (N_10124,N_8055,N_7435);
nand U10125 (N_10125,N_8743,N_7729);
and U10126 (N_10126,N_7840,N_8205);
nor U10127 (N_10127,N_8493,N_7527);
nor U10128 (N_10128,N_7914,N_7482);
nor U10129 (N_10129,N_7895,N_8827);
or U10130 (N_10130,N_7686,N_8110);
nand U10131 (N_10131,N_6370,N_7784);
nor U10132 (N_10132,N_8165,N_6776);
nor U10133 (N_10133,N_7260,N_6255);
and U10134 (N_10134,N_8607,N_7173);
or U10135 (N_10135,N_8399,N_7025);
nand U10136 (N_10136,N_7367,N_6383);
nand U10137 (N_10137,N_8952,N_6619);
or U10138 (N_10138,N_6423,N_7493);
nand U10139 (N_10139,N_6720,N_6854);
and U10140 (N_10140,N_8219,N_7771);
nor U10141 (N_10141,N_7369,N_6887);
xor U10142 (N_10142,N_6672,N_7604);
nor U10143 (N_10143,N_6195,N_7816);
and U10144 (N_10144,N_8051,N_8660);
and U10145 (N_10145,N_8212,N_8356);
nand U10146 (N_10146,N_8863,N_7191);
or U10147 (N_10147,N_8732,N_6660);
or U10148 (N_10148,N_7376,N_7627);
nor U10149 (N_10149,N_7204,N_8107);
nor U10150 (N_10150,N_8186,N_6376);
and U10151 (N_10151,N_6670,N_8926);
and U10152 (N_10152,N_8697,N_6024);
or U10153 (N_10153,N_6513,N_8329);
or U10154 (N_10154,N_8617,N_7543);
nor U10155 (N_10155,N_6957,N_6272);
nor U10156 (N_10156,N_6344,N_7561);
or U10157 (N_10157,N_7485,N_8123);
nor U10158 (N_10158,N_8644,N_8314);
nand U10159 (N_10159,N_6654,N_8315);
or U10160 (N_10160,N_8166,N_8716);
nand U10161 (N_10161,N_7556,N_7626);
or U10162 (N_10162,N_8349,N_7130);
nor U10163 (N_10163,N_6439,N_8184);
nand U10164 (N_10164,N_8025,N_8249);
or U10165 (N_10165,N_6441,N_7801);
nand U10166 (N_10166,N_7711,N_8817);
nand U10167 (N_10167,N_7287,N_8262);
or U10168 (N_10168,N_8258,N_7415);
or U10169 (N_10169,N_7671,N_7588);
or U10170 (N_10170,N_7725,N_7640);
and U10171 (N_10171,N_7016,N_8226);
or U10172 (N_10172,N_8626,N_8532);
and U10173 (N_10173,N_7124,N_8738);
or U10174 (N_10174,N_6085,N_6485);
nand U10175 (N_10175,N_6242,N_8253);
nor U10176 (N_10176,N_7820,N_8886);
nor U10177 (N_10177,N_6804,N_8006);
and U10178 (N_10178,N_6190,N_8566);
and U10179 (N_10179,N_6934,N_6699);
nand U10180 (N_10180,N_8806,N_8594);
or U10181 (N_10181,N_7925,N_8211);
nand U10182 (N_10182,N_6060,N_7444);
nand U10183 (N_10183,N_6695,N_7896);
and U10184 (N_10184,N_7688,N_6791);
and U10185 (N_10185,N_8022,N_8970);
nor U10186 (N_10186,N_6579,N_7824);
nand U10187 (N_10187,N_8824,N_6595);
nor U10188 (N_10188,N_8655,N_8305);
nor U10189 (N_10189,N_7080,N_8150);
and U10190 (N_10190,N_8073,N_7810);
nor U10191 (N_10191,N_6503,N_6681);
nor U10192 (N_10192,N_8770,N_8873);
nand U10193 (N_10193,N_6328,N_8487);
nor U10194 (N_10194,N_6677,N_6903);
nor U10195 (N_10195,N_6771,N_8244);
nor U10196 (N_10196,N_7571,N_8061);
or U10197 (N_10197,N_6426,N_7060);
nand U10198 (N_10198,N_7791,N_6793);
nor U10199 (N_10199,N_7656,N_8505);
or U10200 (N_10200,N_7161,N_8646);
nor U10201 (N_10201,N_6626,N_6502);
nor U10202 (N_10202,N_7238,N_6380);
nand U10203 (N_10203,N_6450,N_6425);
nor U10204 (N_10204,N_6926,N_8709);
nor U10205 (N_10205,N_7833,N_6828);
nor U10206 (N_10206,N_7787,N_8153);
and U10207 (N_10207,N_8694,N_8515);
or U10208 (N_10208,N_8457,N_8794);
nand U10209 (N_10209,N_8642,N_8740);
nand U10210 (N_10210,N_6165,N_8713);
nor U10211 (N_10211,N_8857,N_6743);
and U10212 (N_10212,N_7758,N_8592);
nand U10213 (N_10213,N_8891,N_6650);
nor U10214 (N_10214,N_8768,N_6009);
and U10215 (N_10215,N_7751,N_8203);
nor U10216 (N_10216,N_7680,N_7586);
nor U10217 (N_10217,N_7541,N_6206);
and U10218 (N_10218,N_6876,N_6049);
or U10219 (N_10219,N_8095,N_6759);
nor U10220 (N_10220,N_7763,N_7603);
nor U10221 (N_10221,N_8561,N_6291);
and U10222 (N_10222,N_6448,N_8948);
nor U10223 (N_10223,N_8056,N_6332);
nor U10224 (N_10224,N_6613,N_8375);
or U10225 (N_10225,N_7712,N_6877);
nor U10226 (N_10226,N_6522,N_6110);
nand U10227 (N_10227,N_6180,N_6184);
nand U10228 (N_10228,N_7548,N_8079);
or U10229 (N_10229,N_6978,N_8593);
nor U10230 (N_10230,N_7683,N_8823);
xnor U10231 (N_10231,N_8068,N_6137);
nand U10232 (N_10232,N_8066,N_7174);
or U10233 (N_10233,N_7587,N_8758);
nand U10234 (N_10234,N_7455,N_7759);
and U10235 (N_10235,N_6422,N_8992);
nor U10236 (N_10236,N_7690,N_8999);
or U10237 (N_10237,N_8472,N_8334);
nand U10238 (N_10238,N_7368,N_6737);
nand U10239 (N_10239,N_8058,N_6563);
and U10240 (N_10240,N_6981,N_8444);
and U10241 (N_10241,N_8872,N_8303);
nand U10242 (N_10242,N_7506,N_6545);
and U10243 (N_10243,N_7171,N_6279);
nand U10244 (N_10244,N_8779,N_8240);
and U10245 (N_10245,N_8201,N_6663);
xor U10246 (N_10246,N_6528,N_6932);
or U10247 (N_10247,N_8729,N_7653);
or U10248 (N_10248,N_7737,N_8983);
and U10249 (N_10249,N_6241,N_7024);
nand U10250 (N_10250,N_7460,N_8822);
nor U10251 (N_10251,N_7659,N_8858);
and U10252 (N_10252,N_6136,N_6232);
nor U10253 (N_10253,N_7167,N_6844);
or U10254 (N_10254,N_7699,N_6852);
or U10255 (N_10255,N_7983,N_6105);
nand U10256 (N_10256,N_6127,N_8248);
or U10257 (N_10257,N_8686,N_6816);
and U10258 (N_10258,N_8587,N_6703);
or U10259 (N_10259,N_6580,N_6547);
nand U10260 (N_10260,N_7296,N_8597);
nor U10261 (N_10261,N_8455,N_6213);
nor U10262 (N_10262,N_8267,N_6553);
nor U10263 (N_10263,N_6859,N_8245);
nand U10264 (N_10264,N_6483,N_6109);
nor U10265 (N_10265,N_6801,N_7974);
nand U10266 (N_10266,N_6657,N_8330);
xor U10267 (N_10267,N_7249,N_7685);
nor U10268 (N_10268,N_7938,N_6505);
or U10269 (N_10269,N_6046,N_8185);
nand U10270 (N_10270,N_8031,N_6655);
nand U10271 (N_10271,N_6221,N_8202);
nand U10272 (N_10272,N_6925,N_6484);
nand U10273 (N_10273,N_8871,N_8968);
nor U10274 (N_10274,N_8181,N_8704);
nand U10275 (N_10275,N_7443,N_7142);
or U10276 (N_10276,N_6948,N_7385);
or U10277 (N_10277,N_8156,N_6974);
and U10278 (N_10278,N_7927,N_8261);
nand U10279 (N_10279,N_6041,N_6082);
and U10280 (N_10280,N_8431,N_7007);
nand U10281 (N_10281,N_6160,N_6800);
nand U10282 (N_10282,N_6435,N_6792);
or U10283 (N_10283,N_6004,N_6977);
or U10284 (N_10284,N_6639,N_8528);
or U10285 (N_10285,N_7709,N_6070);
and U10286 (N_10286,N_7241,N_6429);
and U10287 (N_10287,N_6591,N_7356);
nand U10288 (N_10288,N_8121,N_6228);
and U10289 (N_10289,N_8242,N_8130);
nor U10290 (N_10290,N_8947,N_8728);
and U10291 (N_10291,N_6130,N_6787);
nor U10292 (N_10292,N_8715,N_6831);
nor U10293 (N_10293,N_6419,N_8311);
and U10294 (N_10294,N_6516,N_6309);
or U10295 (N_10295,N_8426,N_7647);
nor U10296 (N_10296,N_8925,N_8324);
nor U10297 (N_10297,N_6807,N_6300);
and U10298 (N_10298,N_6245,N_6741);
nand U10299 (N_10299,N_8826,N_6858);
nor U10300 (N_10300,N_7678,N_8556);
nand U10301 (N_10301,N_8811,N_7378);
nand U10302 (N_10302,N_8359,N_7183);
and U10303 (N_10303,N_6713,N_8669);
or U10304 (N_10304,N_7544,N_6539);
and U10305 (N_10305,N_8838,N_7915);
or U10306 (N_10306,N_7484,N_8231);
nor U10307 (N_10307,N_6738,N_7256);
nor U10308 (N_10308,N_6479,N_6431);
or U10309 (N_10309,N_7210,N_7344);
and U10310 (N_10310,N_6002,N_8325);
nor U10311 (N_10311,N_6056,N_6795);
nor U10312 (N_10312,N_8631,N_8397);
nor U10313 (N_10313,N_8227,N_6301);
xnor U10314 (N_10314,N_8736,N_7128);
or U10315 (N_10315,N_7507,N_7691);
and U10316 (N_10316,N_7224,N_6354);
and U10317 (N_10317,N_8338,N_8599);
and U10318 (N_10318,N_8494,N_8252);
or U10319 (N_10319,N_6895,N_8737);
or U10320 (N_10320,N_8480,N_8946);
nand U10321 (N_10321,N_7765,N_6899);
or U10322 (N_10322,N_6253,N_7236);
nor U10323 (N_10323,N_8365,N_8415);
and U10324 (N_10324,N_8560,N_6211);
nand U10325 (N_10325,N_8247,N_8002);
nor U10326 (N_10326,N_8299,N_6746);
and U10327 (N_10327,N_6266,N_6929);
and U10328 (N_10328,N_6525,N_8490);
nor U10329 (N_10329,N_7580,N_6181);
nand U10330 (N_10330,N_8906,N_6225);
nor U10331 (N_10331,N_6840,N_7092);
or U10332 (N_10332,N_6704,N_8675);
nor U10333 (N_10333,N_7723,N_8503);
nor U10334 (N_10334,N_6106,N_7597);
nand U10335 (N_10335,N_7777,N_7501);
nor U10336 (N_10336,N_8394,N_6139);
nor U10337 (N_10337,N_8802,N_6103);
nand U10338 (N_10338,N_8034,N_7498);
nor U10339 (N_10339,N_8290,N_8390);
nor U10340 (N_10340,N_7079,N_8191);
or U10341 (N_10341,N_7615,N_6617);
and U10342 (N_10342,N_6172,N_6813);
nand U10343 (N_10343,N_7767,N_7703);
nand U10344 (N_10344,N_8080,N_6068);
nor U10345 (N_10345,N_6989,N_7361);
nor U10346 (N_10346,N_8256,N_8674);
and U10347 (N_10347,N_8000,N_6393);
and U10348 (N_10348,N_6612,N_7502);
nor U10349 (N_10349,N_6297,N_7797);
nor U10350 (N_10350,N_6177,N_7611);
nor U10351 (N_10351,N_6970,N_6796);
nand U10352 (N_10352,N_6874,N_8388);
or U10353 (N_10353,N_8640,N_8820);
and U10354 (N_10354,N_7635,N_6756);
nand U10355 (N_10355,N_8398,N_7804);
nand U10356 (N_10356,N_8564,N_7197);
nand U10357 (N_10357,N_8845,N_6821);
and U10358 (N_10358,N_7350,N_8661);
nor U10359 (N_10359,N_7134,N_6025);
and U10360 (N_10360,N_6437,N_6262);
and U10361 (N_10361,N_7252,N_6694);
nand U10362 (N_10362,N_6566,N_8091);
nand U10363 (N_10363,N_6818,N_7871);
or U10364 (N_10364,N_8429,N_7220);
nor U10365 (N_10365,N_7154,N_8373);
nand U10366 (N_10366,N_6554,N_7805);
nor U10367 (N_10367,N_7838,N_6214);
nor U10368 (N_10368,N_7097,N_7028);
or U10369 (N_10369,N_7956,N_8351);
nand U10370 (N_10370,N_8955,N_6953);
or U10371 (N_10371,N_8059,N_7339);
nor U10372 (N_10372,N_7293,N_8828);
or U10373 (N_10373,N_8539,N_8747);
or U10374 (N_10374,N_6094,N_8862);
nor U10375 (N_10375,N_6033,N_7071);
nor U10376 (N_10376,N_8474,N_8883);
nor U10377 (N_10377,N_8531,N_8131);
or U10378 (N_10378,N_7792,N_7593);
nor U10379 (N_10379,N_6178,N_8404);
nor U10380 (N_10380,N_8321,N_6433);
nand U10381 (N_10381,N_6946,N_8193);
nor U10382 (N_10382,N_6259,N_8469);
nor U10383 (N_10383,N_6416,N_6097);
and U10384 (N_10384,N_7047,N_8223);
nor U10385 (N_10385,N_8800,N_8934);
or U10386 (N_10386,N_6498,N_7996);
nand U10387 (N_10387,N_7555,N_8347);
nor U10388 (N_10388,N_6805,N_8614);
and U10389 (N_10389,N_8562,N_8143);
or U10390 (N_10390,N_6960,N_7882);
or U10391 (N_10391,N_6394,N_6430);
or U10392 (N_10392,N_8724,N_6905);
or U10393 (N_10393,N_7333,N_7318);
and U10394 (N_10394,N_7885,N_6900);
and U10395 (N_10395,N_7841,N_8029);
and U10396 (N_10396,N_8708,N_8850);
and U10397 (N_10397,N_7939,N_6622);
and U10398 (N_10398,N_6534,N_6661);
nand U10399 (N_10399,N_7404,N_6597);
nor U10400 (N_10400,N_8605,N_7408);
or U10401 (N_10401,N_7425,N_7744);
nor U10402 (N_10402,N_7978,N_8711);
nand U10403 (N_10403,N_7814,N_6740);
or U10404 (N_10404,N_7265,N_7535);
or U10405 (N_10405,N_8912,N_8534);
nor U10406 (N_10406,N_7738,N_7438);
nand U10407 (N_10407,N_8064,N_7479);
and U10408 (N_10408,N_8013,N_8504);
nor U10409 (N_10409,N_7094,N_7329);
and U10410 (N_10410,N_7572,N_7428);
nor U10411 (N_10411,N_7510,N_6488);
and U10412 (N_10412,N_7466,N_8050);
and U10413 (N_10413,N_8216,N_6176);
nor U10414 (N_10414,N_6885,N_8521);
nand U10415 (N_10415,N_6248,N_7421);
or U10416 (N_10416,N_6747,N_8777);
or U10417 (N_10417,N_6862,N_7941);
and U10418 (N_10418,N_6476,N_8865);
or U10419 (N_10419,N_7594,N_6587);
and U10420 (N_10420,N_8788,N_6758);
and U10421 (N_10421,N_7093,N_6040);
nor U10422 (N_10422,N_6578,N_7033);
and U10423 (N_10423,N_7931,N_8384);
and U10424 (N_10424,N_7987,N_6782);
nor U10425 (N_10425,N_7246,N_8263);
nor U10426 (N_10426,N_6099,N_7044);
or U10427 (N_10427,N_6198,N_6693);
or U10428 (N_10428,N_7005,N_6157);
nand U10429 (N_10429,N_8851,N_7642);
nand U10430 (N_10430,N_7162,N_8221);
nor U10431 (N_10431,N_6384,N_6794);
and U10432 (N_10432,N_6656,N_6625);
or U10433 (N_10433,N_6933,N_6806);
or U10434 (N_10434,N_7932,N_7177);
nor U10435 (N_10435,N_6560,N_8549);
nand U10436 (N_10436,N_6113,N_6825);
nand U10437 (N_10437,N_8015,N_6640);
and U10438 (N_10438,N_7508,N_7375);
nand U10439 (N_10439,N_7768,N_7129);
or U10440 (N_10440,N_8009,N_8993);
nand U10441 (N_10441,N_8901,N_8741);
and U10442 (N_10442,N_8183,N_6898);
and U10443 (N_10443,N_6906,N_8780);
nor U10444 (N_10444,N_8998,N_6201);
nand U10445 (N_10445,N_8209,N_7300);
or U10446 (N_10446,N_8555,N_8188);
and U10447 (N_10447,N_6397,N_8074);
and U10448 (N_10448,N_6659,N_8632);
and U10449 (N_10449,N_8392,N_6962);
or U10450 (N_10450,N_6983,N_6101);
nor U10451 (N_10451,N_6543,N_8676);
or U10452 (N_10452,N_7003,N_6915);
nor U10453 (N_10453,N_7453,N_6283);
or U10454 (N_10454,N_7295,N_8761);
and U10455 (N_10455,N_8220,N_6511);
nand U10456 (N_10456,N_6602,N_7778);
or U10457 (N_10457,N_6005,N_7612);
nand U10458 (N_10458,N_7977,N_6442);
nand U10459 (N_10459,N_6599,N_6209);
and U10460 (N_10460,N_8991,N_7698);
nand U10461 (N_10461,N_7529,N_6822);
nand U10462 (N_10462,N_8237,N_7672);
nor U10463 (N_10463,N_6186,N_8584);
and U10464 (N_10464,N_7990,N_6133);
nor U10465 (N_10465,N_8565,N_6188);
nor U10466 (N_10466,N_7059,N_8282);
and U10467 (N_10467,N_8937,N_7670);
nand U10468 (N_10468,N_8204,N_8134);
and U10469 (N_10469,N_7574,N_8122);
nor U10470 (N_10470,N_6562,N_8046);
nor U10471 (N_10471,N_6988,N_7537);
and U10472 (N_10472,N_8440,N_7441);
nor U10473 (N_10473,N_7634,N_7745);
nor U10474 (N_10474,N_7823,N_6508);
nor U10475 (N_10475,N_6086,N_8235);
or U10476 (N_10476,N_8149,N_8520);
nand U10477 (N_10477,N_7628,N_8849);
and U10478 (N_10478,N_7920,N_7492);
and U10479 (N_10479,N_6191,N_7809);
or U10480 (N_10480,N_7554,N_8920);
and U10481 (N_10481,N_8673,N_8550);
nand U10482 (N_10482,N_6636,N_7062);
and U10483 (N_10483,N_8668,N_8198);
nand U10484 (N_10484,N_7437,N_7798);
or U10485 (N_10485,N_6901,N_8471);
nand U10486 (N_10486,N_8496,N_8428);
or U10487 (N_10487,N_8790,N_7740);
nand U10488 (N_10488,N_6312,N_8734);
or U10489 (N_10489,N_6163,N_8255);
or U10490 (N_10490,N_8410,N_6739);
or U10491 (N_10491,N_6750,N_8578);
and U10492 (N_10492,N_6902,N_6406);
nor U10493 (N_10493,N_6080,N_7899);
or U10494 (N_10494,N_8371,N_7280);
nor U10495 (N_10495,N_6273,N_6197);
xor U10496 (N_10496,N_6031,N_7728);
nand U10497 (N_10497,N_7921,N_8395);
nand U10498 (N_10498,N_8168,N_6530);
nand U10499 (N_10499,N_8739,N_6629);
nor U10500 (N_10500,N_7592,N_6580);
and U10501 (N_10501,N_6376,N_7138);
or U10502 (N_10502,N_7760,N_8266);
or U10503 (N_10503,N_8284,N_7951);
and U10504 (N_10504,N_7064,N_8229);
nor U10505 (N_10505,N_7684,N_7971);
nor U10506 (N_10506,N_8432,N_6910);
or U10507 (N_10507,N_7630,N_6918);
or U10508 (N_10508,N_8638,N_7439);
and U10509 (N_10509,N_8524,N_7602);
or U10510 (N_10510,N_6583,N_6054);
nand U10511 (N_10511,N_7433,N_6185);
nand U10512 (N_10512,N_7658,N_8326);
and U10513 (N_10513,N_7571,N_8812);
and U10514 (N_10514,N_7634,N_6532);
and U10515 (N_10515,N_7170,N_8803);
nand U10516 (N_10516,N_8343,N_8822);
nor U10517 (N_10517,N_7561,N_7633);
nor U10518 (N_10518,N_8868,N_8833);
or U10519 (N_10519,N_7311,N_6543);
nor U10520 (N_10520,N_7050,N_8606);
and U10521 (N_10521,N_6215,N_8020);
and U10522 (N_10522,N_8622,N_8809);
nand U10523 (N_10523,N_8423,N_8421);
or U10524 (N_10524,N_8198,N_6682);
nand U10525 (N_10525,N_8480,N_6197);
nand U10526 (N_10526,N_6546,N_8486);
nor U10527 (N_10527,N_8537,N_8507);
or U10528 (N_10528,N_7118,N_8868);
nand U10529 (N_10529,N_7343,N_7722);
or U10530 (N_10530,N_6333,N_8343);
nor U10531 (N_10531,N_7881,N_8615);
and U10532 (N_10532,N_6252,N_6197);
and U10533 (N_10533,N_8403,N_8400);
and U10534 (N_10534,N_7477,N_7203);
nand U10535 (N_10535,N_6164,N_7198);
xor U10536 (N_10536,N_7003,N_8687);
nor U10537 (N_10537,N_6065,N_7091);
or U10538 (N_10538,N_7900,N_8336);
and U10539 (N_10539,N_8874,N_6144);
and U10540 (N_10540,N_6207,N_8523);
nand U10541 (N_10541,N_6214,N_6116);
nor U10542 (N_10542,N_8302,N_6494);
and U10543 (N_10543,N_8808,N_6453);
and U10544 (N_10544,N_8668,N_7695);
nor U10545 (N_10545,N_6326,N_6290);
xor U10546 (N_10546,N_7308,N_6456);
and U10547 (N_10547,N_7588,N_8176);
nand U10548 (N_10548,N_7010,N_6536);
or U10549 (N_10549,N_6070,N_7329);
nand U10550 (N_10550,N_6542,N_8384);
nand U10551 (N_10551,N_7913,N_8015);
nor U10552 (N_10552,N_8393,N_6670);
and U10553 (N_10553,N_7581,N_7315);
nor U10554 (N_10554,N_8509,N_8970);
nand U10555 (N_10555,N_6140,N_7614);
nor U10556 (N_10556,N_8114,N_6470);
nand U10557 (N_10557,N_8901,N_8408);
nor U10558 (N_10558,N_8687,N_7848);
nand U10559 (N_10559,N_6031,N_7365);
nand U10560 (N_10560,N_8807,N_7086);
nor U10561 (N_10561,N_8829,N_7608);
or U10562 (N_10562,N_8572,N_8894);
nor U10563 (N_10563,N_8798,N_6710);
or U10564 (N_10564,N_7591,N_6760);
or U10565 (N_10565,N_6376,N_6667);
nor U10566 (N_10566,N_7781,N_8332);
nand U10567 (N_10567,N_6348,N_7255);
and U10568 (N_10568,N_7480,N_7977);
and U10569 (N_10569,N_7955,N_6223);
or U10570 (N_10570,N_7821,N_8269);
or U10571 (N_10571,N_6976,N_6433);
nor U10572 (N_10572,N_7581,N_6540);
nor U10573 (N_10573,N_8114,N_7191);
nand U10574 (N_10574,N_7951,N_7717);
nand U10575 (N_10575,N_8475,N_8291);
and U10576 (N_10576,N_8139,N_7001);
nand U10577 (N_10577,N_6765,N_7379);
nor U10578 (N_10578,N_6447,N_8637);
nor U10579 (N_10579,N_8135,N_6357);
nand U10580 (N_10580,N_7883,N_7062);
nor U10581 (N_10581,N_8964,N_7500);
or U10582 (N_10582,N_8953,N_8281);
and U10583 (N_10583,N_6537,N_7753);
nor U10584 (N_10584,N_8307,N_6162);
or U10585 (N_10585,N_7011,N_6265);
nand U10586 (N_10586,N_6007,N_7075);
and U10587 (N_10587,N_8087,N_6174);
and U10588 (N_10588,N_6060,N_7611);
nor U10589 (N_10589,N_6772,N_8854);
and U10590 (N_10590,N_8711,N_6514);
or U10591 (N_10591,N_8114,N_6811);
nand U10592 (N_10592,N_6720,N_6299);
or U10593 (N_10593,N_6268,N_7082);
and U10594 (N_10594,N_8952,N_8586);
nand U10595 (N_10595,N_8745,N_6579);
nor U10596 (N_10596,N_7022,N_6840);
nand U10597 (N_10597,N_8391,N_6192);
and U10598 (N_10598,N_7721,N_8430);
or U10599 (N_10599,N_8973,N_8849);
or U10600 (N_10600,N_6225,N_8453);
nor U10601 (N_10601,N_7026,N_7473);
xnor U10602 (N_10602,N_7504,N_8857);
nand U10603 (N_10603,N_7972,N_7308);
nand U10604 (N_10604,N_8805,N_6916);
nor U10605 (N_10605,N_8520,N_7389);
nor U10606 (N_10606,N_8522,N_8436);
nor U10607 (N_10607,N_7139,N_8691);
and U10608 (N_10608,N_8165,N_8892);
nand U10609 (N_10609,N_8290,N_8058);
and U10610 (N_10610,N_8195,N_7175);
nand U10611 (N_10611,N_8000,N_7116);
and U10612 (N_10612,N_6597,N_7333);
and U10613 (N_10613,N_6172,N_7541);
and U10614 (N_10614,N_8164,N_7865);
or U10615 (N_10615,N_7758,N_6324);
nand U10616 (N_10616,N_8931,N_7985);
or U10617 (N_10617,N_7882,N_6929);
nor U10618 (N_10618,N_6249,N_7489);
nand U10619 (N_10619,N_8139,N_7828);
nand U10620 (N_10620,N_7302,N_7797);
nand U10621 (N_10621,N_6973,N_8122);
nand U10622 (N_10622,N_6394,N_8662);
nand U10623 (N_10623,N_6844,N_6104);
and U10624 (N_10624,N_8189,N_6141);
or U10625 (N_10625,N_7497,N_8152);
and U10626 (N_10626,N_8950,N_8124);
nand U10627 (N_10627,N_7251,N_8169);
or U10628 (N_10628,N_6583,N_7027);
nor U10629 (N_10629,N_6235,N_6292);
nor U10630 (N_10630,N_8310,N_8741);
nor U10631 (N_10631,N_8323,N_7828);
nand U10632 (N_10632,N_7805,N_8806);
nand U10633 (N_10633,N_7183,N_8129);
nand U10634 (N_10634,N_6816,N_6049);
or U10635 (N_10635,N_8556,N_6410);
or U10636 (N_10636,N_7853,N_7051);
or U10637 (N_10637,N_7787,N_8867);
nor U10638 (N_10638,N_8526,N_8801);
or U10639 (N_10639,N_8955,N_6312);
nand U10640 (N_10640,N_8841,N_7675);
and U10641 (N_10641,N_8097,N_8973);
or U10642 (N_10642,N_6861,N_6308);
nand U10643 (N_10643,N_7616,N_6241);
nand U10644 (N_10644,N_6177,N_8441);
nand U10645 (N_10645,N_7087,N_8874);
nor U10646 (N_10646,N_6645,N_8163);
nand U10647 (N_10647,N_6270,N_6714);
nand U10648 (N_10648,N_8673,N_6603);
or U10649 (N_10649,N_6565,N_7799);
and U10650 (N_10650,N_7737,N_7648);
or U10651 (N_10651,N_6582,N_7158);
nand U10652 (N_10652,N_7844,N_8914);
and U10653 (N_10653,N_8433,N_6820);
nor U10654 (N_10654,N_8939,N_8842);
and U10655 (N_10655,N_7460,N_7670);
or U10656 (N_10656,N_6605,N_8651);
nand U10657 (N_10657,N_8580,N_8482);
and U10658 (N_10658,N_6498,N_7816);
nand U10659 (N_10659,N_7649,N_6311);
and U10660 (N_10660,N_8704,N_8508);
nor U10661 (N_10661,N_6768,N_6459);
nor U10662 (N_10662,N_8200,N_6373);
nor U10663 (N_10663,N_7050,N_7351);
nand U10664 (N_10664,N_7219,N_6198);
nor U10665 (N_10665,N_6819,N_6318);
or U10666 (N_10666,N_6593,N_6981);
nor U10667 (N_10667,N_7965,N_6084);
nor U10668 (N_10668,N_7625,N_8930);
nand U10669 (N_10669,N_8785,N_7296);
or U10670 (N_10670,N_6217,N_7779);
and U10671 (N_10671,N_7089,N_7003);
and U10672 (N_10672,N_7928,N_8387);
and U10673 (N_10673,N_8394,N_7954);
and U10674 (N_10674,N_7372,N_8289);
or U10675 (N_10675,N_6558,N_7454);
nor U10676 (N_10676,N_8661,N_8304);
nand U10677 (N_10677,N_6343,N_6101);
and U10678 (N_10678,N_6200,N_6090);
nand U10679 (N_10679,N_8243,N_8005);
nor U10680 (N_10680,N_6699,N_6910);
nor U10681 (N_10681,N_6359,N_7494);
or U10682 (N_10682,N_8578,N_6254);
or U10683 (N_10683,N_8163,N_6479);
nand U10684 (N_10684,N_6718,N_8516);
nand U10685 (N_10685,N_7781,N_8308);
and U10686 (N_10686,N_6888,N_6942);
or U10687 (N_10687,N_7444,N_6633);
nand U10688 (N_10688,N_8471,N_7138);
nor U10689 (N_10689,N_7195,N_6312);
and U10690 (N_10690,N_8861,N_8573);
or U10691 (N_10691,N_7780,N_7842);
and U10692 (N_10692,N_6224,N_6512);
nand U10693 (N_10693,N_6576,N_7041);
and U10694 (N_10694,N_7636,N_6133);
or U10695 (N_10695,N_8124,N_6155);
or U10696 (N_10696,N_7894,N_7673);
nor U10697 (N_10697,N_6227,N_7286);
nor U10698 (N_10698,N_8149,N_7436);
nand U10699 (N_10699,N_6569,N_6680);
nand U10700 (N_10700,N_8516,N_8894);
or U10701 (N_10701,N_6749,N_8627);
or U10702 (N_10702,N_7156,N_6414);
nand U10703 (N_10703,N_6610,N_7048);
nor U10704 (N_10704,N_6134,N_6950);
and U10705 (N_10705,N_6882,N_7346);
nor U10706 (N_10706,N_6083,N_7324);
nor U10707 (N_10707,N_7440,N_8046);
or U10708 (N_10708,N_8819,N_7879);
or U10709 (N_10709,N_8220,N_6736);
and U10710 (N_10710,N_8549,N_6486);
and U10711 (N_10711,N_7396,N_7312);
and U10712 (N_10712,N_7320,N_7708);
nor U10713 (N_10713,N_8637,N_6416);
nor U10714 (N_10714,N_7017,N_8035);
and U10715 (N_10715,N_7543,N_7333);
nand U10716 (N_10716,N_8285,N_8476);
nor U10717 (N_10717,N_6798,N_8665);
and U10718 (N_10718,N_8581,N_7578);
nand U10719 (N_10719,N_8829,N_8143);
and U10720 (N_10720,N_6627,N_6643);
nor U10721 (N_10721,N_7824,N_6501);
and U10722 (N_10722,N_7313,N_6020);
nor U10723 (N_10723,N_6924,N_6606);
and U10724 (N_10724,N_8695,N_7288);
nand U10725 (N_10725,N_8255,N_7594);
or U10726 (N_10726,N_7639,N_8248);
nor U10727 (N_10727,N_7703,N_6669);
nand U10728 (N_10728,N_8091,N_7156);
nand U10729 (N_10729,N_7861,N_8296);
and U10730 (N_10730,N_8495,N_6121);
nor U10731 (N_10731,N_8938,N_6111);
nand U10732 (N_10732,N_7408,N_7357);
or U10733 (N_10733,N_7898,N_6347);
nand U10734 (N_10734,N_6537,N_7909);
and U10735 (N_10735,N_7683,N_6428);
and U10736 (N_10736,N_8169,N_6078);
nand U10737 (N_10737,N_6103,N_7319);
or U10738 (N_10738,N_6631,N_7094);
or U10739 (N_10739,N_8172,N_6093);
nor U10740 (N_10740,N_6494,N_8356);
nor U10741 (N_10741,N_7602,N_7911);
or U10742 (N_10742,N_7225,N_7316);
or U10743 (N_10743,N_7409,N_6287);
nand U10744 (N_10744,N_7142,N_6562);
and U10745 (N_10745,N_6561,N_8424);
nor U10746 (N_10746,N_8731,N_8496);
or U10747 (N_10747,N_6163,N_6504);
nand U10748 (N_10748,N_8175,N_6787);
or U10749 (N_10749,N_6713,N_8307);
nor U10750 (N_10750,N_8882,N_7451);
and U10751 (N_10751,N_7966,N_7928);
nand U10752 (N_10752,N_7722,N_7344);
or U10753 (N_10753,N_6591,N_6098);
and U10754 (N_10754,N_7140,N_7731);
or U10755 (N_10755,N_6343,N_6829);
or U10756 (N_10756,N_8004,N_7281);
or U10757 (N_10757,N_7960,N_8962);
and U10758 (N_10758,N_7057,N_7214);
nand U10759 (N_10759,N_6849,N_7640);
or U10760 (N_10760,N_8572,N_8381);
or U10761 (N_10761,N_6772,N_7725);
nor U10762 (N_10762,N_6727,N_6711);
nand U10763 (N_10763,N_8276,N_6672);
nand U10764 (N_10764,N_7942,N_8415);
and U10765 (N_10765,N_6266,N_6372);
nand U10766 (N_10766,N_7400,N_7620);
and U10767 (N_10767,N_8591,N_8633);
nand U10768 (N_10768,N_7926,N_6565);
nand U10769 (N_10769,N_7014,N_8076);
or U10770 (N_10770,N_7762,N_8722);
nand U10771 (N_10771,N_6618,N_6312);
and U10772 (N_10772,N_6567,N_7901);
and U10773 (N_10773,N_6064,N_8349);
or U10774 (N_10774,N_6998,N_6244);
and U10775 (N_10775,N_6506,N_6530);
nor U10776 (N_10776,N_6413,N_7164);
nor U10777 (N_10777,N_6812,N_7331);
or U10778 (N_10778,N_7118,N_7638);
or U10779 (N_10779,N_8384,N_7574);
nor U10780 (N_10780,N_8856,N_7126);
or U10781 (N_10781,N_8819,N_8132);
and U10782 (N_10782,N_6124,N_8606);
nand U10783 (N_10783,N_6832,N_8757);
and U10784 (N_10784,N_6138,N_6924);
or U10785 (N_10785,N_6386,N_7225);
nor U10786 (N_10786,N_6627,N_8065);
and U10787 (N_10787,N_6501,N_7284);
nand U10788 (N_10788,N_8771,N_7436);
and U10789 (N_10789,N_6702,N_6879);
or U10790 (N_10790,N_7790,N_7804);
and U10791 (N_10791,N_8676,N_8326);
nand U10792 (N_10792,N_7608,N_8986);
nand U10793 (N_10793,N_7748,N_8898);
and U10794 (N_10794,N_6603,N_8293);
nand U10795 (N_10795,N_6570,N_8480);
nor U10796 (N_10796,N_7634,N_8414);
and U10797 (N_10797,N_8497,N_8901);
nor U10798 (N_10798,N_6941,N_8504);
nand U10799 (N_10799,N_7158,N_8236);
and U10800 (N_10800,N_7109,N_6430);
xor U10801 (N_10801,N_8824,N_8939);
and U10802 (N_10802,N_6479,N_7098);
and U10803 (N_10803,N_6781,N_8022);
nor U10804 (N_10804,N_8369,N_7168);
and U10805 (N_10805,N_8640,N_6276);
or U10806 (N_10806,N_6293,N_7294);
and U10807 (N_10807,N_7077,N_7257);
or U10808 (N_10808,N_8752,N_7512);
and U10809 (N_10809,N_6936,N_8376);
or U10810 (N_10810,N_7143,N_7489);
or U10811 (N_10811,N_8486,N_7764);
nor U10812 (N_10812,N_7776,N_7107);
or U10813 (N_10813,N_7621,N_7856);
or U10814 (N_10814,N_8606,N_8422);
nand U10815 (N_10815,N_8528,N_6653);
and U10816 (N_10816,N_6385,N_7298);
and U10817 (N_10817,N_7014,N_8415);
nor U10818 (N_10818,N_7479,N_7442);
and U10819 (N_10819,N_7256,N_7131);
nand U10820 (N_10820,N_6711,N_8621);
or U10821 (N_10821,N_7819,N_8908);
nand U10822 (N_10822,N_7569,N_7324);
or U10823 (N_10823,N_6023,N_8455);
nand U10824 (N_10824,N_6177,N_7869);
nor U10825 (N_10825,N_7103,N_6696);
and U10826 (N_10826,N_6486,N_7884);
and U10827 (N_10827,N_7098,N_8945);
or U10828 (N_10828,N_6289,N_7994);
and U10829 (N_10829,N_8551,N_8349);
and U10830 (N_10830,N_7759,N_6109);
and U10831 (N_10831,N_7441,N_7104);
or U10832 (N_10832,N_6708,N_6811);
nand U10833 (N_10833,N_6850,N_6454);
or U10834 (N_10834,N_7297,N_8329);
nor U10835 (N_10835,N_7290,N_8905);
nor U10836 (N_10836,N_8553,N_8831);
and U10837 (N_10837,N_7323,N_7025);
nand U10838 (N_10838,N_6134,N_8715);
or U10839 (N_10839,N_7048,N_7249);
nor U10840 (N_10840,N_6214,N_8747);
nand U10841 (N_10841,N_7351,N_7053);
or U10842 (N_10842,N_8913,N_6981);
or U10843 (N_10843,N_6183,N_6242);
and U10844 (N_10844,N_7894,N_8410);
nand U10845 (N_10845,N_7059,N_8529);
nand U10846 (N_10846,N_8161,N_7199);
or U10847 (N_10847,N_6702,N_7120);
nor U10848 (N_10848,N_7258,N_7688);
or U10849 (N_10849,N_7429,N_7001);
nand U10850 (N_10850,N_8908,N_6049);
or U10851 (N_10851,N_8565,N_7695);
nor U10852 (N_10852,N_6859,N_6661);
nand U10853 (N_10853,N_8777,N_7291);
nand U10854 (N_10854,N_6819,N_7789);
nor U10855 (N_10855,N_8173,N_7763);
xnor U10856 (N_10856,N_8831,N_6723);
nor U10857 (N_10857,N_6206,N_7052);
and U10858 (N_10858,N_6170,N_8074);
and U10859 (N_10859,N_8495,N_6076);
or U10860 (N_10860,N_7518,N_6081);
nor U10861 (N_10861,N_6106,N_8995);
and U10862 (N_10862,N_8705,N_6943);
or U10863 (N_10863,N_7299,N_7750);
and U10864 (N_10864,N_7239,N_7355);
or U10865 (N_10865,N_8373,N_7412);
and U10866 (N_10866,N_8654,N_7196);
or U10867 (N_10867,N_7533,N_6932);
nor U10868 (N_10868,N_6385,N_6931);
or U10869 (N_10869,N_6044,N_6430);
or U10870 (N_10870,N_6702,N_7531);
nor U10871 (N_10871,N_8414,N_6191);
nor U10872 (N_10872,N_8482,N_7475);
or U10873 (N_10873,N_7664,N_6451);
or U10874 (N_10874,N_8805,N_7130);
nor U10875 (N_10875,N_6992,N_8269);
or U10876 (N_10876,N_6152,N_7644);
or U10877 (N_10877,N_6920,N_6273);
xnor U10878 (N_10878,N_8231,N_7323);
or U10879 (N_10879,N_6575,N_8866);
nand U10880 (N_10880,N_8485,N_6947);
or U10881 (N_10881,N_8059,N_7893);
or U10882 (N_10882,N_6362,N_6942);
nand U10883 (N_10883,N_8584,N_6527);
xnor U10884 (N_10884,N_8890,N_7360);
nor U10885 (N_10885,N_6815,N_6991);
and U10886 (N_10886,N_7584,N_8535);
or U10887 (N_10887,N_8311,N_6031);
or U10888 (N_10888,N_6315,N_7041);
xnor U10889 (N_10889,N_6774,N_6581);
and U10890 (N_10890,N_7078,N_6065);
nand U10891 (N_10891,N_8626,N_8768);
or U10892 (N_10892,N_8064,N_6281);
or U10893 (N_10893,N_7368,N_6602);
nand U10894 (N_10894,N_8717,N_8125);
nor U10895 (N_10895,N_6426,N_7176);
nand U10896 (N_10896,N_8309,N_8474);
and U10897 (N_10897,N_6942,N_7815);
nand U10898 (N_10898,N_6815,N_8260);
nand U10899 (N_10899,N_8767,N_7332);
nor U10900 (N_10900,N_6188,N_8277);
or U10901 (N_10901,N_8219,N_6943);
nand U10902 (N_10902,N_8043,N_7057);
nand U10903 (N_10903,N_7137,N_6361);
or U10904 (N_10904,N_7528,N_8842);
nor U10905 (N_10905,N_8393,N_7397);
nand U10906 (N_10906,N_7384,N_8311);
and U10907 (N_10907,N_7830,N_7122);
nor U10908 (N_10908,N_6397,N_7240);
or U10909 (N_10909,N_8254,N_7168);
nand U10910 (N_10910,N_6017,N_8378);
nand U10911 (N_10911,N_7931,N_7287);
or U10912 (N_10912,N_8877,N_8722);
nor U10913 (N_10913,N_7151,N_8764);
and U10914 (N_10914,N_7436,N_7506);
or U10915 (N_10915,N_7081,N_8473);
and U10916 (N_10916,N_7243,N_8695);
and U10917 (N_10917,N_6056,N_6576);
and U10918 (N_10918,N_8420,N_7793);
nor U10919 (N_10919,N_6069,N_7356);
and U10920 (N_10920,N_7062,N_6315);
nand U10921 (N_10921,N_6243,N_8079);
and U10922 (N_10922,N_7549,N_8037);
or U10923 (N_10923,N_8259,N_7761);
nand U10924 (N_10924,N_6889,N_6197);
nor U10925 (N_10925,N_6550,N_8217);
nor U10926 (N_10926,N_7748,N_7970);
nor U10927 (N_10927,N_7066,N_8832);
nor U10928 (N_10928,N_7276,N_6130);
nor U10929 (N_10929,N_6832,N_6882);
and U10930 (N_10930,N_8317,N_6685);
and U10931 (N_10931,N_8621,N_8238);
nand U10932 (N_10932,N_6154,N_6784);
and U10933 (N_10933,N_7257,N_7391);
or U10934 (N_10934,N_7630,N_7071);
nand U10935 (N_10935,N_6244,N_7454);
and U10936 (N_10936,N_8567,N_6284);
nor U10937 (N_10937,N_6309,N_7011);
and U10938 (N_10938,N_8888,N_8939);
nor U10939 (N_10939,N_8063,N_7159);
and U10940 (N_10940,N_7127,N_6199);
or U10941 (N_10941,N_8635,N_8676);
nor U10942 (N_10942,N_7913,N_6047);
nor U10943 (N_10943,N_7373,N_7110);
or U10944 (N_10944,N_7898,N_6427);
or U10945 (N_10945,N_7853,N_6918);
and U10946 (N_10946,N_6523,N_7211);
nand U10947 (N_10947,N_8456,N_8273);
nand U10948 (N_10948,N_8798,N_8502);
nand U10949 (N_10949,N_6104,N_8196);
nor U10950 (N_10950,N_7752,N_6925);
and U10951 (N_10951,N_8555,N_8653);
or U10952 (N_10952,N_8627,N_6789);
and U10953 (N_10953,N_8367,N_7186);
or U10954 (N_10954,N_7581,N_7630);
or U10955 (N_10955,N_7216,N_6703);
nand U10956 (N_10956,N_7670,N_8658);
nand U10957 (N_10957,N_6427,N_7100);
or U10958 (N_10958,N_8159,N_6206);
nand U10959 (N_10959,N_6760,N_6840);
and U10960 (N_10960,N_6715,N_7986);
or U10961 (N_10961,N_7709,N_7734);
or U10962 (N_10962,N_7946,N_7956);
and U10963 (N_10963,N_7365,N_8437);
or U10964 (N_10964,N_6871,N_8768);
nor U10965 (N_10965,N_7102,N_7938);
or U10966 (N_10966,N_7922,N_6360);
nand U10967 (N_10967,N_7687,N_8176);
or U10968 (N_10968,N_8725,N_8468);
and U10969 (N_10969,N_8384,N_8338);
or U10970 (N_10970,N_8883,N_7351);
nand U10971 (N_10971,N_7576,N_7173);
nand U10972 (N_10972,N_8934,N_6718);
nor U10973 (N_10973,N_8978,N_8440);
and U10974 (N_10974,N_6193,N_7778);
and U10975 (N_10975,N_7397,N_7059);
nand U10976 (N_10976,N_8698,N_7930);
or U10977 (N_10977,N_6740,N_7234);
or U10978 (N_10978,N_6762,N_6305);
nand U10979 (N_10979,N_7320,N_7350);
and U10980 (N_10980,N_8176,N_6125);
nand U10981 (N_10981,N_8368,N_7609);
and U10982 (N_10982,N_8041,N_6695);
nand U10983 (N_10983,N_6948,N_8476);
and U10984 (N_10984,N_8830,N_7316);
and U10985 (N_10985,N_6389,N_6977);
nand U10986 (N_10986,N_6318,N_6272);
nor U10987 (N_10987,N_8796,N_8749);
nor U10988 (N_10988,N_8618,N_6791);
and U10989 (N_10989,N_8684,N_8085);
or U10990 (N_10990,N_7557,N_8972);
nor U10991 (N_10991,N_8964,N_7028);
or U10992 (N_10992,N_7091,N_7583);
nand U10993 (N_10993,N_7764,N_7364);
nand U10994 (N_10994,N_6326,N_8457);
nor U10995 (N_10995,N_6058,N_7829);
and U10996 (N_10996,N_6246,N_8525);
and U10997 (N_10997,N_6446,N_7324);
or U10998 (N_10998,N_7156,N_8748);
nand U10999 (N_10999,N_8650,N_6710);
nand U11000 (N_11000,N_7241,N_7070);
nor U11001 (N_11001,N_7136,N_8501);
nand U11002 (N_11002,N_7801,N_8269);
nand U11003 (N_11003,N_6733,N_6482);
or U11004 (N_11004,N_7137,N_8276);
and U11005 (N_11005,N_7055,N_8828);
or U11006 (N_11006,N_8152,N_8606);
nand U11007 (N_11007,N_8545,N_7097);
nor U11008 (N_11008,N_8188,N_6818);
and U11009 (N_11009,N_8079,N_6577);
nor U11010 (N_11010,N_7742,N_6509);
or U11011 (N_11011,N_6353,N_7206);
and U11012 (N_11012,N_7084,N_8909);
nand U11013 (N_11013,N_6301,N_6626);
or U11014 (N_11014,N_7323,N_8686);
or U11015 (N_11015,N_6903,N_6924);
nand U11016 (N_11016,N_6950,N_8972);
nand U11017 (N_11017,N_8422,N_7126);
or U11018 (N_11018,N_6335,N_7902);
xor U11019 (N_11019,N_7561,N_6605);
nand U11020 (N_11020,N_7394,N_7221);
or U11021 (N_11021,N_7292,N_8649);
and U11022 (N_11022,N_8434,N_7621);
and U11023 (N_11023,N_6874,N_7393);
and U11024 (N_11024,N_8705,N_7179);
nand U11025 (N_11025,N_6567,N_8142);
nor U11026 (N_11026,N_6709,N_7348);
and U11027 (N_11027,N_8985,N_7283);
nand U11028 (N_11028,N_7184,N_6945);
nand U11029 (N_11029,N_7980,N_6657);
nand U11030 (N_11030,N_6466,N_6800);
and U11031 (N_11031,N_8664,N_6442);
and U11032 (N_11032,N_6506,N_7505);
and U11033 (N_11033,N_8667,N_7548);
nor U11034 (N_11034,N_8907,N_7362);
nand U11035 (N_11035,N_8277,N_8074);
nor U11036 (N_11036,N_7516,N_7938);
nand U11037 (N_11037,N_7007,N_8730);
and U11038 (N_11038,N_8555,N_6186);
or U11039 (N_11039,N_7523,N_8803);
and U11040 (N_11040,N_7941,N_7030);
or U11041 (N_11041,N_7327,N_7005);
nand U11042 (N_11042,N_7983,N_8277);
nor U11043 (N_11043,N_6490,N_8036);
and U11044 (N_11044,N_6861,N_7193);
nand U11045 (N_11045,N_7316,N_7329);
or U11046 (N_11046,N_8687,N_6722);
or U11047 (N_11047,N_6262,N_8417);
or U11048 (N_11048,N_6993,N_7668);
or U11049 (N_11049,N_8876,N_7457);
and U11050 (N_11050,N_7280,N_6644);
and U11051 (N_11051,N_8319,N_6745);
nand U11052 (N_11052,N_6070,N_7818);
and U11053 (N_11053,N_6764,N_6201);
or U11054 (N_11054,N_8881,N_6175);
or U11055 (N_11055,N_8812,N_8382);
or U11056 (N_11056,N_7256,N_6050);
and U11057 (N_11057,N_7655,N_8415);
and U11058 (N_11058,N_6363,N_7673);
and U11059 (N_11059,N_7052,N_7307);
nand U11060 (N_11060,N_6661,N_6081);
nand U11061 (N_11061,N_6915,N_8262);
or U11062 (N_11062,N_6038,N_7265);
or U11063 (N_11063,N_8845,N_7294);
nor U11064 (N_11064,N_8471,N_6660);
or U11065 (N_11065,N_6061,N_8752);
nor U11066 (N_11066,N_6484,N_8547);
nor U11067 (N_11067,N_7991,N_7208);
or U11068 (N_11068,N_8443,N_7879);
and U11069 (N_11069,N_8207,N_7890);
or U11070 (N_11070,N_8634,N_8016);
nand U11071 (N_11071,N_8811,N_6866);
nor U11072 (N_11072,N_8039,N_7365);
and U11073 (N_11073,N_6262,N_6845);
or U11074 (N_11074,N_7308,N_7253);
or U11075 (N_11075,N_6406,N_8622);
nand U11076 (N_11076,N_7804,N_8202);
and U11077 (N_11077,N_6698,N_6432);
and U11078 (N_11078,N_6461,N_8861);
and U11079 (N_11079,N_8541,N_8906);
and U11080 (N_11080,N_7518,N_7877);
nand U11081 (N_11081,N_6307,N_6303);
nor U11082 (N_11082,N_6679,N_8432);
or U11083 (N_11083,N_6493,N_7138);
and U11084 (N_11084,N_7603,N_8276);
nand U11085 (N_11085,N_7442,N_7853);
nand U11086 (N_11086,N_7572,N_8375);
nand U11087 (N_11087,N_8303,N_7662);
nand U11088 (N_11088,N_6893,N_6116);
and U11089 (N_11089,N_6201,N_6684);
or U11090 (N_11090,N_7066,N_7683);
or U11091 (N_11091,N_8025,N_8929);
and U11092 (N_11092,N_6430,N_8617);
and U11093 (N_11093,N_7540,N_7971);
nand U11094 (N_11094,N_8158,N_6232);
nand U11095 (N_11095,N_7857,N_7656);
and U11096 (N_11096,N_6085,N_8126);
nand U11097 (N_11097,N_7253,N_6222);
and U11098 (N_11098,N_7495,N_7156);
nor U11099 (N_11099,N_8268,N_6182);
or U11100 (N_11100,N_8165,N_8535);
nand U11101 (N_11101,N_7849,N_8927);
nand U11102 (N_11102,N_8985,N_8547);
or U11103 (N_11103,N_8458,N_8961);
nor U11104 (N_11104,N_8112,N_8437);
or U11105 (N_11105,N_7253,N_6522);
nand U11106 (N_11106,N_7124,N_6964);
nand U11107 (N_11107,N_8624,N_6923);
or U11108 (N_11108,N_7663,N_8016);
and U11109 (N_11109,N_8396,N_8656);
nand U11110 (N_11110,N_8236,N_8501);
and U11111 (N_11111,N_7323,N_6654);
or U11112 (N_11112,N_8285,N_7585);
and U11113 (N_11113,N_7292,N_7718);
and U11114 (N_11114,N_7526,N_7168);
nand U11115 (N_11115,N_8196,N_6280);
and U11116 (N_11116,N_6515,N_7312);
and U11117 (N_11117,N_8873,N_8162);
or U11118 (N_11118,N_7907,N_6338);
or U11119 (N_11119,N_8027,N_8668);
or U11120 (N_11120,N_7986,N_7531);
nand U11121 (N_11121,N_6425,N_6030);
nor U11122 (N_11122,N_7257,N_8918);
nor U11123 (N_11123,N_7914,N_6999);
nor U11124 (N_11124,N_6148,N_6779);
nand U11125 (N_11125,N_8325,N_8858);
or U11126 (N_11126,N_6077,N_7294);
and U11127 (N_11127,N_8708,N_6288);
or U11128 (N_11128,N_6622,N_6225);
and U11129 (N_11129,N_6290,N_6859);
and U11130 (N_11130,N_6804,N_8370);
and U11131 (N_11131,N_8926,N_8237);
nand U11132 (N_11132,N_7545,N_7587);
or U11133 (N_11133,N_8152,N_8755);
nand U11134 (N_11134,N_8813,N_8748);
or U11135 (N_11135,N_7158,N_7607);
nand U11136 (N_11136,N_8219,N_7530);
or U11137 (N_11137,N_7233,N_6437);
nand U11138 (N_11138,N_6429,N_6789);
nor U11139 (N_11139,N_8977,N_8199);
or U11140 (N_11140,N_7650,N_8460);
or U11141 (N_11141,N_8917,N_8885);
nand U11142 (N_11142,N_8919,N_7056);
or U11143 (N_11143,N_8668,N_8924);
and U11144 (N_11144,N_6422,N_8488);
or U11145 (N_11145,N_6406,N_7716);
or U11146 (N_11146,N_6312,N_6481);
or U11147 (N_11147,N_7641,N_7024);
nor U11148 (N_11148,N_7902,N_6553);
and U11149 (N_11149,N_7696,N_8732);
nor U11150 (N_11150,N_7499,N_7008);
nand U11151 (N_11151,N_6242,N_8262);
nand U11152 (N_11152,N_6835,N_8122);
and U11153 (N_11153,N_7715,N_7770);
and U11154 (N_11154,N_8220,N_8617);
nand U11155 (N_11155,N_6468,N_6990);
nand U11156 (N_11156,N_6264,N_7427);
or U11157 (N_11157,N_7836,N_7095);
nand U11158 (N_11158,N_7108,N_7342);
and U11159 (N_11159,N_7527,N_6677);
and U11160 (N_11160,N_7037,N_7397);
nor U11161 (N_11161,N_6470,N_7199);
and U11162 (N_11162,N_8556,N_7827);
or U11163 (N_11163,N_8133,N_8488);
nand U11164 (N_11164,N_6102,N_6486);
nor U11165 (N_11165,N_7978,N_8158);
nor U11166 (N_11166,N_6425,N_8019);
nand U11167 (N_11167,N_8238,N_6066);
and U11168 (N_11168,N_7836,N_7433);
or U11169 (N_11169,N_8540,N_6555);
and U11170 (N_11170,N_7720,N_8153);
or U11171 (N_11171,N_6910,N_7086);
and U11172 (N_11172,N_7069,N_7148);
nor U11173 (N_11173,N_7022,N_6857);
or U11174 (N_11174,N_7319,N_6258);
nor U11175 (N_11175,N_8705,N_8039);
nand U11176 (N_11176,N_6662,N_7049);
nor U11177 (N_11177,N_6715,N_8853);
nand U11178 (N_11178,N_6699,N_8499);
or U11179 (N_11179,N_8557,N_6128);
nand U11180 (N_11180,N_8527,N_7810);
and U11181 (N_11181,N_6916,N_7410);
or U11182 (N_11182,N_7146,N_8182);
nor U11183 (N_11183,N_6699,N_6956);
nor U11184 (N_11184,N_7626,N_7336);
and U11185 (N_11185,N_8974,N_8873);
or U11186 (N_11186,N_8141,N_8348);
nor U11187 (N_11187,N_8855,N_6152);
and U11188 (N_11188,N_6328,N_7959);
nand U11189 (N_11189,N_7802,N_7662);
or U11190 (N_11190,N_7248,N_6681);
nand U11191 (N_11191,N_6697,N_7729);
or U11192 (N_11192,N_7874,N_8537);
and U11193 (N_11193,N_7495,N_6194);
nand U11194 (N_11194,N_8812,N_7321);
nor U11195 (N_11195,N_6193,N_7436);
and U11196 (N_11196,N_7896,N_7238);
nor U11197 (N_11197,N_8824,N_6517);
or U11198 (N_11198,N_7022,N_6771);
nand U11199 (N_11199,N_8283,N_7977);
nand U11200 (N_11200,N_7027,N_7368);
nand U11201 (N_11201,N_6363,N_7106);
nor U11202 (N_11202,N_6705,N_6775);
and U11203 (N_11203,N_6951,N_8608);
or U11204 (N_11204,N_6318,N_6844);
nor U11205 (N_11205,N_6613,N_6020);
and U11206 (N_11206,N_8076,N_8736);
and U11207 (N_11207,N_8372,N_8871);
nand U11208 (N_11208,N_8278,N_8417);
nand U11209 (N_11209,N_8223,N_7417);
and U11210 (N_11210,N_8720,N_8609);
and U11211 (N_11211,N_8794,N_6422);
or U11212 (N_11212,N_7104,N_6041);
or U11213 (N_11213,N_7362,N_6578);
and U11214 (N_11214,N_6045,N_6281);
nor U11215 (N_11215,N_6492,N_7015);
nand U11216 (N_11216,N_8153,N_8185);
nand U11217 (N_11217,N_6252,N_8262);
nand U11218 (N_11218,N_6699,N_8089);
nand U11219 (N_11219,N_8238,N_7614);
nor U11220 (N_11220,N_6403,N_7180);
and U11221 (N_11221,N_7108,N_7522);
and U11222 (N_11222,N_6744,N_6705);
and U11223 (N_11223,N_6193,N_7772);
nor U11224 (N_11224,N_6670,N_8219);
or U11225 (N_11225,N_7585,N_8250);
or U11226 (N_11226,N_8378,N_8375);
or U11227 (N_11227,N_6658,N_7233);
nor U11228 (N_11228,N_7820,N_8075);
or U11229 (N_11229,N_6488,N_8276);
and U11230 (N_11230,N_8762,N_6978);
nor U11231 (N_11231,N_6785,N_7827);
and U11232 (N_11232,N_8445,N_7834);
and U11233 (N_11233,N_8423,N_7765);
and U11234 (N_11234,N_8932,N_8749);
nand U11235 (N_11235,N_7168,N_6955);
nor U11236 (N_11236,N_8233,N_8190);
nor U11237 (N_11237,N_8360,N_6757);
or U11238 (N_11238,N_8323,N_8390);
and U11239 (N_11239,N_7343,N_6001);
or U11240 (N_11240,N_7039,N_6842);
and U11241 (N_11241,N_6245,N_7542);
and U11242 (N_11242,N_8438,N_6941);
or U11243 (N_11243,N_7478,N_7570);
or U11244 (N_11244,N_8470,N_7783);
and U11245 (N_11245,N_6358,N_8382);
or U11246 (N_11246,N_8069,N_6364);
and U11247 (N_11247,N_8317,N_6169);
and U11248 (N_11248,N_7794,N_6809);
and U11249 (N_11249,N_8842,N_7569);
nand U11250 (N_11250,N_8408,N_6385);
nor U11251 (N_11251,N_6899,N_6606);
or U11252 (N_11252,N_7490,N_6855);
and U11253 (N_11253,N_7354,N_6816);
nor U11254 (N_11254,N_7093,N_7863);
and U11255 (N_11255,N_8136,N_8637);
nor U11256 (N_11256,N_6510,N_6377);
nand U11257 (N_11257,N_7378,N_7718);
nor U11258 (N_11258,N_7778,N_6831);
or U11259 (N_11259,N_7973,N_8212);
nand U11260 (N_11260,N_8683,N_8918);
nand U11261 (N_11261,N_7533,N_8178);
and U11262 (N_11262,N_8438,N_6181);
nor U11263 (N_11263,N_7534,N_7471);
or U11264 (N_11264,N_8004,N_8818);
and U11265 (N_11265,N_7596,N_8136);
xnor U11266 (N_11266,N_7659,N_6869);
and U11267 (N_11267,N_7581,N_8318);
nor U11268 (N_11268,N_6739,N_6569);
nor U11269 (N_11269,N_7025,N_7419);
and U11270 (N_11270,N_6176,N_7373);
nor U11271 (N_11271,N_6291,N_8296);
nor U11272 (N_11272,N_7895,N_8822);
or U11273 (N_11273,N_8146,N_6814);
or U11274 (N_11274,N_6329,N_8892);
or U11275 (N_11275,N_8487,N_6004);
nor U11276 (N_11276,N_7131,N_7139);
nand U11277 (N_11277,N_7854,N_8105);
nand U11278 (N_11278,N_6616,N_7436);
nand U11279 (N_11279,N_6690,N_6156);
nand U11280 (N_11280,N_8525,N_8708);
nand U11281 (N_11281,N_8332,N_8056);
or U11282 (N_11282,N_7136,N_7509);
and U11283 (N_11283,N_8362,N_6668);
nor U11284 (N_11284,N_6658,N_6036);
nor U11285 (N_11285,N_6581,N_8265);
nor U11286 (N_11286,N_8575,N_7478);
nand U11287 (N_11287,N_6948,N_8880);
or U11288 (N_11288,N_7950,N_8701);
and U11289 (N_11289,N_8871,N_7841);
nand U11290 (N_11290,N_7482,N_6891);
and U11291 (N_11291,N_7070,N_7628);
nor U11292 (N_11292,N_7876,N_7743);
or U11293 (N_11293,N_7538,N_8042);
nor U11294 (N_11294,N_8153,N_7981);
or U11295 (N_11295,N_8346,N_8378);
nor U11296 (N_11296,N_6908,N_7168);
or U11297 (N_11297,N_7973,N_6683);
nor U11298 (N_11298,N_7044,N_6972);
nand U11299 (N_11299,N_6924,N_8818);
nand U11300 (N_11300,N_8120,N_8113);
and U11301 (N_11301,N_8922,N_8596);
nor U11302 (N_11302,N_8042,N_8344);
or U11303 (N_11303,N_8227,N_7447);
xor U11304 (N_11304,N_6721,N_8646);
and U11305 (N_11305,N_8917,N_7547);
nor U11306 (N_11306,N_6245,N_6968);
or U11307 (N_11307,N_7943,N_7746);
nand U11308 (N_11308,N_8131,N_6188);
and U11309 (N_11309,N_6011,N_8333);
or U11310 (N_11310,N_7127,N_7393);
or U11311 (N_11311,N_6210,N_7731);
and U11312 (N_11312,N_6318,N_7589);
or U11313 (N_11313,N_7727,N_8437);
nor U11314 (N_11314,N_6200,N_6093);
nor U11315 (N_11315,N_6040,N_8889);
nand U11316 (N_11316,N_6642,N_7444);
and U11317 (N_11317,N_7405,N_6613);
and U11318 (N_11318,N_8188,N_6316);
nor U11319 (N_11319,N_7470,N_6201);
xnor U11320 (N_11320,N_8858,N_6993);
nand U11321 (N_11321,N_6756,N_6388);
nand U11322 (N_11322,N_7343,N_8347);
nor U11323 (N_11323,N_6659,N_6505);
nand U11324 (N_11324,N_7667,N_6668);
and U11325 (N_11325,N_7538,N_7365);
nand U11326 (N_11326,N_8855,N_8687);
nand U11327 (N_11327,N_8945,N_7241);
nand U11328 (N_11328,N_7730,N_6632);
or U11329 (N_11329,N_8650,N_8262);
or U11330 (N_11330,N_6620,N_6565);
and U11331 (N_11331,N_7291,N_6156);
nor U11332 (N_11332,N_7364,N_6470);
nand U11333 (N_11333,N_7104,N_7648);
nor U11334 (N_11334,N_8326,N_7207);
nor U11335 (N_11335,N_7975,N_6489);
and U11336 (N_11336,N_6014,N_8004);
nand U11337 (N_11337,N_7235,N_6323);
or U11338 (N_11338,N_8397,N_8464);
or U11339 (N_11339,N_8340,N_8915);
nor U11340 (N_11340,N_7155,N_6131);
and U11341 (N_11341,N_6796,N_8726);
and U11342 (N_11342,N_7683,N_7867);
and U11343 (N_11343,N_8851,N_6434);
nor U11344 (N_11344,N_8429,N_8853);
or U11345 (N_11345,N_7455,N_7941);
nand U11346 (N_11346,N_8659,N_6995);
nor U11347 (N_11347,N_6184,N_8898);
nor U11348 (N_11348,N_7916,N_8386);
and U11349 (N_11349,N_7798,N_8627);
nand U11350 (N_11350,N_8315,N_8964);
and U11351 (N_11351,N_8966,N_7809);
nor U11352 (N_11352,N_8601,N_6071);
or U11353 (N_11353,N_7247,N_7761);
and U11354 (N_11354,N_6556,N_6561);
nand U11355 (N_11355,N_7080,N_8051);
nand U11356 (N_11356,N_8530,N_8570);
nand U11357 (N_11357,N_7865,N_7500);
or U11358 (N_11358,N_6392,N_7854);
and U11359 (N_11359,N_8042,N_6809);
nand U11360 (N_11360,N_7950,N_8764);
nand U11361 (N_11361,N_6558,N_6185);
nor U11362 (N_11362,N_7233,N_6300);
nand U11363 (N_11363,N_6210,N_6040);
nand U11364 (N_11364,N_7547,N_6618);
or U11365 (N_11365,N_8004,N_8383);
nand U11366 (N_11366,N_8581,N_6512);
and U11367 (N_11367,N_8636,N_7627);
nor U11368 (N_11368,N_8690,N_6148);
or U11369 (N_11369,N_8742,N_7209);
nor U11370 (N_11370,N_6940,N_7290);
nor U11371 (N_11371,N_7863,N_6651);
nand U11372 (N_11372,N_7521,N_8314);
nand U11373 (N_11373,N_8798,N_8082);
nor U11374 (N_11374,N_8917,N_6647);
or U11375 (N_11375,N_8367,N_6316);
and U11376 (N_11376,N_7053,N_6734);
or U11377 (N_11377,N_8292,N_6931);
nor U11378 (N_11378,N_6567,N_7541);
nor U11379 (N_11379,N_8653,N_7907);
or U11380 (N_11380,N_8538,N_8613);
nand U11381 (N_11381,N_8539,N_7731);
or U11382 (N_11382,N_7998,N_8892);
xnor U11383 (N_11383,N_7538,N_7446);
nor U11384 (N_11384,N_6060,N_7402);
and U11385 (N_11385,N_8344,N_8245);
nand U11386 (N_11386,N_8545,N_7168);
nand U11387 (N_11387,N_6637,N_6901);
nor U11388 (N_11388,N_8186,N_7353);
nor U11389 (N_11389,N_8045,N_7640);
and U11390 (N_11390,N_6866,N_8893);
nand U11391 (N_11391,N_7683,N_8889);
and U11392 (N_11392,N_7427,N_7115);
nand U11393 (N_11393,N_8417,N_8687);
nor U11394 (N_11394,N_7507,N_7543);
xor U11395 (N_11395,N_7325,N_6127);
and U11396 (N_11396,N_8613,N_6350);
or U11397 (N_11397,N_8375,N_7053);
nor U11398 (N_11398,N_8181,N_8004);
nand U11399 (N_11399,N_8076,N_8805);
nand U11400 (N_11400,N_7205,N_6218);
nor U11401 (N_11401,N_6415,N_8049);
and U11402 (N_11402,N_8824,N_7545);
or U11403 (N_11403,N_7214,N_7710);
nor U11404 (N_11404,N_6961,N_8309);
nor U11405 (N_11405,N_7816,N_8974);
nor U11406 (N_11406,N_7848,N_6173);
and U11407 (N_11407,N_8374,N_7036);
nand U11408 (N_11408,N_8337,N_7603);
nor U11409 (N_11409,N_6101,N_7814);
nor U11410 (N_11410,N_6701,N_8812);
and U11411 (N_11411,N_8165,N_8810);
nor U11412 (N_11412,N_7142,N_8277);
nor U11413 (N_11413,N_6832,N_6872);
nand U11414 (N_11414,N_6778,N_6179);
and U11415 (N_11415,N_7137,N_8963);
nand U11416 (N_11416,N_6876,N_7192);
nor U11417 (N_11417,N_6255,N_8830);
nor U11418 (N_11418,N_8436,N_8326);
and U11419 (N_11419,N_8127,N_7739);
nor U11420 (N_11420,N_7601,N_6440);
nor U11421 (N_11421,N_8145,N_8351);
nand U11422 (N_11422,N_7729,N_7483);
nor U11423 (N_11423,N_6456,N_7079);
nand U11424 (N_11424,N_8442,N_8929);
or U11425 (N_11425,N_6180,N_7010);
and U11426 (N_11426,N_7496,N_6024);
nand U11427 (N_11427,N_6670,N_7680);
nand U11428 (N_11428,N_6607,N_8132);
or U11429 (N_11429,N_8848,N_6884);
nand U11430 (N_11430,N_6866,N_8787);
and U11431 (N_11431,N_8072,N_6719);
and U11432 (N_11432,N_6522,N_6530);
nor U11433 (N_11433,N_8788,N_8293);
and U11434 (N_11434,N_7934,N_8464);
nor U11435 (N_11435,N_6113,N_6311);
or U11436 (N_11436,N_7877,N_6680);
nor U11437 (N_11437,N_8766,N_8427);
nor U11438 (N_11438,N_8911,N_8494);
nor U11439 (N_11439,N_6272,N_7322);
nor U11440 (N_11440,N_8892,N_6664);
or U11441 (N_11441,N_8731,N_6861);
nor U11442 (N_11442,N_6174,N_6832);
or U11443 (N_11443,N_8739,N_7414);
nor U11444 (N_11444,N_7642,N_7413);
nor U11445 (N_11445,N_7269,N_8966);
nand U11446 (N_11446,N_7526,N_7476);
nor U11447 (N_11447,N_7806,N_8056);
or U11448 (N_11448,N_8227,N_8629);
nor U11449 (N_11449,N_6113,N_6339);
or U11450 (N_11450,N_7176,N_6646);
nand U11451 (N_11451,N_8734,N_7342);
nor U11452 (N_11452,N_7664,N_7359);
nand U11453 (N_11453,N_8413,N_8112);
nand U11454 (N_11454,N_7447,N_8599);
or U11455 (N_11455,N_8320,N_7184);
or U11456 (N_11456,N_6725,N_7659);
nor U11457 (N_11457,N_8185,N_7913);
or U11458 (N_11458,N_7834,N_7909);
xor U11459 (N_11459,N_8721,N_8105);
nor U11460 (N_11460,N_6291,N_6743);
nand U11461 (N_11461,N_8635,N_7607);
nand U11462 (N_11462,N_6781,N_7282);
nand U11463 (N_11463,N_6542,N_6092);
and U11464 (N_11464,N_8991,N_8786);
nor U11465 (N_11465,N_8805,N_8246);
nor U11466 (N_11466,N_8226,N_7662);
and U11467 (N_11467,N_6018,N_6587);
nand U11468 (N_11468,N_6370,N_6694);
nor U11469 (N_11469,N_8436,N_6557);
and U11470 (N_11470,N_7418,N_7037);
and U11471 (N_11471,N_6151,N_8232);
and U11472 (N_11472,N_6876,N_7452);
nor U11473 (N_11473,N_6127,N_8640);
or U11474 (N_11474,N_8117,N_6161);
and U11475 (N_11475,N_6484,N_6788);
or U11476 (N_11476,N_8019,N_6968);
nor U11477 (N_11477,N_8472,N_8026);
or U11478 (N_11478,N_6171,N_7774);
nor U11479 (N_11479,N_6947,N_6496);
nor U11480 (N_11480,N_6874,N_8634);
nor U11481 (N_11481,N_7105,N_6892);
and U11482 (N_11482,N_7174,N_8116);
and U11483 (N_11483,N_8321,N_6557);
nand U11484 (N_11484,N_8232,N_6447);
or U11485 (N_11485,N_6306,N_7753);
and U11486 (N_11486,N_6369,N_7825);
nand U11487 (N_11487,N_8146,N_7696);
or U11488 (N_11488,N_6407,N_8155);
or U11489 (N_11489,N_7833,N_6125);
and U11490 (N_11490,N_8928,N_8153);
nor U11491 (N_11491,N_8660,N_6196);
nor U11492 (N_11492,N_6012,N_8843);
nand U11493 (N_11493,N_7052,N_8791);
nor U11494 (N_11494,N_7777,N_6135);
and U11495 (N_11495,N_7647,N_8494);
or U11496 (N_11496,N_8690,N_8766);
nor U11497 (N_11497,N_7220,N_6761);
nand U11498 (N_11498,N_6031,N_6852);
or U11499 (N_11499,N_7724,N_6585);
or U11500 (N_11500,N_7669,N_7116);
xor U11501 (N_11501,N_8189,N_8474);
and U11502 (N_11502,N_8383,N_8151);
or U11503 (N_11503,N_7768,N_7868);
nand U11504 (N_11504,N_7028,N_7663);
nand U11505 (N_11505,N_6882,N_8151);
nor U11506 (N_11506,N_8117,N_7273);
nand U11507 (N_11507,N_7145,N_7490);
and U11508 (N_11508,N_6658,N_8543);
nand U11509 (N_11509,N_8756,N_6201);
nand U11510 (N_11510,N_7976,N_6110);
nand U11511 (N_11511,N_7754,N_7182);
or U11512 (N_11512,N_8123,N_8107);
or U11513 (N_11513,N_6838,N_8861);
nor U11514 (N_11514,N_6602,N_8357);
or U11515 (N_11515,N_6632,N_7048);
or U11516 (N_11516,N_8279,N_8021);
and U11517 (N_11517,N_6058,N_8874);
or U11518 (N_11518,N_7788,N_8644);
nand U11519 (N_11519,N_7163,N_8474);
nand U11520 (N_11520,N_8973,N_8563);
nand U11521 (N_11521,N_6595,N_6714);
or U11522 (N_11522,N_7519,N_6568);
and U11523 (N_11523,N_7545,N_6534);
or U11524 (N_11524,N_8336,N_7174);
and U11525 (N_11525,N_8597,N_7074);
nor U11526 (N_11526,N_6224,N_6149);
nor U11527 (N_11527,N_8769,N_8557);
nand U11528 (N_11528,N_6893,N_8345);
and U11529 (N_11529,N_8435,N_8121);
nand U11530 (N_11530,N_6752,N_7289);
and U11531 (N_11531,N_8420,N_7933);
or U11532 (N_11532,N_6642,N_8821);
or U11533 (N_11533,N_6774,N_6717);
nand U11534 (N_11534,N_6213,N_8906);
nor U11535 (N_11535,N_8607,N_7991);
or U11536 (N_11536,N_6264,N_8919);
or U11537 (N_11537,N_8067,N_7102);
and U11538 (N_11538,N_8032,N_7708);
and U11539 (N_11539,N_8379,N_7162);
or U11540 (N_11540,N_6328,N_8158);
nand U11541 (N_11541,N_6766,N_8733);
or U11542 (N_11542,N_8920,N_8889);
and U11543 (N_11543,N_6717,N_6758);
nor U11544 (N_11544,N_7926,N_6611);
or U11545 (N_11545,N_8239,N_8114);
nor U11546 (N_11546,N_6779,N_7690);
and U11547 (N_11547,N_7354,N_7337);
nand U11548 (N_11548,N_6508,N_6337);
and U11549 (N_11549,N_6049,N_8926);
and U11550 (N_11550,N_8280,N_7584);
or U11551 (N_11551,N_7367,N_7556);
and U11552 (N_11552,N_7574,N_8499);
and U11553 (N_11553,N_8654,N_8060);
and U11554 (N_11554,N_7156,N_6182);
nand U11555 (N_11555,N_7051,N_6948);
or U11556 (N_11556,N_6282,N_8440);
nand U11557 (N_11557,N_7677,N_6184);
nand U11558 (N_11558,N_8596,N_6723);
or U11559 (N_11559,N_6677,N_8458);
or U11560 (N_11560,N_8001,N_7903);
and U11561 (N_11561,N_6123,N_7108);
or U11562 (N_11562,N_8902,N_6539);
nand U11563 (N_11563,N_7830,N_8407);
and U11564 (N_11564,N_8513,N_6393);
and U11565 (N_11565,N_6054,N_8551);
nand U11566 (N_11566,N_7483,N_7692);
nand U11567 (N_11567,N_7083,N_7240);
nor U11568 (N_11568,N_6531,N_6226);
and U11569 (N_11569,N_6835,N_6636);
nor U11570 (N_11570,N_7448,N_8419);
nor U11571 (N_11571,N_8118,N_8384);
nand U11572 (N_11572,N_8038,N_6972);
nand U11573 (N_11573,N_8385,N_8052);
nor U11574 (N_11574,N_8923,N_8285);
nand U11575 (N_11575,N_6335,N_6317);
nor U11576 (N_11576,N_8573,N_8436);
nand U11577 (N_11577,N_7246,N_6559);
and U11578 (N_11578,N_6521,N_6613);
nand U11579 (N_11579,N_8162,N_8449);
nand U11580 (N_11580,N_7884,N_6171);
nor U11581 (N_11581,N_6132,N_8771);
nor U11582 (N_11582,N_7605,N_8455);
nand U11583 (N_11583,N_8043,N_7551);
nor U11584 (N_11584,N_7293,N_8205);
and U11585 (N_11585,N_7990,N_6177);
or U11586 (N_11586,N_7979,N_7901);
and U11587 (N_11587,N_8250,N_7004);
and U11588 (N_11588,N_8640,N_8499);
nand U11589 (N_11589,N_7331,N_7228);
or U11590 (N_11590,N_8122,N_7613);
nor U11591 (N_11591,N_6258,N_6409);
nand U11592 (N_11592,N_7781,N_6558);
and U11593 (N_11593,N_6112,N_7824);
or U11594 (N_11594,N_8881,N_8525);
or U11595 (N_11595,N_7789,N_7194);
nor U11596 (N_11596,N_8619,N_8380);
and U11597 (N_11597,N_8877,N_7790);
nand U11598 (N_11598,N_7830,N_6623);
nor U11599 (N_11599,N_8697,N_8484);
and U11600 (N_11600,N_7828,N_7407);
nand U11601 (N_11601,N_7154,N_8757);
and U11602 (N_11602,N_6820,N_7876);
or U11603 (N_11603,N_8572,N_7592);
or U11604 (N_11604,N_7752,N_7907);
and U11605 (N_11605,N_6185,N_7556);
nand U11606 (N_11606,N_6665,N_6448);
nor U11607 (N_11607,N_7459,N_8231);
nor U11608 (N_11608,N_8580,N_8707);
or U11609 (N_11609,N_6175,N_6122);
nor U11610 (N_11610,N_7605,N_6000);
nand U11611 (N_11611,N_8430,N_8879);
and U11612 (N_11612,N_7311,N_7667);
nor U11613 (N_11613,N_7294,N_8912);
and U11614 (N_11614,N_6412,N_6555);
nand U11615 (N_11615,N_7421,N_8406);
nor U11616 (N_11616,N_7914,N_7384);
nor U11617 (N_11617,N_8998,N_7005);
or U11618 (N_11618,N_6745,N_8904);
nor U11619 (N_11619,N_8679,N_7723);
and U11620 (N_11620,N_8173,N_6818);
and U11621 (N_11621,N_7165,N_8558);
and U11622 (N_11622,N_8879,N_7250);
nor U11623 (N_11623,N_6607,N_8615);
nor U11624 (N_11624,N_8587,N_7765);
and U11625 (N_11625,N_6929,N_7811);
nor U11626 (N_11626,N_7389,N_8457);
and U11627 (N_11627,N_7045,N_6018);
or U11628 (N_11628,N_7878,N_6953);
nand U11629 (N_11629,N_7636,N_7894);
nor U11630 (N_11630,N_8833,N_6013);
and U11631 (N_11631,N_6390,N_6614);
nand U11632 (N_11632,N_6123,N_7447);
and U11633 (N_11633,N_6992,N_7271);
and U11634 (N_11634,N_8586,N_6562);
nor U11635 (N_11635,N_8547,N_6967);
and U11636 (N_11636,N_6602,N_7472);
nor U11637 (N_11637,N_6463,N_6039);
and U11638 (N_11638,N_7988,N_7378);
nor U11639 (N_11639,N_6772,N_6417);
or U11640 (N_11640,N_6327,N_7450);
or U11641 (N_11641,N_6938,N_6476);
and U11642 (N_11642,N_7349,N_8916);
nor U11643 (N_11643,N_6641,N_7563);
or U11644 (N_11644,N_7070,N_6958);
or U11645 (N_11645,N_7533,N_7947);
or U11646 (N_11646,N_7725,N_6330);
nor U11647 (N_11647,N_8630,N_6597);
nor U11648 (N_11648,N_6081,N_8214);
and U11649 (N_11649,N_7774,N_7503);
nor U11650 (N_11650,N_7956,N_6217);
nand U11651 (N_11651,N_6710,N_8973);
nand U11652 (N_11652,N_6692,N_7379);
and U11653 (N_11653,N_7290,N_8233);
or U11654 (N_11654,N_8342,N_8892);
nor U11655 (N_11655,N_6206,N_6327);
nor U11656 (N_11656,N_7492,N_6586);
nor U11657 (N_11657,N_6493,N_7390);
nand U11658 (N_11658,N_8173,N_7926);
or U11659 (N_11659,N_6921,N_7257);
and U11660 (N_11660,N_8444,N_8687);
nor U11661 (N_11661,N_8690,N_6598);
nor U11662 (N_11662,N_8266,N_8451);
and U11663 (N_11663,N_6869,N_6434);
xor U11664 (N_11664,N_8354,N_8738);
or U11665 (N_11665,N_6005,N_7631);
and U11666 (N_11666,N_8863,N_6870);
or U11667 (N_11667,N_8073,N_6826);
nand U11668 (N_11668,N_6601,N_7547);
or U11669 (N_11669,N_8089,N_7316);
nor U11670 (N_11670,N_6498,N_6956);
nand U11671 (N_11671,N_6256,N_8004);
and U11672 (N_11672,N_7917,N_8418);
and U11673 (N_11673,N_7721,N_8029);
or U11674 (N_11674,N_6604,N_8689);
nand U11675 (N_11675,N_8733,N_8947);
nor U11676 (N_11676,N_6449,N_6175);
nor U11677 (N_11677,N_6263,N_7514);
nor U11678 (N_11678,N_8999,N_6811);
nor U11679 (N_11679,N_6428,N_6477);
or U11680 (N_11680,N_7193,N_8982);
nor U11681 (N_11681,N_6378,N_8014);
or U11682 (N_11682,N_6916,N_6431);
or U11683 (N_11683,N_7244,N_7917);
nor U11684 (N_11684,N_7172,N_6831);
nor U11685 (N_11685,N_8452,N_8770);
or U11686 (N_11686,N_7953,N_7017);
nor U11687 (N_11687,N_6732,N_7174);
nand U11688 (N_11688,N_7821,N_8193);
and U11689 (N_11689,N_8313,N_6899);
and U11690 (N_11690,N_6330,N_8447);
nor U11691 (N_11691,N_8365,N_8829);
nor U11692 (N_11692,N_8657,N_6125);
and U11693 (N_11693,N_7048,N_8354);
and U11694 (N_11694,N_6258,N_7409);
or U11695 (N_11695,N_8620,N_7738);
nor U11696 (N_11696,N_7754,N_6844);
nor U11697 (N_11697,N_8699,N_6829);
and U11698 (N_11698,N_8600,N_8213);
nand U11699 (N_11699,N_7484,N_6330);
nand U11700 (N_11700,N_7802,N_7109);
nand U11701 (N_11701,N_6794,N_6083);
or U11702 (N_11702,N_7282,N_6725);
or U11703 (N_11703,N_8689,N_6811);
or U11704 (N_11704,N_7385,N_6793);
or U11705 (N_11705,N_7921,N_7116);
and U11706 (N_11706,N_8688,N_7819);
nor U11707 (N_11707,N_6054,N_6275);
nor U11708 (N_11708,N_8883,N_7187);
and U11709 (N_11709,N_7474,N_7368);
nand U11710 (N_11710,N_6210,N_6939);
nor U11711 (N_11711,N_7786,N_6920);
or U11712 (N_11712,N_8546,N_6348);
or U11713 (N_11713,N_6127,N_6662);
or U11714 (N_11714,N_8337,N_7024);
or U11715 (N_11715,N_6356,N_8506);
or U11716 (N_11716,N_8552,N_7015);
nor U11717 (N_11717,N_8781,N_6422);
and U11718 (N_11718,N_6109,N_8166);
and U11719 (N_11719,N_6567,N_6350);
and U11720 (N_11720,N_8344,N_8018);
nor U11721 (N_11721,N_8042,N_8964);
or U11722 (N_11722,N_7052,N_8710);
or U11723 (N_11723,N_8633,N_8336);
and U11724 (N_11724,N_8762,N_8115);
and U11725 (N_11725,N_8379,N_8716);
nand U11726 (N_11726,N_6425,N_6725);
and U11727 (N_11727,N_7470,N_8340);
nand U11728 (N_11728,N_7105,N_8410);
nand U11729 (N_11729,N_6805,N_7133);
nand U11730 (N_11730,N_6870,N_8938);
and U11731 (N_11731,N_6673,N_7778);
nor U11732 (N_11732,N_6253,N_7712);
nor U11733 (N_11733,N_6318,N_6194);
and U11734 (N_11734,N_7215,N_7160);
nor U11735 (N_11735,N_8852,N_8481);
nand U11736 (N_11736,N_8841,N_6661);
or U11737 (N_11737,N_7651,N_6214);
or U11738 (N_11738,N_8609,N_7121);
nand U11739 (N_11739,N_8202,N_8349);
and U11740 (N_11740,N_8950,N_6966);
and U11741 (N_11741,N_7849,N_6596);
nor U11742 (N_11742,N_6715,N_8022);
and U11743 (N_11743,N_8690,N_8148);
or U11744 (N_11744,N_8588,N_7387);
nor U11745 (N_11745,N_6948,N_7837);
nand U11746 (N_11746,N_8787,N_8608);
nor U11747 (N_11747,N_8808,N_8011);
nor U11748 (N_11748,N_8516,N_8264);
or U11749 (N_11749,N_6187,N_7554);
nor U11750 (N_11750,N_8939,N_7138);
or U11751 (N_11751,N_6609,N_8583);
nand U11752 (N_11752,N_6850,N_7513);
nand U11753 (N_11753,N_7974,N_8682);
or U11754 (N_11754,N_8167,N_7749);
and U11755 (N_11755,N_6998,N_7986);
nor U11756 (N_11756,N_8124,N_6418);
or U11757 (N_11757,N_7662,N_7875);
and U11758 (N_11758,N_6836,N_7293);
nor U11759 (N_11759,N_7420,N_7280);
nand U11760 (N_11760,N_7238,N_7786);
or U11761 (N_11761,N_7253,N_7871);
nor U11762 (N_11762,N_8680,N_7419);
and U11763 (N_11763,N_6454,N_7703);
and U11764 (N_11764,N_7358,N_7307);
and U11765 (N_11765,N_7124,N_8074);
nor U11766 (N_11766,N_7779,N_6128);
nand U11767 (N_11767,N_6717,N_7346);
and U11768 (N_11768,N_6502,N_6550);
or U11769 (N_11769,N_8546,N_7712);
or U11770 (N_11770,N_6112,N_8827);
or U11771 (N_11771,N_8612,N_8674);
nor U11772 (N_11772,N_6546,N_8010);
nor U11773 (N_11773,N_6989,N_8420);
nand U11774 (N_11774,N_6044,N_6590);
and U11775 (N_11775,N_8117,N_7351);
nand U11776 (N_11776,N_7398,N_7127);
and U11777 (N_11777,N_8913,N_8689);
nor U11778 (N_11778,N_6532,N_6402);
nand U11779 (N_11779,N_6096,N_8610);
and U11780 (N_11780,N_8966,N_8411);
or U11781 (N_11781,N_7223,N_7746);
and U11782 (N_11782,N_7181,N_6306);
nor U11783 (N_11783,N_7237,N_6257);
and U11784 (N_11784,N_8466,N_7063);
nor U11785 (N_11785,N_8690,N_8389);
and U11786 (N_11786,N_6757,N_6748);
nand U11787 (N_11787,N_8177,N_7558);
and U11788 (N_11788,N_7301,N_6187);
or U11789 (N_11789,N_7095,N_6152);
or U11790 (N_11790,N_6131,N_8334);
nand U11791 (N_11791,N_8320,N_7802);
or U11792 (N_11792,N_7771,N_7918);
nor U11793 (N_11793,N_6228,N_6112);
and U11794 (N_11794,N_6812,N_6615);
nor U11795 (N_11795,N_7797,N_8883);
and U11796 (N_11796,N_6709,N_8519);
nor U11797 (N_11797,N_7228,N_6899);
nand U11798 (N_11798,N_8182,N_8450);
nand U11799 (N_11799,N_8345,N_6069);
and U11800 (N_11800,N_8687,N_7960);
and U11801 (N_11801,N_7808,N_6990);
nor U11802 (N_11802,N_6485,N_6768);
or U11803 (N_11803,N_7651,N_6020);
or U11804 (N_11804,N_6726,N_7513);
and U11805 (N_11805,N_7451,N_7067);
xor U11806 (N_11806,N_8049,N_6326);
or U11807 (N_11807,N_6253,N_7330);
and U11808 (N_11808,N_8960,N_6796);
nand U11809 (N_11809,N_8037,N_7531);
nand U11810 (N_11810,N_7742,N_7183);
or U11811 (N_11811,N_8106,N_7664);
nor U11812 (N_11812,N_7658,N_8772);
or U11813 (N_11813,N_7696,N_7713);
nand U11814 (N_11814,N_6154,N_8175);
nor U11815 (N_11815,N_6298,N_6004);
nor U11816 (N_11816,N_7350,N_7951);
nand U11817 (N_11817,N_6624,N_6399);
or U11818 (N_11818,N_8894,N_7405);
and U11819 (N_11819,N_8117,N_6728);
nand U11820 (N_11820,N_6308,N_6539);
nor U11821 (N_11821,N_7908,N_7859);
or U11822 (N_11822,N_8797,N_8505);
nand U11823 (N_11823,N_8863,N_7785);
and U11824 (N_11824,N_7614,N_7174);
or U11825 (N_11825,N_6180,N_7944);
or U11826 (N_11826,N_7042,N_6363);
or U11827 (N_11827,N_7683,N_6511);
and U11828 (N_11828,N_8995,N_6476);
or U11829 (N_11829,N_6980,N_8755);
and U11830 (N_11830,N_8337,N_7201);
and U11831 (N_11831,N_6106,N_8579);
nor U11832 (N_11832,N_6759,N_7288);
and U11833 (N_11833,N_6639,N_6526);
nor U11834 (N_11834,N_7635,N_7482);
nand U11835 (N_11835,N_8663,N_7834);
nor U11836 (N_11836,N_7840,N_6934);
nand U11837 (N_11837,N_8266,N_6961);
nand U11838 (N_11838,N_7371,N_8806);
or U11839 (N_11839,N_6768,N_8511);
and U11840 (N_11840,N_7337,N_6158);
nor U11841 (N_11841,N_6198,N_6708);
nand U11842 (N_11842,N_6187,N_6812);
nor U11843 (N_11843,N_8381,N_7601);
nand U11844 (N_11844,N_7485,N_8181);
xor U11845 (N_11845,N_6478,N_6724);
or U11846 (N_11846,N_6535,N_8739);
nor U11847 (N_11847,N_7045,N_8221);
and U11848 (N_11848,N_8674,N_6955);
and U11849 (N_11849,N_6417,N_6431);
or U11850 (N_11850,N_8954,N_7552);
and U11851 (N_11851,N_8487,N_7778);
nand U11852 (N_11852,N_8507,N_6056);
and U11853 (N_11853,N_8736,N_8335);
nor U11854 (N_11854,N_6624,N_8869);
nand U11855 (N_11855,N_8159,N_7119);
or U11856 (N_11856,N_6763,N_7696);
and U11857 (N_11857,N_7001,N_6223);
or U11858 (N_11858,N_7826,N_8289);
nand U11859 (N_11859,N_6171,N_8355);
or U11860 (N_11860,N_8845,N_8361);
or U11861 (N_11861,N_6815,N_8454);
nand U11862 (N_11862,N_7459,N_8144);
or U11863 (N_11863,N_7983,N_6025);
and U11864 (N_11864,N_6565,N_7211);
nor U11865 (N_11865,N_6354,N_7147);
nor U11866 (N_11866,N_7863,N_8352);
nor U11867 (N_11867,N_8107,N_6950);
nand U11868 (N_11868,N_8528,N_7126);
nor U11869 (N_11869,N_6900,N_7044);
and U11870 (N_11870,N_7651,N_8819);
or U11871 (N_11871,N_7600,N_6678);
and U11872 (N_11872,N_8449,N_6169);
nand U11873 (N_11873,N_7282,N_7739);
and U11874 (N_11874,N_7805,N_6909);
or U11875 (N_11875,N_6101,N_8142);
or U11876 (N_11876,N_6829,N_6630);
or U11877 (N_11877,N_6956,N_6811);
xnor U11878 (N_11878,N_6644,N_7570);
or U11879 (N_11879,N_8510,N_6379);
or U11880 (N_11880,N_6086,N_6316);
or U11881 (N_11881,N_7437,N_7189);
nand U11882 (N_11882,N_7865,N_8154);
nor U11883 (N_11883,N_8737,N_8602);
or U11884 (N_11884,N_8702,N_8170);
nand U11885 (N_11885,N_6308,N_8623);
nand U11886 (N_11886,N_6797,N_7100);
and U11887 (N_11887,N_7172,N_7971);
or U11888 (N_11888,N_8388,N_6242);
or U11889 (N_11889,N_6986,N_8232);
and U11890 (N_11890,N_8111,N_8984);
nand U11891 (N_11891,N_6247,N_8654);
or U11892 (N_11892,N_8684,N_6517);
and U11893 (N_11893,N_7534,N_6668);
nor U11894 (N_11894,N_6905,N_8196);
or U11895 (N_11895,N_7371,N_8986);
or U11896 (N_11896,N_8728,N_7397);
nand U11897 (N_11897,N_7543,N_8169);
nor U11898 (N_11898,N_7594,N_8061);
nor U11899 (N_11899,N_6022,N_6155);
or U11900 (N_11900,N_7906,N_7794);
and U11901 (N_11901,N_8168,N_7360);
nand U11902 (N_11902,N_8919,N_8961);
or U11903 (N_11903,N_8127,N_6920);
or U11904 (N_11904,N_8875,N_7784);
or U11905 (N_11905,N_6932,N_7999);
and U11906 (N_11906,N_8981,N_6836);
nand U11907 (N_11907,N_8503,N_7596);
nor U11908 (N_11908,N_8644,N_7580);
nand U11909 (N_11909,N_8291,N_6200);
and U11910 (N_11910,N_8266,N_7748);
and U11911 (N_11911,N_6485,N_8187);
nand U11912 (N_11912,N_8908,N_8762);
nand U11913 (N_11913,N_8215,N_7686);
and U11914 (N_11914,N_6127,N_7340);
nand U11915 (N_11915,N_6089,N_6275);
nor U11916 (N_11916,N_6455,N_7441);
or U11917 (N_11917,N_7030,N_8433);
and U11918 (N_11918,N_8915,N_7180);
and U11919 (N_11919,N_6829,N_7420);
or U11920 (N_11920,N_8123,N_7328);
nor U11921 (N_11921,N_8493,N_7417);
and U11922 (N_11922,N_7368,N_8642);
nor U11923 (N_11923,N_7773,N_8365);
nand U11924 (N_11924,N_7094,N_8416);
nand U11925 (N_11925,N_7597,N_8144);
nor U11926 (N_11926,N_8046,N_6686);
and U11927 (N_11927,N_6501,N_7077);
nand U11928 (N_11928,N_8745,N_8705);
and U11929 (N_11929,N_6679,N_8230);
and U11930 (N_11930,N_8838,N_7820);
and U11931 (N_11931,N_8072,N_8971);
nand U11932 (N_11932,N_7787,N_6129);
and U11933 (N_11933,N_7582,N_8648);
xor U11934 (N_11934,N_7216,N_6308);
or U11935 (N_11935,N_6917,N_7021);
and U11936 (N_11936,N_8356,N_7595);
nor U11937 (N_11937,N_7205,N_6090);
or U11938 (N_11938,N_7330,N_6287);
nor U11939 (N_11939,N_6834,N_6114);
and U11940 (N_11940,N_6138,N_7475);
nand U11941 (N_11941,N_8429,N_6450);
nand U11942 (N_11942,N_8537,N_7369);
nor U11943 (N_11943,N_8560,N_6014);
nand U11944 (N_11944,N_8218,N_8283);
or U11945 (N_11945,N_6261,N_7004);
and U11946 (N_11946,N_6371,N_6572);
or U11947 (N_11947,N_6688,N_8058);
or U11948 (N_11948,N_8072,N_8129);
nor U11949 (N_11949,N_7955,N_6911);
nor U11950 (N_11950,N_7966,N_8019);
nor U11951 (N_11951,N_7773,N_8812);
nor U11952 (N_11952,N_6694,N_6251);
nor U11953 (N_11953,N_7427,N_6342);
and U11954 (N_11954,N_7732,N_6726);
nand U11955 (N_11955,N_6544,N_6314);
xor U11956 (N_11956,N_6023,N_6222);
nor U11957 (N_11957,N_8000,N_8193);
and U11958 (N_11958,N_6115,N_7496);
or U11959 (N_11959,N_7602,N_8568);
xnor U11960 (N_11960,N_8583,N_7989);
and U11961 (N_11961,N_6064,N_8489);
and U11962 (N_11962,N_8246,N_7150);
or U11963 (N_11963,N_7487,N_6184);
nand U11964 (N_11964,N_8251,N_6182);
or U11965 (N_11965,N_8844,N_6893);
nor U11966 (N_11966,N_7502,N_6701);
nor U11967 (N_11967,N_8556,N_7469);
nand U11968 (N_11968,N_8485,N_7808);
nand U11969 (N_11969,N_7428,N_8431);
or U11970 (N_11970,N_6449,N_7551);
or U11971 (N_11971,N_6881,N_8864);
and U11972 (N_11972,N_7952,N_8458);
and U11973 (N_11973,N_8164,N_7307);
and U11974 (N_11974,N_7037,N_6197);
nor U11975 (N_11975,N_7814,N_7742);
nand U11976 (N_11976,N_6799,N_6407);
or U11977 (N_11977,N_6461,N_8140);
or U11978 (N_11978,N_8748,N_7904);
and U11979 (N_11979,N_8595,N_6448);
nor U11980 (N_11980,N_6528,N_8441);
or U11981 (N_11981,N_7359,N_6397);
nand U11982 (N_11982,N_6153,N_8130);
or U11983 (N_11983,N_6630,N_6425);
nand U11984 (N_11984,N_6221,N_7505);
nor U11985 (N_11985,N_8517,N_7036);
nand U11986 (N_11986,N_6475,N_6830);
nor U11987 (N_11987,N_6572,N_8445);
or U11988 (N_11988,N_6826,N_6886);
nand U11989 (N_11989,N_6761,N_8136);
or U11990 (N_11990,N_7359,N_7287);
nor U11991 (N_11991,N_8930,N_7280);
nor U11992 (N_11992,N_6524,N_6008);
nor U11993 (N_11993,N_6444,N_8026);
and U11994 (N_11994,N_7687,N_8728);
and U11995 (N_11995,N_7943,N_8752);
or U11996 (N_11996,N_7107,N_8843);
nand U11997 (N_11997,N_6888,N_6997);
nor U11998 (N_11998,N_7507,N_7007);
nand U11999 (N_11999,N_8190,N_6409);
nor U12000 (N_12000,N_11720,N_11514);
nand U12001 (N_12001,N_11815,N_10867);
and U12002 (N_12002,N_10782,N_11869);
and U12003 (N_12003,N_10722,N_11746);
nor U12004 (N_12004,N_10197,N_11049);
nor U12005 (N_12005,N_10961,N_10460);
and U12006 (N_12006,N_10776,N_10034);
nor U12007 (N_12007,N_10304,N_10949);
nor U12008 (N_12008,N_10063,N_11292);
nor U12009 (N_12009,N_9962,N_11429);
or U12010 (N_12010,N_10367,N_10480);
nor U12011 (N_12011,N_11233,N_9023);
and U12012 (N_12012,N_9046,N_9881);
nand U12013 (N_12013,N_11252,N_9696);
or U12014 (N_12014,N_10018,N_9349);
nor U12015 (N_12015,N_9328,N_9010);
nor U12016 (N_12016,N_11597,N_9648);
or U12017 (N_12017,N_10102,N_10195);
or U12018 (N_12018,N_9738,N_11439);
and U12019 (N_12019,N_10507,N_11316);
or U12020 (N_12020,N_11324,N_11772);
nor U12021 (N_12021,N_9047,N_10407);
xnor U12022 (N_12022,N_9975,N_9189);
nor U12023 (N_12023,N_11727,N_9906);
and U12024 (N_12024,N_10096,N_9741);
nand U12025 (N_12025,N_10866,N_9626);
nand U12026 (N_12026,N_11030,N_9569);
nand U12027 (N_12027,N_9753,N_11731);
or U12028 (N_12028,N_10504,N_10033);
nand U12029 (N_12029,N_10157,N_10955);
nor U12030 (N_12030,N_11035,N_10899);
nand U12031 (N_12031,N_11663,N_11793);
or U12032 (N_12032,N_11794,N_10758);
nand U12033 (N_12033,N_11430,N_10086);
or U12034 (N_12034,N_9716,N_9922);
nand U12035 (N_12035,N_11799,N_11064);
nand U12036 (N_12036,N_10750,N_10649);
nor U12037 (N_12037,N_10248,N_9750);
nand U12038 (N_12038,N_11048,N_9791);
or U12039 (N_12039,N_11150,N_11238);
nand U12040 (N_12040,N_11997,N_9462);
or U12041 (N_12041,N_11312,N_10793);
nand U12042 (N_12042,N_9680,N_9173);
nor U12043 (N_12043,N_10516,N_11497);
or U12044 (N_12044,N_11420,N_10419);
and U12045 (N_12045,N_10119,N_11465);
or U12046 (N_12046,N_9637,N_11847);
nand U12047 (N_12047,N_10022,N_9083);
and U12048 (N_12048,N_9100,N_11448);
nand U12049 (N_12049,N_11938,N_10999);
nor U12050 (N_12050,N_10055,N_10360);
nor U12051 (N_12051,N_11025,N_10090);
nand U12052 (N_12052,N_11128,N_11432);
nand U12053 (N_12053,N_11594,N_11929);
nor U12054 (N_12054,N_10801,N_9548);
nor U12055 (N_12055,N_10631,N_9103);
nand U12056 (N_12056,N_11068,N_11528);
or U12057 (N_12057,N_11802,N_11040);
nor U12058 (N_12058,N_11708,N_11754);
or U12059 (N_12059,N_10672,N_9967);
nor U12060 (N_12060,N_10957,N_10006);
nor U12061 (N_12061,N_11995,N_10097);
and U12062 (N_12062,N_9534,N_10797);
and U12063 (N_12063,N_11350,N_9774);
or U12064 (N_12064,N_10436,N_10281);
and U12065 (N_12065,N_9092,N_11970);
nand U12066 (N_12066,N_9447,N_10837);
nor U12067 (N_12067,N_10911,N_9702);
and U12068 (N_12068,N_11879,N_11541);
or U12069 (N_12069,N_10819,N_11954);
and U12070 (N_12070,N_11349,N_9008);
nand U12071 (N_12071,N_9535,N_11018);
xnor U12072 (N_12072,N_10994,N_9979);
nand U12073 (N_12073,N_9235,N_11808);
nor U12074 (N_12074,N_10939,N_9985);
xor U12075 (N_12075,N_10679,N_11575);
nand U12076 (N_12076,N_10421,N_10152);
and U12077 (N_12077,N_11910,N_10240);
nor U12078 (N_12078,N_10310,N_10476);
and U12079 (N_12079,N_11906,N_10379);
and U12080 (N_12080,N_9505,N_11552);
nor U12081 (N_12081,N_10676,N_9486);
and U12082 (N_12082,N_11688,N_9164);
nor U12083 (N_12083,N_11608,N_11096);
or U12084 (N_12084,N_9295,N_10438);
nor U12085 (N_12085,N_9986,N_11494);
and U12086 (N_12086,N_11763,N_10920);
nor U12087 (N_12087,N_10149,N_10875);
or U12088 (N_12088,N_10326,N_11210);
nand U12089 (N_12089,N_10146,N_9617);
nand U12090 (N_12090,N_10049,N_11523);
or U12091 (N_12091,N_11783,N_11409);
nor U12092 (N_12092,N_9554,N_9043);
or U12093 (N_12093,N_9778,N_11681);
or U12094 (N_12094,N_11394,N_9801);
nand U12095 (N_12095,N_9378,N_9921);
and U12096 (N_12096,N_10478,N_10740);
nand U12097 (N_12097,N_11134,N_11299);
nand U12098 (N_12098,N_11640,N_9226);
nand U12099 (N_12099,N_11200,N_10735);
and U12100 (N_12100,N_10854,N_9412);
or U12101 (N_12101,N_11917,N_11185);
nand U12102 (N_12102,N_10617,N_11986);
and U12103 (N_12103,N_10330,N_10571);
nor U12104 (N_12104,N_10641,N_9823);
nand U12105 (N_12105,N_10950,N_11849);
nand U12106 (N_12106,N_9846,N_11726);
nor U12107 (N_12107,N_9983,N_9786);
nand U12108 (N_12108,N_10968,N_11700);
nand U12109 (N_12109,N_10175,N_9803);
or U12110 (N_12110,N_9080,N_9176);
and U12111 (N_12111,N_10675,N_9067);
nor U12112 (N_12112,N_11492,N_11722);
nand U12113 (N_12113,N_9667,N_9491);
nor U12114 (N_12114,N_11736,N_10331);
nand U12115 (N_12115,N_11406,N_10332);
and U12116 (N_12116,N_10491,N_11883);
nor U12117 (N_12117,N_9087,N_11805);
nand U12118 (N_12118,N_10285,N_10524);
or U12119 (N_12119,N_10342,N_10868);
nor U12120 (N_12120,N_9317,N_9198);
nor U12121 (N_12121,N_10825,N_9113);
or U12122 (N_12122,N_9597,N_10302);
nand U12123 (N_12123,N_9210,N_10019);
or U12124 (N_12124,N_11493,N_9136);
or U12125 (N_12125,N_11216,N_9065);
nand U12126 (N_12126,N_9187,N_10349);
or U12127 (N_12127,N_9611,N_11180);
and U12128 (N_12128,N_10630,N_9155);
or U12129 (N_12129,N_10880,N_10468);
nor U12130 (N_12130,N_11126,N_11199);
nor U12131 (N_12131,N_11674,N_11240);
nor U12132 (N_12132,N_10395,N_11551);
nor U12133 (N_12133,N_9666,N_10912);
nor U12134 (N_12134,N_9821,N_11374);
and U12135 (N_12135,N_11670,N_11376);
or U12136 (N_12136,N_11297,N_9790);
or U12137 (N_12137,N_9478,N_11827);
or U12138 (N_12138,N_10351,N_10946);
nand U12139 (N_12139,N_11837,N_9565);
nor U12140 (N_12140,N_9674,N_9576);
nand U12141 (N_12141,N_10665,N_10513);
and U12142 (N_12142,N_9280,N_9722);
nand U12143 (N_12143,N_9853,N_10284);
nor U12144 (N_12144,N_10493,N_9630);
nor U12145 (N_12145,N_10227,N_10970);
or U12146 (N_12146,N_10303,N_9146);
and U12147 (N_12147,N_10600,N_9049);
or U12148 (N_12148,N_10267,N_10864);
nand U12149 (N_12149,N_11217,N_11400);
nor U12150 (N_12150,N_10363,N_10466);
nand U12151 (N_12151,N_11780,N_11739);
nor U12152 (N_12152,N_9956,N_10910);
nand U12153 (N_12153,N_10522,N_9684);
nand U12154 (N_12154,N_11074,N_9813);
and U12155 (N_12155,N_11154,N_10228);
nor U12156 (N_12156,N_10323,N_10652);
or U12157 (N_12157,N_11656,N_9015);
or U12158 (N_12158,N_11358,N_9718);
nand U12159 (N_12159,N_10596,N_11996);
nor U12160 (N_12160,N_9923,N_11286);
nor U12161 (N_12161,N_9446,N_10568);
nand U12162 (N_12162,N_11109,N_9201);
or U12163 (N_12163,N_9608,N_10101);
and U12164 (N_12164,N_11012,N_10039);
nand U12165 (N_12165,N_10014,N_9188);
nor U12166 (N_12166,N_10509,N_11692);
and U12167 (N_12167,N_11595,N_11584);
nor U12168 (N_12168,N_10664,N_10009);
or U12169 (N_12169,N_9581,N_9305);
nor U12170 (N_12170,N_10233,N_11268);
or U12171 (N_12171,N_9732,N_11933);
nand U12172 (N_12172,N_9397,N_11566);
or U12173 (N_12173,N_11717,N_9874);
nand U12174 (N_12174,N_10321,N_10122);
and U12175 (N_12175,N_9913,N_10934);
nor U12176 (N_12176,N_9744,N_10807);
nor U12177 (N_12177,N_11609,N_10889);
or U12178 (N_12178,N_11082,N_10364);
nand U12179 (N_12179,N_9997,N_10184);
and U12180 (N_12180,N_10215,N_11713);
nand U12181 (N_12181,N_9493,N_9658);
nand U12182 (N_12182,N_11352,N_10450);
xor U12183 (N_12183,N_10808,N_9629);
nand U12184 (N_12184,N_9622,N_9589);
nor U12185 (N_12185,N_11866,N_10528);
or U12186 (N_12186,N_10132,N_10291);
and U12187 (N_12187,N_11295,N_11946);
nor U12188 (N_12188,N_9450,N_10757);
nor U12189 (N_12189,N_11673,N_10359);
and U12190 (N_12190,N_10206,N_11577);
nand U12191 (N_12191,N_10441,N_11775);
and U12192 (N_12192,N_10702,N_10668);
or U12193 (N_12193,N_10903,N_9069);
or U12194 (N_12194,N_10451,N_11257);
and U12195 (N_12195,N_10645,N_11657);
nand U12196 (N_12196,N_11949,N_10794);
nor U12197 (N_12197,N_9763,N_10163);
nor U12198 (N_12198,N_9789,N_10106);
nor U12199 (N_12199,N_9935,N_11935);
xor U12200 (N_12200,N_9172,N_9818);
or U12201 (N_12201,N_10979,N_10835);
nand U12202 (N_12202,N_9248,N_11858);
and U12203 (N_12203,N_9945,N_11318);
nand U12204 (N_12204,N_11275,N_10357);
and U12205 (N_12205,N_11481,N_10452);
nor U12206 (N_12206,N_9588,N_11991);
nand U12207 (N_12207,N_9286,N_9640);
and U12208 (N_12208,N_10288,N_9476);
and U12209 (N_12209,N_9503,N_10274);
nand U12210 (N_12210,N_11999,N_10339);
and U12211 (N_12211,N_10658,N_10433);
and U12212 (N_12212,N_9619,N_9518);
nor U12213 (N_12213,N_10943,N_9322);
and U12214 (N_12214,N_9401,N_10691);
or U12215 (N_12215,N_10539,N_10021);
nand U12216 (N_12216,N_9151,N_11852);
nor U12217 (N_12217,N_11186,N_10988);
or U12218 (N_12218,N_10320,N_10335);
nand U12219 (N_12219,N_10148,N_9101);
nand U12220 (N_12220,N_9907,N_10947);
nor U12221 (N_12221,N_9085,N_11690);
nor U12222 (N_12222,N_10851,N_11581);
and U12223 (N_12223,N_10699,N_9794);
or U12224 (N_12224,N_11458,N_10881);
and U12225 (N_12225,N_10246,N_11359);
and U12226 (N_12226,N_10928,N_10677);
nor U12227 (N_12227,N_11002,N_9471);
nand U12228 (N_12228,N_10860,N_9893);
nor U12229 (N_12229,N_11418,N_10254);
and U12230 (N_12230,N_10884,N_10951);
or U12231 (N_12231,N_10412,N_9384);
nor U12232 (N_12232,N_9454,N_11982);
nor U12233 (N_12233,N_10669,N_10511);
or U12234 (N_12234,N_10858,N_10377);
and U12235 (N_12235,N_9185,N_10142);
nand U12236 (N_12236,N_10448,N_11101);
nand U12237 (N_12237,N_11930,N_9810);
nor U12238 (N_12238,N_11983,N_10906);
or U12239 (N_12239,N_11784,N_10814);
or U12240 (N_12240,N_9916,N_11426);
nor U12241 (N_12241,N_9819,N_10065);
xor U12242 (N_12242,N_9020,N_11476);
or U12243 (N_12243,N_10088,N_9017);
nand U12244 (N_12244,N_11165,N_9623);
or U12245 (N_12245,N_9169,N_9636);
xnor U12246 (N_12246,N_9969,N_9053);
or U12247 (N_12247,N_11239,N_10201);
nand U12248 (N_12248,N_9267,N_9281);
nor U12249 (N_12249,N_9138,N_10719);
nor U12250 (N_12250,N_10959,N_9760);
nand U12251 (N_12251,N_9426,N_11554);
and U12252 (N_12252,N_9869,N_11117);
and U12253 (N_12253,N_11561,N_10742);
or U12254 (N_12254,N_11567,N_10888);
or U12255 (N_12255,N_10043,N_10005);
nand U12256 (N_12256,N_11621,N_11188);
nor U12257 (N_12257,N_11612,N_10289);
nand U12258 (N_12258,N_9645,N_9542);
and U12259 (N_12259,N_9770,N_11471);
or U12260 (N_12260,N_11704,N_10116);
nor U12261 (N_12261,N_10817,N_11521);
and U12262 (N_12262,N_11389,N_11994);
nor U12263 (N_12263,N_9217,N_11503);
or U12264 (N_12264,N_9757,N_11797);
or U12265 (N_12265,N_9099,N_11510);
or U12266 (N_12266,N_9521,N_10038);
nor U12267 (N_12267,N_9114,N_9353);
and U12268 (N_12268,N_11496,N_10559);
or U12269 (N_12269,N_9119,N_11593);
and U12270 (N_12270,N_10685,N_9829);
nor U12271 (N_12271,N_11036,N_11236);
or U12272 (N_12272,N_10640,N_10054);
nor U12273 (N_12273,N_10381,N_9929);
nor U12274 (N_12274,N_10371,N_9939);
or U12275 (N_12275,N_9319,N_10185);
nand U12276 (N_12276,N_9894,N_11112);
nand U12277 (N_12277,N_10885,N_9538);
nand U12278 (N_12278,N_10662,N_11789);
nand U12279 (N_12279,N_9954,N_11020);
nand U12280 (N_12280,N_10762,N_9098);
or U12281 (N_12281,N_11029,N_11563);
and U12282 (N_12282,N_9405,N_10208);
or U12283 (N_12283,N_11816,N_11872);
nor U12284 (N_12284,N_10455,N_10538);
nand U12285 (N_12285,N_9650,N_9037);
or U12286 (N_12286,N_9805,N_11054);
nand U12287 (N_12287,N_9867,N_9897);
and U12288 (N_12288,N_10815,N_11332);
or U12289 (N_12289,N_11363,N_11310);
nor U12290 (N_12290,N_9165,N_11960);
and U12291 (N_12291,N_9018,N_10989);
and U12292 (N_12292,N_10060,N_11662);
or U12293 (N_12293,N_11173,N_9734);
and U12294 (N_12294,N_10995,N_11806);
or U12295 (N_12295,N_10399,N_10779);
nor U12296 (N_12296,N_10427,N_9614);
nand U12297 (N_12297,N_11807,N_10047);
nand U12298 (N_12298,N_10874,N_11707);
or U12299 (N_12299,N_10389,N_10481);
nand U12300 (N_12300,N_11078,N_11103);
and U12301 (N_12301,N_10711,N_11027);
nand U12302 (N_12302,N_11072,N_11308);
nand U12303 (N_12303,N_10290,N_9844);
and U12304 (N_12304,N_9501,N_9693);
or U12305 (N_12305,N_10000,N_10615);
or U12306 (N_12306,N_11628,N_10512);
nand U12307 (N_12307,N_11606,N_9232);
or U12308 (N_12308,N_9932,N_9208);
and U12309 (N_12309,N_10158,N_11699);
or U12310 (N_12310,N_9560,N_11513);
nor U12311 (N_12311,N_10373,N_9283);
or U12312 (N_12312,N_10397,N_10456);
nand U12313 (N_12313,N_10414,N_10301);
nor U12314 (N_12314,N_11668,N_11485);
nand U12315 (N_12315,N_10471,N_10523);
nand U12316 (N_12316,N_10527,N_11511);
and U12317 (N_12317,N_11532,N_11742);
nor U12318 (N_12318,N_9377,N_11277);
and U12319 (N_12319,N_10725,N_11287);
and U12320 (N_12320,N_11206,N_10873);
or U12321 (N_12321,N_10869,N_10327);
nand U12322 (N_12322,N_10941,N_10862);
nor U12323 (N_12323,N_9263,N_9701);
and U12324 (N_12324,N_11522,N_10143);
or U12325 (N_12325,N_11665,N_10520);
nor U12326 (N_12326,N_10140,N_11187);
nand U12327 (N_12327,N_11119,N_11826);
and U12328 (N_12328,N_9552,N_11371);
and U12329 (N_12329,N_11417,N_9127);
nand U12330 (N_12330,N_9591,N_9292);
nand U12331 (N_12331,N_10264,N_10804);
and U12332 (N_12332,N_11208,N_9812);
and U12333 (N_12333,N_9120,N_9337);
nor U12334 (N_12334,N_10551,N_9430);
and U12335 (N_12335,N_10565,N_9063);
and U12336 (N_12336,N_10714,N_10077);
nor U12337 (N_12337,N_10969,N_9093);
nor U12338 (N_12338,N_10966,N_11644);
and U12339 (N_12339,N_11907,N_10891);
nand U12340 (N_12340,N_11832,N_9938);
and U12341 (N_12341,N_11570,N_9920);
nor U12342 (N_12342,N_9441,N_10189);
nand U12343 (N_12343,N_9381,N_10883);
and U12344 (N_12344,N_10984,N_9871);
and U12345 (N_12345,N_9129,N_9889);
and U12346 (N_12346,N_9348,N_11223);
and U12347 (N_12347,N_10094,N_11571);
and U12348 (N_12348,N_10907,N_9695);
or U12349 (N_12349,N_10890,N_11242);
nor U12350 (N_12350,N_10960,N_9059);
and U12351 (N_12351,N_10730,N_10775);
and U12352 (N_12352,N_11823,N_10078);
nor U12353 (N_12353,N_11331,N_9032);
nand U12354 (N_12354,N_10701,N_9496);
nor U12355 (N_12355,N_11886,N_10982);
or U12356 (N_12356,N_11464,N_10172);
nor U12357 (N_12357,N_11042,N_9870);
and U12358 (N_12358,N_11122,N_11755);
nand U12359 (N_12359,N_10354,N_10865);
nand U12360 (N_12360,N_11762,N_11667);
or U12361 (N_12361,N_9651,N_11360);
nor U12362 (N_12362,N_9026,N_11655);
or U12363 (N_12363,N_10216,N_10297);
nor U12364 (N_12364,N_9105,N_10820);
nand U12365 (N_12365,N_11305,N_10813);
or U12366 (N_12366,N_10435,N_9536);
nor U12367 (N_12367,N_9302,N_10805);
nor U12368 (N_12368,N_9035,N_11457);
or U12369 (N_12369,N_9665,N_9371);
or U12370 (N_12370,N_9191,N_10278);
and U12371 (N_12371,N_9911,N_9091);
nor U12372 (N_12372,N_9331,N_10341);
and U12373 (N_12373,N_10202,N_10986);
nand U12374 (N_12374,N_9561,N_11769);
nor U12375 (N_12375,N_11824,N_9927);
nor U12376 (N_12376,N_10566,N_11839);
or U12377 (N_12377,N_10235,N_10159);
nand U12378 (N_12378,N_11004,N_10541);
or U12379 (N_12379,N_11431,N_10650);
and U12380 (N_12380,N_10413,N_11683);
nor U12381 (N_12381,N_11424,N_11489);
nor U12382 (N_12382,N_10695,N_9711);
nor U12383 (N_12383,N_11868,N_11467);
or U12384 (N_12384,N_9213,N_9288);
nand U12385 (N_12385,N_11893,N_10895);
or U12386 (N_12386,N_9137,N_11266);
or U12387 (N_12387,N_10325,N_11153);
nor U12388 (N_12388,N_11136,N_9948);
nand U12389 (N_12389,N_10315,N_9679);
nand U12390 (N_12390,N_9346,N_11709);
and U12391 (N_12391,N_9311,N_9316);
and U12392 (N_12392,N_10382,N_9585);
and U12393 (N_12393,N_10603,N_10802);
nand U12394 (N_12394,N_11801,N_11841);
and U12395 (N_12395,N_11250,N_10534);
nor U12396 (N_12396,N_9130,N_10109);
and U12397 (N_12397,N_9815,N_11901);
nand U12398 (N_12398,N_9837,N_11047);
nor U12399 (N_12399,N_10066,N_9743);
nor U12400 (N_12400,N_11618,N_10337);
or U12401 (N_12401,N_10422,N_11081);
or U12402 (N_12402,N_11509,N_9102);
nand U12403 (N_12403,N_10688,N_10863);
nor U12404 (N_12404,N_11386,N_11803);
nor U12405 (N_12405,N_10255,N_11262);
or U12406 (N_12406,N_11085,N_9982);
or U12407 (N_12407,N_9433,N_11759);
nand U12408 (N_12408,N_9395,N_10404);
or U12409 (N_12409,N_11853,N_11582);
nand U12410 (N_12410,N_9659,N_9301);
or U12411 (N_12411,N_9748,N_11412);
or U12412 (N_12412,N_9603,N_10446);
nand U12413 (N_12413,N_11795,N_10760);
nand U12414 (N_12414,N_11747,N_11626);
and U12415 (N_12415,N_10489,N_9804);
or U12416 (N_12416,N_10400,N_11650);
or U12417 (N_12417,N_9708,N_11854);
or U12418 (N_12418,N_9044,N_11272);
nor U12419 (N_12419,N_11647,N_9124);
or U12420 (N_12420,N_11307,N_10169);
or U12421 (N_12421,N_9207,N_11043);
or U12422 (N_12422,N_9831,N_10732);
nor U12423 (N_12423,N_9500,N_11676);
and U12424 (N_12424,N_11169,N_10062);
nand U12425 (N_12425,N_10686,N_10329);
nor U12426 (N_12426,N_9021,N_9469);
nand U12427 (N_12427,N_11550,N_9313);
nor U12428 (N_12428,N_11725,N_11499);
nor U12429 (N_12429,N_9537,N_9704);
and U12430 (N_12430,N_10369,N_11634);
nand U12431 (N_12431,N_10663,N_10362);
nor U12432 (N_12432,N_11190,N_10705);
nor U12433 (N_12433,N_10188,N_11034);
or U12434 (N_12434,N_10661,N_11918);
nor U12435 (N_12435,N_11836,N_9257);
nor U12436 (N_12436,N_9767,N_11974);
nor U12437 (N_12437,N_11988,N_11786);
and U12438 (N_12438,N_9268,N_9957);
or U12439 (N_12439,N_9571,N_9237);
nand U12440 (N_12440,N_9883,N_9783);
or U12441 (N_12441,N_11347,N_11388);
or U12442 (N_12442,N_10145,N_9621);
nor U12443 (N_12443,N_11671,N_10633);
and U12444 (N_12444,N_9074,N_9360);
or U12445 (N_12445,N_10756,N_10785);
and U12446 (N_12446,N_10876,N_10074);
or U12447 (N_12447,N_10120,N_9545);
or U12448 (N_12448,N_9830,N_9190);
or U12449 (N_12449,N_11124,N_9838);
or U12450 (N_12450,N_9073,N_11357);
and U12451 (N_12451,N_11373,N_9625);
nor U12452 (N_12452,N_10870,N_9931);
and U12453 (N_12453,N_11882,N_9612);
and U12454 (N_12454,N_11985,N_11005);
nor U12455 (N_12455,N_10032,N_10938);
or U12456 (N_12456,N_9294,N_10070);
nand U12457 (N_12457,N_10449,N_9332);
nand U12458 (N_12458,N_9031,N_11181);
nor U12459 (N_12459,N_10684,N_9375);
and U12460 (N_12460,N_9641,N_11053);
nand U12461 (N_12461,N_10643,N_9972);
nand U12462 (N_12462,N_9628,N_11301);
nand U12463 (N_12463,N_9559,N_10575);
and U12464 (N_12464,N_10345,N_10953);
or U12465 (N_12465,N_10418,N_11354);
nand U12466 (N_12466,N_9024,N_10271);
nor U12467 (N_12467,N_11139,N_9011);
or U12468 (N_12468,N_9016,N_10457);
nor U12469 (N_12469,N_11055,N_11044);
and U12470 (N_12470,N_9943,N_9772);
or U12471 (N_12471,N_11435,N_11993);
or U12472 (N_12472,N_10061,N_11328);
nand U12473 (N_12473,N_9516,N_9407);
nand U12474 (N_12474,N_9992,N_10080);
or U12475 (N_12475,N_11959,N_10554);
nand U12476 (N_12476,N_9066,N_11218);
nand U12477 (N_12477,N_11751,N_9271);
or U12478 (N_12478,N_11366,N_9363);
nor U12479 (N_12479,N_9109,N_10855);
and U12480 (N_12480,N_9269,N_10075);
or U12481 (N_12481,N_9175,N_11605);
nand U12482 (N_12482,N_10751,N_10731);
nor U12483 (N_12483,N_11107,N_10707);
nand U12484 (N_12484,N_11760,N_9780);
or U12485 (N_12485,N_10234,N_10764);
nor U12486 (N_12486,N_11201,N_10378);
and U12487 (N_12487,N_11890,N_10879);
and U12488 (N_12488,N_10799,N_10886);
or U12489 (N_12489,N_10445,N_9211);
or U12490 (N_12490,N_9682,N_10967);
and U12491 (N_12491,N_11613,N_10597);
nand U12492 (N_12492,N_10123,N_11711);
or U12493 (N_12493,N_10069,N_11964);
or U12494 (N_12494,N_9551,N_11140);
or U12495 (N_12495,N_9714,N_9978);
or U12496 (N_12496,N_10085,N_11876);
nand U12497 (N_12497,N_11540,N_9825);
nand U12498 (N_12498,N_11822,N_9858);
nor U12499 (N_12499,N_11159,N_10626);
nor U12500 (N_12500,N_9509,N_9220);
or U12501 (N_12501,N_11896,N_9596);
nor U12502 (N_12502,N_11838,N_10980);
and U12503 (N_12503,N_11385,N_11131);
nand U12504 (N_12504,N_10526,N_10211);
nor U12505 (N_12505,N_10391,N_9751);
nand U12506 (N_12506,N_10212,N_10518);
or U12507 (N_12507,N_10041,N_10638);
and U12508 (N_12508,N_11192,N_9902);
and U12509 (N_12509,N_10375,N_10564);
nor U12510 (N_12510,N_10150,N_11779);
nand U12511 (N_12511,N_10843,N_11059);
and U12512 (N_12512,N_9064,N_11888);
nor U12513 (N_12513,N_11247,N_10479);
nor U12514 (N_12514,N_11764,N_11977);
or U12515 (N_12515,N_11939,N_10237);
nand U12516 (N_12516,N_9350,N_11283);
nand U12517 (N_12517,N_9343,N_11014);
or U12518 (N_12518,N_10981,N_10525);
nor U12519 (N_12519,N_11061,N_10914);
and U12520 (N_12520,N_9944,N_9951);
xor U12521 (N_12521,N_9996,N_11965);
nor U12522 (N_12522,N_10057,N_11490);
and U12523 (N_12523,N_9181,N_10558);
nand U12524 (N_12524,N_9477,N_11573);
and U12525 (N_12525,N_9006,N_9307);
nor U12526 (N_12526,N_10738,N_11925);
or U12527 (N_12527,N_9246,N_9251);
nor U12528 (N_12528,N_11303,N_10829);
nor U12529 (N_12529,N_9362,N_9076);
nor U12530 (N_12530,N_11298,N_11263);
nor U12531 (N_12531,N_10519,N_9276);
or U12532 (N_12532,N_10919,N_11198);
nor U12533 (N_12533,N_9697,N_9094);
or U12534 (N_12534,N_11241,N_11003);
nor U12535 (N_12535,N_10733,N_10251);
nand U12536 (N_12536,N_10550,N_9358);
nand U12537 (N_12537,N_10347,N_9086);
nand U12538 (N_12538,N_9333,N_9262);
nor U12539 (N_12539,N_9553,N_11407);
or U12540 (N_12540,N_9525,N_9273);
nor U12541 (N_12541,N_9506,N_10680);
and U12542 (N_12542,N_10352,N_11987);
and U12543 (N_12543,N_10887,N_11587);
nand U12544 (N_12544,N_10747,N_9664);
nor U12545 (N_12545,N_11404,N_11845);
and U12546 (N_12546,N_10100,N_9224);
and U12547 (N_12547,N_10739,N_9886);
nand U12548 (N_12548,N_9759,N_9739);
and U12549 (N_12549,N_9583,N_10486);
nand U12550 (N_12550,N_9683,N_9861);
nor U12551 (N_12551,N_9409,N_9703);
and U12552 (N_12552,N_9231,N_9884);
and U12553 (N_12553,N_10763,N_11041);
nor U12554 (N_12554,N_9466,N_10515);
and U12555 (N_12555,N_9013,N_11620);
or U12556 (N_12556,N_11395,N_9866);
and U12557 (N_12557,N_11781,N_10555);
nor U12558 (N_12558,N_10933,N_9199);
nor U12559 (N_12559,N_9678,N_9900);
xnor U12560 (N_12560,N_11744,N_11791);
nor U12561 (N_12561,N_9299,N_11329);
or U12562 (N_12562,N_11314,N_9038);
or U12563 (N_12563,N_11560,N_9108);
or U12564 (N_12564,N_11313,N_11421);
and U12565 (N_12565,N_10687,N_10192);
nand U12566 (N_12566,N_11518,N_9502);
and U12567 (N_12567,N_11543,N_10114);
nand U12568 (N_12568,N_11261,N_11865);
or U12569 (N_12569,N_9475,N_9354);
nor U12570 (N_12570,N_9272,N_11280);
nand U12571 (N_12571,N_10431,N_10095);
nor U12572 (N_12572,N_10259,N_9421);
or U12573 (N_12573,N_11940,N_11231);
nor U12574 (N_12574,N_9781,N_9484);
and U12575 (N_12575,N_11179,N_11790);
or U12576 (N_12576,N_10570,N_11737);
and U12577 (N_12577,N_11377,N_9782);
nor U12578 (N_12578,N_11071,N_10107);
nor U12579 (N_12579,N_11256,N_10923);
and U12580 (N_12580,N_11279,N_11911);
xor U12581 (N_12581,N_10081,N_11056);
nor U12582 (N_12582,N_10050,N_11527);
or U12583 (N_12583,N_10266,N_11170);
and U12584 (N_12584,N_9737,N_9709);
nor U12585 (N_12585,N_10842,N_11952);
nand U12586 (N_12586,N_11583,N_10136);
and U12587 (N_12587,N_10328,N_11163);
nand U12588 (N_12588,N_11856,N_10562);
nor U12589 (N_12589,N_11325,N_9472);
xor U12590 (N_12590,N_10318,N_10585);
nor U12591 (N_12591,N_10286,N_11157);
or U12592 (N_12592,N_11834,N_9132);
nand U12593 (N_12593,N_11601,N_10178);
nor U12594 (N_12594,N_11255,N_11967);
and U12595 (N_12595,N_11133,N_9134);
and U12596 (N_12596,N_10044,N_11477);
and U12597 (N_12597,N_9143,N_9000);
and U12598 (N_12598,N_9895,N_11633);
nand U12599 (N_12599,N_11817,N_10408);
and U12600 (N_12600,N_11648,N_10800);
nand U12601 (N_12601,N_9860,N_10901);
nor U12602 (N_12602,N_10287,N_9994);
nand U12603 (N_12603,N_11719,N_9418);
nand U12604 (N_12604,N_9965,N_10498);
nor U12605 (N_12605,N_10390,N_9592);
or U12606 (N_12606,N_11370,N_11205);
or U12607 (N_12607,N_11638,N_9259);
nor U12608 (N_12608,N_11689,N_9029);
and U12609 (N_12609,N_10488,N_9594);
and U12610 (N_12610,N_11544,N_11909);
or U12611 (N_12611,N_11145,N_10544);
or U12612 (N_12612,N_9710,N_10012);
and U12613 (N_12613,N_11415,N_11158);
or U12614 (N_12614,N_9964,N_11281);
or U12615 (N_12615,N_9556,N_9686);
nand U12616 (N_12616,N_11285,N_11478);
nand U12617 (N_12617,N_9104,N_10791);
or U12618 (N_12618,N_11835,N_11321);
nor U12619 (N_12619,N_9706,N_10844);
or U12620 (N_12620,N_10728,N_11086);
and U12621 (N_12621,N_10716,N_9275);
xnor U12622 (N_12622,N_10548,N_9899);
and U12623 (N_12623,N_9184,N_10221);
and U12624 (N_12624,N_11877,N_11825);
nand U12625 (N_12625,N_11007,N_11968);
or U12626 (N_12626,N_11963,N_10280);
nor U12627 (N_12627,N_9524,N_9121);
xnor U12628 (N_12628,N_11753,N_9885);
and U12629 (N_12629,N_9042,N_10810);
nand U12630 (N_12630,N_11693,N_10141);
or U12631 (N_12631,N_11902,N_11291);
or U12632 (N_12632,N_9601,N_9839);
or U12633 (N_12633,N_10741,N_10001);
and U12634 (N_12634,N_9859,N_10619);
nand U12635 (N_12635,N_11898,N_9590);
and U12636 (N_12636,N_9236,N_10003);
and U12637 (N_12637,N_10678,N_9892);
nand U12638 (N_12638,N_11045,N_11369);
or U12639 (N_12639,N_10586,N_10647);
and U12640 (N_12640,N_11557,N_10265);
and U12641 (N_12641,N_11860,N_9314);
nand U12642 (N_12642,N_11636,N_10016);
and U12643 (N_12643,N_9167,N_11413);
nand U12644 (N_12644,N_10992,N_9009);
or U12645 (N_12645,N_11703,N_10690);
nor U12646 (N_12646,N_10608,N_11748);
nor U12647 (N_12647,N_9959,N_10249);
nor U12648 (N_12648,N_9593,N_11228);
nor U12649 (N_12649,N_10183,N_11927);
nor U12650 (N_12650,N_10004,N_10131);
or U12651 (N_12651,N_10167,N_10913);
nand U12652 (N_12652,N_11782,N_10592);
and U12653 (N_12653,N_11580,N_11483);
or U12654 (N_12654,N_11367,N_10674);
and U12655 (N_12655,N_9652,N_9855);
nand U12656 (N_12656,N_11444,N_11372);
nor U12657 (N_12657,N_9570,N_10872);
and U12658 (N_12658,N_9193,N_10023);
nand U12659 (N_12659,N_9152,N_11479);
and U12660 (N_12660,N_9107,N_11535);
or U12661 (N_12661,N_9321,N_10715);
or U12662 (N_12662,N_10905,N_9225);
nand U12663 (N_12663,N_10926,N_11093);
and U12664 (N_12664,N_9467,N_11491);
nand U12665 (N_12665,N_10774,N_9604);
or U12666 (N_12666,N_11961,N_10365);
and U12667 (N_12667,N_11936,N_10822);
and U12668 (N_12668,N_9765,N_11195);
and U12669 (N_12669,N_9631,N_9394);
xor U12670 (N_12670,N_10637,N_9729);
nand U12671 (N_12671,N_11143,N_11222);
or U12672 (N_12672,N_10179,N_11873);
nor U12673 (N_12673,N_10736,N_10396);
nor U12674 (N_12674,N_10437,N_11658);
nand U12675 (N_12675,N_9730,N_11050);
nand U12676 (N_12676,N_11246,N_10606);
nand U12677 (N_12677,N_9041,N_11379);
or U12678 (N_12678,N_9212,N_11032);
and U12679 (N_12679,N_10282,N_9142);
nor U12680 (N_12680,N_11505,N_11900);
or U12681 (N_12681,N_10092,N_11463);
nor U12682 (N_12682,N_11115,N_10311);
nor U12683 (N_12683,N_10224,N_9925);
nor U12684 (N_12684,N_9963,N_10306);
or U12685 (N_12685,N_11456,N_10958);
nor U12686 (N_12686,N_11941,N_11116);
and U12687 (N_12687,N_11973,N_11113);
or U12688 (N_12688,N_10144,N_10151);
nor U12689 (N_12689,N_10463,N_10726);
nand U12690 (N_12690,N_11320,N_9531);
nor U12691 (N_12691,N_9880,N_10602);
and U12692 (N_12692,N_11226,N_11315);
and U12693 (N_12693,N_9572,N_9533);
or U12694 (N_12694,N_10439,N_11083);
or U12695 (N_12695,N_9488,N_10877);
nand U12696 (N_12696,N_10205,N_11773);
or U12697 (N_12697,N_10587,N_10673);
nand U12698 (N_12698,N_9487,N_11830);
nor U12699 (N_12699,N_9529,N_9079);
nand U12700 (N_12700,N_10852,N_9508);
nor U12701 (N_12701,N_9431,N_11686);
or U12702 (N_12702,N_10079,N_11346);
and U12703 (N_12703,N_10622,N_9973);
nand U12704 (N_12704,N_9117,N_10052);
or U12705 (N_12705,N_10432,N_10115);
nand U12706 (N_12706,N_10557,N_10777);
or U12707 (N_12707,N_9550,N_11684);
or U12708 (N_12708,N_9425,N_11894);
or U12709 (N_12709,N_9544,N_11196);
nor U12710 (N_12710,N_9976,N_11937);
and U12711 (N_12711,N_10729,N_9437);
nand U12712 (N_12712,N_10030,N_11381);
or U12713 (N_12713,N_11339,N_11194);
or U12714 (N_12714,N_10008,N_9473);
nand U12715 (N_12715,N_11160,N_9070);
nor U12716 (N_12716,N_9479,N_11639);
and U12717 (N_12717,N_11144,N_11611);
and U12718 (N_12718,N_10723,N_11230);
nor U12719 (N_12719,N_11480,N_11248);
nor U12720 (N_12720,N_11517,N_9241);
and U12721 (N_12721,N_9158,N_11302);
nor U12722 (N_12722,N_9719,N_10882);
and U12723 (N_12723,N_10036,N_11536);
nor U12724 (N_12724,N_9396,N_9153);
nand U12725 (N_12725,N_11627,N_9244);
nor U12726 (N_12726,N_10308,N_10670);
nand U12727 (N_12727,N_11520,N_11219);
or U12728 (N_12728,N_11235,N_10952);
nand U12729 (N_12729,N_11735,N_9386);
and U12730 (N_12730,N_9499,N_9615);
and U12731 (N_12731,N_10824,N_9415);
and U12732 (N_12732,N_11387,N_10783);
nand U12733 (N_12733,N_11249,N_9312);
nand U12734 (N_12734,N_9879,N_10627);
nor U12735 (N_12735,N_9690,N_10604);
nand U12736 (N_12736,N_9392,N_10168);
and U12737 (N_12737,N_10931,N_11106);
nor U12738 (N_12738,N_10540,N_9937);
xnor U12739 (N_12739,N_9209,N_11436);
and U12740 (N_12740,N_9206,N_10350);
or U12741 (N_12741,N_11928,N_9562);
nor U12742 (N_12742,N_11697,N_11019);
nor U12743 (N_12743,N_11953,N_9197);
or U12744 (N_12744,N_10692,N_10904);
nand U12745 (N_12745,N_11768,N_10402);
nand U12746 (N_12746,N_11530,N_9649);
and U12747 (N_12747,N_9723,N_11065);
and U12748 (N_12748,N_9336,N_10440);
nand U12749 (N_12749,N_9712,N_11449);
or U12750 (N_12750,N_9715,N_9567);
nor U12751 (N_12751,N_10501,N_9688);
nand U12752 (N_12752,N_9318,N_11077);
nand U12753 (N_12753,N_11687,N_10292);
or U12754 (N_12754,N_10770,N_10383);
or U12755 (N_12755,N_11714,N_11951);
or U12756 (N_12756,N_10029,N_9391);
or U12757 (N_12757,N_10588,N_10093);
nor U12758 (N_12758,N_10118,N_10199);
or U12759 (N_12759,N_11138,N_9953);
or U12760 (N_12760,N_9133,N_10312);
or U12761 (N_12761,N_11840,N_9872);
or U12762 (N_12762,N_11956,N_9863);
nor U12763 (N_12763,N_10635,N_9836);
or U12764 (N_12764,N_10693,N_10417);
or U12765 (N_12765,N_10011,N_11623);
and U12766 (N_12766,N_9339,N_9558);
nor U12767 (N_12767,N_10642,N_9404);
and U12768 (N_12768,N_9125,N_9517);
nor U12769 (N_12769,N_9514,N_11813);
nand U12770 (N_12770,N_11677,N_10561);
nor U12771 (N_12771,N_11723,N_10583);
and U12772 (N_12772,N_11089,N_9131);
and U12773 (N_12773,N_10514,N_9355);
nand U12774 (N_12774,N_11009,N_10380);
nand U12775 (N_12775,N_11234,N_11637);
or U12776 (N_12776,N_10262,N_11203);
and U12777 (N_12777,N_10704,N_11462);
nor U12778 (N_12778,N_10181,N_9238);
or U12779 (N_12779,N_10614,N_9324);
nor U12780 (N_12780,N_11984,N_11441);
or U12781 (N_12781,N_10589,N_11335);
nand U12782 (N_12782,N_11899,N_11948);
and U12783 (N_12783,N_11393,N_9254);
nand U12784 (N_12784,N_10241,N_10462);
nand U12785 (N_12785,N_9655,N_9584);
nand U12786 (N_12786,N_9400,N_10577);
nor U12787 (N_12787,N_10406,N_10839);
and U12788 (N_12788,N_11445,N_10494);
or U12789 (N_12789,N_9632,N_11785);
nand U12790 (N_12790,N_11090,N_9671);
or U12791 (N_12791,N_9917,N_9694);
and U12792 (N_12792,N_10620,N_11024);
nand U12793 (N_12793,N_9297,N_9045);
nor U12794 (N_12794,N_9676,N_10076);
nor U12795 (N_12795,N_10346,N_11757);
or U12796 (N_12796,N_10296,N_11271);
nor U12797 (N_12797,N_9423,N_9692);
and U12798 (N_12798,N_9419,N_9361);
or U12799 (N_12799,N_9519,N_10113);
nor U12800 (N_12800,N_10127,N_11645);
or U12801 (N_12801,N_11274,N_10682);
and U12802 (N_12802,N_9183,N_10547);
nor U12803 (N_12803,N_9229,N_9758);
or U12804 (N_12804,N_9618,N_10275);
and U12805 (N_12805,N_11001,N_9128);
nand U12806 (N_12806,N_9657,N_9030);
nand U12807 (N_12807,N_11202,N_11998);
and U12808 (N_12808,N_10103,N_10204);
nand U12809 (N_12809,N_9376,N_10572);
and U12810 (N_12810,N_10017,N_10424);
or U12811 (N_12811,N_9215,N_9947);
or U12812 (N_12812,N_9300,N_11622);
and U12813 (N_12813,N_9984,N_10578);
and U12814 (N_12814,N_11390,N_10260);
nor U12815 (N_12815,N_11957,N_9182);
and U12816 (N_12816,N_10334,N_9370);
or U12817 (N_12817,N_10165,N_11244);
xor U12818 (N_12818,N_9383,N_9141);
nor U12819 (N_12819,N_11337,N_11947);
nand U12820 (N_12820,N_10344,N_11419);
and U12821 (N_12821,N_10200,N_10242);
and U12822 (N_12822,N_11391,N_10761);
nor U12823 (N_12823,N_11733,N_10499);
and U12824 (N_12824,N_10376,N_9609);
nand U12825 (N_12825,N_9194,N_9025);
and U12826 (N_12826,N_10230,N_11745);
nand U12827 (N_12827,N_9862,N_10569);
nand U12828 (N_12828,N_9334,N_10368);
nor U12829 (N_12829,N_9222,N_10198);
or U12830 (N_12830,N_9234,N_11698);
or U12831 (N_12831,N_9736,N_11342);
nand U12832 (N_12832,N_11099,N_9054);
nand U12833 (N_12833,N_10838,N_9352);
nand U12834 (N_12834,N_11501,N_10972);
and U12835 (N_12835,N_11149,N_10117);
nor U12836 (N_12836,N_10164,N_10828);
nand U12837 (N_12837,N_11908,N_11942);
nand U12838 (N_12838,N_11592,N_9344);
or U12839 (N_12839,N_9372,N_11300);
and U12840 (N_12840,N_10269,N_9168);
or U12841 (N_12841,N_11718,N_10826);
nand U12842 (N_12842,N_9490,N_10681);
nor U12843 (N_12843,N_10917,N_10244);
nand U12844 (N_12844,N_9039,N_9161);
or U12845 (N_12845,N_11796,N_9247);
nand U12846 (N_12846,N_10210,N_9582);
nand U12847 (N_12847,N_11539,N_9557);
nand U12848 (N_12848,N_9110,N_9647);
xor U12849 (N_12849,N_9203,N_10229);
and U12850 (N_12850,N_11850,N_10734);
nand U12851 (N_12851,N_10841,N_11486);
nand U12852 (N_12852,N_10849,N_9970);
nor U12853 (N_12853,N_10563,N_10717);
nor U12854 (N_12854,N_10605,N_11069);
nand U12855 (N_12855,N_11559,N_9163);
and U12856 (N_12856,N_10111,N_10581);
xnor U12857 (N_12857,N_9439,N_10694);
nand U12858 (N_12858,N_10648,N_11229);
or U12859 (N_12859,N_9936,N_10987);
or U12860 (N_12860,N_9914,N_9335);
nor U12861 (N_12861,N_9578,N_9898);
nor U12862 (N_12862,N_9512,N_11482);
nor U12863 (N_12863,N_9416,N_9771);
nand U12864 (N_12864,N_11108,N_9798);
nor U12865 (N_12865,N_9062,N_11023);
nand U12866 (N_12866,N_10191,N_10792);
nand U12867 (N_12867,N_10458,N_10483);
nand U12868 (N_12868,N_11147,N_11586);
or U12869 (N_12869,N_9239,N_9792);
and U12870 (N_12870,N_11632,N_9705);
and U12871 (N_12871,N_10225,N_10744);
or U12872 (N_12872,N_10937,N_9465);
nand U12873 (N_12873,N_11411,N_11284);
and U12874 (N_12874,N_10218,N_11152);
or U12875 (N_12875,N_11156,N_11897);
nor U12876 (N_12876,N_9356,N_10710);
or U12877 (N_12877,N_11944,N_11176);
nand U12878 (N_12878,N_10978,N_10372);
nor U12879 (N_12879,N_9481,N_10703);
or U12880 (N_12880,N_9977,N_9574);
and U12881 (N_12881,N_10134,N_11423);
nand U12882 (N_12882,N_9669,N_11504);
or U12883 (N_12883,N_11766,N_11102);
or U12884 (N_12884,N_11410,N_11207);
or U12885 (N_12885,N_11118,N_10556);
or U12886 (N_12886,N_11867,N_10924);
nand U12887 (N_12887,N_9919,N_9788);
nand U12888 (N_12888,N_11260,N_9310);
or U12889 (N_12889,N_9634,N_10549);
and U12890 (N_12890,N_9924,N_11182);
or U12891 (N_12891,N_10461,N_10256);
nor U12892 (N_12892,N_10392,N_11507);
and U12893 (N_12893,N_10473,N_10621);
xnor U12894 (N_12894,N_9001,N_9526);
or U12895 (N_12895,N_10543,N_10156);
nand U12896 (N_12896,N_11414,N_9202);
and U12897 (N_12897,N_11660,N_10700);
nand U12898 (N_12898,N_9449,N_9627);
and U12899 (N_12899,N_9796,N_10598);
nor U12900 (N_12900,N_10051,N_9457);
or U12901 (N_12901,N_11884,N_11610);
nor U12902 (N_12902,N_11549,N_9691);
or U12903 (N_12903,N_10857,N_11761);
or U12904 (N_12904,N_11654,N_11110);
nand U12905 (N_12905,N_9385,N_10759);
and U12906 (N_12906,N_11603,N_9460);
nand U12907 (N_12907,N_10276,N_9834);
nand U12908 (N_12908,N_10222,N_9443);
or U12909 (N_12909,N_11469,N_9891);
or U12910 (N_12910,N_9309,N_10922);
nand U12911 (N_12911,N_10646,N_11776);
and U12912 (N_12912,N_10508,N_10125);
or U12913 (N_12913,N_9205,N_10506);
nor U12914 (N_12914,N_10129,N_9040);
and U12915 (N_12915,N_9698,N_9904);
nand U12916 (N_12916,N_9089,N_11615);
and U12917 (N_12917,N_9341,N_9660);
and U12918 (N_12918,N_10485,N_11576);
xor U12919 (N_12919,N_9369,N_10632);
nor U12920 (N_12920,N_10871,N_11887);
and U12921 (N_12921,N_10530,N_10503);
nor U12922 (N_12922,N_10139,N_9359);
and U12923 (N_12923,N_11079,N_9050);
or U12924 (N_12924,N_9434,N_9726);
nand U12925 (N_12925,N_10816,N_9366);
nand U12926 (N_12926,N_11293,N_11814);
nor U12927 (N_12927,N_9776,N_9265);
or U12928 (N_12928,N_9878,N_10956);
and U12929 (N_12929,N_9284,N_10253);
and U12930 (N_12930,N_10529,N_11063);
xnor U12931 (N_12931,N_11438,N_10985);
and U12932 (N_12932,N_11437,N_9088);
nor U12933 (N_12933,N_10313,N_10712);
nor U12934 (N_12934,N_9799,N_9413);
nor U12935 (N_12935,N_9379,N_10532);
or U12936 (N_12936,N_10916,N_11422);
and U12937 (N_12937,N_9458,N_11111);
or U12938 (N_12938,N_10459,N_10177);
and U12939 (N_12939,N_11015,N_10444);
nand U12940 (N_12940,N_11624,N_11453);
and U12941 (N_12941,N_9461,N_10963);
and U12942 (N_12942,N_10517,N_10624);
nand U12943 (N_12943,N_11604,N_9901);
nor U12944 (N_12944,N_11177,N_9177);
nor U12945 (N_12945,N_9540,N_9797);
and U12946 (N_12946,N_9689,N_11734);
nor U12947 (N_12947,N_11537,N_9068);
and U12948 (N_12948,N_9731,N_9277);
or U12949 (N_12949,N_10803,N_11091);
nand U12950 (N_12950,N_10616,N_10387);
or U12951 (N_12951,N_10028,N_9952);
nor U12952 (N_12952,N_11556,N_11383);
nand U12953 (N_12953,N_10998,N_10239);
and U12954 (N_12954,N_9420,N_10497);
or U12955 (N_12955,N_9139,N_9950);
nor U12956 (N_12956,N_9656,N_10831);
nor U12957 (N_12957,N_11533,N_11842);
nand U12958 (N_12958,N_10671,N_10745);
nand U12959 (N_12959,N_10625,N_10393);
or U12960 (N_12960,N_11625,N_10932);
and U12961 (N_12961,N_9668,N_9847);
nor U12962 (N_12962,N_10464,N_10343);
and U12963 (N_12963,N_10584,N_9532);
and U12964 (N_12964,N_11427,N_9082);
nor U12965 (N_12965,N_11052,N_9995);
nor U12966 (N_12966,N_11778,N_10072);
or U12967 (N_12967,N_11564,N_9057);
or U12968 (N_12968,N_10983,N_9242);
and U12969 (N_12969,N_10697,N_11891);
nand U12970 (N_12970,N_10467,N_10469);
and U12971 (N_12971,N_11710,N_9170);
or U12972 (N_12972,N_10348,N_9260);
and U12973 (N_12973,N_10309,N_11546);
and U12974 (N_12974,N_10366,N_10929);
nand U12975 (N_12975,N_9733,N_11804);
and U12976 (N_12976,N_11500,N_10787);
nor U12977 (N_12977,N_9673,N_9279);
nand U12978 (N_12978,N_11990,N_9303);
nor U12979 (N_12979,N_9856,N_11652);
or U12980 (N_12980,N_10784,N_10429);
nor U12981 (N_12981,N_11617,N_10768);
nand U12982 (N_12982,N_9747,N_11848);
nand U12983 (N_12983,N_11752,N_10628);
nor U12984 (N_12984,N_10618,N_11798);
and U12985 (N_12985,N_9410,N_10537);
and U12986 (N_12986,N_9078,N_11141);
nor U12987 (N_12987,N_10976,N_11919);
nand U12988 (N_12988,N_11545,N_10748);
and U12989 (N_12989,N_11749,N_9749);
nand U12990 (N_12990,N_9325,N_11979);
nor U12991 (N_12991,N_9580,N_11502);
and U12992 (N_12992,N_11696,N_9118);
or U12993 (N_12993,N_10048,N_11016);
and U12994 (N_12994,N_10083,N_9174);
nand U12995 (N_12995,N_9527,N_9218);
or U12996 (N_12996,N_9721,N_10245);
nor U12997 (N_12997,N_11148,N_11716);
and U12998 (N_12998,N_9055,N_10474);
or U12999 (N_12999,N_11408,N_10991);
and U13000 (N_13000,N_10482,N_9809);
and U13001 (N_13001,N_9746,N_11861);
nand U13002 (N_13002,N_11294,N_11010);
or U13003 (N_13003,N_11989,N_11028);
nand U13004 (N_13004,N_11428,N_9483);
nor U13005 (N_13005,N_11905,N_10940);
and U13006 (N_13006,N_9034,N_10836);
nor U13007 (N_13007,N_10500,N_10965);
nand U13008 (N_13008,N_9814,N_9756);
or U13009 (N_13009,N_10182,N_11857);
and U13010 (N_13010,N_10927,N_11811);
nand U13011 (N_13011,N_11895,N_9365);
or U13012 (N_13012,N_10137,N_10338);
nand U13013 (N_13013,N_9824,N_11712);
nor U13014 (N_13014,N_10754,N_9662);
and U13015 (N_13015,N_11819,N_9027);
and U13016 (N_13016,N_9178,N_9785);
nor U13017 (N_13017,N_9700,N_10484);
xnor U13018 (N_13018,N_9252,N_9323);
nand U13019 (N_13019,N_9243,N_11087);
or U13020 (N_13020,N_10655,N_10925);
or U13021 (N_13021,N_9498,N_9802);
nor U13022 (N_13022,N_11588,N_11810);
nor U13023 (N_13023,N_9116,N_9699);
nand U13024 (N_13024,N_11155,N_10812);
nand U13025 (N_13025,N_9735,N_11259);
nand U13026 (N_13026,N_10333,N_11643);
nor U13027 (N_13027,N_11193,N_9566);
nor U13028 (N_13028,N_10948,N_11033);
and U13029 (N_13029,N_10059,N_10138);
or U13030 (N_13030,N_9308,N_10743);
nand U13031 (N_13031,N_10653,N_11715);
nand U13032 (N_13032,N_10993,N_11680);
nand U13033 (N_13033,N_11669,N_11251);
or U13034 (N_13034,N_10238,N_9966);
nor U13035 (N_13035,N_11403,N_11971);
nand U13036 (N_13036,N_11475,N_11730);
nor U13037 (N_13037,N_9515,N_9256);
nor U13038 (N_13038,N_11981,N_11892);
nor U13039 (N_13039,N_9342,N_10426);
nor U13040 (N_13040,N_11646,N_9942);
nand U13041 (N_13041,N_10610,N_10214);
nand U13042 (N_13042,N_9051,N_11599);
nor U13043 (N_13043,N_11721,N_11931);
nor U13044 (N_13044,N_10921,N_9406);
and U13045 (N_13045,N_11472,N_9444);
and U13046 (N_13046,N_11097,N_9071);
and U13047 (N_13047,N_10971,N_11651);
and U13048 (N_13048,N_9523,N_9393);
or U13049 (N_13049,N_9261,N_9980);
nand U13050 (N_13050,N_10718,N_9653);
or U13051 (N_13051,N_9002,N_10567);
nor U13052 (N_13052,N_9522,N_9720);
nor U13053 (N_13053,N_10428,N_11258);
nor U13054 (N_13054,N_11026,N_11237);
xor U13055 (N_13055,N_10040,N_9587);
and U13056 (N_13056,N_10252,N_9289);
nor U13057 (N_13057,N_9849,N_11705);
nand U13058 (N_13058,N_9463,N_11484);
or U13059 (N_13059,N_11653,N_9620);
or U13060 (N_13060,N_9577,N_9005);
nor U13061 (N_13061,N_11166,N_9470);
or U13062 (N_13062,N_9511,N_9250);
nand U13063 (N_13063,N_10798,N_9713);
nor U13064 (N_13064,N_11142,N_10698);
or U13065 (N_13065,N_10861,N_11442);
nor U13066 (N_13066,N_9999,N_11343);
and U13067 (N_13067,N_11675,N_9598);
and U13068 (N_13068,N_10298,N_9724);
nor U13069 (N_13069,N_11701,N_11282);
and U13070 (N_13070,N_11913,N_11060);
nand U13071 (N_13071,N_9828,N_10186);
and U13072 (N_13072,N_10213,N_10071);
and U13073 (N_13073,N_10358,N_11955);
or U13074 (N_13074,N_10846,N_11915);
nand U13075 (N_13075,N_9126,N_10753);
and U13076 (N_13076,N_9253,N_9915);
and U13077 (N_13077,N_11225,N_9605);
nand U13078 (N_13078,N_10636,N_10010);
nor U13079 (N_13079,N_10973,N_11455);
nand U13080 (N_13080,N_10270,N_10243);
nand U13081 (N_13081,N_9115,N_11950);
nor U13082 (N_13082,N_10659,N_9910);
nand U13083 (N_13083,N_9122,N_11945);
nor U13084 (N_13084,N_10654,N_11506);
nand U13085 (N_13085,N_11969,N_11903);
and U13086 (N_13086,N_11057,N_9768);
or U13087 (N_13087,N_10405,N_10859);
and U13088 (N_13088,N_9646,N_9826);
nor U13089 (N_13089,N_11460,N_10223);
and U13090 (N_13090,N_10510,N_9144);
and U13091 (N_13091,N_10015,N_11088);
and U13092 (N_13092,N_11197,N_10896);
or U13093 (N_13093,N_11353,N_10579);
xnor U13094 (N_13094,N_10410,N_11317);
and U13095 (N_13095,N_10027,N_10336);
or U13096 (N_13096,N_9060,N_10031);
and U13097 (N_13097,N_9306,N_10806);
or U13098 (N_13098,N_9547,N_9417);
and U13099 (N_13099,N_10660,N_11934);
or U13100 (N_13100,N_10108,N_11209);
nand U13101 (N_13101,N_10442,N_9852);
nor U13102 (N_13102,N_11253,N_9777);
nand U13103 (N_13103,N_10505,N_9993);
or U13104 (N_13104,N_9166,N_11130);
nor U13105 (N_13105,N_9742,N_10727);
nor U13106 (N_13106,N_11924,N_9599);
nand U13107 (N_13107,N_10112,N_9357);
and U13108 (N_13108,N_9214,N_9677);
and U13109 (N_13109,N_11254,N_10657);
nand U13110 (N_13110,N_10623,N_9873);
nor U13111 (N_13111,N_11062,N_10236);
or U13112 (N_13112,N_10273,N_11356);
nor U13113 (N_13113,N_9149,N_11265);
nor U13114 (N_13114,N_9934,N_11525);
nand U13115 (N_13115,N_9095,N_10385);
or U13116 (N_13116,N_9793,N_9981);
nor U13117 (N_13117,N_9270,N_9876);
and U13118 (N_13118,N_11364,N_9338);
and U13119 (N_13119,N_11831,N_10299);
and U13120 (N_13120,N_10394,N_9480);
nand U13121 (N_13121,N_9440,N_11598);
nor U13122 (N_13122,N_11120,N_9255);
nor U13123 (N_13123,N_11073,N_9200);
nand U13124 (N_13124,N_9048,N_11000);
or U13125 (N_13125,N_11355,N_9171);
or U13126 (N_13126,N_11425,N_10219);
nor U13127 (N_13127,N_9579,N_10611);
and U13128 (N_13128,N_9961,N_10316);
nand U13129 (N_13129,N_9084,N_11800);
or U13130 (N_13130,N_11508,N_11017);
nor U13131 (N_13131,N_9875,N_11365);
nor U13132 (N_13132,N_10560,N_10133);
or U13133 (N_13133,N_9912,N_11596);
or U13134 (N_13134,N_9422,N_10068);
nand U13135 (N_13135,N_11450,N_9452);
and U13136 (N_13136,N_9816,N_11512);
or U13137 (N_13137,N_11770,N_9635);
nand U13138 (N_13138,N_10667,N_11641);
nor U13139 (N_13139,N_9278,N_10025);
nor U13140 (N_13140,N_11191,N_10856);
or U13141 (N_13141,N_9670,N_9740);
nand U13142 (N_13142,N_11498,N_10789);
nor U13143 (N_13143,N_10037,N_11590);
nand U13144 (N_13144,N_11125,N_11932);
and U13145 (N_13145,N_11614,N_9233);
nor U13146 (N_13146,N_11975,N_9004);
or U13147 (N_13147,N_10477,N_10490);
or U13148 (N_13148,N_11843,N_10599);
and U13149 (N_13149,N_9075,N_11267);
and U13150 (N_13150,N_10317,N_9795);
or U13151 (N_13151,N_10780,N_11447);
nor U13152 (N_13152,N_11818,N_9779);
and U13153 (N_13153,N_10170,N_10277);
nand U13154 (N_13154,N_10990,N_10531);
nor U13155 (N_13155,N_10207,N_9468);
nand U13156 (N_13156,N_11105,N_9033);
or U13157 (N_13157,N_9946,N_10892);
nand U13158 (N_13158,N_9482,N_10261);
and U13159 (N_13159,N_11943,N_11750);
nor U13160 (N_13160,N_9787,N_10110);
nand U13161 (N_13161,N_9345,N_9492);
nor U13162 (N_13162,N_9287,N_10067);
nand U13163 (N_13163,N_9219,N_10795);
and U13164 (N_13164,N_9061,N_9014);
nand U13165 (N_13165,N_10809,N_11920);
and U13166 (N_13166,N_10900,N_11051);
nand U13167 (N_13167,N_11558,N_9968);
nor U13168 (N_13168,N_10171,N_11132);
nand U13169 (N_13169,N_9304,N_10574);
nand U13170 (N_13170,N_9228,N_10974);
nand U13171 (N_13171,N_10293,N_9685);
and U13172 (N_13172,N_9402,N_10295);
or U13173 (N_13173,N_10492,N_11870);
nand U13174 (N_13174,N_9390,N_9864);
or U13175 (N_13175,N_9600,N_11487);
or U13176 (N_13176,N_10778,N_11137);
or U13177 (N_13177,N_11591,N_10082);
or U13178 (N_13178,N_11164,N_10465);
nand U13179 (N_13179,N_11812,N_9909);
nor U13180 (N_13180,N_9148,N_11066);
or U13181 (N_13181,N_10977,N_9150);
or U13182 (N_13182,N_9728,N_11288);
nand U13183 (N_13183,N_10834,N_9848);
and U13184 (N_13184,N_9192,N_10893);
and U13185 (N_13185,N_9613,N_10105);
nor U13186 (N_13186,N_9845,N_9933);
and U13187 (N_13187,N_9808,N_11264);
or U13188 (N_13188,N_9293,N_11829);
nand U13189 (N_13189,N_9282,N_11741);
and U13190 (N_13190,N_11777,N_9882);
or U13191 (N_13191,N_10821,N_10696);
nor U13192 (N_13192,N_11702,N_11104);
nand U13193 (N_13193,N_10160,N_10945);
or U13194 (N_13194,N_10053,N_11972);
and U13195 (N_13195,N_9347,N_10823);
nand U13196 (N_13196,N_9160,N_9835);
nor U13197 (N_13197,N_9806,N_9290);
nor U13198 (N_13198,N_9717,N_10840);
or U13199 (N_13199,N_11098,N_11529);
and U13200 (N_13200,N_11011,N_9364);
or U13201 (N_13201,N_9435,N_10594);
or U13202 (N_13202,N_9564,N_11454);
or U13203 (N_13203,N_9497,N_9974);
nand U13204 (N_13204,N_10573,N_10769);
nor U13205 (N_13205,N_10388,N_10135);
and U13206 (N_13206,N_9227,N_9081);
nor U13207 (N_13207,N_9530,N_10546);
and U13208 (N_13208,N_11958,N_11183);
or U13209 (N_13209,N_9546,N_10850);
nand U13210 (N_13210,N_10162,N_10833);
or U13211 (N_13211,N_11340,N_11338);
nand U13212 (N_13212,N_9340,N_11311);
nand U13213 (N_13213,N_11495,N_11863);
nand U13214 (N_13214,N_11273,N_11333);
nand U13215 (N_13215,N_11466,N_9820);
xor U13216 (N_13216,N_9903,N_9007);
or U13217 (N_13217,N_11738,N_10613);
or U13218 (N_13218,N_9513,N_10294);
or U13219 (N_13219,N_10322,N_11322);
or U13220 (N_13220,N_10897,N_11341);
nor U13221 (N_13221,N_9389,N_10024);
or U13222 (N_13222,N_9725,N_10788);
and U13223 (N_13223,N_9195,N_10104);
nor U13224 (N_13224,N_11672,N_9543);
nand U13225 (N_13225,N_9438,N_9106);
and U13226 (N_13226,N_9949,N_11167);
nand U13227 (N_13227,N_11526,N_10355);
nand U13228 (N_13228,N_11821,N_9643);
or U13229 (N_13229,N_11562,N_11129);
nand U13230 (N_13230,N_9291,N_10374);
nand U13231 (N_13231,N_9573,N_11021);
or U13232 (N_13232,N_9327,N_10535);
nor U13233 (N_13233,N_11875,N_10443);
and U13234 (N_13234,N_10580,N_9058);
or U13235 (N_13235,N_11889,N_10121);
or U13236 (N_13236,N_11740,N_11080);
nor U13237 (N_13237,N_9773,N_9817);
and U13238 (N_13238,N_11220,N_11362);
or U13239 (N_13239,N_11926,N_11921);
or U13240 (N_13240,N_9811,N_10257);
or U13241 (N_13241,N_11095,N_10708);
nand U13242 (N_13242,N_9451,N_11309);
nand U13243 (N_13243,N_9941,N_9003);
nor U13244 (N_13244,N_9541,N_11459);
or U13245 (N_13245,N_11914,N_10401);
nor U13246 (N_13246,N_11859,N_11323);
nand U13247 (N_13247,N_10629,N_10997);
and U13248 (N_13248,N_11844,N_9162);
nor U13249 (N_13249,N_9330,N_9382);
nor U13250 (N_13250,N_10607,N_9575);
nand U13251 (N_13251,N_9274,N_9285);
nor U13252 (N_13252,N_9624,N_11168);
or U13253 (N_13253,N_11547,N_10176);
and U13254 (N_13254,N_9987,N_10190);
nor U13255 (N_13255,N_10830,N_9456);
nand U13256 (N_13256,N_10724,N_9752);
or U13257 (N_13257,N_11276,N_10454);
or U13258 (N_13258,N_10936,N_11416);
or U13259 (N_13259,N_11765,N_11630);
xnor U13260 (N_13260,N_10942,N_11820);
nand U13261 (N_13261,N_11473,N_9850);
or U13262 (N_13262,N_9960,N_10709);
or U13263 (N_13263,N_9097,N_9464);
nand U13264 (N_13264,N_10644,N_9663);
nor U13265 (N_13265,N_11022,N_9926);
and U13266 (N_13266,N_11978,N_9494);
nand U13267 (N_13267,N_10766,N_9595);
and U13268 (N_13268,N_10666,N_10084);
and U13269 (N_13269,N_11678,N_10124);
and U13270 (N_13270,N_10612,N_11270);
and U13271 (N_13271,N_11855,N_11174);
and U13272 (N_13272,N_11211,N_11232);
nor U13273 (N_13273,N_10247,N_9654);
nor U13274 (N_13274,N_10848,N_9754);
and U13275 (N_13275,N_11306,N_9822);
nand U13276 (N_13276,N_11574,N_11524);
nor U13277 (N_13277,N_11904,N_11384);
xnor U13278 (N_13278,N_10796,N_11452);
and U13279 (N_13279,N_10425,N_11146);
nand U13280 (N_13280,N_11290,N_9428);
nor U13281 (N_13281,N_10553,N_11579);
nor U13282 (N_13282,N_9056,N_9022);
or U13283 (N_13283,N_11382,N_11642);
or U13284 (N_13284,N_10781,N_9448);
nor U13285 (N_13285,N_9414,N_10771);
nand U13286 (N_13286,N_10166,N_10898);
and U13287 (N_13287,N_9877,N_9928);
or U13288 (N_13288,N_10656,N_9320);
nor U13289 (N_13289,N_9495,N_9607);
nand U13290 (N_13290,N_11706,N_11070);
nand U13291 (N_13291,N_11871,N_9135);
nand U13292 (N_13292,N_11694,N_10020);
or U13293 (N_13293,N_11569,N_10307);
nor U13294 (N_13294,N_10174,N_9453);
nor U13295 (N_13295,N_9800,N_9179);
or U13296 (N_13296,N_10749,N_10447);
nor U13297 (N_13297,N_10361,N_9887);
and U13298 (N_13298,N_9520,N_9930);
nand U13299 (N_13299,N_9221,N_10786);
nor U13300 (N_13300,N_10153,N_9633);
xnor U13301 (N_13301,N_11966,N_9638);
or U13302 (N_13302,N_9971,N_11774);
and U13303 (N_13303,N_9489,N_11851);
and U13304 (N_13304,N_11515,N_9958);
nor U13305 (N_13305,N_10073,N_9586);
nor U13306 (N_13306,N_11649,N_11607);
nand U13307 (N_13307,N_9245,N_11361);
and U13308 (N_13308,N_9896,N_10430);
or U13309 (N_13309,N_9832,N_9147);
and U13310 (N_13310,N_9373,N_9264);
nand U13311 (N_13311,N_10324,N_11162);
nand U13312 (N_13312,N_11151,N_11685);
or U13313 (N_13313,N_11100,N_9549);
nand U13314 (N_13314,N_10409,N_10002);
or U13315 (N_13315,N_11589,N_10415);
nand U13316 (N_13316,N_9258,N_11401);
nor U13317 (N_13317,N_9841,N_11008);
nor U13318 (N_13318,N_10283,N_11006);
and U13319 (N_13319,N_11470,N_10193);
nor U13320 (N_13320,N_10263,N_11172);
nor U13321 (N_13321,N_11345,N_10818);
and U13322 (N_13322,N_11214,N_10147);
or U13323 (N_13323,N_11916,N_9775);
xnor U13324 (N_13324,N_10591,N_10962);
nor U13325 (N_13325,N_10220,N_10827);
or U13326 (N_13326,N_11585,N_9296);
and U13327 (N_13327,N_10305,N_11787);
or U13328 (N_13328,N_10026,N_9675);
or U13329 (N_13329,N_10915,N_9762);
and U13330 (N_13330,N_10706,N_11878);
nand U13331 (N_13331,N_11468,N_11534);
or U13332 (N_13332,N_10737,N_11600);
and U13333 (N_13333,N_10582,N_11213);
or U13334 (N_13334,N_11123,N_11013);
or U13335 (N_13335,N_9988,N_10056);
xnor U13336 (N_13336,N_9672,N_11923);
or U13337 (N_13337,N_11474,N_10416);
nand U13338 (N_13338,N_11568,N_11161);
and U13339 (N_13339,N_9555,N_10154);
nand U13340 (N_13340,N_11862,N_11992);
nor U13341 (N_13341,N_10209,N_9368);
nand U13342 (N_13342,N_11398,N_9761);
or U13343 (N_13343,N_11334,N_9240);
or U13344 (N_13344,N_11178,N_11771);
and U13345 (N_13345,N_9851,N_11269);
and U13346 (N_13346,N_9012,N_9833);
nand U13347 (N_13347,N_11542,N_11402);
nor U13348 (N_13348,N_11405,N_11661);
nor U13349 (N_13349,N_9388,N_9455);
or U13350 (N_13350,N_11788,N_11695);
nand U13351 (N_13351,N_11031,N_9266);
nand U13352 (N_13352,N_11538,N_11531);
nand U13353 (N_13353,N_11204,N_9606);
nor U13354 (N_13354,N_10811,N_9857);
nor U13355 (N_13355,N_9769,N_9351);
nor U13356 (N_13356,N_10944,N_10064);
or U13357 (N_13357,N_10384,N_10272);
or U13358 (N_13358,N_9156,N_9681);
or U13359 (N_13359,N_10908,N_11135);
and U13360 (N_13360,N_11092,N_9186);
and U13361 (N_13361,N_11885,N_11397);
or U13362 (N_13362,N_10790,N_9329);
nand U13363 (N_13363,N_9940,N_11962);
and U13364 (N_13364,N_10098,N_9991);
nor U13365 (N_13365,N_10902,N_11215);
nor U13366 (N_13366,N_11732,N_10845);
and U13367 (N_13367,N_10472,N_11221);
or U13368 (N_13368,N_10356,N_10964);
and U13369 (N_13369,N_9216,N_9028);
or U13370 (N_13370,N_10423,N_11171);
nand U13371 (N_13371,N_10089,N_10126);
or U13372 (N_13372,N_9807,N_11729);
and U13373 (N_13373,N_10087,N_9644);
or U13374 (N_13374,N_11319,N_11076);
and U13375 (N_13375,N_11336,N_9510);
or U13376 (N_13376,N_10975,N_10155);
and U13377 (N_13377,N_11516,N_9842);
or U13378 (N_13378,N_9230,N_10411);
and U13379 (N_13379,N_11555,N_10720);
nand U13380 (N_13380,N_10226,N_10128);
nor U13381 (N_13381,N_10130,N_10045);
or U13382 (N_13382,N_10930,N_10542);
nor U13383 (N_13383,N_10217,N_9642);
and U13384 (N_13384,N_10058,N_10258);
or U13385 (N_13385,N_10609,N_10300);
or U13386 (N_13386,N_9387,N_11121);
and U13387 (N_13387,N_9019,N_9827);
nand U13388 (N_13388,N_10007,N_9474);
or U13389 (N_13389,N_11572,N_10832);
nand U13390 (N_13390,N_10194,N_10370);
and U13391 (N_13391,N_10590,N_11664);
or U13392 (N_13392,N_10713,N_11278);
nand U13393 (N_13393,N_9843,N_10918);
or U13394 (N_13394,N_10639,N_10894);
nor U13395 (N_13395,N_11446,N_10772);
and U13396 (N_13396,N_9639,N_11724);
and U13397 (N_13397,N_11304,N_10042);
nor U13398 (N_13398,N_9112,N_11289);
nand U13399 (N_13399,N_9602,N_9052);
nand U13400 (N_13400,N_9123,N_9111);
and U13401 (N_13401,N_10475,N_10502);
nor U13402 (N_13402,N_9399,N_9223);
and U13403 (N_13403,N_11912,N_10013);
and U13404 (N_13404,N_9908,N_9459);
nor U13405 (N_13405,N_10954,N_11809);
and U13406 (N_13406,N_10386,N_10434);
or U13407 (N_13407,N_11629,N_11619);
nor U13408 (N_13408,N_10545,N_11058);
or U13409 (N_13409,N_10773,N_10268);
or U13410 (N_13410,N_10314,N_11682);
or U13411 (N_13411,N_11833,N_11378);
or U13412 (N_13412,N_10487,N_11189);
nand U13413 (N_13413,N_9687,N_11296);
nand U13414 (N_13414,N_11094,N_11758);
nor U13415 (N_13415,N_10161,N_11756);
or U13416 (N_13416,N_11922,N_10847);
nor U13417 (N_13417,N_9157,N_11828);
and U13418 (N_13418,N_9854,N_10495);
nand U13419 (N_13419,N_9315,N_11881);
nor U13420 (N_13420,N_9140,N_10595);
and U13421 (N_13421,N_11224,N_11792);
nor U13422 (N_13422,N_10470,N_10935);
or U13423 (N_13423,N_10521,N_10187);
or U13424 (N_13424,N_10353,N_9204);
or U13425 (N_13425,N_9090,N_11375);
and U13426 (N_13426,N_11433,N_11616);
nand U13427 (N_13427,N_9989,N_11067);
nand U13428 (N_13428,N_9036,N_9436);
nor U13429 (N_13429,N_11980,N_10746);
nor U13430 (N_13430,N_11326,N_11368);
nor U13431 (N_13431,N_9568,N_11519);
or U13432 (N_13432,N_11659,N_9424);
or U13433 (N_13433,N_9154,N_9249);
or U13434 (N_13434,N_11553,N_10420);
nor U13435 (N_13435,N_11635,N_9507);
nand U13436 (N_13436,N_10319,N_9784);
or U13437 (N_13437,N_11245,N_9196);
and U13438 (N_13438,N_9905,N_9764);
nor U13439 (N_13439,N_11114,N_11046);
nor U13440 (N_13440,N_9918,N_9072);
or U13441 (N_13441,N_11864,N_9840);
or U13442 (N_13442,N_9442,N_11846);
nand U13443 (N_13443,N_9610,N_11602);
nor U13444 (N_13444,N_10091,N_11039);
nand U13445 (N_13445,N_9868,N_10180);
and U13446 (N_13446,N_10035,N_9727);
nand U13447 (N_13447,N_11631,N_11874);
nand U13448 (N_13448,N_9367,N_10576);
or U13449 (N_13449,N_9398,N_11976);
nand U13450 (N_13450,N_9955,N_10634);
nor U13451 (N_13451,N_11440,N_9403);
or U13452 (N_13452,N_9326,N_11488);
and U13453 (N_13453,N_9380,N_10651);
and U13454 (N_13454,N_11243,N_10196);
or U13455 (N_13455,N_11451,N_11743);
nor U13456 (N_13456,N_11075,N_11038);
nand U13457 (N_13457,N_10046,N_10279);
nand U13458 (N_13458,N_11578,N_9411);
nand U13459 (N_13459,N_9096,N_10552);
nor U13460 (N_13460,N_9485,N_11327);
nand U13461 (N_13461,N_11175,N_11443);
and U13462 (N_13462,N_10536,N_10232);
nand U13463 (N_13463,N_10721,N_11767);
nor U13464 (N_13464,N_11679,N_10689);
and U13465 (N_13465,N_10496,N_9888);
nor U13466 (N_13466,N_10996,N_11351);
nand U13467 (N_13467,N_10099,N_9298);
nor U13468 (N_13468,N_11565,N_11392);
nor U13469 (N_13469,N_10203,N_9145);
nor U13470 (N_13470,N_9755,N_10755);
and U13471 (N_13471,N_9766,N_10683);
nand U13472 (N_13472,N_9563,N_11084);
and U13473 (N_13473,N_10250,N_9707);
nor U13474 (N_13474,N_10752,N_10231);
nand U13475 (N_13475,N_10767,N_10403);
and U13476 (N_13476,N_9661,N_11396);
and U13477 (N_13477,N_9180,N_9745);
and U13478 (N_13478,N_9616,N_9990);
and U13479 (N_13479,N_9504,N_10593);
nand U13480 (N_13480,N_10601,N_11434);
nand U13481 (N_13481,N_11184,N_11380);
or U13482 (N_13482,N_9890,N_9445);
and U13483 (N_13483,N_10853,N_10340);
and U13484 (N_13484,N_10453,N_11348);
or U13485 (N_13485,N_11728,N_9077);
nand U13486 (N_13486,N_9408,N_11344);
and U13487 (N_13487,N_10533,N_10398);
nor U13488 (N_13488,N_11227,N_11691);
nor U13489 (N_13489,N_11666,N_9528);
nand U13490 (N_13490,N_11330,N_11880);
and U13491 (N_13491,N_11399,N_9159);
and U13492 (N_13492,N_11212,N_9539);
nor U13493 (N_13493,N_9432,N_10878);
and U13494 (N_13494,N_11037,N_9998);
and U13495 (N_13495,N_11548,N_10765);
nor U13496 (N_13496,N_9427,N_9374);
nand U13497 (N_13497,N_9429,N_10909);
nor U13498 (N_13498,N_9865,N_10173);
nor U13499 (N_13499,N_11461,N_11127);
nor U13500 (N_13500,N_11728,N_10360);
nor U13501 (N_13501,N_11786,N_11327);
or U13502 (N_13502,N_10358,N_11908);
nand U13503 (N_13503,N_9550,N_11209);
nor U13504 (N_13504,N_11221,N_9754);
nor U13505 (N_13505,N_11117,N_11157);
or U13506 (N_13506,N_11527,N_9053);
and U13507 (N_13507,N_11777,N_11186);
or U13508 (N_13508,N_11316,N_10232);
nand U13509 (N_13509,N_10668,N_10369);
and U13510 (N_13510,N_10238,N_10900);
and U13511 (N_13511,N_11780,N_9760);
nor U13512 (N_13512,N_11522,N_10024);
or U13513 (N_13513,N_11328,N_9306);
nand U13514 (N_13514,N_11806,N_10473);
nand U13515 (N_13515,N_10366,N_9951);
or U13516 (N_13516,N_9024,N_11417);
or U13517 (N_13517,N_10695,N_9831);
nor U13518 (N_13518,N_11456,N_11725);
or U13519 (N_13519,N_9805,N_9651);
or U13520 (N_13520,N_11270,N_11167);
and U13521 (N_13521,N_10080,N_10626);
nand U13522 (N_13522,N_10513,N_9863);
and U13523 (N_13523,N_11456,N_9123);
and U13524 (N_13524,N_11758,N_11465);
nand U13525 (N_13525,N_10266,N_9094);
and U13526 (N_13526,N_11887,N_11254);
nor U13527 (N_13527,N_10119,N_10294);
and U13528 (N_13528,N_11203,N_10812);
nor U13529 (N_13529,N_10380,N_9671);
or U13530 (N_13530,N_9830,N_10802);
and U13531 (N_13531,N_11575,N_9363);
xor U13532 (N_13532,N_9732,N_9782);
and U13533 (N_13533,N_9009,N_10502);
and U13534 (N_13534,N_10941,N_11990);
nor U13535 (N_13535,N_10558,N_10310);
and U13536 (N_13536,N_9537,N_11601);
or U13537 (N_13537,N_11097,N_11373);
and U13538 (N_13538,N_9848,N_9155);
nand U13539 (N_13539,N_9604,N_11428);
or U13540 (N_13540,N_9840,N_11123);
nand U13541 (N_13541,N_11494,N_11872);
nor U13542 (N_13542,N_9783,N_9917);
nand U13543 (N_13543,N_9879,N_11167);
and U13544 (N_13544,N_11216,N_11130);
nand U13545 (N_13545,N_10220,N_10200);
and U13546 (N_13546,N_10529,N_9561);
nand U13547 (N_13547,N_9361,N_9076);
and U13548 (N_13548,N_10076,N_9640);
or U13549 (N_13549,N_9739,N_11218);
or U13550 (N_13550,N_9261,N_9945);
or U13551 (N_13551,N_10538,N_9859);
nand U13552 (N_13552,N_11494,N_9898);
and U13553 (N_13553,N_11198,N_11908);
nand U13554 (N_13554,N_9699,N_10710);
or U13555 (N_13555,N_10746,N_9214);
nor U13556 (N_13556,N_9156,N_9857);
and U13557 (N_13557,N_11616,N_10923);
or U13558 (N_13558,N_10684,N_11210);
and U13559 (N_13559,N_9849,N_10212);
or U13560 (N_13560,N_9300,N_10576);
nor U13561 (N_13561,N_11477,N_11147);
and U13562 (N_13562,N_11753,N_11825);
nand U13563 (N_13563,N_11876,N_9993);
nand U13564 (N_13564,N_11779,N_9172);
nor U13565 (N_13565,N_11328,N_11715);
nor U13566 (N_13566,N_9410,N_9215);
nand U13567 (N_13567,N_9983,N_10580);
nand U13568 (N_13568,N_11607,N_11356);
nor U13569 (N_13569,N_9475,N_9491);
or U13570 (N_13570,N_9156,N_10201);
or U13571 (N_13571,N_10480,N_11246);
nand U13572 (N_13572,N_9092,N_11384);
nand U13573 (N_13573,N_10496,N_9519);
and U13574 (N_13574,N_11459,N_10561);
and U13575 (N_13575,N_9624,N_10687);
and U13576 (N_13576,N_10541,N_11461);
and U13577 (N_13577,N_11102,N_9167);
nor U13578 (N_13578,N_11696,N_10934);
and U13579 (N_13579,N_11033,N_11757);
and U13580 (N_13580,N_9425,N_11134);
nand U13581 (N_13581,N_11640,N_10374);
or U13582 (N_13582,N_10606,N_11632);
nor U13583 (N_13583,N_10574,N_10131);
or U13584 (N_13584,N_9070,N_10258);
and U13585 (N_13585,N_10100,N_9881);
nand U13586 (N_13586,N_11531,N_10825);
nand U13587 (N_13587,N_10095,N_11958);
and U13588 (N_13588,N_10999,N_10421);
and U13589 (N_13589,N_10951,N_9668);
or U13590 (N_13590,N_9767,N_9211);
nand U13591 (N_13591,N_9075,N_11784);
and U13592 (N_13592,N_9992,N_10503);
and U13593 (N_13593,N_10015,N_10476);
or U13594 (N_13594,N_9343,N_10326);
and U13595 (N_13595,N_10708,N_11024);
nand U13596 (N_13596,N_10261,N_11358);
or U13597 (N_13597,N_10273,N_9066);
or U13598 (N_13598,N_11553,N_11661);
nor U13599 (N_13599,N_10449,N_10618);
nand U13600 (N_13600,N_11845,N_9596);
xnor U13601 (N_13601,N_9662,N_9638);
and U13602 (N_13602,N_10515,N_11664);
nor U13603 (N_13603,N_11074,N_9929);
xnor U13604 (N_13604,N_10882,N_9173);
nand U13605 (N_13605,N_9700,N_10915);
or U13606 (N_13606,N_9488,N_9332);
nand U13607 (N_13607,N_11475,N_10432);
or U13608 (N_13608,N_11231,N_10178);
and U13609 (N_13609,N_9923,N_11104);
and U13610 (N_13610,N_11713,N_11751);
nand U13611 (N_13611,N_9709,N_9357);
nor U13612 (N_13612,N_9254,N_11147);
or U13613 (N_13613,N_9058,N_10477);
nand U13614 (N_13614,N_11337,N_11888);
and U13615 (N_13615,N_11906,N_9378);
nor U13616 (N_13616,N_11868,N_10303);
or U13617 (N_13617,N_10671,N_11135);
nand U13618 (N_13618,N_10630,N_10777);
nand U13619 (N_13619,N_11353,N_11571);
and U13620 (N_13620,N_9175,N_10372);
nor U13621 (N_13621,N_10204,N_9415);
nand U13622 (N_13622,N_10147,N_9916);
nor U13623 (N_13623,N_11606,N_10121);
nand U13624 (N_13624,N_9611,N_10159);
and U13625 (N_13625,N_11184,N_10059);
nor U13626 (N_13626,N_9426,N_9071);
and U13627 (N_13627,N_9028,N_9390);
nor U13628 (N_13628,N_11666,N_11891);
or U13629 (N_13629,N_9444,N_9967);
nand U13630 (N_13630,N_10932,N_9396);
or U13631 (N_13631,N_11706,N_10647);
or U13632 (N_13632,N_9628,N_9319);
nor U13633 (N_13633,N_9941,N_9667);
nor U13634 (N_13634,N_10659,N_10383);
nor U13635 (N_13635,N_11309,N_11358);
or U13636 (N_13636,N_11977,N_9704);
nand U13637 (N_13637,N_10041,N_10090);
or U13638 (N_13638,N_10347,N_11582);
nand U13639 (N_13639,N_11734,N_11226);
or U13640 (N_13640,N_9707,N_9161);
nor U13641 (N_13641,N_11083,N_10395);
or U13642 (N_13642,N_9776,N_9929);
nand U13643 (N_13643,N_11007,N_10567);
nand U13644 (N_13644,N_9896,N_11276);
nor U13645 (N_13645,N_10956,N_11592);
and U13646 (N_13646,N_10047,N_10389);
or U13647 (N_13647,N_11761,N_10928);
or U13648 (N_13648,N_11967,N_11769);
or U13649 (N_13649,N_11348,N_9657);
and U13650 (N_13650,N_9704,N_9499);
nor U13651 (N_13651,N_10597,N_11453);
or U13652 (N_13652,N_11179,N_9142);
or U13653 (N_13653,N_9420,N_11428);
nor U13654 (N_13654,N_10195,N_9946);
and U13655 (N_13655,N_9474,N_9036);
and U13656 (N_13656,N_10620,N_10160);
and U13657 (N_13657,N_9939,N_10462);
and U13658 (N_13658,N_11351,N_11036);
and U13659 (N_13659,N_11536,N_10440);
and U13660 (N_13660,N_11439,N_10329);
nand U13661 (N_13661,N_11865,N_10860);
nor U13662 (N_13662,N_11489,N_9668);
nor U13663 (N_13663,N_9894,N_10457);
and U13664 (N_13664,N_9476,N_11579);
nand U13665 (N_13665,N_11418,N_9104);
and U13666 (N_13666,N_9930,N_10770);
nand U13667 (N_13667,N_9086,N_11997);
or U13668 (N_13668,N_9063,N_11208);
xnor U13669 (N_13669,N_11995,N_10199);
and U13670 (N_13670,N_10221,N_11521);
and U13671 (N_13671,N_11529,N_10208);
nand U13672 (N_13672,N_9608,N_10535);
nor U13673 (N_13673,N_10341,N_10942);
and U13674 (N_13674,N_9558,N_10004);
nand U13675 (N_13675,N_11933,N_9752);
or U13676 (N_13676,N_9486,N_11235);
and U13677 (N_13677,N_11188,N_10267);
nor U13678 (N_13678,N_11342,N_11890);
and U13679 (N_13679,N_9510,N_9770);
nor U13680 (N_13680,N_10626,N_9380);
xor U13681 (N_13681,N_11867,N_11536);
nor U13682 (N_13682,N_9332,N_11852);
and U13683 (N_13683,N_9777,N_10150);
nor U13684 (N_13684,N_10988,N_10584);
and U13685 (N_13685,N_11336,N_10809);
or U13686 (N_13686,N_9968,N_9265);
or U13687 (N_13687,N_9591,N_10507);
nand U13688 (N_13688,N_9462,N_9977);
xnor U13689 (N_13689,N_11261,N_9229);
xor U13690 (N_13690,N_9562,N_9092);
and U13691 (N_13691,N_11114,N_11098);
nor U13692 (N_13692,N_9141,N_9765);
nand U13693 (N_13693,N_10798,N_10304);
nor U13694 (N_13694,N_9867,N_10921);
or U13695 (N_13695,N_11957,N_9920);
nor U13696 (N_13696,N_11813,N_9714);
or U13697 (N_13697,N_11443,N_11648);
or U13698 (N_13698,N_11833,N_10460);
and U13699 (N_13699,N_11534,N_11672);
or U13700 (N_13700,N_9593,N_11888);
nand U13701 (N_13701,N_9076,N_11059);
nor U13702 (N_13702,N_9066,N_11929);
or U13703 (N_13703,N_9156,N_11323);
or U13704 (N_13704,N_9075,N_10312);
and U13705 (N_13705,N_11171,N_9521);
and U13706 (N_13706,N_10875,N_9097);
or U13707 (N_13707,N_11568,N_11932);
nand U13708 (N_13708,N_10817,N_11441);
and U13709 (N_13709,N_11463,N_10154);
or U13710 (N_13710,N_9684,N_10486);
nand U13711 (N_13711,N_10708,N_9406);
and U13712 (N_13712,N_11480,N_10007);
nor U13713 (N_13713,N_9767,N_10231);
nand U13714 (N_13714,N_11124,N_11587);
and U13715 (N_13715,N_10348,N_10938);
or U13716 (N_13716,N_10670,N_9915);
nand U13717 (N_13717,N_10352,N_9142);
and U13718 (N_13718,N_10612,N_11031);
nor U13719 (N_13719,N_10583,N_10214);
or U13720 (N_13720,N_10877,N_11224);
nand U13721 (N_13721,N_9442,N_9800);
nand U13722 (N_13722,N_9778,N_11427);
xnor U13723 (N_13723,N_11135,N_11622);
nand U13724 (N_13724,N_11481,N_9373);
nor U13725 (N_13725,N_11594,N_11784);
nor U13726 (N_13726,N_11078,N_9541);
and U13727 (N_13727,N_10278,N_9015);
or U13728 (N_13728,N_11729,N_10464);
nand U13729 (N_13729,N_10817,N_11054);
nor U13730 (N_13730,N_10981,N_11851);
or U13731 (N_13731,N_9739,N_9040);
nor U13732 (N_13732,N_11965,N_11668);
or U13733 (N_13733,N_10395,N_10600);
or U13734 (N_13734,N_11920,N_9867);
and U13735 (N_13735,N_11557,N_9454);
nor U13736 (N_13736,N_11128,N_11044);
and U13737 (N_13737,N_11935,N_11135);
and U13738 (N_13738,N_9884,N_9954);
nand U13739 (N_13739,N_10113,N_11485);
nand U13740 (N_13740,N_10069,N_9365);
nand U13741 (N_13741,N_10661,N_9233);
nor U13742 (N_13742,N_10180,N_10757);
nand U13743 (N_13743,N_9427,N_11679);
and U13744 (N_13744,N_10118,N_9084);
or U13745 (N_13745,N_11655,N_10152);
nand U13746 (N_13746,N_9040,N_9655);
nor U13747 (N_13747,N_11710,N_9886);
and U13748 (N_13748,N_11800,N_9352);
and U13749 (N_13749,N_10425,N_10708);
nand U13750 (N_13750,N_10326,N_11423);
and U13751 (N_13751,N_10024,N_11995);
and U13752 (N_13752,N_11827,N_10978);
and U13753 (N_13753,N_11708,N_11721);
or U13754 (N_13754,N_11661,N_10643);
nor U13755 (N_13755,N_10729,N_11691);
nand U13756 (N_13756,N_11958,N_9741);
nor U13757 (N_13757,N_11140,N_11213);
nor U13758 (N_13758,N_11779,N_10064);
nand U13759 (N_13759,N_10349,N_11995);
nand U13760 (N_13760,N_11727,N_9575);
and U13761 (N_13761,N_11417,N_9919);
or U13762 (N_13762,N_10052,N_10393);
and U13763 (N_13763,N_9229,N_9342);
nand U13764 (N_13764,N_9348,N_9968);
or U13765 (N_13765,N_11078,N_10449);
or U13766 (N_13766,N_10561,N_9891);
and U13767 (N_13767,N_9042,N_10166);
nor U13768 (N_13768,N_9676,N_10589);
and U13769 (N_13769,N_10416,N_9910);
nand U13770 (N_13770,N_9012,N_10986);
or U13771 (N_13771,N_9823,N_9549);
or U13772 (N_13772,N_11069,N_9004);
or U13773 (N_13773,N_9113,N_11087);
and U13774 (N_13774,N_10060,N_9895);
nand U13775 (N_13775,N_10407,N_11106);
nand U13776 (N_13776,N_9439,N_9528);
xor U13777 (N_13777,N_11283,N_10604);
nand U13778 (N_13778,N_9183,N_11667);
nor U13779 (N_13779,N_10282,N_9052);
nor U13780 (N_13780,N_10786,N_10501);
nor U13781 (N_13781,N_9655,N_10435);
nor U13782 (N_13782,N_10124,N_11839);
xnor U13783 (N_13783,N_9440,N_9974);
and U13784 (N_13784,N_10060,N_9088);
nor U13785 (N_13785,N_11196,N_11152);
or U13786 (N_13786,N_10506,N_10022);
and U13787 (N_13787,N_10618,N_10056);
and U13788 (N_13788,N_10123,N_11735);
nand U13789 (N_13789,N_11086,N_11863);
nand U13790 (N_13790,N_9555,N_9710);
nand U13791 (N_13791,N_11523,N_9057);
and U13792 (N_13792,N_9421,N_11312);
or U13793 (N_13793,N_10942,N_11999);
nor U13794 (N_13794,N_9995,N_10506);
nand U13795 (N_13795,N_9864,N_10430);
nand U13796 (N_13796,N_9830,N_9110);
or U13797 (N_13797,N_10424,N_9411);
nand U13798 (N_13798,N_9493,N_11591);
nand U13799 (N_13799,N_10877,N_9015);
or U13800 (N_13800,N_11553,N_9049);
or U13801 (N_13801,N_10029,N_9164);
nor U13802 (N_13802,N_11537,N_10809);
nand U13803 (N_13803,N_9376,N_10097);
or U13804 (N_13804,N_9879,N_11472);
nor U13805 (N_13805,N_9923,N_10736);
nand U13806 (N_13806,N_11131,N_9095);
nand U13807 (N_13807,N_9289,N_9602);
nand U13808 (N_13808,N_9340,N_10363);
nand U13809 (N_13809,N_11293,N_10244);
and U13810 (N_13810,N_9173,N_11763);
nor U13811 (N_13811,N_10841,N_9124);
and U13812 (N_13812,N_10649,N_9887);
nor U13813 (N_13813,N_11921,N_11917);
or U13814 (N_13814,N_9100,N_11935);
and U13815 (N_13815,N_9174,N_11851);
and U13816 (N_13816,N_10901,N_9789);
and U13817 (N_13817,N_9520,N_11981);
and U13818 (N_13818,N_9168,N_9843);
or U13819 (N_13819,N_11533,N_10683);
or U13820 (N_13820,N_9481,N_9889);
nor U13821 (N_13821,N_10585,N_10663);
nor U13822 (N_13822,N_9133,N_9618);
or U13823 (N_13823,N_10967,N_10370);
nor U13824 (N_13824,N_11251,N_10716);
nor U13825 (N_13825,N_10330,N_10147);
or U13826 (N_13826,N_9119,N_10212);
nand U13827 (N_13827,N_10079,N_11106);
nand U13828 (N_13828,N_11006,N_11584);
nand U13829 (N_13829,N_9641,N_11420);
and U13830 (N_13830,N_9569,N_9928);
nand U13831 (N_13831,N_9285,N_10048);
and U13832 (N_13832,N_10331,N_10467);
or U13833 (N_13833,N_10892,N_9629);
and U13834 (N_13834,N_11399,N_10675);
and U13835 (N_13835,N_10311,N_10743);
or U13836 (N_13836,N_11134,N_9528);
nand U13837 (N_13837,N_9450,N_10781);
or U13838 (N_13838,N_11283,N_9417);
nand U13839 (N_13839,N_9115,N_9109);
or U13840 (N_13840,N_11279,N_11562);
nor U13841 (N_13841,N_10617,N_9827);
nor U13842 (N_13842,N_9186,N_9303);
and U13843 (N_13843,N_10718,N_10680);
nor U13844 (N_13844,N_9197,N_10197);
nor U13845 (N_13845,N_9852,N_11703);
nand U13846 (N_13846,N_10545,N_10961);
nor U13847 (N_13847,N_10156,N_9964);
nor U13848 (N_13848,N_11391,N_9178);
or U13849 (N_13849,N_10536,N_10451);
or U13850 (N_13850,N_9649,N_10813);
nand U13851 (N_13851,N_10045,N_11590);
or U13852 (N_13852,N_11864,N_9781);
nor U13853 (N_13853,N_9899,N_10218);
nor U13854 (N_13854,N_10736,N_11153);
nor U13855 (N_13855,N_10500,N_10857);
nor U13856 (N_13856,N_10307,N_10847);
nor U13857 (N_13857,N_10221,N_11076);
or U13858 (N_13858,N_10114,N_10367);
nor U13859 (N_13859,N_9924,N_10567);
or U13860 (N_13860,N_10350,N_10734);
nand U13861 (N_13861,N_10513,N_11227);
nand U13862 (N_13862,N_9771,N_9189);
or U13863 (N_13863,N_10671,N_9230);
or U13864 (N_13864,N_11787,N_9946);
nand U13865 (N_13865,N_9569,N_11947);
nand U13866 (N_13866,N_11973,N_11920);
nand U13867 (N_13867,N_9292,N_10784);
or U13868 (N_13868,N_10756,N_10278);
and U13869 (N_13869,N_11970,N_11530);
nand U13870 (N_13870,N_10376,N_9842);
and U13871 (N_13871,N_9430,N_11902);
or U13872 (N_13872,N_11250,N_10005);
or U13873 (N_13873,N_10846,N_10753);
and U13874 (N_13874,N_10491,N_9758);
and U13875 (N_13875,N_11353,N_10153);
and U13876 (N_13876,N_10088,N_11361);
nor U13877 (N_13877,N_10613,N_11544);
nor U13878 (N_13878,N_9778,N_11612);
or U13879 (N_13879,N_9436,N_9627);
nand U13880 (N_13880,N_11856,N_11326);
nand U13881 (N_13881,N_11041,N_9772);
nand U13882 (N_13882,N_10712,N_10579);
or U13883 (N_13883,N_11424,N_11551);
and U13884 (N_13884,N_10915,N_9489);
or U13885 (N_13885,N_9084,N_11003);
or U13886 (N_13886,N_9553,N_9030);
nor U13887 (N_13887,N_10428,N_9041);
and U13888 (N_13888,N_10040,N_9612);
or U13889 (N_13889,N_10900,N_9611);
or U13890 (N_13890,N_10445,N_11701);
or U13891 (N_13891,N_9644,N_10565);
and U13892 (N_13892,N_10958,N_10695);
nor U13893 (N_13893,N_11352,N_11940);
nor U13894 (N_13894,N_11405,N_10383);
nor U13895 (N_13895,N_11520,N_11104);
nor U13896 (N_13896,N_11925,N_11562);
or U13897 (N_13897,N_10272,N_11882);
nand U13898 (N_13898,N_10858,N_9160);
and U13899 (N_13899,N_10283,N_10540);
or U13900 (N_13900,N_11968,N_11100);
and U13901 (N_13901,N_9456,N_10918);
nand U13902 (N_13902,N_10372,N_11038);
nor U13903 (N_13903,N_11827,N_10817);
or U13904 (N_13904,N_11345,N_11112);
and U13905 (N_13905,N_10191,N_9422);
nand U13906 (N_13906,N_11359,N_10768);
or U13907 (N_13907,N_11551,N_11855);
or U13908 (N_13908,N_11254,N_11754);
nand U13909 (N_13909,N_11340,N_9832);
nor U13910 (N_13910,N_9800,N_10175);
nand U13911 (N_13911,N_10299,N_9313);
and U13912 (N_13912,N_9113,N_11308);
nor U13913 (N_13913,N_9986,N_11986);
and U13914 (N_13914,N_10973,N_11223);
nor U13915 (N_13915,N_10444,N_10761);
and U13916 (N_13916,N_9527,N_10571);
and U13917 (N_13917,N_11850,N_9815);
nand U13918 (N_13918,N_10911,N_9999);
and U13919 (N_13919,N_11282,N_9522);
or U13920 (N_13920,N_11349,N_9934);
nor U13921 (N_13921,N_9719,N_10205);
nand U13922 (N_13922,N_10289,N_10883);
nand U13923 (N_13923,N_10675,N_9294);
nand U13924 (N_13924,N_10966,N_10831);
or U13925 (N_13925,N_10224,N_11492);
and U13926 (N_13926,N_9389,N_11128);
and U13927 (N_13927,N_9135,N_10891);
and U13928 (N_13928,N_10607,N_9157);
nand U13929 (N_13929,N_11587,N_9085);
and U13930 (N_13930,N_9871,N_9439);
or U13931 (N_13931,N_10734,N_9842);
nand U13932 (N_13932,N_9817,N_10098);
and U13933 (N_13933,N_9917,N_9693);
nand U13934 (N_13934,N_10428,N_9795);
nand U13935 (N_13935,N_9085,N_9950);
and U13936 (N_13936,N_10422,N_10047);
nor U13937 (N_13937,N_11922,N_11783);
nor U13938 (N_13938,N_9146,N_10336);
nor U13939 (N_13939,N_9268,N_11642);
and U13940 (N_13940,N_9101,N_9715);
nor U13941 (N_13941,N_10845,N_10540);
nor U13942 (N_13942,N_10608,N_10692);
or U13943 (N_13943,N_10703,N_9306);
or U13944 (N_13944,N_11886,N_9418);
nand U13945 (N_13945,N_10508,N_9141);
nand U13946 (N_13946,N_9298,N_10467);
or U13947 (N_13947,N_11765,N_10980);
and U13948 (N_13948,N_10822,N_10151);
or U13949 (N_13949,N_10434,N_10169);
and U13950 (N_13950,N_9291,N_11755);
or U13951 (N_13951,N_10514,N_9195);
nand U13952 (N_13952,N_10429,N_9462);
and U13953 (N_13953,N_9474,N_9550);
and U13954 (N_13954,N_11004,N_9025);
and U13955 (N_13955,N_9183,N_9738);
and U13956 (N_13956,N_9981,N_11773);
nand U13957 (N_13957,N_10680,N_11059);
and U13958 (N_13958,N_9635,N_10627);
nor U13959 (N_13959,N_11280,N_11356);
nor U13960 (N_13960,N_9600,N_9606);
and U13961 (N_13961,N_11187,N_9661);
nor U13962 (N_13962,N_9871,N_10081);
nand U13963 (N_13963,N_9491,N_9608);
and U13964 (N_13964,N_10262,N_9290);
or U13965 (N_13965,N_9355,N_11526);
and U13966 (N_13966,N_9535,N_9913);
and U13967 (N_13967,N_10460,N_10021);
and U13968 (N_13968,N_11366,N_9252);
nor U13969 (N_13969,N_9722,N_10214);
nor U13970 (N_13970,N_9761,N_10459);
nor U13971 (N_13971,N_11033,N_10798);
and U13972 (N_13972,N_9195,N_10111);
or U13973 (N_13973,N_10902,N_11880);
or U13974 (N_13974,N_10874,N_10231);
nor U13975 (N_13975,N_11348,N_11929);
nand U13976 (N_13976,N_9280,N_11826);
nor U13977 (N_13977,N_10931,N_11776);
nand U13978 (N_13978,N_10789,N_9707);
nor U13979 (N_13979,N_9763,N_9168);
or U13980 (N_13980,N_9836,N_11317);
or U13981 (N_13981,N_9233,N_10744);
nand U13982 (N_13982,N_10545,N_11651);
nor U13983 (N_13983,N_11447,N_9474);
nand U13984 (N_13984,N_11736,N_11611);
xnor U13985 (N_13985,N_10681,N_11287);
or U13986 (N_13986,N_11689,N_10853);
nand U13987 (N_13987,N_9150,N_9885);
and U13988 (N_13988,N_10514,N_10560);
or U13989 (N_13989,N_11422,N_9912);
and U13990 (N_13990,N_11083,N_10071);
or U13991 (N_13991,N_9604,N_10520);
nand U13992 (N_13992,N_11231,N_10061);
or U13993 (N_13993,N_11773,N_9909);
and U13994 (N_13994,N_10260,N_9848);
and U13995 (N_13995,N_11354,N_9448);
or U13996 (N_13996,N_9956,N_9504);
nand U13997 (N_13997,N_11318,N_9942);
nand U13998 (N_13998,N_10074,N_9664);
or U13999 (N_13999,N_10692,N_11715);
nand U14000 (N_14000,N_9730,N_9333);
nand U14001 (N_14001,N_9615,N_10913);
and U14002 (N_14002,N_10207,N_11975);
nand U14003 (N_14003,N_10806,N_9654);
nor U14004 (N_14004,N_11862,N_9280);
nor U14005 (N_14005,N_10168,N_9848);
nand U14006 (N_14006,N_9336,N_10890);
nand U14007 (N_14007,N_9878,N_10683);
and U14008 (N_14008,N_11493,N_10181);
and U14009 (N_14009,N_11113,N_10594);
nand U14010 (N_14010,N_11783,N_10384);
and U14011 (N_14011,N_9824,N_11819);
and U14012 (N_14012,N_11086,N_11591);
nor U14013 (N_14013,N_10186,N_10671);
nor U14014 (N_14014,N_11432,N_10809);
or U14015 (N_14015,N_9716,N_11083);
xor U14016 (N_14016,N_10121,N_11411);
and U14017 (N_14017,N_9636,N_10301);
or U14018 (N_14018,N_10897,N_10934);
nand U14019 (N_14019,N_9092,N_9277);
nor U14020 (N_14020,N_11784,N_11532);
nand U14021 (N_14021,N_11820,N_9805);
nand U14022 (N_14022,N_11570,N_11049);
and U14023 (N_14023,N_9268,N_9552);
nor U14024 (N_14024,N_10411,N_9500);
and U14025 (N_14025,N_11716,N_9418);
and U14026 (N_14026,N_10985,N_11214);
nor U14027 (N_14027,N_10176,N_11670);
and U14028 (N_14028,N_9718,N_9202);
and U14029 (N_14029,N_9194,N_9348);
nand U14030 (N_14030,N_9908,N_11320);
and U14031 (N_14031,N_9344,N_10176);
or U14032 (N_14032,N_9916,N_9078);
nor U14033 (N_14033,N_11965,N_9465);
nor U14034 (N_14034,N_11386,N_9674);
nor U14035 (N_14035,N_11822,N_9369);
or U14036 (N_14036,N_9258,N_11238);
or U14037 (N_14037,N_10787,N_10018);
or U14038 (N_14038,N_10810,N_9102);
nor U14039 (N_14039,N_9547,N_11673);
or U14040 (N_14040,N_10750,N_10488);
and U14041 (N_14041,N_11081,N_10727);
or U14042 (N_14042,N_10080,N_9586);
or U14043 (N_14043,N_9136,N_11894);
xor U14044 (N_14044,N_9370,N_9098);
or U14045 (N_14045,N_10544,N_11039);
nand U14046 (N_14046,N_11330,N_11226);
nor U14047 (N_14047,N_10920,N_11057);
nor U14048 (N_14048,N_11058,N_9892);
or U14049 (N_14049,N_9708,N_11438);
or U14050 (N_14050,N_10577,N_10409);
nor U14051 (N_14051,N_10958,N_10906);
nand U14052 (N_14052,N_11119,N_9799);
nor U14053 (N_14053,N_11673,N_9553);
nand U14054 (N_14054,N_10488,N_9927);
nand U14055 (N_14055,N_9979,N_9263);
or U14056 (N_14056,N_10488,N_10405);
and U14057 (N_14057,N_11373,N_9271);
or U14058 (N_14058,N_11168,N_10514);
and U14059 (N_14059,N_11201,N_11977);
and U14060 (N_14060,N_11772,N_10469);
or U14061 (N_14061,N_10430,N_10208);
nor U14062 (N_14062,N_11089,N_10438);
or U14063 (N_14063,N_9078,N_10150);
or U14064 (N_14064,N_11381,N_9213);
nand U14065 (N_14065,N_11161,N_11207);
nor U14066 (N_14066,N_9829,N_9641);
and U14067 (N_14067,N_9916,N_11385);
nor U14068 (N_14068,N_11404,N_11429);
or U14069 (N_14069,N_9620,N_9371);
and U14070 (N_14070,N_11427,N_11991);
nand U14071 (N_14071,N_10267,N_10414);
nor U14072 (N_14072,N_10287,N_11969);
or U14073 (N_14073,N_11874,N_9948);
nand U14074 (N_14074,N_11423,N_9968);
or U14075 (N_14075,N_9179,N_11682);
nand U14076 (N_14076,N_10829,N_11094);
nand U14077 (N_14077,N_11074,N_10296);
or U14078 (N_14078,N_9608,N_10316);
nor U14079 (N_14079,N_11574,N_10562);
nor U14080 (N_14080,N_11232,N_9138);
or U14081 (N_14081,N_9358,N_11844);
nand U14082 (N_14082,N_10193,N_10242);
nor U14083 (N_14083,N_10273,N_9748);
nand U14084 (N_14084,N_10579,N_9797);
nand U14085 (N_14085,N_11682,N_11292);
nor U14086 (N_14086,N_11830,N_10411);
nand U14087 (N_14087,N_11065,N_11806);
or U14088 (N_14088,N_11879,N_10748);
or U14089 (N_14089,N_9305,N_11048);
nor U14090 (N_14090,N_11448,N_11279);
nor U14091 (N_14091,N_11220,N_10199);
nor U14092 (N_14092,N_11977,N_9837);
nor U14093 (N_14093,N_10472,N_11973);
or U14094 (N_14094,N_10329,N_9711);
and U14095 (N_14095,N_11310,N_9322);
and U14096 (N_14096,N_10882,N_9733);
nand U14097 (N_14097,N_11456,N_10531);
or U14098 (N_14098,N_9754,N_10084);
and U14099 (N_14099,N_11935,N_11785);
nor U14100 (N_14100,N_9183,N_9592);
nand U14101 (N_14101,N_10497,N_10416);
nand U14102 (N_14102,N_11080,N_10547);
or U14103 (N_14103,N_9027,N_11562);
and U14104 (N_14104,N_10435,N_9842);
and U14105 (N_14105,N_11529,N_10617);
or U14106 (N_14106,N_9856,N_9651);
nand U14107 (N_14107,N_10893,N_10212);
nand U14108 (N_14108,N_11798,N_11232);
or U14109 (N_14109,N_11164,N_10223);
or U14110 (N_14110,N_9203,N_9063);
and U14111 (N_14111,N_10211,N_11905);
and U14112 (N_14112,N_11990,N_11136);
nand U14113 (N_14113,N_11096,N_9697);
or U14114 (N_14114,N_11128,N_9006);
nand U14115 (N_14115,N_10987,N_11788);
or U14116 (N_14116,N_11301,N_9062);
nor U14117 (N_14117,N_9675,N_9135);
and U14118 (N_14118,N_11667,N_10941);
and U14119 (N_14119,N_9864,N_11821);
or U14120 (N_14120,N_9467,N_11691);
nor U14121 (N_14121,N_10978,N_10899);
nor U14122 (N_14122,N_10228,N_9286);
nand U14123 (N_14123,N_11007,N_9458);
nor U14124 (N_14124,N_10516,N_9568);
nand U14125 (N_14125,N_9839,N_10293);
and U14126 (N_14126,N_11232,N_11317);
and U14127 (N_14127,N_10946,N_10612);
and U14128 (N_14128,N_11287,N_10676);
and U14129 (N_14129,N_11268,N_10740);
nand U14130 (N_14130,N_11744,N_11947);
nand U14131 (N_14131,N_9931,N_9281);
and U14132 (N_14132,N_9032,N_11406);
nor U14133 (N_14133,N_11031,N_11146);
or U14134 (N_14134,N_11320,N_10092);
or U14135 (N_14135,N_9918,N_11290);
or U14136 (N_14136,N_11853,N_10106);
and U14137 (N_14137,N_11926,N_9190);
nand U14138 (N_14138,N_10303,N_11492);
or U14139 (N_14139,N_10296,N_10408);
nor U14140 (N_14140,N_11363,N_11338);
nand U14141 (N_14141,N_10193,N_9315);
or U14142 (N_14142,N_9693,N_10723);
or U14143 (N_14143,N_11113,N_10801);
and U14144 (N_14144,N_10269,N_9942);
nand U14145 (N_14145,N_9405,N_11790);
nand U14146 (N_14146,N_11987,N_9454);
and U14147 (N_14147,N_9897,N_9890);
and U14148 (N_14148,N_10567,N_11595);
nor U14149 (N_14149,N_9097,N_10818);
or U14150 (N_14150,N_11353,N_9141);
and U14151 (N_14151,N_11118,N_9263);
and U14152 (N_14152,N_9902,N_9574);
nand U14153 (N_14153,N_10240,N_9157);
or U14154 (N_14154,N_9900,N_11872);
and U14155 (N_14155,N_11932,N_11666);
and U14156 (N_14156,N_9801,N_10573);
nand U14157 (N_14157,N_9587,N_9604);
nor U14158 (N_14158,N_11699,N_11125);
nand U14159 (N_14159,N_11033,N_9233);
nor U14160 (N_14160,N_9352,N_11931);
nand U14161 (N_14161,N_11128,N_11782);
nand U14162 (N_14162,N_10574,N_9694);
nand U14163 (N_14163,N_10199,N_10011);
and U14164 (N_14164,N_9960,N_9777);
or U14165 (N_14165,N_11361,N_10242);
and U14166 (N_14166,N_11443,N_9490);
nor U14167 (N_14167,N_10097,N_10264);
nand U14168 (N_14168,N_9313,N_10143);
nor U14169 (N_14169,N_11575,N_11314);
nor U14170 (N_14170,N_10065,N_11057);
nor U14171 (N_14171,N_9026,N_11585);
nor U14172 (N_14172,N_10656,N_10840);
and U14173 (N_14173,N_11778,N_10386);
and U14174 (N_14174,N_11959,N_10169);
nand U14175 (N_14175,N_9409,N_11414);
nor U14176 (N_14176,N_10882,N_10198);
and U14177 (N_14177,N_9909,N_11017);
nand U14178 (N_14178,N_10610,N_9929);
and U14179 (N_14179,N_11089,N_10648);
nand U14180 (N_14180,N_11155,N_9434);
nand U14181 (N_14181,N_9041,N_9251);
and U14182 (N_14182,N_9981,N_11092);
or U14183 (N_14183,N_9235,N_11436);
nand U14184 (N_14184,N_10897,N_9903);
nand U14185 (N_14185,N_11497,N_9699);
nand U14186 (N_14186,N_10636,N_9078);
and U14187 (N_14187,N_10014,N_11337);
nand U14188 (N_14188,N_9789,N_11989);
or U14189 (N_14189,N_9908,N_9230);
or U14190 (N_14190,N_11165,N_10536);
and U14191 (N_14191,N_11037,N_11934);
nand U14192 (N_14192,N_11543,N_10099);
nor U14193 (N_14193,N_9793,N_10883);
nand U14194 (N_14194,N_11260,N_10955);
and U14195 (N_14195,N_10800,N_9565);
nand U14196 (N_14196,N_11079,N_10227);
nor U14197 (N_14197,N_11290,N_10641);
or U14198 (N_14198,N_11809,N_10053);
and U14199 (N_14199,N_11424,N_9013);
and U14200 (N_14200,N_11511,N_10070);
and U14201 (N_14201,N_11515,N_11548);
nor U14202 (N_14202,N_9397,N_11408);
nand U14203 (N_14203,N_11817,N_9696);
or U14204 (N_14204,N_10583,N_10740);
or U14205 (N_14205,N_11118,N_9044);
or U14206 (N_14206,N_11494,N_11325);
nor U14207 (N_14207,N_10475,N_10347);
nand U14208 (N_14208,N_11941,N_11979);
nor U14209 (N_14209,N_11249,N_9051);
or U14210 (N_14210,N_9961,N_9057);
nor U14211 (N_14211,N_10799,N_9991);
and U14212 (N_14212,N_10905,N_11607);
nand U14213 (N_14213,N_10940,N_11097);
nor U14214 (N_14214,N_10522,N_11534);
and U14215 (N_14215,N_10042,N_9810);
nor U14216 (N_14216,N_11039,N_10006);
nand U14217 (N_14217,N_11150,N_11932);
or U14218 (N_14218,N_11036,N_10396);
and U14219 (N_14219,N_10029,N_9053);
nand U14220 (N_14220,N_9122,N_10074);
nand U14221 (N_14221,N_10449,N_9324);
nor U14222 (N_14222,N_9867,N_9511);
nand U14223 (N_14223,N_11577,N_11556);
nor U14224 (N_14224,N_10194,N_11689);
and U14225 (N_14225,N_9297,N_10244);
or U14226 (N_14226,N_10420,N_11567);
or U14227 (N_14227,N_11616,N_11994);
or U14228 (N_14228,N_9807,N_9870);
nor U14229 (N_14229,N_10746,N_11328);
and U14230 (N_14230,N_9595,N_11846);
nand U14231 (N_14231,N_9320,N_11019);
nand U14232 (N_14232,N_10206,N_10920);
and U14233 (N_14233,N_11794,N_9713);
or U14234 (N_14234,N_10343,N_11280);
and U14235 (N_14235,N_9404,N_11030);
nor U14236 (N_14236,N_9970,N_9652);
and U14237 (N_14237,N_10561,N_11962);
and U14238 (N_14238,N_9276,N_10044);
nor U14239 (N_14239,N_9831,N_10677);
nor U14240 (N_14240,N_11688,N_11651);
nand U14241 (N_14241,N_10074,N_9986);
nor U14242 (N_14242,N_11384,N_9901);
and U14243 (N_14243,N_10482,N_10633);
or U14244 (N_14244,N_10321,N_10898);
nor U14245 (N_14245,N_9147,N_9960);
nor U14246 (N_14246,N_9804,N_10473);
nand U14247 (N_14247,N_11753,N_11106);
and U14248 (N_14248,N_11764,N_10449);
nor U14249 (N_14249,N_9843,N_9409);
nor U14250 (N_14250,N_10515,N_11622);
or U14251 (N_14251,N_11516,N_11678);
and U14252 (N_14252,N_10597,N_9644);
and U14253 (N_14253,N_11618,N_10138);
nor U14254 (N_14254,N_9997,N_9838);
nand U14255 (N_14255,N_11790,N_9991);
and U14256 (N_14256,N_9199,N_9597);
nand U14257 (N_14257,N_10688,N_9357);
nand U14258 (N_14258,N_9399,N_11153);
and U14259 (N_14259,N_9900,N_9520);
or U14260 (N_14260,N_11523,N_10677);
nor U14261 (N_14261,N_11857,N_10810);
nand U14262 (N_14262,N_10458,N_9608);
or U14263 (N_14263,N_10856,N_10195);
nor U14264 (N_14264,N_9452,N_11307);
nor U14265 (N_14265,N_9204,N_11419);
nand U14266 (N_14266,N_11551,N_10865);
and U14267 (N_14267,N_9275,N_11445);
or U14268 (N_14268,N_10949,N_11221);
nor U14269 (N_14269,N_9149,N_10313);
and U14270 (N_14270,N_9243,N_10389);
nand U14271 (N_14271,N_10110,N_9309);
and U14272 (N_14272,N_11670,N_11843);
xor U14273 (N_14273,N_10020,N_9437);
or U14274 (N_14274,N_9864,N_9428);
or U14275 (N_14275,N_11472,N_9730);
nand U14276 (N_14276,N_11381,N_11713);
or U14277 (N_14277,N_11086,N_9996);
nor U14278 (N_14278,N_9098,N_11183);
nand U14279 (N_14279,N_11841,N_9070);
nand U14280 (N_14280,N_9071,N_10819);
and U14281 (N_14281,N_9583,N_10842);
nand U14282 (N_14282,N_11795,N_11934);
or U14283 (N_14283,N_10225,N_10767);
nand U14284 (N_14284,N_9537,N_9777);
or U14285 (N_14285,N_9306,N_9842);
and U14286 (N_14286,N_10134,N_9049);
nand U14287 (N_14287,N_10330,N_10661);
nor U14288 (N_14288,N_9006,N_10651);
or U14289 (N_14289,N_10162,N_11891);
or U14290 (N_14290,N_10251,N_11260);
or U14291 (N_14291,N_9666,N_10162);
or U14292 (N_14292,N_11418,N_11158);
nor U14293 (N_14293,N_11150,N_9921);
nor U14294 (N_14294,N_11829,N_11060);
or U14295 (N_14295,N_10048,N_10648);
nor U14296 (N_14296,N_10828,N_10833);
nand U14297 (N_14297,N_10308,N_11594);
nand U14298 (N_14298,N_9945,N_11270);
nand U14299 (N_14299,N_10383,N_9906);
nor U14300 (N_14300,N_11846,N_10387);
nor U14301 (N_14301,N_9002,N_10253);
or U14302 (N_14302,N_10796,N_11680);
nand U14303 (N_14303,N_9445,N_11270);
and U14304 (N_14304,N_9914,N_9600);
and U14305 (N_14305,N_11027,N_9316);
xnor U14306 (N_14306,N_10235,N_9430);
nand U14307 (N_14307,N_10999,N_9262);
and U14308 (N_14308,N_10756,N_10250);
nand U14309 (N_14309,N_10183,N_11349);
nand U14310 (N_14310,N_9547,N_10193);
and U14311 (N_14311,N_9655,N_11978);
and U14312 (N_14312,N_10486,N_10282);
and U14313 (N_14313,N_11108,N_10006);
nor U14314 (N_14314,N_9431,N_9341);
or U14315 (N_14315,N_11736,N_11935);
nand U14316 (N_14316,N_11675,N_11511);
nand U14317 (N_14317,N_10204,N_11925);
xnor U14318 (N_14318,N_11280,N_11809);
nand U14319 (N_14319,N_11288,N_9433);
or U14320 (N_14320,N_11651,N_10473);
or U14321 (N_14321,N_11804,N_9146);
or U14322 (N_14322,N_10590,N_9574);
and U14323 (N_14323,N_10582,N_9091);
nand U14324 (N_14324,N_9761,N_10209);
nand U14325 (N_14325,N_9217,N_11652);
nor U14326 (N_14326,N_11708,N_9646);
or U14327 (N_14327,N_10077,N_10148);
or U14328 (N_14328,N_10925,N_11051);
and U14329 (N_14329,N_9601,N_10878);
nand U14330 (N_14330,N_11447,N_10271);
nor U14331 (N_14331,N_10059,N_9821);
and U14332 (N_14332,N_11451,N_9120);
nor U14333 (N_14333,N_11629,N_11511);
nand U14334 (N_14334,N_11737,N_9479);
or U14335 (N_14335,N_11981,N_10525);
or U14336 (N_14336,N_10864,N_11765);
nor U14337 (N_14337,N_10122,N_9002);
or U14338 (N_14338,N_9673,N_10049);
and U14339 (N_14339,N_9478,N_11155);
and U14340 (N_14340,N_9530,N_10488);
or U14341 (N_14341,N_11690,N_10930);
and U14342 (N_14342,N_10554,N_11543);
or U14343 (N_14343,N_9269,N_10890);
nand U14344 (N_14344,N_11078,N_10095);
and U14345 (N_14345,N_10043,N_11917);
nand U14346 (N_14346,N_10777,N_10853);
nand U14347 (N_14347,N_11982,N_11981);
and U14348 (N_14348,N_9762,N_9496);
and U14349 (N_14349,N_9532,N_9286);
nand U14350 (N_14350,N_9389,N_9091);
nor U14351 (N_14351,N_10272,N_11411);
or U14352 (N_14352,N_11089,N_10510);
nor U14353 (N_14353,N_10673,N_9090);
nor U14354 (N_14354,N_9371,N_11604);
nand U14355 (N_14355,N_11700,N_10352);
nor U14356 (N_14356,N_9524,N_9429);
and U14357 (N_14357,N_10219,N_9312);
xnor U14358 (N_14358,N_9069,N_10277);
nand U14359 (N_14359,N_10295,N_11123);
nand U14360 (N_14360,N_10231,N_10598);
nand U14361 (N_14361,N_11842,N_9190);
and U14362 (N_14362,N_9884,N_11655);
and U14363 (N_14363,N_10460,N_9799);
and U14364 (N_14364,N_10018,N_11065);
xnor U14365 (N_14365,N_9080,N_9614);
nor U14366 (N_14366,N_11870,N_11077);
or U14367 (N_14367,N_11658,N_10882);
and U14368 (N_14368,N_9396,N_11968);
nand U14369 (N_14369,N_10674,N_9442);
nand U14370 (N_14370,N_11424,N_10932);
and U14371 (N_14371,N_9964,N_10285);
nand U14372 (N_14372,N_10940,N_10975);
nand U14373 (N_14373,N_11196,N_9532);
or U14374 (N_14374,N_9609,N_9578);
or U14375 (N_14375,N_10228,N_11143);
or U14376 (N_14376,N_9022,N_10607);
nor U14377 (N_14377,N_10900,N_9806);
nor U14378 (N_14378,N_10553,N_11208);
or U14379 (N_14379,N_11041,N_11390);
nor U14380 (N_14380,N_9445,N_10198);
and U14381 (N_14381,N_10815,N_11303);
nand U14382 (N_14382,N_11835,N_10663);
nand U14383 (N_14383,N_9530,N_9799);
nand U14384 (N_14384,N_9292,N_11582);
nor U14385 (N_14385,N_9708,N_11896);
and U14386 (N_14386,N_9069,N_11712);
nand U14387 (N_14387,N_11873,N_10687);
or U14388 (N_14388,N_9976,N_10985);
and U14389 (N_14389,N_9718,N_11565);
or U14390 (N_14390,N_9252,N_10563);
nor U14391 (N_14391,N_11344,N_10437);
and U14392 (N_14392,N_11037,N_10494);
or U14393 (N_14393,N_10794,N_9957);
nor U14394 (N_14394,N_11262,N_11614);
nor U14395 (N_14395,N_11333,N_11561);
nand U14396 (N_14396,N_11690,N_10803);
nor U14397 (N_14397,N_10578,N_10633);
nor U14398 (N_14398,N_11264,N_11705);
nand U14399 (N_14399,N_9399,N_11686);
nand U14400 (N_14400,N_10924,N_10343);
nand U14401 (N_14401,N_9249,N_9711);
and U14402 (N_14402,N_9232,N_10965);
or U14403 (N_14403,N_11709,N_10826);
nand U14404 (N_14404,N_9016,N_11875);
and U14405 (N_14405,N_10046,N_9962);
or U14406 (N_14406,N_11746,N_10711);
xor U14407 (N_14407,N_10442,N_10237);
nor U14408 (N_14408,N_11632,N_10884);
nand U14409 (N_14409,N_10067,N_9722);
nor U14410 (N_14410,N_11763,N_9578);
xnor U14411 (N_14411,N_11569,N_11982);
or U14412 (N_14412,N_11334,N_11859);
nand U14413 (N_14413,N_11865,N_10667);
or U14414 (N_14414,N_10257,N_10423);
nor U14415 (N_14415,N_11465,N_9272);
nor U14416 (N_14416,N_11379,N_10798);
or U14417 (N_14417,N_10743,N_10004);
nand U14418 (N_14418,N_9797,N_10896);
nor U14419 (N_14419,N_10971,N_10312);
or U14420 (N_14420,N_10365,N_9507);
and U14421 (N_14421,N_11361,N_11966);
nand U14422 (N_14422,N_9511,N_11362);
and U14423 (N_14423,N_10332,N_11065);
or U14424 (N_14424,N_11137,N_10448);
and U14425 (N_14425,N_11100,N_9004);
nor U14426 (N_14426,N_10900,N_9969);
and U14427 (N_14427,N_11543,N_9634);
nor U14428 (N_14428,N_11039,N_9191);
nand U14429 (N_14429,N_9168,N_9810);
nand U14430 (N_14430,N_9103,N_10398);
nor U14431 (N_14431,N_9753,N_9349);
and U14432 (N_14432,N_9713,N_10891);
or U14433 (N_14433,N_9821,N_9626);
and U14434 (N_14434,N_11204,N_11485);
nand U14435 (N_14435,N_11968,N_9239);
and U14436 (N_14436,N_9207,N_9719);
nand U14437 (N_14437,N_10988,N_9161);
nand U14438 (N_14438,N_10004,N_10864);
and U14439 (N_14439,N_11197,N_10924);
or U14440 (N_14440,N_10571,N_9206);
and U14441 (N_14441,N_9012,N_10253);
nor U14442 (N_14442,N_9029,N_10205);
nand U14443 (N_14443,N_9456,N_10730);
nor U14444 (N_14444,N_11242,N_9089);
and U14445 (N_14445,N_9097,N_9088);
nand U14446 (N_14446,N_10877,N_10133);
and U14447 (N_14447,N_10193,N_10422);
nand U14448 (N_14448,N_9905,N_10863);
or U14449 (N_14449,N_11530,N_9645);
nor U14450 (N_14450,N_9592,N_11407);
nand U14451 (N_14451,N_9708,N_11385);
nand U14452 (N_14452,N_11911,N_11418);
or U14453 (N_14453,N_11087,N_9554);
or U14454 (N_14454,N_9703,N_9170);
nand U14455 (N_14455,N_11383,N_11182);
nand U14456 (N_14456,N_9448,N_10124);
nand U14457 (N_14457,N_9550,N_9980);
nor U14458 (N_14458,N_11274,N_10834);
and U14459 (N_14459,N_10757,N_9771);
or U14460 (N_14460,N_10049,N_10980);
nand U14461 (N_14461,N_11160,N_10218);
or U14462 (N_14462,N_11894,N_11999);
nand U14463 (N_14463,N_10217,N_9109);
and U14464 (N_14464,N_11810,N_10319);
and U14465 (N_14465,N_9307,N_11213);
or U14466 (N_14466,N_11850,N_10951);
nor U14467 (N_14467,N_10036,N_10789);
nand U14468 (N_14468,N_11870,N_10200);
nand U14469 (N_14469,N_11628,N_10247);
or U14470 (N_14470,N_10182,N_11197);
and U14471 (N_14471,N_9356,N_11005);
and U14472 (N_14472,N_9029,N_9980);
nor U14473 (N_14473,N_9466,N_10608);
or U14474 (N_14474,N_11083,N_11370);
and U14475 (N_14475,N_11330,N_9612);
nand U14476 (N_14476,N_9657,N_10473);
nand U14477 (N_14477,N_10570,N_11688);
nor U14478 (N_14478,N_11764,N_10731);
nand U14479 (N_14479,N_10802,N_11013);
or U14480 (N_14480,N_9752,N_9329);
or U14481 (N_14481,N_10582,N_10862);
nand U14482 (N_14482,N_9058,N_10650);
or U14483 (N_14483,N_11729,N_9065);
nand U14484 (N_14484,N_9646,N_11616);
or U14485 (N_14485,N_10099,N_9000);
or U14486 (N_14486,N_11423,N_9055);
or U14487 (N_14487,N_11533,N_9635);
nand U14488 (N_14488,N_11158,N_11377);
or U14489 (N_14489,N_11024,N_11427);
and U14490 (N_14490,N_10824,N_11144);
nor U14491 (N_14491,N_9182,N_9991);
nor U14492 (N_14492,N_11441,N_11126);
or U14493 (N_14493,N_10615,N_11371);
or U14494 (N_14494,N_10787,N_10623);
and U14495 (N_14495,N_9462,N_11334);
nand U14496 (N_14496,N_11676,N_10905);
nand U14497 (N_14497,N_11583,N_11250);
or U14498 (N_14498,N_9814,N_10085);
nor U14499 (N_14499,N_10253,N_11669);
nor U14500 (N_14500,N_9409,N_11925);
or U14501 (N_14501,N_9214,N_9189);
nand U14502 (N_14502,N_10223,N_9585);
or U14503 (N_14503,N_9556,N_10924);
nor U14504 (N_14504,N_10007,N_10051);
nand U14505 (N_14505,N_9960,N_10021);
xnor U14506 (N_14506,N_11320,N_9550);
nor U14507 (N_14507,N_10294,N_9880);
nor U14508 (N_14508,N_10193,N_10861);
and U14509 (N_14509,N_11917,N_11077);
and U14510 (N_14510,N_11330,N_9350);
or U14511 (N_14511,N_9157,N_10962);
nand U14512 (N_14512,N_9677,N_10318);
or U14513 (N_14513,N_9951,N_9748);
nand U14514 (N_14514,N_9871,N_9284);
nor U14515 (N_14515,N_11705,N_11348);
or U14516 (N_14516,N_10596,N_10094);
and U14517 (N_14517,N_9894,N_10398);
or U14518 (N_14518,N_9735,N_10673);
nand U14519 (N_14519,N_10932,N_9260);
or U14520 (N_14520,N_9336,N_10520);
nor U14521 (N_14521,N_9119,N_10273);
and U14522 (N_14522,N_10109,N_11718);
or U14523 (N_14523,N_11126,N_11266);
or U14524 (N_14524,N_11945,N_9241);
nor U14525 (N_14525,N_10718,N_10691);
nand U14526 (N_14526,N_10979,N_11483);
or U14527 (N_14527,N_10912,N_10507);
nand U14528 (N_14528,N_11292,N_10067);
nand U14529 (N_14529,N_10951,N_11733);
xor U14530 (N_14530,N_11010,N_11442);
nand U14531 (N_14531,N_9225,N_10220);
and U14532 (N_14532,N_11020,N_11927);
or U14533 (N_14533,N_9576,N_10069);
and U14534 (N_14534,N_10420,N_11944);
nor U14535 (N_14535,N_10173,N_10101);
nand U14536 (N_14536,N_11468,N_11906);
or U14537 (N_14537,N_10666,N_11265);
and U14538 (N_14538,N_11429,N_9865);
nand U14539 (N_14539,N_10572,N_9070);
and U14540 (N_14540,N_9302,N_9030);
nor U14541 (N_14541,N_10777,N_11147);
and U14542 (N_14542,N_10650,N_11329);
nor U14543 (N_14543,N_10872,N_11200);
or U14544 (N_14544,N_10420,N_11176);
and U14545 (N_14545,N_9758,N_10533);
or U14546 (N_14546,N_11082,N_9944);
and U14547 (N_14547,N_9693,N_9349);
or U14548 (N_14548,N_11971,N_9436);
nand U14549 (N_14549,N_11717,N_11147);
or U14550 (N_14550,N_10416,N_11869);
or U14551 (N_14551,N_11126,N_9592);
nand U14552 (N_14552,N_10536,N_10598);
nor U14553 (N_14553,N_9753,N_11064);
nand U14554 (N_14554,N_11157,N_9628);
nor U14555 (N_14555,N_10795,N_9879);
nand U14556 (N_14556,N_9028,N_11767);
nor U14557 (N_14557,N_10082,N_9765);
nor U14558 (N_14558,N_11890,N_11478);
nand U14559 (N_14559,N_10165,N_10147);
nand U14560 (N_14560,N_9733,N_9729);
nor U14561 (N_14561,N_11474,N_11427);
and U14562 (N_14562,N_9824,N_9847);
nor U14563 (N_14563,N_11915,N_9708);
or U14564 (N_14564,N_10587,N_11187);
nand U14565 (N_14565,N_9117,N_11653);
and U14566 (N_14566,N_9527,N_9750);
nor U14567 (N_14567,N_9575,N_9184);
or U14568 (N_14568,N_9357,N_10693);
or U14569 (N_14569,N_10695,N_9138);
nor U14570 (N_14570,N_11123,N_10417);
and U14571 (N_14571,N_9241,N_10692);
nand U14572 (N_14572,N_9155,N_11740);
and U14573 (N_14573,N_10375,N_11343);
nand U14574 (N_14574,N_9180,N_10568);
and U14575 (N_14575,N_10417,N_9058);
and U14576 (N_14576,N_11413,N_9895);
nand U14577 (N_14577,N_9386,N_11697);
nand U14578 (N_14578,N_10075,N_11714);
and U14579 (N_14579,N_11444,N_9599);
and U14580 (N_14580,N_10766,N_10633);
or U14581 (N_14581,N_9489,N_10406);
nor U14582 (N_14582,N_11647,N_11491);
and U14583 (N_14583,N_10310,N_9815);
and U14584 (N_14584,N_9217,N_11748);
nor U14585 (N_14585,N_9800,N_11076);
or U14586 (N_14586,N_9236,N_11584);
nor U14587 (N_14587,N_10951,N_9343);
nor U14588 (N_14588,N_11855,N_10267);
and U14589 (N_14589,N_11756,N_10172);
nand U14590 (N_14590,N_10202,N_10327);
nand U14591 (N_14591,N_9538,N_11720);
xnor U14592 (N_14592,N_9778,N_11160);
or U14593 (N_14593,N_11735,N_9029);
nor U14594 (N_14594,N_11422,N_10232);
nor U14595 (N_14595,N_11373,N_10739);
nand U14596 (N_14596,N_9120,N_10909);
nand U14597 (N_14597,N_11110,N_10250);
nor U14598 (N_14598,N_11841,N_9971);
nand U14599 (N_14599,N_9541,N_10546);
nand U14600 (N_14600,N_9706,N_9608);
xor U14601 (N_14601,N_10758,N_10254);
nand U14602 (N_14602,N_9209,N_11695);
nor U14603 (N_14603,N_9264,N_11619);
nand U14604 (N_14604,N_10308,N_9374);
nor U14605 (N_14605,N_10335,N_9292);
or U14606 (N_14606,N_10131,N_9849);
or U14607 (N_14607,N_10829,N_11054);
and U14608 (N_14608,N_11686,N_9753);
and U14609 (N_14609,N_11782,N_9291);
nor U14610 (N_14610,N_11920,N_9173);
and U14611 (N_14611,N_10159,N_11446);
nor U14612 (N_14612,N_9197,N_9490);
and U14613 (N_14613,N_10069,N_11772);
or U14614 (N_14614,N_9499,N_10225);
or U14615 (N_14615,N_10455,N_11284);
or U14616 (N_14616,N_11335,N_10114);
and U14617 (N_14617,N_10389,N_9554);
and U14618 (N_14618,N_11531,N_11627);
and U14619 (N_14619,N_11487,N_9973);
nor U14620 (N_14620,N_9570,N_11442);
nand U14621 (N_14621,N_9245,N_9472);
or U14622 (N_14622,N_10790,N_9596);
and U14623 (N_14623,N_11706,N_11116);
nor U14624 (N_14624,N_11609,N_10220);
or U14625 (N_14625,N_9657,N_10878);
nand U14626 (N_14626,N_9704,N_9782);
nand U14627 (N_14627,N_9648,N_11793);
nor U14628 (N_14628,N_10956,N_9461);
or U14629 (N_14629,N_10022,N_9476);
or U14630 (N_14630,N_11434,N_9403);
and U14631 (N_14631,N_10517,N_9690);
nand U14632 (N_14632,N_10441,N_10427);
or U14633 (N_14633,N_11166,N_9656);
nand U14634 (N_14634,N_10554,N_11259);
nor U14635 (N_14635,N_10748,N_10736);
nand U14636 (N_14636,N_10208,N_11765);
nor U14637 (N_14637,N_11697,N_9724);
nor U14638 (N_14638,N_11623,N_11021);
and U14639 (N_14639,N_9138,N_10258);
or U14640 (N_14640,N_11492,N_10085);
nor U14641 (N_14641,N_10600,N_11318);
or U14642 (N_14642,N_11966,N_10400);
nand U14643 (N_14643,N_11923,N_10505);
or U14644 (N_14644,N_11847,N_10560);
or U14645 (N_14645,N_9083,N_9639);
or U14646 (N_14646,N_11212,N_11677);
or U14647 (N_14647,N_10399,N_10742);
and U14648 (N_14648,N_9962,N_11347);
nor U14649 (N_14649,N_10384,N_9094);
and U14650 (N_14650,N_9774,N_11229);
and U14651 (N_14651,N_9984,N_10817);
or U14652 (N_14652,N_10426,N_10329);
or U14653 (N_14653,N_9806,N_9395);
or U14654 (N_14654,N_9788,N_11776);
nand U14655 (N_14655,N_10092,N_9306);
or U14656 (N_14656,N_9067,N_10108);
nor U14657 (N_14657,N_10027,N_11295);
nand U14658 (N_14658,N_11944,N_10613);
nand U14659 (N_14659,N_11729,N_11637);
or U14660 (N_14660,N_9459,N_10270);
nor U14661 (N_14661,N_9981,N_11547);
or U14662 (N_14662,N_10984,N_11860);
nand U14663 (N_14663,N_9675,N_10407);
nor U14664 (N_14664,N_11569,N_9690);
nor U14665 (N_14665,N_10304,N_9505);
nor U14666 (N_14666,N_11887,N_9832);
and U14667 (N_14667,N_10751,N_11353);
nand U14668 (N_14668,N_9794,N_9285);
nand U14669 (N_14669,N_10022,N_11852);
and U14670 (N_14670,N_9604,N_10701);
nand U14671 (N_14671,N_10499,N_11681);
nand U14672 (N_14672,N_9366,N_9123);
nor U14673 (N_14673,N_11163,N_11002);
nor U14674 (N_14674,N_11493,N_10029);
nor U14675 (N_14675,N_10192,N_9600);
nor U14676 (N_14676,N_10658,N_9284);
nand U14677 (N_14677,N_11216,N_11327);
and U14678 (N_14678,N_9549,N_9778);
nand U14679 (N_14679,N_11860,N_10620);
nand U14680 (N_14680,N_11561,N_11087);
and U14681 (N_14681,N_9586,N_9321);
and U14682 (N_14682,N_10874,N_11565);
nor U14683 (N_14683,N_9650,N_11550);
nor U14684 (N_14684,N_11507,N_9256);
nor U14685 (N_14685,N_11681,N_11806);
or U14686 (N_14686,N_10617,N_10793);
nand U14687 (N_14687,N_9603,N_10790);
nor U14688 (N_14688,N_10144,N_11095);
and U14689 (N_14689,N_9298,N_11889);
nand U14690 (N_14690,N_11620,N_10771);
and U14691 (N_14691,N_10969,N_11462);
and U14692 (N_14692,N_9003,N_9203);
or U14693 (N_14693,N_11800,N_11312);
nor U14694 (N_14694,N_11681,N_10216);
nor U14695 (N_14695,N_9673,N_10692);
or U14696 (N_14696,N_9686,N_10113);
nand U14697 (N_14697,N_9870,N_9177);
nor U14698 (N_14698,N_11486,N_10743);
nor U14699 (N_14699,N_10126,N_11909);
and U14700 (N_14700,N_9162,N_9689);
nand U14701 (N_14701,N_11378,N_9967);
and U14702 (N_14702,N_10467,N_11445);
nor U14703 (N_14703,N_10323,N_11499);
or U14704 (N_14704,N_9101,N_9807);
nor U14705 (N_14705,N_11790,N_11822);
nor U14706 (N_14706,N_9794,N_9885);
nand U14707 (N_14707,N_9794,N_11580);
and U14708 (N_14708,N_9806,N_11797);
or U14709 (N_14709,N_9289,N_10040);
nand U14710 (N_14710,N_10443,N_10798);
and U14711 (N_14711,N_9469,N_10164);
nand U14712 (N_14712,N_10831,N_10815);
or U14713 (N_14713,N_11911,N_9408);
nor U14714 (N_14714,N_9042,N_9556);
nand U14715 (N_14715,N_11993,N_10177);
nand U14716 (N_14716,N_9433,N_10982);
and U14717 (N_14717,N_11536,N_10693);
xor U14718 (N_14718,N_10947,N_9488);
nand U14719 (N_14719,N_10587,N_10974);
nand U14720 (N_14720,N_10791,N_10091);
nand U14721 (N_14721,N_10412,N_9253);
nor U14722 (N_14722,N_10031,N_11239);
nor U14723 (N_14723,N_11623,N_11353);
nor U14724 (N_14724,N_10873,N_11702);
or U14725 (N_14725,N_10634,N_11986);
nand U14726 (N_14726,N_10769,N_9462);
or U14727 (N_14727,N_11715,N_11920);
and U14728 (N_14728,N_11473,N_10318);
nor U14729 (N_14729,N_11336,N_11881);
nor U14730 (N_14730,N_9522,N_11636);
or U14731 (N_14731,N_9196,N_10084);
nor U14732 (N_14732,N_11370,N_9403);
nand U14733 (N_14733,N_10682,N_11111);
or U14734 (N_14734,N_11103,N_9147);
nor U14735 (N_14735,N_9907,N_9925);
or U14736 (N_14736,N_11338,N_10246);
nor U14737 (N_14737,N_10261,N_11913);
nand U14738 (N_14738,N_10506,N_11323);
nand U14739 (N_14739,N_9695,N_10192);
nand U14740 (N_14740,N_11381,N_9440);
nor U14741 (N_14741,N_10562,N_10246);
nand U14742 (N_14742,N_9482,N_11355);
or U14743 (N_14743,N_11750,N_9377);
nor U14744 (N_14744,N_9424,N_10292);
nor U14745 (N_14745,N_9804,N_10019);
and U14746 (N_14746,N_9070,N_10463);
and U14747 (N_14747,N_10932,N_11577);
nor U14748 (N_14748,N_9915,N_11849);
nand U14749 (N_14749,N_9265,N_11864);
nor U14750 (N_14750,N_10976,N_10176);
or U14751 (N_14751,N_9774,N_9808);
and U14752 (N_14752,N_9746,N_11510);
or U14753 (N_14753,N_11095,N_9022);
nor U14754 (N_14754,N_11164,N_11807);
xnor U14755 (N_14755,N_9434,N_11556);
or U14756 (N_14756,N_11859,N_9452);
nand U14757 (N_14757,N_10564,N_10546);
nor U14758 (N_14758,N_9196,N_9507);
or U14759 (N_14759,N_11491,N_11985);
and U14760 (N_14760,N_11661,N_10200);
or U14761 (N_14761,N_11557,N_11461);
and U14762 (N_14762,N_9672,N_11361);
nand U14763 (N_14763,N_9443,N_10676);
nand U14764 (N_14764,N_9447,N_11742);
nand U14765 (N_14765,N_11458,N_10835);
nand U14766 (N_14766,N_9590,N_9855);
or U14767 (N_14767,N_10034,N_10769);
and U14768 (N_14768,N_11536,N_11918);
nor U14769 (N_14769,N_9227,N_10392);
nand U14770 (N_14770,N_11335,N_9586);
nand U14771 (N_14771,N_9364,N_10240);
nand U14772 (N_14772,N_9264,N_11484);
nand U14773 (N_14773,N_10127,N_10659);
nand U14774 (N_14774,N_11182,N_10593);
nor U14775 (N_14775,N_11532,N_10837);
nand U14776 (N_14776,N_10558,N_9201);
nand U14777 (N_14777,N_10397,N_10347);
or U14778 (N_14778,N_11435,N_10565);
nor U14779 (N_14779,N_11476,N_11114);
or U14780 (N_14780,N_10696,N_9345);
xnor U14781 (N_14781,N_10516,N_10561);
nor U14782 (N_14782,N_11396,N_9741);
xor U14783 (N_14783,N_9215,N_9312);
nor U14784 (N_14784,N_9011,N_11545);
or U14785 (N_14785,N_10970,N_10881);
and U14786 (N_14786,N_9565,N_11054);
nand U14787 (N_14787,N_11187,N_9142);
nor U14788 (N_14788,N_11567,N_11394);
or U14789 (N_14789,N_11766,N_10287);
or U14790 (N_14790,N_11544,N_11882);
and U14791 (N_14791,N_11425,N_11289);
xnor U14792 (N_14792,N_10459,N_10219);
or U14793 (N_14793,N_10042,N_9989);
nor U14794 (N_14794,N_11933,N_10472);
nand U14795 (N_14795,N_10216,N_10000);
nor U14796 (N_14796,N_11397,N_11844);
xnor U14797 (N_14797,N_9809,N_11988);
nand U14798 (N_14798,N_10996,N_10911);
or U14799 (N_14799,N_11267,N_10531);
nand U14800 (N_14800,N_9568,N_11842);
or U14801 (N_14801,N_11005,N_9304);
nor U14802 (N_14802,N_9248,N_11443);
nand U14803 (N_14803,N_9436,N_11152);
and U14804 (N_14804,N_9305,N_9875);
and U14805 (N_14805,N_10168,N_11502);
and U14806 (N_14806,N_11192,N_11018);
and U14807 (N_14807,N_9290,N_11008);
or U14808 (N_14808,N_11527,N_10785);
or U14809 (N_14809,N_10150,N_10766);
or U14810 (N_14810,N_9032,N_10574);
nor U14811 (N_14811,N_11934,N_10694);
or U14812 (N_14812,N_10811,N_11031);
and U14813 (N_14813,N_11683,N_11874);
or U14814 (N_14814,N_11981,N_9316);
nand U14815 (N_14815,N_9118,N_10234);
nor U14816 (N_14816,N_9088,N_9851);
or U14817 (N_14817,N_11738,N_11508);
nand U14818 (N_14818,N_11346,N_11307);
and U14819 (N_14819,N_9923,N_11071);
or U14820 (N_14820,N_11769,N_9751);
nor U14821 (N_14821,N_11629,N_9890);
or U14822 (N_14822,N_10466,N_11524);
nor U14823 (N_14823,N_10848,N_9175);
and U14824 (N_14824,N_10220,N_9116);
nor U14825 (N_14825,N_11283,N_9855);
and U14826 (N_14826,N_10242,N_9901);
nor U14827 (N_14827,N_11572,N_11064);
nand U14828 (N_14828,N_11550,N_11352);
xor U14829 (N_14829,N_10027,N_11481);
and U14830 (N_14830,N_10446,N_10674);
nor U14831 (N_14831,N_11515,N_10103);
and U14832 (N_14832,N_11757,N_10447);
nand U14833 (N_14833,N_11015,N_9201);
nor U14834 (N_14834,N_11953,N_10627);
and U14835 (N_14835,N_11729,N_11951);
and U14836 (N_14836,N_11634,N_11014);
or U14837 (N_14837,N_9154,N_9793);
nor U14838 (N_14838,N_11618,N_10066);
and U14839 (N_14839,N_11884,N_11162);
nor U14840 (N_14840,N_11482,N_10598);
nor U14841 (N_14841,N_10346,N_10652);
and U14842 (N_14842,N_10650,N_11836);
or U14843 (N_14843,N_11938,N_11976);
nor U14844 (N_14844,N_9323,N_10905);
nand U14845 (N_14845,N_9172,N_10659);
nor U14846 (N_14846,N_10326,N_9220);
nand U14847 (N_14847,N_10003,N_9015);
or U14848 (N_14848,N_9535,N_9235);
or U14849 (N_14849,N_9235,N_11474);
nand U14850 (N_14850,N_10021,N_11028);
nand U14851 (N_14851,N_10514,N_11070);
and U14852 (N_14852,N_11982,N_10118);
or U14853 (N_14853,N_10608,N_9539);
nor U14854 (N_14854,N_11763,N_9528);
or U14855 (N_14855,N_9368,N_11737);
or U14856 (N_14856,N_9244,N_9527);
nand U14857 (N_14857,N_9447,N_10857);
nor U14858 (N_14858,N_10732,N_9219);
nand U14859 (N_14859,N_11499,N_9886);
and U14860 (N_14860,N_9468,N_9484);
or U14861 (N_14861,N_9465,N_11698);
nor U14862 (N_14862,N_10810,N_10661);
nand U14863 (N_14863,N_11408,N_9455);
nor U14864 (N_14864,N_11195,N_10861);
and U14865 (N_14865,N_9093,N_9770);
nand U14866 (N_14866,N_10277,N_10699);
xor U14867 (N_14867,N_11962,N_10044);
nand U14868 (N_14868,N_11243,N_11383);
and U14869 (N_14869,N_11943,N_9486);
and U14870 (N_14870,N_11223,N_10487);
or U14871 (N_14871,N_10768,N_10570);
or U14872 (N_14872,N_9709,N_9599);
nor U14873 (N_14873,N_11747,N_11091);
nor U14874 (N_14874,N_9392,N_10456);
nor U14875 (N_14875,N_11980,N_9244);
nor U14876 (N_14876,N_11555,N_11002);
nor U14877 (N_14877,N_9475,N_11065);
nand U14878 (N_14878,N_10295,N_10100);
or U14879 (N_14879,N_9207,N_9605);
and U14880 (N_14880,N_11722,N_11623);
nor U14881 (N_14881,N_11846,N_9496);
nand U14882 (N_14882,N_10367,N_9104);
nor U14883 (N_14883,N_11833,N_10148);
or U14884 (N_14884,N_11621,N_10672);
and U14885 (N_14885,N_10824,N_10507);
or U14886 (N_14886,N_11994,N_11379);
and U14887 (N_14887,N_10680,N_10002);
and U14888 (N_14888,N_10726,N_9718);
and U14889 (N_14889,N_11177,N_10278);
nor U14890 (N_14890,N_10920,N_9524);
and U14891 (N_14891,N_9962,N_10201);
nor U14892 (N_14892,N_9512,N_9819);
nand U14893 (N_14893,N_10567,N_10281);
or U14894 (N_14894,N_10388,N_10971);
nand U14895 (N_14895,N_10923,N_10397);
nor U14896 (N_14896,N_10089,N_9049);
nor U14897 (N_14897,N_11766,N_11187);
nand U14898 (N_14898,N_9730,N_11131);
nand U14899 (N_14899,N_10243,N_9410);
or U14900 (N_14900,N_10078,N_10502);
and U14901 (N_14901,N_11307,N_11856);
and U14902 (N_14902,N_10916,N_10754);
and U14903 (N_14903,N_9926,N_9131);
and U14904 (N_14904,N_9255,N_10376);
nand U14905 (N_14905,N_10773,N_9992);
xnor U14906 (N_14906,N_10165,N_10175);
or U14907 (N_14907,N_10495,N_9556);
nor U14908 (N_14908,N_10897,N_9199);
or U14909 (N_14909,N_9218,N_10946);
and U14910 (N_14910,N_11781,N_10497);
nor U14911 (N_14911,N_10177,N_10274);
or U14912 (N_14912,N_11662,N_11098);
or U14913 (N_14913,N_9956,N_9281);
or U14914 (N_14914,N_10630,N_11961);
or U14915 (N_14915,N_9795,N_10534);
or U14916 (N_14916,N_10708,N_10040);
nor U14917 (N_14917,N_11336,N_11218);
nand U14918 (N_14918,N_9243,N_11136);
or U14919 (N_14919,N_9409,N_9624);
nand U14920 (N_14920,N_11212,N_10873);
or U14921 (N_14921,N_11527,N_10800);
and U14922 (N_14922,N_10366,N_10965);
nand U14923 (N_14923,N_11813,N_10587);
or U14924 (N_14924,N_10184,N_10524);
nand U14925 (N_14925,N_10732,N_11526);
or U14926 (N_14926,N_9495,N_10452);
nand U14927 (N_14927,N_9825,N_10029);
and U14928 (N_14928,N_11463,N_10257);
or U14929 (N_14929,N_9126,N_11399);
nand U14930 (N_14930,N_9493,N_11596);
or U14931 (N_14931,N_11844,N_9512);
and U14932 (N_14932,N_9757,N_10210);
or U14933 (N_14933,N_9391,N_10991);
nor U14934 (N_14934,N_10907,N_11579);
nor U14935 (N_14935,N_11428,N_9071);
nand U14936 (N_14936,N_11308,N_11520);
and U14937 (N_14937,N_10613,N_11372);
and U14938 (N_14938,N_9387,N_10646);
or U14939 (N_14939,N_9158,N_10626);
nor U14940 (N_14940,N_11179,N_9514);
xor U14941 (N_14941,N_11811,N_11386);
nor U14942 (N_14942,N_10290,N_10238);
nand U14943 (N_14943,N_10519,N_10621);
nand U14944 (N_14944,N_11063,N_9888);
nor U14945 (N_14945,N_9435,N_9955);
nor U14946 (N_14946,N_10544,N_10944);
nand U14947 (N_14947,N_10602,N_10998);
nor U14948 (N_14948,N_11238,N_9180);
and U14949 (N_14949,N_10699,N_10683);
and U14950 (N_14950,N_11341,N_10945);
and U14951 (N_14951,N_10115,N_9681);
xnor U14952 (N_14952,N_9588,N_11839);
nand U14953 (N_14953,N_10110,N_9410);
nand U14954 (N_14954,N_9440,N_10571);
and U14955 (N_14955,N_10045,N_11447);
and U14956 (N_14956,N_9978,N_11485);
or U14957 (N_14957,N_11342,N_10052);
nand U14958 (N_14958,N_11267,N_11837);
nor U14959 (N_14959,N_11096,N_11853);
nor U14960 (N_14960,N_9851,N_9318);
nor U14961 (N_14961,N_11178,N_11363);
nor U14962 (N_14962,N_10146,N_11670);
nor U14963 (N_14963,N_10975,N_10149);
and U14964 (N_14964,N_9904,N_9046);
and U14965 (N_14965,N_11530,N_11798);
and U14966 (N_14966,N_10468,N_9588);
or U14967 (N_14967,N_10158,N_9316);
nand U14968 (N_14968,N_10321,N_9846);
and U14969 (N_14969,N_10837,N_11332);
and U14970 (N_14970,N_11492,N_11738);
or U14971 (N_14971,N_10012,N_10498);
nand U14972 (N_14972,N_10539,N_9519);
and U14973 (N_14973,N_11849,N_10749);
or U14974 (N_14974,N_9864,N_11477);
and U14975 (N_14975,N_10379,N_11494);
and U14976 (N_14976,N_11696,N_11843);
nand U14977 (N_14977,N_9619,N_10521);
nor U14978 (N_14978,N_9579,N_9167);
nor U14979 (N_14979,N_11803,N_11787);
or U14980 (N_14980,N_11426,N_9647);
and U14981 (N_14981,N_10717,N_11057);
and U14982 (N_14982,N_9090,N_9656);
nand U14983 (N_14983,N_9420,N_9403);
or U14984 (N_14984,N_11499,N_10034);
and U14985 (N_14985,N_9008,N_9394);
and U14986 (N_14986,N_9039,N_10738);
or U14987 (N_14987,N_11227,N_9407);
nor U14988 (N_14988,N_10439,N_10351);
and U14989 (N_14989,N_10155,N_10099);
and U14990 (N_14990,N_10572,N_9185);
nor U14991 (N_14991,N_10775,N_9080);
nor U14992 (N_14992,N_10352,N_9683);
or U14993 (N_14993,N_9865,N_9921);
xor U14994 (N_14994,N_9098,N_10772);
nor U14995 (N_14995,N_11809,N_11812);
and U14996 (N_14996,N_10541,N_9082);
nor U14997 (N_14997,N_10532,N_11231);
nor U14998 (N_14998,N_9466,N_11108);
nor U14999 (N_14999,N_11405,N_9115);
nand UO_0 (O_0,N_13039,N_14899);
and UO_1 (O_1,N_14383,N_12663);
or UO_2 (O_2,N_12773,N_13774);
nand UO_3 (O_3,N_12085,N_12385);
nand UO_4 (O_4,N_12243,N_12553);
nor UO_5 (O_5,N_13825,N_14653);
nand UO_6 (O_6,N_12734,N_14168);
and UO_7 (O_7,N_14799,N_12602);
and UO_8 (O_8,N_13016,N_13734);
or UO_9 (O_9,N_14576,N_14635);
or UO_10 (O_10,N_12544,N_12560);
nor UO_11 (O_11,N_13741,N_12273);
and UO_12 (O_12,N_13682,N_13376);
nor UO_13 (O_13,N_12499,N_14546);
nand UO_14 (O_14,N_14138,N_14311);
and UO_15 (O_15,N_12726,N_14361);
nor UO_16 (O_16,N_12383,N_13539);
nand UO_17 (O_17,N_13501,N_12762);
nand UO_18 (O_18,N_12526,N_14292);
or UO_19 (O_19,N_14795,N_14433);
and UO_20 (O_20,N_13425,N_14780);
or UO_21 (O_21,N_14785,N_13094);
nand UO_22 (O_22,N_14389,N_14086);
and UO_23 (O_23,N_13577,N_13752);
and UO_24 (O_24,N_13731,N_14186);
or UO_25 (O_25,N_12057,N_12906);
or UO_26 (O_26,N_14758,N_13700);
and UO_27 (O_27,N_14166,N_12873);
nor UO_28 (O_28,N_12805,N_13944);
or UO_29 (O_29,N_13581,N_14956);
or UO_30 (O_30,N_14732,N_13138);
nand UO_31 (O_31,N_14497,N_12005);
nor UO_32 (O_32,N_14434,N_12113);
nor UO_33 (O_33,N_12994,N_13664);
nor UO_34 (O_34,N_14084,N_12502);
or UO_35 (O_35,N_12914,N_13690);
and UO_36 (O_36,N_13086,N_14170);
nand UO_37 (O_37,N_12742,N_14530);
or UO_38 (O_38,N_12096,N_12911);
and UO_39 (O_39,N_12839,N_14938);
nand UO_40 (O_40,N_14187,N_14588);
or UO_41 (O_41,N_12686,N_14744);
and UO_42 (O_42,N_14599,N_14879);
and UO_43 (O_43,N_12451,N_14997);
nand UO_44 (O_44,N_14723,N_13781);
and UO_45 (O_45,N_14487,N_14027);
or UO_46 (O_46,N_14387,N_13544);
and UO_47 (O_47,N_14976,N_14334);
nand UO_48 (O_48,N_12006,N_13365);
nand UO_49 (O_49,N_12014,N_14812);
nand UO_50 (O_50,N_13630,N_12258);
nor UO_51 (O_51,N_14451,N_12951);
and UO_52 (O_52,N_14330,N_14686);
and UO_53 (O_53,N_14637,N_12139);
nor UO_54 (O_54,N_14132,N_14660);
nand UO_55 (O_55,N_14774,N_13896);
nor UO_56 (O_56,N_14565,N_14306);
nand UO_57 (O_57,N_14531,N_14738);
nor UO_58 (O_58,N_13089,N_13048);
nand UO_59 (O_59,N_14188,N_14100);
nand UO_60 (O_60,N_12459,N_14566);
or UO_61 (O_61,N_12819,N_14199);
nor UO_62 (O_62,N_14855,N_12938);
nand UO_63 (O_63,N_12484,N_13477);
nor UO_64 (O_64,N_13267,N_13108);
or UO_65 (O_65,N_13214,N_12832);
or UO_66 (O_66,N_14690,N_13785);
xnor UO_67 (O_67,N_14789,N_12775);
or UO_68 (O_68,N_13804,N_12838);
and UO_69 (O_69,N_12927,N_13322);
nand UO_70 (O_70,N_12293,N_13132);
or UO_71 (O_71,N_12292,N_14849);
or UO_72 (O_72,N_12272,N_12260);
nand UO_73 (O_73,N_13388,N_14563);
nand UO_74 (O_74,N_12487,N_13657);
and UO_75 (O_75,N_13836,N_13768);
and UO_76 (O_76,N_12188,N_12635);
nor UO_77 (O_77,N_12376,N_12818);
nand UO_78 (O_78,N_13950,N_13171);
or UO_79 (O_79,N_12572,N_13380);
nand UO_80 (O_80,N_13585,N_12262);
or UO_81 (O_81,N_14721,N_12545);
or UO_82 (O_82,N_12104,N_14307);
xnor UO_83 (O_83,N_14549,N_13508);
or UO_84 (O_84,N_14864,N_12285);
and UO_85 (O_85,N_13715,N_12929);
or UO_86 (O_86,N_12406,N_14274);
nor UO_87 (O_87,N_13337,N_14413);
nor UO_88 (O_88,N_13260,N_14952);
or UO_89 (O_89,N_12398,N_12250);
nand UO_90 (O_90,N_14631,N_12696);
and UO_91 (O_91,N_12346,N_12470);
and UO_92 (O_92,N_13351,N_13824);
nand UO_93 (O_93,N_14619,N_14324);
or UO_94 (O_94,N_13517,N_12909);
nor UO_95 (O_95,N_13255,N_13426);
nor UO_96 (O_96,N_13166,N_12195);
or UO_97 (O_97,N_12965,N_14740);
nor UO_98 (O_98,N_13056,N_14582);
and UO_99 (O_99,N_12147,N_12310);
and UO_100 (O_100,N_14459,N_14702);
nand UO_101 (O_101,N_13583,N_13869);
nand UO_102 (O_102,N_12920,N_13343);
nor UO_103 (O_103,N_13188,N_12971);
nor UO_104 (O_104,N_13724,N_14435);
or UO_105 (O_105,N_13937,N_13582);
and UO_106 (O_106,N_12714,N_13943);
or UO_107 (O_107,N_12193,N_12855);
nand UO_108 (O_108,N_14421,N_12543);
or UO_109 (O_109,N_14480,N_14505);
and UO_110 (O_110,N_13125,N_13933);
or UO_111 (O_111,N_13156,N_14816);
xnor UO_112 (O_112,N_12858,N_13586);
and UO_113 (O_113,N_13604,N_14634);
and UO_114 (O_114,N_12180,N_13503);
nand UO_115 (O_115,N_12444,N_12606);
or UO_116 (O_116,N_14075,N_14983);
or UO_117 (O_117,N_12809,N_12004);
nor UO_118 (O_118,N_14820,N_14913);
nor UO_119 (O_119,N_13140,N_14044);
nand UO_120 (O_120,N_14578,N_13936);
and UO_121 (O_121,N_14171,N_12440);
nor UO_122 (O_122,N_13284,N_14162);
nand UO_123 (O_123,N_13952,N_13970);
and UO_124 (O_124,N_12549,N_14126);
nor UO_125 (O_125,N_14408,N_14496);
nor UO_126 (O_126,N_12901,N_13311);
nand UO_127 (O_127,N_14607,N_14600);
and UO_128 (O_128,N_13961,N_13318);
nor UO_129 (O_129,N_13221,N_12083);
and UO_130 (O_130,N_12569,N_14798);
and UO_131 (O_131,N_12844,N_12322);
nor UO_132 (O_132,N_14458,N_13231);
or UO_133 (O_133,N_13120,N_13018);
and UO_134 (O_134,N_13282,N_12640);
nor UO_135 (O_135,N_14895,N_14537);
nor UO_136 (O_136,N_13256,N_13122);
or UO_137 (O_137,N_13017,N_12015);
xor UO_138 (O_138,N_12656,N_12883);
and UO_139 (O_139,N_12660,N_12941);
and UO_140 (O_140,N_13098,N_12593);
nor UO_141 (O_141,N_12515,N_13840);
nand UO_142 (O_142,N_13168,N_12067);
nand UO_143 (O_143,N_13817,N_13654);
nand UO_144 (O_144,N_13207,N_13356);
or UO_145 (O_145,N_14392,N_12054);
and UO_146 (O_146,N_13325,N_14127);
nor UO_147 (O_147,N_13321,N_14289);
or UO_148 (O_148,N_14805,N_14338);
nor UO_149 (O_149,N_12366,N_13521);
nand UO_150 (O_150,N_13746,N_13025);
nor UO_151 (O_151,N_13885,N_14329);
or UO_152 (O_152,N_14046,N_13903);
nand UO_153 (O_153,N_14065,N_14058);
or UO_154 (O_154,N_14131,N_13536);
and UO_155 (O_155,N_12367,N_12771);
and UO_156 (O_156,N_12063,N_13195);
or UO_157 (O_157,N_12280,N_14181);
or UO_158 (O_158,N_12763,N_12348);
nand UO_159 (O_159,N_13241,N_14315);
nand UO_160 (O_160,N_12282,N_14129);
nor UO_161 (O_161,N_12021,N_13244);
nand UO_162 (O_162,N_13106,N_14230);
or UO_163 (O_163,N_14196,N_13819);
nand UO_164 (O_164,N_13934,N_14484);
and UO_165 (O_165,N_14834,N_13623);
nor UO_166 (O_166,N_13798,N_14647);
nor UO_167 (O_167,N_12103,N_14352);
and UO_168 (O_168,N_13530,N_14542);
nor UO_169 (O_169,N_13219,N_12616);
or UO_170 (O_170,N_13008,N_13850);
and UO_171 (O_171,N_13526,N_12425);
or UO_172 (O_172,N_13767,N_12071);
nor UO_173 (O_173,N_13485,N_13002);
and UO_174 (O_174,N_12482,N_14845);
and UO_175 (O_175,N_12979,N_12202);
nor UO_176 (O_176,N_14861,N_14406);
or UO_177 (O_177,N_14095,N_12680);
nand UO_178 (O_178,N_13917,N_14840);
nor UO_179 (O_179,N_14909,N_12027);
nor UO_180 (O_180,N_13161,N_13225);
xnor UO_181 (O_181,N_12806,N_12955);
nor UO_182 (O_182,N_13352,N_14357);
nand UO_183 (O_183,N_13829,N_12613);
or UO_184 (O_184,N_12298,N_12749);
and UO_185 (O_185,N_14907,N_12521);
or UO_186 (O_186,N_13736,N_14050);
or UO_187 (O_187,N_14355,N_14667);
nand UO_188 (O_188,N_12768,N_12893);
and UO_189 (O_189,N_12304,N_13513);
or UO_190 (O_190,N_13876,N_14376);
nand UO_191 (O_191,N_12752,N_12853);
nand UO_192 (O_192,N_13883,N_12415);
nor UO_193 (O_193,N_14949,N_13803);
nor UO_194 (O_194,N_12825,N_13424);
nand UO_195 (O_195,N_12991,N_14625);
and UO_196 (O_196,N_14892,N_14471);
nand UO_197 (O_197,N_13441,N_14632);
nor UO_198 (O_198,N_14950,N_12795);
nand UO_199 (O_199,N_14349,N_14499);
nand UO_200 (O_200,N_13651,N_13858);
nand UO_201 (O_201,N_14978,N_13766);
and UO_202 (O_202,N_12240,N_14322);
and UO_203 (O_203,N_12181,N_13958);
or UO_204 (O_204,N_12099,N_12120);
nor UO_205 (O_205,N_14124,N_13440);
and UO_206 (O_206,N_14219,N_13043);
nor UO_207 (O_207,N_14428,N_13831);
nor UO_208 (O_208,N_12141,N_12224);
nand UO_209 (O_209,N_14431,N_14846);
or UO_210 (O_210,N_13925,N_12158);
or UO_211 (O_211,N_14716,N_12769);
nand UO_212 (O_212,N_13872,N_14457);
or UO_213 (O_213,N_13710,N_12932);
and UO_214 (O_214,N_13624,N_13049);
and UO_215 (O_215,N_12408,N_12291);
nand UO_216 (O_216,N_12600,N_13929);
nand UO_217 (O_217,N_13681,N_13986);
or UO_218 (O_218,N_12748,N_14368);
or UO_219 (O_219,N_14140,N_14426);
and UO_220 (O_220,N_14222,N_14227);
or UO_221 (O_221,N_14103,N_14544);
nand UO_222 (O_222,N_14034,N_13190);
or UO_223 (O_223,N_12238,N_13044);
nand UO_224 (O_224,N_14904,N_12361);
nor UO_225 (O_225,N_13749,N_12305);
and UO_226 (O_226,N_13495,N_12102);
nand UO_227 (O_227,N_12698,N_13704);
or UO_228 (O_228,N_13652,N_14807);
and UO_229 (O_229,N_14013,N_13626);
nand UO_230 (O_230,N_12179,N_14609);
nand UO_231 (O_231,N_13598,N_13780);
and UO_232 (O_232,N_13887,N_12118);
nor UO_233 (O_233,N_13727,N_12319);
and UO_234 (O_234,N_14614,N_14948);
nor UO_235 (O_235,N_13891,N_14291);
and UO_236 (O_236,N_12232,N_14994);
and UO_237 (O_237,N_12245,N_14351);
nand UO_238 (O_238,N_14098,N_13870);
nor UO_239 (O_239,N_12985,N_12491);
nor UO_240 (O_240,N_14060,N_13402);
nor UO_241 (O_241,N_13571,N_12090);
nand UO_242 (O_242,N_12791,N_12064);
nor UO_243 (O_243,N_13471,N_12710);
and UO_244 (O_244,N_13665,N_14183);
nor UO_245 (O_245,N_12641,N_14698);
nor UO_246 (O_246,N_14813,N_13689);
nor UO_247 (O_247,N_13150,N_12435);
and UO_248 (O_248,N_14118,N_13488);
nor UO_249 (O_249,N_12998,N_12581);
nor UO_250 (O_250,N_14601,N_14377);
nand UO_251 (O_251,N_14247,N_12928);
nand UO_252 (O_252,N_13875,N_12325);
or UO_253 (O_253,N_13867,N_14198);
and UO_254 (O_254,N_13229,N_14955);
nand UO_255 (O_255,N_12599,N_12974);
or UO_256 (O_256,N_14704,N_12295);
nand UO_257 (O_257,N_13423,N_12207);
nor UO_258 (O_258,N_12508,N_14932);
and UO_259 (O_259,N_13786,N_13320);
and UO_260 (O_260,N_14397,N_14741);
and UO_261 (O_261,N_13186,N_13733);
nor UO_262 (O_262,N_12454,N_12667);
or UO_263 (O_263,N_12815,N_13923);
and UO_264 (O_264,N_12342,N_14485);
nand UO_265 (O_265,N_12664,N_12199);
nor UO_266 (O_266,N_13595,N_12221);
or UO_267 (O_267,N_13643,N_13900);
nor UO_268 (O_268,N_14763,N_13182);
and UO_269 (O_269,N_12317,N_12442);
nand UO_270 (O_270,N_13069,N_14827);
and UO_271 (O_271,N_12392,N_12166);
or UO_272 (O_272,N_14231,N_13930);
nand UO_273 (O_273,N_12650,N_12165);
or UO_274 (O_274,N_13893,N_13844);
nor UO_275 (O_275,N_14179,N_12558);
or UO_276 (O_276,N_12235,N_14016);
nor UO_277 (O_277,N_13742,N_14176);
nand UO_278 (O_278,N_13249,N_12903);
and UO_279 (O_279,N_13789,N_12935);
nand UO_280 (O_280,N_14562,N_14500);
nand UO_281 (O_281,N_12958,N_13871);
nor UO_282 (O_282,N_14865,N_13748);
and UO_283 (O_283,N_13985,N_12862);
or UO_284 (O_284,N_13790,N_13111);
nand UO_285 (O_285,N_13174,N_14266);
and UO_286 (O_286,N_14854,N_14374);
nand UO_287 (O_287,N_14178,N_13014);
or UO_288 (O_288,N_13594,N_14271);
nand UO_289 (O_289,N_12737,N_13747);
nor UO_290 (O_290,N_13841,N_12702);
or UO_291 (O_291,N_12441,N_13183);
and UO_292 (O_292,N_14282,N_13864);
nor UO_293 (O_293,N_12643,N_13969);
and UO_294 (O_294,N_13979,N_14725);
nor UO_295 (O_295,N_14919,N_12793);
or UO_296 (O_296,N_12175,N_14669);
nor UO_297 (O_297,N_12024,N_14220);
and UO_298 (O_298,N_12916,N_13147);
nand UO_299 (O_299,N_12945,N_14398);
or UO_300 (O_300,N_13187,N_13511);
or UO_301 (O_301,N_12419,N_13035);
nand UO_302 (O_302,N_12725,N_12143);
nor UO_303 (O_303,N_12570,N_13019);
or UO_304 (O_304,N_12041,N_13631);
and UO_305 (O_305,N_13305,N_12625);
nor UO_306 (O_306,N_13890,N_12492);
nor UO_307 (O_307,N_13579,N_12003);
xor UO_308 (O_308,N_13336,N_12318);
and UO_309 (O_309,N_13576,N_14708);
nor UO_310 (O_310,N_14111,N_13496);
nor UO_311 (O_311,N_13981,N_12939);
nor UO_312 (O_312,N_12984,N_14203);
and UO_313 (O_313,N_14482,N_13597);
and UO_314 (O_314,N_14825,N_13644);
or UO_315 (O_315,N_12327,N_13713);
nor UO_316 (O_316,N_13063,N_13638);
and UO_317 (O_317,N_14216,N_14536);
nand UO_318 (O_318,N_12896,N_12607);
nor UO_319 (O_319,N_12471,N_14474);
nor UO_320 (O_320,N_14073,N_14999);
and UO_321 (O_321,N_13419,N_14346);
or UO_322 (O_322,N_13239,N_12833);
or UO_323 (O_323,N_14185,N_12138);
nor UO_324 (O_324,N_14101,N_14359);
or UO_325 (O_325,N_14273,N_14224);
and UO_326 (O_326,N_14063,N_12403);
nand UO_327 (O_327,N_14262,N_12445);
and UO_328 (O_328,N_12628,N_12448);
or UO_329 (O_329,N_13418,N_14108);
or UO_330 (O_330,N_12764,N_14942);
nand UO_331 (O_331,N_14621,N_12247);
and UO_332 (O_332,N_14069,N_14573);
or UO_333 (O_333,N_12452,N_14200);
nor UO_334 (O_334,N_12146,N_14739);
nor UO_335 (O_335,N_12174,N_12925);
or UO_336 (O_336,N_13332,N_14509);
or UO_337 (O_337,N_12168,N_12511);
nor UO_338 (O_338,N_12644,N_12533);
nor UO_339 (O_339,N_13180,N_14654);
nand UO_340 (O_340,N_13611,N_12183);
nor UO_341 (O_341,N_13148,N_12388);
nor UO_342 (O_342,N_14819,N_12156);
nand UO_343 (O_343,N_12275,N_12759);
or UO_344 (O_344,N_12144,N_14571);
xor UO_345 (O_345,N_12414,N_13059);
nand UO_346 (O_346,N_14844,N_13153);
and UO_347 (O_347,N_14501,N_13309);
nand UO_348 (O_348,N_12861,N_12042);
nand UO_349 (O_349,N_14303,N_12200);
nand UO_350 (O_350,N_13264,N_12326);
nor UO_351 (O_351,N_13915,N_13678);
nor UO_352 (O_352,N_13022,N_13191);
or UO_353 (O_353,N_12384,N_12897);
or UO_354 (O_354,N_14888,N_13660);
nor UO_355 (O_355,N_13026,N_14305);
or UO_356 (O_356,N_12196,N_12501);
nor UO_357 (O_357,N_14745,N_13942);
nor UO_358 (O_358,N_13967,N_13912);
and UO_359 (O_359,N_13340,N_13708);
or UO_360 (O_360,N_12251,N_12595);
and UO_361 (O_361,N_14350,N_13298);
nor UO_362 (O_362,N_12946,N_12962);
nor UO_363 (O_363,N_14028,N_12031);
or UO_364 (O_364,N_13009,N_14335);
and UO_365 (O_365,N_14513,N_13116);
and UO_366 (O_366,N_13762,N_12178);
nand UO_367 (O_367,N_14048,N_12720);
and UO_368 (O_368,N_12401,N_12343);
or UO_369 (O_369,N_14523,N_14277);
nand UO_370 (O_370,N_12337,N_13091);
nand UO_371 (O_371,N_14823,N_14014);
or UO_372 (O_372,N_13199,N_14256);
and UO_373 (O_373,N_12541,N_12489);
nor UO_374 (O_374,N_14233,N_12056);
and UO_375 (O_375,N_14596,N_13811);
nor UO_376 (O_376,N_14891,N_14011);
nor UO_377 (O_377,N_14232,N_12687);
and UO_378 (O_378,N_12476,N_14842);
nand UO_379 (O_379,N_12461,N_14608);
or UO_380 (O_380,N_12070,N_12007);
and UO_381 (O_381,N_13721,N_14666);
nand UO_382 (O_382,N_12802,N_13692);
and UO_383 (O_383,N_13232,N_13353);
or UO_384 (O_384,N_12624,N_13647);
nand UO_385 (O_385,N_14701,N_13550);
nand UO_386 (O_386,N_12923,N_12697);
nor UO_387 (O_387,N_14156,N_12344);
and UO_388 (O_388,N_14279,N_13629);
nor UO_389 (O_389,N_12821,N_13552);
or UO_390 (O_390,N_13765,N_12430);
or UO_391 (O_391,N_13141,N_14285);
nand UO_392 (O_392,N_12807,N_12836);
and UO_393 (O_393,N_12049,N_12101);
nor UO_394 (O_394,N_12980,N_12259);
or UO_395 (O_395,N_14677,N_14452);
nand UO_396 (O_396,N_14979,N_12707);
nor UO_397 (O_397,N_13245,N_14929);
nor UO_398 (O_398,N_13650,N_14894);
nor UO_399 (O_399,N_12271,N_13294);
nand UO_400 (O_400,N_12605,N_13348);
or UO_401 (O_401,N_13907,N_13978);
and UO_402 (O_402,N_13744,N_12222);
nand UO_403 (O_403,N_12803,N_13416);
nand UO_404 (O_404,N_13888,N_14354);
nand UO_405 (O_405,N_13874,N_13154);
nand UO_406 (O_406,N_13655,N_12885);
and UO_407 (O_407,N_13432,N_13822);
nor UO_408 (O_408,N_14991,N_14042);
nand UO_409 (O_409,N_14281,N_14877);
or UO_410 (O_410,N_12869,N_13984);
nor UO_411 (O_411,N_13545,N_12842);
and UO_412 (O_412,N_13490,N_12400);
and UO_413 (O_413,N_13843,N_14438);
nand UO_414 (O_414,N_13658,N_12485);
or UO_415 (O_415,N_14278,N_12283);
or UO_416 (O_416,N_12418,N_14441);
nor UO_417 (O_417,N_14193,N_14752);
nor UO_418 (O_418,N_12865,N_12647);
or UO_419 (O_419,N_13673,N_13818);
or UO_420 (O_420,N_14080,N_12431);
or UO_421 (O_421,N_12094,N_13115);
or UO_422 (O_422,N_14293,N_13683);
or UO_423 (O_423,N_13442,N_14314);
nand UO_424 (O_424,N_12886,N_14436);
nand UO_425 (O_425,N_14460,N_13670);
or UO_426 (O_426,N_13770,N_12525);
and UO_427 (O_427,N_12693,N_14524);
and UO_428 (O_428,N_12703,N_13235);
or UO_429 (O_429,N_13460,N_12249);
nand UO_430 (O_430,N_12131,N_13411);
or UO_431 (O_431,N_13935,N_12876);
or UO_432 (O_432,N_12948,N_12827);
nand UO_433 (O_433,N_14520,N_13753);
or UO_434 (O_434,N_12469,N_14286);
nand UO_435 (O_435,N_12128,N_13566);
or UO_436 (O_436,N_14810,N_14419);
nand UO_437 (O_437,N_13385,N_14870);
nand UO_438 (O_438,N_12604,N_13620);
and UO_439 (O_439,N_13760,N_13007);
and UO_440 (O_440,N_14665,N_14859);
or UO_441 (O_441,N_13688,N_13773);
and UO_442 (O_442,N_13719,N_14308);
nor UO_443 (O_443,N_13557,N_12753);
nor UO_444 (O_444,N_14477,N_14339);
or UO_445 (O_445,N_14372,N_14673);
nand UO_446 (O_446,N_12025,N_12859);
nor UO_447 (O_447,N_12652,N_13527);
or UO_448 (O_448,N_13792,N_14139);
nand UO_449 (O_449,N_12566,N_13030);
nor UO_450 (O_450,N_14478,N_13213);
and UO_451 (O_451,N_14730,N_13354);
nand UO_452 (O_452,N_13522,N_12117);
or UO_453 (O_453,N_13757,N_13962);
nor UO_454 (O_454,N_13013,N_14679);
and UO_455 (O_455,N_12591,N_12637);
nand UO_456 (O_456,N_12576,N_12691);
or UO_457 (O_457,N_14990,N_14089);
xor UO_458 (O_458,N_14194,N_14159);
nand UO_459 (O_459,N_12642,N_14618);
nor UO_460 (O_460,N_14803,N_12648);
or UO_461 (O_461,N_13344,N_13834);
nor UO_462 (O_462,N_14328,N_12472);
nor UO_463 (O_463,N_12162,N_14402);
or UO_464 (O_464,N_13389,N_13662);
or UO_465 (O_465,N_14963,N_12864);
nor UO_466 (O_466,N_12206,N_13333);
or UO_467 (O_467,N_12402,N_14033);
nor UO_468 (O_468,N_12187,N_14589);
nand UO_469 (O_469,N_12574,N_13203);
nor UO_470 (O_470,N_12931,N_14117);
nor UO_471 (O_471,N_14411,N_14295);
nor UO_472 (O_472,N_14786,N_12785);
xor UO_473 (O_473,N_14229,N_14056);
and UO_474 (O_474,N_13973,N_13377);
and UO_475 (O_475,N_12449,N_12133);
or UO_476 (O_476,N_12550,N_13467);
nor UO_477 (O_477,N_13291,N_12443);
nand UO_478 (O_478,N_14733,N_12790);
or UO_479 (O_479,N_14779,N_13073);
nor UO_480 (O_480,N_14041,N_13737);
nor UO_481 (O_481,N_13756,N_12378);
nor UO_482 (O_482,N_14047,N_14751);
and UO_483 (O_483,N_12226,N_12329);
nand UO_484 (O_484,N_12436,N_14863);
or UO_485 (O_485,N_13479,N_14757);
nor UO_486 (O_486,N_12288,N_12227);
or UO_487 (O_487,N_13437,N_14724);
nand UO_488 (O_488,N_12333,N_12405);
or UO_489 (O_489,N_13999,N_12672);
nor UO_490 (O_490,N_14450,N_13649);
or UO_491 (O_491,N_14756,N_12908);
or UO_492 (O_492,N_13134,N_14353);
nor UO_493 (O_493,N_14380,N_12137);
nor UO_494 (O_494,N_12368,N_12562);
or UO_495 (O_495,N_13555,N_12142);
nand UO_496 (O_496,N_12524,N_12789);
or UO_497 (O_497,N_14128,N_14195);
or UO_498 (O_498,N_14212,N_12173);
nand UO_499 (O_499,N_13295,N_12347);
or UO_500 (O_500,N_13103,N_14465);
and UO_501 (O_501,N_13093,N_12301);
nand UO_502 (O_502,N_12062,N_12437);
nand UO_503 (O_503,N_13457,N_14663);
or UO_504 (O_504,N_12052,N_12638);
or UO_505 (O_505,N_13474,N_14826);
or UO_506 (O_506,N_13945,N_13990);
and UO_507 (O_507,N_12706,N_13832);
nor UO_508 (O_508,N_14604,N_14746);
and UO_509 (O_509,N_14694,N_13669);
nor UO_510 (O_510,N_14720,N_13310);
and UO_511 (O_511,N_13248,N_13211);
and UO_512 (O_512,N_12309,N_14209);
or UO_513 (O_513,N_14936,N_13184);
and UO_514 (O_514,N_12364,N_12567);
nand UO_515 (O_515,N_14284,N_12194);
nor UO_516 (O_516,N_13464,N_12395);
and UO_517 (O_517,N_12701,N_13684);
nand UO_518 (O_518,N_12084,N_12252);
nor UO_519 (O_519,N_12912,N_14481);
nor UO_520 (O_520,N_14313,N_13395);
or UO_521 (O_521,N_12051,N_14903);
and UO_522 (O_522,N_13468,N_14550);
nor UO_523 (O_523,N_13393,N_13596);
nand UO_524 (O_524,N_13033,N_14053);
or UO_525 (O_525,N_12959,N_13699);
nor UO_526 (O_526,N_14633,N_14945);
nor UO_527 (O_527,N_12675,N_14268);
and UO_528 (O_528,N_12716,N_13081);
nand UO_529 (O_529,N_13677,N_14561);
nand UO_530 (O_530,N_12766,N_13208);
nor UO_531 (O_531,N_12510,N_13516);
and UO_532 (O_532,N_14759,N_14259);
nand UO_533 (O_533,N_12503,N_13809);
and UO_534 (O_534,N_14885,N_12040);
and UO_535 (O_535,N_13777,N_14533);
nand UO_536 (O_536,N_14331,N_12394);
nor UO_537 (O_537,N_14897,N_12032);
nor UO_538 (O_538,N_12812,N_13612);
nand UO_539 (O_539,N_13640,N_13105);
nand UO_540 (O_540,N_13163,N_12776);
nor UO_541 (O_541,N_13642,N_14163);
and UO_542 (O_542,N_14985,N_13286);
nor UO_543 (O_543,N_14773,N_12059);
nand UO_544 (O_544,N_14081,N_14753);
nand UO_545 (O_545,N_12692,N_12996);
and UO_546 (O_546,N_12881,N_12080);
nand UO_547 (O_547,N_14624,N_12268);
nor UO_548 (O_548,N_13121,N_12741);
nand UO_549 (O_549,N_12241,N_12314);
or UO_550 (O_550,N_14023,N_13603);
or UO_551 (O_551,N_12846,N_13641);
nor UO_552 (O_552,N_14747,N_14680);
and UO_553 (O_553,N_12111,N_12170);
or UO_554 (O_554,N_14772,N_14119);
or UO_555 (O_555,N_12784,N_13075);
and UO_556 (O_556,N_14876,N_14922);
or UO_557 (O_557,N_13838,N_12256);
nand UO_558 (O_558,N_13347,N_14797);
nor UO_559 (O_559,N_14177,N_13205);
or UO_560 (O_560,N_13608,N_12622);
nand UO_561 (O_561,N_14943,N_14364);
and UO_562 (O_562,N_14783,N_12705);
nor UO_563 (O_563,N_14043,N_14926);
and UO_564 (O_564,N_13548,N_13856);
and UO_565 (O_565,N_13610,N_12538);
and UO_566 (O_566,N_14371,N_13862);
nor UO_567 (O_567,N_13820,N_13178);
nor UO_568 (O_568,N_14228,N_13728);
or UO_569 (O_569,N_12300,N_12770);
nand UO_570 (O_570,N_12801,N_13443);
nand UO_571 (O_571,N_14257,N_13633);
and UO_572 (O_572,N_13123,N_14587);
nand UO_573 (O_573,N_12708,N_14822);
or UO_574 (O_574,N_13735,N_14538);
nor UO_575 (O_575,N_12646,N_12761);
nand UO_576 (O_576,N_12756,N_13455);
nand UO_577 (O_577,N_13551,N_13288);
or UO_578 (O_578,N_12596,N_13927);
and UO_579 (O_579,N_12584,N_13158);
or UO_580 (O_580,N_14557,N_14092);
or UO_581 (O_581,N_12270,N_13117);
or UO_582 (O_582,N_12717,N_12255);
or UO_583 (O_583,N_12214,N_12087);
nand UO_584 (O_584,N_13564,N_14367);
and UO_585 (O_585,N_14323,N_12100);
nor UO_586 (O_586,N_13941,N_14464);
nand UO_587 (O_587,N_12788,N_13435);
nor UO_588 (O_588,N_13082,N_12840);
or UO_589 (O_589,N_12189,N_14172);
and UO_590 (O_590,N_13863,N_14400);
nand UO_591 (O_591,N_14540,N_13529);
nand UO_592 (O_592,N_13114,N_12197);
nand UO_593 (O_593,N_13242,N_14373);
or UO_594 (O_594,N_12185,N_14466);
and UO_595 (O_595,N_14336,N_13361);
and UO_596 (O_596,N_14057,N_14115);
and UO_597 (O_597,N_13370,N_12877);
nor UO_598 (O_598,N_13589,N_14296);
and UO_599 (O_599,N_14064,N_14644);
or UO_600 (O_600,N_14341,N_13053);
nand UO_601 (O_601,N_12234,N_12774);
nor UO_602 (O_602,N_12612,N_12152);
and UO_603 (O_603,N_12653,N_13279);
nor UO_604 (O_604,N_13278,N_12580);
and UO_605 (O_605,N_14096,N_13601);
nand UO_606 (O_606,N_14717,N_13360);
nand UO_607 (O_607,N_14569,N_14409);
nor UO_608 (O_608,N_12108,N_13717);
or UO_609 (O_609,N_13124,N_14927);
or UO_610 (O_610,N_13963,N_13478);
nand UO_611 (O_611,N_12001,N_13261);
nand UO_612 (O_612,N_13901,N_14365);
and UO_613 (O_613,N_13918,N_12230);
or UO_614 (O_614,N_14283,N_13051);
and UO_615 (O_615,N_14715,N_14964);
and UO_616 (O_616,N_13625,N_14532);
nor UO_617 (O_617,N_14189,N_14051);
or UO_618 (O_618,N_13909,N_14815);
nand UO_619 (O_619,N_13782,N_13632);
and UO_620 (O_620,N_12715,N_13165);
and UO_621 (O_621,N_13702,N_13143);
or UO_622 (O_622,N_14937,N_14527);
or UO_623 (O_623,N_13454,N_14630);
or UO_624 (O_624,N_12016,N_13331);
nand UO_625 (O_625,N_14275,N_12396);
nand UO_626 (O_626,N_13216,N_14210);
nand UO_627 (O_627,N_13461,N_14239);
or UO_628 (O_628,N_13619,N_14560);
nor UO_629 (O_629,N_13271,N_14022);
nand UO_630 (O_630,N_12330,N_14959);
or UO_631 (O_631,N_13397,N_13796);
and UO_632 (O_632,N_12588,N_13367);
or UO_633 (O_633,N_12422,N_14029);
nand UO_634 (O_634,N_12498,N_12012);
or UO_635 (O_635,N_12603,N_12617);
nand UO_636 (O_636,N_12532,N_13797);
and UO_637 (O_637,N_13057,N_13519);
and UO_638 (O_638,N_14440,N_14568);
nor UO_639 (O_639,N_13068,N_14886);
nor UO_640 (O_640,N_12548,N_12302);
and UO_641 (O_641,N_12353,N_14574);
or UO_642 (O_642,N_12380,N_14290);
and UO_643 (O_643,N_12129,N_13592);
and UO_644 (O_644,N_14018,N_14731);
nor UO_645 (O_645,N_14264,N_14676);
and UO_646 (O_646,N_13515,N_13405);
or UO_647 (O_647,N_14122,N_12246);
and UO_648 (O_648,N_12306,N_14143);
or UO_649 (O_649,N_14150,N_13252);
or UO_650 (O_650,N_13563,N_13299);
nor UO_651 (O_651,N_14984,N_14152);
or UO_652 (O_652,N_14824,N_13494);
xor UO_653 (O_653,N_13701,N_12046);
nor UO_654 (O_654,N_14390,N_12516);
or UO_655 (O_655,N_13480,N_12944);
or UO_656 (O_656,N_13429,N_14605);
or UO_657 (O_657,N_13860,N_13543);
nor UO_658 (O_658,N_14862,N_14900);
and UO_659 (O_659,N_13032,N_13324);
and UO_660 (O_660,N_12694,N_13714);
nor UO_661 (O_661,N_13413,N_14005);
nand UO_662 (O_662,N_13730,N_12621);
xnor UO_663 (O_663,N_13940,N_14893);
nand UO_664 (O_664,N_12954,N_13745);
nor UO_665 (O_665,N_14363,N_13865);
or UO_666 (O_666,N_13989,N_13559);
nand UO_667 (O_667,N_13088,N_13868);
nor UO_668 (O_668,N_14602,N_14727);
and UO_669 (O_669,N_14083,N_12536);
nor UO_670 (O_670,N_12719,N_12136);
nand UO_671 (O_671,N_13991,N_13290);
nor UO_672 (O_672,N_12870,N_12736);
nor UO_673 (O_673,N_14489,N_12816);
nand UO_674 (O_674,N_13371,N_14302);
nor UO_675 (O_675,N_13645,N_14896);
nor UO_676 (O_676,N_14914,N_13304);
or UO_677 (O_677,N_13109,N_13220);
nand UO_678 (O_678,N_13812,N_13137);
nor UO_679 (O_679,N_13146,N_14719);
or UO_680 (O_680,N_14197,N_12279);
nor UO_681 (O_681,N_14002,N_12947);
or UO_682 (O_682,N_13622,N_13977);
and UO_683 (O_683,N_12649,N_14378);
or UO_684 (O_684,N_13217,N_14711);
or UO_685 (O_685,N_13070,N_12554);
or UO_686 (O_686,N_14917,N_14572);
nand UO_687 (O_687,N_13924,N_13897);
nand UO_688 (O_688,N_14417,N_13857);
nand UO_689 (O_689,N_13821,N_14078);
nand UO_690 (O_690,N_13483,N_14215);
nand UO_691 (O_691,N_14828,N_13466);
or UO_692 (O_692,N_13816,N_13335);
and UO_693 (O_693,N_13189,N_12020);
nor UO_694 (O_694,N_12239,N_13497);
or UO_695 (O_695,N_13584,N_12982);
and UO_696 (O_696,N_14468,N_14790);
nor UO_697 (O_697,N_12857,N_14503);
and UO_698 (O_698,N_14792,N_12655);
or UO_699 (O_699,N_13541,N_13698);
or UO_700 (O_700,N_14971,N_13027);
or UO_701 (O_701,N_13470,N_12835);
nand UO_702 (O_702,N_12438,N_13637);
or UO_703 (O_703,N_14424,N_12389);
and UO_704 (O_704,N_14652,N_14399);
nand UO_705 (O_705,N_13313,N_12072);
nor UO_706 (O_706,N_12311,N_12217);
nand UO_707 (O_707,N_14661,N_12287);
and UO_708 (O_708,N_14356,N_13772);
and UO_709 (O_709,N_14941,N_14547);
or UO_710 (O_710,N_14366,N_14299);
or UO_711 (O_711,N_12154,N_14309);
nor UO_712 (O_712,N_14184,N_12145);
nand UO_713 (O_713,N_12284,N_14890);
nand UO_714 (O_714,N_13492,N_12760);
nor UO_715 (O_715,N_12918,N_13590);
nor UO_716 (O_716,N_12514,N_14930);
nor UO_717 (O_717,N_12799,N_12804);
nor UO_718 (O_718,N_14407,N_13446);
and UO_719 (O_719,N_13755,N_13675);
nand UO_720 (O_720,N_13855,N_14954);
and UO_721 (O_721,N_13880,N_13301);
nor UO_722 (O_722,N_12848,N_14507);
or UO_723 (O_723,N_14981,N_14836);
nor UO_724 (O_724,N_13157,N_14067);
nor UO_725 (O_725,N_12190,N_12248);
and UO_726 (O_726,N_14650,N_13499);
nor UO_727 (O_727,N_14771,N_14035);
xor UO_728 (O_728,N_13036,N_13133);
nand UO_729 (O_729,N_12420,N_14074);
or UO_730 (O_730,N_12608,N_12357);
and UO_731 (O_731,N_14947,N_13374);
nor UO_732 (O_732,N_13671,N_12689);
or UO_733 (O_733,N_12778,N_13562);
nand UO_734 (O_734,N_13826,N_13258);
or UO_735 (O_735,N_13761,N_14734);
xnor UO_736 (O_736,N_13297,N_14645);
nor UO_737 (O_737,N_14902,N_12631);
nor UO_738 (O_738,N_14688,N_13080);
or UO_739 (O_739,N_13006,N_13653);
or UO_740 (O_740,N_14970,N_13170);
and UO_741 (O_741,N_12598,N_14493);
or UO_742 (O_742,N_12009,N_12978);
nand UO_743 (O_743,N_14025,N_12375);
and UO_744 (O_744,N_12618,N_12261);
or UO_745 (O_745,N_14444,N_14764);
or UO_746 (O_746,N_12462,N_13759);
or UO_747 (O_747,N_13277,N_12999);
and UO_748 (O_748,N_12172,N_12547);
and UO_749 (O_749,N_14627,N_13709);
or UO_750 (O_750,N_12729,N_14248);
nor UO_751 (O_751,N_13328,N_13046);
and UO_752 (O_752,N_12699,N_12155);
nor UO_753 (O_753,N_14343,N_14748);
nor UO_754 (O_754,N_12856,N_14052);
or UO_755 (O_755,N_14395,N_13421);
and UO_756 (O_756,N_12738,N_14455);
nor UO_757 (O_757,N_12630,N_14375);
nor UO_758 (O_758,N_12460,N_12614);
nand UO_759 (O_759,N_14583,N_13078);
nand UO_760 (O_760,N_14781,N_12851);
or UO_761 (O_761,N_14495,N_13458);
nor UO_762 (O_762,N_14591,N_12623);
nand UO_763 (O_763,N_14884,N_14422);
or UO_764 (O_764,N_14967,N_13666);
nor UO_765 (O_765,N_13453,N_12830);
nor UO_766 (O_766,N_12429,N_14486);
nand UO_767 (O_767,N_13040,N_14072);
nor UO_768 (O_768,N_14423,N_12213);
nor UO_769 (O_769,N_13906,N_12077);
and UO_770 (O_770,N_14996,N_12975);
nor UO_771 (O_771,N_13591,N_12455);
nand UO_772 (O_772,N_14213,N_12875);
and UO_773 (O_773,N_14358,N_13206);
nor UO_774 (O_774,N_14993,N_13061);
or UO_775 (O_775,N_14946,N_14674);
or UO_776 (O_776,N_14412,N_14534);
or UO_777 (O_777,N_13489,N_14622);
or UO_778 (O_778,N_14965,N_14137);
nor UO_779 (O_779,N_14575,N_13902);
and UO_780 (O_780,N_12477,N_12130);
nor UO_781 (O_781,N_13621,N_14850);
nor UO_782 (O_782,N_14208,N_14332);
or UO_783 (O_783,N_12223,N_13672);
nor UO_784 (O_784,N_14418,N_14180);
nand UO_785 (O_785,N_14610,N_14553);
and UO_786 (O_786,N_14347,N_14467);
or UO_787 (O_787,N_14326,N_14966);
nand UO_788 (O_788,N_12530,N_13661);
nor UO_789 (O_789,N_12186,N_12810);
and UO_790 (O_790,N_14640,N_12294);
and UO_791 (O_791,N_14001,N_13546);
nand UO_792 (O_792,N_13386,N_14592);
nor UO_793 (O_793,N_14449,N_14304);
xnor UO_794 (O_794,N_14791,N_12850);
or UO_795 (O_795,N_12331,N_13238);
nand UO_796 (O_796,N_12321,N_14294);
or UO_797 (O_797,N_13269,N_13427);
and UO_798 (O_798,N_13995,N_14515);
and UO_799 (O_799,N_12953,N_12892);
or UO_800 (O_800,N_14829,N_12668);
or UO_801 (O_801,N_13813,N_13247);
nor UO_802 (O_802,N_13417,N_14838);
nor UO_803 (O_803,N_14671,N_12157);
or UO_804 (O_804,N_12229,N_14852);
or UO_805 (O_805,N_13707,N_12907);
or UO_806 (O_806,N_14445,N_13407);
nand UO_807 (O_807,N_12627,N_13272);
and UO_808 (O_808,N_12828,N_13445);
or UO_809 (O_809,N_13218,N_13634);
or UO_810 (O_810,N_12546,N_12561);
and UO_811 (O_811,N_12468,N_13129);
and UO_812 (O_812,N_12552,N_12732);
nor UO_813 (O_813,N_12163,N_13280);
or UO_814 (O_814,N_14379,N_12814);
and UO_815 (O_815,N_12727,N_13932);
and UO_816 (O_816,N_13274,N_14910);
nor UO_817 (O_817,N_14858,N_13020);
nand UO_818 (O_818,N_12709,N_14476);
and UO_819 (O_819,N_13646,N_14327);
nand UO_820 (O_820,N_13635,N_13212);
nor UO_821 (O_821,N_12535,N_12556);
or UO_822 (O_822,N_14288,N_13788);
or UO_823 (O_823,N_14794,N_14975);
nand UO_824 (O_824,N_13830,N_14251);
nor UO_825 (O_825,N_14867,N_14488);
and UO_826 (O_826,N_12000,N_12363);
or UO_827 (O_827,N_14742,N_13778);
or UO_828 (O_828,N_13743,N_14683);
or UO_829 (O_829,N_14154,N_14019);
nor UO_830 (O_830,N_12589,N_12467);
and UO_831 (O_831,N_13276,N_12088);
and UO_832 (O_832,N_12116,N_13916);
nand UO_833 (O_833,N_13775,N_13845);
or UO_834 (O_834,N_14254,N_12743);
nor UO_835 (O_835,N_14218,N_12659);
or UO_836 (O_836,N_13848,N_12488);
nand UO_837 (O_837,N_13119,N_12028);
and UO_838 (O_838,N_12244,N_14026);
xnor UO_839 (O_839,N_13167,N_13066);
nor UO_840 (O_840,N_14603,N_14728);
and UO_841 (O_841,N_13096,N_12266);
nor UO_842 (O_842,N_12757,N_12841);
nand UO_843 (O_843,N_14918,N_12296);
and UO_844 (O_844,N_14818,N_13266);
nor UO_845 (O_845,N_12845,N_14657);
nor UO_846 (O_846,N_12434,N_13330);
or UO_847 (O_847,N_14519,N_14113);
nand UO_848 (O_848,N_13600,N_12496);
or UO_849 (O_849,N_13283,N_13507);
nand UO_850 (O_850,N_14225,N_14007);
nand UO_851 (O_851,N_12531,N_14944);
nor UO_852 (O_852,N_12798,N_13270);
or UO_853 (O_853,N_12993,N_14814);
or UO_854 (O_854,N_13381,N_12231);
nor UO_855 (O_855,N_12479,N_12215);
nor UO_856 (O_856,N_14204,N_12781);
nand UO_857 (O_857,N_14755,N_14526);
or UO_858 (O_858,N_14242,N_14032);
or UO_859 (O_859,N_14453,N_14830);
nor UO_860 (O_860,N_14808,N_13636);
nand UO_861 (O_861,N_13783,N_13691);
or UO_862 (O_862,N_14040,N_13064);
nor UO_863 (O_863,N_13285,N_14595);
nor UO_864 (O_864,N_14161,N_13988);
or UO_865 (O_865,N_14427,N_14469);
or UO_866 (O_866,N_13378,N_14887);
xor UO_867 (O_867,N_13136,N_12055);
and UO_868 (O_868,N_14386,N_14000);
or UO_869 (O_869,N_13750,N_13695);
and UO_870 (O_870,N_12824,N_14167);
or UO_871 (O_871,N_14804,N_14082);
nand UO_872 (O_872,N_12466,N_14020);
nor UO_873 (O_873,N_13487,N_12677);
or UO_874 (O_874,N_14062,N_12493);
nand UO_875 (O_875,N_12332,N_14866);
nand UO_876 (O_876,N_14689,N_12029);
or UO_877 (O_877,N_14425,N_13083);
and UO_878 (O_878,N_13465,N_12695);
or UO_879 (O_879,N_14590,N_13732);
nand UO_880 (O_880,N_13823,N_12095);
and UO_881 (O_881,N_13565,N_12820);
or UO_882 (O_882,N_12711,N_14681);
or UO_883 (O_883,N_14009,N_12204);
xnor UO_884 (O_884,N_14236,N_13431);
or UO_885 (O_885,N_14839,N_12160);
nor UO_886 (O_886,N_13326,N_13175);
and UO_887 (O_887,N_14388,N_14656);
and UO_888 (O_888,N_13410,N_14898);
or UO_889 (O_889,N_13914,N_12540);
nand UO_890 (O_890,N_12447,N_14528);
or UO_891 (O_891,N_12149,N_14017);
nand UO_892 (O_892,N_13300,N_14420);
and UO_893 (O_893,N_13209,N_14085);
and UO_894 (O_894,N_12529,N_14015);
nor UO_895 (O_895,N_12577,N_13938);
and UO_896 (O_896,N_12661,N_13142);
and UO_897 (O_897,N_14049,N_12413);
nor UO_898 (O_898,N_12457,N_13805);
nand UO_899 (O_899,N_13892,N_12888);
nand UO_900 (O_900,N_14933,N_14319);
nand UO_901 (O_901,N_13296,N_14470);
or UO_902 (O_902,N_13574,N_12404);
or UO_903 (O_903,N_12373,N_12023);
or UO_904 (O_904,N_14787,N_12594);
nor UO_905 (O_905,N_13268,N_14916);
and UO_906 (O_906,N_14340,N_12135);
or UO_907 (O_907,N_13965,N_12973);
and UO_908 (O_908,N_13685,N_12030);
and UO_909 (O_909,N_14136,N_12936);
or UO_910 (O_910,N_12690,N_13273);
or UO_911 (O_911,N_12362,N_13100);
nand UO_912 (O_912,N_14982,N_14874);
or UO_913 (O_913,N_12182,N_12126);
nand UO_914 (O_914,N_12619,N_13837);
nor UO_915 (O_915,N_12963,N_12369);
and UO_916 (O_916,N_14345,N_12787);
nor UO_917 (O_917,N_14141,N_12219);
or UO_918 (O_918,N_14658,N_12191);
nor UO_919 (O_919,N_12061,N_12542);
nor UO_920 (O_920,N_14087,N_13145);
nor UO_921 (O_921,N_13428,N_14134);
nand UO_922 (O_922,N_14506,N_13606);
nand UO_923 (O_923,N_13375,N_13392);
nand UO_924 (O_924,N_14906,N_12208);
or UO_925 (O_925,N_12098,N_13537);
nor UO_926 (O_926,N_13162,N_13993);
nand UO_927 (O_927,N_13102,N_12289);
and UO_928 (O_928,N_12184,N_14258);
or UO_929 (O_929,N_14403,N_12264);
nand UO_930 (O_930,N_13315,N_13814);
nand UO_931 (O_931,N_14381,N_14695);
and UO_932 (O_932,N_14726,N_12730);
nor UO_933 (O_933,N_12303,N_12887);
nand UO_934 (O_934,N_14995,N_13481);
and UO_935 (O_935,N_12528,N_13262);
and UO_936 (O_936,N_13415,N_12359);
or UO_937 (O_937,N_13987,N_12341);
nor UO_938 (O_938,N_13449,N_12427);
and UO_939 (O_939,N_14784,N_13379);
nor UO_940 (O_940,N_12209,N_13345);
and UO_941 (O_941,N_14461,N_12013);
and UO_942 (O_942,N_14693,N_12465);
nand UO_943 (O_943,N_13835,N_14174);
and UO_944 (O_944,N_12940,N_13575);
or UO_945 (O_945,N_12125,N_14234);
nor UO_946 (O_946,N_14754,N_12751);
nand UO_947 (O_947,N_13236,N_13362);
or UO_948 (O_948,N_12386,N_12237);
and UO_949 (O_949,N_13323,N_14099);
nand UO_950 (O_950,N_12728,N_14931);
and UO_951 (O_951,N_12633,N_12069);
nand UO_952 (O_952,N_14123,N_14853);
xor UO_953 (O_953,N_13886,N_13135);
nand UO_954 (O_954,N_13853,N_13502);
nand UO_955 (O_955,N_12997,N_14249);
nor UO_956 (O_956,N_13317,N_12092);
xnor UO_957 (O_957,N_13567,N_13038);
or UO_958 (O_958,N_14169,N_12336);
or UO_959 (O_959,N_12731,N_13023);
nand UO_960 (O_960,N_12712,N_13253);
nand UO_961 (O_961,N_14243,N_13827);
and UO_962 (O_962,N_14318,N_12349);
nand UO_963 (O_963,N_12076,N_14325);
or UO_964 (O_964,N_13055,N_13227);
nor UO_965 (O_965,N_12210,N_12783);
or UO_966 (O_966,N_12977,N_14404);
nand UO_967 (O_967,N_12225,N_13725);
xor UO_968 (O_968,N_12866,N_14010);
nand UO_969 (O_969,N_14697,N_14793);
or UO_970 (O_970,N_14908,N_13104);
and UO_971 (O_971,N_14564,N_12937);
and UO_972 (O_972,N_13972,N_13946);
nor UO_973 (O_973,N_13346,N_13289);
or UO_974 (O_974,N_14512,N_13609);
and UO_975 (O_975,N_12700,N_13028);
and UO_976 (O_976,N_12390,N_14102);
nor UO_977 (O_977,N_14401,N_12474);
nor UO_978 (O_978,N_13177,N_12253);
and UO_979 (O_979,N_14905,N_12713);
and UO_980 (O_980,N_14068,N_13561);
nand UO_981 (O_981,N_13338,N_13438);
or UO_982 (O_982,N_13486,N_13959);
and UO_983 (O_983,N_14655,N_12475);
nor UO_984 (O_984,N_12350,N_12354);
nand UO_985 (O_985,N_14516,N_12423);
or UO_986 (O_986,N_12579,N_12863);
nand UO_987 (O_987,N_13003,N_14939);
and UO_988 (O_988,N_14121,N_12074);
or UO_989 (O_989,N_12662,N_14491);
nor UO_990 (O_990,N_14039,N_14396);
nand UO_991 (O_991,N_13257,N_12777);
and UO_992 (O_992,N_12504,N_13740);
nor UO_993 (O_993,N_14911,N_13139);
nor UO_994 (O_994,N_14510,N_14071);
nor UO_995 (O_995,N_12220,N_14662);
or UO_996 (O_996,N_14472,N_12114);
nand UO_997 (O_997,N_14703,N_13854);
nor UO_998 (O_998,N_12704,N_13920);
nand UO_999 (O_999,N_12609,N_12817);
or UO_1000 (O_1000,N_12639,N_12148);
nand UO_1001 (O_1001,N_13996,N_12473);
nand UO_1002 (O_1002,N_14454,N_12632);
and UO_1003 (O_1003,N_13693,N_12339);
or UO_1004 (O_1004,N_12026,N_12500);
nand UO_1005 (O_1005,N_12212,N_13334);
nor UO_1006 (O_1006,N_14806,N_14255);
nand UO_1007 (O_1007,N_13314,N_14437);
nand UO_1008 (O_1008,N_13616,N_14969);
nor UO_1009 (O_1009,N_13193,N_14475);
and UO_1010 (O_1010,N_12290,N_14837);
nor UO_1011 (O_1011,N_12328,N_13130);
or UO_1012 (O_1012,N_13847,N_13668);
xor UO_1013 (O_1013,N_14066,N_12421);
nand UO_1014 (O_1014,N_12456,N_12274);
nor UO_1015 (O_1015,N_12987,N_12926);
nand UO_1016 (O_1016,N_12159,N_14415);
nand UO_1017 (O_1017,N_13045,N_13472);
nor UO_1018 (O_1018,N_14164,N_14692);
nand UO_1019 (O_1019,N_13580,N_13366);
nor UO_1020 (O_1020,N_14687,N_14263);
or UO_1021 (O_1021,N_12676,N_12043);
and UO_1022 (O_1022,N_14817,N_13339);
nor UO_1023 (O_1023,N_14511,N_13307);
and UO_1024 (O_1024,N_13452,N_12988);
and UO_1025 (O_1025,N_13350,N_12093);
nand UO_1026 (O_1026,N_13215,N_13953);
or UO_1027 (O_1027,N_13160,N_12433);
nor UO_1028 (O_1028,N_12826,N_14038);
nand UO_1029 (O_1029,N_13112,N_12112);
nand UO_1030 (O_1030,N_14593,N_13430);
or UO_1031 (O_1031,N_12483,N_13077);
nor UO_1032 (O_1032,N_14252,N_14240);
and UO_1033 (O_1033,N_14442,N_14843);
or UO_1034 (O_1034,N_12990,N_13951);
or UO_1035 (O_1035,N_14796,N_13042);
nand UO_1036 (O_1036,N_13372,N_14393);
or UO_1037 (O_1037,N_12849,N_13087);
or UO_1038 (O_1038,N_12002,N_12735);
and UO_1039 (O_1039,N_14492,N_13763);
or UO_1040 (O_1040,N_13172,N_13394);
nor UO_1041 (O_1041,N_14713,N_14091);
nand UO_1042 (O_1042,N_12943,N_13911);
nand UO_1043 (O_1043,N_14989,N_12079);
nand UO_1044 (O_1044,N_13308,N_12365);
or UO_1045 (O_1045,N_12575,N_13021);
nor UO_1046 (O_1046,N_12681,N_14462);
or UO_1047 (O_1047,N_12960,N_13359);
nand UO_1048 (O_1048,N_13092,N_12276);
nor UO_1049 (O_1049,N_14165,N_13198);
or UO_1050 (O_1050,N_14097,N_14191);
or UO_1051 (O_1051,N_14616,N_14155);
and UO_1052 (O_1052,N_14148,N_13784);
or UO_1053 (O_1053,N_12010,N_14962);
or UO_1054 (O_1054,N_13233,N_13573);
and UO_1055 (O_1055,N_13568,N_12913);
and UO_1056 (O_1056,N_14749,N_12463);
nor UO_1057 (O_1057,N_12582,N_14643);
nand UO_1058 (O_1058,N_13396,N_14130);
nor UO_1059 (O_1059,N_12409,N_13444);
and UO_1060 (O_1060,N_14831,N_13484);
and UO_1061 (O_1061,N_12132,N_14076);
nor UO_1062 (O_1062,N_12334,N_13050);
nor UO_1063 (O_1063,N_12439,N_14077);
or UO_1064 (O_1064,N_13113,N_14923);
and UO_1065 (O_1065,N_12045,N_12629);
and UO_1066 (O_1066,N_14664,N_12522);
nand UO_1067 (O_1067,N_13185,N_12416);
nand UO_1068 (O_1068,N_12315,N_14951);
nand UO_1069 (O_1069,N_13358,N_12381);
or UO_1070 (O_1070,N_12755,N_14394);
nand UO_1071 (O_1071,N_12352,N_13680);
and UO_1072 (O_1072,N_14414,N_12986);
nor UO_1073 (O_1073,N_12889,N_12424);
or UO_1074 (O_1074,N_12312,N_13808);
nor UO_1075 (O_1075,N_13982,N_13639);
or UO_1076 (O_1076,N_13012,N_13910);
nand UO_1077 (O_1077,N_14972,N_14205);
and UO_1078 (O_1078,N_14646,N_12961);
nand UO_1079 (O_1079,N_14736,N_12122);
or UO_1080 (O_1080,N_14260,N_13599);
and UO_1081 (O_1081,N_14934,N_14545);
nor UO_1082 (O_1082,N_14628,N_13197);
and UO_1083 (O_1083,N_13194,N_14743);
nand UO_1084 (O_1084,N_14638,N_13771);
and UO_1085 (O_1085,N_12615,N_14525);
nand UO_1086 (O_1086,N_13794,N_14105);
or UO_1087 (O_1087,N_14031,N_13828);
nand UO_1088 (O_1088,N_12744,N_14847);
and UO_1089 (O_1089,N_14712,N_13922);
nor UO_1090 (O_1090,N_14521,N_13506);
nand UO_1091 (O_1091,N_14777,N_13980);
xnor UO_1092 (O_1092,N_12198,N_13459);
nand UO_1093 (O_1093,N_12019,N_12573);
xor UO_1094 (O_1094,N_13237,N_13776);
or UO_1095 (O_1095,N_13703,N_13751);
nor UO_1096 (O_1096,N_14782,N_13005);
or UO_1097 (O_1097,N_12203,N_14301);
nor UO_1098 (O_1098,N_12882,N_13974);
or UO_1099 (O_1099,N_13807,N_12950);
or UO_1100 (O_1100,N_12746,N_13787);
or UO_1101 (O_1101,N_14901,N_12497);
nor UO_1102 (O_1102,N_12121,N_12519);
and UO_1103 (O_1103,N_14217,N_14775);
or UO_1104 (O_1104,N_13884,N_13534);
nand UO_1105 (O_1105,N_14636,N_12382);
and UO_1106 (O_1106,N_12890,N_12078);
nand UO_1107 (O_1107,N_12037,N_14811);
or UO_1108 (O_1108,N_13240,N_12399);
and UO_1109 (O_1109,N_14924,N_14998);
and UO_1110 (O_1110,N_12278,N_12254);
nand UO_1111 (O_1111,N_13895,N_13615);
and UO_1112 (O_1112,N_14543,N_14448);
nor UO_1113 (O_1113,N_12171,N_14135);
and UO_1114 (O_1114,N_14253,N_13390);
and UO_1115 (O_1115,N_12654,N_13947);
nand UO_1116 (O_1116,N_12011,N_12837);
nor UO_1117 (O_1117,N_14337,N_13034);
nor UO_1118 (O_1118,N_13793,N_13931);
and UO_1119 (O_1119,N_14316,N_13224);
nand UO_1120 (O_1120,N_12393,N_12917);
nor UO_1121 (O_1121,N_14809,N_14778);
nand UO_1122 (O_1122,N_13060,N_12379);
nor UO_1123 (O_1123,N_14718,N_12086);
and UO_1124 (O_1124,N_13052,N_13364);
nand UO_1125 (O_1125,N_12286,N_13169);
and UO_1126 (O_1126,N_12458,N_14432);
nand UO_1127 (O_1127,N_14173,N_14832);
nor UO_1128 (O_1128,N_12898,N_12324);
or UO_1129 (O_1129,N_14555,N_14244);
nor UO_1130 (O_1130,N_12518,N_13877);
or UO_1131 (O_1131,N_12930,N_14860);
nor UO_1132 (O_1132,N_14093,N_14988);
or UO_1133 (O_1133,N_14977,N_14522);
nand UO_1134 (O_1134,N_12739,N_13512);
or UO_1135 (O_1135,N_12658,N_12517);
and UO_1136 (O_1136,N_14802,N_12765);
or UO_1137 (O_1137,N_14160,N_13329);
nand UO_1138 (O_1138,N_12796,N_13697);
and UO_1139 (O_1139,N_12666,N_12355);
nor UO_1140 (O_1140,N_13228,N_14928);
nand UO_1141 (O_1141,N_14548,N_14585);
nand UO_1142 (O_1142,N_13090,N_14490);
or UO_1143 (O_1143,N_14974,N_14735);
or UO_1144 (O_1144,N_12486,N_12107);
and UO_1145 (O_1145,N_14710,N_13729);
nand UO_1146 (O_1146,N_13058,N_14848);
nor UO_1147 (O_1147,N_12780,N_12537);
or UO_1148 (O_1148,N_14245,N_14430);
or UO_1149 (O_1149,N_13578,N_13509);
and UO_1150 (O_1150,N_12047,N_14986);
or UO_1151 (O_1151,N_13382,N_13547);
nand UO_1152 (O_1152,N_14344,N_13202);
or UO_1153 (O_1153,N_13164,N_14079);
nor UO_1154 (O_1154,N_12320,N_14447);
and UO_1155 (O_1155,N_14157,N_13839);
nand UO_1156 (O_1156,N_14586,N_12428);
or UO_1157 (O_1157,N_13833,N_12834);
nor UO_1158 (O_1158,N_14514,N_12902);
xnor UO_1159 (O_1159,N_13204,N_14237);
nand UO_1160 (O_1160,N_13674,N_13882);
and UO_1161 (O_1161,N_14767,N_14882);
nand UO_1162 (O_1162,N_12831,N_12391);
and UO_1163 (O_1163,N_13861,N_13614);
nand UO_1164 (O_1164,N_14873,N_13451);
and UO_1165 (O_1165,N_14594,N_13726);
or UO_1166 (O_1166,N_13037,N_14706);
or UO_1167 (O_1167,N_14508,N_13196);
or UO_1168 (O_1168,N_14149,N_12626);
or UO_1169 (O_1169,N_13505,N_14112);
and UO_1170 (O_1170,N_12089,N_14606);
nor UO_1171 (O_1171,N_12880,N_14762);
and UO_1172 (O_1172,N_13878,N_14880);
and UO_1173 (O_1173,N_14558,N_13694);
or UO_1174 (O_1174,N_13738,N_13316);
or UO_1175 (O_1175,N_13815,N_13155);
or UO_1176 (O_1176,N_13928,N_12808);
nand UO_1177 (O_1177,N_14321,N_14729);
nand UO_1178 (O_1178,N_13349,N_12620);
or UO_1179 (O_1179,N_12682,N_12651);
or UO_1180 (O_1180,N_14856,N_13200);
and UO_1181 (O_1181,N_12722,N_12036);
and UO_1182 (O_1182,N_14584,N_14570);
and UO_1183 (O_1183,N_12192,N_14705);
nand UO_1184 (O_1184,N_12679,N_12340);
nor UO_1185 (O_1185,N_12060,N_13399);
nand UO_1186 (O_1186,N_12257,N_13259);
or UO_1187 (O_1187,N_13712,N_13948);
nand UO_1188 (O_1188,N_13476,N_14504);
and UO_1189 (O_1189,N_13179,N_12665);
and UO_1190 (O_1190,N_12211,N_12610);
or UO_1191 (O_1191,N_14003,N_13960);
and UO_1192 (O_1192,N_13409,N_14333);
or UO_1193 (O_1193,N_13341,N_14142);
nand UO_1194 (O_1194,N_13605,N_12177);
nand UO_1195 (O_1195,N_14707,N_14714);
and UO_1196 (O_1196,N_13287,N_13739);
nor UO_1197 (O_1197,N_13983,N_12688);
or UO_1198 (O_1198,N_14265,N_12081);
or UO_1199 (O_1199,N_12134,N_13799);
and UO_1200 (O_1200,N_14269,N_14012);
nand UO_1201 (O_1201,N_14611,N_12407);
and UO_1202 (O_1202,N_13533,N_13434);
or UO_1203 (O_1203,N_14276,N_12981);
nor UO_1204 (O_1204,N_12847,N_14881);
nor UO_1205 (O_1205,N_14973,N_12265);
nand UO_1206 (O_1206,N_14006,N_14883);
or UO_1207 (O_1207,N_14391,N_12674);
nor UO_1208 (O_1208,N_13384,N_13905);
and UO_1209 (O_1209,N_14766,N_13447);
or UO_1210 (O_1210,N_12412,N_13491);
or UO_1211 (O_1211,N_12800,N_12371);
nor UO_1212 (O_1212,N_13067,N_13842);
nand UO_1213 (O_1213,N_13613,N_13711);
or UO_1214 (O_1214,N_13176,N_13720);
nand UO_1215 (O_1215,N_13899,N_13439);
nand UO_1216 (O_1216,N_13975,N_13957);
and UO_1217 (O_1217,N_14416,N_13101);
and UO_1218 (O_1218,N_14059,N_12724);
xnor UO_1219 (O_1219,N_14737,N_12316);
nor UO_1220 (O_1220,N_12335,N_13998);
nor UO_1221 (O_1221,N_12411,N_12269);
and UO_1222 (O_1222,N_14801,N_12822);
and UO_1223 (O_1223,N_14317,N_12685);
nor UO_1224 (O_1224,N_12377,N_13696);
nor UO_1225 (O_1225,N_13412,N_14090);
nand UO_1226 (O_1226,N_14221,N_14612);
or UO_1227 (O_1227,N_12075,N_14670);
or UO_1228 (O_1228,N_12218,N_12657);
and UO_1229 (O_1229,N_13085,N_14559);
nor UO_1230 (O_1230,N_12905,N_14145);
nor UO_1231 (O_1231,N_12464,N_12509);
and UO_1232 (O_1232,N_13327,N_13939);
or UO_1233 (O_1233,N_13754,N_13549);
nand UO_1234 (O_1234,N_12073,N_14158);
nor UO_1235 (O_1235,N_13716,N_14250);
or UO_1236 (O_1236,N_12586,N_13553);
nand UO_1237 (O_1237,N_14684,N_13525);
nand UO_1238 (O_1238,N_12048,N_14770);
and UO_1239 (O_1239,N_12995,N_13926);
and UO_1240 (O_1240,N_13031,N_13254);
and UO_1241 (O_1241,N_12754,N_12351);
nand UO_1242 (O_1242,N_13722,N_12058);
and UO_1243 (O_1243,N_13723,N_14921);
nor UO_1244 (O_1244,N_12372,N_13556);
or UO_1245 (O_1245,N_12983,N_13482);
and UO_1246 (O_1246,N_12852,N_13246);
and UO_1247 (O_1247,N_14211,N_14147);
and UO_1248 (O_1248,N_13226,N_12097);
nand UO_1249 (O_1249,N_13475,N_12894);
or UO_1250 (O_1250,N_12453,N_13992);
or UO_1251 (O_1251,N_12563,N_13968);
or UO_1252 (O_1252,N_14498,N_14070);
or UO_1253 (O_1253,N_12559,N_12745);
nand UO_1254 (O_1254,N_14675,N_12564);
nor UO_1255 (O_1255,N_13011,N_12871);
nor UO_1256 (O_1256,N_13802,N_12109);
or UO_1257 (O_1257,N_14107,N_13071);
and UO_1258 (O_1258,N_12426,N_13679);
or UO_1259 (O_1259,N_13997,N_14045);
or UO_1260 (O_1260,N_13964,N_12164);
nor UO_1261 (O_1261,N_12038,N_13851);
nor UO_1262 (O_1262,N_13004,N_13588);
nor UO_1263 (O_1263,N_12611,N_14114);
and UO_1264 (O_1264,N_14579,N_12216);
xnor UO_1265 (O_1265,N_14598,N_13041);
nand UO_1266 (O_1266,N_13015,N_12035);
nand UO_1267 (O_1267,N_14875,N_12813);
nand UO_1268 (O_1268,N_13448,N_12153);
and UO_1269 (O_1269,N_14960,N_13904);
and UO_1270 (O_1270,N_12150,N_13663);
nor UO_1271 (O_1271,N_13949,N_14235);
or UO_1272 (O_1272,N_14722,N_12992);
nor UO_1273 (O_1273,N_13956,N_12039);
and UO_1274 (O_1274,N_12555,N_12053);
nand UO_1275 (O_1275,N_14800,N_14153);
nor UO_1276 (O_1276,N_12527,N_13342);
or UO_1277 (O_1277,N_12904,N_14226);
nor UO_1278 (O_1278,N_13265,N_14146);
nor UO_1279 (O_1279,N_12968,N_14362);
or UO_1280 (O_1280,N_14109,N_14940);
and UO_1281 (O_1281,N_12205,N_13976);
nand UO_1282 (O_1282,N_12557,N_14699);
or UO_1283 (O_1283,N_13149,N_12297);
or UO_1284 (O_1284,N_13391,N_14851);
nand UO_1285 (O_1285,N_12590,N_14958);
and UO_1286 (O_1286,N_14104,N_13062);
nor UO_1287 (O_1287,N_12843,N_13450);
nor UO_1288 (O_1288,N_12176,N_13234);
nand UO_1289 (O_1289,N_13686,N_13128);
nand UO_1290 (O_1290,N_14369,N_14691);
nor UO_1291 (O_1291,N_12050,N_14750);
or UO_1292 (O_1292,N_13422,N_13971);
and UO_1293 (O_1293,N_12970,N_12481);
nor UO_1294 (O_1294,N_13538,N_12115);
or UO_1295 (O_1295,N_12167,N_12360);
nor UO_1296 (O_1296,N_14246,N_14443);
nor UO_1297 (O_1297,N_12868,N_14517);
and UO_1298 (O_1298,N_12884,N_12972);
or UO_1299 (O_1299,N_13894,N_14768);
nor UO_1300 (O_1300,N_14668,N_14577);
or UO_1301 (O_1301,N_13493,N_14925);
or UO_1302 (O_1302,N_12964,N_12921);
nand UO_1303 (O_1303,N_14761,N_13800);
or UO_1304 (O_1304,N_14685,N_12082);
nand UO_1305 (O_1305,N_13126,N_12140);
and UO_1306 (O_1306,N_14535,N_14241);
and UO_1307 (O_1307,N_13357,N_12969);
or UO_1308 (O_1308,N_12891,N_14297);
nand UO_1309 (O_1309,N_14054,N_12587);
or UO_1310 (O_1310,N_13602,N_12065);
and UO_1311 (O_1311,N_12033,N_13420);
and UO_1312 (O_1312,N_14298,N_13097);
nor UO_1313 (O_1313,N_12673,N_14580);
xor UO_1314 (O_1314,N_14175,N_14629);
or UO_1315 (O_1315,N_13368,N_12008);
nor UO_1316 (O_1316,N_13074,N_13433);
nor UO_1317 (O_1317,N_13306,N_13192);
nor UO_1318 (O_1318,N_14429,N_14287);
nand UO_1319 (O_1319,N_13029,N_14872);
or UO_1320 (O_1320,N_14871,N_13414);
nand UO_1321 (O_1321,N_14659,N_12267);
or UO_1322 (O_1322,N_14021,N_14456);
nand UO_1323 (O_1323,N_13363,N_14641);
nand UO_1324 (O_1324,N_12758,N_12967);
or UO_1325 (O_1325,N_12636,N_14868);
nand UO_1326 (O_1326,N_14620,N_14267);
and UO_1327 (O_1327,N_12539,N_14502);
nor UO_1328 (O_1328,N_12767,N_14835);
nand UO_1329 (O_1329,N_13151,N_12900);
nand UO_1330 (O_1330,N_14494,N_14342);
nor UO_1331 (O_1331,N_14700,N_14672);
nand UO_1332 (O_1332,N_12017,N_14151);
or UO_1333 (O_1333,N_13510,N_13473);
and UO_1334 (O_1334,N_12919,N_14144);
and UO_1335 (O_1335,N_12338,N_14037);
or UO_1336 (O_1336,N_12592,N_12358);
nand UO_1337 (O_1337,N_12956,N_12233);
nor UO_1338 (O_1338,N_13540,N_13404);
or UO_1339 (O_1339,N_14617,N_13570);
xor UO_1340 (O_1340,N_13524,N_12811);
nor UO_1341 (O_1341,N_14270,N_14125);
or UO_1342 (O_1342,N_13801,N_13628);
nand UO_1343 (O_1343,N_14463,N_13250);
nor UO_1344 (O_1344,N_14206,N_12578);
nand UO_1345 (O_1345,N_13201,N_13520);
or UO_1346 (O_1346,N_14682,N_13000);
and UO_1347 (O_1347,N_14987,N_12151);
or UO_1348 (O_1348,N_13889,N_12922);
and UO_1349 (O_1349,N_12568,N_14889);
or UO_1350 (O_1350,N_12874,N_12684);
and UO_1351 (O_1351,N_14405,N_13764);
nand UO_1352 (O_1352,N_13373,N_13994);
nor UO_1353 (O_1353,N_13355,N_13118);
nand UO_1354 (O_1354,N_12161,N_14857);
nand UO_1355 (O_1355,N_12585,N_14190);
and UO_1356 (O_1356,N_14980,N_12201);
nor UO_1357 (O_1357,N_13791,N_13558);
and UO_1358 (O_1358,N_13528,N_13159);
nor UO_1359 (O_1359,N_13618,N_13076);
nor UO_1360 (O_1360,N_12933,N_12512);
xnor UO_1361 (O_1361,N_13810,N_13251);
nand UO_1362 (O_1362,N_12867,N_14623);
nand UO_1363 (O_1363,N_12478,N_14055);
and UO_1364 (O_1364,N_13500,N_13001);
nor UO_1365 (O_1365,N_13554,N_14348);
xnor UO_1366 (O_1366,N_12523,N_14961);
and UO_1367 (O_1367,N_14552,N_13263);
nor UO_1368 (O_1368,N_14788,N_13302);
or UO_1369 (O_1369,N_13535,N_14518);
or UO_1370 (O_1370,N_13627,N_14004);
nand UO_1371 (O_1371,N_13593,N_14869);
or UO_1372 (O_1372,N_13065,N_12397);
or UO_1373 (O_1373,N_12281,N_13010);
nand UO_1374 (O_1374,N_14106,N_14439);
or UO_1375 (O_1375,N_12323,N_14207);
or UO_1376 (O_1376,N_12387,N_14310);
or UO_1377 (O_1377,N_13072,N_14272);
nor UO_1378 (O_1378,N_14841,N_12718);
nor UO_1379 (O_1379,N_12313,N_14821);
nand UO_1380 (O_1380,N_14696,N_13542);
or UO_1381 (O_1381,N_13369,N_13406);
and UO_1382 (O_1382,N_13498,N_13401);
nand UO_1383 (O_1383,N_12683,N_13687);
or UO_1384 (O_1384,N_13462,N_12976);
xor UO_1385 (O_1385,N_13095,N_13181);
nand UO_1386 (O_1386,N_12942,N_14651);
nor UO_1387 (O_1387,N_13210,N_12308);
nand UO_1388 (O_1388,N_12669,N_12878);
or UO_1389 (O_1389,N_12169,N_12105);
and UO_1390 (O_1390,N_14551,N_13898);
nand UO_1391 (O_1391,N_13560,N_12670);
or UO_1392 (O_1392,N_14567,N_13152);
and UO_1393 (O_1393,N_14642,N_14648);
and UO_1394 (O_1394,N_14935,N_12370);
nor UO_1395 (O_1395,N_12356,N_13398);
nand UO_1396 (O_1396,N_12506,N_14384);
nand UO_1397 (O_1397,N_14223,N_14312);
nor UO_1398 (O_1398,N_12127,N_12417);
and UO_1399 (O_1399,N_13293,N_12782);
nor UO_1400 (O_1400,N_14088,N_14300);
or UO_1401 (O_1401,N_12733,N_12723);
nand UO_1402 (O_1402,N_14554,N_13523);
nor UO_1403 (O_1403,N_12678,N_12091);
nor UO_1404 (O_1404,N_12915,N_12513);
and UO_1405 (O_1405,N_14776,N_13456);
or UO_1406 (O_1406,N_13312,N_12934);
nand UO_1407 (O_1407,N_12571,N_12236);
nor UO_1408 (O_1408,N_13852,N_12106);
and UO_1409 (O_1409,N_13587,N_12494);
nor UO_1410 (O_1410,N_12446,N_13676);
or UO_1411 (O_1411,N_14370,N_14182);
nand UO_1412 (O_1412,N_12242,N_14280);
and UO_1413 (O_1413,N_12634,N_13518);
or UO_1414 (O_1414,N_13569,N_12779);
nor UO_1415 (O_1415,N_13383,N_13955);
and UO_1416 (O_1416,N_12895,N_14120);
nand UO_1417 (O_1417,N_12495,N_12721);
and UO_1418 (O_1418,N_12228,N_12034);
and UO_1419 (O_1419,N_12966,N_14678);
nand UO_1420 (O_1420,N_12989,N_13230);
or UO_1421 (O_1421,N_12671,N_12645);
and UO_1422 (O_1422,N_13222,N_14920);
or UO_1423 (O_1423,N_12792,N_12823);
nor UO_1424 (O_1424,N_12786,N_12307);
or UO_1425 (O_1425,N_13849,N_12583);
nand UO_1426 (O_1426,N_14769,N_13846);
nor UO_1427 (O_1427,N_13110,N_12450);
and UO_1428 (O_1428,N_13243,N_14094);
and UO_1429 (O_1429,N_14912,N_12068);
nand UO_1430 (O_1430,N_14382,N_12505);
nand UO_1431 (O_1431,N_13127,N_14201);
or UO_1432 (O_1432,N_14968,N_13047);
nor UO_1433 (O_1433,N_13532,N_13469);
nor UO_1434 (O_1434,N_13173,N_13319);
nor UO_1435 (O_1435,N_13387,N_13866);
nor UO_1436 (O_1436,N_13806,N_14765);
nand UO_1437 (O_1437,N_13504,N_14615);
nand UO_1438 (O_1438,N_12022,N_12910);
xnor UO_1439 (O_1439,N_14385,N_14957);
or UO_1440 (O_1440,N_12740,N_13403);
nand UO_1441 (O_1441,N_14483,N_12044);
nand UO_1442 (O_1442,N_14539,N_13879);
nor UO_1443 (O_1443,N_12872,N_12432);
nand UO_1444 (O_1444,N_13705,N_13795);
nor UO_1445 (O_1445,N_14360,N_12565);
nor UO_1446 (O_1446,N_12124,N_14953);
or UO_1447 (O_1447,N_12277,N_13084);
or UO_1448 (O_1448,N_12772,N_12551);
and UO_1449 (O_1449,N_14556,N_13292);
or UO_1450 (O_1450,N_14992,N_13514);
or UO_1451 (O_1451,N_13913,N_13659);
nor UO_1452 (O_1452,N_13779,N_14541);
nor UO_1453 (O_1453,N_14238,N_13572);
nand UO_1454 (O_1454,N_12924,N_13718);
nand UO_1455 (O_1455,N_14024,N_13107);
nand UO_1456 (O_1456,N_14192,N_12534);
nor UO_1457 (O_1457,N_14214,N_13131);
nor UO_1458 (O_1458,N_13408,N_13908);
nor UO_1459 (O_1459,N_14581,N_14915);
and UO_1460 (O_1460,N_14878,N_12374);
and UO_1461 (O_1461,N_13223,N_13079);
nand UO_1462 (O_1462,N_13648,N_14030);
or UO_1463 (O_1463,N_13099,N_14410);
nor UO_1464 (O_1464,N_12123,N_14473);
or UO_1465 (O_1465,N_13954,N_13921);
nor UO_1466 (O_1466,N_14613,N_12854);
and UO_1467 (O_1467,N_13303,N_12797);
or UO_1468 (O_1468,N_14626,N_12957);
nor UO_1469 (O_1469,N_14320,N_14833);
nand UO_1470 (O_1470,N_14760,N_13436);
and UO_1471 (O_1471,N_12794,N_12110);
or UO_1472 (O_1472,N_12879,N_12899);
or UO_1473 (O_1473,N_12490,N_14639);
nand UO_1474 (O_1474,N_13966,N_12601);
nor UO_1475 (O_1475,N_14061,N_13463);
nor UO_1476 (O_1476,N_14133,N_12952);
and UO_1477 (O_1477,N_12747,N_12345);
and UO_1478 (O_1478,N_12018,N_13656);
nand UO_1479 (O_1479,N_14008,N_13873);
nor UO_1480 (O_1480,N_12949,N_13919);
or UO_1481 (O_1481,N_12480,N_13144);
nor UO_1482 (O_1482,N_12410,N_13706);
nor UO_1483 (O_1483,N_14649,N_13607);
nor UO_1484 (O_1484,N_13024,N_14110);
or UO_1485 (O_1485,N_12507,N_12066);
nor UO_1486 (O_1486,N_14446,N_12829);
nand UO_1487 (O_1487,N_12597,N_13531);
nor UO_1488 (O_1488,N_13281,N_14479);
and UO_1489 (O_1489,N_14709,N_13758);
or UO_1490 (O_1490,N_13275,N_14261);
nand UO_1491 (O_1491,N_13667,N_13054);
nor UO_1492 (O_1492,N_13881,N_12299);
and UO_1493 (O_1493,N_14529,N_14036);
nand UO_1494 (O_1494,N_12119,N_12750);
nand UO_1495 (O_1495,N_12860,N_12263);
nor UO_1496 (O_1496,N_13400,N_14116);
nand UO_1497 (O_1497,N_12520,N_14597);
and UO_1498 (O_1498,N_14202,N_13769);
and UO_1499 (O_1499,N_13617,N_13859);
nor UO_1500 (O_1500,N_13094,N_12570);
nor UO_1501 (O_1501,N_12641,N_12652);
and UO_1502 (O_1502,N_12248,N_13610);
nand UO_1503 (O_1503,N_13950,N_14997);
nand UO_1504 (O_1504,N_14034,N_12848);
and UO_1505 (O_1505,N_12071,N_12419);
nand UO_1506 (O_1506,N_13499,N_14442);
and UO_1507 (O_1507,N_13677,N_13988);
nand UO_1508 (O_1508,N_14409,N_14128);
or UO_1509 (O_1509,N_12802,N_14810);
nand UO_1510 (O_1510,N_12282,N_14096);
or UO_1511 (O_1511,N_13540,N_13050);
xnor UO_1512 (O_1512,N_14541,N_12931);
nor UO_1513 (O_1513,N_12263,N_12581);
nor UO_1514 (O_1514,N_12643,N_12058);
nand UO_1515 (O_1515,N_13572,N_13965);
nand UO_1516 (O_1516,N_12490,N_12676);
nand UO_1517 (O_1517,N_14079,N_14217);
and UO_1518 (O_1518,N_12885,N_14233);
nor UO_1519 (O_1519,N_14544,N_12853);
nor UO_1520 (O_1520,N_12400,N_14325);
nand UO_1521 (O_1521,N_14470,N_13303);
nor UO_1522 (O_1522,N_13987,N_14747);
nand UO_1523 (O_1523,N_14243,N_13848);
nand UO_1524 (O_1524,N_14224,N_13872);
nor UO_1525 (O_1525,N_14897,N_14313);
and UO_1526 (O_1526,N_12580,N_12125);
nor UO_1527 (O_1527,N_14436,N_13467);
nand UO_1528 (O_1528,N_12574,N_13340);
nor UO_1529 (O_1529,N_14084,N_13418);
or UO_1530 (O_1530,N_12120,N_14922);
nor UO_1531 (O_1531,N_12936,N_12070);
or UO_1532 (O_1532,N_13497,N_14345);
nand UO_1533 (O_1533,N_13322,N_14906);
nand UO_1534 (O_1534,N_12671,N_14364);
or UO_1535 (O_1535,N_12574,N_14538);
and UO_1536 (O_1536,N_14130,N_13876);
nand UO_1537 (O_1537,N_13131,N_13280);
and UO_1538 (O_1538,N_14704,N_14816);
nor UO_1539 (O_1539,N_12482,N_14666);
nor UO_1540 (O_1540,N_13562,N_14165);
nand UO_1541 (O_1541,N_14312,N_12922);
nand UO_1542 (O_1542,N_14877,N_14992);
or UO_1543 (O_1543,N_12881,N_12217);
nand UO_1544 (O_1544,N_14129,N_12631);
nor UO_1545 (O_1545,N_13228,N_12388);
nand UO_1546 (O_1546,N_12383,N_14197);
nor UO_1547 (O_1547,N_14989,N_12873);
nand UO_1548 (O_1548,N_12946,N_14078);
nand UO_1549 (O_1549,N_12821,N_12604);
nand UO_1550 (O_1550,N_14770,N_14375);
or UO_1551 (O_1551,N_14458,N_13616);
and UO_1552 (O_1552,N_12638,N_13301);
nor UO_1553 (O_1553,N_13115,N_13387);
and UO_1554 (O_1554,N_13137,N_12190);
and UO_1555 (O_1555,N_12275,N_13536);
nand UO_1556 (O_1556,N_14812,N_14552);
nor UO_1557 (O_1557,N_12781,N_13061);
nor UO_1558 (O_1558,N_12897,N_13559);
or UO_1559 (O_1559,N_13872,N_12463);
and UO_1560 (O_1560,N_14514,N_12005);
xnor UO_1561 (O_1561,N_12650,N_12181);
and UO_1562 (O_1562,N_12616,N_14568);
or UO_1563 (O_1563,N_13975,N_12915);
nor UO_1564 (O_1564,N_14811,N_14890);
nor UO_1565 (O_1565,N_13787,N_12703);
or UO_1566 (O_1566,N_12304,N_13117);
and UO_1567 (O_1567,N_13725,N_14986);
nand UO_1568 (O_1568,N_14749,N_12170);
nor UO_1569 (O_1569,N_14285,N_12824);
and UO_1570 (O_1570,N_12588,N_12545);
nor UO_1571 (O_1571,N_12627,N_12688);
nor UO_1572 (O_1572,N_12818,N_14646);
nor UO_1573 (O_1573,N_12930,N_12621);
nor UO_1574 (O_1574,N_14492,N_14171);
and UO_1575 (O_1575,N_12164,N_14985);
nor UO_1576 (O_1576,N_12857,N_14239);
or UO_1577 (O_1577,N_14511,N_14751);
nand UO_1578 (O_1578,N_14181,N_12499);
nor UO_1579 (O_1579,N_14907,N_13488);
nor UO_1580 (O_1580,N_12318,N_13280);
or UO_1581 (O_1581,N_12819,N_12237);
or UO_1582 (O_1582,N_12909,N_12541);
or UO_1583 (O_1583,N_14469,N_14683);
and UO_1584 (O_1584,N_12009,N_13828);
nor UO_1585 (O_1585,N_12386,N_14601);
nor UO_1586 (O_1586,N_13369,N_14410);
nor UO_1587 (O_1587,N_12286,N_12666);
and UO_1588 (O_1588,N_14088,N_13390);
nand UO_1589 (O_1589,N_13289,N_14908);
nor UO_1590 (O_1590,N_13404,N_14745);
nor UO_1591 (O_1591,N_13449,N_12039);
and UO_1592 (O_1592,N_12711,N_12047);
and UO_1593 (O_1593,N_14739,N_13930);
or UO_1594 (O_1594,N_12102,N_12147);
nor UO_1595 (O_1595,N_13121,N_12435);
or UO_1596 (O_1596,N_12730,N_13630);
nand UO_1597 (O_1597,N_12620,N_12393);
and UO_1598 (O_1598,N_14451,N_12454);
and UO_1599 (O_1599,N_12142,N_12686);
nor UO_1600 (O_1600,N_14266,N_13036);
nor UO_1601 (O_1601,N_14232,N_14312);
nand UO_1602 (O_1602,N_12712,N_14764);
nor UO_1603 (O_1603,N_14198,N_14990);
and UO_1604 (O_1604,N_13575,N_14312);
or UO_1605 (O_1605,N_12373,N_12367);
or UO_1606 (O_1606,N_12670,N_12338);
and UO_1607 (O_1607,N_13653,N_13056);
and UO_1608 (O_1608,N_13573,N_14765);
nor UO_1609 (O_1609,N_12732,N_12124);
nand UO_1610 (O_1610,N_14826,N_13230);
or UO_1611 (O_1611,N_12590,N_14796);
nand UO_1612 (O_1612,N_14716,N_13145);
and UO_1613 (O_1613,N_12321,N_13963);
or UO_1614 (O_1614,N_12959,N_13523);
or UO_1615 (O_1615,N_13387,N_14407);
nor UO_1616 (O_1616,N_12918,N_13498);
nor UO_1617 (O_1617,N_14991,N_14798);
or UO_1618 (O_1618,N_13776,N_13768);
and UO_1619 (O_1619,N_13595,N_12513);
or UO_1620 (O_1620,N_12877,N_13194);
or UO_1621 (O_1621,N_13647,N_14112);
or UO_1622 (O_1622,N_13203,N_13223);
nand UO_1623 (O_1623,N_14100,N_14200);
nor UO_1624 (O_1624,N_12480,N_14595);
or UO_1625 (O_1625,N_12944,N_12171);
or UO_1626 (O_1626,N_12120,N_13391);
nor UO_1627 (O_1627,N_12311,N_14671);
nor UO_1628 (O_1628,N_14360,N_12951);
nand UO_1629 (O_1629,N_12581,N_14114);
nand UO_1630 (O_1630,N_13382,N_14538);
nor UO_1631 (O_1631,N_13622,N_14652);
or UO_1632 (O_1632,N_13797,N_13296);
nor UO_1633 (O_1633,N_12632,N_14613);
nand UO_1634 (O_1634,N_12780,N_14741);
nand UO_1635 (O_1635,N_14353,N_13202);
or UO_1636 (O_1636,N_12566,N_13277);
and UO_1637 (O_1637,N_14689,N_14169);
nand UO_1638 (O_1638,N_12531,N_14217);
or UO_1639 (O_1639,N_14220,N_12615);
nand UO_1640 (O_1640,N_14937,N_13900);
and UO_1641 (O_1641,N_13774,N_14204);
or UO_1642 (O_1642,N_14050,N_13167);
nor UO_1643 (O_1643,N_14708,N_14050);
nor UO_1644 (O_1644,N_12586,N_14230);
or UO_1645 (O_1645,N_13784,N_12246);
and UO_1646 (O_1646,N_13614,N_13212);
and UO_1647 (O_1647,N_13580,N_12229);
nor UO_1648 (O_1648,N_14145,N_13851);
and UO_1649 (O_1649,N_14295,N_12819);
and UO_1650 (O_1650,N_12778,N_12618);
and UO_1651 (O_1651,N_12098,N_13571);
nor UO_1652 (O_1652,N_13262,N_12826);
or UO_1653 (O_1653,N_14444,N_12134);
or UO_1654 (O_1654,N_12196,N_13261);
nor UO_1655 (O_1655,N_14268,N_12144);
and UO_1656 (O_1656,N_12025,N_13511);
and UO_1657 (O_1657,N_13978,N_12168);
and UO_1658 (O_1658,N_12319,N_12617);
and UO_1659 (O_1659,N_12865,N_14073);
and UO_1660 (O_1660,N_13269,N_13633);
and UO_1661 (O_1661,N_12440,N_13506);
nand UO_1662 (O_1662,N_13290,N_14947);
or UO_1663 (O_1663,N_14401,N_12565);
and UO_1664 (O_1664,N_12261,N_12944);
or UO_1665 (O_1665,N_12065,N_14330);
xnor UO_1666 (O_1666,N_14619,N_14518);
nand UO_1667 (O_1667,N_12211,N_14019);
nor UO_1668 (O_1668,N_13915,N_14065);
or UO_1669 (O_1669,N_12199,N_12703);
and UO_1670 (O_1670,N_14051,N_13563);
nor UO_1671 (O_1671,N_14206,N_14260);
nor UO_1672 (O_1672,N_13218,N_12878);
nor UO_1673 (O_1673,N_12395,N_12706);
or UO_1674 (O_1674,N_14265,N_13936);
and UO_1675 (O_1675,N_13436,N_12110);
nand UO_1676 (O_1676,N_12684,N_14032);
or UO_1677 (O_1677,N_14607,N_13436);
and UO_1678 (O_1678,N_14031,N_12648);
nor UO_1679 (O_1679,N_13968,N_14456);
or UO_1680 (O_1680,N_12787,N_12936);
and UO_1681 (O_1681,N_12979,N_12019);
nor UO_1682 (O_1682,N_14239,N_12163);
and UO_1683 (O_1683,N_14935,N_13534);
nor UO_1684 (O_1684,N_14765,N_14973);
or UO_1685 (O_1685,N_13720,N_14356);
nand UO_1686 (O_1686,N_14469,N_13353);
nand UO_1687 (O_1687,N_12905,N_12388);
or UO_1688 (O_1688,N_14090,N_13157);
nand UO_1689 (O_1689,N_14041,N_14811);
or UO_1690 (O_1690,N_13712,N_14749);
and UO_1691 (O_1691,N_12178,N_14378);
or UO_1692 (O_1692,N_14028,N_14516);
nand UO_1693 (O_1693,N_14996,N_13258);
and UO_1694 (O_1694,N_12434,N_12577);
nand UO_1695 (O_1695,N_12605,N_14890);
nor UO_1696 (O_1696,N_12169,N_12542);
and UO_1697 (O_1697,N_13301,N_14413);
or UO_1698 (O_1698,N_13452,N_12770);
nand UO_1699 (O_1699,N_14150,N_14098);
nand UO_1700 (O_1700,N_14003,N_14374);
or UO_1701 (O_1701,N_12295,N_12149);
and UO_1702 (O_1702,N_13293,N_14343);
nor UO_1703 (O_1703,N_13004,N_14309);
nor UO_1704 (O_1704,N_13311,N_13082);
nor UO_1705 (O_1705,N_12228,N_12977);
xnor UO_1706 (O_1706,N_13127,N_12345);
and UO_1707 (O_1707,N_12948,N_12613);
nor UO_1708 (O_1708,N_14904,N_13399);
nand UO_1709 (O_1709,N_14152,N_14397);
nand UO_1710 (O_1710,N_12825,N_14110);
xor UO_1711 (O_1711,N_12825,N_13457);
nand UO_1712 (O_1712,N_13574,N_12167);
nor UO_1713 (O_1713,N_14463,N_14138);
nor UO_1714 (O_1714,N_12893,N_13724);
nor UO_1715 (O_1715,N_14815,N_12922);
or UO_1716 (O_1716,N_13185,N_12629);
and UO_1717 (O_1717,N_12185,N_12312);
or UO_1718 (O_1718,N_12269,N_14855);
nor UO_1719 (O_1719,N_13839,N_13512);
nor UO_1720 (O_1720,N_14502,N_13287);
nor UO_1721 (O_1721,N_13567,N_14826);
nor UO_1722 (O_1722,N_13923,N_14205);
and UO_1723 (O_1723,N_14181,N_12334);
or UO_1724 (O_1724,N_13210,N_14182);
or UO_1725 (O_1725,N_13296,N_13750);
nor UO_1726 (O_1726,N_14773,N_13373);
and UO_1727 (O_1727,N_13233,N_14806);
nand UO_1728 (O_1728,N_12382,N_13964);
or UO_1729 (O_1729,N_13178,N_12361);
and UO_1730 (O_1730,N_14479,N_13537);
or UO_1731 (O_1731,N_12652,N_13672);
or UO_1732 (O_1732,N_13716,N_13247);
or UO_1733 (O_1733,N_12550,N_14431);
nor UO_1734 (O_1734,N_13164,N_13889);
nor UO_1735 (O_1735,N_14442,N_12937);
nand UO_1736 (O_1736,N_12016,N_13641);
or UO_1737 (O_1737,N_13065,N_14548);
nand UO_1738 (O_1738,N_13949,N_13807);
or UO_1739 (O_1739,N_13997,N_14656);
or UO_1740 (O_1740,N_14266,N_12489);
nand UO_1741 (O_1741,N_12548,N_14854);
or UO_1742 (O_1742,N_12821,N_13327);
and UO_1743 (O_1743,N_14701,N_12836);
nor UO_1744 (O_1744,N_14629,N_12484);
or UO_1745 (O_1745,N_13804,N_12416);
and UO_1746 (O_1746,N_14316,N_14714);
and UO_1747 (O_1747,N_12128,N_13347);
xor UO_1748 (O_1748,N_14244,N_14438);
or UO_1749 (O_1749,N_12172,N_13194);
nand UO_1750 (O_1750,N_12340,N_14395);
and UO_1751 (O_1751,N_13802,N_13983);
nor UO_1752 (O_1752,N_12990,N_12769);
nor UO_1753 (O_1753,N_14327,N_13560);
nor UO_1754 (O_1754,N_13321,N_12537);
and UO_1755 (O_1755,N_13209,N_12085);
nor UO_1756 (O_1756,N_13400,N_14257);
and UO_1757 (O_1757,N_14477,N_14175);
or UO_1758 (O_1758,N_14985,N_12459);
nor UO_1759 (O_1759,N_13368,N_13449);
or UO_1760 (O_1760,N_14234,N_13617);
nand UO_1761 (O_1761,N_13586,N_12200);
or UO_1762 (O_1762,N_12990,N_14672);
nor UO_1763 (O_1763,N_14965,N_12855);
and UO_1764 (O_1764,N_13866,N_13064);
or UO_1765 (O_1765,N_13609,N_14745);
or UO_1766 (O_1766,N_14537,N_13535);
and UO_1767 (O_1767,N_13782,N_12245);
nand UO_1768 (O_1768,N_13019,N_14536);
or UO_1769 (O_1769,N_13146,N_12277);
or UO_1770 (O_1770,N_14643,N_12067);
and UO_1771 (O_1771,N_13854,N_14575);
and UO_1772 (O_1772,N_13045,N_14999);
nand UO_1773 (O_1773,N_14526,N_12720);
or UO_1774 (O_1774,N_12639,N_13080);
and UO_1775 (O_1775,N_13749,N_13551);
and UO_1776 (O_1776,N_14553,N_12980);
and UO_1777 (O_1777,N_13055,N_12401);
and UO_1778 (O_1778,N_13980,N_14793);
nand UO_1779 (O_1779,N_12967,N_14578);
nand UO_1780 (O_1780,N_14286,N_14256);
and UO_1781 (O_1781,N_13621,N_13941);
and UO_1782 (O_1782,N_12175,N_12265);
nor UO_1783 (O_1783,N_14531,N_14409);
nand UO_1784 (O_1784,N_14080,N_13604);
or UO_1785 (O_1785,N_13068,N_13612);
and UO_1786 (O_1786,N_13861,N_14308);
and UO_1787 (O_1787,N_14998,N_12917);
and UO_1788 (O_1788,N_14869,N_13078);
nor UO_1789 (O_1789,N_14655,N_13117);
nand UO_1790 (O_1790,N_12071,N_12232);
and UO_1791 (O_1791,N_12195,N_12569);
nand UO_1792 (O_1792,N_13310,N_14269);
and UO_1793 (O_1793,N_12030,N_12253);
or UO_1794 (O_1794,N_14797,N_14806);
and UO_1795 (O_1795,N_14600,N_14428);
or UO_1796 (O_1796,N_13290,N_12892);
nand UO_1797 (O_1797,N_12373,N_12835);
or UO_1798 (O_1798,N_14070,N_13907);
nor UO_1799 (O_1799,N_13424,N_14330);
nand UO_1800 (O_1800,N_13778,N_13228);
nand UO_1801 (O_1801,N_12843,N_14933);
and UO_1802 (O_1802,N_12990,N_12294);
or UO_1803 (O_1803,N_14515,N_14045);
or UO_1804 (O_1804,N_13786,N_12417);
nor UO_1805 (O_1805,N_12510,N_13544);
and UO_1806 (O_1806,N_12280,N_13807);
nor UO_1807 (O_1807,N_13725,N_12466);
and UO_1808 (O_1808,N_12915,N_12149);
nor UO_1809 (O_1809,N_13893,N_12533);
or UO_1810 (O_1810,N_12814,N_13646);
nor UO_1811 (O_1811,N_14740,N_13060);
nor UO_1812 (O_1812,N_13700,N_12705);
nand UO_1813 (O_1813,N_12244,N_14340);
nand UO_1814 (O_1814,N_13637,N_12049);
nor UO_1815 (O_1815,N_13917,N_13604);
and UO_1816 (O_1816,N_12555,N_13522);
nor UO_1817 (O_1817,N_13438,N_13417);
and UO_1818 (O_1818,N_14166,N_14525);
or UO_1819 (O_1819,N_14103,N_13372);
nand UO_1820 (O_1820,N_13211,N_14218);
and UO_1821 (O_1821,N_12834,N_13776);
nand UO_1822 (O_1822,N_13909,N_12759);
and UO_1823 (O_1823,N_14094,N_14469);
nor UO_1824 (O_1824,N_13289,N_12960);
or UO_1825 (O_1825,N_12890,N_12350);
or UO_1826 (O_1826,N_13287,N_12045);
or UO_1827 (O_1827,N_13203,N_12126);
and UO_1828 (O_1828,N_12753,N_12760);
or UO_1829 (O_1829,N_14849,N_13415);
and UO_1830 (O_1830,N_14584,N_13147);
nand UO_1831 (O_1831,N_12572,N_12319);
or UO_1832 (O_1832,N_14970,N_12652);
nor UO_1833 (O_1833,N_14120,N_14520);
nand UO_1834 (O_1834,N_12184,N_14883);
nand UO_1835 (O_1835,N_12327,N_12024);
or UO_1836 (O_1836,N_14002,N_14312);
nand UO_1837 (O_1837,N_12280,N_14880);
or UO_1838 (O_1838,N_14666,N_14892);
or UO_1839 (O_1839,N_13128,N_13068);
nand UO_1840 (O_1840,N_14219,N_12627);
nor UO_1841 (O_1841,N_13083,N_14091);
nor UO_1842 (O_1842,N_12635,N_12664);
nor UO_1843 (O_1843,N_14443,N_12430);
nand UO_1844 (O_1844,N_12242,N_14676);
or UO_1845 (O_1845,N_13240,N_14648);
nor UO_1846 (O_1846,N_14792,N_13093);
and UO_1847 (O_1847,N_13690,N_13474);
and UO_1848 (O_1848,N_14902,N_12586);
or UO_1849 (O_1849,N_13043,N_13381);
or UO_1850 (O_1850,N_13933,N_14651);
and UO_1851 (O_1851,N_12012,N_13679);
nor UO_1852 (O_1852,N_12960,N_13809);
nor UO_1853 (O_1853,N_14008,N_14287);
and UO_1854 (O_1854,N_14840,N_12215);
and UO_1855 (O_1855,N_13589,N_12436);
or UO_1856 (O_1856,N_12098,N_14390);
xor UO_1857 (O_1857,N_14612,N_12164);
or UO_1858 (O_1858,N_14322,N_12990);
nor UO_1859 (O_1859,N_13462,N_12482);
nand UO_1860 (O_1860,N_14681,N_13007);
and UO_1861 (O_1861,N_13974,N_12071);
or UO_1862 (O_1862,N_13180,N_13938);
nor UO_1863 (O_1863,N_12200,N_13705);
and UO_1864 (O_1864,N_12136,N_12196);
nor UO_1865 (O_1865,N_12515,N_13376);
or UO_1866 (O_1866,N_14406,N_13155);
nand UO_1867 (O_1867,N_13597,N_12978);
and UO_1868 (O_1868,N_12964,N_12563);
nand UO_1869 (O_1869,N_14623,N_12575);
or UO_1870 (O_1870,N_12362,N_12342);
nand UO_1871 (O_1871,N_14495,N_14859);
and UO_1872 (O_1872,N_12000,N_14348);
nand UO_1873 (O_1873,N_14807,N_13897);
nand UO_1874 (O_1874,N_12687,N_14950);
or UO_1875 (O_1875,N_12431,N_12555);
nand UO_1876 (O_1876,N_13133,N_14230);
and UO_1877 (O_1877,N_13047,N_13751);
and UO_1878 (O_1878,N_14545,N_14165);
or UO_1879 (O_1879,N_14312,N_14678);
and UO_1880 (O_1880,N_14238,N_13175);
nand UO_1881 (O_1881,N_14450,N_12007);
or UO_1882 (O_1882,N_14752,N_14470);
and UO_1883 (O_1883,N_12278,N_12849);
and UO_1884 (O_1884,N_14478,N_13365);
or UO_1885 (O_1885,N_13478,N_13124);
nor UO_1886 (O_1886,N_12594,N_14042);
or UO_1887 (O_1887,N_13171,N_12523);
nor UO_1888 (O_1888,N_12895,N_13974);
nor UO_1889 (O_1889,N_13135,N_13176);
nor UO_1890 (O_1890,N_13321,N_13295);
and UO_1891 (O_1891,N_13602,N_14811);
or UO_1892 (O_1892,N_12044,N_14360);
or UO_1893 (O_1893,N_14180,N_14360);
or UO_1894 (O_1894,N_14164,N_14855);
and UO_1895 (O_1895,N_13132,N_12887);
and UO_1896 (O_1896,N_14477,N_14518);
nand UO_1897 (O_1897,N_13917,N_12290);
nor UO_1898 (O_1898,N_12972,N_14630);
or UO_1899 (O_1899,N_13060,N_13916);
or UO_1900 (O_1900,N_12111,N_14338);
nand UO_1901 (O_1901,N_13378,N_14870);
nor UO_1902 (O_1902,N_12890,N_14865);
or UO_1903 (O_1903,N_13359,N_14642);
nor UO_1904 (O_1904,N_13373,N_14276);
or UO_1905 (O_1905,N_12600,N_12289);
nor UO_1906 (O_1906,N_13449,N_13597);
and UO_1907 (O_1907,N_13043,N_13119);
nor UO_1908 (O_1908,N_13833,N_14674);
nand UO_1909 (O_1909,N_12720,N_13951);
or UO_1910 (O_1910,N_12063,N_13135);
nor UO_1911 (O_1911,N_13385,N_12907);
nand UO_1912 (O_1912,N_12730,N_14246);
nand UO_1913 (O_1913,N_12391,N_14929);
or UO_1914 (O_1914,N_14327,N_12881);
nand UO_1915 (O_1915,N_12171,N_12618);
or UO_1916 (O_1916,N_13247,N_12187);
nor UO_1917 (O_1917,N_12231,N_13432);
and UO_1918 (O_1918,N_13825,N_12135);
or UO_1919 (O_1919,N_13631,N_14648);
or UO_1920 (O_1920,N_13805,N_13498);
nor UO_1921 (O_1921,N_14240,N_12916);
and UO_1922 (O_1922,N_14575,N_13220);
or UO_1923 (O_1923,N_13279,N_12684);
nand UO_1924 (O_1924,N_12890,N_13806);
and UO_1925 (O_1925,N_12988,N_13993);
nand UO_1926 (O_1926,N_12816,N_13098);
or UO_1927 (O_1927,N_13668,N_12278);
or UO_1928 (O_1928,N_14505,N_14960);
nand UO_1929 (O_1929,N_13353,N_12854);
nor UO_1930 (O_1930,N_14319,N_14623);
nor UO_1931 (O_1931,N_13732,N_12582);
nor UO_1932 (O_1932,N_13275,N_14696);
nor UO_1933 (O_1933,N_14178,N_12811);
nand UO_1934 (O_1934,N_14374,N_12257);
nand UO_1935 (O_1935,N_13574,N_13233);
or UO_1936 (O_1936,N_12375,N_14965);
nand UO_1937 (O_1937,N_13757,N_12079);
or UO_1938 (O_1938,N_13393,N_12643);
and UO_1939 (O_1939,N_14780,N_12846);
and UO_1940 (O_1940,N_14940,N_14917);
nor UO_1941 (O_1941,N_14285,N_13728);
or UO_1942 (O_1942,N_13623,N_14809);
or UO_1943 (O_1943,N_13291,N_14787);
or UO_1944 (O_1944,N_12221,N_12682);
nand UO_1945 (O_1945,N_13201,N_13414);
and UO_1946 (O_1946,N_14043,N_12007);
nand UO_1947 (O_1947,N_14532,N_12141);
nor UO_1948 (O_1948,N_13326,N_12711);
nand UO_1949 (O_1949,N_12788,N_12322);
or UO_1950 (O_1950,N_13967,N_12564);
and UO_1951 (O_1951,N_12430,N_14890);
nand UO_1952 (O_1952,N_14806,N_14118);
or UO_1953 (O_1953,N_12621,N_14867);
or UO_1954 (O_1954,N_14044,N_12860);
or UO_1955 (O_1955,N_14804,N_13167);
nor UO_1956 (O_1956,N_13886,N_13166);
nand UO_1957 (O_1957,N_12642,N_14915);
or UO_1958 (O_1958,N_13753,N_14422);
nor UO_1959 (O_1959,N_14109,N_12169);
nand UO_1960 (O_1960,N_13758,N_13888);
or UO_1961 (O_1961,N_14702,N_14590);
or UO_1962 (O_1962,N_12070,N_12440);
or UO_1963 (O_1963,N_14111,N_14797);
or UO_1964 (O_1964,N_12461,N_12521);
nand UO_1965 (O_1965,N_14590,N_13462);
nand UO_1966 (O_1966,N_14746,N_14154);
and UO_1967 (O_1967,N_13269,N_12079);
nor UO_1968 (O_1968,N_14983,N_14436);
and UO_1969 (O_1969,N_14457,N_14742);
and UO_1970 (O_1970,N_13273,N_12023);
nand UO_1971 (O_1971,N_14659,N_14069);
and UO_1972 (O_1972,N_12167,N_14454);
nor UO_1973 (O_1973,N_13476,N_12525);
and UO_1974 (O_1974,N_12539,N_14786);
nor UO_1975 (O_1975,N_12319,N_12871);
or UO_1976 (O_1976,N_13112,N_12285);
and UO_1977 (O_1977,N_13602,N_12847);
or UO_1978 (O_1978,N_13609,N_14148);
nand UO_1979 (O_1979,N_12418,N_13618);
and UO_1980 (O_1980,N_12299,N_13795);
or UO_1981 (O_1981,N_12116,N_12076);
or UO_1982 (O_1982,N_12241,N_14348);
xor UO_1983 (O_1983,N_13271,N_14533);
or UO_1984 (O_1984,N_14248,N_12454);
and UO_1985 (O_1985,N_14171,N_13025);
nor UO_1986 (O_1986,N_13237,N_14119);
and UO_1987 (O_1987,N_13025,N_13457);
or UO_1988 (O_1988,N_13328,N_12097);
xnor UO_1989 (O_1989,N_14272,N_13971);
nand UO_1990 (O_1990,N_13997,N_14458);
and UO_1991 (O_1991,N_13661,N_13306);
and UO_1992 (O_1992,N_14131,N_13896);
and UO_1993 (O_1993,N_12263,N_12477);
and UO_1994 (O_1994,N_12595,N_13340);
nor UO_1995 (O_1995,N_14476,N_13914);
or UO_1996 (O_1996,N_12824,N_14180);
or UO_1997 (O_1997,N_12065,N_13333);
and UO_1998 (O_1998,N_14459,N_14375);
and UO_1999 (O_1999,N_12678,N_12987);
endmodule