module basic_500_3000_500_50_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_163,In_144);
nand U1 (N_1,In_211,In_134);
nand U2 (N_2,In_269,In_8);
and U3 (N_3,In_478,In_101);
nand U4 (N_4,In_242,In_26);
and U5 (N_5,In_128,In_328);
and U6 (N_6,In_32,In_202);
nand U7 (N_7,In_84,In_477);
and U8 (N_8,In_323,In_456);
or U9 (N_9,In_44,In_117);
nor U10 (N_10,In_196,In_153);
or U11 (N_11,In_77,In_332);
nor U12 (N_12,In_7,In_1);
nor U13 (N_13,In_124,In_222);
nor U14 (N_14,In_57,In_14);
xnor U15 (N_15,In_105,In_413);
or U16 (N_16,In_427,In_240);
and U17 (N_17,In_418,In_194);
and U18 (N_18,In_38,In_436);
nor U19 (N_19,In_291,In_268);
or U20 (N_20,In_86,In_238);
nand U21 (N_21,In_56,In_348);
or U22 (N_22,In_419,In_435);
or U23 (N_23,In_394,In_90);
or U24 (N_24,In_213,In_361);
or U25 (N_25,In_283,In_476);
nor U26 (N_26,In_472,In_145);
nand U27 (N_27,In_335,In_341);
and U28 (N_28,In_480,In_95);
and U29 (N_29,In_489,In_364);
nand U30 (N_30,In_343,In_299);
or U31 (N_31,In_251,In_140);
or U32 (N_32,In_19,In_239);
nor U33 (N_33,In_308,In_146);
or U34 (N_34,In_200,In_10);
nor U35 (N_35,In_162,In_305);
nand U36 (N_36,In_241,In_390);
and U37 (N_37,In_142,In_41);
nand U38 (N_38,In_298,In_199);
or U39 (N_39,In_284,In_416);
nor U40 (N_40,In_404,In_442);
and U41 (N_41,In_6,In_383);
xor U42 (N_42,In_319,In_382);
and U43 (N_43,In_420,In_141);
and U44 (N_44,In_387,In_18);
nor U45 (N_45,In_326,In_176);
and U46 (N_46,In_143,In_498);
nor U47 (N_47,In_206,In_374);
nor U48 (N_48,In_78,In_278);
or U49 (N_49,In_203,In_155);
nor U50 (N_50,In_345,In_169);
nor U51 (N_51,In_330,In_454);
and U52 (N_52,In_233,In_130);
nand U53 (N_53,In_360,In_290);
nand U54 (N_54,In_149,In_452);
and U55 (N_55,In_71,In_223);
xor U56 (N_56,In_131,In_17);
and U57 (N_57,In_386,In_102);
and U58 (N_58,In_373,In_349);
or U59 (N_59,In_257,In_98);
nor U60 (N_60,In_367,In_111);
or U61 (N_61,In_258,In_220);
nor U62 (N_62,In_85,N_47);
nor U63 (N_63,In_350,In_83);
and U64 (N_64,In_168,In_174);
xnor U65 (N_65,In_42,In_39);
nor U66 (N_66,In_475,In_380);
and U67 (N_67,In_219,In_62);
nor U68 (N_68,In_499,In_92);
nor U69 (N_69,N_38,In_253);
and U70 (N_70,In_487,In_372);
nor U71 (N_71,In_256,In_27);
and U72 (N_72,In_497,In_226);
nand U73 (N_73,In_368,In_282);
or U74 (N_74,In_422,In_186);
or U75 (N_75,In_228,In_33);
or U76 (N_76,In_66,In_362);
and U77 (N_77,N_42,In_285);
and U78 (N_78,In_188,In_354);
nor U79 (N_79,In_403,In_231);
nor U80 (N_80,In_371,In_112);
nand U81 (N_81,In_352,In_279);
and U82 (N_82,In_451,In_75);
or U83 (N_83,In_316,In_133);
xnor U84 (N_84,In_304,In_310);
xor U85 (N_85,In_224,In_467);
or U86 (N_86,In_407,In_457);
or U87 (N_87,In_209,In_230);
or U88 (N_88,In_204,N_14);
or U89 (N_89,In_333,In_346);
or U90 (N_90,In_395,In_152);
nor U91 (N_91,In_63,In_470);
nor U92 (N_92,In_82,In_287);
nand U93 (N_93,In_358,In_214);
or U94 (N_94,In_150,In_439);
xor U95 (N_95,In_347,In_400);
nor U96 (N_96,In_106,In_414);
xnor U97 (N_97,In_138,In_81);
and U98 (N_98,In_313,In_197);
nor U99 (N_99,In_23,In_3);
and U100 (N_100,In_312,In_119);
nor U101 (N_101,In_227,In_356);
nor U102 (N_102,In_170,In_154);
xnor U103 (N_103,In_329,N_28);
or U104 (N_104,In_402,In_384);
nand U105 (N_105,In_183,N_43);
and U106 (N_106,In_51,In_421);
nor U107 (N_107,In_307,In_125);
or U108 (N_108,In_173,In_243);
nor U109 (N_109,In_317,N_48);
nand U110 (N_110,In_482,In_496);
nand U111 (N_111,In_463,In_392);
and U112 (N_112,In_201,In_192);
xor U113 (N_113,In_359,In_261);
or U114 (N_114,In_453,In_431);
and U115 (N_115,In_184,N_59);
or U116 (N_116,N_49,In_22);
nor U117 (N_117,In_178,N_31);
and U118 (N_118,In_266,In_129);
nand U119 (N_119,N_23,In_55);
and U120 (N_120,In_486,In_275);
xor U121 (N_121,In_52,In_409);
nand U122 (N_122,In_303,In_492);
or U123 (N_123,In_68,In_47);
nand U124 (N_124,In_417,In_73);
and U125 (N_125,In_179,N_79);
and U126 (N_126,In_339,In_260);
or U127 (N_127,N_102,In_491);
nor U128 (N_128,In_462,In_110);
nor U129 (N_129,In_271,In_259);
and U130 (N_130,N_58,N_88);
or U131 (N_131,In_447,In_137);
and U132 (N_132,In_324,In_363);
nor U133 (N_133,In_208,In_195);
and U134 (N_134,In_429,In_446);
nand U135 (N_135,N_85,In_393);
nand U136 (N_136,In_236,In_99);
xor U137 (N_137,In_425,In_444);
nor U138 (N_138,In_296,In_272);
or U139 (N_139,In_250,N_29);
nor U140 (N_140,In_325,In_198);
nor U141 (N_141,In_189,In_495);
nor U142 (N_142,In_61,In_469);
nor U143 (N_143,In_247,N_117);
nand U144 (N_144,In_97,In_177);
nor U145 (N_145,N_108,In_79);
and U146 (N_146,In_280,In_29);
nand U147 (N_147,N_87,N_27);
nand U148 (N_148,N_97,In_397);
nor U149 (N_149,In_432,In_72);
nor U150 (N_150,In_88,In_232);
or U151 (N_151,N_61,In_434);
or U152 (N_152,In_375,In_334);
nor U153 (N_153,N_105,In_385);
xor U154 (N_154,In_428,In_118);
or U155 (N_155,In_460,N_69);
nand U156 (N_156,N_113,In_221);
or U157 (N_157,In_338,N_6);
and U158 (N_158,In_25,In_406);
nand U159 (N_159,N_32,N_98);
and U160 (N_160,In_139,N_109);
nor U161 (N_161,In_315,In_379);
nand U162 (N_162,In_262,In_210);
nand U163 (N_163,N_40,In_411);
nand U164 (N_164,In_54,In_289);
nor U165 (N_165,In_252,In_336);
or U166 (N_166,In_295,In_351);
nor U167 (N_167,In_474,N_63);
and U168 (N_168,N_17,In_158);
nor U169 (N_169,In_292,N_82);
or U170 (N_170,In_331,In_255);
and U171 (N_171,In_301,In_342);
or U172 (N_172,In_48,In_215);
and U173 (N_173,In_69,N_5);
xor U174 (N_174,N_75,N_104);
nand U175 (N_175,In_225,N_91);
and U176 (N_176,In_355,In_415);
and U177 (N_177,In_217,In_126);
nand U178 (N_178,N_101,N_116);
nor U179 (N_179,N_50,N_77);
or U180 (N_180,In_13,N_1);
or U181 (N_181,N_26,N_3);
or U182 (N_182,N_2,N_74);
and U183 (N_183,N_65,In_156);
and U184 (N_184,In_180,N_144);
nor U185 (N_185,In_193,In_235);
nor U186 (N_186,N_66,N_67);
and U187 (N_187,N_127,In_166);
nand U188 (N_188,N_141,In_31);
and U189 (N_189,N_4,In_264);
nand U190 (N_190,In_485,In_481);
xnor U191 (N_191,In_59,In_391);
or U192 (N_192,N_20,N_84);
nor U193 (N_193,N_94,In_24);
and U194 (N_194,In_80,In_74);
nand U195 (N_195,N_100,In_276);
xnor U196 (N_196,In_450,N_107);
or U197 (N_197,N_121,In_160);
and U198 (N_198,N_80,In_16);
nor U199 (N_199,N_164,In_167);
and U200 (N_200,N_78,N_150);
or U201 (N_201,In_396,In_340);
nand U202 (N_202,N_35,In_5);
xnor U203 (N_203,In_365,In_314);
nand U204 (N_204,In_322,N_155);
and U205 (N_205,N_138,In_286);
nand U206 (N_206,N_71,In_245);
nand U207 (N_207,N_11,In_104);
nor U208 (N_208,N_151,N_86);
or U209 (N_209,N_92,N_115);
and U210 (N_210,N_37,N_54);
and U211 (N_211,In_107,N_154);
xnor U212 (N_212,In_440,N_153);
nand U213 (N_213,N_122,In_114);
or U214 (N_214,In_490,In_108);
or U215 (N_215,In_164,In_50);
and U216 (N_216,In_132,N_30);
nor U217 (N_217,N_55,In_116);
nand U218 (N_218,N_93,N_19);
or U219 (N_219,N_139,N_143);
or U220 (N_220,In_465,In_357);
nor U221 (N_221,In_2,In_58);
nor U222 (N_222,In_76,N_64);
nand U223 (N_223,In_493,N_18);
nor U224 (N_224,N_0,In_40);
or U225 (N_225,In_165,N_132);
nor U226 (N_226,In_468,In_473);
or U227 (N_227,In_185,In_34);
nand U228 (N_228,N_118,In_494);
nor U229 (N_229,In_237,In_294);
nor U230 (N_230,In_378,In_127);
nand U231 (N_231,N_33,In_91);
nand U232 (N_232,In_94,N_22);
xnor U233 (N_233,In_65,In_229);
nand U234 (N_234,N_158,In_426);
nor U235 (N_235,In_376,N_177);
nor U236 (N_236,In_484,In_35);
nand U237 (N_237,N_56,In_263);
xor U238 (N_238,In_274,N_172);
nand U239 (N_239,In_265,In_399);
nand U240 (N_240,N_159,In_190);
and U241 (N_241,N_12,In_122);
or U242 (N_242,N_45,In_311);
or U243 (N_243,N_205,N_187);
and U244 (N_244,N_169,N_76);
xor U245 (N_245,N_137,N_156);
or U246 (N_246,In_423,N_60);
nor U247 (N_247,In_438,N_7);
and U248 (N_248,In_248,In_120);
nand U249 (N_249,N_175,N_185);
nor U250 (N_250,N_224,In_175);
xor U251 (N_251,In_254,N_214);
nand U252 (N_252,N_148,In_9);
nand U253 (N_253,N_57,N_53);
and U254 (N_254,N_41,In_205);
xor U255 (N_255,In_318,N_216);
xor U256 (N_256,In_320,N_128);
nand U257 (N_257,N_176,N_190);
nor U258 (N_258,N_119,In_369);
or U259 (N_259,N_210,In_366);
or U260 (N_260,N_174,N_220);
nand U261 (N_261,N_162,N_209);
and U262 (N_262,N_89,In_464);
nand U263 (N_263,In_21,In_103);
nand U264 (N_264,In_353,In_389);
nor U265 (N_265,N_9,In_60);
nand U266 (N_266,In_70,In_45);
or U267 (N_267,In_53,In_159);
and U268 (N_268,In_433,N_181);
or U269 (N_269,N_166,N_44);
xnor U270 (N_270,In_147,In_445);
nand U271 (N_271,In_448,In_161);
or U272 (N_272,In_89,N_160);
or U273 (N_273,N_163,N_183);
xnor U274 (N_274,In_151,In_37);
or U275 (N_275,N_200,N_24);
or U276 (N_276,In_302,In_187);
nand U277 (N_277,In_244,In_466);
or U278 (N_278,In_381,N_145);
or U279 (N_279,N_232,In_20);
and U280 (N_280,N_140,In_267);
or U281 (N_281,In_424,N_96);
nand U282 (N_282,N_72,N_152);
and U283 (N_283,In_4,In_293);
and U284 (N_284,In_93,In_0);
and U285 (N_285,N_189,N_62);
nor U286 (N_286,In_288,In_136);
nand U287 (N_287,In_471,N_147);
or U288 (N_288,N_197,N_182);
and U289 (N_289,In_12,In_408);
nor U290 (N_290,N_239,N_120);
and U291 (N_291,N_168,N_15);
or U292 (N_292,N_136,N_112);
nor U293 (N_293,In_458,N_81);
xor U294 (N_294,N_218,In_28);
nand U295 (N_295,N_178,In_483);
nor U296 (N_296,In_437,N_211);
nor U297 (N_297,In_157,N_180);
nand U298 (N_298,In_441,In_344);
nor U299 (N_299,In_171,In_370);
or U300 (N_300,N_293,N_213);
nand U301 (N_301,N_236,In_115);
and U302 (N_302,N_184,N_217);
and U303 (N_303,N_292,N_279);
and U304 (N_304,N_16,N_283);
xor U305 (N_305,N_258,N_262);
nand U306 (N_306,In_270,N_99);
nor U307 (N_307,In_123,N_242);
nor U308 (N_308,In_172,N_111);
or U309 (N_309,In_49,N_204);
nand U310 (N_310,N_249,N_257);
nor U311 (N_311,In_306,N_248);
nor U312 (N_312,In_181,N_126);
and U313 (N_313,In_30,N_68);
and U314 (N_314,N_266,N_260);
nand U315 (N_315,N_229,N_268);
nor U316 (N_316,In_461,N_246);
nor U317 (N_317,N_106,N_51);
nor U318 (N_318,In_67,N_165);
or U319 (N_319,In_488,N_256);
and U320 (N_320,In_309,N_295);
or U321 (N_321,In_459,N_10);
nand U322 (N_322,In_277,In_15);
or U323 (N_323,N_226,In_100);
or U324 (N_324,N_206,N_125);
nand U325 (N_325,N_238,N_286);
and U326 (N_326,N_179,N_25);
and U327 (N_327,N_240,In_216);
and U328 (N_328,N_288,N_244);
nor U329 (N_329,In_410,N_124);
nor U330 (N_330,N_52,N_272);
and U331 (N_331,N_161,In_249);
xor U332 (N_332,In_443,N_250);
nand U333 (N_333,N_253,N_36);
or U334 (N_334,N_247,N_241);
nand U335 (N_335,In_36,In_148);
and U336 (N_336,In_11,In_455);
or U337 (N_337,N_235,N_270);
and U338 (N_338,N_21,N_228);
and U339 (N_339,N_289,N_191);
nor U340 (N_340,N_269,In_449);
or U341 (N_341,N_114,N_223);
nand U342 (N_342,N_274,In_234);
and U343 (N_343,N_103,In_191);
and U344 (N_344,In_182,N_142);
and U345 (N_345,N_215,N_198);
and U346 (N_346,N_280,N_199);
nand U347 (N_347,N_230,N_73);
and U348 (N_348,N_90,In_297);
nand U349 (N_349,N_70,N_278);
and U350 (N_350,N_243,In_64);
nand U351 (N_351,N_261,N_188);
xor U352 (N_352,N_271,In_401);
or U353 (N_353,N_277,N_131);
and U354 (N_354,N_290,N_34);
nand U355 (N_355,N_297,N_255);
and U356 (N_356,N_173,N_234);
and U357 (N_357,In_337,In_96);
or U358 (N_358,N_251,In_135);
or U359 (N_359,N_273,N_193);
and U360 (N_360,N_133,N_170);
nand U361 (N_361,N_357,N_225);
nand U362 (N_362,N_324,N_304);
or U363 (N_363,N_291,N_344);
nor U364 (N_364,In_430,N_334);
and U365 (N_365,N_110,N_300);
nor U366 (N_366,N_319,N_8);
nand U367 (N_367,N_310,In_405);
nor U368 (N_368,In_273,In_87);
and U369 (N_369,N_284,N_346);
nand U370 (N_370,N_46,N_302);
and U371 (N_371,N_338,In_109);
or U372 (N_372,In_321,N_358);
nor U373 (N_373,N_233,N_345);
or U374 (N_374,N_339,N_39);
and U375 (N_375,N_314,N_352);
and U376 (N_376,N_303,N_331);
nand U377 (N_377,N_327,N_135);
nor U378 (N_378,N_212,N_315);
or U379 (N_379,N_326,In_300);
or U380 (N_380,N_196,N_353);
nand U381 (N_381,N_157,N_354);
and U382 (N_382,N_207,N_307);
nor U383 (N_383,N_254,N_313);
nor U384 (N_384,N_312,N_231);
and U385 (N_385,N_343,N_306);
nor U386 (N_386,N_309,N_146);
nor U387 (N_387,N_336,N_351);
nor U388 (N_388,N_237,N_192);
and U389 (N_389,N_203,N_13);
xor U390 (N_390,N_123,In_218);
nor U391 (N_391,In_327,N_328);
or U392 (N_392,N_275,N_347);
nand U393 (N_393,N_134,N_311);
xnor U394 (N_394,N_350,N_359);
nor U395 (N_395,In_46,N_333);
nor U396 (N_396,N_340,In_43);
xor U397 (N_397,N_149,N_130);
or U398 (N_398,N_227,N_342);
nor U399 (N_399,N_348,N_282);
nand U400 (N_400,N_355,N_83);
or U401 (N_401,N_171,N_323);
or U402 (N_402,N_95,N_267);
or U403 (N_403,N_335,N_330);
or U404 (N_404,N_298,N_186);
and U405 (N_405,N_305,N_222);
nand U406 (N_406,N_202,N_265);
or U407 (N_407,N_294,N_285);
nand U408 (N_408,In_398,N_318);
nand U409 (N_409,N_356,N_221);
or U410 (N_410,N_259,N_263);
and U411 (N_411,N_167,N_320);
nand U412 (N_412,In_246,N_208);
nor U413 (N_413,N_276,N_317);
xor U414 (N_414,N_325,N_252);
nor U415 (N_415,N_301,N_299);
or U416 (N_416,N_332,In_121);
and U417 (N_417,In_377,N_341);
nand U418 (N_418,N_349,N_219);
or U419 (N_419,N_264,N_194);
nor U420 (N_420,N_195,N_417);
nand U421 (N_421,N_374,N_407);
or U422 (N_422,N_296,N_404);
xor U423 (N_423,N_408,In_207);
nor U424 (N_424,N_367,N_129);
and U425 (N_425,N_402,N_380);
nor U426 (N_426,N_375,In_479);
or U427 (N_427,N_383,N_403);
nor U428 (N_428,N_370,N_384);
and U429 (N_429,N_413,N_391);
nor U430 (N_430,N_414,N_373);
xor U431 (N_431,N_410,N_376);
nand U432 (N_432,N_379,In_281);
and U433 (N_433,N_395,N_308);
nor U434 (N_434,N_401,N_419);
nand U435 (N_435,N_389,N_418);
nor U436 (N_436,N_337,N_378);
or U437 (N_437,N_281,N_386);
nand U438 (N_438,In_113,N_397);
and U439 (N_439,N_287,N_363);
nand U440 (N_440,N_394,N_369);
or U441 (N_441,N_392,N_415);
and U442 (N_442,N_322,N_371);
or U443 (N_443,N_366,N_390);
and U444 (N_444,N_361,N_412);
nand U445 (N_445,N_316,In_388);
and U446 (N_446,N_362,N_388);
nand U447 (N_447,N_399,N_321);
xor U448 (N_448,N_372,N_387);
and U449 (N_449,N_368,N_381);
nor U450 (N_450,N_411,N_201);
or U451 (N_451,N_416,N_398);
or U452 (N_452,N_406,N_245);
xor U453 (N_453,N_365,In_412);
nor U454 (N_454,N_405,N_382);
nor U455 (N_455,N_393,N_400);
nor U456 (N_456,In_212,N_329);
xor U457 (N_457,N_377,N_360);
nor U458 (N_458,N_396,N_385);
xor U459 (N_459,N_409,N_364);
and U460 (N_460,In_281,N_360);
or U461 (N_461,N_415,N_322);
nor U462 (N_462,In_479,In_212);
nand U463 (N_463,N_308,N_408);
nand U464 (N_464,N_396,In_207);
nor U465 (N_465,In_412,N_409);
nand U466 (N_466,N_394,N_376);
or U467 (N_467,N_418,N_412);
xor U468 (N_468,N_369,N_372);
nor U469 (N_469,N_362,N_398);
or U470 (N_470,N_374,N_409);
nand U471 (N_471,N_390,N_281);
and U472 (N_472,N_389,N_417);
or U473 (N_473,N_371,N_364);
nor U474 (N_474,N_380,N_413);
nand U475 (N_475,N_366,N_316);
xnor U476 (N_476,N_308,N_374);
nand U477 (N_477,N_414,N_337);
or U478 (N_478,In_207,N_373);
or U479 (N_479,N_281,N_373);
and U480 (N_480,N_470,N_472);
and U481 (N_481,N_444,N_478);
or U482 (N_482,N_425,N_438);
and U483 (N_483,N_429,N_466);
nor U484 (N_484,N_463,N_422);
nor U485 (N_485,N_423,N_439);
and U486 (N_486,N_433,N_424);
or U487 (N_487,N_426,N_437);
nor U488 (N_488,N_476,N_462);
nand U489 (N_489,N_454,N_446);
nor U490 (N_490,N_427,N_461);
or U491 (N_491,N_474,N_468);
and U492 (N_492,N_445,N_456);
or U493 (N_493,N_464,N_451);
and U494 (N_494,N_440,N_449);
nor U495 (N_495,N_471,N_479);
nor U496 (N_496,N_475,N_443);
nand U497 (N_497,N_460,N_448);
and U498 (N_498,N_421,N_436);
and U499 (N_499,N_435,N_469);
or U500 (N_500,N_431,N_473);
nand U501 (N_501,N_477,N_459);
or U502 (N_502,N_455,N_434);
nor U503 (N_503,N_450,N_441);
and U504 (N_504,N_467,N_453);
nor U505 (N_505,N_447,N_430);
or U506 (N_506,N_432,N_465);
and U507 (N_507,N_428,N_457);
xor U508 (N_508,N_452,N_442);
nand U509 (N_509,N_458,N_420);
and U510 (N_510,N_458,N_450);
nand U511 (N_511,N_479,N_439);
and U512 (N_512,N_428,N_461);
nand U513 (N_513,N_454,N_473);
nand U514 (N_514,N_458,N_466);
and U515 (N_515,N_436,N_428);
nor U516 (N_516,N_469,N_448);
nor U517 (N_517,N_476,N_429);
nand U518 (N_518,N_473,N_442);
and U519 (N_519,N_431,N_476);
nor U520 (N_520,N_441,N_467);
nand U521 (N_521,N_450,N_422);
or U522 (N_522,N_436,N_460);
xor U523 (N_523,N_479,N_422);
and U524 (N_524,N_478,N_479);
and U525 (N_525,N_437,N_428);
nand U526 (N_526,N_433,N_459);
nor U527 (N_527,N_454,N_435);
or U528 (N_528,N_446,N_458);
nor U529 (N_529,N_431,N_438);
or U530 (N_530,N_466,N_474);
nor U531 (N_531,N_471,N_437);
nor U532 (N_532,N_443,N_454);
or U533 (N_533,N_423,N_464);
and U534 (N_534,N_459,N_432);
nand U535 (N_535,N_440,N_463);
nor U536 (N_536,N_464,N_439);
nor U537 (N_537,N_475,N_462);
nor U538 (N_538,N_425,N_433);
nor U539 (N_539,N_442,N_474);
nand U540 (N_540,N_493,N_495);
or U541 (N_541,N_526,N_498);
nand U542 (N_542,N_531,N_488);
or U543 (N_543,N_483,N_529);
and U544 (N_544,N_520,N_521);
nand U545 (N_545,N_514,N_527);
nor U546 (N_546,N_510,N_504);
nor U547 (N_547,N_512,N_518);
or U548 (N_548,N_528,N_496);
nand U549 (N_549,N_513,N_494);
and U550 (N_550,N_534,N_524);
nand U551 (N_551,N_486,N_537);
nand U552 (N_552,N_523,N_482);
and U553 (N_553,N_502,N_505);
xor U554 (N_554,N_517,N_538);
nor U555 (N_555,N_491,N_532);
xnor U556 (N_556,N_503,N_480);
nand U557 (N_557,N_508,N_497);
nor U558 (N_558,N_533,N_511);
and U559 (N_559,N_507,N_499);
or U560 (N_560,N_509,N_492);
or U561 (N_561,N_485,N_484);
nor U562 (N_562,N_515,N_519);
and U563 (N_563,N_536,N_490);
nor U564 (N_564,N_525,N_522);
and U565 (N_565,N_481,N_500);
xnor U566 (N_566,N_487,N_501);
and U567 (N_567,N_539,N_489);
nand U568 (N_568,N_530,N_516);
nor U569 (N_569,N_535,N_506);
and U570 (N_570,N_535,N_510);
nand U571 (N_571,N_498,N_496);
or U572 (N_572,N_505,N_481);
and U573 (N_573,N_496,N_525);
nor U574 (N_574,N_512,N_497);
or U575 (N_575,N_532,N_527);
xnor U576 (N_576,N_529,N_512);
xor U577 (N_577,N_533,N_498);
or U578 (N_578,N_513,N_536);
xnor U579 (N_579,N_504,N_527);
and U580 (N_580,N_495,N_503);
nor U581 (N_581,N_514,N_499);
nor U582 (N_582,N_506,N_537);
nand U583 (N_583,N_490,N_480);
nand U584 (N_584,N_536,N_538);
nand U585 (N_585,N_510,N_532);
nor U586 (N_586,N_490,N_509);
or U587 (N_587,N_510,N_505);
and U588 (N_588,N_521,N_499);
nor U589 (N_589,N_495,N_538);
nor U590 (N_590,N_525,N_499);
nor U591 (N_591,N_515,N_530);
or U592 (N_592,N_480,N_517);
nor U593 (N_593,N_483,N_499);
nor U594 (N_594,N_493,N_489);
and U595 (N_595,N_515,N_496);
or U596 (N_596,N_528,N_530);
nand U597 (N_597,N_497,N_484);
and U598 (N_598,N_501,N_497);
nor U599 (N_599,N_483,N_480);
and U600 (N_600,N_566,N_571);
or U601 (N_601,N_581,N_540);
nand U602 (N_602,N_575,N_579);
xor U603 (N_603,N_546,N_592);
and U604 (N_604,N_565,N_599);
nor U605 (N_605,N_591,N_578);
nand U606 (N_606,N_589,N_577);
nor U607 (N_607,N_552,N_559);
and U608 (N_608,N_593,N_542);
nand U609 (N_609,N_588,N_586);
or U610 (N_610,N_580,N_585);
and U611 (N_611,N_556,N_550);
and U612 (N_612,N_595,N_553);
and U613 (N_613,N_554,N_545);
and U614 (N_614,N_567,N_557);
or U615 (N_615,N_597,N_549);
or U616 (N_616,N_570,N_555);
nor U617 (N_617,N_574,N_598);
and U618 (N_618,N_564,N_551);
and U619 (N_619,N_582,N_583);
xor U620 (N_620,N_587,N_576);
xor U621 (N_621,N_569,N_541);
and U622 (N_622,N_558,N_547);
nand U623 (N_623,N_584,N_543);
nor U624 (N_624,N_544,N_573);
and U625 (N_625,N_596,N_590);
nand U626 (N_626,N_594,N_563);
and U627 (N_627,N_561,N_568);
nor U628 (N_628,N_548,N_562);
and U629 (N_629,N_572,N_560);
nor U630 (N_630,N_588,N_569);
and U631 (N_631,N_554,N_591);
or U632 (N_632,N_572,N_592);
and U633 (N_633,N_551,N_585);
and U634 (N_634,N_581,N_587);
or U635 (N_635,N_565,N_580);
and U636 (N_636,N_594,N_557);
and U637 (N_637,N_560,N_575);
nand U638 (N_638,N_546,N_553);
and U639 (N_639,N_559,N_571);
or U640 (N_640,N_554,N_574);
or U641 (N_641,N_563,N_595);
nand U642 (N_642,N_540,N_554);
or U643 (N_643,N_542,N_596);
or U644 (N_644,N_568,N_545);
or U645 (N_645,N_546,N_545);
nand U646 (N_646,N_592,N_573);
xnor U647 (N_647,N_549,N_558);
and U648 (N_648,N_591,N_569);
nand U649 (N_649,N_577,N_596);
nor U650 (N_650,N_544,N_577);
and U651 (N_651,N_583,N_590);
or U652 (N_652,N_592,N_542);
and U653 (N_653,N_568,N_588);
xor U654 (N_654,N_581,N_562);
nand U655 (N_655,N_563,N_574);
xnor U656 (N_656,N_560,N_568);
xnor U657 (N_657,N_569,N_566);
and U658 (N_658,N_547,N_582);
xnor U659 (N_659,N_559,N_596);
or U660 (N_660,N_633,N_628);
nand U661 (N_661,N_617,N_645);
nand U662 (N_662,N_631,N_606);
or U663 (N_663,N_651,N_620);
and U664 (N_664,N_619,N_637);
or U665 (N_665,N_648,N_604);
and U666 (N_666,N_658,N_639);
and U667 (N_667,N_647,N_638);
nor U668 (N_668,N_600,N_622);
and U669 (N_669,N_607,N_643);
nand U670 (N_670,N_603,N_653);
and U671 (N_671,N_608,N_624);
nor U672 (N_672,N_618,N_646);
nand U673 (N_673,N_642,N_635);
nor U674 (N_674,N_605,N_656);
and U675 (N_675,N_652,N_632);
or U676 (N_676,N_625,N_615);
and U677 (N_677,N_629,N_601);
or U678 (N_678,N_611,N_609);
or U679 (N_679,N_614,N_644);
nor U680 (N_680,N_640,N_657);
nor U681 (N_681,N_623,N_654);
and U682 (N_682,N_659,N_616);
nor U683 (N_683,N_630,N_621);
or U684 (N_684,N_627,N_634);
xor U685 (N_685,N_613,N_602);
nand U686 (N_686,N_626,N_655);
nand U687 (N_687,N_612,N_650);
and U688 (N_688,N_610,N_649);
or U689 (N_689,N_641,N_636);
and U690 (N_690,N_644,N_647);
and U691 (N_691,N_649,N_601);
and U692 (N_692,N_609,N_642);
nand U693 (N_693,N_620,N_626);
nand U694 (N_694,N_655,N_639);
and U695 (N_695,N_654,N_651);
or U696 (N_696,N_659,N_635);
or U697 (N_697,N_601,N_658);
or U698 (N_698,N_607,N_617);
nor U699 (N_699,N_639,N_603);
nand U700 (N_700,N_652,N_610);
and U701 (N_701,N_609,N_631);
or U702 (N_702,N_658,N_644);
nand U703 (N_703,N_645,N_629);
and U704 (N_704,N_612,N_639);
xor U705 (N_705,N_648,N_654);
nand U706 (N_706,N_600,N_656);
and U707 (N_707,N_604,N_642);
or U708 (N_708,N_658,N_625);
and U709 (N_709,N_615,N_635);
or U710 (N_710,N_600,N_605);
nand U711 (N_711,N_601,N_648);
or U712 (N_712,N_648,N_621);
nor U713 (N_713,N_621,N_623);
or U714 (N_714,N_603,N_656);
xnor U715 (N_715,N_657,N_617);
and U716 (N_716,N_647,N_616);
xnor U717 (N_717,N_602,N_612);
or U718 (N_718,N_615,N_630);
nand U719 (N_719,N_610,N_650);
or U720 (N_720,N_715,N_710);
nand U721 (N_721,N_670,N_668);
and U722 (N_722,N_662,N_675);
and U723 (N_723,N_689,N_687);
xnor U724 (N_724,N_700,N_661);
nor U725 (N_725,N_717,N_719);
xnor U726 (N_726,N_669,N_708);
and U727 (N_727,N_678,N_693);
xor U728 (N_728,N_716,N_694);
and U729 (N_729,N_697,N_671);
nand U730 (N_730,N_680,N_695);
nand U731 (N_731,N_696,N_709);
xnor U732 (N_732,N_673,N_685);
nor U733 (N_733,N_683,N_704);
or U734 (N_734,N_672,N_698);
and U735 (N_735,N_677,N_682);
nand U736 (N_736,N_713,N_674);
or U737 (N_737,N_664,N_665);
and U738 (N_738,N_688,N_711);
or U739 (N_739,N_681,N_692);
xnor U740 (N_740,N_701,N_691);
xnor U741 (N_741,N_686,N_690);
nand U742 (N_742,N_660,N_714);
nor U743 (N_743,N_718,N_699);
or U744 (N_744,N_667,N_707);
and U745 (N_745,N_666,N_702);
or U746 (N_746,N_684,N_706);
xor U747 (N_747,N_703,N_712);
and U748 (N_748,N_679,N_705);
nor U749 (N_749,N_663,N_676);
and U750 (N_750,N_679,N_712);
and U751 (N_751,N_667,N_662);
nand U752 (N_752,N_687,N_703);
and U753 (N_753,N_698,N_663);
or U754 (N_754,N_705,N_712);
nor U755 (N_755,N_716,N_677);
nor U756 (N_756,N_661,N_662);
and U757 (N_757,N_662,N_665);
xnor U758 (N_758,N_708,N_675);
and U759 (N_759,N_675,N_707);
and U760 (N_760,N_685,N_711);
or U761 (N_761,N_680,N_706);
or U762 (N_762,N_666,N_713);
or U763 (N_763,N_711,N_670);
and U764 (N_764,N_668,N_719);
nand U765 (N_765,N_673,N_687);
or U766 (N_766,N_688,N_717);
nor U767 (N_767,N_712,N_664);
nand U768 (N_768,N_691,N_660);
nor U769 (N_769,N_705,N_717);
or U770 (N_770,N_696,N_703);
or U771 (N_771,N_708,N_681);
and U772 (N_772,N_690,N_715);
or U773 (N_773,N_715,N_719);
xor U774 (N_774,N_704,N_705);
xor U775 (N_775,N_707,N_689);
nand U776 (N_776,N_682,N_698);
or U777 (N_777,N_704,N_692);
or U778 (N_778,N_702,N_670);
nand U779 (N_779,N_693,N_683);
xor U780 (N_780,N_764,N_761);
or U781 (N_781,N_738,N_753);
or U782 (N_782,N_735,N_778);
nor U783 (N_783,N_746,N_745);
and U784 (N_784,N_768,N_772);
nand U785 (N_785,N_739,N_736);
or U786 (N_786,N_759,N_725);
and U787 (N_787,N_773,N_747);
and U788 (N_788,N_730,N_765);
and U789 (N_789,N_771,N_727);
and U790 (N_790,N_779,N_750);
or U791 (N_791,N_751,N_720);
or U792 (N_792,N_726,N_763);
nor U793 (N_793,N_743,N_742);
or U794 (N_794,N_766,N_758);
nand U795 (N_795,N_754,N_769);
or U796 (N_796,N_741,N_752);
and U797 (N_797,N_757,N_733);
or U798 (N_798,N_731,N_777);
nand U799 (N_799,N_755,N_775);
nand U800 (N_800,N_722,N_723);
nor U801 (N_801,N_776,N_721);
and U802 (N_802,N_767,N_734);
nor U803 (N_803,N_740,N_732);
or U804 (N_804,N_760,N_756);
xnor U805 (N_805,N_729,N_728);
or U806 (N_806,N_744,N_737);
and U807 (N_807,N_770,N_748);
nand U808 (N_808,N_762,N_724);
nand U809 (N_809,N_749,N_774);
xnor U810 (N_810,N_742,N_751);
and U811 (N_811,N_766,N_767);
or U812 (N_812,N_740,N_733);
and U813 (N_813,N_766,N_733);
nand U814 (N_814,N_755,N_779);
nand U815 (N_815,N_750,N_774);
xor U816 (N_816,N_759,N_776);
nand U817 (N_817,N_751,N_775);
nand U818 (N_818,N_736,N_749);
nor U819 (N_819,N_744,N_766);
or U820 (N_820,N_770,N_766);
xor U821 (N_821,N_767,N_723);
and U822 (N_822,N_770,N_776);
nand U823 (N_823,N_768,N_766);
xor U824 (N_824,N_776,N_774);
nand U825 (N_825,N_771,N_726);
nand U826 (N_826,N_731,N_727);
or U827 (N_827,N_741,N_742);
xnor U828 (N_828,N_776,N_743);
or U829 (N_829,N_730,N_769);
or U830 (N_830,N_776,N_763);
or U831 (N_831,N_743,N_768);
nor U832 (N_832,N_733,N_738);
xor U833 (N_833,N_758,N_741);
and U834 (N_834,N_752,N_726);
nor U835 (N_835,N_760,N_735);
and U836 (N_836,N_768,N_725);
nor U837 (N_837,N_743,N_762);
or U838 (N_838,N_742,N_779);
nand U839 (N_839,N_724,N_776);
and U840 (N_840,N_804,N_814);
nand U841 (N_841,N_787,N_803);
nor U842 (N_842,N_833,N_789);
nand U843 (N_843,N_824,N_794);
or U844 (N_844,N_829,N_802);
nand U845 (N_845,N_792,N_795);
or U846 (N_846,N_810,N_821);
nand U847 (N_847,N_785,N_817);
and U848 (N_848,N_826,N_819);
or U849 (N_849,N_784,N_832);
nor U850 (N_850,N_812,N_791);
nand U851 (N_851,N_835,N_823);
nor U852 (N_852,N_797,N_822);
nor U853 (N_853,N_834,N_790);
and U854 (N_854,N_808,N_793);
nor U855 (N_855,N_838,N_830);
and U856 (N_856,N_813,N_831);
nand U857 (N_857,N_806,N_825);
nor U858 (N_858,N_801,N_796);
xor U859 (N_859,N_783,N_839);
nand U860 (N_860,N_781,N_828);
nor U861 (N_861,N_837,N_788);
nand U862 (N_862,N_799,N_780);
nor U863 (N_863,N_782,N_827);
nand U864 (N_864,N_836,N_816);
and U865 (N_865,N_818,N_786);
nand U866 (N_866,N_811,N_820);
xnor U867 (N_867,N_798,N_807);
and U868 (N_868,N_800,N_805);
or U869 (N_869,N_809,N_815);
and U870 (N_870,N_824,N_833);
nand U871 (N_871,N_794,N_814);
or U872 (N_872,N_808,N_817);
nor U873 (N_873,N_781,N_837);
nand U874 (N_874,N_829,N_812);
nor U875 (N_875,N_814,N_792);
nand U876 (N_876,N_821,N_809);
nor U877 (N_877,N_805,N_798);
xor U878 (N_878,N_792,N_838);
nand U879 (N_879,N_831,N_838);
nand U880 (N_880,N_837,N_814);
xnor U881 (N_881,N_825,N_791);
nand U882 (N_882,N_818,N_813);
and U883 (N_883,N_805,N_808);
or U884 (N_884,N_793,N_780);
or U885 (N_885,N_822,N_816);
and U886 (N_886,N_813,N_819);
and U887 (N_887,N_815,N_791);
or U888 (N_888,N_838,N_794);
xnor U889 (N_889,N_802,N_831);
or U890 (N_890,N_790,N_828);
and U891 (N_891,N_791,N_828);
nand U892 (N_892,N_792,N_823);
nand U893 (N_893,N_830,N_822);
or U894 (N_894,N_822,N_835);
or U895 (N_895,N_822,N_811);
nor U896 (N_896,N_815,N_803);
nor U897 (N_897,N_797,N_807);
and U898 (N_898,N_802,N_788);
or U899 (N_899,N_802,N_821);
nand U900 (N_900,N_841,N_889);
or U901 (N_901,N_869,N_866);
nor U902 (N_902,N_857,N_886);
nor U903 (N_903,N_854,N_859);
nand U904 (N_904,N_868,N_893);
or U905 (N_905,N_850,N_875);
nor U906 (N_906,N_882,N_880);
xnor U907 (N_907,N_876,N_845);
nor U908 (N_908,N_883,N_887);
nand U909 (N_909,N_852,N_871);
nand U910 (N_910,N_844,N_878);
xor U911 (N_911,N_896,N_860);
nand U912 (N_912,N_867,N_899);
and U913 (N_913,N_897,N_856);
or U914 (N_914,N_894,N_851);
nor U915 (N_915,N_873,N_858);
nor U916 (N_916,N_884,N_879);
xnor U917 (N_917,N_853,N_898);
or U918 (N_918,N_872,N_849);
nand U919 (N_919,N_890,N_888);
nand U920 (N_920,N_862,N_870);
nand U921 (N_921,N_874,N_861);
or U922 (N_922,N_855,N_847);
nor U923 (N_923,N_865,N_877);
and U924 (N_924,N_846,N_848);
xor U925 (N_925,N_842,N_843);
nor U926 (N_926,N_881,N_885);
or U927 (N_927,N_840,N_892);
nor U928 (N_928,N_895,N_864);
nor U929 (N_929,N_863,N_891);
and U930 (N_930,N_863,N_879);
or U931 (N_931,N_891,N_852);
nand U932 (N_932,N_850,N_881);
nand U933 (N_933,N_855,N_846);
nand U934 (N_934,N_853,N_879);
nand U935 (N_935,N_868,N_843);
and U936 (N_936,N_892,N_878);
nor U937 (N_937,N_881,N_841);
nor U938 (N_938,N_872,N_843);
xnor U939 (N_939,N_870,N_885);
xnor U940 (N_940,N_848,N_867);
or U941 (N_941,N_882,N_892);
nor U942 (N_942,N_864,N_861);
nor U943 (N_943,N_883,N_863);
nor U944 (N_944,N_872,N_885);
nor U945 (N_945,N_865,N_895);
nor U946 (N_946,N_846,N_898);
xnor U947 (N_947,N_840,N_869);
and U948 (N_948,N_876,N_879);
nand U949 (N_949,N_890,N_851);
or U950 (N_950,N_845,N_878);
or U951 (N_951,N_875,N_841);
xor U952 (N_952,N_864,N_859);
and U953 (N_953,N_850,N_852);
or U954 (N_954,N_872,N_857);
or U955 (N_955,N_844,N_874);
or U956 (N_956,N_894,N_896);
or U957 (N_957,N_885,N_877);
nor U958 (N_958,N_862,N_851);
or U959 (N_959,N_867,N_847);
nor U960 (N_960,N_923,N_936);
and U961 (N_961,N_946,N_951);
nor U962 (N_962,N_925,N_903);
or U963 (N_963,N_931,N_954);
nor U964 (N_964,N_929,N_959);
nor U965 (N_965,N_932,N_926);
and U966 (N_966,N_913,N_952);
and U967 (N_967,N_921,N_953);
nor U968 (N_968,N_956,N_918);
nand U969 (N_969,N_912,N_927);
and U970 (N_970,N_920,N_906);
and U971 (N_971,N_904,N_922);
nor U972 (N_972,N_949,N_928);
nand U973 (N_973,N_910,N_930);
nand U974 (N_974,N_942,N_940);
or U975 (N_975,N_924,N_943);
nand U976 (N_976,N_937,N_945);
xnor U977 (N_977,N_911,N_957);
nand U978 (N_978,N_948,N_938);
and U979 (N_979,N_947,N_958);
xor U980 (N_980,N_914,N_909);
nand U981 (N_981,N_916,N_917);
nand U982 (N_982,N_939,N_919);
nand U983 (N_983,N_908,N_934);
and U984 (N_984,N_915,N_933);
nand U985 (N_985,N_900,N_905);
nor U986 (N_986,N_902,N_901);
or U987 (N_987,N_944,N_935);
nand U988 (N_988,N_950,N_955);
nor U989 (N_989,N_907,N_941);
and U990 (N_990,N_908,N_902);
or U991 (N_991,N_913,N_930);
or U992 (N_992,N_953,N_959);
nor U993 (N_993,N_953,N_908);
or U994 (N_994,N_950,N_902);
or U995 (N_995,N_914,N_955);
xnor U996 (N_996,N_951,N_908);
nor U997 (N_997,N_944,N_955);
xor U998 (N_998,N_919,N_922);
nand U999 (N_999,N_931,N_919);
nand U1000 (N_1000,N_942,N_958);
nor U1001 (N_1001,N_915,N_954);
nor U1002 (N_1002,N_934,N_902);
or U1003 (N_1003,N_923,N_940);
and U1004 (N_1004,N_959,N_933);
or U1005 (N_1005,N_945,N_958);
and U1006 (N_1006,N_953,N_944);
and U1007 (N_1007,N_926,N_928);
nor U1008 (N_1008,N_903,N_906);
or U1009 (N_1009,N_921,N_917);
nand U1010 (N_1010,N_952,N_919);
nor U1011 (N_1011,N_950,N_942);
nor U1012 (N_1012,N_941,N_959);
and U1013 (N_1013,N_935,N_934);
or U1014 (N_1014,N_959,N_956);
or U1015 (N_1015,N_937,N_946);
and U1016 (N_1016,N_937,N_943);
nor U1017 (N_1017,N_924,N_957);
or U1018 (N_1018,N_908,N_955);
or U1019 (N_1019,N_924,N_903);
nand U1020 (N_1020,N_966,N_1000);
nand U1021 (N_1021,N_1006,N_992);
or U1022 (N_1022,N_999,N_1013);
nor U1023 (N_1023,N_970,N_1009);
or U1024 (N_1024,N_998,N_967);
or U1025 (N_1025,N_974,N_1004);
or U1026 (N_1026,N_987,N_989);
nor U1027 (N_1027,N_982,N_986);
or U1028 (N_1028,N_962,N_961);
and U1029 (N_1029,N_971,N_969);
nor U1030 (N_1030,N_1016,N_1018);
nor U1031 (N_1031,N_1012,N_996);
nor U1032 (N_1032,N_1014,N_1008);
nor U1033 (N_1033,N_1011,N_980);
or U1034 (N_1034,N_984,N_988);
nand U1035 (N_1035,N_977,N_1003);
and U1036 (N_1036,N_975,N_968);
and U1037 (N_1037,N_1005,N_979);
nor U1038 (N_1038,N_1017,N_990);
or U1039 (N_1039,N_994,N_1010);
nor U1040 (N_1040,N_1007,N_1002);
nand U1041 (N_1041,N_963,N_993);
nand U1042 (N_1042,N_995,N_997);
and U1043 (N_1043,N_985,N_964);
xnor U1044 (N_1044,N_991,N_978);
nand U1045 (N_1045,N_983,N_965);
or U1046 (N_1046,N_1001,N_1015);
and U1047 (N_1047,N_976,N_973);
and U1048 (N_1048,N_1019,N_972);
or U1049 (N_1049,N_960,N_981);
nand U1050 (N_1050,N_960,N_987);
nor U1051 (N_1051,N_966,N_987);
or U1052 (N_1052,N_1010,N_987);
nand U1053 (N_1053,N_1007,N_1013);
xnor U1054 (N_1054,N_960,N_980);
nand U1055 (N_1055,N_1006,N_1004);
nand U1056 (N_1056,N_999,N_968);
nor U1057 (N_1057,N_1002,N_987);
and U1058 (N_1058,N_987,N_986);
nand U1059 (N_1059,N_1016,N_971);
or U1060 (N_1060,N_973,N_979);
nor U1061 (N_1061,N_1011,N_978);
nor U1062 (N_1062,N_969,N_994);
nor U1063 (N_1063,N_966,N_986);
or U1064 (N_1064,N_974,N_1019);
nand U1065 (N_1065,N_1019,N_1002);
and U1066 (N_1066,N_983,N_995);
xnor U1067 (N_1067,N_974,N_976);
nand U1068 (N_1068,N_1004,N_1008);
or U1069 (N_1069,N_1013,N_992);
xor U1070 (N_1070,N_1013,N_985);
nor U1071 (N_1071,N_994,N_980);
nand U1072 (N_1072,N_1019,N_988);
or U1073 (N_1073,N_970,N_969);
or U1074 (N_1074,N_988,N_1002);
nand U1075 (N_1075,N_965,N_975);
or U1076 (N_1076,N_977,N_1001);
and U1077 (N_1077,N_1007,N_960);
and U1078 (N_1078,N_1007,N_963);
nor U1079 (N_1079,N_988,N_1003);
and U1080 (N_1080,N_1041,N_1047);
xor U1081 (N_1081,N_1075,N_1063);
or U1082 (N_1082,N_1072,N_1064);
nand U1083 (N_1083,N_1051,N_1028);
nand U1084 (N_1084,N_1050,N_1026);
nor U1085 (N_1085,N_1037,N_1024);
nor U1086 (N_1086,N_1071,N_1045);
nand U1087 (N_1087,N_1049,N_1065);
xor U1088 (N_1088,N_1079,N_1061);
or U1089 (N_1089,N_1032,N_1067);
or U1090 (N_1090,N_1076,N_1056);
or U1091 (N_1091,N_1020,N_1031);
and U1092 (N_1092,N_1044,N_1035);
and U1093 (N_1093,N_1030,N_1069);
and U1094 (N_1094,N_1074,N_1027);
and U1095 (N_1095,N_1034,N_1052);
or U1096 (N_1096,N_1033,N_1021);
or U1097 (N_1097,N_1059,N_1040);
nor U1098 (N_1098,N_1048,N_1078);
xor U1099 (N_1099,N_1058,N_1068);
nor U1100 (N_1100,N_1070,N_1038);
nand U1101 (N_1101,N_1066,N_1029);
or U1102 (N_1102,N_1060,N_1043);
xor U1103 (N_1103,N_1073,N_1042);
nor U1104 (N_1104,N_1054,N_1055);
nor U1105 (N_1105,N_1039,N_1077);
or U1106 (N_1106,N_1023,N_1036);
nand U1107 (N_1107,N_1053,N_1057);
and U1108 (N_1108,N_1062,N_1022);
or U1109 (N_1109,N_1025,N_1046);
or U1110 (N_1110,N_1034,N_1056);
nor U1111 (N_1111,N_1029,N_1027);
xor U1112 (N_1112,N_1066,N_1049);
xnor U1113 (N_1113,N_1038,N_1060);
and U1114 (N_1114,N_1036,N_1040);
nand U1115 (N_1115,N_1027,N_1063);
nor U1116 (N_1116,N_1070,N_1034);
nor U1117 (N_1117,N_1067,N_1063);
nand U1118 (N_1118,N_1027,N_1052);
or U1119 (N_1119,N_1078,N_1044);
and U1120 (N_1120,N_1069,N_1036);
or U1121 (N_1121,N_1021,N_1072);
or U1122 (N_1122,N_1034,N_1043);
and U1123 (N_1123,N_1043,N_1054);
nor U1124 (N_1124,N_1068,N_1061);
nor U1125 (N_1125,N_1074,N_1055);
and U1126 (N_1126,N_1065,N_1048);
nor U1127 (N_1127,N_1057,N_1027);
xnor U1128 (N_1128,N_1076,N_1023);
nand U1129 (N_1129,N_1023,N_1033);
nand U1130 (N_1130,N_1041,N_1045);
xnor U1131 (N_1131,N_1060,N_1036);
nand U1132 (N_1132,N_1035,N_1022);
nand U1133 (N_1133,N_1037,N_1047);
nor U1134 (N_1134,N_1057,N_1046);
nor U1135 (N_1135,N_1035,N_1036);
or U1136 (N_1136,N_1076,N_1062);
and U1137 (N_1137,N_1075,N_1024);
nand U1138 (N_1138,N_1047,N_1077);
nor U1139 (N_1139,N_1039,N_1040);
nor U1140 (N_1140,N_1119,N_1082);
nor U1141 (N_1141,N_1135,N_1106);
xnor U1142 (N_1142,N_1136,N_1080);
xor U1143 (N_1143,N_1120,N_1132);
xor U1144 (N_1144,N_1095,N_1110);
or U1145 (N_1145,N_1090,N_1091);
or U1146 (N_1146,N_1118,N_1098);
and U1147 (N_1147,N_1117,N_1125);
nor U1148 (N_1148,N_1139,N_1130);
or U1149 (N_1149,N_1123,N_1114);
and U1150 (N_1150,N_1122,N_1133);
nand U1151 (N_1151,N_1083,N_1087);
nor U1152 (N_1152,N_1116,N_1081);
xnor U1153 (N_1153,N_1129,N_1124);
and U1154 (N_1154,N_1097,N_1134);
nor U1155 (N_1155,N_1102,N_1109);
nand U1156 (N_1156,N_1131,N_1085);
and U1157 (N_1157,N_1100,N_1089);
nor U1158 (N_1158,N_1101,N_1137);
and U1159 (N_1159,N_1108,N_1121);
nand U1160 (N_1160,N_1113,N_1104);
and U1161 (N_1161,N_1084,N_1094);
xor U1162 (N_1162,N_1138,N_1115);
xnor U1163 (N_1163,N_1127,N_1088);
xor U1164 (N_1164,N_1099,N_1111);
and U1165 (N_1165,N_1107,N_1105);
or U1166 (N_1166,N_1112,N_1128);
nand U1167 (N_1167,N_1092,N_1096);
nand U1168 (N_1168,N_1093,N_1103);
or U1169 (N_1169,N_1086,N_1126);
nand U1170 (N_1170,N_1123,N_1118);
nor U1171 (N_1171,N_1115,N_1135);
nand U1172 (N_1172,N_1133,N_1124);
and U1173 (N_1173,N_1092,N_1083);
nand U1174 (N_1174,N_1117,N_1127);
or U1175 (N_1175,N_1097,N_1112);
nand U1176 (N_1176,N_1088,N_1123);
nand U1177 (N_1177,N_1092,N_1093);
nand U1178 (N_1178,N_1104,N_1121);
nor U1179 (N_1179,N_1131,N_1134);
and U1180 (N_1180,N_1109,N_1092);
and U1181 (N_1181,N_1093,N_1082);
nand U1182 (N_1182,N_1136,N_1139);
nor U1183 (N_1183,N_1136,N_1086);
xnor U1184 (N_1184,N_1128,N_1123);
or U1185 (N_1185,N_1093,N_1124);
or U1186 (N_1186,N_1113,N_1099);
and U1187 (N_1187,N_1118,N_1086);
or U1188 (N_1188,N_1127,N_1085);
nor U1189 (N_1189,N_1081,N_1125);
nand U1190 (N_1190,N_1088,N_1095);
and U1191 (N_1191,N_1112,N_1127);
or U1192 (N_1192,N_1090,N_1100);
or U1193 (N_1193,N_1095,N_1126);
nand U1194 (N_1194,N_1101,N_1112);
nand U1195 (N_1195,N_1124,N_1105);
nand U1196 (N_1196,N_1096,N_1118);
nand U1197 (N_1197,N_1132,N_1102);
nor U1198 (N_1198,N_1113,N_1137);
nor U1199 (N_1199,N_1110,N_1104);
nor U1200 (N_1200,N_1168,N_1182);
and U1201 (N_1201,N_1175,N_1158);
or U1202 (N_1202,N_1177,N_1164);
nor U1203 (N_1203,N_1155,N_1150);
nand U1204 (N_1204,N_1156,N_1157);
nand U1205 (N_1205,N_1189,N_1179);
nor U1206 (N_1206,N_1161,N_1183);
and U1207 (N_1207,N_1174,N_1140);
nor U1208 (N_1208,N_1197,N_1187);
or U1209 (N_1209,N_1198,N_1159);
xnor U1210 (N_1210,N_1166,N_1148);
and U1211 (N_1211,N_1192,N_1143);
or U1212 (N_1212,N_1176,N_1195);
nor U1213 (N_1213,N_1173,N_1191);
nor U1214 (N_1214,N_1170,N_1149);
nor U1215 (N_1215,N_1146,N_1162);
or U1216 (N_1216,N_1178,N_1145);
nand U1217 (N_1217,N_1142,N_1172);
nor U1218 (N_1218,N_1180,N_1190);
nand U1219 (N_1219,N_1194,N_1199);
or U1220 (N_1220,N_1154,N_1184);
or U1221 (N_1221,N_1171,N_1196);
nor U1222 (N_1222,N_1188,N_1160);
nand U1223 (N_1223,N_1151,N_1181);
nand U1224 (N_1224,N_1165,N_1185);
or U1225 (N_1225,N_1167,N_1144);
and U1226 (N_1226,N_1141,N_1147);
or U1227 (N_1227,N_1153,N_1186);
or U1228 (N_1228,N_1152,N_1163);
nor U1229 (N_1229,N_1169,N_1193);
and U1230 (N_1230,N_1172,N_1197);
and U1231 (N_1231,N_1195,N_1171);
and U1232 (N_1232,N_1154,N_1177);
nor U1233 (N_1233,N_1153,N_1159);
and U1234 (N_1234,N_1185,N_1175);
nor U1235 (N_1235,N_1196,N_1181);
and U1236 (N_1236,N_1176,N_1169);
or U1237 (N_1237,N_1188,N_1180);
and U1238 (N_1238,N_1156,N_1162);
nand U1239 (N_1239,N_1160,N_1164);
nor U1240 (N_1240,N_1159,N_1162);
or U1241 (N_1241,N_1167,N_1154);
or U1242 (N_1242,N_1146,N_1168);
and U1243 (N_1243,N_1178,N_1152);
nor U1244 (N_1244,N_1198,N_1195);
or U1245 (N_1245,N_1146,N_1185);
and U1246 (N_1246,N_1189,N_1163);
or U1247 (N_1247,N_1144,N_1179);
nand U1248 (N_1248,N_1149,N_1152);
and U1249 (N_1249,N_1167,N_1169);
or U1250 (N_1250,N_1168,N_1177);
nand U1251 (N_1251,N_1141,N_1157);
nor U1252 (N_1252,N_1168,N_1171);
or U1253 (N_1253,N_1158,N_1190);
nand U1254 (N_1254,N_1174,N_1154);
nand U1255 (N_1255,N_1156,N_1196);
or U1256 (N_1256,N_1197,N_1183);
or U1257 (N_1257,N_1151,N_1171);
nand U1258 (N_1258,N_1171,N_1170);
nand U1259 (N_1259,N_1176,N_1152);
nor U1260 (N_1260,N_1232,N_1225);
nand U1261 (N_1261,N_1207,N_1201);
or U1262 (N_1262,N_1251,N_1218);
and U1263 (N_1263,N_1244,N_1249);
and U1264 (N_1264,N_1226,N_1213);
and U1265 (N_1265,N_1215,N_1212);
and U1266 (N_1266,N_1217,N_1255);
and U1267 (N_1267,N_1200,N_1258);
nor U1268 (N_1268,N_1242,N_1246);
nand U1269 (N_1269,N_1211,N_1245);
nor U1270 (N_1270,N_1238,N_1220);
or U1271 (N_1271,N_1219,N_1229);
and U1272 (N_1272,N_1252,N_1202);
xor U1273 (N_1273,N_1214,N_1234);
or U1274 (N_1274,N_1236,N_1247);
and U1275 (N_1275,N_1203,N_1254);
nor U1276 (N_1276,N_1209,N_1235);
and U1277 (N_1277,N_1223,N_1250);
nand U1278 (N_1278,N_1205,N_1253);
nand U1279 (N_1279,N_1243,N_1231);
or U1280 (N_1280,N_1228,N_1248);
and U1281 (N_1281,N_1224,N_1239);
xnor U1282 (N_1282,N_1206,N_1241);
or U1283 (N_1283,N_1233,N_1222);
or U1284 (N_1284,N_1208,N_1216);
and U1285 (N_1285,N_1240,N_1204);
nand U1286 (N_1286,N_1221,N_1256);
xor U1287 (N_1287,N_1227,N_1259);
and U1288 (N_1288,N_1210,N_1257);
nand U1289 (N_1289,N_1237,N_1230);
and U1290 (N_1290,N_1236,N_1232);
and U1291 (N_1291,N_1212,N_1219);
xnor U1292 (N_1292,N_1214,N_1227);
nor U1293 (N_1293,N_1212,N_1220);
nand U1294 (N_1294,N_1229,N_1234);
xnor U1295 (N_1295,N_1221,N_1251);
nand U1296 (N_1296,N_1244,N_1245);
nand U1297 (N_1297,N_1221,N_1254);
and U1298 (N_1298,N_1255,N_1209);
nor U1299 (N_1299,N_1249,N_1200);
nor U1300 (N_1300,N_1239,N_1230);
or U1301 (N_1301,N_1237,N_1217);
nor U1302 (N_1302,N_1257,N_1252);
xnor U1303 (N_1303,N_1230,N_1202);
nor U1304 (N_1304,N_1235,N_1206);
and U1305 (N_1305,N_1236,N_1239);
nor U1306 (N_1306,N_1228,N_1200);
or U1307 (N_1307,N_1257,N_1215);
nand U1308 (N_1308,N_1243,N_1230);
nor U1309 (N_1309,N_1248,N_1245);
and U1310 (N_1310,N_1248,N_1204);
nor U1311 (N_1311,N_1239,N_1256);
and U1312 (N_1312,N_1203,N_1216);
or U1313 (N_1313,N_1212,N_1206);
nor U1314 (N_1314,N_1230,N_1256);
and U1315 (N_1315,N_1220,N_1217);
and U1316 (N_1316,N_1241,N_1224);
or U1317 (N_1317,N_1230,N_1211);
nand U1318 (N_1318,N_1227,N_1239);
nand U1319 (N_1319,N_1201,N_1219);
and U1320 (N_1320,N_1276,N_1275);
and U1321 (N_1321,N_1282,N_1260);
nor U1322 (N_1322,N_1307,N_1304);
xnor U1323 (N_1323,N_1311,N_1286);
nand U1324 (N_1324,N_1301,N_1317);
nand U1325 (N_1325,N_1262,N_1313);
nor U1326 (N_1326,N_1294,N_1271);
and U1327 (N_1327,N_1278,N_1303);
or U1328 (N_1328,N_1279,N_1280);
or U1329 (N_1329,N_1298,N_1316);
or U1330 (N_1330,N_1269,N_1305);
nand U1331 (N_1331,N_1285,N_1300);
or U1332 (N_1332,N_1264,N_1295);
xnor U1333 (N_1333,N_1288,N_1291);
or U1334 (N_1334,N_1266,N_1293);
or U1335 (N_1335,N_1310,N_1263);
nand U1336 (N_1336,N_1272,N_1277);
and U1337 (N_1337,N_1267,N_1284);
or U1338 (N_1338,N_1314,N_1309);
or U1339 (N_1339,N_1281,N_1268);
and U1340 (N_1340,N_1297,N_1261);
nor U1341 (N_1341,N_1265,N_1289);
nand U1342 (N_1342,N_1296,N_1302);
nor U1343 (N_1343,N_1270,N_1306);
and U1344 (N_1344,N_1290,N_1274);
and U1345 (N_1345,N_1299,N_1315);
and U1346 (N_1346,N_1283,N_1273);
nor U1347 (N_1347,N_1312,N_1292);
nand U1348 (N_1348,N_1319,N_1318);
and U1349 (N_1349,N_1287,N_1308);
or U1350 (N_1350,N_1311,N_1279);
nand U1351 (N_1351,N_1264,N_1278);
nand U1352 (N_1352,N_1294,N_1268);
or U1353 (N_1353,N_1285,N_1319);
and U1354 (N_1354,N_1284,N_1300);
nand U1355 (N_1355,N_1298,N_1288);
and U1356 (N_1356,N_1309,N_1262);
nor U1357 (N_1357,N_1294,N_1289);
or U1358 (N_1358,N_1311,N_1292);
nand U1359 (N_1359,N_1276,N_1268);
and U1360 (N_1360,N_1266,N_1284);
and U1361 (N_1361,N_1274,N_1285);
nand U1362 (N_1362,N_1286,N_1266);
nor U1363 (N_1363,N_1313,N_1291);
or U1364 (N_1364,N_1305,N_1297);
nor U1365 (N_1365,N_1274,N_1272);
or U1366 (N_1366,N_1304,N_1302);
and U1367 (N_1367,N_1293,N_1319);
or U1368 (N_1368,N_1317,N_1271);
and U1369 (N_1369,N_1296,N_1285);
or U1370 (N_1370,N_1276,N_1298);
or U1371 (N_1371,N_1266,N_1305);
nor U1372 (N_1372,N_1270,N_1265);
nand U1373 (N_1373,N_1292,N_1262);
or U1374 (N_1374,N_1281,N_1270);
or U1375 (N_1375,N_1301,N_1283);
xnor U1376 (N_1376,N_1281,N_1302);
nor U1377 (N_1377,N_1319,N_1286);
or U1378 (N_1378,N_1280,N_1300);
nor U1379 (N_1379,N_1260,N_1310);
xnor U1380 (N_1380,N_1353,N_1379);
nand U1381 (N_1381,N_1344,N_1358);
xor U1382 (N_1382,N_1357,N_1340);
nand U1383 (N_1383,N_1332,N_1327);
and U1384 (N_1384,N_1337,N_1326);
and U1385 (N_1385,N_1361,N_1331);
and U1386 (N_1386,N_1378,N_1376);
xor U1387 (N_1387,N_1338,N_1330);
or U1388 (N_1388,N_1370,N_1374);
nor U1389 (N_1389,N_1350,N_1354);
xor U1390 (N_1390,N_1321,N_1364);
and U1391 (N_1391,N_1372,N_1329);
nor U1392 (N_1392,N_1328,N_1371);
nand U1393 (N_1393,N_1373,N_1334);
nor U1394 (N_1394,N_1342,N_1368);
nor U1395 (N_1395,N_1362,N_1367);
or U1396 (N_1396,N_1346,N_1360);
nor U1397 (N_1397,N_1345,N_1341);
nor U1398 (N_1398,N_1356,N_1363);
or U1399 (N_1399,N_1366,N_1320);
nand U1400 (N_1400,N_1325,N_1377);
nor U1401 (N_1401,N_1339,N_1351);
and U1402 (N_1402,N_1348,N_1333);
xor U1403 (N_1403,N_1349,N_1352);
xor U1404 (N_1404,N_1375,N_1322);
nor U1405 (N_1405,N_1335,N_1323);
nor U1406 (N_1406,N_1324,N_1355);
nor U1407 (N_1407,N_1359,N_1365);
and U1408 (N_1408,N_1336,N_1347);
nor U1409 (N_1409,N_1369,N_1343);
nor U1410 (N_1410,N_1372,N_1345);
nor U1411 (N_1411,N_1322,N_1343);
nand U1412 (N_1412,N_1352,N_1377);
or U1413 (N_1413,N_1330,N_1336);
nand U1414 (N_1414,N_1362,N_1343);
or U1415 (N_1415,N_1342,N_1369);
and U1416 (N_1416,N_1340,N_1333);
nand U1417 (N_1417,N_1326,N_1356);
nand U1418 (N_1418,N_1341,N_1354);
nor U1419 (N_1419,N_1326,N_1371);
nor U1420 (N_1420,N_1320,N_1342);
xor U1421 (N_1421,N_1348,N_1362);
nor U1422 (N_1422,N_1321,N_1346);
nor U1423 (N_1423,N_1320,N_1371);
or U1424 (N_1424,N_1344,N_1339);
and U1425 (N_1425,N_1368,N_1327);
nand U1426 (N_1426,N_1328,N_1350);
nor U1427 (N_1427,N_1323,N_1369);
xnor U1428 (N_1428,N_1337,N_1352);
nand U1429 (N_1429,N_1344,N_1329);
nand U1430 (N_1430,N_1362,N_1325);
nand U1431 (N_1431,N_1344,N_1340);
nand U1432 (N_1432,N_1355,N_1366);
or U1433 (N_1433,N_1322,N_1350);
nand U1434 (N_1434,N_1377,N_1356);
and U1435 (N_1435,N_1349,N_1334);
nand U1436 (N_1436,N_1348,N_1327);
or U1437 (N_1437,N_1348,N_1364);
or U1438 (N_1438,N_1349,N_1354);
xnor U1439 (N_1439,N_1353,N_1372);
and U1440 (N_1440,N_1426,N_1411);
nand U1441 (N_1441,N_1410,N_1399);
nor U1442 (N_1442,N_1394,N_1391);
and U1443 (N_1443,N_1390,N_1420);
and U1444 (N_1444,N_1428,N_1421);
nor U1445 (N_1445,N_1424,N_1423);
nor U1446 (N_1446,N_1401,N_1415);
nand U1447 (N_1447,N_1407,N_1404);
xor U1448 (N_1448,N_1400,N_1432);
nand U1449 (N_1449,N_1405,N_1402);
or U1450 (N_1450,N_1385,N_1425);
and U1451 (N_1451,N_1431,N_1389);
nand U1452 (N_1452,N_1436,N_1384);
nand U1453 (N_1453,N_1388,N_1435);
nand U1454 (N_1454,N_1403,N_1419);
nand U1455 (N_1455,N_1406,N_1416);
nand U1456 (N_1456,N_1414,N_1433);
nand U1457 (N_1457,N_1437,N_1439);
and U1458 (N_1458,N_1383,N_1430);
or U1459 (N_1459,N_1387,N_1427);
nor U1460 (N_1460,N_1393,N_1408);
and U1461 (N_1461,N_1398,N_1395);
and U1462 (N_1462,N_1413,N_1438);
xor U1463 (N_1463,N_1397,N_1417);
and U1464 (N_1464,N_1409,N_1412);
or U1465 (N_1465,N_1396,N_1429);
or U1466 (N_1466,N_1381,N_1422);
and U1467 (N_1467,N_1380,N_1386);
and U1468 (N_1468,N_1418,N_1392);
nand U1469 (N_1469,N_1382,N_1434);
and U1470 (N_1470,N_1381,N_1401);
and U1471 (N_1471,N_1404,N_1431);
nand U1472 (N_1472,N_1389,N_1422);
or U1473 (N_1473,N_1409,N_1389);
nand U1474 (N_1474,N_1387,N_1401);
nand U1475 (N_1475,N_1428,N_1407);
xnor U1476 (N_1476,N_1398,N_1382);
nor U1477 (N_1477,N_1424,N_1434);
or U1478 (N_1478,N_1409,N_1393);
xor U1479 (N_1479,N_1402,N_1401);
nand U1480 (N_1480,N_1389,N_1406);
nand U1481 (N_1481,N_1408,N_1438);
or U1482 (N_1482,N_1412,N_1415);
nor U1483 (N_1483,N_1435,N_1415);
xor U1484 (N_1484,N_1438,N_1383);
or U1485 (N_1485,N_1397,N_1410);
or U1486 (N_1486,N_1417,N_1434);
nor U1487 (N_1487,N_1414,N_1387);
nand U1488 (N_1488,N_1402,N_1389);
nand U1489 (N_1489,N_1407,N_1398);
or U1490 (N_1490,N_1389,N_1404);
xor U1491 (N_1491,N_1424,N_1385);
xor U1492 (N_1492,N_1383,N_1425);
nor U1493 (N_1493,N_1434,N_1385);
or U1494 (N_1494,N_1392,N_1429);
xnor U1495 (N_1495,N_1384,N_1418);
and U1496 (N_1496,N_1426,N_1433);
nor U1497 (N_1497,N_1431,N_1391);
nand U1498 (N_1498,N_1395,N_1383);
nand U1499 (N_1499,N_1400,N_1424);
and U1500 (N_1500,N_1450,N_1467);
or U1501 (N_1501,N_1458,N_1463);
xor U1502 (N_1502,N_1454,N_1472);
and U1503 (N_1503,N_1497,N_1477);
nand U1504 (N_1504,N_1480,N_1493);
or U1505 (N_1505,N_1496,N_1452);
or U1506 (N_1506,N_1498,N_1494);
nand U1507 (N_1507,N_1475,N_1487);
xor U1508 (N_1508,N_1441,N_1446);
or U1509 (N_1509,N_1453,N_1462);
nand U1510 (N_1510,N_1444,N_1492);
and U1511 (N_1511,N_1499,N_1466);
nor U1512 (N_1512,N_1461,N_1442);
or U1513 (N_1513,N_1473,N_1485);
or U1514 (N_1514,N_1495,N_1449);
or U1515 (N_1515,N_1479,N_1464);
xnor U1516 (N_1516,N_1468,N_1476);
nor U1517 (N_1517,N_1471,N_1456);
or U1518 (N_1518,N_1457,N_1491);
nand U1519 (N_1519,N_1469,N_1474);
and U1520 (N_1520,N_1447,N_1470);
nor U1521 (N_1521,N_1445,N_1488);
or U1522 (N_1522,N_1478,N_1465);
or U1523 (N_1523,N_1483,N_1486);
or U1524 (N_1524,N_1460,N_1484);
or U1525 (N_1525,N_1490,N_1489);
nand U1526 (N_1526,N_1440,N_1443);
nand U1527 (N_1527,N_1482,N_1455);
nor U1528 (N_1528,N_1448,N_1451);
and U1529 (N_1529,N_1459,N_1481);
or U1530 (N_1530,N_1466,N_1443);
nor U1531 (N_1531,N_1477,N_1464);
xor U1532 (N_1532,N_1490,N_1462);
and U1533 (N_1533,N_1475,N_1454);
and U1534 (N_1534,N_1448,N_1440);
xor U1535 (N_1535,N_1465,N_1441);
or U1536 (N_1536,N_1478,N_1486);
xor U1537 (N_1537,N_1476,N_1444);
nand U1538 (N_1538,N_1484,N_1475);
nor U1539 (N_1539,N_1444,N_1454);
and U1540 (N_1540,N_1482,N_1475);
nor U1541 (N_1541,N_1474,N_1488);
and U1542 (N_1542,N_1484,N_1452);
xor U1543 (N_1543,N_1473,N_1483);
nor U1544 (N_1544,N_1460,N_1473);
nor U1545 (N_1545,N_1481,N_1490);
or U1546 (N_1546,N_1446,N_1487);
nand U1547 (N_1547,N_1499,N_1470);
or U1548 (N_1548,N_1482,N_1483);
nor U1549 (N_1549,N_1461,N_1462);
xnor U1550 (N_1550,N_1455,N_1462);
nor U1551 (N_1551,N_1487,N_1482);
nor U1552 (N_1552,N_1497,N_1485);
xnor U1553 (N_1553,N_1487,N_1494);
or U1554 (N_1554,N_1485,N_1460);
nor U1555 (N_1555,N_1456,N_1490);
or U1556 (N_1556,N_1454,N_1489);
nand U1557 (N_1557,N_1482,N_1474);
or U1558 (N_1558,N_1483,N_1460);
nor U1559 (N_1559,N_1479,N_1494);
or U1560 (N_1560,N_1521,N_1524);
nand U1561 (N_1561,N_1531,N_1508);
nor U1562 (N_1562,N_1504,N_1530);
and U1563 (N_1563,N_1536,N_1554);
and U1564 (N_1564,N_1505,N_1526);
nand U1565 (N_1565,N_1546,N_1552);
and U1566 (N_1566,N_1532,N_1529);
nor U1567 (N_1567,N_1544,N_1512);
nor U1568 (N_1568,N_1543,N_1517);
nor U1569 (N_1569,N_1500,N_1547);
or U1570 (N_1570,N_1539,N_1520);
nand U1571 (N_1571,N_1557,N_1537);
nor U1572 (N_1572,N_1556,N_1516);
nand U1573 (N_1573,N_1511,N_1527);
nand U1574 (N_1574,N_1506,N_1549);
nor U1575 (N_1575,N_1535,N_1501);
and U1576 (N_1576,N_1514,N_1513);
and U1577 (N_1577,N_1559,N_1545);
xor U1578 (N_1578,N_1548,N_1555);
nor U1579 (N_1579,N_1502,N_1558);
nor U1580 (N_1580,N_1528,N_1541);
or U1581 (N_1581,N_1534,N_1510);
and U1582 (N_1582,N_1503,N_1522);
nor U1583 (N_1583,N_1518,N_1519);
xnor U1584 (N_1584,N_1553,N_1550);
xnor U1585 (N_1585,N_1507,N_1542);
nor U1586 (N_1586,N_1540,N_1509);
and U1587 (N_1587,N_1533,N_1523);
nor U1588 (N_1588,N_1515,N_1551);
nand U1589 (N_1589,N_1538,N_1525);
nor U1590 (N_1590,N_1550,N_1514);
or U1591 (N_1591,N_1558,N_1504);
and U1592 (N_1592,N_1541,N_1516);
nand U1593 (N_1593,N_1523,N_1522);
nor U1594 (N_1594,N_1553,N_1514);
and U1595 (N_1595,N_1546,N_1506);
nand U1596 (N_1596,N_1509,N_1526);
or U1597 (N_1597,N_1502,N_1505);
nand U1598 (N_1598,N_1535,N_1537);
and U1599 (N_1599,N_1524,N_1508);
or U1600 (N_1600,N_1521,N_1543);
nor U1601 (N_1601,N_1516,N_1543);
and U1602 (N_1602,N_1518,N_1528);
nand U1603 (N_1603,N_1523,N_1501);
or U1604 (N_1604,N_1532,N_1552);
and U1605 (N_1605,N_1533,N_1500);
nand U1606 (N_1606,N_1550,N_1508);
and U1607 (N_1607,N_1506,N_1508);
and U1608 (N_1608,N_1547,N_1535);
xor U1609 (N_1609,N_1525,N_1516);
and U1610 (N_1610,N_1502,N_1503);
or U1611 (N_1611,N_1521,N_1530);
nand U1612 (N_1612,N_1550,N_1524);
or U1613 (N_1613,N_1556,N_1526);
and U1614 (N_1614,N_1544,N_1502);
nor U1615 (N_1615,N_1546,N_1525);
xnor U1616 (N_1616,N_1541,N_1512);
or U1617 (N_1617,N_1541,N_1534);
nor U1618 (N_1618,N_1517,N_1539);
nor U1619 (N_1619,N_1536,N_1509);
nor U1620 (N_1620,N_1565,N_1560);
nor U1621 (N_1621,N_1579,N_1583);
nand U1622 (N_1622,N_1593,N_1569);
nand U1623 (N_1623,N_1577,N_1568);
and U1624 (N_1624,N_1605,N_1561);
or U1625 (N_1625,N_1570,N_1590);
nor U1626 (N_1626,N_1607,N_1611);
nand U1627 (N_1627,N_1609,N_1566);
or U1628 (N_1628,N_1571,N_1600);
nand U1629 (N_1629,N_1602,N_1585);
or U1630 (N_1630,N_1610,N_1581);
nand U1631 (N_1631,N_1586,N_1604);
or U1632 (N_1632,N_1563,N_1598);
and U1633 (N_1633,N_1573,N_1589);
nor U1634 (N_1634,N_1584,N_1576);
or U1635 (N_1635,N_1617,N_1608);
or U1636 (N_1636,N_1580,N_1603);
or U1637 (N_1637,N_1596,N_1615);
or U1638 (N_1638,N_1618,N_1562);
or U1639 (N_1639,N_1614,N_1594);
and U1640 (N_1640,N_1564,N_1613);
xnor U1641 (N_1641,N_1616,N_1572);
and U1642 (N_1642,N_1595,N_1597);
nand U1643 (N_1643,N_1574,N_1567);
nand U1644 (N_1644,N_1588,N_1599);
nand U1645 (N_1645,N_1591,N_1612);
nand U1646 (N_1646,N_1575,N_1592);
nor U1647 (N_1647,N_1601,N_1578);
nor U1648 (N_1648,N_1582,N_1606);
and U1649 (N_1649,N_1619,N_1587);
xnor U1650 (N_1650,N_1563,N_1612);
nor U1651 (N_1651,N_1563,N_1578);
xnor U1652 (N_1652,N_1585,N_1606);
nand U1653 (N_1653,N_1565,N_1589);
or U1654 (N_1654,N_1604,N_1560);
and U1655 (N_1655,N_1573,N_1569);
xnor U1656 (N_1656,N_1567,N_1565);
or U1657 (N_1657,N_1560,N_1567);
and U1658 (N_1658,N_1585,N_1610);
and U1659 (N_1659,N_1579,N_1586);
or U1660 (N_1660,N_1582,N_1577);
nand U1661 (N_1661,N_1604,N_1583);
nand U1662 (N_1662,N_1566,N_1589);
xor U1663 (N_1663,N_1606,N_1570);
nand U1664 (N_1664,N_1564,N_1584);
or U1665 (N_1665,N_1570,N_1595);
xor U1666 (N_1666,N_1598,N_1612);
nand U1667 (N_1667,N_1587,N_1576);
or U1668 (N_1668,N_1611,N_1568);
and U1669 (N_1669,N_1608,N_1578);
or U1670 (N_1670,N_1581,N_1594);
or U1671 (N_1671,N_1574,N_1615);
xnor U1672 (N_1672,N_1613,N_1618);
nor U1673 (N_1673,N_1616,N_1611);
or U1674 (N_1674,N_1593,N_1589);
and U1675 (N_1675,N_1608,N_1606);
or U1676 (N_1676,N_1578,N_1597);
or U1677 (N_1677,N_1578,N_1605);
and U1678 (N_1678,N_1576,N_1580);
nor U1679 (N_1679,N_1605,N_1576);
nand U1680 (N_1680,N_1673,N_1628);
or U1681 (N_1681,N_1649,N_1632);
xnor U1682 (N_1682,N_1631,N_1651);
or U1683 (N_1683,N_1624,N_1662);
nand U1684 (N_1684,N_1636,N_1650);
nor U1685 (N_1685,N_1653,N_1664);
nand U1686 (N_1686,N_1626,N_1674);
nand U1687 (N_1687,N_1676,N_1622);
and U1688 (N_1688,N_1655,N_1641);
xor U1689 (N_1689,N_1668,N_1658);
nand U1690 (N_1690,N_1675,N_1669);
nor U1691 (N_1691,N_1635,N_1640);
and U1692 (N_1692,N_1679,N_1678);
or U1693 (N_1693,N_1644,N_1638);
and U1694 (N_1694,N_1625,N_1659);
or U1695 (N_1695,N_1657,N_1630);
nand U1696 (N_1696,N_1670,N_1656);
or U1697 (N_1697,N_1661,N_1633);
and U1698 (N_1698,N_1627,N_1620);
nor U1699 (N_1699,N_1643,N_1648);
nand U1700 (N_1700,N_1634,N_1665);
and U1701 (N_1701,N_1637,N_1621);
or U1702 (N_1702,N_1671,N_1646);
nor U1703 (N_1703,N_1642,N_1645);
or U1704 (N_1704,N_1667,N_1639);
nand U1705 (N_1705,N_1654,N_1647);
nor U1706 (N_1706,N_1677,N_1663);
nor U1707 (N_1707,N_1660,N_1629);
nand U1708 (N_1708,N_1652,N_1623);
and U1709 (N_1709,N_1672,N_1666);
or U1710 (N_1710,N_1639,N_1636);
and U1711 (N_1711,N_1662,N_1675);
nor U1712 (N_1712,N_1628,N_1631);
or U1713 (N_1713,N_1656,N_1653);
or U1714 (N_1714,N_1675,N_1626);
nand U1715 (N_1715,N_1671,N_1630);
and U1716 (N_1716,N_1646,N_1634);
xor U1717 (N_1717,N_1666,N_1621);
or U1718 (N_1718,N_1637,N_1620);
or U1719 (N_1719,N_1656,N_1671);
or U1720 (N_1720,N_1670,N_1679);
nand U1721 (N_1721,N_1675,N_1636);
and U1722 (N_1722,N_1641,N_1639);
nand U1723 (N_1723,N_1648,N_1678);
and U1724 (N_1724,N_1641,N_1663);
nor U1725 (N_1725,N_1642,N_1629);
nor U1726 (N_1726,N_1658,N_1622);
or U1727 (N_1727,N_1653,N_1674);
and U1728 (N_1728,N_1648,N_1630);
nand U1729 (N_1729,N_1643,N_1624);
and U1730 (N_1730,N_1635,N_1672);
or U1731 (N_1731,N_1632,N_1648);
nor U1732 (N_1732,N_1636,N_1630);
xnor U1733 (N_1733,N_1640,N_1657);
and U1734 (N_1734,N_1643,N_1620);
or U1735 (N_1735,N_1631,N_1620);
and U1736 (N_1736,N_1624,N_1657);
nand U1737 (N_1737,N_1657,N_1652);
xnor U1738 (N_1738,N_1674,N_1665);
or U1739 (N_1739,N_1649,N_1654);
or U1740 (N_1740,N_1705,N_1703);
nand U1741 (N_1741,N_1715,N_1712);
nand U1742 (N_1742,N_1735,N_1700);
nor U1743 (N_1743,N_1718,N_1734);
nor U1744 (N_1744,N_1682,N_1719);
nand U1745 (N_1745,N_1683,N_1710);
nor U1746 (N_1746,N_1707,N_1680);
xnor U1747 (N_1747,N_1696,N_1685);
or U1748 (N_1748,N_1697,N_1692);
nor U1749 (N_1749,N_1691,N_1732);
nor U1750 (N_1750,N_1727,N_1731);
or U1751 (N_1751,N_1686,N_1716);
xor U1752 (N_1752,N_1699,N_1693);
and U1753 (N_1753,N_1725,N_1724);
nand U1754 (N_1754,N_1730,N_1690);
nand U1755 (N_1755,N_1739,N_1706);
nor U1756 (N_1756,N_1688,N_1709);
xor U1757 (N_1757,N_1684,N_1698);
xor U1758 (N_1758,N_1736,N_1713);
xnor U1759 (N_1759,N_1701,N_1704);
and U1760 (N_1760,N_1689,N_1694);
nand U1761 (N_1761,N_1738,N_1726);
and U1762 (N_1762,N_1729,N_1728);
and U1763 (N_1763,N_1723,N_1681);
or U1764 (N_1764,N_1717,N_1720);
nand U1765 (N_1765,N_1737,N_1687);
or U1766 (N_1766,N_1714,N_1722);
and U1767 (N_1767,N_1702,N_1711);
and U1768 (N_1768,N_1695,N_1708);
or U1769 (N_1769,N_1733,N_1721);
or U1770 (N_1770,N_1690,N_1733);
nor U1771 (N_1771,N_1695,N_1703);
nand U1772 (N_1772,N_1731,N_1693);
or U1773 (N_1773,N_1697,N_1708);
and U1774 (N_1774,N_1718,N_1729);
or U1775 (N_1775,N_1695,N_1680);
or U1776 (N_1776,N_1686,N_1702);
nand U1777 (N_1777,N_1717,N_1701);
nand U1778 (N_1778,N_1708,N_1702);
nand U1779 (N_1779,N_1703,N_1715);
xor U1780 (N_1780,N_1723,N_1696);
xnor U1781 (N_1781,N_1693,N_1702);
or U1782 (N_1782,N_1704,N_1680);
nand U1783 (N_1783,N_1738,N_1724);
nand U1784 (N_1784,N_1694,N_1721);
and U1785 (N_1785,N_1680,N_1715);
or U1786 (N_1786,N_1703,N_1697);
nand U1787 (N_1787,N_1705,N_1682);
and U1788 (N_1788,N_1711,N_1719);
and U1789 (N_1789,N_1691,N_1683);
nand U1790 (N_1790,N_1684,N_1688);
xor U1791 (N_1791,N_1686,N_1727);
xnor U1792 (N_1792,N_1732,N_1719);
nor U1793 (N_1793,N_1729,N_1683);
or U1794 (N_1794,N_1719,N_1710);
and U1795 (N_1795,N_1688,N_1714);
or U1796 (N_1796,N_1724,N_1707);
nor U1797 (N_1797,N_1735,N_1720);
nor U1798 (N_1798,N_1682,N_1730);
and U1799 (N_1799,N_1733,N_1718);
and U1800 (N_1800,N_1787,N_1788);
and U1801 (N_1801,N_1757,N_1777);
nand U1802 (N_1802,N_1795,N_1740);
or U1803 (N_1803,N_1774,N_1741);
or U1804 (N_1804,N_1796,N_1743);
nand U1805 (N_1805,N_1749,N_1750);
xor U1806 (N_1806,N_1752,N_1747);
and U1807 (N_1807,N_1793,N_1746);
and U1808 (N_1808,N_1790,N_1759);
nand U1809 (N_1809,N_1754,N_1764);
nor U1810 (N_1810,N_1789,N_1748);
and U1811 (N_1811,N_1771,N_1791);
or U1812 (N_1812,N_1799,N_1753);
and U1813 (N_1813,N_1762,N_1772);
and U1814 (N_1814,N_1770,N_1767);
and U1815 (N_1815,N_1784,N_1758);
nand U1816 (N_1816,N_1780,N_1792);
nor U1817 (N_1817,N_1742,N_1773);
nand U1818 (N_1818,N_1745,N_1778);
nor U1819 (N_1819,N_1751,N_1775);
nor U1820 (N_1820,N_1744,N_1798);
or U1821 (N_1821,N_1776,N_1763);
xor U1822 (N_1822,N_1765,N_1782);
or U1823 (N_1823,N_1756,N_1794);
xnor U1824 (N_1824,N_1760,N_1761);
nand U1825 (N_1825,N_1779,N_1766);
nand U1826 (N_1826,N_1786,N_1785);
nor U1827 (N_1827,N_1781,N_1783);
and U1828 (N_1828,N_1768,N_1797);
nor U1829 (N_1829,N_1769,N_1755);
or U1830 (N_1830,N_1772,N_1744);
nand U1831 (N_1831,N_1748,N_1773);
and U1832 (N_1832,N_1763,N_1749);
or U1833 (N_1833,N_1784,N_1770);
or U1834 (N_1834,N_1756,N_1773);
and U1835 (N_1835,N_1798,N_1758);
nand U1836 (N_1836,N_1750,N_1747);
nand U1837 (N_1837,N_1790,N_1781);
xnor U1838 (N_1838,N_1756,N_1772);
and U1839 (N_1839,N_1745,N_1788);
or U1840 (N_1840,N_1787,N_1799);
and U1841 (N_1841,N_1751,N_1758);
nor U1842 (N_1842,N_1761,N_1778);
nand U1843 (N_1843,N_1783,N_1771);
or U1844 (N_1844,N_1757,N_1749);
nand U1845 (N_1845,N_1768,N_1796);
nor U1846 (N_1846,N_1781,N_1756);
and U1847 (N_1847,N_1782,N_1791);
or U1848 (N_1848,N_1752,N_1760);
or U1849 (N_1849,N_1764,N_1782);
and U1850 (N_1850,N_1743,N_1790);
xnor U1851 (N_1851,N_1762,N_1757);
nor U1852 (N_1852,N_1741,N_1779);
or U1853 (N_1853,N_1752,N_1743);
nor U1854 (N_1854,N_1782,N_1774);
nor U1855 (N_1855,N_1756,N_1748);
nor U1856 (N_1856,N_1756,N_1750);
nand U1857 (N_1857,N_1798,N_1782);
and U1858 (N_1858,N_1770,N_1758);
xnor U1859 (N_1859,N_1771,N_1779);
nand U1860 (N_1860,N_1848,N_1819);
or U1861 (N_1861,N_1852,N_1818);
nand U1862 (N_1862,N_1830,N_1847);
nor U1863 (N_1863,N_1810,N_1859);
nor U1864 (N_1864,N_1839,N_1833);
xnor U1865 (N_1865,N_1858,N_1812);
nor U1866 (N_1866,N_1820,N_1829);
nand U1867 (N_1867,N_1807,N_1804);
and U1868 (N_1868,N_1806,N_1809);
nor U1869 (N_1869,N_1803,N_1801);
nor U1870 (N_1870,N_1821,N_1813);
or U1871 (N_1871,N_1814,N_1842);
nor U1872 (N_1872,N_1849,N_1853);
or U1873 (N_1873,N_1822,N_1824);
nand U1874 (N_1874,N_1838,N_1836);
nor U1875 (N_1875,N_1834,N_1855);
xor U1876 (N_1876,N_1840,N_1811);
and U1877 (N_1877,N_1844,N_1856);
nand U1878 (N_1878,N_1846,N_1800);
nor U1879 (N_1879,N_1851,N_1808);
and U1880 (N_1880,N_1835,N_1845);
xor U1881 (N_1881,N_1843,N_1857);
and U1882 (N_1882,N_1827,N_1825);
and U1883 (N_1883,N_1837,N_1826);
or U1884 (N_1884,N_1832,N_1831);
and U1885 (N_1885,N_1805,N_1816);
nor U1886 (N_1886,N_1841,N_1854);
and U1887 (N_1887,N_1817,N_1815);
and U1888 (N_1888,N_1823,N_1828);
or U1889 (N_1889,N_1802,N_1850);
or U1890 (N_1890,N_1811,N_1802);
or U1891 (N_1891,N_1807,N_1826);
nand U1892 (N_1892,N_1821,N_1822);
nand U1893 (N_1893,N_1829,N_1847);
nand U1894 (N_1894,N_1815,N_1841);
nor U1895 (N_1895,N_1810,N_1843);
nand U1896 (N_1896,N_1839,N_1827);
nor U1897 (N_1897,N_1842,N_1848);
nand U1898 (N_1898,N_1813,N_1825);
or U1899 (N_1899,N_1807,N_1800);
and U1900 (N_1900,N_1820,N_1833);
or U1901 (N_1901,N_1810,N_1813);
and U1902 (N_1902,N_1802,N_1854);
nand U1903 (N_1903,N_1839,N_1844);
nor U1904 (N_1904,N_1818,N_1849);
nor U1905 (N_1905,N_1857,N_1848);
and U1906 (N_1906,N_1820,N_1809);
and U1907 (N_1907,N_1819,N_1805);
or U1908 (N_1908,N_1820,N_1841);
nor U1909 (N_1909,N_1805,N_1800);
nor U1910 (N_1910,N_1823,N_1843);
nor U1911 (N_1911,N_1858,N_1851);
nor U1912 (N_1912,N_1842,N_1836);
nand U1913 (N_1913,N_1816,N_1828);
or U1914 (N_1914,N_1808,N_1826);
xnor U1915 (N_1915,N_1843,N_1807);
or U1916 (N_1916,N_1801,N_1854);
nor U1917 (N_1917,N_1814,N_1820);
or U1918 (N_1918,N_1817,N_1852);
or U1919 (N_1919,N_1845,N_1811);
xor U1920 (N_1920,N_1885,N_1916);
xor U1921 (N_1921,N_1896,N_1917);
nor U1922 (N_1922,N_1882,N_1900);
nand U1923 (N_1923,N_1912,N_1863);
and U1924 (N_1924,N_1918,N_1879);
and U1925 (N_1925,N_1899,N_1864);
nor U1926 (N_1926,N_1908,N_1867);
nor U1927 (N_1927,N_1889,N_1870);
xor U1928 (N_1928,N_1868,N_1888);
nand U1929 (N_1929,N_1874,N_1890);
nand U1930 (N_1930,N_1895,N_1903);
and U1931 (N_1931,N_1913,N_1872);
nor U1932 (N_1932,N_1919,N_1907);
or U1933 (N_1933,N_1876,N_1881);
xnor U1934 (N_1934,N_1898,N_1894);
or U1935 (N_1935,N_1884,N_1914);
or U1936 (N_1936,N_1891,N_1862);
nor U1937 (N_1937,N_1911,N_1880);
nand U1938 (N_1938,N_1873,N_1906);
nor U1939 (N_1939,N_1861,N_1902);
nand U1940 (N_1940,N_1886,N_1893);
and U1941 (N_1941,N_1905,N_1883);
and U1942 (N_1942,N_1915,N_1877);
nand U1943 (N_1943,N_1897,N_1910);
and U1944 (N_1944,N_1860,N_1875);
and U1945 (N_1945,N_1901,N_1871);
nand U1946 (N_1946,N_1865,N_1887);
nand U1947 (N_1947,N_1878,N_1869);
nor U1948 (N_1948,N_1892,N_1904);
nor U1949 (N_1949,N_1866,N_1909);
nor U1950 (N_1950,N_1913,N_1884);
nor U1951 (N_1951,N_1903,N_1907);
or U1952 (N_1952,N_1886,N_1904);
and U1953 (N_1953,N_1891,N_1880);
nor U1954 (N_1954,N_1901,N_1861);
nor U1955 (N_1955,N_1870,N_1875);
nand U1956 (N_1956,N_1877,N_1878);
or U1957 (N_1957,N_1873,N_1882);
and U1958 (N_1958,N_1902,N_1872);
nor U1959 (N_1959,N_1891,N_1871);
or U1960 (N_1960,N_1872,N_1877);
nand U1961 (N_1961,N_1860,N_1916);
nor U1962 (N_1962,N_1879,N_1896);
or U1963 (N_1963,N_1899,N_1907);
or U1964 (N_1964,N_1883,N_1910);
xnor U1965 (N_1965,N_1863,N_1883);
nor U1966 (N_1966,N_1891,N_1876);
nand U1967 (N_1967,N_1913,N_1918);
or U1968 (N_1968,N_1892,N_1891);
or U1969 (N_1969,N_1881,N_1888);
or U1970 (N_1970,N_1916,N_1871);
or U1971 (N_1971,N_1865,N_1889);
or U1972 (N_1972,N_1880,N_1871);
nor U1973 (N_1973,N_1868,N_1886);
nor U1974 (N_1974,N_1918,N_1863);
nand U1975 (N_1975,N_1866,N_1888);
and U1976 (N_1976,N_1868,N_1873);
nor U1977 (N_1977,N_1870,N_1903);
nand U1978 (N_1978,N_1910,N_1903);
or U1979 (N_1979,N_1902,N_1919);
nor U1980 (N_1980,N_1936,N_1941);
and U1981 (N_1981,N_1946,N_1923);
and U1982 (N_1982,N_1933,N_1934);
nor U1983 (N_1983,N_1974,N_1954);
nand U1984 (N_1984,N_1953,N_1945);
nand U1985 (N_1985,N_1968,N_1966);
nand U1986 (N_1986,N_1972,N_1926);
nand U1987 (N_1987,N_1927,N_1958);
nor U1988 (N_1988,N_1931,N_1967);
nand U1989 (N_1989,N_1952,N_1962);
nand U1990 (N_1990,N_1938,N_1957);
and U1991 (N_1991,N_1955,N_1947);
and U1992 (N_1992,N_1930,N_1956);
nor U1993 (N_1993,N_1963,N_1970);
or U1994 (N_1994,N_1940,N_1929);
or U1995 (N_1995,N_1921,N_1965);
nor U1996 (N_1996,N_1979,N_1975);
nand U1997 (N_1997,N_1937,N_1977);
or U1998 (N_1998,N_1976,N_1924);
nor U1999 (N_1999,N_1960,N_1973);
nor U2000 (N_2000,N_1942,N_1935);
nand U2001 (N_2001,N_1943,N_1944);
and U2002 (N_2002,N_1932,N_1961);
xnor U2003 (N_2003,N_1928,N_1948);
and U2004 (N_2004,N_1978,N_1951);
nor U2005 (N_2005,N_1922,N_1939);
and U2006 (N_2006,N_1925,N_1964);
nor U2007 (N_2007,N_1971,N_1959);
and U2008 (N_2008,N_1950,N_1920);
nand U2009 (N_2009,N_1969,N_1949);
or U2010 (N_2010,N_1952,N_1932);
nand U2011 (N_2011,N_1975,N_1959);
nand U2012 (N_2012,N_1943,N_1929);
nand U2013 (N_2013,N_1933,N_1971);
and U2014 (N_2014,N_1961,N_1970);
nand U2015 (N_2015,N_1954,N_1933);
nand U2016 (N_2016,N_1930,N_1929);
and U2017 (N_2017,N_1964,N_1950);
and U2018 (N_2018,N_1942,N_1974);
and U2019 (N_2019,N_1939,N_1956);
nand U2020 (N_2020,N_1924,N_1949);
or U2021 (N_2021,N_1969,N_1921);
nand U2022 (N_2022,N_1955,N_1963);
nor U2023 (N_2023,N_1943,N_1938);
or U2024 (N_2024,N_1962,N_1936);
nand U2025 (N_2025,N_1940,N_1958);
nor U2026 (N_2026,N_1927,N_1968);
nand U2027 (N_2027,N_1960,N_1953);
nand U2028 (N_2028,N_1968,N_1955);
or U2029 (N_2029,N_1974,N_1958);
nor U2030 (N_2030,N_1973,N_1966);
nor U2031 (N_2031,N_1959,N_1943);
xnor U2032 (N_2032,N_1970,N_1957);
and U2033 (N_2033,N_1939,N_1934);
and U2034 (N_2034,N_1947,N_1961);
and U2035 (N_2035,N_1920,N_1976);
and U2036 (N_2036,N_1946,N_1928);
xor U2037 (N_2037,N_1957,N_1926);
or U2038 (N_2038,N_1921,N_1940);
or U2039 (N_2039,N_1954,N_1945);
or U2040 (N_2040,N_1983,N_2019);
nand U2041 (N_2041,N_2038,N_2007);
or U2042 (N_2042,N_2001,N_1990);
nand U2043 (N_2043,N_1991,N_1998);
nand U2044 (N_2044,N_2005,N_2022);
nand U2045 (N_2045,N_2037,N_1997);
and U2046 (N_2046,N_1989,N_2013);
nor U2047 (N_2047,N_1985,N_2000);
xor U2048 (N_2048,N_1999,N_2021);
nor U2049 (N_2049,N_1993,N_2024);
or U2050 (N_2050,N_2025,N_1992);
nor U2051 (N_2051,N_1984,N_2026);
and U2052 (N_2052,N_1986,N_1994);
and U2053 (N_2053,N_2006,N_1995);
or U2054 (N_2054,N_1987,N_2008);
or U2055 (N_2055,N_2018,N_2012);
nand U2056 (N_2056,N_2020,N_2023);
nand U2057 (N_2057,N_1981,N_2039);
nand U2058 (N_2058,N_2004,N_2009);
nand U2059 (N_2059,N_2027,N_1982);
nor U2060 (N_2060,N_2010,N_2031);
or U2061 (N_2061,N_2034,N_1980);
and U2062 (N_2062,N_2036,N_1988);
or U2063 (N_2063,N_2030,N_2016);
and U2064 (N_2064,N_2035,N_2029);
and U2065 (N_2065,N_2003,N_1996);
or U2066 (N_2066,N_2028,N_2014);
nand U2067 (N_2067,N_2033,N_2032);
or U2068 (N_2068,N_2017,N_2015);
and U2069 (N_2069,N_2002,N_2011);
nor U2070 (N_2070,N_2022,N_1993);
nor U2071 (N_2071,N_1990,N_2005);
and U2072 (N_2072,N_2039,N_1980);
or U2073 (N_2073,N_1984,N_2015);
nand U2074 (N_2074,N_2034,N_2012);
nor U2075 (N_2075,N_1998,N_1981);
nand U2076 (N_2076,N_2039,N_2038);
nand U2077 (N_2077,N_2033,N_2038);
xor U2078 (N_2078,N_1995,N_1990);
and U2079 (N_2079,N_1992,N_2030);
or U2080 (N_2080,N_2002,N_2016);
nand U2081 (N_2081,N_2006,N_1999);
or U2082 (N_2082,N_2025,N_2036);
and U2083 (N_2083,N_1999,N_2019);
nor U2084 (N_2084,N_2021,N_2009);
and U2085 (N_2085,N_2028,N_1993);
nand U2086 (N_2086,N_2015,N_2001);
xor U2087 (N_2087,N_2035,N_1982);
xor U2088 (N_2088,N_2038,N_2016);
xnor U2089 (N_2089,N_2012,N_2025);
nor U2090 (N_2090,N_2020,N_2001);
or U2091 (N_2091,N_2029,N_2018);
and U2092 (N_2092,N_1985,N_2002);
or U2093 (N_2093,N_2037,N_2030);
nand U2094 (N_2094,N_2020,N_2033);
or U2095 (N_2095,N_1987,N_1992);
xnor U2096 (N_2096,N_1989,N_1997);
nor U2097 (N_2097,N_2015,N_1987);
nand U2098 (N_2098,N_2012,N_1983);
and U2099 (N_2099,N_1980,N_2024);
and U2100 (N_2100,N_2087,N_2060);
nor U2101 (N_2101,N_2085,N_2067);
or U2102 (N_2102,N_2096,N_2057);
or U2103 (N_2103,N_2075,N_2099);
xor U2104 (N_2104,N_2040,N_2058);
nand U2105 (N_2105,N_2050,N_2063);
nand U2106 (N_2106,N_2093,N_2077);
and U2107 (N_2107,N_2041,N_2084);
or U2108 (N_2108,N_2079,N_2090);
or U2109 (N_2109,N_2048,N_2051);
nand U2110 (N_2110,N_2054,N_2052);
nand U2111 (N_2111,N_2043,N_2049);
nand U2112 (N_2112,N_2064,N_2097);
nand U2113 (N_2113,N_2055,N_2094);
xnor U2114 (N_2114,N_2092,N_2076);
or U2115 (N_2115,N_2053,N_2073);
and U2116 (N_2116,N_2069,N_2062);
nor U2117 (N_2117,N_2088,N_2066);
and U2118 (N_2118,N_2068,N_2047);
and U2119 (N_2119,N_2046,N_2059);
and U2120 (N_2120,N_2074,N_2056);
nor U2121 (N_2121,N_2045,N_2095);
and U2122 (N_2122,N_2083,N_2082);
nor U2123 (N_2123,N_2098,N_2065);
nand U2124 (N_2124,N_2044,N_2081);
or U2125 (N_2125,N_2061,N_2071);
nand U2126 (N_2126,N_2086,N_2089);
nand U2127 (N_2127,N_2091,N_2080);
and U2128 (N_2128,N_2078,N_2042);
nor U2129 (N_2129,N_2070,N_2072);
nor U2130 (N_2130,N_2061,N_2055);
or U2131 (N_2131,N_2089,N_2079);
and U2132 (N_2132,N_2084,N_2080);
nor U2133 (N_2133,N_2064,N_2096);
or U2134 (N_2134,N_2053,N_2046);
nor U2135 (N_2135,N_2048,N_2081);
nand U2136 (N_2136,N_2061,N_2043);
and U2137 (N_2137,N_2074,N_2050);
or U2138 (N_2138,N_2062,N_2065);
xnor U2139 (N_2139,N_2053,N_2076);
and U2140 (N_2140,N_2040,N_2068);
and U2141 (N_2141,N_2069,N_2074);
nand U2142 (N_2142,N_2055,N_2091);
xnor U2143 (N_2143,N_2076,N_2067);
nand U2144 (N_2144,N_2062,N_2071);
nand U2145 (N_2145,N_2055,N_2077);
nor U2146 (N_2146,N_2086,N_2099);
and U2147 (N_2147,N_2084,N_2086);
nand U2148 (N_2148,N_2046,N_2049);
and U2149 (N_2149,N_2054,N_2047);
nand U2150 (N_2150,N_2042,N_2060);
nor U2151 (N_2151,N_2081,N_2045);
or U2152 (N_2152,N_2092,N_2061);
nand U2153 (N_2153,N_2045,N_2057);
or U2154 (N_2154,N_2066,N_2073);
nand U2155 (N_2155,N_2047,N_2050);
or U2156 (N_2156,N_2080,N_2094);
xor U2157 (N_2157,N_2087,N_2066);
or U2158 (N_2158,N_2067,N_2056);
nor U2159 (N_2159,N_2090,N_2042);
or U2160 (N_2160,N_2154,N_2131);
nand U2161 (N_2161,N_2148,N_2155);
xnor U2162 (N_2162,N_2142,N_2100);
nand U2163 (N_2163,N_2116,N_2127);
and U2164 (N_2164,N_2106,N_2103);
xor U2165 (N_2165,N_2123,N_2130);
and U2166 (N_2166,N_2151,N_2110);
nand U2167 (N_2167,N_2129,N_2115);
nor U2168 (N_2168,N_2125,N_2114);
and U2169 (N_2169,N_2146,N_2128);
xor U2170 (N_2170,N_2135,N_2150);
nand U2171 (N_2171,N_2136,N_2139);
nand U2172 (N_2172,N_2159,N_2144);
nand U2173 (N_2173,N_2117,N_2140);
or U2174 (N_2174,N_2101,N_2111);
nor U2175 (N_2175,N_2137,N_2107);
or U2176 (N_2176,N_2119,N_2138);
and U2177 (N_2177,N_2126,N_2104);
nand U2178 (N_2178,N_2108,N_2118);
and U2179 (N_2179,N_2156,N_2147);
nand U2180 (N_2180,N_2105,N_2112);
or U2181 (N_2181,N_2122,N_2124);
and U2182 (N_2182,N_2149,N_2141);
or U2183 (N_2183,N_2102,N_2120);
or U2184 (N_2184,N_2145,N_2158);
nand U2185 (N_2185,N_2153,N_2132);
nand U2186 (N_2186,N_2134,N_2113);
nor U2187 (N_2187,N_2152,N_2121);
nor U2188 (N_2188,N_2133,N_2157);
nand U2189 (N_2189,N_2109,N_2143);
or U2190 (N_2190,N_2104,N_2112);
or U2191 (N_2191,N_2104,N_2137);
or U2192 (N_2192,N_2135,N_2128);
or U2193 (N_2193,N_2106,N_2126);
nand U2194 (N_2194,N_2159,N_2134);
and U2195 (N_2195,N_2101,N_2119);
or U2196 (N_2196,N_2148,N_2156);
xor U2197 (N_2197,N_2107,N_2151);
or U2198 (N_2198,N_2159,N_2101);
nor U2199 (N_2199,N_2144,N_2140);
xor U2200 (N_2200,N_2150,N_2151);
and U2201 (N_2201,N_2126,N_2112);
and U2202 (N_2202,N_2113,N_2118);
and U2203 (N_2203,N_2154,N_2137);
and U2204 (N_2204,N_2102,N_2107);
and U2205 (N_2205,N_2147,N_2152);
or U2206 (N_2206,N_2139,N_2111);
or U2207 (N_2207,N_2104,N_2132);
nand U2208 (N_2208,N_2147,N_2121);
or U2209 (N_2209,N_2108,N_2137);
nand U2210 (N_2210,N_2156,N_2127);
and U2211 (N_2211,N_2103,N_2148);
nand U2212 (N_2212,N_2138,N_2115);
or U2213 (N_2213,N_2116,N_2121);
nor U2214 (N_2214,N_2141,N_2112);
or U2215 (N_2215,N_2140,N_2128);
or U2216 (N_2216,N_2140,N_2124);
and U2217 (N_2217,N_2116,N_2154);
or U2218 (N_2218,N_2134,N_2136);
nand U2219 (N_2219,N_2158,N_2131);
and U2220 (N_2220,N_2194,N_2201);
nand U2221 (N_2221,N_2184,N_2165);
nor U2222 (N_2222,N_2161,N_2182);
and U2223 (N_2223,N_2213,N_2195);
and U2224 (N_2224,N_2215,N_2198);
nand U2225 (N_2225,N_2200,N_2212);
or U2226 (N_2226,N_2205,N_2203);
or U2227 (N_2227,N_2207,N_2210);
and U2228 (N_2228,N_2173,N_2206);
and U2229 (N_2229,N_2180,N_2190);
nand U2230 (N_2230,N_2187,N_2167);
and U2231 (N_2231,N_2193,N_2181);
xor U2232 (N_2232,N_2197,N_2192);
or U2233 (N_2233,N_2164,N_2162);
and U2234 (N_2234,N_2174,N_2175);
nor U2235 (N_2235,N_2177,N_2218);
and U2236 (N_2236,N_2208,N_2179);
and U2237 (N_2237,N_2199,N_2202);
or U2238 (N_2238,N_2219,N_2183);
nand U2239 (N_2239,N_2172,N_2191);
or U2240 (N_2240,N_2185,N_2166);
xnor U2241 (N_2241,N_2168,N_2196);
or U2242 (N_2242,N_2217,N_2178);
or U2243 (N_2243,N_2169,N_2186);
nand U2244 (N_2244,N_2163,N_2170);
xnor U2245 (N_2245,N_2188,N_2176);
and U2246 (N_2246,N_2214,N_2216);
and U2247 (N_2247,N_2171,N_2209);
nand U2248 (N_2248,N_2189,N_2204);
nor U2249 (N_2249,N_2160,N_2211);
xnor U2250 (N_2250,N_2166,N_2189);
or U2251 (N_2251,N_2183,N_2198);
xor U2252 (N_2252,N_2186,N_2180);
nor U2253 (N_2253,N_2199,N_2204);
nor U2254 (N_2254,N_2209,N_2176);
xor U2255 (N_2255,N_2208,N_2202);
or U2256 (N_2256,N_2161,N_2162);
nor U2257 (N_2257,N_2217,N_2162);
nand U2258 (N_2258,N_2206,N_2188);
and U2259 (N_2259,N_2214,N_2190);
and U2260 (N_2260,N_2176,N_2175);
nor U2261 (N_2261,N_2191,N_2193);
and U2262 (N_2262,N_2195,N_2218);
nor U2263 (N_2263,N_2160,N_2173);
nor U2264 (N_2264,N_2202,N_2182);
nand U2265 (N_2265,N_2173,N_2163);
nor U2266 (N_2266,N_2183,N_2215);
nand U2267 (N_2267,N_2166,N_2209);
nand U2268 (N_2268,N_2161,N_2180);
nand U2269 (N_2269,N_2166,N_2183);
nor U2270 (N_2270,N_2200,N_2181);
or U2271 (N_2271,N_2179,N_2173);
nor U2272 (N_2272,N_2176,N_2214);
or U2273 (N_2273,N_2190,N_2211);
and U2274 (N_2274,N_2180,N_2187);
nor U2275 (N_2275,N_2194,N_2165);
or U2276 (N_2276,N_2192,N_2171);
xnor U2277 (N_2277,N_2213,N_2196);
nor U2278 (N_2278,N_2205,N_2186);
nand U2279 (N_2279,N_2205,N_2214);
nor U2280 (N_2280,N_2228,N_2269);
nand U2281 (N_2281,N_2263,N_2251);
nand U2282 (N_2282,N_2265,N_2227);
nand U2283 (N_2283,N_2247,N_2256);
and U2284 (N_2284,N_2236,N_2229);
or U2285 (N_2285,N_2230,N_2224);
or U2286 (N_2286,N_2246,N_2225);
xor U2287 (N_2287,N_2242,N_2261);
or U2288 (N_2288,N_2276,N_2240);
nor U2289 (N_2289,N_2239,N_2270);
and U2290 (N_2290,N_2254,N_2253);
nor U2291 (N_2291,N_2258,N_2257);
or U2292 (N_2292,N_2275,N_2248);
or U2293 (N_2293,N_2235,N_2278);
and U2294 (N_2294,N_2272,N_2259);
nor U2295 (N_2295,N_2268,N_2232);
or U2296 (N_2296,N_2250,N_2226);
nand U2297 (N_2297,N_2262,N_2244);
nand U2298 (N_2298,N_2231,N_2233);
or U2299 (N_2299,N_2277,N_2249);
or U2300 (N_2300,N_2274,N_2264);
or U2301 (N_2301,N_2234,N_2273);
and U2302 (N_2302,N_2237,N_2267);
and U2303 (N_2303,N_2222,N_2260);
nor U2304 (N_2304,N_2241,N_2245);
nor U2305 (N_2305,N_2221,N_2223);
and U2306 (N_2306,N_2255,N_2266);
and U2307 (N_2307,N_2243,N_2220);
or U2308 (N_2308,N_2238,N_2279);
or U2309 (N_2309,N_2252,N_2271);
nand U2310 (N_2310,N_2257,N_2238);
nor U2311 (N_2311,N_2255,N_2271);
nand U2312 (N_2312,N_2250,N_2265);
or U2313 (N_2313,N_2244,N_2229);
nand U2314 (N_2314,N_2225,N_2257);
or U2315 (N_2315,N_2244,N_2263);
nand U2316 (N_2316,N_2277,N_2256);
and U2317 (N_2317,N_2224,N_2265);
and U2318 (N_2318,N_2259,N_2228);
nor U2319 (N_2319,N_2257,N_2252);
and U2320 (N_2320,N_2262,N_2257);
or U2321 (N_2321,N_2237,N_2231);
nor U2322 (N_2322,N_2253,N_2279);
nor U2323 (N_2323,N_2252,N_2234);
nor U2324 (N_2324,N_2255,N_2248);
nor U2325 (N_2325,N_2275,N_2220);
xnor U2326 (N_2326,N_2257,N_2245);
xnor U2327 (N_2327,N_2264,N_2235);
nor U2328 (N_2328,N_2229,N_2246);
and U2329 (N_2329,N_2248,N_2274);
nor U2330 (N_2330,N_2245,N_2242);
nand U2331 (N_2331,N_2244,N_2246);
nand U2332 (N_2332,N_2274,N_2236);
or U2333 (N_2333,N_2254,N_2276);
or U2334 (N_2334,N_2264,N_2258);
nor U2335 (N_2335,N_2269,N_2255);
xnor U2336 (N_2336,N_2235,N_2257);
and U2337 (N_2337,N_2230,N_2240);
nor U2338 (N_2338,N_2245,N_2237);
or U2339 (N_2339,N_2273,N_2228);
xnor U2340 (N_2340,N_2293,N_2291);
and U2341 (N_2341,N_2320,N_2282);
nor U2342 (N_2342,N_2289,N_2295);
and U2343 (N_2343,N_2331,N_2296);
nor U2344 (N_2344,N_2321,N_2300);
and U2345 (N_2345,N_2317,N_2327);
or U2346 (N_2346,N_2308,N_2284);
and U2347 (N_2347,N_2310,N_2319);
nor U2348 (N_2348,N_2322,N_2339);
or U2349 (N_2349,N_2337,N_2287);
and U2350 (N_2350,N_2285,N_2335);
nor U2351 (N_2351,N_2297,N_2318);
and U2352 (N_2352,N_2336,N_2311);
xor U2353 (N_2353,N_2301,N_2326);
xnor U2354 (N_2354,N_2332,N_2304);
or U2355 (N_2355,N_2329,N_2288);
nor U2356 (N_2356,N_2314,N_2328);
or U2357 (N_2357,N_2323,N_2281);
nor U2358 (N_2358,N_2333,N_2313);
and U2359 (N_2359,N_2330,N_2316);
nand U2360 (N_2360,N_2324,N_2298);
xnor U2361 (N_2361,N_2303,N_2290);
nand U2362 (N_2362,N_2299,N_2283);
xor U2363 (N_2363,N_2307,N_2292);
and U2364 (N_2364,N_2286,N_2338);
nor U2365 (N_2365,N_2312,N_2280);
nor U2366 (N_2366,N_2294,N_2309);
xor U2367 (N_2367,N_2325,N_2305);
xor U2368 (N_2368,N_2302,N_2306);
and U2369 (N_2369,N_2334,N_2315);
nand U2370 (N_2370,N_2301,N_2313);
nand U2371 (N_2371,N_2309,N_2293);
nand U2372 (N_2372,N_2290,N_2329);
and U2373 (N_2373,N_2313,N_2319);
and U2374 (N_2374,N_2320,N_2308);
and U2375 (N_2375,N_2305,N_2308);
nor U2376 (N_2376,N_2337,N_2320);
nor U2377 (N_2377,N_2330,N_2318);
or U2378 (N_2378,N_2321,N_2329);
nand U2379 (N_2379,N_2323,N_2287);
xnor U2380 (N_2380,N_2291,N_2330);
nor U2381 (N_2381,N_2323,N_2325);
or U2382 (N_2382,N_2329,N_2313);
nand U2383 (N_2383,N_2305,N_2301);
and U2384 (N_2384,N_2296,N_2325);
and U2385 (N_2385,N_2311,N_2315);
and U2386 (N_2386,N_2321,N_2320);
nor U2387 (N_2387,N_2313,N_2298);
or U2388 (N_2388,N_2315,N_2295);
nand U2389 (N_2389,N_2333,N_2287);
and U2390 (N_2390,N_2326,N_2282);
nand U2391 (N_2391,N_2335,N_2290);
or U2392 (N_2392,N_2291,N_2298);
xor U2393 (N_2393,N_2321,N_2283);
and U2394 (N_2394,N_2308,N_2299);
and U2395 (N_2395,N_2288,N_2304);
nand U2396 (N_2396,N_2300,N_2308);
xor U2397 (N_2397,N_2297,N_2339);
nor U2398 (N_2398,N_2330,N_2301);
and U2399 (N_2399,N_2306,N_2303);
and U2400 (N_2400,N_2357,N_2399);
and U2401 (N_2401,N_2379,N_2352);
nand U2402 (N_2402,N_2365,N_2366);
xnor U2403 (N_2403,N_2354,N_2393);
and U2404 (N_2404,N_2389,N_2390);
nor U2405 (N_2405,N_2351,N_2343);
nor U2406 (N_2406,N_2381,N_2384);
nand U2407 (N_2407,N_2367,N_2377);
nand U2408 (N_2408,N_2347,N_2342);
and U2409 (N_2409,N_2341,N_2340);
nand U2410 (N_2410,N_2353,N_2383);
or U2411 (N_2411,N_2360,N_2375);
or U2412 (N_2412,N_2382,N_2372);
nand U2413 (N_2413,N_2361,N_2386);
nand U2414 (N_2414,N_2394,N_2395);
or U2415 (N_2415,N_2368,N_2355);
nor U2416 (N_2416,N_2380,N_2345);
or U2417 (N_2417,N_2397,N_2376);
and U2418 (N_2418,N_2359,N_2348);
and U2419 (N_2419,N_2387,N_2370);
and U2420 (N_2420,N_2388,N_2349);
nor U2421 (N_2421,N_2378,N_2398);
or U2422 (N_2422,N_2364,N_2344);
or U2423 (N_2423,N_2371,N_2358);
and U2424 (N_2424,N_2350,N_2392);
or U2425 (N_2425,N_2374,N_2391);
and U2426 (N_2426,N_2396,N_2346);
or U2427 (N_2427,N_2385,N_2362);
nand U2428 (N_2428,N_2373,N_2356);
nand U2429 (N_2429,N_2369,N_2363);
and U2430 (N_2430,N_2394,N_2378);
xnor U2431 (N_2431,N_2352,N_2374);
or U2432 (N_2432,N_2362,N_2397);
nor U2433 (N_2433,N_2384,N_2342);
nand U2434 (N_2434,N_2358,N_2389);
nand U2435 (N_2435,N_2359,N_2349);
and U2436 (N_2436,N_2396,N_2353);
and U2437 (N_2437,N_2397,N_2379);
or U2438 (N_2438,N_2360,N_2354);
or U2439 (N_2439,N_2385,N_2347);
and U2440 (N_2440,N_2363,N_2352);
and U2441 (N_2441,N_2393,N_2343);
and U2442 (N_2442,N_2355,N_2382);
xnor U2443 (N_2443,N_2394,N_2388);
or U2444 (N_2444,N_2374,N_2356);
nand U2445 (N_2445,N_2393,N_2377);
nand U2446 (N_2446,N_2389,N_2372);
and U2447 (N_2447,N_2358,N_2341);
and U2448 (N_2448,N_2364,N_2379);
or U2449 (N_2449,N_2392,N_2378);
nand U2450 (N_2450,N_2360,N_2371);
nor U2451 (N_2451,N_2388,N_2361);
nand U2452 (N_2452,N_2361,N_2369);
nand U2453 (N_2453,N_2375,N_2346);
nand U2454 (N_2454,N_2347,N_2362);
nand U2455 (N_2455,N_2354,N_2387);
or U2456 (N_2456,N_2348,N_2360);
nand U2457 (N_2457,N_2372,N_2398);
xnor U2458 (N_2458,N_2354,N_2369);
nand U2459 (N_2459,N_2352,N_2366);
nand U2460 (N_2460,N_2436,N_2451);
or U2461 (N_2461,N_2432,N_2457);
nor U2462 (N_2462,N_2454,N_2414);
xnor U2463 (N_2463,N_2453,N_2458);
nor U2464 (N_2464,N_2433,N_2448);
and U2465 (N_2465,N_2411,N_2434);
nor U2466 (N_2466,N_2442,N_2417);
or U2467 (N_2467,N_2437,N_2455);
nand U2468 (N_2468,N_2428,N_2450);
or U2469 (N_2469,N_2427,N_2430);
nor U2470 (N_2470,N_2401,N_2459);
xnor U2471 (N_2471,N_2408,N_2400);
or U2472 (N_2472,N_2452,N_2421);
nor U2473 (N_2473,N_2439,N_2456);
nand U2474 (N_2474,N_2415,N_2413);
nor U2475 (N_2475,N_2422,N_2423);
and U2476 (N_2476,N_2420,N_2444);
nand U2477 (N_2477,N_2443,N_2431);
xor U2478 (N_2478,N_2418,N_2405);
nor U2479 (N_2479,N_2404,N_2424);
or U2480 (N_2480,N_2412,N_2449);
xnor U2481 (N_2481,N_2409,N_2416);
nand U2482 (N_2482,N_2402,N_2426);
nand U2483 (N_2483,N_2425,N_2410);
and U2484 (N_2484,N_2440,N_2446);
or U2485 (N_2485,N_2438,N_2406);
or U2486 (N_2486,N_2429,N_2403);
nor U2487 (N_2487,N_2435,N_2419);
nor U2488 (N_2488,N_2445,N_2407);
or U2489 (N_2489,N_2441,N_2447);
and U2490 (N_2490,N_2451,N_2456);
nand U2491 (N_2491,N_2443,N_2407);
and U2492 (N_2492,N_2433,N_2415);
and U2493 (N_2493,N_2431,N_2402);
or U2494 (N_2494,N_2415,N_2420);
xnor U2495 (N_2495,N_2423,N_2424);
and U2496 (N_2496,N_2456,N_2414);
and U2497 (N_2497,N_2444,N_2435);
or U2498 (N_2498,N_2449,N_2400);
xor U2499 (N_2499,N_2403,N_2407);
nor U2500 (N_2500,N_2431,N_2439);
or U2501 (N_2501,N_2442,N_2456);
nor U2502 (N_2502,N_2404,N_2443);
nand U2503 (N_2503,N_2456,N_2411);
and U2504 (N_2504,N_2401,N_2435);
nand U2505 (N_2505,N_2429,N_2421);
and U2506 (N_2506,N_2447,N_2437);
or U2507 (N_2507,N_2459,N_2433);
nand U2508 (N_2508,N_2418,N_2415);
or U2509 (N_2509,N_2405,N_2414);
nand U2510 (N_2510,N_2444,N_2445);
and U2511 (N_2511,N_2438,N_2425);
xor U2512 (N_2512,N_2432,N_2403);
nand U2513 (N_2513,N_2414,N_2453);
nand U2514 (N_2514,N_2454,N_2446);
xor U2515 (N_2515,N_2417,N_2428);
xnor U2516 (N_2516,N_2423,N_2405);
or U2517 (N_2517,N_2408,N_2430);
or U2518 (N_2518,N_2423,N_2446);
and U2519 (N_2519,N_2411,N_2412);
or U2520 (N_2520,N_2503,N_2471);
or U2521 (N_2521,N_2509,N_2491);
or U2522 (N_2522,N_2485,N_2475);
or U2523 (N_2523,N_2497,N_2513);
nor U2524 (N_2524,N_2494,N_2518);
or U2525 (N_2525,N_2469,N_2473);
nand U2526 (N_2526,N_2508,N_2488);
and U2527 (N_2527,N_2492,N_2490);
or U2528 (N_2528,N_2504,N_2510);
nand U2529 (N_2529,N_2479,N_2499);
nor U2530 (N_2530,N_2487,N_2496);
nand U2531 (N_2531,N_2461,N_2498);
or U2532 (N_2532,N_2517,N_2468);
xor U2533 (N_2533,N_2462,N_2495);
nand U2534 (N_2534,N_2477,N_2505);
xor U2535 (N_2535,N_2511,N_2516);
nand U2536 (N_2536,N_2486,N_2502);
nand U2537 (N_2537,N_2472,N_2466);
and U2538 (N_2538,N_2515,N_2467);
nor U2539 (N_2539,N_2460,N_2474);
and U2540 (N_2540,N_2478,N_2501);
and U2541 (N_2541,N_2463,N_2476);
or U2542 (N_2542,N_2481,N_2483);
xnor U2543 (N_2543,N_2465,N_2519);
nand U2544 (N_2544,N_2500,N_2506);
nor U2545 (N_2545,N_2470,N_2484);
and U2546 (N_2546,N_2480,N_2512);
and U2547 (N_2547,N_2507,N_2489);
xnor U2548 (N_2548,N_2493,N_2464);
and U2549 (N_2549,N_2482,N_2514);
or U2550 (N_2550,N_2501,N_2482);
or U2551 (N_2551,N_2462,N_2468);
or U2552 (N_2552,N_2504,N_2499);
or U2553 (N_2553,N_2504,N_2517);
nand U2554 (N_2554,N_2476,N_2494);
nor U2555 (N_2555,N_2515,N_2503);
or U2556 (N_2556,N_2476,N_2464);
nand U2557 (N_2557,N_2490,N_2486);
or U2558 (N_2558,N_2477,N_2481);
nor U2559 (N_2559,N_2463,N_2489);
or U2560 (N_2560,N_2511,N_2487);
nand U2561 (N_2561,N_2482,N_2475);
and U2562 (N_2562,N_2507,N_2514);
or U2563 (N_2563,N_2518,N_2478);
nor U2564 (N_2564,N_2493,N_2473);
nor U2565 (N_2565,N_2496,N_2499);
or U2566 (N_2566,N_2511,N_2463);
or U2567 (N_2567,N_2494,N_2491);
nor U2568 (N_2568,N_2507,N_2481);
or U2569 (N_2569,N_2484,N_2499);
nand U2570 (N_2570,N_2486,N_2470);
or U2571 (N_2571,N_2518,N_2489);
nand U2572 (N_2572,N_2478,N_2507);
nand U2573 (N_2573,N_2498,N_2515);
and U2574 (N_2574,N_2485,N_2503);
nand U2575 (N_2575,N_2509,N_2514);
or U2576 (N_2576,N_2491,N_2506);
or U2577 (N_2577,N_2474,N_2504);
nand U2578 (N_2578,N_2480,N_2511);
nor U2579 (N_2579,N_2500,N_2515);
nand U2580 (N_2580,N_2574,N_2553);
nor U2581 (N_2581,N_2559,N_2537);
nor U2582 (N_2582,N_2530,N_2568);
or U2583 (N_2583,N_2523,N_2547);
or U2584 (N_2584,N_2577,N_2536);
and U2585 (N_2585,N_2543,N_2551);
or U2586 (N_2586,N_2550,N_2570);
nand U2587 (N_2587,N_2531,N_2549);
and U2588 (N_2588,N_2557,N_2548);
xnor U2589 (N_2589,N_2524,N_2535);
and U2590 (N_2590,N_2562,N_2555);
xor U2591 (N_2591,N_2563,N_2522);
nand U2592 (N_2592,N_2527,N_2541);
and U2593 (N_2593,N_2539,N_2569);
nand U2594 (N_2594,N_2532,N_2521);
nor U2595 (N_2595,N_2565,N_2579);
nand U2596 (N_2596,N_2533,N_2566);
nand U2597 (N_2597,N_2571,N_2520);
or U2598 (N_2598,N_2526,N_2538);
nand U2599 (N_2599,N_2573,N_2578);
or U2600 (N_2600,N_2552,N_2558);
nand U2601 (N_2601,N_2564,N_2554);
nor U2602 (N_2602,N_2576,N_2560);
nand U2603 (N_2603,N_2534,N_2528);
nand U2604 (N_2604,N_2529,N_2575);
nor U2605 (N_2605,N_2542,N_2525);
nor U2606 (N_2606,N_2572,N_2567);
or U2607 (N_2607,N_2546,N_2561);
nand U2608 (N_2608,N_2544,N_2545);
nor U2609 (N_2609,N_2556,N_2540);
nor U2610 (N_2610,N_2533,N_2576);
nand U2611 (N_2611,N_2524,N_2567);
or U2612 (N_2612,N_2561,N_2544);
nand U2613 (N_2613,N_2543,N_2545);
or U2614 (N_2614,N_2564,N_2573);
or U2615 (N_2615,N_2550,N_2573);
or U2616 (N_2616,N_2574,N_2529);
nand U2617 (N_2617,N_2522,N_2552);
nor U2618 (N_2618,N_2551,N_2523);
nor U2619 (N_2619,N_2535,N_2570);
and U2620 (N_2620,N_2537,N_2524);
nand U2621 (N_2621,N_2520,N_2553);
and U2622 (N_2622,N_2550,N_2527);
nor U2623 (N_2623,N_2536,N_2560);
xnor U2624 (N_2624,N_2537,N_2530);
or U2625 (N_2625,N_2551,N_2553);
nand U2626 (N_2626,N_2571,N_2563);
and U2627 (N_2627,N_2548,N_2576);
xor U2628 (N_2628,N_2541,N_2535);
or U2629 (N_2629,N_2554,N_2529);
and U2630 (N_2630,N_2546,N_2577);
or U2631 (N_2631,N_2566,N_2536);
or U2632 (N_2632,N_2542,N_2557);
and U2633 (N_2633,N_2552,N_2521);
or U2634 (N_2634,N_2525,N_2561);
and U2635 (N_2635,N_2564,N_2548);
nand U2636 (N_2636,N_2562,N_2522);
or U2637 (N_2637,N_2577,N_2535);
nor U2638 (N_2638,N_2560,N_2550);
nor U2639 (N_2639,N_2555,N_2547);
or U2640 (N_2640,N_2583,N_2616);
and U2641 (N_2641,N_2632,N_2625);
or U2642 (N_2642,N_2634,N_2614);
xnor U2643 (N_2643,N_2626,N_2596);
nand U2644 (N_2644,N_2620,N_2612);
xor U2645 (N_2645,N_2585,N_2601);
and U2646 (N_2646,N_2619,N_2624);
nor U2647 (N_2647,N_2635,N_2627);
xnor U2648 (N_2648,N_2591,N_2608);
nor U2649 (N_2649,N_2630,N_2581);
and U2650 (N_2650,N_2602,N_2582);
and U2651 (N_2651,N_2609,N_2586);
xnor U2652 (N_2652,N_2584,N_2603);
nor U2653 (N_2653,N_2606,N_2607);
nand U2654 (N_2654,N_2622,N_2617);
or U2655 (N_2655,N_2631,N_2633);
and U2656 (N_2656,N_2638,N_2618);
or U2657 (N_2657,N_2595,N_2613);
and U2658 (N_2658,N_2594,N_2598);
nand U2659 (N_2659,N_2628,N_2611);
nand U2660 (N_2660,N_2636,N_2589);
and U2661 (N_2661,N_2599,N_2580);
or U2662 (N_2662,N_2621,N_2597);
nand U2663 (N_2663,N_2615,N_2593);
or U2664 (N_2664,N_2605,N_2637);
and U2665 (N_2665,N_2639,N_2604);
nand U2666 (N_2666,N_2600,N_2629);
xnor U2667 (N_2667,N_2623,N_2592);
nor U2668 (N_2668,N_2588,N_2587);
nand U2669 (N_2669,N_2610,N_2590);
or U2670 (N_2670,N_2608,N_2636);
nor U2671 (N_2671,N_2603,N_2639);
nand U2672 (N_2672,N_2592,N_2636);
nand U2673 (N_2673,N_2593,N_2610);
and U2674 (N_2674,N_2614,N_2608);
and U2675 (N_2675,N_2616,N_2585);
or U2676 (N_2676,N_2638,N_2633);
nor U2677 (N_2677,N_2621,N_2598);
nor U2678 (N_2678,N_2638,N_2600);
and U2679 (N_2679,N_2620,N_2592);
nand U2680 (N_2680,N_2604,N_2583);
xnor U2681 (N_2681,N_2588,N_2607);
nand U2682 (N_2682,N_2596,N_2586);
or U2683 (N_2683,N_2617,N_2593);
xnor U2684 (N_2684,N_2612,N_2586);
nor U2685 (N_2685,N_2599,N_2597);
or U2686 (N_2686,N_2625,N_2582);
nand U2687 (N_2687,N_2620,N_2582);
nor U2688 (N_2688,N_2599,N_2601);
xor U2689 (N_2689,N_2616,N_2620);
nor U2690 (N_2690,N_2613,N_2612);
nor U2691 (N_2691,N_2588,N_2627);
nand U2692 (N_2692,N_2619,N_2585);
nand U2693 (N_2693,N_2585,N_2604);
or U2694 (N_2694,N_2601,N_2613);
xnor U2695 (N_2695,N_2582,N_2619);
nor U2696 (N_2696,N_2598,N_2614);
nor U2697 (N_2697,N_2592,N_2594);
xnor U2698 (N_2698,N_2598,N_2624);
and U2699 (N_2699,N_2584,N_2626);
or U2700 (N_2700,N_2693,N_2646);
or U2701 (N_2701,N_2695,N_2689);
and U2702 (N_2702,N_2641,N_2643);
xor U2703 (N_2703,N_2677,N_2662);
nor U2704 (N_2704,N_2681,N_2655);
nand U2705 (N_2705,N_2674,N_2667);
xor U2706 (N_2706,N_2668,N_2664);
nand U2707 (N_2707,N_2675,N_2658);
or U2708 (N_2708,N_2673,N_2644);
or U2709 (N_2709,N_2642,N_2651);
nor U2710 (N_2710,N_2640,N_2680);
nor U2711 (N_2711,N_2650,N_2649);
nor U2712 (N_2712,N_2694,N_2661);
and U2713 (N_2713,N_2648,N_2670);
and U2714 (N_2714,N_2688,N_2665);
nor U2715 (N_2715,N_2686,N_2663);
nor U2716 (N_2716,N_2653,N_2678);
or U2717 (N_2717,N_2699,N_2697);
and U2718 (N_2718,N_2659,N_2696);
nand U2719 (N_2719,N_2690,N_2660);
nand U2720 (N_2720,N_2676,N_2652);
and U2721 (N_2721,N_2684,N_2669);
and U2722 (N_2722,N_2672,N_2698);
nor U2723 (N_2723,N_2656,N_2685);
or U2724 (N_2724,N_2647,N_2645);
nand U2725 (N_2725,N_2682,N_2679);
nand U2726 (N_2726,N_2687,N_2683);
xnor U2727 (N_2727,N_2692,N_2654);
nor U2728 (N_2728,N_2671,N_2666);
nand U2729 (N_2729,N_2657,N_2691);
and U2730 (N_2730,N_2692,N_2684);
and U2731 (N_2731,N_2691,N_2655);
nand U2732 (N_2732,N_2640,N_2681);
or U2733 (N_2733,N_2673,N_2667);
or U2734 (N_2734,N_2689,N_2661);
and U2735 (N_2735,N_2672,N_2640);
nor U2736 (N_2736,N_2691,N_2662);
xnor U2737 (N_2737,N_2696,N_2661);
xnor U2738 (N_2738,N_2647,N_2682);
or U2739 (N_2739,N_2687,N_2664);
nor U2740 (N_2740,N_2649,N_2676);
nor U2741 (N_2741,N_2693,N_2673);
nor U2742 (N_2742,N_2690,N_2670);
nand U2743 (N_2743,N_2696,N_2664);
or U2744 (N_2744,N_2644,N_2692);
and U2745 (N_2745,N_2670,N_2643);
or U2746 (N_2746,N_2692,N_2672);
or U2747 (N_2747,N_2691,N_2698);
and U2748 (N_2748,N_2670,N_2655);
xnor U2749 (N_2749,N_2685,N_2667);
and U2750 (N_2750,N_2685,N_2679);
nand U2751 (N_2751,N_2655,N_2697);
or U2752 (N_2752,N_2659,N_2655);
nand U2753 (N_2753,N_2640,N_2654);
nand U2754 (N_2754,N_2699,N_2684);
nor U2755 (N_2755,N_2674,N_2675);
and U2756 (N_2756,N_2679,N_2653);
or U2757 (N_2757,N_2691,N_2645);
and U2758 (N_2758,N_2665,N_2661);
or U2759 (N_2759,N_2646,N_2643);
nor U2760 (N_2760,N_2751,N_2744);
nor U2761 (N_2761,N_2758,N_2721);
and U2762 (N_2762,N_2705,N_2703);
or U2763 (N_2763,N_2740,N_2746);
nor U2764 (N_2764,N_2755,N_2700);
nor U2765 (N_2765,N_2726,N_2757);
nand U2766 (N_2766,N_2747,N_2716);
xnor U2767 (N_2767,N_2712,N_2714);
nand U2768 (N_2768,N_2736,N_2733);
or U2769 (N_2769,N_2731,N_2715);
or U2770 (N_2770,N_2725,N_2732);
or U2771 (N_2771,N_2708,N_2730);
and U2772 (N_2772,N_2741,N_2748);
nand U2773 (N_2773,N_2734,N_2759);
and U2774 (N_2774,N_2711,N_2723);
xor U2775 (N_2775,N_2752,N_2717);
and U2776 (N_2776,N_2743,N_2724);
and U2777 (N_2777,N_2735,N_2713);
nor U2778 (N_2778,N_2719,N_2722);
nand U2779 (N_2779,N_2737,N_2739);
nor U2780 (N_2780,N_2709,N_2745);
or U2781 (N_2781,N_2749,N_2701);
and U2782 (N_2782,N_2710,N_2756);
and U2783 (N_2783,N_2706,N_2754);
nor U2784 (N_2784,N_2750,N_2727);
nand U2785 (N_2785,N_2729,N_2720);
xor U2786 (N_2786,N_2753,N_2738);
nor U2787 (N_2787,N_2728,N_2702);
and U2788 (N_2788,N_2718,N_2707);
or U2789 (N_2789,N_2704,N_2742);
nand U2790 (N_2790,N_2749,N_2714);
nor U2791 (N_2791,N_2741,N_2736);
and U2792 (N_2792,N_2708,N_2735);
xor U2793 (N_2793,N_2736,N_2711);
and U2794 (N_2794,N_2712,N_2752);
or U2795 (N_2795,N_2740,N_2700);
nand U2796 (N_2796,N_2731,N_2723);
and U2797 (N_2797,N_2733,N_2725);
or U2798 (N_2798,N_2758,N_2733);
or U2799 (N_2799,N_2740,N_2704);
nor U2800 (N_2800,N_2746,N_2754);
or U2801 (N_2801,N_2706,N_2725);
and U2802 (N_2802,N_2759,N_2717);
or U2803 (N_2803,N_2746,N_2715);
or U2804 (N_2804,N_2740,N_2713);
nor U2805 (N_2805,N_2722,N_2734);
and U2806 (N_2806,N_2744,N_2757);
nor U2807 (N_2807,N_2759,N_2711);
and U2808 (N_2808,N_2742,N_2759);
nor U2809 (N_2809,N_2741,N_2729);
nor U2810 (N_2810,N_2712,N_2704);
nand U2811 (N_2811,N_2703,N_2740);
or U2812 (N_2812,N_2737,N_2757);
or U2813 (N_2813,N_2751,N_2718);
nor U2814 (N_2814,N_2705,N_2750);
nor U2815 (N_2815,N_2711,N_2742);
nor U2816 (N_2816,N_2730,N_2726);
nor U2817 (N_2817,N_2756,N_2736);
nand U2818 (N_2818,N_2702,N_2754);
and U2819 (N_2819,N_2752,N_2706);
nor U2820 (N_2820,N_2778,N_2775);
xnor U2821 (N_2821,N_2797,N_2802);
or U2822 (N_2822,N_2806,N_2788);
nand U2823 (N_2823,N_2817,N_2804);
and U2824 (N_2824,N_2809,N_2780);
nand U2825 (N_2825,N_2807,N_2794);
nor U2826 (N_2826,N_2767,N_2761);
xor U2827 (N_2827,N_2782,N_2812);
or U2828 (N_2828,N_2811,N_2810);
nand U2829 (N_2829,N_2770,N_2771);
nor U2830 (N_2830,N_2808,N_2800);
nand U2831 (N_2831,N_2814,N_2777);
and U2832 (N_2832,N_2774,N_2764);
xnor U2833 (N_2833,N_2765,N_2762);
nand U2834 (N_2834,N_2787,N_2789);
nand U2835 (N_2835,N_2813,N_2773);
xor U2836 (N_2836,N_2763,N_2816);
nand U2837 (N_2837,N_2779,N_2818);
or U2838 (N_2838,N_2785,N_2790);
nor U2839 (N_2839,N_2805,N_2798);
nand U2840 (N_2840,N_2781,N_2793);
or U2841 (N_2841,N_2760,N_2815);
and U2842 (N_2842,N_2799,N_2768);
nand U2843 (N_2843,N_2776,N_2783);
or U2844 (N_2844,N_2791,N_2766);
and U2845 (N_2845,N_2819,N_2801);
nor U2846 (N_2846,N_2786,N_2792);
nand U2847 (N_2847,N_2796,N_2803);
and U2848 (N_2848,N_2795,N_2784);
and U2849 (N_2849,N_2772,N_2769);
nand U2850 (N_2850,N_2779,N_2791);
or U2851 (N_2851,N_2809,N_2777);
nand U2852 (N_2852,N_2781,N_2819);
and U2853 (N_2853,N_2771,N_2802);
nand U2854 (N_2854,N_2812,N_2780);
and U2855 (N_2855,N_2808,N_2766);
and U2856 (N_2856,N_2791,N_2764);
nor U2857 (N_2857,N_2798,N_2803);
nand U2858 (N_2858,N_2797,N_2780);
and U2859 (N_2859,N_2802,N_2781);
xnor U2860 (N_2860,N_2811,N_2794);
nand U2861 (N_2861,N_2808,N_2813);
nand U2862 (N_2862,N_2783,N_2764);
nand U2863 (N_2863,N_2783,N_2775);
nor U2864 (N_2864,N_2801,N_2807);
nand U2865 (N_2865,N_2785,N_2806);
nand U2866 (N_2866,N_2809,N_2781);
or U2867 (N_2867,N_2803,N_2762);
nor U2868 (N_2868,N_2760,N_2795);
and U2869 (N_2869,N_2784,N_2767);
nor U2870 (N_2870,N_2774,N_2771);
or U2871 (N_2871,N_2799,N_2780);
or U2872 (N_2872,N_2801,N_2792);
and U2873 (N_2873,N_2802,N_2816);
nor U2874 (N_2874,N_2766,N_2793);
nor U2875 (N_2875,N_2816,N_2793);
and U2876 (N_2876,N_2775,N_2788);
or U2877 (N_2877,N_2776,N_2760);
and U2878 (N_2878,N_2806,N_2765);
nand U2879 (N_2879,N_2805,N_2765);
xnor U2880 (N_2880,N_2822,N_2837);
or U2881 (N_2881,N_2872,N_2849);
xnor U2882 (N_2882,N_2853,N_2842);
nor U2883 (N_2883,N_2867,N_2829);
and U2884 (N_2884,N_2836,N_2823);
nand U2885 (N_2885,N_2877,N_2863);
and U2886 (N_2886,N_2856,N_2868);
and U2887 (N_2887,N_2848,N_2846);
xnor U2888 (N_2888,N_2879,N_2865);
nand U2889 (N_2889,N_2831,N_2860);
and U2890 (N_2890,N_2861,N_2852);
nor U2891 (N_2891,N_2878,N_2838);
or U2892 (N_2892,N_2828,N_2876);
or U2893 (N_2893,N_2843,N_2871);
nor U2894 (N_2894,N_2873,N_2866);
and U2895 (N_2895,N_2858,N_2820);
nand U2896 (N_2896,N_2875,N_2825);
nand U2897 (N_2897,N_2832,N_2826);
and U2898 (N_2898,N_2827,N_2862);
nor U2899 (N_2899,N_2839,N_2855);
or U2900 (N_2900,N_2824,N_2830);
and U2901 (N_2901,N_2851,N_2857);
nand U2902 (N_2902,N_2869,N_2850);
or U2903 (N_2903,N_2844,N_2859);
or U2904 (N_2904,N_2847,N_2870);
xnor U2905 (N_2905,N_2845,N_2864);
nand U2906 (N_2906,N_2821,N_2874);
nor U2907 (N_2907,N_2835,N_2833);
nand U2908 (N_2908,N_2834,N_2854);
nand U2909 (N_2909,N_2840,N_2841);
nor U2910 (N_2910,N_2868,N_2839);
or U2911 (N_2911,N_2845,N_2823);
nand U2912 (N_2912,N_2834,N_2866);
and U2913 (N_2913,N_2830,N_2834);
nor U2914 (N_2914,N_2846,N_2824);
and U2915 (N_2915,N_2859,N_2873);
nor U2916 (N_2916,N_2861,N_2831);
and U2917 (N_2917,N_2836,N_2844);
nor U2918 (N_2918,N_2823,N_2833);
or U2919 (N_2919,N_2825,N_2848);
or U2920 (N_2920,N_2878,N_2879);
nor U2921 (N_2921,N_2857,N_2836);
xnor U2922 (N_2922,N_2827,N_2840);
nor U2923 (N_2923,N_2860,N_2849);
xor U2924 (N_2924,N_2830,N_2833);
nor U2925 (N_2925,N_2849,N_2858);
nor U2926 (N_2926,N_2868,N_2850);
nand U2927 (N_2927,N_2841,N_2834);
or U2928 (N_2928,N_2835,N_2854);
nand U2929 (N_2929,N_2833,N_2824);
nor U2930 (N_2930,N_2849,N_2833);
or U2931 (N_2931,N_2829,N_2863);
and U2932 (N_2932,N_2855,N_2865);
and U2933 (N_2933,N_2872,N_2845);
nor U2934 (N_2934,N_2860,N_2876);
nand U2935 (N_2935,N_2827,N_2830);
or U2936 (N_2936,N_2857,N_2835);
nand U2937 (N_2937,N_2857,N_2876);
xor U2938 (N_2938,N_2820,N_2825);
nor U2939 (N_2939,N_2844,N_2840);
or U2940 (N_2940,N_2930,N_2883);
and U2941 (N_2941,N_2922,N_2901);
nor U2942 (N_2942,N_2912,N_2929);
nand U2943 (N_2943,N_2925,N_2928);
nand U2944 (N_2944,N_2884,N_2916);
xnor U2945 (N_2945,N_2937,N_2935);
nand U2946 (N_2946,N_2933,N_2895);
nor U2947 (N_2947,N_2911,N_2924);
and U2948 (N_2948,N_2905,N_2891);
nand U2949 (N_2949,N_2939,N_2906);
xor U2950 (N_2950,N_2923,N_2896);
nand U2951 (N_2951,N_2921,N_2913);
nor U2952 (N_2952,N_2934,N_2885);
nand U2953 (N_2953,N_2882,N_2917);
nor U2954 (N_2954,N_2888,N_2907);
or U2955 (N_2955,N_2931,N_2914);
or U2956 (N_2956,N_2920,N_2881);
nand U2957 (N_2957,N_2900,N_2902);
or U2958 (N_2958,N_2938,N_2919);
nand U2959 (N_2959,N_2894,N_2889);
nor U2960 (N_2960,N_2880,N_2897);
or U2961 (N_2961,N_2915,N_2892);
nor U2962 (N_2962,N_2926,N_2898);
and U2963 (N_2963,N_2903,N_2887);
nor U2964 (N_2964,N_2899,N_2890);
nand U2965 (N_2965,N_2936,N_2918);
and U2966 (N_2966,N_2909,N_2910);
xor U2967 (N_2967,N_2904,N_2927);
nor U2968 (N_2968,N_2893,N_2908);
or U2969 (N_2969,N_2932,N_2886);
nor U2970 (N_2970,N_2918,N_2930);
or U2971 (N_2971,N_2885,N_2899);
nor U2972 (N_2972,N_2895,N_2911);
nand U2973 (N_2973,N_2907,N_2900);
and U2974 (N_2974,N_2896,N_2895);
xor U2975 (N_2975,N_2933,N_2919);
and U2976 (N_2976,N_2896,N_2904);
and U2977 (N_2977,N_2920,N_2882);
nor U2978 (N_2978,N_2888,N_2926);
xor U2979 (N_2979,N_2915,N_2938);
and U2980 (N_2980,N_2929,N_2932);
nand U2981 (N_2981,N_2919,N_2917);
nor U2982 (N_2982,N_2939,N_2916);
nor U2983 (N_2983,N_2921,N_2928);
and U2984 (N_2984,N_2927,N_2899);
nand U2985 (N_2985,N_2903,N_2922);
or U2986 (N_2986,N_2906,N_2913);
nand U2987 (N_2987,N_2885,N_2919);
and U2988 (N_2988,N_2922,N_2936);
or U2989 (N_2989,N_2889,N_2936);
xor U2990 (N_2990,N_2910,N_2884);
or U2991 (N_2991,N_2903,N_2904);
nand U2992 (N_2992,N_2887,N_2886);
or U2993 (N_2993,N_2920,N_2880);
and U2994 (N_2994,N_2901,N_2929);
nor U2995 (N_2995,N_2919,N_2883);
nand U2996 (N_2996,N_2924,N_2899);
and U2997 (N_2997,N_2890,N_2934);
nand U2998 (N_2998,N_2927,N_2920);
and U2999 (N_2999,N_2930,N_2925);
nand UO_0 (O_0,N_2950,N_2953);
nor UO_1 (O_1,N_2949,N_2985);
or UO_2 (O_2,N_2986,N_2961);
nor UO_3 (O_3,N_2982,N_2979);
nor UO_4 (O_4,N_2992,N_2998);
nor UO_5 (O_5,N_2997,N_2968);
nand UO_6 (O_6,N_2942,N_2999);
nand UO_7 (O_7,N_2940,N_2943);
nor UO_8 (O_8,N_2994,N_2973);
and UO_9 (O_9,N_2981,N_2988);
nor UO_10 (O_10,N_2990,N_2974);
nor UO_11 (O_11,N_2956,N_2957);
or UO_12 (O_12,N_2960,N_2947);
and UO_13 (O_13,N_2996,N_2955);
xor UO_14 (O_14,N_2983,N_2970);
nor UO_15 (O_15,N_2972,N_2975);
and UO_16 (O_16,N_2984,N_2995);
nor UO_17 (O_17,N_2944,N_2966);
and UO_18 (O_18,N_2980,N_2952);
nand UO_19 (O_19,N_2965,N_2969);
and UO_20 (O_20,N_2958,N_2959);
or UO_21 (O_21,N_2962,N_2967);
xor UO_22 (O_22,N_2978,N_2954);
and UO_23 (O_23,N_2971,N_2987);
or UO_24 (O_24,N_2964,N_2946);
and UO_25 (O_25,N_2977,N_2951);
or UO_26 (O_26,N_2989,N_2991);
nand UO_27 (O_27,N_2941,N_2945);
nor UO_28 (O_28,N_2976,N_2993);
or UO_29 (O_29,N_2963,N_2948);
nor UO_30 (O_30,N_2976,N_2989);
xnor UO_31 (O_31,N_2993,N_2981);
nor UO_32 (O_32,N_2948,N_2992);
nand UO_33 (O_33,N_2952,N_2990);
and UO_34 (O_34,N_2993,N_2978);
xnor UO_35 (O_35,N_2973,N_2959);
nor UO_36 (O_36,N_2956,N_2965);
nor UO_37 (O_37,N_2949,N_2943);
xnor UO_38 (O_38,N_2976,N_2958);
or UO_39 (O_39,N_2993,N_2949);
nand UO_40 (O_40,N_2942,N_2985);
and UO_41 (O_41,N_2986,N_2995);
xor UO_42 (O_42,N_2978,N_2952);
nor UO_43 (O_43,N_2944,N_2965);
xor UO_44 (O_44,N_2962,N_2954);
and UO_45 (O_45,N_2959,N_2991);
nor UO_46 (O_46,N_2986,N_2999);
nand UO_47 (O_47,N_2963,N_2986);
and UO_48 (O_48,N_2957,N_2994);
nand UO_49 (O_49,N_2979,N_2970);
nand UO_50 (O_50,N_2958,N_2991);
and UO_51 (O_51,N_2990,N_2987);
nor UO_52 (O_52,N_2971,N_2995);
and UO_53 (O_53,N_2961,N_2973);
or UO_54 (O_54,N_2999,N_2988);
and UO_55 (O_55,N_2992,N_2951);
nand UO_56 (O_56,N_2944,N_2949);
and UO_57 (O_57,N_2971,N_2964);
nand UO_58 (O_58,N_2968,N_2985);
nand UO_59 (O_59,N_2987,N_2956);
or UO_60 (O_60,N_2954,N_2995);
nor UO_61 (O_61,N_2977,N_2948);
and UO_62 (O_62,N_2991,N_2992);
nand UO_63 (O_63,N_2956,N_2992);
and UO_64 (O_64,N_2966,N_2995);
or UO_65 (O_65,N_2961,N_2982);
and UO_66 (O_66,N_2993,N_2972);
and UO_67 (O_67,N_2991,N_2956);
nand UO_68 (O_68,N_2950,N_2947);
or UO_69 (O_69,N_2992,N_2995);
nor UO_70 (O_70,N_2997,N_2985);
nand UO_71 (O_71,N_2959,N_2979);
or UO_72 (O_72,N_2988,N_2959);
and UO_73 (O_73,N_2956,N_2998);
and UO_74 (O_74,N_2969,N_2964);
nor UO_75 (O_75,N_2997,N_2982);
nor UO_76 (O_76,N_2946,N_2973);
xor UO_77 (O_77,N_2990,N_2983);
and UO_78 (O_78,N_2967,N_2940);
and UO_79 (O_79,N_2966,N_2985);
or UO_80 (O_80,N_2996,N_2989);
nand UO_81 (O_81,N_2963,N_2985);
or UO_82 (O_82,N_2959,N_2961);
nand UO_83 (O_83,N_2972,N_2947);
and UO_84 (O_84,N_2972,N_2963);
nor UO_85 (O_85,N_2957,N_2976);
or UO_86 (O_86,N_2974,N_2941);
nor UO_87 (O_87,N_2952,N_2976);
xor UO_88 (O_88,N_2975,N_2970);
nor UO_89 (O_89,N_2969,N_2998);
xor UO_90 (O_90,N_2970,N_2956);
nand UO_91 (O_91,N_2998,N_2993);
and UO_92 (O_92,N_2960,N_2946);
or UO_93 (O_93,N_2954,N_2961);
xnor UO_94 (O_94,N_2949,N_2995);
or UO_95 (O_95,N_2956,N_2994);
nor UO_96 (O_96,N_2950,N_2986);
nor UO_97 (O_97,N_2990,N_2946);
and UO_98 (O_98,N_2989,N_2967);
and UO_99 (O_99,N_2958,N_2950);
nand UO_100 (O_100,N_2945,N_2947);
and UO_101 (O_101,N_2959,N_2945);
nand UO_102 (O_102,N_2979,N_2983);
or UO_103 (O_103,N_2957,N_2984);
nand UO_104 (O_104,N_2987,N_2994);
xor UO_105 (O_105,N_2952,N_2989);
or UO_106 (O_106,N_2977,N_2958);
or UO_107 (O_107,N_2971,N_2965);
or UO_108 (O_108,N_2942,N_2992);
or UO_109 (O_109,N_2963,N_2949);
nor UO_110 (O_110,N_2946,N_2995);
nand UO_111 (O_111,N_2949,N_2971);
xor UO_112 (O_112,N_2981,N_2980);
or UO_113 (O_113,N_2965,N_2952);
or UO_114 (O_114,N_2971,N_2966);
or UO_115 (O_115,N_2971,N_2985);
xnor UO_116 (O_116,N_2972,N_2954);
or UO_117 (O_117,N_2963,N_2980);
or UO_118 (O_118,N_2955,N_2972);
or UO_119 (O_119,N_2990,N_2998);
nor UO_120 (O_120,N_2940,N_2964);
and UO_121 (O_121,N_2994,N_2959);
xnor UO_122 (O_122,N_2959,N_2993);
xnor UO_123 (O_123,N_2967,N_2948);
and UO_124 (O_124,N_2976,N_2985);
and UO_125 (O_125,N_2974,N_2972);
nand UO_126 (O_126,N_2943,N_2946);
nor UO_127 (O_127,N_2952,N_2969);
or UO_128 (O_128,N_2997,N_2965);
nor UO_129 (O_129,N_2962,N_2981);
xnor UO_130 (O_130,N_2954,N_2998);
nand UO_131 (O_131,N_2985,N_2984);
nor UO_132 (O_132,N_2968,N_2952);
nand UO_133 (O_133,N_2957,N_2963);
nand UO_134 (O_134,N_2991,N_2970);
nand UO_135 (O_135,N_2942,N_2959);
nor UO_136 (O_136,N_2991,N_2964);
and UO_137 (O_137,N_2995,N_2945);
or UO_138 (O_138,N_2964,N_2955);
nor UO_139 (O_139,N_2994,N_2949);
nor UO_140 (O_140,N_2979,N_2996);
or UO_141 (O_141,N_2965,N_2974);
or UO_142 (O_142,N_2993,N_2967);
and UO_143 (O_143,N_2954,N_2964);
nor UO_144 (O_144,N_2970,N_2994);
and UO_145 (O_145,N_2951,N_2964);
or UO_146 (O_146,N_2966,N_2959);
nand UO_147 (O_147,N_2994,N_2955);
nand UO_148 (O_148,N_2964,N_2973);
nor UO_149 (O_149,N_2966,N_2947);
nor UO_150 (O_150,N_2994,N_2969);
or UO_151 (O_151,N_2988,N_2977);
or UO_152 (O_152,N_2993,N_2964);
nand UO_153 (O_153,N_2941,N_2977);
nand UO_154 (O_154,N_2978,N_2989);
nor UO_155 (O_155,N_2942,N_2996);
and UO_156 (O_156,N_2969,N_2980);
nor UO_157 (O_157,N_2952,N_2958);
nor UO_158 (O_158,N_2968,N_2944);
or UO_159 (O_159,N_2984,N_2946);
nand UO_160 (O_160,N_2986,N_2970);
or UO_161 (O_161,N_2982,N_2995);
or UO_162 (O_162,N_2950,N_2985);
and UO_163 (O_163,N_2946,N_2953);
nand UO_164 (O_164,N_2962,N_2998);
or UO_165 (O_165,N_2968,N_2941);
or UO_166 (O_166,N_2994,N_2964);
xor UO_167 (O_167,N_2973,N_2981);
and UO_168 (O_168,N_2986,N_2944);
nor UO_169 (O_169,N_2968,N_2950);
nand UO_170 (O_170,N_2982,N_2999);
xor UO_171 (O_171,N_2979,N_2957);
xnor UO_172 (O_172,N_2997,N_2996);
and UO_173 (O_173,N_2940,N_2970);
nand UO_174 (O_174,N_2951,N_2944);
or UO_175 (O_175,N_2963,N_2966);
or UO_176 (O_176,N_2967,N_2977);
and UO_177 (O_177,N_2995,N_2961);
nor UO_178 (O_178,N_2940,N_2976);
and UO_179 (O_179,N_2984,N_2979);
and UO_180 (O_180,N_2975,N_2985);
nand UO_181 (O_181,N_2975,N_2991);
or UO_182 (O_182,N_2941,N_2979);
nand UO_183 (O_183,N_2941,N_2962);
and UO_184 (O_184,N_2997,N_2963);
xnor UO_185 (O_185,N_2974,N_2977);
nand UO_186 (O_186,N_2946,N_2950);
and UO_187 (O_187,N_2967,N_2946);
xnor UO_188 (O_188,N_2972,N_2942);
or UO_189 (O_189,N_2951,N_2941);
nor UO_190 (O_190,N_2952,N_2949);
nor UO_191 (O_191,N_2961,N_2983);
or UO_192 (O_192,N_2972,N_2945);
and UO_193 (O_193,N_2948,N_2966);
nor UO_194 (O_194,N_2948,N_2999);
or UO_195 (O_195,N_2990,N_2982);
nand UO_196 (O_196,N_2960,N_2958);
and UO_197 (O_197,N_2973,N_2998);
and UO_198 (O_198,N_2983,N_2960);
and UO_199 (O_199,N_2988,N_2943);
and UO_200 (O_200,N_2979,N_2942);
xor UO_201 (O_201,N_2941,N_2944);
nor UO_202 (O_202,N_2967,N_2975);
xor UO_203 (O_203,N_2962,N_2972);
or UO_204 (O_204,N_2976,N_2962);
or UO_205 (O_205,N_2953,N_2947);
or UO_206 (O_206,N_2993,N_2997);
and UO_207 (O_207,N_2992,N_2949);
or UO_208 (O_208,N_2949,N_2969);
nor UO_209 (O_209,N_2993,N_2996);
nor UO_210 (O_210,N_2987,N_2995);
nor UO_211 (O_211,N_2945,N_2964);
nand UO_212 (O_212,N_2978,N_2969);
xor UO_213 (O_213,N_2957,N_2968);
nand UO_214 (O_214,N_2956,N_2988);
and UO_215 (O_215,N_2997,N_2995);
nand UO_216 (O_216,N_2989,N_2987);
nand UO_217 (O_217,N_2983,N_2963);
nand UO_218 (O_218,N_2977,N_2947);
nand UO_219 (O_219,N_2958,N_2965);
or UO_220 (O_220,N_2945,N_2967);
nand UO_221 (O_221,N_2999,N_2952);
nor UO_222 (O_222,N_2966,N_2953);
xnor UO_223 (O_223,N_2942,N_2975);
and UO_224 (O_224,N_2984,N_2990);
nor UO_225 (O_225,N_2983,N_2985);
or UO_226 (O_226,N_2974,N_2992);
nand UO_227 (O_227,N_2950,N_2993);
nand UO_228 (O_228,N_2950,N_2998);
and UO_229 (O_229,N_2992,N_2964);
nor UO_230 (O_230,N_2953,N_2941);
or UO_231 (O_231,N_2959,N_2997);
nor UO_232 (O_232,N_2944,N_2973);
or UO_233 (O_233,N_2979,N_2994);
or UO_234 (O_234,N_2973,N_2976);
and UO_235 (O_235,N_2964,N_2943);
nand UO_236 (O_236,N_2991,N_2980);
and UO_237 (O_237,N_2957,N_2998);
xor UO_238 (O_238,N_2967,N_2979);
or UO_239 (O_239,N_2983,N_2945);
nor UO_240 (O_240,N_2943,N_2998);
and UO_241 (O_241,N_2996,N_2994);
or UO_242 (O_242,N_2997,N_2952);
nor UO_243 (O_243,N_2946,N_2942);
and UO_244 (O_244,N_2967,N_2986);
or UO_245 (O_245,N_2965,N_2990);
or UO_246 (O_246,N_2977,N_2986);
nor UO_247 (O_247,N_2969,N_2941);
nand UO_248 (O_248,N_2983,N_2952);
or UO_249 (O_249,N_2950,N_2971);
nand UO_250 (O_250,N_2987,N_2996);
nor UO_251 (O_251,N_2986,N_2964);
or UO_252 (O_252,N_2970,N_2985);
nor UO_253 (O_253,N_2992,N_2984);
nand UO_254 (O_254,N_2975,N_2982);
nand UO_255 (O_255,N_2991,N_2998);
or UO_256 (O_256,N_2947,N_2990);
and UO_257 (O_257,N_2966,N_2986);
nor UO_258 (O_258,N_2984,N_2997);
nor UO_259 (O_259,N_2942,N_2963);
nor UO_260 (O_260,N_2944,N_2984);
and UO_261 (O_261,N_2965,N_2983);
and UO_262 (O_262,N_2992,N_2996);
nor UO_263 (O_263,N_2950,N_2944);
nand UO_264 (O_264,N_2953,N_2945);
nand UO_265 (O_265,N_2944,N_2940);
xnor UO_266 (O_266,N_2995,N_2979);
nor UO_267 (O_267,N_2957,N_2989);
nor UO_268 (O_268,N_2989,N_2943);
xor UO_269 (O_269,N_2975,N_2962);
or UO_270 (O_270,N_2952,N_2984);
nor UO_271 (O_271,N_2995,N_2977);
or UO_272 (O_272,N_2982,N_2976);
and UO_273 (O_273,N_2966,N_2982);
and UO_274 (O_274,N_2951,N_2974);
xor UO_275 (O_275,N_2958,N_2954);
nand UO_276 (O_276,N_2968,N_2965);
nand UO_277 (O_277,N_2993,N_2957);
or UO_278 (O_278,N_2965,N_2982);
and UO_279 (O_279,N_2958,N_2942);
or UO_280 (O_280,N_2984,N_2958);
nand UO_281 (O_281,N_2960,N_2991);
nor UO_282 (O_282,N_2943,N_2987);
nor UO_283 (O_283,N_2979,N_2976);
or UO_284 (O_284,N_2968,N_2954);
nand UO_285 (O_285,N_2951,N_2988);
nand UO_286 (O_286,N_2966,N_2996);
nor UO_287 (O_287,N_2955,N_2953);
xor UO_288 (O_288,N_2963,N_2994);
xor UO_289 (O_289,N_2967,N_2950);
or UO_290 (O_290,N_2978,N_2946);
and UO_291 (O_291,N_2976,N_2960);
or UO_292 (O_292,N_2983,N_2978);
or UO_293 (O_293,N_2971,N_2989);
or UO_294 (O_294,N_2997,N_2940);
nor UO_295 (O_295,N_2955,N_2970);
xnor UO_296 (O_296,N_2980,N_2966);
nor UO_297 (O_297,N_2949,N_2968);
nand UO_298 (O_298,N_2972,N_2985);
nor UO_299 (O_299,N_2967,N_2981);
nand UO_300 (O_300,N_2991,N_2981);
and UO_301 (O_301,N_2983,N_2944);
nor UO_302 (O_302,N_2971,N_2959);
nor UO_303 (O_303,N_2980,N_2962);
nor UO_304 (O_304,N_2966,N_2961);
and UO_305 (O_305,N_2944,N_2974);
nand UO_306 (O_306,N_2951,N_2999);
and UO_307 (O_307,N_2975,N_2989);
nand UO_308 (O_308,N_2961,N_2977);
nor UO_309 (O_309,N_2973,N_2941);
nor UO_310 (O_310,N_2958,N_2994);
xor UO_311 (O_311,N_2975,N_2978);
nor UO_312 (O_312,N_2971,N_2956);
nand UO_313 (O_313,N_2955,N_2952);
or UO_314 (O_314,N_2962,N_2978);
or UO_315 (O_315,N_2953,N_2998);
and UO_316 (O_316,N_2960,N_2951);
or UO_317 (O_317,N_2967,N_2963);
nand UO_318 (O_318,N_2976,N_2972);
and UO_319 (O_319,N_2953,N_2948);
or UO_320 (O_320,N_2966,N_2991);
nor UO_321 (O_321,N_2951,N_2969);
and UO_322 (O_322,N_2966,N_2968);
or UO_323 (O_323,N_2976,N_2959);
or UO_324 (O_324,N_2979,N_2974);
and UO_325 (O_325,N_2959,N_2948);
and UO_326 (O_326,N_2968,N_2974);
or UO_327 (O_327,N_2944,N_2978);
or UO_328 (O_328,N_2985,N_2941);
nor UO_329 (O_329,N_2977,N_2981);
nand UO_330 (O_330,N_2966,N_2994);
nand UO_331 (O_331,N_2958,N_2987);
and UO_332 (O_332,N_2972,N_2984);
and UO_333 (O_333,N_2988,N_2964);
and UO_334 (O_334,N_2985,N_2974);
nand UO_335 (O_335,N_2998,N_2976);
nor UO_336 (O_336,N_2966,N_2962);
nand UO_337 (O_337,N_2980,N_2961);
or UO_338 (O_338,N_2985,N_2992);
or UO_339 (O_339,N_2941,N_2989);
nor UO_340 (O_340,N_2960,N_2984);
and UO_341 (O_341,N_2992,N_2970);
or UO_342 (O_342,N_2990,N_2954);
and UO_343 (O_343,N_2967,N_2982);
nor UO_344 (O_344,N_2991,N_2947);
nor UO_345 (O_345,N_2973,N_2966);
and UO_346 (O_346,N_2979,N_2988);
nand UO_347 (O_347,N_2983,N_2967);
or UO_348 (O_348,N_2971,N_2984);
or UO_349 (O_349,N_2979,N_2981);
or UO_350 (O_350,N_2999,N_2965);
nor UO_351 (O_351,N_2951,N_2995);
or UO_352 (O_352,N_2951,N_2986);
or UO_353 (O_353,N_2951,N_2998);
nand UO_354 (O_354,N_2980,N_2990);
and UO_355 (O_355,N_2970,N_2977);
and UO_356 (O_356,N_2947,N_2957);
and UO_357 (O_357,N_2981,N_2969);
nand UO_358 (O_358,N_2955,N_2974);
nand UO_359 (O_359,N_2945,N_2960);
nand UO_360 (O_360,N_2974,N_2980);
nor UO_361 (O_361,N_2965,N_2976);
or UO_362 (O_362,N_2981,N_2956);
or UO_363 (O_363,N_2971,N_2958);
and UO_364 (O_364,N_2974,N_2940);
or UO_365 (O_365,N_2953,N_2986);
or UO_366 (O_366,N_2967,N_2999);
nand UO_367 (O_367,N_2987,N_2948);
and UO_368 (O_368,N_2953,N_2984);
and UO_369 (O_369,N_2966,N_2951);
nor UO_370 (O_370,N_2972,N_2995);
nand UO_371 (O_371,N_2990,N_2995);
or UO_372 (O_372,N_2958,N_2981);
and UO_373 (O_373,N_2942,N_2966);
nand UO_374 (O_374,N_2983,N_2953);
or UO_375 (O_375,N_2961,N_2972);
nor UO_376 (O_376,N_2991,N_2942);
nand UO_377 (O_377,N_2963,N_2973);
nor UO_378 (O_378,N_2989,N_2962);
nand UO_379 (O_379,N_2949,N_2965);
nand UO_380 (O_380,N_2985,N_2956);
nor UO_381 (O_381,N_2940,N_2956);
and UO_382 (O_382,N_2993,N_2977);
or UO_383 (O_383,N_2977,N_2979);
xor UO_384 (O_384,N_2960,N_2987);
or UO_385 (O_385,N_2993,N_2955);
and UO_386 (O_386,N_2991,N_2995);
and UO_387 (O_387,N_2996,N_2945);
nand UO_388 (O_388,N_2972,N_2953);
or UO_389 (O_389,N_2999,N_2953);
nor UO_390 (O_390,N_2983,N_2972);
or UO_391 (O_391,N_2960,N_2978);
or UO_392 (O_392,N_2990,N_2993);
xnor UO_393 (O_393,N_2947,N_2942);
and UO_394 (O_394,N_2956,N_2990);
or UO_395 (O_395,N_2956,N_2974);
nor UO_396 (O_396,N_2942,N_2952);
and UO_397 (O_397,N_2941,N_2965);
and UO_398 (O_398,N_2977,N_2975);
and UO_399 (O_399,N_2952,N_2994);
nand UO_400 (O_400,N_2993,N_2983);
nor UO_401 (O_401,N_2989,N_2966);
nor UO_402 (O_402,N_2996,N_2967);
nor UO_403 (O_403,N_2967,N_2968);
or UO_404 (O_404,N_2985,N_2965);
xor UO_405 (O_405,N_2967,N_2941);
and UO_406 (O_406,N_2963,N_2991);
nor UO_407 (O_407,N_2956,N_2980);
nand UO_408 (O_408,N_2982,N_2971);
nor UO_409 (O_409,N_2951,N_2957);
xnor UO_410 (O_410,N_2981,N_2965);
and UO_411 (O_411,N_2942,N_2973);
nor UO_412 (O_412,N_2980,N_2954);
nand UO_413 (O_413,N_2976,N_2981);
xnor UO_414 (O_414,N_2951,N_2993);
or UO_415 (O_415,N_2998,N_2960);
or UO_416 (O_416,N_2987,N_2979);
nand UO_417 (O_417,N_2963,N_2984);
and UO_418 (O_418,N_2961,N_2963);
nand UO_419 (O_419,N_2992,N_2955);
and UO_420 (O_420,N_2984,N_2998);
nand UO_421 (O_421,N_2953,N_2949);
nand UO_422 (O_422,N_2950,N_2988);
or UO_423 (O_423,N_2951,N_2983);
nor UO_424 (O_424,N_2965,N_2942);
nand UO_425 (O_425,N_2953,N_2951);
xnor UO_426 (O_426,N_2976,N_2964);
nand UO_427 (O_427,N_2959,N_2983);
nand UO_428 (O_428,N_2975,N_2956);
or UO_429 (O_429,N_2979,N_2964);
nand UO_430 (O_430,N_2960,N_2954);
nor UO_431 (O_431,N_2941,N_2970);
and UO_432 (O_432,N_2973,N_2967);
nand UO_433 (O_433,N_2981,N_2950);
and UO_434 (O_434,N_2987,N_2978);
xnor UO_435 (O_435,N_2966,N_2969);
nand UO_436 (O_436,N_2992,N_2969);
or UO_437 (O_437,N_2996,N_2946);
nand UO_438 (O_438,N_2976,N_2986);
nand UO_439 (O_439,N_2977,N_2960);
nand UO_440 (O_440,N_2987,N_2993);
and UO_441 (O_441,N_2982,N_2951);
nand UO_442 (O_442,N_2979,N_2943);
nor UO_443 (O_443,N_2960,N_2972);
nand UO_444 (O_444,N_2985,N_2994);
and UO_445 (O_445,N_2963,N_2971);
nor UO_446 (O_446,N_2953,N_2997);
and UO_447 (O_447,N_2975,N_2958);
nor UO_448 (O_448,N_2975,N_2994);
and UO_449 (O_449,N_2984,N_2943);
and UO_450 (O_450,N_2963,N_2981);
nand UO_451 (O_451,N_2954,N_2986);
or UO_452 (O_452,N_2985,N_2957);
and UO_453 (O_453,N_2967,N_2995);
or UO_454 (O_454,N_2992,N_2980);
nand UO_455 (O_455,N_2973,N_2968);
nor UO_456 (O_456,N_2993,N_2947);
xor UO_457 (O_457,N_2952,N_2971);
nand UO_458 (O_458,N_2985,N_2951);
nor UO_459 (O_459,N_2948,N_2947);
nor UO_460 (O_460,N_2961,N_2940);
and UO_461 (O_461,N_2981,N_2947);
and UO_462 (O_462,N_2992,N_2990);
nand UO_463 (O_463,N_2949,N_2954);
xnor UO_464 (O_464,N_2973,N_2952);
nand UO_465 (O_465,N_2991,N_2974);
nor UO_466 (O_466,N_2961,N_2945);
xor UO_467 (O_467,N_2941,N_2966);
nor UO_468 (O_468,N_2984,N_2961);
xnor UO_469 (O_469,N_2969,N_2988);
nor UO_470 (O_470,N_2993,N_2975);
or UO_471 (O_471,N_2970,N_2957);
or UO_472 (O_472,N_2950,N_2995);
nor UO_473 (O_473,N_2942,N_2984);
or UO_474 (O_474,N_2963,N_2977);
nand UO_475 (O_475,N_2970,N_2996);
nor UO_476 (O_476,N_2965,N_2953);
and UO_477 (O_477,N_2962,N_2977);
nand UO_478 (O_478,N_2987,N_2944);
xor UO_479 (O_479,N_2977,N_2956);
nand UO_480 (O_480,N_2940,N_2945);
nand UO_481 (O_481,N_2950,N_2977);
nor UO_482 (O_482,N_2955,N_2947);
nand UO_483 (O_483,N_2997,N_2999);
nand UO_484 (O_484,N_2941,N_2997);
nor UO_485 (O_485,N_2962,N_2986);
or UO_486 (O_486,N_2988,N_2992);
and UO_487 (O_487,N_2946,N_2945);
nor UO_488 (O_488,N_2974,N_2952);
nor UO_489 (O_489,N_2984,N_2970);
and UO_490 (O_490,N_2970,N_2949);
xnor UO_491 (O_491,N_2973,N_2949);
xor UO_492 (O_492,N_2999,N_2940);
or UO_493 (O_493,N_2993,N_2956);
and UO_494 (O_494,N_2986,N_2940);
and UO_495 (O_495,N_2968,N_2948);
nor UO_496 (O_496,N_2946,N_2971);
nor UO_497 (O_497,N_2978,N_2984);
nor UO_498 (O_498,N_2945,N_2994);
or UO_499 (O_499,N_2999,N_2941);
endmodule