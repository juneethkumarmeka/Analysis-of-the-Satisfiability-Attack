module basic_2000_20000_2500_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_348,In_178);
or U1 (N_1,In_936,In_376);
nor U2 (N_2,In_1182,In_949);
and U3 (N_3,In_1581,In_56);
or U4 (N_4,In_529,In_94);
and U5 (N_5,In_1906,In_946);
nand U6 (N_6,In_1884,In_570);
or U7 (N_7,In_711,In_267);
and U8 (N_8,In_1837,In_709);
xor U9 (N_9,In_7,In_350);
nor U10 (N_10,In_1529,In_1000);
and U11 (N_11,In_277,In_117);
or U12 (N_12,In_1517,In_27);
and U13 (N_13,In_1457,In_822);
or U14 (N_14,In_1808,In_55);
xor U15 (N_15,In_1342,In_1344);
and U16 (N_16,In_1520,In_1999);
nand U17 (N_17,In_1634,In_1192);
or U18 (N_18,In_640,In_1735);
or U19 (N_19,In_1672,In_1785);
and U20 (N_20,In_1227,In_1459);
or U21 (N_21,In_1461,In_1867);
and U22 (N_22,In_1251,In_406);
nand U23 (N_23,In_351,In_1299);
and U24 (N_24,In_1932,In_1430);
nand U25 (N_25,In_420,In_1080);
xor U26 (N_26,In_1900,In_1352);
nor U27 (N_27,In_942,In_1774);
nor U28 (N_28,In_375,In_1198);
nand U29 (N_29,In_1945,In_576);
and U30 (N_30,In_928,In_229);
or U31 (N_31,In_400,In_1268);
nor U32 (N_32,In_980,In_768);
nor U33 (N_33,In_825,In_1249);
nand U34 (N_34,In_740,In_22);
nor U35 (N_35,In_1982,In_251);
xor U36 (N_36,In_392,In_1348);
nand U37 (N_37,In_1909,In_509);
or U38 (N_38,In_1812,In_1143);
nand U39 (N_39,In_829,In_585);
nor U40 (N_40,In_362,In_368);
or U41 (N_41,In_1665,In_1689);
xnor U42 (N_42,In_1066,In_1212);
xnor U43 (N_43,In_1781,In_1081);
nor U44 (N_44,In_1990,In_272);
and U45 (N_45,In_1599,In_632);
or U46 (N_46,In_74,In_702);
nor U47 (N_47,In_235,In_1978);
or U48 (N_48,In_811,In_1720);
nor U49 (N_49,In_525,In_1264);
nor U50 (N_50,In_1893,In_1061);
and U51 (N_51,In_138,In_107);
and U52 (N_52,In_46,In_1545);
nand U53 (N_53,In_1663,In_1283);
and U54 (N_54,In_372,In_1569);
nor U55 (N_55,In_1676,In_605);
and U56 (N_56,In_387,In_1436);
nor U57 (N_57,In_1358,In_1379);
or U58 (N_58,In_18,In_360);
and U59 (N_59,In_1841,In_1071);
and U60 (N_60,In_1836,In_1832);
xor U61 (N_61,In_757,In_165);
nand U62 (N_62,In_32,In_540);
nand U63 (N_63,In_494,In_662);
and U64 (N_64,In_1910,In_727);
or U65 (N_65,In_381,In_1626);
and U66 (N_66,In_672,In_1340);
or U67 (N_67,In_54,In_1141);
nor U68 (N_68,In_900,In_1522);
nand U69 (N_69,In_451,In_769);
nand U70 (N_70,In_1127,In_436);
nand U71 (N_71,In_1632,In_1038);
and U72 (N_72,In_1482,In_526);
or U73 (N_73,In_1547,In_992);
nand U74 (N_74,In_1651,In_135);
xor U75 (N_75,In_1871,In_1579);
and U76 (N_76,In_1662,In_732);
nand U77 (N_77,In_814,In_1408);
nor U78 (N_78,In_1318,In_1470);
and U79 (N_79,In_1012,In_613);
nor U80 (N_80,In_1953,In_1537);
nand U81 (N_81,In_23,In_579);
nand U82 (N_82,In_661,In_432);
nand U83 (N_83,In_296,In_523);
nand U84 (N_84,In_885,In_798);
and U85 (N_85,In_1388,In_1915);
xor U86 (N_86,In_256,In_1869);
and U87 (N_87,In_608,In_1438);
xnor U88 (N_88,In_1412,In_1823);
and U89 (N_89,In_1493,In_1715);
nor U90 (N_90,In_1842,In_1395);
or U91 (N_91,In_1698,In_1306);
nand U92 (N_92,In_158,In_857);
xor U93 (N_93,In_404,In_448);
and U94 (N_94,In_847,In_993);
and U95 (N_95,In_995,In_111);
nor U96 (N_96,In_1356,In_1446);
nand U97 (N_97,In_344,In_1428);
nor U98 (N_98,In_1743,In_1969);
or U99 (N_99,In_64,In_845);
xnor U100 (N_100,In_685,In_345);
nand U101 (N_101,In_1683,In_1445);
or U102 (N_102,In_934,In_1788);
or U103 (N_103,In_1267,In_527);
and U104 (N_104,In_1319,In_1189);
nor U105 (N_105,In_1309,In_602);
nand U106 (N_106,In_1116,In_1548);
and U107 (N_107,In_561,In_726);
xnor U108 (N_108,In_1901,In_1986);
or U109 (N_109,In_1184,In_385);
nor U110 (N_110,In_790,In_1233);
nand U111 (N_111,In_1684,In_1668);
and U112 (N_112,In_374,In_37);
and U113 (N_113,In_952,In_1584);
xor U114 (N_114,In_285,In_1010);
nor U115 (N_115,In_88,In_991);
or U116 (N_116,In_1571,In_164);
and U117 (N_117,In_500,In_245);
xor U118 (N_118,In_850,In_909);
nand U119 (N_119,In_1918,In_1941);
nand U120 (N_120,In_156,In_987);
and U121 (N_121,In_13,In_854);
or U122 (N_122,In_1670,In_622);
and U123 (N_123,In_276,In_1312);
nand U124 (N_124,In_1708,In_1142);
or U125 (N_125,In_1732,In_1594);
or U126 (N_126,In_904,In_736);
xor U127 (N_127,In_1937,In_532);
or U128 (N_128,In_1096,In_1508);
xor U129 (N_129,In_79,In_1544);
nor U130 (N_130,In_872,In_1677);
xnor U131 (N_131,In_1382,In_471);
nand U132 (N_132,In_1336,In_1642);
xnor U133 (N_133,In_1043,In_1039);
nor U134 (N_134,In_69,In_1567);
nand U135 (N_135,In_1629,In_102);
nand U136 (N_136,In_1343,In_421);
or U137 (N_137,In_748,In_817);
or U138 (N_138,In_265,In_259);
or U139 (N_139,In_324,In_1403);
nor U140 (N_140,In_1576,In_1657);
or U141 (N_141,In_468,In_1717);
nand U142 (N_142,In_631,In_180);
nand U143 (N_143,In_865,In_78);
nor U144 (N_144,In_1916,In_1917);
nor U145 (N_145,In_271,In_758);
nand U146 (N_146,In_1624,In_396);
and U147 (N_147,In_14,In_86);
nor U148 (N_148,In_1664,In_1751);
nor U149 (N_149,In_288,In_1484);
and U150 (N_150,In_1056,In_505);
and U151 (N_151,In_589,In_137);
or U152 (N_152,In_1686,In_827);
nor U153 (N_153,In_1321,In_452);
nand U154 (N_154,In_331,In_690);
nor U155 (N_155,In_1583,In_1165);
or U156 (N_156,In_333,In_53);
xnor U157 (N_157,In_1313,In_1351);
nor U158 (N_158,In_1682,In_1580);
xor U159 (N_159,In_1123,In_1852);
xnor U160 (N_160,In_475,In_1844);
and U161 (N_161,In_1749,In_1475);
xor U162 (N_162,In_1089,In_1033);
nand U163 (N_163,In_1185,In_985);
or U164 (N_164,In_314,In_515);
and U165 (N_165,In_352,In_628);
xor U166 (N_166,In_1350,In_1469);
nor U167 (N_167,In_29,In_1865);
xnor U168 (N_168,In_734,In_967);
nor U169 (N_169,In_1144,In_1125);
nor U170 (N_170,In_950,In_1013);
nor U171 (N_171,In_994,In_506);
xor U172 (N_172,In_1830,In_1654);
or U173 (N_173,In_104,In_582);
and U174 (N_174,In_724,In_1526);
nand U175 (N_175,In_1070,In_1007);
nor U176 (N_176,In_710,In_329);
nor U177 (N_177,In_1647,In_116);
nor U178 (N_178,In_1222,In_433);
and U179 (N_179,In_974,In_1725);
and U180 (N_180,In_1181,In_1064);
and U181 (N_181,In_407,In_260);
and U182 (N_182,In_1896,In_1001);
and U183 (N_183,In_1878,In_1887);
nor U184 (N_184,In_678,In_39);
xor U185 (N_185,In_1736,In_982);
xnor U186 (N_186,In_1699,In_299);
or U187 (N_187,In_1118,In_1965);
and U188 (N_188,In_1962,In_236);
xor U189 (N_189,In_804,In_999);
or U190 (N_190,In_1546,In_848);
xnor U191 (N_191,In_888,In_1169);
xnor U192 (N_192,In_282,In_1967);
nand U193 (N_193,In_1577,In_1630);
xnor U194 (N_194,In_1330,In_391);
and U195 (N_195,In_187,In_1147);
xor U196 (N_196,In_651,In_204);
nor U197 (N_197,In_818,In_1092);
nor U198 (N_198,In_1863,In_336);
nor U199 (N_199,In_1153,In_513);
and U200 (N_200,In_571,In_1199);
or U201 (N_201,In_1968,In_988);
xor U202 (N_202,In_1220,In_645);
xnor U203 (N_203,In_565,In_205);
or U204 (N_204,In_1922,In_1609);
nand U205 (N_205,In_76,In_1427);
nand U206 (N_206,In_114,In_971);
nor U207 (N_207,In_1053,In_130);
or U208 (N_208,In_1806,In_522);
and U209 (N_209,In_1140,In_856);
nand U210 (N_210,In_11,In_887);
and U211 (N_211,In_1180,In_428);
or U212 (N_212,In_340,In_925);
xnor U213 (N_213,In_1897,In_612);
nor U214 (N_214,In_166,In_1478);
or U215 (N_215,In_84,In_1462);
and U216 (N_216,In_1355,In_1276);
or U217 (N_217,In_1491,In_170);
nor U218 (N_218,In_1300,In_1560);
and U219 (N_219,In_1762,In_1757);
nor U220 (N_220,In_1138,In_318);
nor U221 (N_221,In_1973,In_152);
or U222 (N_222,In_1471,In_780);
and U223 (N_223,In_761,In_639);
nand U224 (N_224,In_1173,In_1880);
and U225 (N_225,In_1800,In_466);
nand U226 (N_226,In_370,In_849);
nor U227 (N_227,In_77,In_1022);
nor U228 (N_228,In_1155,In_714);
nor U229 (N_229,In_125,In_830);
nor U230 (N_230,In_1817,In_1995);
nand U231 (N_231,In_160,In_603);
xor U232 (N_232,In_241,In_721);
xnor U233 (N_233,In_250,In_1373);
and U234 (N_234,In_313,In_590);
xor U235 (N_235,In_1332,In_292);
xnor U236 (N_236,In_1819,In_1543);
or U237 (N_237,In_749,In_781);
nor U238 (N_238,In_203,In_363);
nand U239 (N_239,In_1855,In_1858);
and U240 (N_240,In_1111,In_408);
or U241 (N_241,In_666,In_1727);
nor U242 (N_242,In_1710,In_207);
nand U243 (N_243,In_869,In_40);
xor U244 (N_244,In_1246,In_1667);
xnor U245 (N_245,In_1316,In_1456);
and U246 (N_246,In_587,In_504);
nor U247 (N_247,In_816,In_866);
nand U248 (N_248,In_550,In_1929);
and U249 (N_249,In_596,In_334);
nor U250 (N_250,In_1661,In_1447);
or U251 (N_251,In_927,In_723);
and U252 (N_252,In_1981,In_939);
and U253 (N_253,In_1602,In_1016);
and U254 (N_254,In_948,In_71);
and U255 (N_255,In_1082,In_1091);
xnor U256 (N_256,In_1151,In_1020);
nand U257 (N_257,In_442,In_28);
and U258 (N_258,In_703,In_1210);
or U259 (N_259,In_1886,In_1881);
xnor U260 (N_260,In_384,In_636);
or U261 (N_261,In_87,In_933);
xor U262 (N_262,In_127,In_80);
or U263 (N_263,In_239,In_1317);
nand U264 (N_264,In_653,In_255);
nand U265 (N_265,In_1390,In_1158);
and U266 (N_266,In_1791,In_1925);
nor U267 (N_267,In_1253,In_446);
or U268 (N_268,In_96,In_1364);
or U269 (N_269,In_218,In_543);
or U270 (N_270,In_1051,In_1879);
nor U271 (N_271,In_1617,In_258);
nor U272 (N_272,In_1902,In_891);
or U273 (N_273,In_1248,In_367);
and U274 (N_274,In_1899,In_1231);
and U275 (N_275,In_737,In_1154);
or U276 (N_276,In_1818,In_57);
nand U277 (N_277,In_1095,In_133);
or U278 (N_278,In_1301,In_1174);
and U279 (N_279,In_1345,In_641);
xor U280 (N_280,In_917,In_903);
xnor U281 (N_281,In_1333,In_1826);
or U282 (N_282,In_1988,In_1741);
and U283 (N_283,In_283,In_747);
or U284 (N_284,In_1025,In_968);
and U285 (N_285,In_1553,In_693);
xor U286 (N_286,In_1961,In_1401);
nor U287 (N_287,In_530,In_253);
or U288 (N_288,In_172,In_754);
and U289 (N_289,In_325,In_915);
nor U290 (N_290,In_932,In_521);
nor U291 (N_291,In_581,In_1705);
nand U292 (N_292,In_1372,In_1843);
xnor U293 (N_293,In_1407,In_1566);
nor U294 (N_294,In_1132,In_435);
nand U295 (N_295,In_580,In_669);
nor U296 (N_296,In_517,In_615);
or U297 (N_297,In_183,In_1644);
xor U298 (N_298,In_63,In_139);
nand U299 (N_299,In_713,In_2);
nor U300 (N_300,In_1112,In_1744);
nor U301 (N_301,In_1964,In_1816);
nand U302 (N_302,In_1604,In_695);
or U303 (N_303,In_38,In_518);
xor U304 (N_304,In_1850,In_1448);
nand U305 (N_305,In_1019,In_1883);
nand U306 (N_306,In_588,In_1513);
or U307 (N_307,In_177,In_1308);
nand U308 (N_308,In_1337,In_873);
nand U309 (N_309,In_427,In_91);
nand U310 (N_310,In_1347,In_1534);
xnor U311 (N_311,In_1422,In_257);
xnor U312 (N_312,In_1911,In_1799);
xor U313 (N_313,In_564,In_1055);
and U314 (N_314,In_1149,In_1633);
nand U315 (N_315,In_1671,In_692);
nand U316 (N_316,In_1835,In_1655);
nand U317 (N_317,In_1261,In_499);
and U318 (N_318,In_592,In_677);
nor U319 (N_319,In_943,In_547);
nand U320 (N_320,In_3,In_1714);
or U321 (N_321,In_658,In_1083);
nand U322 (N_322,In_1814,In_1801);
xor U323 (N_323,In_356,In_49);
or U324 (N_324,In_246,In_567);
nand U325 (N_325,In_686,In_1240);
xor U326 (N_326,In_846,In_1483);
nor U327 (N_327,In_263,In_1845);
nand U328 (N_328,In_275,In_575);
and U329 (N_329,In_1955,In_1769);
and U330 (N_330,In_227,In_868);
xor U331 (N_331,In_1110,In_614);
nand U332 (N_332,In_231,In_935);
and U333 (N_333,In_1938,In_182);
nand U334 (N_334,In_377,In_434);
or U335 (N_335,In_1612,In_121);
xor U336 (N_336,In_1550,In_1585);
xor U337 (N_337,In_1891,In_365);
and U338 (N_338,In_1172,In_896);
and U339 (N_339,In_910,In_1338);
and U340 (N_340,In_689,In_202);
and U341 (N_341,In_284,In_1875);
nand U342 (N_342,In_1572,In_890);
xnor U343 (N_343,In_1223,In_1414);
nor U344 (N_344,In_520,In_1178);
nand U345 (N_345,In_1608,In_1591);
xnor U346 (N_346,In_1856,In_1564);
or U347 (N_347,In_621,In_1040);
nand U348 (N_348,In_1215,In_1587);
nor U349 (N_349,In_1693,In_269);
and U350 (N_350,In_1979,In_712);
nand U351 (N_351,In_624,In_1479);
and U352 (N_352,In_663,In_1574);
nor U353 (N_353,In_1256,In_1179);
xnor U354 (N_354,In_337,In_338);
or U355 (N_355,In_1614,In_112);
or U356 (N_356,In_1488,In_1079);
xnor U357 (N_357,In_1429,In_842);
xor U358 (N_358,In_1985,In_1695);
nor U359 (N_359,In_62,In_198);
nor U360 (N_360,In_1512,In_820);
and U361 (N_361,In_1650,In_461);
nor U362 (N_362,In_1864,In_1870);
nand U363 (N_363,In_278,In_293);
xor U364 (N_364,In_1077,In_1966);
xnor U365 (N_365,In_349,In_1728);
nand U366 (N_366,In_1600,In_1226);
or U367 (N_367,In_99,In_1868);
or U368 (N_368,In_836,In_1556);
or U369 (N_369,In_1764,In_771);
nand U370 (N_370,In_501,In_1669);
and U371 (N_371,In_1031,In_1775);
xnor U372 (N_372,In_1573,In_766);
xnor U373 (N_373,In_361,In_1252);
nand U374 (N_374,In_1829,In_1723);
nor U375 (N_375,In_1217,In_1521);
xor U376 (N_376,In_1653,In_457);
nand U377 (N_377,In_248,In_167);
xor U378 (N_378,In_1726,In_149);
nor U379 (N_379,In_1489,In_1058);
nand U380 (N_380,In_752,In_1778);
nand U381 (N_381,In_1273,In_1375);
and U382 (N_382,In_358,In_477);
xnor U383 (N_383,In_1416,In_717);
xnor U384 (N_384,In_431,In_469);
nand U385 (N_385,In_1797,In_1136);
or U386 (N_386,In_261,In_1063);
and U387 (N_387,In_1700,In_153);
or U388 (N_388,In_1497,In_220);
nor U389 (N_389,In_735,In_774);
xnor U390 (N_390,In_719,In_1767);
and U391 (N_391,In_792,In_1378);
xor U392 (N_392,In_1558,In_196);
xor U393 (N_393,In_1100,In_24);
xnor U394 (N_394,In_58,In_1354);
or U395 (N_395,In_577,In_146);
nand U396 (N_396,In_45,In_1511);
and U397 (N_397,In_459,In_716);
nand U398 (N_398,In_1825,In_1674);
xnor U399 (N_399,In_535,In_1224);
xnor U400 (N_400,In_249,In_660);
and U401 (N_401,In_1152,In_1833);
and U402 (N_402,In_136,In_775);
nand U403 (N_403,In_1235,In_1162);
or U404 (N_404,In_311,In_1464);
nor U405 (N_405,In_819,In_1376);
xnor U406 (N_406,In_50,In_1627);
or U407 (N_407,In_1384,In_1716);
or U408 (N_408,In_807,In_1324);
xnor U409 (N_409,In_414,In_1588);
and U410 (N_410,In_493,In_1204);
or U411 (N_411,In_1646,In_607);
or U412 (N_412,In_1385,In_439);
xor U413 (N_413,In_274,In_357);
nand U414 (N_414,In_1921,In_1292);
nor U415 (N_415,In_528,In_1903);
or U416 (N_416,In_295,In_1828);
xnor U417 (N_417,In_430,In_455);
and U418 (N_418,In_1398,In_566);
and U419 (N_419,In_1258,In_899);
xor U420 (N_420,In_560,In_1768);
and U421 (N_421,In_1940,In_1059);
xor U422 (N_422,In_83,In_98);
and U423 (N_423,In_1150,In_682);
nand U424 (N_424,In_97,In_657);
nor U425 (N_425,In_225,In_75);
nor U426 (N_426,In_958,In_1387);
or U427 (N_427,In_123,In_534);
xnor U428 (N_428,In_1259,In_1976);
nand U429 (N_429,In_1820,In_676);
xnor U430 (N_430,In_1983,In_597);
nand U431 (N_431,In_1196,In_655);
nor U432 (N_432,In_1054,In_1107);
nor U433 (N_433,In_569,In_463);
and U434 (N_434,In_929,In_1792);
nor U435 (N_435,In_1796,In_1255);
and U436 (N_436,In_1514,In_1989);
and U437 (N_437,In_35,In_1718);
nor U438 (N_438,In_1085,In_397);
and U439 (N_439,In_1625,In_926);
and U440 (N_440,In_963,In_728);
or U441 (N_441,In_892,In_1197);
or U442 (N_442,In_186,In_1);
nor U443 (N_443,In_524,In_1076);
nor U444 (N_444,In_1238,In_415);
nand U445 (N_445,In_833,In_1994);
nand U446 (N_446,In_252,In_1302);
nor U447 (N_447,In_1562,In_1113);
xor U448 (N_448,In_492,In_1425);
nand U449 (N_449,In_1750,In_411);
or U450 (N_450,In_889,In_744);
and U451 (N_451,In_1367,In_268);
nand U452 (N_452,In_986,In_326);
nor U453 (N_453,In_1130,In_619);
or U454 (N_454,In_1810,In_1164);
or U455 (N_455,In_1017,In_1274);
and U456 (N_456,In_1139,In_1790);
xor U457 (N_457,In_1963,In_905);
or U458 (N_458,In_650,In_611);
or U459 (N_459,In_1601,In_1244);
nand U460 (N_460,In_1305,In_1729);
xor U461 (N_461,In_131,In_595);
xnor U462 (N_462,In_1314,In_1702);
or U463 (N_463,In_1277,In_806);
or U464 (N_464,In_1450,In_1760);
and U465 (N_465,In_609,In_1296);
nand U466 (N_466,In_1538,In_1894);
nor U467 (N_467,In_481,In_1948);
xnor U468 (N_468,In_1115,In_1861);
nand U469 (N_469,In_214,In_698);
and U470 (N_470,In_1697,In_1463);
nor U471 (N_471,In_1129,In_541);
nor U472 (N_472,In_1639,In_1809);
nor U473 (N_473,In_147,In_209);
or U474 (N_474,In_1128,In_959);
nand U475 (N_475,In_1822,In_199);
and U476 (N_476,In_777,In_1752);
nand U477 (N_477,In_332,In_1106);
or U478 (N_478,In_454,In_1005);
or U479 (N_479,In_1168,In_1758);
nand U480 (N_480,In_1593,In_1794);
xnor U481 (N_481,In_70,In_1440);
nor U482 (N_482,In_839,In_1687);
and U483 (N_483,In_844,In_48);
nor U484 (N_484,In_1563,In_1023);
nand U485 (N_485,In_1417,In_977);
nand U486 (N_486,In_1200,In_502);
and U487 (N_487,In_545,In_1203);
nor U488 (N_488,In_1166,In_584);
nor U489 (N_489,In_1090,In_210);
nor U490 (N_490,In_1289,In_549);
and U491 (N_491,In_1160,In_1008);
and U492 (N_492,In_573,In_1952);
xnor U493 (N_493,In_1439,In_1854);
or U494 (N_494,In_1939,In_232);
nor U495 (N_495,In_1782,In_1539);
or U496 (N_496,In_1673,In_65);
or U497 (N_497,In_141,In_1451);
and U498 (N_498,In_859,In_169);
xnor U499 (N_499,In_1786,In_1536);
or U500 (N_500,In_1377,In_756);
nor U501 (N_501,In_1631,In_812);
nand U502 (N_502,In_9,In_443);
nand U503 (N_503,In_34,In_1021);
nand U504 (N_504,In_593,In_416);
nand U505 (N_505,In_67,In_1097);
nand U506 (N_506,In_1487,In_490);
nand U507 (N_507,In_1949,In_36);
or U508 (N_508,In_1892,In_322);
nand U509 (N_509,In_185,In_1024);
or U510 (N_510,In_776,In_1685);
nor U511 (N_511,In_1177,In_42);
nor U512 (N_512,In_1777,In_343);
or U513 (N_513,In_1862,In_895);
or U514 (N_514,In_1831,In_307);
nand U515 (N_515,In_234,In_906);
xor U516 (N_516,In_1122,In_1610);
nor U517 (N_517,In_161,In_617);
or U518 (N_518,In_4,In_824);
nand U519 (N_519,In_1286,In_1265);
or U520 (N_520,In_557,In_51);
nand U521 (N_521,In_106,In_742);
nor U522 (N_522,In_6,In_1230);
and U523 (N_523,In_1485,In_200);
nor U524 (N_524,In_870,In_423);
nor U525 (N_525,In_1065,In_1392);
and U526 (N_526,In_1984,In_1191);
or U527 (N_527,In_305,In_1303);
nand U528 (N_528,In_1291,In_841);
and U529 (N_529,In_516,In_1003);
and U530 (N_530,In_1114,In_862);
nor U531 (N_531,In_563,In_1552);
and U532 (N_532,In_132,In_1467);
xnor U533 (N_533,In_262,In_1641);
nor U534 (N_534,In_938,In_976);
and U535 (N_535,In_1795,In_786);
or U536 (N_536,In_1103,In_539);
and U537 (N_537,In_1015,In_355);
xor U538 (N_538,In_770,In_1409);
nand U539 (N_539,In_1014,In_1557);
xor U540 (N_540,In_941,In_855);
nand U541 (N_541,In_1549,In_763);
and U542 (N_542,In_201,In_1201);
nand U543 (N_543,In_918,In_1346);
and U544 (N_544,In_1435,In_1688);
xnor U545 (N_545,In_1270,In_449);
xnor U546 (N_546,In_953,In_1369);
nand U547 (N_547,In_1997,In_996);
or U548 (N_548,In_1027,In_243);
or U549 (N_549,In_1293,In_1272);
xor U550 (N_550,In_89,In_683);
nor U551 (N_551,In_1592,In_637);
nor U552 (N_552,In_705,In_1241);
or U553 (N_553,In_1047,In_1466);
or U554 (N_554,In_667,In_1045);
nand U555 (N_555,In_171,In_674);
nor U556 (N_556,In_1254,In_1525);
and U557 (N_557,In_1171,In_1516);
nor U558 (N_558,In_1205,In_1737);
and U559 (N_559,In_90,In_1857);
and U560 (N_560,In_552,In_730);
nor U561 (N_561,In_1243,In_1481);
and U562 (N_562,In_330,In_1357);
and U563 (N_563,In_1402,In_898);
and U564 (N_564,In_778,In_1490);
and U565 (N_565,In_1783,In_93);
or U566 (N_566,In_1944,In_1619);
xor U567 (N_567,In_731,In_1618);
and U568 (N_568,In_670,In_955);
xor U569 (N_569,In_497,In_984);
or U570 (N_570,In_1959,In_19);
xor U571 (N_571,In_1405,In_1499);
nand U572 (N_572,In_583,In_956);
or U573 (N_573,In_1780,In_598);
or U574 (N_574,In_1960,In_386);
and U575 (N_575,In_1060,In_779);
nand U576 (N_576,In_1441,In_1946);
nand U577 (N_577,In_542,In_796);
xnor U578 (N_578,In_441,In_460);
nand U579 (N_579,In_572,In_894);
nor U580 (N_580,In_979,In_718);
nand U581 (N_581,In_217,In_456);
xnor U582 (N_582,In_558,In_840);
nor U583 (N_583,In_883,In_864);
xnor U584 (N_584,In_1104,In_861);
nor U585 (N_585,In_1044,In_1094);
nand U586 (N_586,In_1635,In_491);
or U587 (N_587,In_1658,In_1515);
or U588 (N_588,In_725,In_1186);
nor U589 (N_589,In_41,In_12);
and U590 (N_590,In_1360,In_279);
xor U591 (N_591,In_25,In_823);
nor U592 (N_592,In_405,In_1393);
or U593 (N_593,In_66,In_1742);
nor U594 (N_594,In_838,In_1889);
or U595 (N_595,In_422,In_916);
xor U596 (N_596,In_1413,In_708);
and U597 (N_597,In_1611,In_244);
xor U598 (N_598,In_1518,In_1032);
xor U599 (N_599,In_881,In_1914);
nand U600 (N_600,In_638,In_867);
nor U601 (N_601,In_301,In_664);
xor U602 (N_602,In_364,In_1386);
and U603 (N_603,In_1190,In_1410);
or U604 (N_604,In_223,In_21);
nor U605 (N_605,In_1209,In_195);
and U606 (N_606,In_1187,In_1406);
or U607 (N_607,In_1009,In_1018);
or U608 (N_608,In_1334,In_1006);
or U609 (N_609,In_495,In_1322);
nand U610 (N_610,In_1500,In_1146);
xnor U611 (N_611,In_1363,In_110);
or U612 (N_612,In_179,In_242);
nor U613 (N_613,In_733,In_1062);
or U614 (N_614,In_1640,In_1126);
xnor U615 (N_615,In_1802,In_81);
xor U616 (N_616,In_880,In_1444);
and U617 (N_617,In_1958,In_1298);
or U618 (N_618,In_1805,In_1389);
nor U619 (N_619,In_1559,In_794);
and U620 (N_620,In_1072,In_458);
or U621 (N_621,In_1991,In_813);
and U622 (N_622,In_1331,In_373);
or U623 (N_623,In_315,In_618);
or U624 (N_624,In_1766,In_450);
nand U625 (N_625,In_1052,In_1637);
or U626 (N_626,In_148,In_1613);
nand U627 (N_627,In_599,In_1380);
and U628 (N_628,In_480,In_1362);
nor U629 (N_629,In_1279,In_1509);
and U630 (N_630,In_924,In_1297);
and U631 (N_631,In_126,In_652);
and U632 (N_632,In_1747,In_1904);
xnor U633 (N_633,In_961,In_1636);
nor U634 (N_634,In_1603,In_1565);
or U635 (N_635,In_962,In_1753);
nand U636 (N_636,In_1815,In_473);
nor U637 (N_637,In_983,In_403);
nand U638 (N_638,In_1211,In_1311);
or U639 (N_639,In_82,In_1099);
or U640 (N_640,In_1163,In_767);
nor U641 (N_641,In_797,In_317);
nor U642 (N_642,In_1824,In_341);
nor U643 (N_643,In_1993,In_1908);
and U644 (N_644,In_750,In_1692);
xnor U645 (N_645,In_510,In_828);
xnor U646 (N_646,In_1418,In_810);
or U647 (N_647,In_378,In_393);
xnor U648 (N_648,In_772,In_783);
xnor U649 (N_649,In_383,In_1895);
nor U650 (N_650,In_1652,In_1229);
xor U651 (N_651,In_1523,In_675);
xnor U652 (N_652,In_1763,In_1504);
nand U653 (N_653,In_1535,In_1067);
or U654 (N_654,In_1453,In_1420);
or U655 (N_655,In_142,In_1454);
or U656 (N_656,In_1175,In_688);
nand U657 (N_657,In_1415,In_1934);
xor U658 (N_658,In_1847,In_1771);
nor U659 (N_659,In_1505,In_1349);
nand U660 (N_660,In_1383,In_419);
nor U661 (N_661,In_438,In_291);
and U662 (N_662,In_237,In_831);
nor U663 (N_663,In_635,In_1590);
and U664 (N_664,In_1218,In_1507);
or U665 (N_665,In_1145,In_26);
nor U666 (N_666,In_118,In_1159);
xor U667 (N_667,In_739,In_1754);
xor U668 (N_668,In_1659,In_809);
nand U669 (N_669,In_175,In_1029);
xor U670 (N_670,In_852,In_327);
xnor U671 (N_671,In_1882,In_591);
nor U672 (N_672,In_1848,In_700);
nand U673 (N_673,In_551,In_1531);
nand U674 (N_674,In_462,In_1931);
and U675 (N_675,In_1711,In_1872);
or U676 (N_676,In_1761,In_1074);
nor U677 (N_677,In_467,In_646);
and U678 (N_678,In_1046,In_1473);
nand U679 (N_679,In_447,In_1068);
nor U680 (N_680,In_1370,In_1779);
or U681 (N_681,In_1853,In_417);
nor U682 (N_682,In_893,In_902);
nand U683 (N_683,In_379,In_464);
and U684 (N_684,In_803,In_445);
xor U685 (N_685,In_219,In_907);
nor U686 (N_686,In_951,In_537);
nor U687 (N_687,In_858,In_649);
and U688 (N_688,In_1712,In_47);
nor U689 (N_689,In_1266,In_1492);
nor U690 (N_690,In_371,In_1148);
and U691 (N_691,In_554,In_1616);
nor U692 (N_692,In_173,In_553);
nand U693 (N_693,In_323,In_20);
and U694 (N_694,In_1216,In_476);
xnor U695 (N_695,In_1325,In_233);
and U696 (N_696,In_287,In_1339);
nand U697 (N_697,In_208,In_206);
and U698 (N_698,In_681,In_1936);
xnor U699 (N_699,In_101,In_1834);
and U700 (N_700,In_1411,In_878);
xor U701 (N_701,In_656,In_1620);
nor U702 (N_702,In_1933,In_784);
nor U703 (N_703,In_1998,In_115);
xor U704 (N_704,In_212,In_1666);
and U705 (N_705,In_1078,In_1706);
nand U706 (N_706,In_1368,In_821);
and U707 (N_707,In_930,In_230);
or U708 (N_708,In_793,In_1004);
nand U709 (N_709,In_155,In_1912);
xnor U710 (N_710,In_743,In_538);
xor U711 (N_711,In_879,In_1798);
nand U712 (N_712,In_1117,In_1956);
or U713 (N_713,In_1789,In_1102);
or U714 (N_714,In_312,In_759);
nand U715 (N_715,In_1101,In_286);
and U716 (N_716,In_751,In_181);
xnor U717 (N_717,In_1260,In_145);
xor U718 (N_718,In_399,In_59);
xor U719 (N_719,In_1787,In_871);
or U720 (N_720,In_496,In_425);
and U721 (N_721,In_701,In_800);
or U722 (N_722,In_696,In_228);
or U723 (N_723,In_308,In_1704);
or U724 (N_724,In_548,In_514);
xnor U725 (N_725,In_531,In_1381);
or U726 (N_726,In_508,In_465);
xor U727 (N_727,In_707,In_1502);
and U728 (N_728,In_908,In_5);
and U729 (N_729,In_85,In_799);
or U730 (N_730,In_1207,In_1776);
xnor U731 (N_731,In_1399,In_1759);
or U732 (N_732,In_555,In_321);
or U733 (N_733,In_290,In_388);
nor U734 (N_734,In_1236,In_1951);
xor U735 (N_735,In_1746,In_100);
and U736 (N_736,In_1935,In_832);
or U737 (N_737,In_1028,In_1161);
xor U738 (N_738,In_1694,In_1073);
xor U739 (N_739,In_401,In_1284);
xnor U740 (N_740,In_347,In_1443);
nand U741 (N_741,In_1851,In_654);
xnor U742 (N_742,In_1554,In_762);
nor U743 (N_743,In_969,In_1898);
or U744 (N_744,In_886,In_1294);
or U745 (N_745,In_1838,In_874);
or U746 (N_746,In_1885,In_474);
nand U747 (N_747,In_215,In_1335);
nand U748 (N_748,In_1086,In_302);
and U749 (N_749,In_1943,In_1503);
nand U750 (N_750,In_310,In_973);
and U751 (N_751,In_273,In_746);
nand U752 (N_752,In_1452,In_1860);
and U753 (N_753,In_913,In_211);
or U754 (N_754,In_1645,In_1221);
nand U755 (N_755,In_1755,In_536);
nor U756 (N_756,In_1036,In_1075);
xnor U757 (N_757,In_1873,In_978);
xor U758 (N_758,In_1426,In_604);
nand U759 (N_759,In_1119,In_1980);
and U760 (N_760,In_1734,In_479);
nor U761 (N_761,In_1359,In_745);
nor U762 (N_762,In_630,In_1905);
nor U763 (N_763,In_1920,In_1807);
nand U764 (N_764,In_1206,In_489);
nand U765 (N_765,In_954,In_1188);
nor U766 (N_766,In_1011,In_1468);
and U767 (N_767,In_163,In_1121);
xor U768 (N_768,In_788,In_1374);
and U769 (N_769,In_1605,In_544);
xnor U770 (N_770,In_159,In_1719);
and U771 (N_771,In_168,In_339);
xor U772 (N_772,In_1972,In_1225);
nand U773 (N_773,In_722,In_1578);
nand U774 (N_774,In_964,In_1275);
or U775 (N_775,In_140,In_95);
or U776 (N_776,In_1304,In_741);
nor U777 (N_777,In_782,In_1323);
or U778 (N_778,In_1432,In_998);
nor U779 (N_779,In_1282,In_193);
nand U780 (N_780,In_1105,In_1195);
and U781 (N_781,In_911,In_1495);
and U782 (N_782,In_1568,In_1315);
or U783 (N_783,In_715,In_1437);
nor U784 (N_784,In_1239,In_860);
nor U785 (N_785,In_1738,In_981);
or U786 (N_786,In_1476,In_1480);
nand U787 (N_787,In_304,In_300);
xnor U788 (N_788,In_691,In_1219);
nor U789 (N_789,In_426,In_395);
xnor U790 (N_790,In_1607,In_1524);
xnor U791 (N_791,In_1278,In_31);
xnor U792 (N_792,In_328,In_1134);
nor U793 (N_793,In_1245,In_194);
or U794 (N_794,In_60,In_72);
nand U795 (N_795,In_247,In_174);
xor U796 (N_796,In_1739,In_1721);
nor U797 (N_797,In_1713,In_1449);
or U798 (N_798,In_912,In_787);
or U799 (N_799,In_346,In_568);
and U800 (N_800,In_546,In_1722);
xnor U801 (N_801,In_923,In_1551);
xor U802 (N_802,In_1923,In_738);
nor U803 (N_803,In_151,In_1257);
and U804 (N_804,In_629,In_1193);
and U805 (N_805,In_1326,In_1035);
nor U806 (N_806,In_221,In_940);
and U807 (N_807,In_240,In_627);
and U808 (N_808,In_1866,In_306);
nand U809 (N_809,In_1271,In_1397);
nand U810 (N_810,In_488,In_1606);
xnor U811 (N_811,In_398,In_487);
nor U812 (N_812,In_150,In_1400);
xnor U813 (N_813,In_128,In_1773);
nor U814 (N_814,In_1486,In_1532);
nor U815 (N_815,In_1108,In_366);
xor U816 (N_816,In_478,In_143);
xnor U817 (N_817,In_1846,In_1396);
and U818 (N_818,In_1170,In_483);
and U819 (N_819,In_1530,In_484);
nand U820 (N_820,In_922,In_919);
xnor U821 (N_821,In_1628,In_1057);
nor U822 (N_822,In_1597,In_877);
and U823 (N_823,In_1703,In_1947);
nand U824 (N_824,In_808,In_625);
xor U825 (N_825,In_390,In_972);
nand U826 (N_826,In_642,In_1030);
xnor U827 (N_827,In_556,In_498);
and U828 (N_828,In_1131,In_753);
and U829 (N_829,In_1109,In_1623);
and U830 (N_830,In_586,In_1034);
nor U831 (N_831,In_1924,In_1269);
and U832 (N_832,In_1496,In_1026);
xor U833 (N_833,In_1733,In_297);
xnor U834 (N_834,In_801,In_1840);
nor U835 (N_835,In_512,In_1974);
nor U836 (N_836,In_1877,In_380);
and U837 (N_837,In_1156,In_644);
or U838 (N_838,In_1849,In_197);
or U839 (N_839,In_1926,In_440);
nand U840 (N_840,In_990,In_1093);
and U841 (N_841,In_697,In_1542);
nand U842 (N_842,In_760,In_1098);
xnor U843 (N_843,In_188,In_1048);
xnor U844 (N_844,In_945,In_1731);
and U845 (N_845,In_1069,In_1555);
nand U846 (N_846,In_16,In_1307);
and U847 (N_847,In_680,In_1088);
nor U848 (N_848,In_947,In_213);
xor U849 (N_849,In_1859,In_389);
xnor U850 (N_850,In_989,In_1970);
nand U851 (N_851,In_1730,In_626);
xnor U852 (N_852,In_1678,In_129);
xnor U853 (N_853,In_157,In_1615);
or U854 (N_854,In_289,In_402);
nor U855 (N_855,In_1784,In_342);
and U856 (N_856,In_1950,In_1680);
and U857 (N_857,In_511,In_353);
and U858 (N_858,In_1242,In_1421);
nand U859 (N_859,In_134,In_1954);
nand U860 (N_860,In_1194,In_1701);
and U861 (N_861,In_1084,In_1745);
nand U862 (N_862,In_931,In_1295);
xor U863 (N_863,In_453,In_1595);
xor U864 (N_864,In_533,In_1281);
or U865 (N_865,In_1120,In_144);
nand U866 (N_866,In_1656,In_960);
nor U867 (N_867,In_1527,In_73);
xnor U868 (N_868,In_190,In_835);
xor U869 (N_869,In_578,In_966);
xnor U870 (N_870,In_1287,In_162);
nand U871 (N_871,In_1002,In_382);
or U872 (N_872,In_562,In_1498);
xor U873 (N_873,In_429,In_1575);
and U874 (N_874,In_1582,In_1213);
nand U875 (N_875,In_1460,In_1208);
or U876 (N_876,In_394,In_610);
and U877 (N_877,In_805,In_1975);
nor U878 (N_878,In_1472,In_875);
or U879 (N_879,In_965,In_1971);
or U880 (N_880,In_643,In_1285);
nand U881 (N_881,In_1811,In_1157);
and U882 (N_882,In_222,In_1176);
or U883 (N_883,In_668,In_1827);
and U884 (N_884,In_1124,In_1740);
nor U885 (N_885,In_1280,In_620);
nor U886 (N_886,In_1087,In_17);
nand U887 (N_887,In_684,In_785);
xnor U888 (N_888,In_1433,In_1050);
nor U889 (N_889,In_1167,In_1262);
and U890 (N_890,In_1528,In_472);
xnor U891 (N_891,In_1391,In_192);
and U892 (N_892,In_826,In_1638);
or U893 (N_893,In_103,In_413);
nand U894 (N_894,In_1648,In_294);
and U895 (N_895,In_1765,In_975);
xnor U896 (N_896,In_280,In_1310);
xnor U897 (N_897,In_1533,In_1477);
nand U898 (N_898,In_412,In_43);
or U899 (N_899,In_1681,In_937);
nor U900 (N_900,In_1996,In_1183);
or U901 (N_901,In_1394,In_113);
and U902 (N_902,In_503,In_1803);
xor U903 (N_903,In_1928,In_1135);
nor U904 (N_904,In_837,In_154);
or U905 (N_905,In_706,In_1361);
and U906 (N_906,In_1237,In_687);
and U907 (N_907,In_921,In_1458);
nor U908 (N_908,In_226,In_1561);
xnor U909 (N_909,In_15,In_1540);
xnor U910 (N_910,In_671,In_815);
nor U911 (N_911,In_30,In_1622);
or U912 (N_912,In_720,In_694);
nor U913 (N_913,In_789,In_264);
xor U914 (N_914,In_369,In_120);
nand U915 (N_915,In_1709,In_108);
or U916 (N_916,In_1598,In_486);
xnor U917 (N_917,In_470,In_623);
xor U918 (N_918,In_68,In_1890);
nand U919 (N_919,In_1992,In_834);
or U920 (N_920,In_1234,In_1494);
nor U921 (N_921,In_1930,In_409);
or U922 (N_922,In_359,In_1813);
and U923 (N_923,In_1793,In_764);
nor U924 (N_924,In_1041,In_1501);
xnor U925 (N_925,In_1247,In_1250);
nand U926 (N_926,In_270,In_1366);
nand U927 (N_927,In_1442,In_802);
xnor U928 (N_928,In_1724,In_309);
and U929 (N_929,In_673,In_1772);
and U930 (N_930,In_606,In_1570);
nand U931 (N_931,In_1596,In_1756);
nor U932 (N_932,In_1455,In_485);
and U933 (N_933,In_1649,In_997);
or U934 (N_934,In_424,In_319);
nand U935 (N_935,In_897,In_1696);
or U936 (N_936,In_298,In_970);
xor U937 (N_937,In_1137,In_1821);
nor U938 (N_938,In_1707,In_791);
xor U939 (N_939,In_44,In_184);
xor U940 (N_940,In_679,In_1874);
or U941 (N_941,In_1353,In_1037);
nand U942 (N_942,In_1804,In_52);
nand U943 (N_943,In_189,In_119);
nand U944 (N_944,In_1927,In_884);
nor U945 (N_945,In_1621,In_105);
nor U946 (N_946,In_843,In_1474);
xor U947 (N_947,In_944,In_600);
nand U948 (N_948,In_755,In_559);
nor U949 (N_949,In_1519,In_699);
and U950 (N_950,In_1691,In_1839);
or U951 (N_951,In_1690,In_8);
nand U952 (N_952,In_124,In_1328);
xnor U953 (N_953,In_335,In_574);
or U954 (N_954,In_1424,In_1365);
xnor U955 (N_955,In_1232,In_1263);
xor U956 (N_956,In_773,In_704);
and U957 (N_957,In_1679,In_1876);
or U958 (N_958,In_1913,In_354);
and U959 (N_959,In_729,In_1748);
nor U960 (N_960,In_61,In_1431);
or U961 (N_961,In_957,In_1320);
and U962 (N_962,In_418,In_1419);
nor U963 (N_963,In_1434,In_901);
nand U964 (N_964,In_1643,In_882);
and U965 (N_965,In_109,In_224);
xnor U966 (N_966,In_1919,In_216);
xnor U967 (N_967,In_594,In_191);
xor U968 (N_968,In_482,In_1290);
or U969 (N_969,In_1202,In_519);
nand U970 (N_970,In_665,In_238);
nor U971 (N_971,In_320,In_1506);
or U972 (N_972,In_876,In_437);
xnor U973 (N_973,In_1327,In_647);
nor U974 (N_974,In_303,In_10);
nand U975 (N_975,In_122,In_1228);
nor U976 (N_976,In_1942,In_1660);
or U977 (N_977,In_33,In_316);
nor U978 (N_978,In_1770,In_254);
xnor U979 (N_979,In_863,In_659);
xnor U980 (N_980,In_765,In_616);
nor U981 (N_981,In_1987,In_795);
and U982 (N_982,In_1977,In_1049);
or U983 (N_983,In_920,In_1541);
nor U984 (N_984,In_1465,In_1888);
xnor U985 (N_985,In_266,In_851);
or U986 (N_986,In_1510,In_1371);
nand U987 (N_987,In_1589,In_1907);
or U988 (N_988,In_1675,In_1042);
nand U989 (N_989,In_410,In_648);
nor U990 (N_990,In_853,In_176);
xor U991 (N_991,In_1586,In_1423);
nor U992 (N_992,In_281,In_634);
nand U993 (N_993,In_1404,In_507);
and U994 (N_994,In_1133,In_633);
nor U995 (N_995,In_444,In_601);
or U996 (N_996,In_914,In_0);
xor U997 (N_997,In_1329,In_92);
xor U998 (N_998,In_1214,In_1957);
xor U999 (N_999,In_1288,In_1341);
nand U1000 (N_1000,N_249,N_850);
or U1001 (N_1001,N_728,N_558);
xnor U1002 (N_1002,N_654,N_800);
nand U1003 (N_1003,N_910,N_669);
nor U1004 (N_1004,N_582,N_770);
nor U1005 (N_1005,N_356,N_458);
and U1006 (N_1006,N_532,N_312);
and U1007 (N_1007,N_331,N_834);
or U1008 (N_1008,N_391,N_430);
or U1009 (N_1009,N_671,N_417);
and U1010 (N_1010,N_831,N_165);
nor U1011 (N_1011,N_560,N_682);
or U1012 (N_1012,N_970,N_849);
or U1013 (N_1013,N_343,N_824);
and U1014 (N_1014,N_194,N_542);
nand U1015 (N_1015,N_746,N_347);
and U1016 (N_1016,N_647,N_466);
and U1017 (N_1017,N_424,N_315);
nand U1018 (N_1018,N_164,N_118);
nor U1019 (N_1019,N_125,N_620);
or U1020 (N_1020,N_609,N_155);
and U1021 (N_1021,N_179,N_695);
and U1022 (N_1022,N_174,N_392);
nand U1023 (N_1023,N_825,N_998);
and U1024 (N_1024,N_222,N_767);
and U1025 (N_1025,N_461,N_984);
nor U1026 (N_1026,N_758,N_992);
or U1027 (N_1027,N_749,N_148);
nor U1028 (N_1028,N_28,N_205);
nor U1029 (N_1029,N_23,N_862);
and U1030 (N_1030,N_891,N_570);
nor U1031 (N_1031,N_720,N_122);
nand U1032 (N_1032,N_738,N_11);
nand U1033 (N_1033,N_597,N_150);
and U1034 (N_1034,N_324,N_463);
or U1035 (N_1035,N_903,N_261);
and U1036 (N_1036,N_665,N_18);
or U1037 (N_1037,N_655,N_785);
xor U1038 (N_1038,N_224,N_12);
xnor U1039 (N_1039,N_818,N_188);
xor U1040 (N_1040,N_622,N_844);
nand U1041 (N_1041,N_57,N_691);
nand U1042 (N_1042,N_816,N_983);
xor U1043 (N_1043,N_580,N_931);
nand U1044 (N_1044,N_523,N_246);
nor U1045 (N_1045,N_43,N_395);
xor U1046 (N_1046,N_82,N_64);
nor U1047 (N_1047,N_940,N_923);
and U1048 (N_1048,N_83,N_907);
and U1049 (N_1049,N_355,N_928);
nor U1050 (N_1050,N_379,N_81);
or U1051 (N_1051,N_562,N_288);
or U1052 (N_1052,N_846,N_278);
or U1053 (N_1053,N_673,N_555);
nor U1054 (N_1054,N_804,N_988);
or U1055 (N_1055,N_748,N_25);
xor U1056 (N_1056,N_453,N_892);
xnor U1057 (N_1057,N_149,N_27);
and U1058 (N_1058,N_877,N_590);
and U1059 (N_1059,N_740,N_19);
xnor U1060 (N_1060,N_888,N_672);
or U1061 (N_1061,N_185,N_366);
nand U1062 (N_1062,N_163,N_207);
nand U1063 (N_1063,N_668,N_530);
and U1064 (N_1064,N_329,N_566);
nand U1065 (N_1065,N_295,N_635);
or U1066 (N_1066,N_166,N_886);
nor U1067 (N_1067,N_72,N_496);
and U1068 (N_1068,N_629,N_321);
xor U1069 (N_1069,N_994,N_743);
and U1070 (N_1070,N_364,N_779);
nand U1071 (N_1071,N_337,N_821);
or U1072 (N_1072,N_917,N_58);
nand U1073 (N_1073,N_982,N_771);
xor U1074 (N_1074,N_275,N_432);
and U1075 (N_1075,N_349,N_426);
nand U1076 (N_1076,N_946,N_525);
nand U1077 (N_1077,N_652,N_958);
xnor U1078 (N_1078,N_773,N_86);
nor U1079 (N_1079,N_739,N_658);
nor U1080 (N_1080,N_35,N_693);
nand U1081 (N_1081,N_881,N_236);
and U1082 (N_1082,N_156,N_692);
and U1083 (N_1083,N_649,N_414);
xor U1084 (N_1084,N_133,N_536);
nor U1085 (N_1085,N_522,N_814);
or U1086 (N_1086,N_554,N_400);
or U1087 (N_1087,N_833,N_248);
xor U1088 (N_1088,N_240,N_279);
and U1089 (N_1089,N_995,N_911);
or U1090 (N_1090,N_412,N_482);
xor U1091 (N_1091,N_782,N_196);
nand U1092 (N_1092,N_607,N_146);
or U1093 (N_1093,N_679,N_657);
xnor U1094 (N_1094,N_398,N_987);
nand U1095 (N_1095,N_322,N_718);
and U1096 (N_1096,N_380,N_914);
nor U1097 (N_1097,N_500,N_419);
and U1098 (N_1098,N_901,N_713);
and U1099 (N_1099,N_698,N_596);
xor U1100 (N_1100,N_485,N_625);
nor U1101 (N_1101,N_386,N_613);
nor U1102 (N_1102,N_534,N_504);
or U1103 (N_1103,N_896,N_178);
nand U1104 (N_1104,N_587,N_55);
nor U1105 (N_1105,N_884,N_367);
or U1106 (N_1106,N_880,N_66);
and U1107 (N_1107,N_707,N_422);
or U1108 (N_1108,N_553,N_399);
xor U1109 (N_1109,N_368,N_683);
nand U1110 (N_1110,N_722,N_733);
xor U1111 (N_1111,N_611,N_344);
nand U1112 (N_1112,N_448,N_688);
xor U1113 (N_1113,N_650,N_478);
or U1114 (N_1114,N_213,N_203);
xor U1115 (N_1115,N_280,N_798);
nor U1116 (N_1116,N_427,N_599);
and U1117 (N_1117,N_670,N_385);
xnor U1118 (N_1118,N_631,N_703);
and U1119 (N_1119,N_784,N_826);
or U1120 (N_1120,N_169,N_114);
nand U1121 (N_1121,N_702,N_936);
and U1122 (N_1122,N_52,N_215);
nand U1123 (N_1123,N_885,N_853);
or U1124 (N_1124,N_511,N_598);
and U1125 (N_1125,N_787,N_320);
nand U1126 (N_1126,N_841,N_586);
nand U1127 (N_1127,N_193,N_510);
nor U1128 (N_1128,N_492,N_488);
or U1129 (N_1129,N_281,N_745);
nor U1130 (N_1130,N_541,N_709);
xor U1131 (N_1131,N_856,N_131);
xnor U1132 (N_1132,N_699,N_471);
nand U1133 (N_1133,N_381,N_545);
nor U1134 (N_1134,N_479,N_137);
nand U1135 (N_1135,N_232,N_817);
and U1136 (N_1136,N_211,N_128);
and U1137 (N_1137,N_662,N_512);
nand U1138 (N_1138,N_80,N_247);
and U1139 (N_1139,N_859,N_161);
or U1140 (N_1140,N_490,N_108);
and U1141 (N_1141,N_102,N_780);
nor U1142 (N_1142,N_5,N_667);
and U1143 (N_1143,N_2,N_802);
and U1144 (N_1144,N_456,N_666);
nand U1145 (N_1145,N_198,N_34);
nor U1146 (N_1146,N_741,N_302);
and U1147 (N_1147,N_243,N_38);
or U1148 (N_1148,N_450,N_441);
or U1149 (N_1149,N_949,N_483);
nand U1150 (N_1150,N_628,N_84);
xnor U1151 (N_1151,N_228,N_172);
nand U1152 (N_1152,N_291,N_975);
nand U1153 (N_1153,N_956,N_806);
and U1154 (N_1154,N_601,N_934);
xor U1155 (N_1155,N_799,N_990);
nor U1156 (N_1156,N_761,N_362);
or U1157 (N_1157,N_837,N_795);
xor U1158 (N_1158,N_363,N_993);
nor U1159 (N_1159,N_285,N_168);
and U1160 (N_1160,N_209,N_793);
and U1161 (N_1161,N_251,N_869);
and U1162 (N_1162,N_747,N_421);
and U1163 (N_1163,N_835,N_867);
or U1164 (N_1164,N_369,N_332);
nor U1165 (N_1165,N_439,N_565);
xnor U1166 (N_1166,N_933,N_201);
nor U1167 (N_1167,N_696,N_435);
nor U1168 (N_1168,N_348,N_978);
and U1169 (N_1169,N_230,N_516);
nor U1170 (N_1170,N_811,N_572);
nand U1171 (N_1171,N_764,N_687);
nand U1172 (N_1172,N_106,N_78);
and U1173 (N_1173,N_781,N_253);
nand U1174 (N_1174,N_14,N_883);
or U1175 (N_1175,N_100,N_468);
nor U1176 (N_1176,N_95,N_50);
xor U1177 (N_1177,N_723,N_543);
or U1178 (N_1178,N_527,N_508);
xor U1179 (N_1179,N_769,N_897);
nand U1180 (N_1180,N_651,N_403);
xor U1181 (N_1181,N_942,N_415);
xor U1182 (N_1182,N_229,N_845);
and U1183 (N_1183,N_44,N_431);
nand U1184 (N_1184,N_182,N_474);
nor U1185 (N_1185,N_199,N_396);
and U1186 (N_1186,N_751,N_464);
xor U1187 (N_1187,N_305,N_101);
xnor U1188 (N_1188,N_985,N_85);
or U1189 (N_1189,N_88,N_1);
nand U1190 (N_1190,N_204,N_443);
nor U1191 (N_1191,N_955,N_685);
xnor U1192 (N_1192,N_333,N_792);
xnor U1193 (N_1193,N_142,N_971);
or U1194 (N_1194,N_925,N_377);
or U1195 (N_1195,N_328,N_342);
xor U1196 (N_1196,N_216,N_575);
or U1197 (N_1197,N_710,N_812);
nor U1198 (N_1198,N_730,N_96);
nand U1199 (N_1199,N_898,N_56);
nand U1200 (N_1200,N_564,N_53);
nand U1201 (N_1201,N_873,N_346);
and U1202 (N_1202,N_950,N_171);
and U1203 (N_1203,N_308,N_290);
and U1204 (N_1204,N_405,N_581);
nand U1205 (N_1205,N_41,N_531);
and U1206 (N_1206,N_314,N_513);
nand U1207 (N_1207,N_937,N_255);
xnor U1208 (N_1208,N_663,N_929);
or U1209 (N_1209,N_71,N_217);
or U1210 (N_1210,N_518,N_296);
nor U1211 (N_1211,N_98,N_617);
xnor U1212 (N_1212,N_976,N_865);
xor U1213 (N_1213,N_103,N_42);
or U1214 (N_1214,N_621,N_552);
nor U1215 (N_1215,N_449,N_353);
nand U1216 (N_1216,N_220,N_8);
or U1217 (N_1217,N_803,N_231);
or U1218 (N_1218,N_69,N_158);
or U1219 (N_1219,N_105,N_365);
nand U1220 (N_1220,N_538,N_979);
and U1221 (N_1221,N_498,N_729);
nand U1222 (N_1222,N_961,N_828);
nand U1223 (N_1223,N_74,N_31);
xnor U1224 (N_1224,N_571,N_645);
nor U1225 (N_1225,N_537,N_752);
and U1226 (N_1226,N_579,N_547);
and U1227 (N_1227,N_473,N_310);
or U1228 (N_1228,N_943,N_868);
nand U1229 (N_1229,N_476,N_820);
nor U1230 (N_1230,N_775,N_638);
nor U1231 (N_1231,N_912,N_65);
and U1232 (N_1232,N_319,N_813);
and U1233 (N_1233,N_866,N_777);
or U1234 (N_1234,N_339,N_960);
nor U1235 (N_1235,N_115,N_445);
and U1236 (N_1236,N_274,N_964);
nand U1237 (N_1237,N_765,N_766);
nand U1238 (N_1238,N_402,N_890);
nor U1239 (N_1239,N_616,N_16);
nor U1240 (N_1240,N_306,N_551);
or U1241 (N_1241,N_801,N_167);
nor U1242 (N_1242,N_966,N_499);
xnor U1243 (N_1243,N_899,N_848);
or U1244 (N_1244,N_284,N_92);
xnor U1245 (N_1245,N_411,N_953);
xnor U1246 (N_1246,N_875,N_548);
and U1247 (N_1247,N_300,N_89);
nor U1248 (N_1248,N_197,N_134);
and U1249 (N_1249,N_996,N_378);
nand U1250 (N_1250,N_20,N_756);
nand U1251 (N_1251,N_639,N_593);
or U1252 (N_1252,N_352,N_574);
and U1253 (N_1253,N_10,N_0);
or U1254 (N_1254,N_721,N_546);
xnor U1255 (N_1255,N_678,N_797);
nand U1256 (N_1256,N_521,N_726);
nand U1257 (N_1257,N_111,N_21);
or U1258 (N_1258,N_872,N_176);
and U1259 (N_1259,N_939,N_186);
nand U1260 (N_1260,N_47,N_623);
xnor U1261 (N_1261,N_408,N_947);
xor U1262 (N_1262,N_123,N_615);
or U1263 (N_1263,N_874,N_404);
nor U1264 (N_1264,N_59,N_68);
xnor U1265 (N_1265,N_736,N_573);
xnor U1266 (N_1266,N_141,N_762);
nor U1267 (N_1267,N_594,N_79);
xnor U1268 (N_1268,N_282,N_37);
xnor U1269 (N_1269,N_140,N_719);
nand U1270 (N_1270,N_67,N_265);
nand U1271 (N_1271,N_603,N_717);
nor U1272 (N_1272,N_132,N_529);
nor U1273 (N_1273,N_371,N_656);
or U1274 (N_1274,N_429,N_624);
nand U1275 (N_1275,N_535,N_180);
xnor U1276 (N_1276,N_303,N_409);
xor U1277 (N_1277,N_838,N_87);
nand U1278 (N_1278,N_459,N_842);
nand U1279 (N_1279,N_863,N_494);
nand U1280 (N_1280,N_735,N_876);
and U1281 (N_1281,N_653,N_48);
and U1282 (N_1282,N_569,N_641);
or U1283 (N_1283,N_714,N_160);
and U1284 (N_1284,N_840,N_268);
nor U1285 (N_1285,N_602,N_153);
nor U1286 (N_1286,N_577,N_805);
or U1287 (N_1287,N_30,N_906);
nand U1288 (N_1288,N_24,N_920);
nor U1289 (N_1289,N_299,N_588);
or U1290 (N_1290,N_460,N_341);
and U1291 (N_1291,N_823,N_822);
nor U1292 (N_1292,N_452,N_585);
nand U1293 (N_1293,N_786,N_847);
nor U1294 (N_1294,N_918,N_681);
xor U1295 (N_1295,N_212,N_446);
nand U1296 (N_1296,N_152,N_980);
nor U1297 (N_1297,N_472,N_744);
nand U1298 (N_1298,N_237,N_287);
xnor U1299 (N_1299,N_338,N_326);
nor U1300 (N_1300,N_410,N_317);
and U1301 (N_1301,N_245,N_694);
xor U1302 (N_1302,N_304,N_219);
and U1303 (N_1303,N_829,N_286);
and U1304 (N_1304,N_690,N_170);
nand U1305 (N_1305,N_447,N_852);
nand U1306 (N_1306,N_126,N_17);
xnor U1307 (N_1307,N_514,N_680);
xnor U1308 (N_1308,N_659,N_433);
or U1309 (N_1309,N_361,N_894);
and U1310 (N_1310,N_425,N_359);
and U1311 (N_1311,N_605,N_878);
nand U1312 (N_1312,N_908,N_904);
nand U1313 (N_1313,N_94,N_578);
nor U1314 (N_1314,N_854,N_965);
xor U1315 (N_1315,N_388,N_614);
xnor U1316 (N_1316,N_33,N_819);
nand U1317 (N_1317,N_855,N_660);
or U1318 (N_1318,N_619,N_40);
xnor U1319 (N_1319,N_423,N_489);
nand U1320 (N_1320,N_708,N_832);
and U1321 (N_1321,N_794,N_705);
and U1322 (N_1322,N_157,N_484);
or U1323 (N_1323,N_725,N_857);
nor U1324 (N_1324,N_242,N_843);
nand U1325 (N_1325,N_807,N_589);
nor U1326 (N_1326,N_418,N_354);
xnor U1327 (N_1327,N_768,N_632);
xor U1328 (N_1328,N_357,N_241);
and U1329 (N_1329,N_238,N_208);
nor U1330 (N_1330,N_454,N_610);
or U1331 (N_1331,N_393,N_75);
and U1332 (N_1332,N_345,N_351);
and U1333 (N_1333,N_627,N_776);
nor U1334 (N_1334,N_135,N_93);
nor U1335 (N_1335,N_63,N_922);
nor U1336 (N_1336,N_734,N_416);
xnor U1337 (N_1337,N_189,N_307);
and U1338 (N_1338,N_959,N_99);
and U1339 (N_1339,N_675,N_60);
or U1340 (N_1340,N_187,N_376);
xnor U1341 (N_1341,N_384,N_467);
nand U1342 (N_1342,N_154,N_138);
or U1343 (N_1343,N_634,N_259);
nand U1344 (N_1344,N_600,N_495);
nand U1345 (N_1345,N_916,N_120);
xor U1346 (N_1346,N_316,N_390);
xnor U1347 (N_1347,N_151,N_921);
xor U1348 (N_1348,N_202,N_686);
and U1349 (N_1349,N_190,N_113);
nor U1350 (N_1350,N_477,N_962);
nor U1351 (N_1351,N_754,N_475);
and U1352 (N_1352,N_177,N_497);
or U1353 (N_1353,N_774,N_544);
xnor U1354 (N_1354,N_557,N_646);
nor U1355 (N_1355,N_382,N_272);
nand U1356 (N_1356,N_389,N_76);
nor U1357 (N_1357,N_712,N_129);
or U1358 (N_1358,N_62,N_227);
or U1359 (N_1359,N_860,N_206);
nand U1360 (N_1360,N_32,N_977);
nand U1361 (N_1361,N_968,N_591);
nor U1362 (N_1362,N_989,N_526);
xnor U1363 (N_1363,N_277,N_517);
xnor U1364 (N_1364,N_858,N_919);
nor U1365 (N_1365,N_257,N_991);
or U1366 (N_1366,N_250,N_335);
or U1367 (N_1367,N_997,N_791);
or U1368 (N_1368,N_839,N_932);
nand U1369 (N_1369,N_643,N_974);
xnor U1370 (N_1370,N_394,N_13);
nor U1371 (N_1371,N_706,N_372);
xor U1372 (N_1372,N_969,N_294);
or U1373 (N_1373,N_871,N_608);
nand U1374 (N_1374,N_732,N_15);
and U1375 (N_1375,N_935,N_116);
and U1376 (N_1376,N_413,N_271);
nor U1377 (N_1377,N_469,N_505);
xnor U1378 (N_1378,N_273,N_887);
xnor U1379 (N_1379,N_563,N_195);
nand U1380 (N_1380,N_674,N_39);
and U1381 (N_1381,N_254,N_112);
nand U1382 (N_1382,N_436,N_486);
nor U1383 (N_1383,N_963,N_515);
or U1384 (N_1384,N_861,N_926);
nor U1385 (N_1385,N_104,N_130);
nor U1386 (N_1386,N_539,N_124);
xor U1387 (N_1387,N_192,N_815);
and U1388 (N_1388,N_350,N_292);
nand U1389 (N_1389,N_684,N_716);
or U1390 (N_1390,N_986,N_127);
and U1391 (N_1391,N_938,N_759);
nand U1392 (N_1392,N_256,N_3);
xor U1393 (N_1393,N_397,N_298);
nand U1394 (N_1394,N_233,N_642);
nand U1395 (N_1395,N_263,N_509);
and U1396 (N_1396,N_143,N_905);
or U1397 (N_1397,N_900,N_4);
or U1398 (N_1398,N_309,N_550);
xor U1399 (N_1399,N_913,N_51);
and U1400 (N_1400,N_715,N_387);
nor U1401 (N_1401,N_325,N_612);
nor U1402 (N_1402,N_827,N_540);
nand U1403 (N_1403,N_297,N_6);
nand U1404 (N_1404,N_677,N_701);
xor U1405 (N_1405,N_119,N_370);
and U1406 (N_1406,N_221,N_957);
xor U1407 (N_1407,N_270,N_451);
or U1408 (N_1408,N_606,N_864);
or U1409 (N_1409,N_45,N_136);
or U1410 (N_1410,N_336,N_967);
xor U1411 (N_1411,N_9,N_267);
nand U1412 (N_1412,N_311,N_323);
xor U1413 (N_1413,N_70,N_22);
nor U1414 (N_1414,N_258,N_879);
nor U1415 (N_1415,N_533,N_375);
or U1416 (N_1416,N_173,N_301);
nand U1417 (N_1417,N_330,N_465);
nor U1418 (N_1418,N_262,N_561);
or U1419 (N_1419,N_318,N_457);
nor U1420 (N_1420,N_568,N_637);
nor U1421 (N_1421,N_470,N_549);
nor U1422 (N_1422,N_954,N_556);
nor U1423 (N_1423,N_438,N_948);
and U1424 (N_1424,N_358,N_7);
or U1425 (N_1425,N_809,N_783);
nor U1426 (N_1426,N_524,N_97);
xnor U1427 (N_1427,N_944,N_595);
or U1428 (N_1428,N_640,N_895);
nor U1429 (N_1429,N_373,N_491);
and U1430 (N_1430,N_239,N_235);
nand U1431 (N_1431,N_506,N_428);
xnor U1432 (N_1432,N_742,N_147);
nor U1433 (N_1433,N_407,N_117);
nor U1434 (N_1434,N_283,N_727);
and U1435 (N_1435,N_54,N_503);
or U1436 (N_1436,N_440,N_252);
and U1437 (N_1437,N_592,N_401);
or U1438 (N_1438,N_711,N_528);
nand U1439 (N_1439,N_244,N_210);
xnor U1440 (N_1440,N_882,N_162);
nand U1441 (N_1441,N_49,N_90);
or U1442 (N_1442,N_583,N_636);
nor U1443 (N_1443,N_851,N_260);
nand U1444 (N_1444,N_648,N_406);
or U1445 (N_1445,N_360,N_893);
and U1446 (N_1446,N_755,N_234);
nor U1447 (N_1447,N_915,N_214);
and U1448 (N_1448,N_999,N_633);
nand U1449 (N_1449,N_788,N_289);
xor U1450 (N_1450,N_789,N_313);
or U1451 (N_1451,N_374,N_481);
xor U1452 (N_1452,N_973,N_644);
nor U1453 (N_1453,N_36,N_808);
xor U1454 (N_1454,N_200,N_559);
nor U1455 (N_1455,N_661,N_731);
or U1456 (N_1456,N_704,N_576);
and U1457 (N_1457,N_264,N_327);
nor U1458 (N_1458,N_753,N_225);
and U1459 (N_1459,N_29,N_909);
xor U1460 (N_1460,N_760,N_226);
or U1461 (N_1461,N_266,N_145);
and U1462 (N_1462,N_630,N_269);
and U1463 (N_1463,N_383,N_757);
xor U1464 (N_1464,N_502,N_689);
nand U1465 (N_1465,N_889,N_972);
nor U1466 (N_1466,N_750,N_737);
or U1467 (N_1467,N_724,N_184);
or U1468 (N_1468,N_444,N_772);
xor U1469 (N_1469,N_437,N_697);
and U1470 (N_1470,N_434,N_191);
nor U1471 (N_1471,N_941,N_46);
nand U1472 (N_1472,N_110,N_618);
or U1473 (N_1473,N_664,N_77);
nor U1474 (N_1474,N_501,N_924);
xnor U1475 (N_1475,N_626,N_836);
or U1476 (N_1476,N_507,N_73);
and U1477 (N_1477,N_293,N_159);
and U1478 (N_1478,N_420,N_810);
xnor U1479 (N_1479,N_830,N_520);
nor U1480 (N_1480,N_763,N_790);
or U1481 (N_1481,N_567,N_584);
nor U1482 (N_1482,N_778,N_175);
and U1483 (N_1483,N_870,N_442);
nand U1484 (N_1484,N_796,N_144);
nand U1485 (N_1485,N_952,N_462);
xnor U1486 (N_1486,N_676,N_700);
and U1487 (N_1487,N_181,N_945);
and U1488 (N_1488,N_223,N_183);
or U1489 (N_1489,N_493,N_109);
or U1490 (N_1490,N_480,N_61);
nor U1491 (N_1491,N_121,N_276);
or U1492 (N_1492,N_951,N_218);
xnor U1493 (N_1493,N_487,N_930);
or U1494 (N_1494,N_107,N_604);
nand U1495 (N_1495,N_91,N_340);
nand U1496 (N_1496,N_139,N_334);
nor U1497 (N_1497,N_981,N_902);
nor U1498 (N_1498,N_927,N_519);
nor U1499 (N_1499,N_455,N_26);
xor U1500 (N_1500,N_927,N_31);
nand U1501 (N_1501,N_937,N_749);
nand U1502 (N_1502,N_128,N_971);
nor U1503 (N_1503,N_271,N_593);
nor U1504 (N_1504,N_228,N_380);
nand U1505 (N_1505,N_337,N_971);
nand U1506 (N_1506,N_319,N_323);
xnor U1507 (N_1507,N_819,N_908);
nor U1508 (N_1508,N_793,N_411);
nor U1509 (N_1509,N_376,N_823);
nor U1510 (N_1510,N_172,N_592);
nor U1511 (N_1511,N_145,N_287);
xor U1512 (N_1512,N_314,N_183);
or U1513 (N_1513,N_612,N_584);
and U1514 (N_1514,N_386,N_848);
and U1515 (N_1515,N_4,N_426);
nand U1516 (N_1516,N_768,N_7);
nor U1517 (N_1517,N_517,N_17);
nor U1518 (N_1518,N_304,N_757);
or U1519 (N_1519,N_10,N_172);
nor U1520 (N_1520,N_767,N_519);
xnor U1521 (N_1521,N_593,N_891);
or U1522 (N_1522,N_616,N_955);
and U1523 (N_1523,N_826,N_333);
nand U1524 (N_1524,N_880,N_907);
or U1525 (N_1525,N_391,N_51);
or U1526 (N_1526,N_347,N_79);
or U1527 (N_1527,N_356,N_308);
nand U1528 (N_1528,N_997,N_159);
and U1529 (N_1529,N_957,N_316);
nand U1530 (N_1530,N_200,N_965);
nor U1531 (N_1531,N_708,N_904);
nand U1532 (N_1532,N_936,N_31);
xnor U1533 (N_1533,N_164,N_553);
xnor U1534 (N_1534,N_381,N_674);
nand U1535 (N_1535,N_335,N_894);
xnor U1536 (N_1536,N_422,N_125);
or U1537 (N_1537,N_805,N_732);
nor U1538 (N_1538,N_592,N_849);
or U1539 (N_1539,N_107,N_557);
nor U1540 (N_1540,N_342,N_496);
nand U1541 (N_1541,N_820,N_71);
nor U1542 (N_1542,N_628,N_844);
and U1543 (N_1543,N_927,N_43);
nor U1544 (N_1544,N_62,N_718);
nor U1545 (N_1545,N_66,N_189);
xor U1546 (N_1546,N_650,N_987);
xnor U1547 (N_1547,N_459,N_859);
xor U1548 (N_1548,N_572,N_955);
or U1549 (N_1549,N_458,N_8);
nand U1550 (N_1550,N_860,N_976);
and U1551 (N_1551,N_571,N_753);
xnor U1552 (N_1552,N_188,N_170);
xor U1553 (N_1553,N_245,N_408);
or U1554 (N_1554,N_917,N_361);
and U1555 (N_1555,N_326,N_671);
nand U1556 (N_1556,N_829,N_871);
and U1557 (N_1557,N_648,N_230);
or U1558 (N_1558,N_119,N_318);
and U1559 (N_1559,N_136,N_737);
xor U1560 (N_1560,N_813,N_620);
or U1561 (N_1561,N_544,N_920);
nor U1562 (N_1562,N_478,N_745);
xor U1563 (N_1563,N_216,N_595);
nand U1564 (N_1564,N_89,N_977);
and U1565 (N_1565,N_976,N_796);
or U1566 (N_1566,N_818,N_59);
and U1567 (N_1567,N_693,N_501);
and U1568 (N_1568,N_185,N_468);
or U1569 (N_1569,N_797,N_296);
nand U1570 (N_1570,N_445,N_871);
or U1571 (N_1571,N_23,N_751);
or U1572 (N_1572,N_180,N_401);
nand U1573 (N_1573,N_947,N_757);
or U1574 (N_1574,N_695,N_978);
xnor U1575 (N_1575,N_795,N_788);
nor U1576 (N_1576,N_820,N_659);
nor U1577 (N_1577,N_311,N_875);
xnor U1578 (N_1578,N_368,N_412);
and U1579 (N_1579,N_515,N_1);
and U1580 (N_1580,N_140,N_668);
nor U1581 (N_1581,N_199,N_599);
or U1582 (N_1582,N_870,N_558);
or U1583 (N_1583,N_336,N_270);
and U1584 (N_1584,N_927,N_619);
nand U1585 (N_1585,N_229,N_326);
xnor U1586 (N_1586,N_542,N_560);
and U1587 (N_1587,N_600,N_506);
nand U1588 (N_1588,N_478,N_202);
nor U1589 (N_1589,N_774,N_422);
xor U1590 (N_1590,N_731,N_220);
xor U1591 (N_1591,N_306,N_858);
nand U1592 (N_1592,N_687,N_57);
xnor U1593 (N_1593,N_557,N_974);
xnor U1594 (N_1594,N_408,N_608);
xnor U1595 (N_1595,N_766,N_379);
nand U1596 (N_1596,N_165,N_76);
nand U1597 (N_1597,N_786,N_618);
nand U1598 (N_1598,N_201,N_102);
or U1599 (N_1599,N_86,N_378);
xnor U1600 (N_1600,N_733,N_288);
nor U1601 (N_1601,N_899,N_491);
xnor U1602 (N_1602,N_467,N_224);
or U1603 (N_1603,N_247,N_630);
xor U1604 (N_1604,N_146,N_886);
xor U1605 (N_1605,N_533,N_471);
nand U1606 (N_1606,N_651,N_399);
and U1607 (N_1607,N_659,N_237);
or U1608 (N_1608,N_486,N_670);
or U1609 (N_1609,N_857,N_919);
nor U1610 (N_1610,N_854,N_765);
and U1611 (N_1611,N_464,N_549);
or U1612 (N_1612,N_365,N_94);
nor U1613 (N_1613,N_110,N_257);
nand U1614 (N_1614,N_129,N_48);
nor U1615 (N_1615,N_840,N_527);
xor U1616 (N_1616,N_429,N_345);
nand U1617 (N_1617,N_285,N_287);
and U1618 (N_1618,N_676,N_453);
nor U1619 (N_1619,N_548,N_140);
and U1620 (N_1620,N_813,N_725);
nand U1621 (N_1621,N_189,N_521);
nand U1622 (N_1622,N_883,N_761);
and U1623 (N_1623,N_969,N_928);
nor U1624 (N_1624,N_377,N_756);
xor U1625 (N_1625,N_442,N_880);
nor U1626 (N_1626,N_302,N_452);
and U1627 (N_1627,N_625,N_821);
nand U1628 (N_1628,N_432,N_269);
or U1629 (N_1629,N_732,N_919);
xnor U1630 (N_1630,N_161,N_423);
nand U1631 (N_1631,N_928,N_424);
nor U1632 (N_1632,N_521,N_72);
and U1633 (N_1633,N_937,N_34);
and U1634 (N_1634,N_244,N_966);
or U1635 (N_1635,N_998,N_185);
nor U1636 (N_1636,N_105,N_902);
nor U1637 (N_1637,N_953,N_767);
nor U1638 (N_1638,N_188,N_590);
nand U1639 (N_1639,N_121,N_222);
and U1640 (N_1640,N_126,N_380);
nor U1641 (N_1641,N_185,N_801);
and U1642 (N_1642,N_921,N_952);
nand U1643 (N_1643,N_572,N_726);
xor U1644 (N_1644,N_895,N_24);
nand U1645 (N_1645,N_595,N_10);
and U1646 (N_1646,N_259,N_877);
nand U1647 (N_1647,N_330,N_804);
xor U1648 (N_1648,N_551,N_470);
nand U1649 (N_1649,N_346,N_109);
xor U1650 (N_1650,N_563,N_393);
nand U1651 (N_1651,N_869,N_560);
or U1652 (N_1652,N_256,N_642);
xnor U1653 (N_1653,N_688,N_416);
and U1654 (N_1654,N_703,N_740);
xor U1655 (N_1655,N_611,N_251);
xor U1656 (N_1656,N_985,N_322);
nand U1657 (N_1657,N_135,N_934);
nor U1658 (N_1658,N_157,N_408);
nand U1659 (N_1659,N_801,N_766);
or U1660 (N_1660,N_699,N_974);
nor U1661 (N_1661,N_312,N_327);
nand U1662 (N_1662,N_266,N_940);
nor U1663 (N_1663,N_286,N_798);
or U1664 (N_1664,N_908,N_439);
nor U1665 (N_1665,N_741,N_742);
nor U1666 (N_1666,N_713,N_37);
or U1667 (N_1667,N_531,N_835);
and U1668 (N_1668,N_564,N_207);
nor U1669 (N_1669,N_544,N_272);
xnor U1670 (N_1670,N_919,N_381);
nor U1671 (N_1671,N_462,N_1);
or U1672 (N_1672,N_931,N_364);
nor U1673 (N_1673,N_567,N_879);
xor U1674 (N_1674,N_783,N_357);
nand U1675 (N_1675,N_31,N_45);
nand U1676 (N_1676,N_814,N_202);
xor U1677 (N_1677,N_0,N_433);
nand U1678 (N_1678,N_253,N_618);
or U1679 (N_1679,N_927,N_865);
nor U1680 (N_1680,N_487,N_665);
and U1681 (N_1681,N_489,N_305);
and U1682 (N_1682,N_113,N_839);
and U1683 (N_1683,N_239,N_736);
or U1684 (N_1684,N_751,N_727);
and U1685 (N_1685,N_267,N_504);
nor U1686 (N_1686,N_530,N_368);
and U1687 (N_1687,N_176,N_540);
nand U1688 (N_1688,N_361,N_945);
nand U1689 (N_1689,N_138,N_81);
and U1690 (N_1690,N_753,N_889);
xnor U1691 (N_1691,N_924,N_937);
nand U1692 (N_1692,N_578,N_155);
or U1693 (N_1693,N_531,N_969);
nor U1694 (N_1694,N_355,N_436);
or U1695 (N_1695,N_756,N_363);
nand U1696 (N_1696,N_267,N_646);
nand U1697 (N_1697,N_838,N_837);
and U1698 (N_1698,N_989,N_63);
nand U1699 (N_1699,N_996,N_461);
and U1700 (N_1700,N_572,N_591);
or U1701 (N_1701,N_775,N_334);
xnor U1702 (N_1702,N_255,N_755);
xnor U1703 (N_1703,N_479,N_46);
nor U1704 (N_1704,N_308,N_235);
xnor U1705 (N_1705,N_449,N_142);
and U1706 (N_1706,N_797,N_782);
nand U1707 (N_1707,N_892,N_685);
nand U1708 (N_1708,N_627,N_316);
nor U1709 (N_1709,N_8,N_414);
or U1710 (N_1710,N_598,N_251);
nand U1711 (N_1711,N_807,N_859);
or U1712 (N_1712,N_701,N_724);
and U1713 (N_1713,N_895,N_701);
and U1714 (N_1714,N_960,N_940);
nor U1715 (N_1715,N_836,N_586);
or U1716 (N_1716,N_798,N_89);
xor U1717 (N_1717,N_586,N_453);
or U1718 (N_1718,N_470,N_31);
and U1719 (N_1719,N_405,N_565);
nand U1720 (N_1720,N_227,N_728);
nand U1721 (N_1721,N_186,N_362);
xnor U1722 (N_1722,N_543,N_18);
nor U1723 (N_1723,N_401,N_728);
nand U1724 (N_1724,N_401,N_764);
and U1725 (N_1725,N_971,N_713);
xor U1726 (N_1726,N_595,N_447);
xor U1727 (N_1727,N_420,N_958);
or U1728 (N_1728,N_354,N_372);
and U1729 (N_1729,N_880,N_380);
xnor U1730 (N_1730,N_505,N_478);
and U1731 (N_1731,N_993,N_388);
nor U1732 (N_1732,N_296,N_898);
xor U1733 (N_1733,N_978,N_555);
nor U1734 (N_1734,N_896,N_676);
and U1735 (N_1735,N_62,N_342);
or U1736 (N_1736,N_922,N_692);
or U1737 (N_1737,N_0,N_986);
nand U1738 (N_1738,N_216,N_685);
xor U1739 (N_1739,N_958,N_827);
or U1740 (N_1740,N_514,N_405);
nor U1741 (N_1741,N_734,N_806);
or U1742 (N_1742,N_21,N_848);
or U1743 (N_1743,N_756,N_244);
nand U1744 (N_1744,N_194,N_33);
nor U1745 (N_1745,N_637,N_232);
nor U1746 (N_1746,N_271,N_269);
or U1747 (N_1747,N_811,N_315);
xnor U1748 (N_1748,N_191,N_624);
xnor U1749 (N_1749,N_41,N_598);
nand U1750 (N_1750,N_254,N_156);
or U1751 (N_1751,N_697,N_678);
xor U1752 (N_1752,N_517,N_338);
nor U1753 (N_1753,N_674,N_281);
nand U1754 (N_1754,N_512,N_525);
xor U1755 (N_1755,N_66,N_79);
and U1756 (N_1756,N_827,N_331);
nand U1757 (N_1757,N_734,N_579);
and U1758 (N_1758,N_398,N_971);
and U1759 (N_1759,N_331,N_688);
nor U1760 (N_1760,N_875,N_221);
nand U1761 (N_1761,N_648,N_494);
or U1762 (N_1762,N_646,N_634);
or U1763 (N_1763,N_774,N_704);
and U1764 (N_1764,N_712,N_294);
nand U1765 (N_1765,N_347,N_560);
nor U1766 (N_1766,N_980,N_396);
nor U1767 (N_1767,N_557,N_229);
or U1768 (N_1768,N_858,N_512);
or U1769 (N_1769,N_877,N_685);
xnor U1770 (N_1770,N_101,N_58);
and U1771 (N_1771,N_336,N_278);
xor U1772 (N_1772,N_588,N_405);
xor U1773 (N_1773,N_909,N_178);
nor U1774 (N_1774,N_61,N_320);
xor U1775 (N_1775,N_730,N_558);
and U1776 (N_1776,N_238,N_339);
xor U1777 (N_1777,N_856,N_481);
nand U1778 (N_1778,N_742,N_702);
or U1779 (N_1779,N_819,N_453);
and U1780 (N_1780,N_721,N_398);
or U1781 (N_1781,N_393,N_461);
or U1782 (N_1782,N_759,N_823);
nor U1783 (N_1783,N_828,N_793);
or U1784 (N_1784,N_328,N_671);
and U1785 (N_1785,N_732,N_512);
nand U1786 (N_1786,N_217,N_89);
xor U1787 (N_1787,N_478,N_33);
nor U1788 (N_1788,N_371,N_789);
nand U1789 (N_1789,N_733,N_172);
xnor U1790 (N_1790,N_986,N_926);
and U1791 (N_1791,N_275,N_582);
xnor U1792 (N_1792,N_36,N_707);
xnor U1793 (N_1793,N_992,N_626);
and U1794 (N_1794,N_76,N_973);
and U1795 (N_1795,N_686,N_544);
or U1796 (N_1796,N_165,N_554);
and U1797 (N_1797,N_221,N_120);
nor U1798 (N_1798,N_377,N_458);
nand U1799 (N_1799,N_623,N_532);
or U1800 (N_1800,N_327,N_384);
nand U1801 (N_1801,N_535,N_553);
xnor U1802 (N_1802,N_293,N_617);
xnor U1803 (N_1803,N_39,N_943);
xnor U1804 (N_1804,N_649,N_380);
nor U1805 (N_1805,N_869,N_85);
and U1806 (N_1806,N_633,N_136);
nand U1807 (N_1807,N_606,N_683);
and U1808 (N_1808,N_943,N_347);
xnor U1809 (N_1809,N_323,N_789);
nand U1810 (N_1810,N_171,N_664);
nor U1811 (N_1811,N_845,N_535);
nand U1812 (N_1812,N_132,N_611);
nand U1813 (N_1813,N_269,N_743);
nor U1814 (N_1814,N_409,N_717);
xor U1815 (N_1815,N_235,N_627);
or U1816 (N_1816,N_32,N_570);
xor U1817 (N_1817,N_107,N_823);
or U1818 (N_1818,N_355,N_609);
and U1819 (N_1819,N_719,N_999);
nand U1820 (N_1820,N_356,N_90);
nor U1821 (N_1821,N_9,N_257);
and U1822 (N_1822,N_530,N_477);
or U1823 (N_1823,N_127,N_676);
nor U1824 (N_1824,N_593,N_396);
or U1825 (N_1825,N_394,N_909);
nor U1826 (N_1826,N_962,N_135);
xor U1827 (N_1827,N_764,N_259);
xor U1828 (N_1828,N_161,N_836);
or U1829 (N_1829,N_930,N_688);
nand U1830 (N_1830,N_253,N_664);
xor U1831 (N_1831,N_837,N_299);
nor U1832 (N_1832,N_600,N_894);
xnor U1833 (N_1833,N_817,N_272);
or U1834 (N_1834,N_925,N_744);
or U1835 (N_1835,N_678,N_767);
nor U1836 (N_1836,N_548,N_29);
nor U1837 (N_1837,N_203,N_642);
and U1838 (N_1838,N_37,N_79);
nand U1839 (N_1839,N_429,N_275);
and U1840 (N_1840,N_112,N_792);
nor U1841 (N_1841,N_371,N_802);
nand U1842 (N_1842,N_714,N_936);
or U1843 (N_1843,N_519,N_893);
or U1844 (N_1844,N_756,N_17);
nor U1845 (N_1845,N_552,N_788);
nor U1846 (N_1846,N_652,N_310);
xnor U1847 (N_1847,N_786,N_933);
and U1848 (N_1848,N_391,N_828);
nand U1849 (N_1849,N_989,N_114);
nand U1850 (N_1850,N_253,N_21);
nor U1851 (N_1851,N_353,N_576);
xnor U1852 (N_1852,N_124,N_403);
nor U1853 (N_1853,N_509,N_317);
or U1854 (N_1854,N_465,N_840);
or U1855 (N_1855,N_292,N_474);
nor U1856 (N_1856,N_167,N_468);
nor U1857 (N_1857,N_362,N_663);
nor U1858 (N_1858,N_616,N_274);
and U1859 (N_1859,N_111,N_386);
xnor U1860 (N_1860,N_579,N_890);
nor U1861 (N_1861,N_569,N_181);
and U1862 (N_1862,N_670,N_569);
or U1863 (N_1863,N_50,N_343);
and U1864 (N_1864,N_602,N_75);
nand U1865 (N_1865,N_253,N_431);
nor U1866 (N_1866,N_379,N_593);
xor U1867 (N_1867,N_962,N_217);
or U1868 (N_1868,N_952,N_384);
xor U1869 (N_1869,N_688,N_328);
nand U1870 (N_1870,N_827,N_121);
xnor U1871 (N_1871,N_12,N_35);
nand U1872 (N_1872,N_287,N_788);
or U1873 (N_1873,N_930,N_414);
and U1874 (N_1874,N_149,N_900);
and U1875 (N_1875,N_149,N_726);
nor U1876 (N_1876,N_212,N_915);
nand U1877 (N_1877,N_672,N_518);
nor U1878 (N_1878,N_694,N_964);
nor U1879 (N_1879,N_902,N_514);
or U1880 (N_1880,N_198,N_227);
xnor U1881 (N_1881,N_575,N_72);
xor U1882 (N_1882,N_824,N_294);
or U1883 (N_1883,N_290,N_445);
nor U1884 (N_1884,N_973,N_677);
and U1885 (N_1885,N_525,N_344);
nor U1886 (N_1886,N_89,N_301);
nor U1887 (N_1887,N_745,N_19);
and U1888 (N_1888,N_778,N_577);
nor U1889 (N_1889,N_844,N_169);
nand U1890 (N_1890,N_773,N_914);
or U1891 (N_1891,N_228,N_726);
and U1892 (N_1892,N_710,N_282);
nor U1893 (N_1893,N_934,N_368);
or U1894 (N_1894,N_688,N_514);
nor U1895 (N_1895,N_157,N_205);
nor U1896 (N_1896,N_153,N_151);
nand U1897 (N_1897,N_868,N_535);
nor U1898 (N_1898,N_652,N_996);
xnor U1899 (N_1899,N_750,N_591);
or U1900 (N_1900,N_873,N_852);
xor U1901 (N_1901,N_532,N_558);
nand U1902 (N_1902,N_53,N_221);
nand U1903 (N_1903,N_495,N_764);
nor U1904 (N_1904,N_143,N_835);
nor U1905 (N_1905,N_559,N_500);
and U1906 (N_1906,N_821,N_122);
or U1907 (N_1907,N_787,N_559);
or U1908 (N_1908,N_213,N_123);
or U1909 (N_1909,N_592,N_16);
nor U1910 (N_1910,N_869,N_848);
nand U1911 (N_1911,N_151,N_547);
nor U1912 (N_1912,N_161,N_203);
xnor U1913 (N_1913,N_933,N_339);
nand U1914 (N_1914,N_477,N_353);
xor U1915 (N_1915,N_745,N_397);
xnor U1916 (N_1916,N_296,N_960);
and U1917 (N_1917,N_385,N_964);
xor U1918 (N_1918,N_95,N_252);
xnor U1919 (N_1919,N_395,N_5);
nand U1920 (N_1920,N_303,N_292);
nor U1921 (N_1921,N_110,N_877);
nand U1922 (N_1922,N_33,N_812);
nor U1923 (N_1923,N_911,N_336);
nand U1924 (N_1924,N_679,N_135);
and U1925 (N_1925,N_614,N_390);
or U1926 (N_1926,N_165,N_328);
nand U1927 (N_1927,N_786,N_884);
or U1928 (N_1928,N_845,N_509);
and U1929 (N_1929,N_771,N_806);
xnor U1930 (N_1930,N_217,N_681);
nor U1931 (N_1931,N_269,N_539);
nand U1932 (N_1932,N_669,N_123);
xnor U1933 (N_1933,N_308,N_392);
nor U1934 (N_1934,N_381,N_176);
xor U1935 (N_1935,N_527,N_629);
nand U1936 (N_1936,N_905,N_909);
nand U1937 (N_1937,N_2,N_594);
and U1938 (N_1938,N_799,N_4);
and U1939 (N_1939,N_876,N_711);
and U1940 (N_1940,N_379,N_574);
nand U1941 (N_1941,N_669,N_745);
nor U1942 (N_1942,N_368,N_863);
and U1943 (N_1943,N_805,N_145);
and U1944 (N_1944,N_219,N_357);
xor U1945 (N_1945,N_681,N_518);
xor U1946 (N_1946,N_695,N_900);
nand U1947 (N_1947,N_802,N_847);
xnor U1948 (N_1948,N_928,N_971);
nor U1949 (N_1949,N_933,N_290);
and U1950 (N_1950,N_665,N_153);
xor U1951 (N_1951,N_589,N_596);
and U1952 (N_1952,N_890,N_280);
nor U1953 (N_1953,N_131,N_82);
xnor U1954 (N_1954,N_866,N_242);
nand U1955 (N_1955,N_22,N_988);
nand U1956 (N_1956,N_589,N_926);
or U1957 (N_1957,N_57,N_621);
nor U1958 (N_1958,N_406,N_317);
nor U1959 (N_1959,N_284,N_866);
xor U1960 (N_1960,N_926,N_387);
and U1961 (N_1961,N_984,N_409);
and U1962 (N_1962,N_844,N_496);
xor U1963 (N_1963,N_63,N_897);
and U1964 (N_1964,N_347,N_56);
nor U1965 (N_1965,N_204,N_620);
xor U1966 (N_1966,N_11,N_443);
xnor U1967 (N_1967,N_136,N_506);
xor U1968 (N_1968,N_132,N_432);
or U1969 (N_1969,N_96,N_200);
nand U1970 (N_1970,N_743,N_199);
and U1971 (N_1971,N_548,N_148);
nand U1972 (N_1972,N_777,N_929);
or U1973 (N_1973,N_700,N_977);
nor U1974 (N_1974,N_502,N_282);
nand U1975 (N_1975,N_50,N_537);
nor U1976 (N_1976,N_968,N_986);
nand U1977 (N_1977,N_279,N_484);
or U1978 (N_1978,N_36,N_31);
nand U1979 (N_1979,N_77,N_411);
nor U1980 (N_1980,N_317,N_691);
or U1981 (N_1981,N_998,N_456);
and U1982 (N_1982,N_753,N_856);
nor U1983 (N_1983,N_937,N_881);
or U1984 (N_1984,N_891,N_513);
and U1985 (N_1985,N_768,N_725);
or U1986 (N_1986,N_899,N_404);
nand U1987 (N_1987,N_182,N_252);
xor U1988 (N_1988,N_291,N_82);
nand U1989 (N_1989,N_139,N_225);
or U1990 (N_1990,N_612,N_960);
nand U1991 (N_1991,N_714,N_603);
or U1992 (N_1992,N_302,N_137);
or U1993 (N_1993,N_984,N_502);
xor U1994 (N_1994,N_595,N_167);
and U1995 (N_1995,N_805,N_516);
and U1996 (N_1996,N_950,N_460);
or U1997 (N_1997,N_934,N_777);
nand U1998 (N_1998,N_287,N_215);
nand U1999 (N_1999,N_460,N_650);
or U2000 (N_2000,N_1115,N_1464);
xor U2001 (N_2001,N_1881,N_1357);
nor U2002 (N_2002,N_1310,N_1356);
nand U2003 (N_2003,N_1706,N_1619);
xnor U2004 (N_2004,N_1034,N_1102);
nor U2005 (N_2005,N_1506,N_1334);
and U2006 (N_2006,N_1387,N_1795);
xnor U2007 (N_2007,N_1892,N_1610);
and U2008 (N_2008,N_1197,N_1308);
nand U2009 (N_2009,N_1471,N_1518);
nor U2010 (N_2010,N_1755,N_1317);
xnor U2011 (N_2011,N_1072,N_1523);
xnor U2012 (N_2012,N_1534,N_1314);
nor U2013 (N_2013,N_1887,N_1675);
nand U2014 (N_2014,N_1753,N_1634);
nand U2015 (N_2015,N_1535,N_1039);
nand U2016 (N_2016,N_1407,N_1873);
xnor U2017 (N_2017,N_1144,N_1744);
and U2018 (N_2018,N_1950,N_1816);
nor U2019 (N_2019,N_1544,N_1394);
or U2020 (N_2020,N_1882,N_1424);
xor U2021 (N_2021,N_1948,N_1525);
and U2022 (N_2022,N_1746,N_1351);
nor U2023 (N_2023,N_1078,N_1332);
or U2024 (N_2024,N_1716,N_1161);
and U2025 (N_2025,N_1999,N_1509);
nand U2026 (N_2026,N_1839,N_1520);
nand U2027 (N_2027,N_1925,N_1994);
xnor U2028 (N_2028,N_1231,N_1673);
and U2029 (N_2029,N_1081,N_1902);
xnor U2030 (N_2030,N_1597,N_1215);
nand U2031 (N_2031,N_1353,N_1193);
xor U2032 (N_2032,N_1777,N_1549);
nand U2033 (N_2033,N_1919,N_1167);
nand U2034 (N_2034,N_1604,N_1896);
nand U2035 (N_2035,N_1048,N_1089);
nand U2036 (N_2036,N_1488,N_1561);
nor U2037 (N_2037,N_1894,N_1271);
nor U2038 (N_2038,N_1517,N_1642);
and U2039 (N_2039,N_1079,N_1192);
xnor U2040 (N_2040,N_1715,N_1934);
or U2041 (N_2041,N_1758,N_1773);
xnor U2042 (N_2042,N_1339,N_1216);
nor U2043 (N_2043,N_1043,N_1020);
or U2044 (N_2044,N_1587,N_1009);
nor U2045 (N_2045,N_1266,N_1275);
nand U2046 (N_2046,N_1786,N_1166);
nand U2047 (N_2047,N_1062,N_1131);
or U2048 (N_2048,N_1446,N_1451);
nor U2049 (N_2049,N_1309,N_1973);
or U2050 (N_2050,N_1616,N_1124);
nor U2051 (N_2051,N_1123,N_1729);
and U2052 (N_2052,N_1511,N_1465);
and U2053 (N_2053,N_1472,N_1190);
nor U2054 (N_2054,N_1432,N_1418);
nand U2055 (N_2055,N_1319,N_1686);
or U2056 (N_2056,N_1248,N_1836);
xor U2057 (N_2057,N_1297,N_1987);
and U2058 (N_2058,N_1855,N_1083);
and U2059 (N_2059,N_1195,N_1459);
nand U2060 (N_2060,N_1321,N_1515);
or U2061 (N_2061,N_1212,N_1402);
and U2062 (N_2062,N_1390,N_1245);
nand U2063 (N_2063,N_1347,N_1117);
nor U2064 (N_2064,N_1552,N_1848);
or U2065 (N_2065,N_1875,N_1400);
nor U2066 (N_2066,N_1947,N_1110);
or U2067 (N_2067,N_1200,N_1572);
xor U2068 (N_2068,N_1399,N_1198);
or U2069 (N_2069,N_1186,N_1533);
nor U2070 (N_2070,N_1085,N_1447);
and U2071 (N_2071,N_1139,N_1766);
nor U2072 (N_2072,N_1921,N_1255);
or U2073 (N_2073,N_1132,N_1305);
or U2074 (N_2074,N_1259,N_1141);
and U2075 (N_2075,N_1538,N_1933);
nor U2076 (N_2076,N_1752,N_1573);
nand U2077 (N_2077,N_1799,N_1431);
or U2078 (N_2078,N_1863,N_1218);
nor U2079 (N_2079,N_1233,N_1364);
nand U2080 (N_2080,N_1564,N_1981);
nand U2081 (N_2081,N_1098,N_1494);
nor U2082 (N_2082,N_1849,N_1907);
nor U2083 (N_2083,N_1286,N_1016);
and U2084 (N_2084,N_1809,N_1363);
nand U2085 (N_2085,N_1213,N_1513);
nand U2086 (N_2086,N_1789,N_1926);
nand U2087 (N_2087,N_1700,N_1938);
and U2088 (N_2088,N_1965,N_1852);
or U2089 (N_2089,N_1183,N_1064);
nand U2090 (N_2090,N_1847,N_1895);
xor U2091 (N_2091,N_1159,N_1874);
nor U2092 (N_2092,N_1976,N_1268);
xnor U2093 (N_2093,N_1282,N_1893);
and U2094 (N_2094,N_1983,N_1223);
nor U2095 (N_2095,N_1270,N_1949);
nor U2096 (N_2096,N_1810,N_1140);
and U2097 (N_2097,N_1194,N_1612);
nand U2098 (N_2098,N_1519,N_1466);
and U2099 (N_2099,N_1898,N_1316);
or U2100 (N_2100,N_1011,N_1367);
or U2101 (N_2101,N_1550,N_1574);
and U2102 (N_2102,N_1929,N_1204);
xnor U2103 (N_2103,N_1804,N_1137);
nand U2104 (N_2104,N_1916,N_1555);
nand U2105 (N_2105,N_1236,N_1001);
and U2106 (N_2106,N_1554,N_1829);
and U2107 (N_2107,N_1486,N_1153);
nor U2108 (N_2108,N_1412,N_1005);
nand U2109 (N_2109,N_1253,N_1670);
and U2110 (N_2110,N_1735,N_1671);
nor U2111 (N_2111,N_1207,N_1764);
nand U2112 (N_2112,N_1485,N_1570);
or U2113 (N_2113,N_1521,N_1802);
and U2114 (N_2114,N_1010,N_1608);
nand U2115 (N_2115,N_1522,N_1780);
nand U2116 (N_2116,N_1368,N_1313);
or U2117 (N_2117,N_1172,N_1638);
xor U2118 (N_2118,N_1743,N_1229);
nor U2119 (N_2119,N_1073,N_1811);
and U2120 (N_2120,N_1120,N_1346);
nand U2121 (N_2121,N_1427,N_1377);
xor U2122 (N_2122,N_1345,N_1644);
nand U2123 (N_2123,N_1021,N_1258);
xor U2124 (N_2124,N_1737,N_1489);
nand U2125 (N_2125,N_1329,N_1684);
or U2126 (N_2126,N_1415,N_1196);
and U2127 (N_2127,N_1374,N_1910);
xor U2128 (N_2128,N_1114,N_1033);
and U2129 (N_2129,N_1868,N_1813);
or U2130 (N_2130,N_1458,N_1646);
xor U2131 (N_2131,N_1361,N_1678);
or U2132 (N_2132,N_1179,N_1870);
or U2133 (N_2133,N_1841,N_1862);
nor U2134 (N_2134,N_1834,N_1877);
nor U2135 (N_2135,N_1843,N_1280);
nor U2136 (N_2136,N_1918,N_1805);
and U2137 (N_2137,N_1854,N_1049);
or U2138 (N_2138,N_1911,N_1923);
or U2139 (N_2139,N_1695,N_1201);
nor U2140 (N_2140,N_1118,N_1145);
xor U2141 (N_2141,N_1080,N_1974);
or U2142 (N_2142,N_1298,N_1734);
nor U2143 (N_2143,N_1955,N_1842);
nand U2144 (N_2144,N_1264,N_1864);
nand U2145 (N_2145,N_1661,N_1288);
and U2146 (N_2146,N_1508,N_1337);
nand U2147 (N_2147,N_1566,N_1585);
nor U2148 (N_2148,N_1222,N_1782);
and U2149 (N_2149,N_1605,N_1476);
nor U2150 (N_2150,N_1691,N_1512);
or U2151 (N_2151,N_1252,N_1146);
or U2152 (N_2152,N_1582,N_1539);
or U2153 (N_2153,N_1262,N_1577);
or U2154 (N_2154,N_1107,N_1939);
xor U2155 (N_2155,N_1354,N_1026);
xor U2156 (N_2156,N_1722,N_1928);
and U2157 (N_2157,N_1617,N_1532);
nor U2158 (N_2158,N_1395,N_1831);
or U2159 (N_2159,N_1074,N_1589);
nor U2160 (N_2160,N_1699,N_1108);
nand U2161 (N_2161,N_1372,N_1667);
or U2162 (N_2162,N_1155,N_1036);
nand U2163 (N_2163,N_1358,N_1503);
or U2164 (N_2164,N_1244,N_1593);
nand U2165 (N_2165,N_1177,N_1794);
and U2166 (N_2166,N_1819,N_1866);
or U2167 (N_2167,N_1952,N_1590);
and U2168 (N_2168,N_1507,N_1293);
nor U2169 (N_2169,N_1478,N_1677);
and U2170 (N_2170,N_1912,N_1065);
nor U2171 (N_2171,N_1980,N_1059);
or U2172 (N_2172,N_1500,N_1635);
or U2173 (N_2173,N_1676,N_1430);
nand U2174 (N_2174,N_1833,N_1360);
nand U2175 (N_2175,N_1013,N_1891);
or U2176 (N_2176,N_1449,N_1787);
xnor U2177 (N_2177,N_1633,N_1575);
xnor U2178 (N_2178,N_1246,N_1793);
or U2179 (N_2179,N_1164,N_1596);
or U2180 (N_2180,N_1627,N_1355);
or U2181 (N_2181,N_1982,N_1487);
nor U2182 (N_2182,N_1998,N_1714);
and U2183 (N_2183,N_1710,N_1312);
xor U2184 (N_2184,N_1111,N_1728);
and U2185 (N_2185,N_1901,N_1409);
and U2186 (N_2186,N_1042,N_1694);
nor U2187 (N_2187,N_1740,N_1239);
nor U2188 (N_2188,N_1171,N_1457);
nand U2189 (N_2189,N_1630,N_1628);
or U2190 (N_2190,N_1030,N_1133);
nor U2191 (N_2191,N_1814,N_1014);
nand U2192 (N_2192,N_1289,N_1654);
and U2193 (N_2193,N_1495,N_1708);
xnor U2194 (N_2194,N_1304,N_1128);
nand U2195 (N_2195,N_1584,N_1019);
and U2196 (N_2196,N_1051,N_1301);
or U2197 (N_2197,N_1975,N_1050);
xnor U2198 (N_2198,N_1170,N_1576);
or U2199 (N_2199,N_1398,N_1504);
nand U2200 (N_2200,N_1324,N_1851);
nand U2201 (N_2201,N_1696,N_1456);
or U2202 (N_2202,N_1669,N_1165);
and U2203 (N_2203,N_1025,N_1417);
nor U2204 (N_2204,N_1443,N_1338);
nor U2205 (N_2205,N_1817,N_1429);
or U2206 (N_2206,N_1341,N_1029);
nand U2207 (N_2207,N_1067,N_1422);
or U2208 (N_2208,N_1547,N_1269);
nand U2209 (N_2209,N_1420,N_1665);
and U2210 (N_2210,N_1733,N_1148);
xnor U2211 (N_2211,N_1749,N_1524);
nand U2212 (N_2212,N_1636,N_1031);
xnor U2213 (N_2213,N_1732,N_1084);
or U2214 (N_2214,N_1045,N_1869);
nor U2215 (N_2215,N_1040,N_1299);
or U2216 (N_2216,N_1725,N_1778);
or U2217 (N_2217,N_1662,N_1154);
nand U2218 (N_2218,N_1857,N_1536);
or U2219 (N_2219,N_1796,N_1625);
or U2220 (N_2220,N_1100,N_1598);
xnor U2221 (N_2221,N_1242,N_1191);
and U2222 (N_2222,N_1052,N_1529);
xor U2223 (N_2223,N_1762,N_1185);
nor U2224 (N_2224,N_1047,N_1707);
or U2225 (N_2225,N_1203,N_1054);
nor U2226 (N_2226,N_1614,N_1463);
and U2227 (N_2227,N_1666,N_1878);
and U2228 (N_2228,N_1688,N_1373);
nand U2229 (N_2229,N_1546,N_1228);
or U2230 (N_2230,N_1462,N_1276);
nor U2231 (N_2231,N_1344,N_1643);
nor U2232 (N_2232,N_1375,N_1718);
nand U2233 (N_2233,N_1989,N_1087);
or U2234 (N_2234,N_1467,N_1122);
nand U2235 (N_2235,N_1292,N_1105);
nand U2236 (N_2236,N_1091,N_1370);
or U2237 (N_2237,N_1189,N_1953);
nor U2238 (N_2238,N_1856,N_1664);
or U2239 (N_2239,N_1580,N_1116);
or U2240 (N_2240,N_1499,N_1571);
or U2241 (N_2241,N_1249,N_1908);
nand U2242 (N_2242,N_1143,N_1531);
xnor U2243 (N_2243,N_1038,N_1438);
nor U2244 (N_2244,N_1406,N_1602);
nand U2245 (N_2245,N_1053,N_1993);
or U2246 (N_2246,N_1915,N_1129);
and U2247 (N_2247,N_1704,N_1035);
nor U2248 (N_2248,N_1682,N_1077);
xnor U2249 (N_2249,N_1188,N_1689);
nor U2250 (N_2250,N_1626,N_1711);
nand U2251 (N_2251,N_1526,N_1460);
nor U2252 (N_2252,N_1224,N_1359);
nor U2253 (N_2253,N_1880,N_1530);
xor U2254 (N_2254,N_1741,N_1932);
nor U2255 (N_2255,N_1624,N_1865);
and U2256 (N_2256,N_1962,N_1379);
nand U2257 (N_2257,N_1303,N_1647);
and U2258 (N_2258,N_1261,N_1541);
xor U2259 (N_2259,N_1340,N_1232);
nand U2260 (N_2260,N_1563,N_1992);
nor U2261 (N_2261,N_1342,N_1957);
nor U2262 (N_2262,N_1540,N_1477);
xnor U2263 (N_2263,N_1798,N_1685);
xnor U2264 (N_2264,N_1437,N_1180);
xnor U2265 (N_2265,N_1972,N_1637);
and U2266 (N_2266,N_1937,N_1979);
or U2267 (N_2267,N_1595,N_1690);
or U2268 (N_2268,N_1588,N_1227);
or U2269 (N_2269,N_1365,N_1768);
nand U2270 (N_2270,N_1138,N_1060);
xnor U2271 (N_2271,N_1480,N_1581);
nand U2272 (N_2272,N_1158,N_1075);
or U2273 (N_2273,N_1335,N_1498);
and U2274 (N_2274,N_1328,N_1182);
or U2275 (N_2275,N_1788,N_1510);
or U2276 (N_2276,N_1209,N_1296);
nor U2277 (N_2277,N_1803,N_1012);
nand U2278 (N_2278,N_1943,N_1199);
nand U2279 (N_2279,N_1959,N_1243);
nor U2280 (N_2280,N_1672,N_1703);
xnor U2281 (N_2281,N_1986,N_1835);
and U2282 (N_2282,N_1184,N_1931);
nand U2283 (N_2283,N_1210,N_1705);
nor U2284 (N_2284,N_1006,N_1300);
or U2285 (N_2285,N_1860,N_1086);
nor U2286 (N_2286,N_1285,N_1076);
or U2287 (N_2287,N_1542,N_1712);
or U2288 (N_2288,N_1969,N_1645);
nor U2289 (N_2289,N_1388,N_1230);
nand U2290 (N_2290,N_1769,N_1846);
xor U2291 (N_2291,N_1996,N_1004);
nor U2292 (N_2292,N_1022,N_1825);
nor U2293 (N_2293,N_1679,N_1558);
nand U2294 (N_2294,N_1927,N_1069);
xnor U2295 (N_2295,N_1149,N_1641);
or U2296 (N_2296,N_1325,N_1058);
and U2297 (N_2297,N_1473,N_1537);
and U2298 (N_2298,N_1823,N_1263);
nor U2299 (N_2299,N_1482,N_1656);
nand U2300 (N_2300,N_1444,N_1294);
xnor U2301 (N_2301,N_1790,N_1632);
xor U2302 (N_2302,N_1991,N_1883);
nor U2303 (N_2303,N_1423,N_1090);
or U2304 (N_2304,N_1267,N_1454);
nand U2305 (N_2305,N_1562,N_1237);
xnor U2306 (N_2306,N_1886,N_1640);
or U2307 (N_2307,N_1828,N_1904);
nor U2308 (N_2308,N_1369,N_1941);
or U2309 (N_2309,N_1384,N_1234);
nor U2310 (N_2310,N_1772,N_1832);
and U2311 (N_2311,N_1015,N_1436);
nand U2312 (N_2312,N_1757,N_1343);
and U2313 (N_2313,N_1615,N_1968);
nand U2314 (N_2314,N_1859,N_1717);
nand U2315 (N_2315,N_1469,N_1751);
nor U2316 (N_2316,N_1046,N_1560);
nand U2317 (N_2317,N_1770,N_1651);
xnor U2318 (N_2318,N_1924,N_1428);
or U2319 (N_2319,N_1917,N_1386);
nand U2320 (N_2320,N_1844,N_1609);
nor U2321 (N_2321,N_1125,N_1988);
or U2322 (N_2322,N_1861,N_1997);
nor U2323 (N_2323,N_1378,N_1779);
nand U2324 (N_2324,N_1553,N_1173);
xor U2325 (N_2325,N_1273,N_1951);
or U2326 (N_2326,N_1238,N_1748);
or U2327 (N_2327,N_1027,N_1502);
nor U2328 (N_2328,N_1657,N_1956);
and U2329 (N_2329,N_1389,N_1362);
xnor U2330 (N_2330,N_1884,N_1401);
nand U2331 (N_2331,N_1063,N_1984);
and U2332 (N_2332,N_1961,N_1876);
and U2333 (N_2333,N_1442,N_1135);
xnor U2334 (N_2334,N_1385,N_1954);
nand U2335 (N_2335,N_1254,N_1600);
nor U2336 (N_2336,N_1958,N_1410);
or U2337 (N_2337,N_1291,N_1692);
nor U2338 (N_2338,N_1336,N_1514);
nor U2339 (N_2339,N_1995,N_1761);
nand U2340 (N_2340,N_1693,N_1320);
nor U2341 (N_2341,N_1622,N_1147);
nor U2342 (N_2342,N_1601,N_1548);
nor U2343 (N_2343,N_1709,N_1942);
nor U2344 (N_2344,N_1414,N_1061);
xnor U2345 (N_2345,N_1352,N_1441);
and U2346 (N_2346,N_1070,N_1157);
nor U2347 (N_2347,N_1785,N_1897);
nand U2348 (N_2348,N_1491,N_1629);
nand U2349 (N_2349,N_1606,N_1127);
or U2350 (N_2350,N_1806,N_1724);
and U2351 (N_2351,N_1871,N_1411);
nor U2352 (N_2352,N_1408,N_1240);
nand U2353 (N_2353,N_1327,N_1745);
and U2354 (N_2354,N_1002,N_1284);
nor U2355 (N_2355,N_1885,N_1440);
nand U2356 (N_2356,N_1217,N_1134);
xnor U2357 (N_2357,N_1879,N_1611);
xor U2358 (N_2358,N_1037,N_1713);
or U2359 (N_2359,N_1505,N_1381);
nand U2360 (N_2360,N_1426,N_1750);
xnor U2361 (N_2361,N_1822,N_1742);
xor U2362 (N_2362,N_1760,N_1490);
nand U2363 (N_2363,N_1028,N_1136);
xor U2364 (N_2364,N_1583,N_1413);
xor U2365 (N_2365,N_1944,N_1660);
xor U2366 (N_2366,N_1702,N_1315);
nand U2367 (N_2367,N_1727,N_1815);
nor U2368 (N_2368,N_1088,N_1936);
and U2369 (N_2369,N_1392,N_1251);
nand U2370 (N_2370,N_1985,N_1383);
xor U2371 (N_2371,N_1175,N_1720);
and U2372 (N_2372,N_1888,N_1445);
nand U2373 (N_2373,N_1150,N_1791);
nand U2374 (N_2374,N_1774,N_1763);
and U2375 (N_2375,N_1812,N_1208);
xor U2376 (N_2376,N_1739,N_1754);
and U2377 (N_2377,N_1631,N_1701);
and U2378 (N_2378,N_1225,N_1781);
nand U2379 (N_2379,N_1648,N_1698);
nor U2380 (N_2380,N_1680,N_1820);
and U2381 (N_2381,N_1516,N_1113);
nand U2382 (N_2382,N_1784,N_1738);
or U2383 (N_2383,N_1187,N_1913);
and U2384 (N_2384,N_1565,N_1845);
nor U2385 (N_2385,N_1567,N_1290);
xor U2386 (N_2386,N_1265,N_1331);
xor U2387 (N_2387,N_1101,N_1579);
and U2388 (N_2388,N_1000,N_1801);
nor U2389 (N_2389,N_1808,N_1545);
nor U2390 (N_2390,N_1056,N_1591);
nand U2391 (N_2391,N_1905,N_1821);
xor U2392 (N_2392,N_1211,N_1481);
and U2393 (N_2393,N_1007,N_1017);
and U2394 (N_2394,N_1468,N_1668);
and U2395 (N_2395,N_1311,N_1241);
nor U2396 (N_2396,N_1160,N_1152);
nand U2397 (N_2397,N_1250,N_1326);
nand U2398 (N_2398,N_1569,N_1322);
and U2399 (N_2399,N_1055,N_1277);
nand U2400 (N_2400,N_1439,N_1448);
nor U2401 (N_2401,N_1169,N_1226);
nand U2402 (N_2402,N_1099,N_1475);
nor U2403 (N_2403,N_1650,N_1391);
nand U2404 (N_2404,N_1119,N_1221);
nor U2405 (N_2405,N_1840,N_1966);
nor U2406 (N_2406,N_1097,N_1623);
and U2407 (N_2407,N_1930,N_1556);
xnor U2408 (N_2408,N_1235,N_1247);
nand U2409 (N_2409,N_1178,N_1559);
nor U2410 (N_2410,N_1093,N_1274);
xor U2411 (N_2411,N_1607,N_1658);
nor U2412 (N_2412,N_1205,N_1453);
or U2413 (N_2413,N_1800,N_1492);
nor U2414 (N_2414,N_1106,N_1963);
nand U2415 (N_2415,N_1371,N_1202);
xor U2416 (N_2416,N_1594,N_1071);
nor U2417 (N_2417,N_1162,N_1543);
nor U2418 (N_2418,N_1260,N_1747);
xor U2419 (N_2419,N_1659,N_1528);
and U2420 (N_2420,N_1653,N_1434);
or U2421 (N_2421,N_1283,N_1403);
or U2422 (N_2422,N_1142,N_1257);
or U2423 (N_2423,N_1586,N_1920);
xor U2424 (N_2424,N_1797,N_1032);
nor U2425 (N_2425,N_1978,N_1655);
and U2426 (N_2426,N_1104,N_1922);
nor U2427 (N_2427,N_1838,N_1396);
nor U2428 (N_2428,N_1767,N_1421);
or U2429 (N_2429,N_1867,N_1350);
nand U2430 (N_2430,N_1461,N_1765);
xnor U2431 (N_2431,N_1783,N_1419);
xnor U2432 (N_2432,N_1771,N_1450);
nand U2433 (N_2433,N_1620,N_1474);
or U2434 (N_2434,N_1066,N_1501);
xor U2435 (N_2435,N_1163,N_1404);
nor U2436 (N_2436,N_1455,N_1826);
xnor U2437 (N_2437,N_1775,N_1082);
nand U2438 (N_2438,N_1307,N_1726);
and U2439 (N_2439,N_1618,N_1484);
xnor U2440 (N_2440,N_1425,N_1220);
and U2441 (N_2441,N_1174,N_1008);
and U2442 (N_2442,N_1302,N_1397);
and U2443 (N_2443,N_1730,N_1736);
nor U2444 (N_2444,N_1935,N_1914);
nand U2445 (N_2445,N_1452,N_1899);
or U2446 (N_2446,N_1687,N_1112);
or U2447 (N_2447,N_1721,N_1756);
and U2448 (N_2448,N_1057,N_1483);
nand U2449 (N_2449,N_1323,N_1126);
nand U2450 (N_2450,N_1094,N_1318);
nand U2451 (N_2451,N_1493,N_1940);
or U2452 (N_2452,N_1807,N_1333);
nand U2453 (N_2453,N_1044,N_1853);
xor U2454 (N_2454,N_1272,N_1470);
and U2455 (N_2455,N_1281,N_1971);
nand U2456 (N_2456,N_1792,N_1946);
nor U2457 (N_2457,N_1719,N_1977);
xnor U2458 (N_2458,N_1723,N_1818);
and U2459 (N_2459,N_1092,N_1003);
nand U2460 (N_2460,N_1776,N_1121);
xor U2461 (N_2461,N_1393,N_1970);
or U2462 (N_2462,N_1759,N_1023);
nor U2463 (N_2463,N_1578,N_1568);
xnor U2464 (N_2464,N_1900,N_1603);
nand U2465 (N_2465,N_1206,N_1903);
nor U2466 (N_2466,N_1681,N_1683);
nor U2467 (N_2467,N_1599,N_1279);
or U2468 (N_2468,N_1592,N_1479);
nand U2469 (N_2469,N_1176,N_1109);
nor U2470 (N_2470,N_1278,N_1433);
nand U2471 (N_2471,N_1639,N_1024);
and U2472 (N_2472,N_1731,N_1416);
or U2473 (N_2473,N_1380,N_1967);
and U2474 (N_2474,N_1376,N_1068);
xnor U2475 (N_2475,N_1287,N_1837);
and U2476 (N_2476,N_1830,N_1613);
and U2477 (N_2477,N_1496,N_1348);
nand U2478 (N_2478,N_1041,N_1960);
and U2479 (N_2479,N_1827,N_1497);
nor U2480 (N_2480,N_1295,N_1909);
or U2481 (N_2481,N_1366,N_1621);
nor U2482 (N_2482,N_1652,N_1349);
and U2483 (N_2483,N_1945,N_1306);
nand U2484 (N_2484,N_1964,N_1663);
or U2485 (N_2485,N_1697,N_1527);
nand U2486 (N_2486,N_1435,N_1557);
xnor U2487 (N_2487,N_1130,N_1824);
or U2488 (N_2488,N_1850,N_1181);
and U2489 (N_2489,N_1890,N_1156);
xor U2490 (N_2490,N_1095,N_1858);
nor U2491 (N_2491,N_1382,N_1872);
and U2492 (N_2492,N_1214,N_1103);
xor U2493 (N_2493,N_1256,N_1096);
nand U2494 (N_2494,N_1649,N_1219);
and U2495 (N_2495,N_1151,N_1168);
nand U2496 (N_2496,N_1330,N_1674);
xor U2497 (N_2497,N_1906,N_1990);
or U2498 (N_2498,N_1018,N_1405);
xnor U2499 (N_2499,N_1889,N_1551);
nor U2500 (N_2500,N_1776,N_1190);
and U2501 (N_2501,N_1700,N_1238);
and U2502 (N_2502,N_1332,N_1357);
xor U2503 (N_2503,N_1909,N_1277);
nor U2504 (N_2504,N_1445,N_1921);
and U2505 (N_2505,N_1327,N_1821);
nand U2506 (N_2506,N_1744,N_1410);
and U2507 (N_2507,N_1181,N_1340);
nand U2508 (N_2508,N_1265,N_1225);
or U2509 (N_2509,N_1548,N_1783);
and U2510 (N_2510,N_1940,N_1570);
and U2511 (N_2511,N_1950,N_1070);
or U2512 (N_2512,N_1403,N_1082);
or U2513 (N_2513,N_1091,N_1675);
nor U2514 (N_2514,N_1999,N_1840);
and U2515 (N_2515,N_1597,N_1112);
nand U2516 (N_2516,N_1420,N_1806);
xor U2517 (N_2517,N_1400,N_1395);
nor U2518 (N_2518,N_1900,N_1741);
and U2519 (N_2519,N_1907,N_1918);
nand U2520 (N_2520,N_1944,N_1977);
or U2521 (N_2521,N_1066,N_1549);
nand U2522 (N_2522,N_1604,N_1092);
or U2523 (N_2523,N_1328,N_1198);
nand U2524 (N_2524,N_1398,N_1468);
and U2525 (N_2525,N_1501,N_1419);
xnor U2526 (N_2526,N_1351,N_1848);
and U2527 (N_2527,N_1143,N_1378);
nor U2528 (N_2528,N_1859,N_1205);
xor U2529 (N_2529,N_1235,N_1974);
and U2530 (N_2530,N_1063,N_1609);
and U2531 (N_2531,N_1304,N_1713);
nor U2532 (N_2532,N_1191,N_1395);
and U2533 (N_2533,N_1019,N_1216);
xnor U2534 (N_2534,N_1418,N_1914);
or U2535 (N_2535,N_1544,N_1550);
xor U2536 (N_2536,N_1262,N_1936);
xor U2537 (N_2537,N_1112,N_1093);
nor U2538 (N_2538,N_1570,N_1442);
and U2539 (N_2539,N_1009,N_1948);
xnor U2540 (N_2540,N_1481,N_1137);
nand U2541 (N_2541,N_1923,N_1082);
xor U2542 (N_2542,N_1101,N_1526);
or U2543 (N_2543,N_1662,N_1760);
and U2544 (N_2544,N_1956,N_1327);
xnor U2545 (N_2545,N_1735,N_1230);
xor U2546 (N_2546,N_1029,N_1274);
nand U2547 (N_2547,N_1804,N_1647);
and U2548 (N_2548,N_1290,N_1703);
nand U2549 (N_2549,N_1216,N_1285);
xor U2550 (N_2550,N_1819,N_1999);
or U2551 (N_2551,N_1151,N_1308);
nand U2552 (N_2552,N_1324,N_1326);
xor U2553 (N_2553,N_1096,N_1473);
nand U2554 (N_2554,N_1119,N_1124);
nor U2555 (N_2555,N_1258,N_1608);
nor U2556 (N_2556,N_1392,N_1471);
xnor U2557 (N_2557,N_1352,N_1550);
nand U2558 (N_2558,N_1413,N_1477);
xor U2559 (N_2559,N_1470,N_1908);
xor U2560 (N_2560,N_1980,N_1141);
or U2561 (N_2561,N_1191,N_1434);
and U2562 (N_2562,N_1852,N_1894);
or U2563 (N_2563,N_1121,N_1945);
or U2564 (N_2564,N_1061,N_1513);
nand U2565 (N_2565,N_1779,N_1047);
and U2566 (N_2566,N_1059,N_1883);
and U2567 (N_2567,N_1434,N_1912);
nor U2568 (N_2568,N_1771,N_1874);
xnor U2569 (N_2569,N_1936,N_1996);
or U2570 (N_2570,N_1627,N_1873);
nor U2571 (N_2571,N_1173,N_1404);
and U2572 (N_2572,N_1677,N_1437);
xor U2573 (N_2573,N_1615,N_1010);
nor U2574 (N_2574,N_1705,N_1328);
nor U2575 (N_2575,N_1858,N_1256);
nor U2576 (N_2576,N_1803,N_1582);
nor U2577 (N_2577,N_1853,N_1028);
nor U2578 (N_2578,N_1246,N_1917);
nand U2579 (N_2579,N_1826,N_1362);
xnor U2580 (N_2580,N_1774,N_1027);
and U2581 (N_2581,N_1597,N_1220);
xnor U2582 (N_2582,N_1370,N_1075);
xnor U2583 (N_2583,N_1799,N_1661);
and U2584 (N_2584,N_1047,N_1339);
nor U2585 (N_2585,N_1544,N_1917);
or U2586 (N_2586,N_1763,N_1748);
nand U2587 (N_2587,N_1496,N_1419);
nor U2588 (N_2588,N_1474,N_1733);
and U2589 (N_2589,N_1484,N_1490);
nand U2590 (N_2590,N_1780,N_1178);
xnor U2591 (N_2591,N_1503,N_1663);
and U2592 (N_2592,N_1263,N_1349);
nor U2593 (N_2593,N_1908,N_1902);
and U2594 (N_2594,N_1785,N_1797);
nor U2595 (N_2595,N_1064,N_1716);
or U2596 (N_2596,N_1352,N_1388);
nor U2597 (N_2597,N_1387,N_1042);
or U2598 (N_2598,N_1566,N_1507);
nor U2599 (N_2599,N_1444,N_1139);
or U2600 (N_2600,N_1273,N_1345);
or U2601 (N_2601,N_1766,N_1592);
nor U2602 (N_2602,N_1547,N_1346);
and U2603 (N_2603,N_1922,N_1224);
xor U2604 (N_2604,N_1092,N_1331);
or U2605 (N_2605,N_1574,N_1338);
and U2606 (N_2606,N_1189,N_1802);
nand U2607 (N_2607,N_1567,N_1011);
or U2608 (N_2608,N_1740,N_1899);
nor U2609 (N_2609,N_1892,N_1782);
or U2610 (N_2610,N_1058,N_1090);
or U2611 (N_2611,N_1483,N_1839);
or U2612 (N_2612,N_1534,N_1614);
nor U2613 (N_2613,N_1095,N_1424);
and U2614 (N_2614,N_1431,N_1057);
xor U2615 (N_2615,N_1058,N_1133);
xor U2616 (N_2616,N_1598,N_1182);
or U2617 (N_2617,N_1742,N_1593);
xor U2618 (N_2618,N_1332,N_1002);
xnor U2619 (N_2619,N_1541,N_1458);
xor U2620 (N_2620,N_1603,N_1990);
nor U2621 (N_2621,N_1886,N_1238);
or U2622 (N_2622,N_1577,N_1042);
and U2623 (N_2623,N_1487,N_1184);
and U2624 (N_2624,N_1381,N_1168);
and U2625 (N_2625,N_1967,N_1025);
xnor U2626 (N_2626,N_1300,N_1583);
or U2627 (N_2627,N_1839,N_1845);
xnor U2628 (N_2628,N_1769,N_1808);
xnor U2629 (N_2629,N_1428,N_1503);
or U2630 (N_2630,N_1429,N_1339);
and U2631 (N_2631,N_1748,N_1798);
and U2632 (N_2632,N_1243,N_1981);
and U2633 (N_2633,N_1372,N_1776);
nor U2634 (N_2634,N_1961,N_1814);
and U2635 (N_2635,N_1621,N_1787);
nor U2636 (N_2636,N_1512,N_1145);
nand U2637 (N_2637,N_1836,N_1579);
xor U2638 (N_2638,N_1840,N_1515);
nor U2639 (N_2639,N_1071,N_1742);
xor U2640 (N_2640,N_1528,N_1679);
or U2641 (N_2641,N_1659,N_1225);
nor U2642 (N_2642,N_1780,N_1636);
nand U2643 (N_2643,N_1971,N_1708);
xor U2644 (N_2644,N_1943,N_1710);
or U2645 (N_2645,N_1059,N_1690);
xor U2646 (N_2646,N_1882,N_1082);
or U2647 (N_2647,N_1640,N_1921);
xnor U2648 (N_2648,N_1927,N_1542);
xnor U2649 (N_2649,N_1699,N_1641);
nand U2650 (N_2650,N_1753,N_1016);
xor U2651 (N_2651,N_1451,N_1180);
nand U2652 (N_2652,N_1810,N_1051);
and U2653 (N_2653,N_1437,N_1986);
or U2654 (N_2654,N_1579,N_1152);
xnor U2655 (N_2655,N_1810,N_1296);
or U2656 (N_2656,N_1703,N_1567);
nor U2657 (N_2657,N_1352,N_1419);
nor U2658 (N_2658,N_1687,N_1991);
nand U2659 (N_2659,N_1154,N_1639);
nand U2660 (N_2660,N_1821,N_1341);
or U2661 (N_2661,N_1572,N_1058);
xnor U2662 (N_2662,N_1134,N_1264);
or U2663 (N_2663,N_1070,N_1307);
xor U2664 (N_2664,N_1896,N_1376);
and U2665 (N_2665,N_1500,N_1106);
xnor U2666 (N_2666,N_1867,N_1320);
or U2667 (N_2667,N_1629,N_1205);
and U2668 (N_2668,N_1038,N_1078);
nand U2669 (N_2669,N_1215,N_1461);
or U2670 (N_2670,N_1147,N_1106);
xor U2671 (N_2671,N_1347,N_1912);
nor U2672 (N_2672,N_1547,N_1978);
nor U2673 (N_2673,N_1210,N_1692);
xnor U2674 (N_2674,N_1746,N_1019);
and U2675 (N_2675,N_1676,N_1150);
or U2676 (N_2676,N_1006,N_1111);
nand U2677 (N_2677,N_1745,N_1591);
xor U2678 (N_2678,N_1012,N_1218);
or U2679 (N_2679,N_1468,N_1646);
or U2680 (N_2680,N_1915,N_1208);
and U2681 (N_2681,N_1998,N_1721);
or U2682 (N_2682,N_1637,N_1315);
and U2683 (N_2683,N_1611,N_1350);
and U2684 (N_2684,N_1321,N_1410);
nor U2685 (N_2685,N_1143,N_1075);
xor U2686 (N_2686,N_1856,N_1540);
nand U2687 (N_2687,N_1258,N_1406);
nand U2688 (N_2688,N_1337,N_1568);
or U2689 (N_2689,N_1876,N_1516);
nor U2690 (N_2690,N_1410,N_1275);
nor U2691 (N_2691,N_1415,N_1392);
and U2692 (N_2692,N_1876,N_1317);
nand U2693 (N_2693,N_1745,N_1723);
and U2694 (N_2694,N_1902,N_1050);
nand U2695 (N_2695,N_1402,N_1851);
or U2696 (N_2696,N_1232,N_1590);
nor U2697 (N_2697,N_1783,N_1345);
nor U2698 (N_2698,N_1514,N_1707);
xor U2699 (N_2699,N_1859,N_1143);
or U2700 (N_2700,N_1680,N_1924);
and U2701 (N_2701,N_1310,N_1186);
nand U2702 (N_2702,N_1202,N_1133);
or U2703 (N_2703,N_1093,N_1252);
or U2704 (N_2704,N_1509,N_1953);
nand U2705 (N_2705,N_1442,N_1835);
and U2706 (N_2706,N_1524,N_1876);
and U2707 (N_2707,N_1599,N_1720);
or U2708 (N_2708,N_1302,N_1414);
nor U2709 (N_2709,N_1745,N_1702);
nor U2710 (N_2710,N_1776,N_1601);
or U2711 (N_2711,N_1288,N_1015);
nor U2712 (N_2712,N_1757,N_1860);
xor U2713 (N_2713,N_1632,N_1654);
nand U2714 (N_2714,N_1885,N_1614);
nor U2715 (N_2715,N_1729,N_1322);
nor U2716 (N_2716,N_1071,N_1830);
xnor U2717 (N_2717,N_1108,N_1348);
nand U2718 (N_2718,N_1548,N_1985);
and U2719 (N_2719,N_1275,N_1916);
xor U2720 (N_2720,N_1711,N_1946);
or U2721 (N_2721,N_1854,N_1152);
xor U2722 (N_2722,N_1388,N_1385);
and U2723 (N_2723,N_1698,N_1338);
or U2724 (N_2724,N_1743,N_1933);
nor U2725 (N_2725,N_1226,N_1715);
and U2726 (N_2726,N_1606,N_1731);
nand U2727 (N_2727,N_1158,N_1220);
or U2728 (N_2728,N_1906,N_1760);
xnor U2729 (N_2729,N_1847,N_1155);
nor U2730 (N_2730,N_1199,N_1236);
nand U2731 (N_2731,N_1060,N_1292);
nand U2732 (N_2732,N_1129,N_1160);
and U2733 (N_2733,N_1504,N_1188);
or U2734 (N_2734,N_1200,N_1354);
and U2735 (N_2735,N_1513,N_1292);
nand U2736 (N_2736,N_1954,N_1060);
xnor U2737 (N_2737,N_1915,N_1259);
nand U2738 (N_2738,N_1429,N_1112);
nor U2739 (N_2739,N_1092,N_1658);
nor U2740 (N_2740,N_1095,N_1661);
and U2741 (N_2741,N_1879,N_1708);
xor U2742 (N_2742,N_1407,N_1374);
nand U2743 (N_2743,N_1083,N_1806);
nand U2744 (N_2744,N_1912,N_1156);
nor U2745 (N_2745,N_1964,N_1496);
or U2746 (N_2746,N_1494,N_1008);
nand U2747 (N_2747,N_1361,N_1901);
or U2748 (N_2748,N_1765,N_1016);
and U2749 (N_2749,N_1541,N_1155);
nand U2750 (N_2750,N_1184,N_1295);
xnor U2751 (N_2751,N_1587,N_1741);
or U2752 (N_2752,N_1404,N_1211);
nor U2753 (N_2753,N_1334,N_1541);
and U2754 (N_2754,N_1052,N_1041);
nand U2755 (N_2755,N_1917,N_1280);
nor U2756 (N_2756,N_1345,N_1449);
nor U2757 (N_2757,N_1975,N_1137);
nor U2758 (N_2758,N_1629,N_1428);
xnor U2759 (N_2759,N_1520,N_1135);
and U2760 (N_2760,N_1861,N_1314);
and U2761 (N_2761,N_1344,N_1700);
nor U2762 (N_2762,N_1935,N_1445);
nand U2763 (N_2763,N_1044,N_1402);
nor U2764 (N_2764,N_1419,N_1172);
and U2765 (N_2765,N_1636,N_1849);
or U2766 (N_2766,N_1783,N_1685);
nor U2767 (N_2767,N_1145,N_1811);
xor U2768 (N_2768,N_1848,N_1521);
xor U2769 (N_2769,N_1162,N_1335);
xor U2770 (N_2770,N_1049,N_1613);
nor U2771 (N_2771,N_1630,N_1016);
or U2772 (N_2772,N_1098,N_1485);
and U2773 (N_2773,N_1210,N_1552);
and U2774 (N_2774,N_1574,N_1295);
nor U2775 (N_2775,N_1981,N_1548);
and U2776 (N_2776,N_1214,N_1863);
nand U2777 (N_2777,N_1348,N_1249);
xor U2778 (N_2778,N_1658,N_1148);
or U2779 (N_2779,N_1880,N_1623);
or U2780 (N_2780,N_1704,N_1349);
or U2781 (N_2781,N_1875,N_1587);
or U2782 (N_2782,N_1355,N_1204);
or U2783 (N_2783,N_1404,N_1950);
or U2784 (N_2784,N_1095,N_1954);
xnor U2785 (N_2785,N_1545,N_1670);
and U2786 (N_2786,N_1132,N_1803);
xnor U2787 (N_2787,N_1678,N_1255);
nor U2788 (N_2788,N_1788,N_1246);
xor U2789 (N_2789,N_1392,N_1555);
nor U2790 (N_2790,N_1435,N_1750);
nand U2791 (N_2791,N_1212,N_1328);
and U2792 (N_2792,N_1324,N_1537);
and U2793 (N_2793,N_1137,N_1040);
xnor U2794 (N_2794,N_1992,N_1539);
xnor U2795 (N_2795,N_1035,N_1386);
xor U2796 (N_2796,N_1037,N_1220);
xor U2797 (N_2797,N_1551,N_1425);
nor U2798 (N_2798,N_1464,N_1030);
nand U2799 (N_2799,N_1777,N_1915);
xnor U2800 (N_2800,N_1295,N_1903);
and U2801 (N_2801,N_1640,N_1750);
nor U2802 (N_2802,N_1971,N_1122);
and U2803 (N_2803,N_1435,N_1776);
or U2804 (N_2804,N_1710,N_1054);
nor U2805 (N_2805,N_1589,N_1611);
or U2806 (N_2806,N_1859,N_1824);
or U2807 (N_2807,N_1514,N_1520);
nand U2808 (N_2808,N_1698,N_1393);
nand U2809 (N_2809,N_1830,N_1801);
xor U2810 (N_2810,N_1153,N_1584);
or U2811 (N_2811,N_1423,N_1973);
nor U2812 (N_2812,N_1077,N_1613);
nor U2813 (N_2813,N_1066,N_1261);
or U2814 (N_2814,N_1823,N_1371);
and U2815 (N_2815,N_1153,N_1270);
xor U2816 (N_2816,N_1202,N_1777);
xor U2817 (N_2817,N_1318,N_1177);
nor U2818 (N_2818,N_1365,N_1104);
and U2819 (N_2819,N_1323,N_1723);
nand U2820 (N_2820,N_1623,N_1384);
nor U2821 (N_2821,N_1745,N_1262);
xor U2822 (N_2822,N_1850,N_1264);
xnor U2823 (N_2823,N_1468,N_1479);
or U2824 (N_2824,N_1671,N_1038);
nand U2825 (N_2825,N_1159,N_1992);
or U2826 (N_2826,N_1493,N_1983);
nor U2827 (N_2827,N_1127,N_1477);
and U2828 (N_2828,N_1108,N_1969);
or U2829 (N_2829,N_1256,N_1324);
nand U2830 (N_2830,N_1495,N_1634);
or U2831 (N_2831,N_1379,N_1790);
nand U2832 (N_2832,N_1394,N_1942);
and U2833 (N_2833,N_1984,N_1769);
and U2834 (N_2834,N_1590,N_1919);
nand U2835 (N_2835,N_1442,N_1201);
and U2836 (N_2836,N_1086,N_1613);
nor U2837 (N_2837,N_1184,N_1728);
nand U2838 (N_2838,N_1195,N_1658);
xor U2839 (N_2839,N_1228,N_1995);
xor U2840 (N_2840,N_1590,N_1392);
xnor U2841 (N_2841,N_1513,N_1831);
nor U2842 (N_2842,N_1320,N_1146);
or U2843 (N_2843,N_1012,N_1672);
and U2844 (N_2844,N_1210,N_1880);
xor U2845 (N_2845,N_1851,N_1869);
and U2846 (N_2846,N_1686,N_1309);
nor U2847 (N_2847,N_1979,N_1075);
nor U2848 (N_2848,N_1116,N_1863);
nand U2849 (N_2849,N_1589,N_1499);
nor U2850 (N_2850,N_1446,N_1263);
or U2851 (N_2851,N_1618,N_1250);
xnor U2852 (N_2852,N_1300,N_1147);
xor U2853 (N_2853,N_1174,N_1445);
nand U2854 (N_2854,N_1139,N_1304);
nand U2855 (N_2855,N_1922,N_1400);
nor U2856 (N_2856,N_1175,N_1502);
xnor U2857 (N_2857,N_1107,N_1275);
or U2858 (N_2858,N_1558,N_1426);
xnor U2859 (N_2859,N_1626,N_1545);
or U2860 (N_2860,N_1081,N_1023);
and U2861 (N_2861,N_1347,N_1818);
xnor U2862 (N_2862,N_1366,N_1719);
and U2863 (N_2863,N_1687,N_1423);
nand U2864 (N_2864,N_1152,N_1932);
xor U2865 (N_2865,N_1435,N_1971);
nor U2866 (N_2866,N_1391,N_1856);
xnor U2867 (N_2867,N_1289,N_1968);
and U2868 (N_2868,N_1845,N_1636);
xnor U2869 (N_2869,N_1678,N_1943);
and U2870 (N_2870,N_1489,N_1890);
and U2871 (N_2871,N_1559,N_1791);
xor U2872 (N_2872,N_1811,N_1675);
and U2873 (N_2873,N_1614,N_1298);
nand U2874 (N_2874,N_1865,N_1279);
xnor U2875 (N_2875,N_1709,N_1278);
and U2876 (N_2876,N_1941,N_1613);
nand U2877 (N_2877,N_1276,N_1354);
nand U2878 (N_2878,N_1126,N_1411);
xnor U2879 (N_2879,N_1706,N_1708);
nand U2880 (N_2880,N_1445,N_1169);
xor U2881 (N_2881,N_1127,N_1888);
or U2882 (N_2882,N_1041,N_1807);
nor U2883 (N_2883,N_1664,N_1386);
xor U2884 (N_2884,N_1251,N_1203);
nand U2885 (N_2885,N_1876,N_1515);
and U2886 (N_2886,N_1413,N_1941);
xnor U2887 (N_2887,N_1673,N_1169);
nand U2888 (N_2888,N_1534,N_1447);
nor U2889 (N_2889,N_1150,N_1215);
or U2890 (N_2890,N_1679,N_1381);
nor U2891 (N_2891,N_1675,N_1666);
and U2892 (N_2892,N_1314,N_1119);
and U2893 (N_2893,N_1840,N_1157);
or U2894 (N_2894,N_1326,N_1287);
and U2895 (N_2895,N_1180,N_1736);
nor U2896 (N_2896,N_1603,N_1425);
or U2897 (N_2897,N_1746,N_1979);
and U2898 (N_2898,N_1521,N_1089);
nand U2899 (N_2899,N_1797,N_1230);
or U2900 (N_2900,N_1250,N_1694);
or U2901 (N_2901,N_1567,N_1280);
xnor U2902 (N_2902,N_1690,N_1079);
or U2903 (N_2903,N_1185,N_1075);
and U2904 (N_2904,N_1315,N_1511);
or U2905 (N_2905,N_1327,N_1573);
nand U2906 (N_2906,N_1022,N_1904);
or U2907 (N_2907,N_1825,N_1380);
xnor U2908 (N_2908,N_1287,N_1937);
and U2909 (N_2909,N_1428,N_1339);
or U2910 (N_2910,N_1656,N_1818);
nand U2911 (N_2911,N_1135,N_1942);
or U2912 (N_2912,N_1905,N_1563);
nor U2913 (N_2913,N_1246,N_1572);
nand U2914 (N_2914,N_1874,N_1521);
or U2915 (N_2915,N_1967,N_1957);
nand U2916 (N_2916,N_1813,N_1433);
nand U2917 (N_2917,N_1704,N_1046);
or U2918 (N_2918,N_1314,N_1964);
nand U2919 (N_2919,N_1657,N_1350);
xnor U2920 (N_2920,N_1336,N_1897);
nand U2921 (N_2921,N_1047,N_1130);
xnor U2922 (N_2922,N_1719,N_1437);
nand U2923 (N_2923,N_1318,N_1341);
nand U2924 (N_2924,N_1068,N_1087);
nor U2925 (N_2925,N_1466,N_1319);
nand U2926 (N_2926,N_1024,N_1121);
nor U2927 (N_2927,N_1511,N_1189);
or U2928 (N_2928,N_1257,N_1060);
nand U2929 (N_2929,N_1315,N_1888);
nor U2930 (N_2930,N_1567,N_1978);
nor U2931 (N_2931,N_1089,N_1565);
nand U2932 (N_2932,N_1234,N_1231);
and U2933 (N_2933,N_1339,N_1686);
xor U2934 (N_2934,N_1619,N_1713);
and U2935 (N_2935,N_1757,N_1418);
xnor U2936 (N_2936,N_1078,N_1224);
nand U2937 (N_2937,N_1078,N_1655);
and U2938 (N_2938,N_1008,N_1630);
and U2939 (N_2939,N_1570,N_1927);
xor U2940 (N_2940,N_1769,N_1258);
and U2941 (N_2941,N_1100,N_1807);
and U2942 (N_2942,N_1630,N_1007);
xnor U2943 (N_2943,N_1830,N_1945);
or U2944 (N_2944,N_1813,N_1181);
xnor U2945 (N_2945,N_1304,N_1726);
nor U2946 (N_2946,N_1873,N_1951);
nand U2947 (N_2947,N_1051,N_1873);
and U2948 (N_2948,N_1448,N_1284);
nand U2949 (N_2949,N_1703,N_1619);
nor U2950 (N_2950,N_1965,N_1654);
nand U2951 (N_2951,N_1251,N_1903);
nand U2952 (N_2952,N_1469,N_1483);
and U2953 (N_2953,N_1682,N_1700);
or U2954 (N_2954,N_1674,N_1746);
and U2955 (N_2955,N_1594,N_1807);
and U2956 (N_2956,N_1956,N_1859);
and U2957 (N_2957,N_1954,N_1106);
or U2958 (N_2958,N_1747,N_1700);
and U2959 (N_2959,N_1848,N_1654);
nor U2960 (N_2960,N_1297,N_1574);
nand U2961 (N_2961,N_1259,N_1572);
nand U2962 (N_2962,N_1121,N_1523);
xnor U2963 (N_2963,N_1270,N_1380);
or U2964 (N_2964,N_1944,N_1770);
and U2965 (N_2965,N_1352,N_1919);
or U2966 (N_2966,N_1494,N_1382);
xnor U2967 (N_2967,N_1238,N_1807);
or U2968 (N_2968,N_1420,N_1637);
nor U2969 (N_2969,N_1524,N_1841);
nand U2970 (N_2970,N_1053,N_1339);
nand U2971 (N_2971,N_1010,N_1749);
xor U2972 (N_2972,N_1950,N_1608);
or U2973 (N_2973,N_1867,N_1373);
xor U2974 (N_2974,N_1577,N_1229);
nand U2975 (N_2975,N_1865,N_1718);
and U2976 (N_2976,N_1667,N_1828);
nor U2977 (N_2977,N_1438,N_1436);
nor U2978 (N_2978,N_1858,N_1876);
xor U2979 (N_2979,N_1583,N_1262);
nand U2980 (N_2980,N_1049,N_1257);
nor U2981 (N_2981,N_1127,N_1883);
or U2982 (N_2982,N_1427,N_1216);
xnor U2983 (N_2983,N_1266,N_1121);
nand U2984 (N_2984,N_1071,N_1843);
nand U2985 (N_2985,N_1890,N_1137);
and U2986 (N_2986,N_1676,N_1594);
nand U2987 (N_2987,N_1740,N_1770);
xor U2988 (N_2988,N_1689,N_1088);
nor U2989 (N_2989,N_1207,N_1070);
nor U2990 (N_2990,N_1807,N_1401);
or U2991 (N_2991,N_1071,N_1520);
nor U2992 (N_2992,N_1362,N_1317);
nand U2993 (N_2993,N_1225,N_1336);
xnor U2994 (N_2994,N_1469,N_1569);
xnor U2995 (N_2995,N_1233,N_1827);
or U2996 (N_2996,N_1227,N_1796);
or U2997 (N_2997,N_1077,N_1981);
or U2998 (N_2998,N_1294,N_1334);
and U2999 (N_2999,N_1468,N_1786);
or U3000 (N_3000,N_2079,N_2455);
nand U3001 (N_3001,N_2735,N_2649);
nand U3002 (N_3002,N_2543,N_2774);
xnor U3003 (N_3003,N_2744,N_2768);
nor U3004 (N_3004,N_2662,N_2444);
or U3005 (N_3005,N_2131,N_2199);
and U3006 (N_3006,N_2177,N_2992);
nand U3007 (N_3007,N_2099,N_2695);
and U3008 (N_3008,N_2874,N_2640);
nand U3009 (N_3009,N_2164,N_2779);
xnor U3010 (N_3010,N_2610,N_2959);
and U3011 (N_3011,N_2669,N_2214);
nand U3012 (N_3012,N_2514,N_2036);
nand U3013 (N_3013,N_2712,N_2435);
or U3014 (N_3014,N_2719,N_2069);
nand U3015 (N_3015,N_2900,N_2832);
or U3016 (N_3016,N_2644,N_2458);
xor U3017 (N_3017,N_2805,N_2667);
nor U3018 (N_3018,N_2839,N_2833);
nor U3019 (N_3019,N_2933,N_2072);
nor U3020 (N_3020,N_2464,N_2869);
nor U3021 (N_3021,N_2271,N_2870);
or U3022 (N_3022,N_2357,N_2246);
nor U3023 (N_3023,N_2120,N_2741);
nor U3024 (N_3024,N_2310,N_2687);
or U3025 (N_3025,N_2705,N_2141);
and U3026 (N_3026,N_2736,N_2003);
and U3027 (N_3027,N_2658,N_2809);
or U3028 (N_3028,N_2866,N_2278);
or U3029 (N_3029,N_2180,N_2293);
and U3030 (N_3030,N_2476,N_2620);
or U3031 (N_3031,N_2556,N_2063);
or U3032 (N_3032,N_2415,N_2044);
nor U3033 (N_3033,N_2088,N_2244);
or U3034 (N_3034,N_2264,N_2351);
xnor U3035 (N_3035,N_2837,N_2742);
or U3036 (N_3036,N_2269,N_2300);
nand U3037 (N_3037,N_2161,N_2289);
or U3038 (N_3038,N_2489,N_2134);
nand U3039 (N_3039,N_2263,N_2892);
or U3040 (N_3040,N_2818,N_2864);
xnor U3041 (N_3041,N_2188,N_2802);
nand U3042 (N_3042,N_2976,N_2600);
xor U3043 (N_3043,N_2137,N_2077);
and U3044 (N_3044,N_2296,N_2970);
nand U3045 (N_3045,N_2674,N_2206);
nand U3046 (N_3046,N_2852,N_2017);
nand U3047 (N_3047,N_2442,N_2248);
xnor U3048 (N_3048,N_2362,N_2910);
or U3049 (N_3049,N_2738,N_2021);
and U3050 (N_3050,N_2974,N_2569);
nor U3051 (N_3051,N_2957,N_2292);
or U3052 (N_3052,N_2367,N_2086);
or U3053 (N_3053,N_2273,N_2630);
nor U3054 (N_3054,N_2418,N_2405);
xor U3055 (N_3055,N_2345,N_2189);
xor U3056 (N_3056,N_2265,N_2672);
nand U3057 (N_3057,N_2865,N_2225);
xor U3058 (N_3058,N_2522,N_2568);
or U3059 (N_3059,N_2924,N_2819);
nand U3060 (N_3060,N_2806,N_2731);
and U3061 (N_3061,N_2893,N_2043);
and U3062 (N_3062,N_2814,N_2033);
and U3063 (N_3063,N_2082,N_2022);
nor U3064 (N_3064,N_2335,N_2563);
nor U3065 (N_3065,N_2666,N_2315);
and U3066 (N_3066,N_2626,N_2845);
xnor U3067 (N_3067,N_2966,N_2130);
nor U3068 (N_3068,N_2450,N_2208);
nand U3069 (N_3069,N_2571,N_2723);
or U3070 (N_3070,N_2734,N_2322);
nand U3071 (N_3071,N_2955,N_2162);
nand U3072 (N_3072,N_2570,N_2813);
or U3073 (N_3073,N_2872,N_2118);
or U3074 (N_3074,N_2449,N_2122);
nand U3075 (N_3075,N_2715,N_2011);
nand U3076 (N_3076,N_2673,N_2235);
or U3077 (N_3077,N_2283,N_2634);
and U3078 (N_3078,N_2958,N_2877);
or U3079 (N_3079,N_2429,N_2690);
xnor U3080 (N_3080,N_2201,N_2601);
nand U3081 (N_3081,N_2093,N_2237);
and U3082 (N_3082,N_2477,N_2932);
nor U3083 (N_3083,N_2124,N_2778);
or U3084 (N_3084,N_2875,N_2725);
xor U3085 (N_3085,N_2332,N_2797);
nand U3086 (N_3086,N_2226,N_2227);
nand U3087 (N_3087,N_2890,N_2680);
nor U3088 (N_3088,N_2420,N_2045);
and U3089 (N_3089,N_2516,N_2711);
nand U3090 (N_3090,N_2037,N_2821);
nor U3091 (N_3091,N_2119,N_2920);
nand U3092 (N_3092,N_2395,N_2615);
or U3093 (N_3093,N_2193,N_2421);
nor U3094 (N_3094,N_2625,N_2907);
and U3095 (N_3095,N_2732,N_2996);
or U3096 (N_3096,N_2758,N_2721);
xor U3097 (N_3097,N_2396,N_2105);
and U3098 (N_3098,N_2685,N_2575);
nand U3099 (N_3099,N_2102,N_2187);
nand U3100 (N_3100,N_2001,N_2139);
xor U3101 (N_3101,N_2585,N_2050);
or U3102 (N_3102,N_2384,N_2720);
xor U3103 (N_3103,N_2297,N_2236);
and U3104 (N_3104,N_2880,N_2794);
xnor U3105 (N_3105,N_2340,N_2174);
or U3106 (N_3106,N_2851,N_2535);
nand U3107 (N_3107,N_2902,N_2453);
xor U3108 (N_3108,N_2937,N_2987);
or U3109 (N_3109,N_2229,N_2196);
nor U3110 (N_3110,N_2915,N_2785);
nor U3111 (N_3111,N_2066,N_2787);
nor U3112 (N_3112,N_2084,N_2372);
xnor U3113 (N_3113,N_2126,N_2588);
or U3114 (N_3114,N_2936,N_2288);
and U3115 (N_3115,N_2995,N_2727);
and U3116 (N_3116,N_2682,N_2906);
or U3117 (N_3117,N_2903,N_2982);
and U3118 (N_3118,N_2109,N_2655);
nor U3119 (N_3119,N_2166,N_2980);
nor U3120 (N_3120,N_2761,N_2108);
xnor U3121 (N_3121,N_2143,N_2954);
or U3122 (N_3122,N_2185,N_2191);
nor U3123 (N_3123,N_2307,N_2078);
nor U3124 (N_3124,N_2049,N_2159);
or U3125 (N_3125,N_2317,N_2309);
and U3126 (N_3126,N_2026,N_2485);
nand U3127 (N_3127,N_2468,N_2402);
nor U3128 (N_3128,N_2800,N_2660);
nor U3129 (N_3129,N_2276,N_2960);
nand U3130 (N_3130,N_2346,N_2117);
nor U3131 (N_3131,N_2073,N_2323);
nor U3132 (N_3132,N_2553,N_2925);
and U3133 (N_3133,N_2128,N_2927);
nand U3134 (N_3134,N_2934,N_2632);
xnor U3135 (N_3135,N_2614,N_2047);
or U3136 (N_3136,N_2243,N_2039);
nand U3137 (N_3137,N_2827,N_2422);
nand U3138 (N_3138,N_2978,N_2055);
or U3139 (N_3139,N_2268,N_2176);
nand U3140 (N_3140,N_2152,N_2546);
xnor U3141 (N_3141,N_2849,N_2540);
nand U3142 (N_3142,N_2173,N_2587);
and U3143 (N_3143,N_2737,N_2425);
and U3144 (N_3144,N_2847,N_2138);
xor U3145 (N_3145,N_2772,N_2071);
or U3146 (N_3146,N_2492,N_2863);
and U3147 (N_3147,N_2270,N_2356);
nand U3148 (N_3148,N_2834,N_2261);
nor U3149 (N_3149,N_2990,N_2596);
xor U3150 (N_3150,N_2984,N_2245);
xnor U3151 (N_3151,N_2502,N_2562);
nor U3152 (N_3152,N_2368,N_2469);
nand U3153 (N_3153,N_2290,N_2080);
nand U3154 (N_3154,N_2500,N_2360);
nor U3155 (N_3155,N_2838,N_2359);
nand U3156 (N_3156,N_2439,N_2697);
or U3157 (N_3157,N_2217,N_2803);
or U3158 (N_3158,N_2733,N_2700);
and U3159 (N_3159,N_2950,N_2272);
xor U3160 (N_3160,N_2320,N_2378);
or U3161 (N_3161,N_2791,N_2266);
nor U3162 (N_3162,N_2058,N_2560);
nor U3163 (N_3163,N_2341,N_2145);
xnor U3164 (N_3164,N_2365,N_2651);
or U3165 (N_3165,N_2090,N_2081);
and U3166 (N_3166,N_2817,N_2679);
or U3167 (N_3167,N_2179,N_2052);
and U3168 (N_3168,N_2490,N_2886);
nor U3169 (N_3169,N_2799,N_2221);
xor U3170 (N_3170,N_2324,N_2197);
and U3171 (N_3171,N_2146,N_2523);
xor U3172 (N_3172,N_2617,N_2621);
and U3173 (N_3173,N_2355,N_2548);
nand U3174 (N_3174,N_2115,N_2487);
and U3175 (N_3175,N_2509,N_2153);
xor U3176 (N_3176,N_2371,N_2859);
and U3177 (N_3177,N_2537,N_2336);
nor U3178 (N_3178,N_2748,N_2815);
nand U3179 (N_3179,N_2769,N_2504);
nor U3180 (N_3180,N_2417,N_2867);
nor U3181 (N_3181,N_2607,N_2408);
and U3182 (N_3182,N_2498,N_2089);
xnor U3183 (N_3183,N_2035,N_2505);
xnor U3184 (N_3184,N_2897,N_2076);
nand U3185 (N_3185,N_2445,N_2949);
nor U3186 (N_3186,N_2671,N_2220);
or U3187 (N_3187,N_2965,N_2401);
nor U3188 (N_3188,N_2777,N_2521);
nor U3189 (N_3189,N_2593,N_2083);
nand U3190 (N_3190,N_2653,N_2232);
xnor U3191 (N_3191,N_2148,N_2528);
nor U3192 (N_3192,N_2413,N_2136);
nand U3193 (N_3193,N_2380,N_2993);
and U3194 (N_3194,N_2430,N_2370);
nand U3195 (N_3195,N_2631,N_2150);
xor U3196 (N_3196,N_2692,N_2098);
or U3197 (N_3197,N_2070,N_2746);
and U3198 (N_3198,N_2530,N_2762);
nor U3199 (N_3199,N_2773,N_2002);
and U3200 (N_3200,N_2251,N_2767);
nand U3201 (N_3201,N_2896,N_2539);
nand U3202 (N_3202,N_2414,N_2030);
nand U3203 (N_3203,N_2018,N_2943);
nor U3204 (N_3204,N_2260,N_2501);
nor U3205 (N_3205,N_2064,N_2280);
xnor U3206 (N_3206,N_2824,N_2754);
nand U3207 (N_3207,N_2178,N_2633);
xnor U3208 (N_3208,N_2602,N_2301);
nand U3209 (N_3209,N_2740,N_2096);
nor U3210 (N_3210,N_2274,N_2545);
and U3211 (N_3211,N_2254,N_2598);
nor U3212 (N_3212,N_2807,N_2713);
or U3213 (N_3213,N_2855,N_2888);
nand U3214 (N_3214,N_2029,N_2125);
nand U3215 (N_3215,N_2067,N_2279);
nor U3216 (N_3216,N_2574,N_2042);
nor U3217 (N_3217,N_2525,N_2060);
or U3218 (N_3218,N_2912,N_2929);
nor U3219 (N_3219,N_2836,N_2510);
nor U3220 (N_3220,N_2032,N_2316);
nand U3221 (N_3221,N_2419,N_2603);
and U3222 (N_3222,N_2314,N_2739);
xnor U3223 (N_3223,N_2350,N_2358);
and U3224 (N_3224,N_2004,N_2503);
nor U3225 (N_3225,N_2506,N_2580);
and U3226 (N_3226,N_2432,N_2515);
and U3227 (N_3227,N_2224,N_2526);
xor U3228 (N_3228,N_2823,N_2804);
or U3229 (N_3229,N_2258,N_2928);
nor U3230 (N_3230,N_2592,N_2776);
xnor U3231 (N_3231,N_2696,N_2133);
or U3232 (N_3232,N_2945,N_2282);
nand U3233 (N_3233,N_2559,N_2461);
xnor U3234 (N_3234,N_2648,N_2218);
or U3235 (N_3235,N_2973,N_2961);
or U3236 (N_3236,N_2686,N_2544);
and U3237 (N_3237,N_2423,N_2828);
and U3238 (N_3238,N_2765,N_2230);
nand U3239 (N_3239,N_2325,N_2895);
nor U3240 (N_3240,N_2142,N_2750);
and U3241 (N_3241,N_2684,N_2262);
xor U3242 (N_3242,N_2062,N_2578);
xor U3243 (N_3243,N_2930,N_2239);
xor U3244 (N_3244,N_2749,N_2013);
nor U3245 (N_3245,N_2678,N_2056);
nand U3246 (N_3246,N_2205,N_2411);
nand U3247 (N_3247,N_2222,N_2657);
and U3248 (N_3248,N_2914,N_2840);
and U3249 (N_3249,N_2154,N_2998);
xnor U3250 (N_3250,N_2312,N_2329);
and U3251 (N_3251,N_2557,N_2707);
nor U3252 (N_3252,N_2726,N_2348);
xnor U3253 (N_3253,N_2894,N_2202);
or U3254 (N_3254,N_2114,N_2475);
and U3255 (N_3255,N_2665,N_2710);
and U3256 (N_3256,N_2443,N_2829);
or U3257 (N_3257,N_2028,N_2170);
or U3258 (N_3258,N_2428,N_2618);
and U3259 (N_3259,N_2688,N_2977);
or U3260 (N_3260,N_2844,N_2377);
nand U3261 (N_3261,N_2353,N_2110);
nand U3262 (N_3262,N_2092,N_2755);
or U3263 (N_3263,N_2223,N_2853);
and U3264 (N_3264,N_2645,N_2167);
or U3265 (N_3265,N_2406,N_2403);
and U3266 (N_3266,N_2520,N_2994);
nand U3267 (N_3267,N_2303,N_2190);
or U3268 (N_3268,N_2459,N_2386);
or U3269 (N_3269,N_2616,N_2472);
and U3270 (N_3270,N_2165,N_2216);
and U3271 (N_3271,N_2000,N_2228);
or U3272 (N_3272,N_2871,N_2519);
and U3273 (N_3273,N_2005,N_2656);
or U3274 (N_3274,N_2463,N_2363);
or U3275 (N_3275,N_2612,N_2287);
nor U3276 (N_3276,N_2771,N_2786);
and U3277 (N_3277,N_2479,N_2156);
and U3278 (N_3278,N_2701,N_2605);
and U3279 (N_3279,N_2862,N_2623);
xnor U3280 (N_3280,N_2583,N_2532);
nand U3281 (N_3281,N_2184,N_2100);
nand U3282 (N_3282,N_2462,N_2249);
xor U3283 (N_3283,N_2981,N_2327);
nand U3284 (N_3284,N_2780,N_2252);
xor U3285 (N_3285,N_2843,N_2926);
and U3286 (N_3286,N_2466,N_2410);
or U3287 (N_3287,N_2881,N_2820);
nand U3288 (N_3288,N_2121,N_2913);
or U3289 (N_3289,N_2714,N_2399);
xnor U3290 (N_3290,N_2347,N_2048);
xnor U3291 (N_3291,N_2650,N_2275);
nor U3292 (N_3292,N_2016,N_2751);
and U3293 (N_3293,N_2057,N_2259);
nor U3294 (N_3294,N_2584,N_2473);
xnor U3295 (N_3295,N_2899,N_2878);
or U3296 (N_3296,N_2416,N_2564);
or U3297 (N_3297,N_2438,N_2361);
or U3298 (N_3298,N_2447,N_2012);
or U3299 (N_3299,N_2319,N_2116);
xnor U3300 (N_3300,N_2664,N_2364);
nand U3301 (N_3301,N_2683,N_2511);
nand U3302 (N_3302,N_2135,N_2209);
and U3303 (N_3303,N_2085,N_2675);
or U3304 (N_3304,N_2397,N_2549);
or U3305 (N_3305,N_2808,N_2195);
and U3306 (N_3306,N_2536,N_2385);
nand U3307 (N_3307,N_2795,N_2497);
nand U3308 (N_3308,N_2677,N_2181);
nor U3309 (N_3309,N_2285,N_2997);
xor U3310 (N_3310,N_2242,N_2728);
nor U3311 (N_3311,N_2972,N_2281);
and U3312 (N_3312,N_2835,N_2919);
or U3313 (N_3313,N_2952,N_2962);
or U3314 (N_3314,N_2956,N_2611);
nand U3315 (N_3315,N_2305,N_2983);
nand U3316 (N_3316,N_2433,N_2101);
and U3317 (N_3317,N_2652,N_2594);
nand U3318 (N_3318,N_2277,N_2172);
and U3319 (N_3319,N_2151,N_2321);
nand U3320 (N_3320,N_2424,N_2451);
nor U3321 (N_3321,N_2512,N_2149);
nor U3322 (N_3322,N_2127,N_2963);
nand U3323 (N_3323,N_2533,N_2582);
nor U3324 (N_3324,N_2339,N_2129);
xor U3325 (N_3325,N_2638,N_2784);
or U3326 (N_3326,N_2752,N_2822);
or U3327 (N_3327,N_2111,N_2901);
and U3328 (N_3328,N_2635,N_2801);
nor U3329 (N_3329,N_2456,N_2391);
or U3330 (N_3330,N_2757,N_2857);
and U3331 (N_3331,N_2534,N_2448);
nor U3332 (N_3332,N_2889,N_2495);
xor U3333 (N_3333,N_2724,N_2494);
and U3334 (N_3334,N_2091,N_2953);
or U3335 (N_3335,N_2046,N_2891);
nand U3336 (N_3336,N_2722,N_2613);
nand U3337 (N_3337,N_2948,N_2038);
and U3338 (N_3338,N_2699,N_2812);
or U3339 (N_3339,N_2203,N_2192);
or U3340 (N_3340,N_2471,N_2729);
nand U3341 (N_3341,N_2663,N_2441);
or U3342 (N_3342,N_2483,N_2373);
xnor U3343 (N_3343,N_2331,N_2499);
nand U3344 (N_3344,N_2668,N_2622);
nand U3345 (N_3345,N_2693,N_2789);
and U3346 (N_3346,N_2440,N_2846);
and U3347 (N_3347,N_2393,N_2213);
nor U3348 (N_3348,N_2826,N_2104);
or U3349 (N_3349,N_2898,N_2163);
and U3350 (N_3350,N_2541,N_2027);
or U3351 (N_3351,N_2020,N_2198);
nor U3352 (N_3352,N_2019,N_2550);
nand U3353 (N_3353,N_2861,N_2676);
and U3354 (N_3354,N_2169,N_2766);
or U3355 (N_3355,N_2294,N_2654);
nand U3356 (N_3356,N_2770,N_2302);
xor U3357 (N_3357,N_2454,N_2641);
and U3358 (N_3358,N_2581,N_2873);
nand U3359 (N_3359,N_2968,N_2642);
xnor U3360 (N_3360,N_2379,N_2383);
or U3361 (N_3361,N_2392,N_2908);
nand U3362 (N_3362,N_2053,N_2031);
xnor U3363 (N_3363,N_2969,N_2627);
xor U3364 (N_3364,N_2606,N_2389);
or U3365 (N_3365,N_2160,N_2527);
nor U3366 (N_3366,N_2186,N_2524);
nand U3367 (N_3367,N_2661,N_2681);
nor U3368 (N_3368,N_2764,N_2918);
nor U3369 (N_3369,N_2369,N_2484);
nand U3370 (N_3370,N_2007,N_2942);
xor U3371 (N_3371,N_2061,N_2298);
nand U3372 (N_3372,N_2552,N_2474);
or U3373 (N_3373,N_2183,N_2210);
nor U3374 (N_3374,N_2200,N_2646);
xnor U3375 (N_3375,N_2911,N_2882);
or U3376 (N_3376,N_2879,N_2106);
xor U3377 (N_3377,N_2702,N_2999);
or U3378 (N_3378,N_2374,N_2986);
or U3379 (N_3379,N_2338,N_2481);
or U3380 (N_3380,N_2542,N_2470);
xnor U3381 (N_3381,N_2830,N_2006);
nand U3382 (N_3382,N_2604,N_2561);
or U3383 (N_3383,N_2009,N_2486);
or U3384 (N_3384,N_2436,N_2366);
nand U3385 (N_3385,N_2376,N_2572);
nand U3386 (N_3386,N_2427,N_2842);
nand U3387 (N_3387,N_2286,N_2493);
xnor U3388 (N_3388,N_2619,N_2887);
and U3389 (N_3389,N_2586,N_2591);
and U3390 (N_3390,N_2306,N_2344);
nor U3391 (N_3391,N_2354,N_2790);
xnor U3392 (N_3392,N_2793,N_2551);
and U3393 (N_3393,N_2975,N_2015);
nand U3394 (N_3394,N_2792,N_2446);
xor U3395 (N_3395,N_2989,N_2608);
xor U3396 (N_3396,N_2308,N_2040);
xnor U3397 (N_3397,N_2964,N_2437);
and U3398 (N_3398,N_2388,N_2951);
or U3399 (N_3399,N_2629,N_2760);
nand U3400 (N_3400,N_2946,N_2132);
nor U3401 (N_3401,N_2291,N_2831);
nand U3402 (N_3402,N_2670,N_2054);
and U3403 (N_3403,N_2759,N_2343);
and U3404 (N_3404,N_2904,N_2508);
nor U3405 (N_3405,N_2387,N_2311);
xor U3406 (N_3406,N_2008,N_2923);
nand U3407 (N_3407,N_2788,N_2706);
nor U3408 (N_3408,N_2491,N_2775);
xnor U3409 (N_3409,N_2753,N_2637);
xor U3410 (N_3410,N_2240,N_2390);
nand U3411 (N_3411,N_2457,N_2643);
nor U3412 (N_3412,N_2971,N_2434);
nand U3413 (N_3413,N_2478,N_2330);
nand U3414 (N_3414,N_2255,N_2182);
nand U3415 (N_3415,N_2337,N_2783);
xnor U3416 (N_3416,N_2595,N_2909);
nor U3417 (N_3417,N_2407,N_2938);
nand U3418 (N_3418,N_2916,N_2798);
nor U3419 (N_3419,N_2988,N_2328);
and U3420 (N_3420,N_2400,N_2636);
nor U3421 (N_3421,N_2075,N_2333);
nand U3422 (N_3422,N_2639,N_2985);
and U3423 (N_3423,N_2905,N_2858);
xor U3424 (N_3424,N_2231,N_2597);
xnor U3425 (N_3425,N_2628,N_2496);
or U3426 (N_3426,N_2991,N_2024);
or U3427 (N_3427,N_2810,N_2940);
nor U3428 (N_3428,N_2691,N_2647);
xnor U3429 (N_3429,N_2747,N_2531);
xnor U3430 (N_3430,N_2730,N_2065);
nand U3431 (N_3431,N_2219,N_2482);
and U3432 (N_3432,N_2781,N_2194);
nor U3433 (N_3433,N_2488,N_2967);
nand U3434 (N_3434,N_2059,N_2460);
nor U3435 (N_3435,N_2404,N_2233);
nor U3436 (N_3436,N_2095,N_2211);
nand U3437 (N_3437,N_2342,N_2941);
or U3438 (N_3438,N_2841,N_2207);
and U3439 (N_3439,N_2659,N_2375);
xnor U3440 (N_3440,N_2763,N_2935);
nor U3441 (N_3441,N_2782,N_2480);
and U3442 (N_3442,N_2257,N_2010);
nor U3443 (N_3443,N_2253,N_2155);
or U3444 (N_3444,N_2576,N_2171);
nor U3445 (N_3445,N_2979,N_2168);
nand U3446 (N_3446,N_2465,N_2624);
xor U3447 (N_3447,N_2051,N_2579);
nand U3448 (N_3448,N_2034,N_2609);
xnor U3449 (N_3449,N_2326,N_2944);
and U3450 (N_3450,N_2868,N_2709);
nand U3451 (N_3451,N_2398,N_2241);
xnor U3452 (N_3452,N_2382,N_2097);
nand U3453 (N_3453,N_2939,N_2745);
and U3454 (N_3454,N_2068,N_2547);
xnor U3455 (N_3455,N_2860,N_2204);
nor U3456 (N_3456,N_2883,N_2518);
xor U3457 (N_3457,N_2885,N_2452);
xnor U3458 (N_3458,N_2513,N_2123);
xnor U3459 (N_3459,N_2811,N_2094);
xnor U3460 (N_3460,N_2238,N_2334);
nand U3461 (N_3461,N_2717,N_2107);
xnor U3462 (N_3462,N_2884,N_2074);
and U3463 (N_3463,N_2394,N_2112);
xor U3464 (N_3464,N_2816,N_2538);
nor U3465 (N_3465,N_2467,N_2215);
and U3466 (N_3466,N_2144,N_2284);
xor U3467 (N_3467,N_2025,N_2158);
and U3468 (N_3468,N_2147,N_2087);
xor U3469 (N_3469,N_2318,N_2431);
or U3470 (N_3470,N_2825,N_2694);
or U3471 (N_3471,N_2234,N_2555);
nand U3472 (N_3472,N_2850,N_2599);
nand U3473 (N_3473,N_2756,N_2704);
and U3474 (N_3474,N_2304,N_2567);
or U3475 (N_3475,N_2256,N_2349);
or U3476 (N_3476,N_2381,N_2565);
nor U3477 (N_3477,N_2250,N_2573);
nor U3478 (N_3478,N_2577,N_2103);
nor U3479 (N_3479,N_2566,N_2157);
xnor U3480 (N_3480,N_2590,N_2212);
or U3481 (N_3481,N_2698,N_2917);
or U3482 (N_3482,N_2299,N_2554);
nand U3483 (N_3483,N_2352,N_2295);
xor U3484 (N_3484,N_2517,N_2412);
and U3485 (N_3485,N_2113,N_2854);
xnor U3486 (N_3486,N_2023,N_2718);
or U3487 (N_3487,N_2409,N_2743);
or U3488 (N_3488,N_2716,N_2921);
xnor U3489 (N_3489,N_2507,N_2931);
nand U3490 (N_3490,N_2529,N_2014);
nand U3491 (N_3491,N_2689,N_2589);
and U3492 (N_3492,N_2796,N_2876);
and U3493 (N_3493,N_2703,N_2558);
or U3494 (N_3494,N_2856,N_2947);
or U3495 (N_3495,N_2267,N_2247);
nor U3496 (N_3496,N_2313,N_2426);
and U3497 (N_3497,N_2175,N_2848);
or U3498 (N_3498,N_2922,N_2708);
nor U3499 (N_3499,N_2140,N_2041);
xnor U3500 (N_3500,N_2539,N_2981);
and U3501 (N_3501,N_2715,N_2512);
nor U3502 (N_3502,N_2279,N_2972);
nor U3503 (N_3503,N_2656,N_2345);
xor U3504 (N_3504,N_2457,N_2603);
xnor U3505 (N_3505,N_2001,N_2271);
nand U3506 (N_3506,N_2102,N_2609);
or U3507 (N_3507,N_2905,N_2327);
xor U3508 (N_3508,N_2359,N_2737);
xor U3509 (N_3509,N_2073,N_2487);
xnor U3510 (N_3510,N_2369,N_2396);
xor U3511 (N_3511,N_2143,N_2212);
nand U3512 (N_3512,N_2789,N_2397);
xor U3513 (N_3513,N_2827,N_2696);
nor U3514 (N_3514,N_2106,N_2064);
nor U3515 (N_3515,N_2346,N_2989);
xnor U3516 (N_3516,N_2140,N_2366);
and U3517 (N_3517,N_2516,N_2649);
xor U3518 (N_3518,N_2358,N_2400);
or U3519 (N_3519,N_2626,N_2811);
nand U3520 (N_3520,N_2790,N_2333);
xnor U3521 (N_3521,N_2952,N_2197);
xnor U3522 (N_3522,N_2518,N_2685);
and U3523 (N_3523,N_2031,N_2404);
or U3524 (N_3524,N_2461,N_2708);
xnor U3525 (N_3525,N_2175,N_2904);
or U3526 (N_3526,N_2819,N_2915);
nor U3527 (N_3527,N_2662,N_2830);
nand U3528 (N_3528,N_2662,N_2931);
nor U3529 (N_3529,N_2400,N_2428);
nand U3530 (N_3530,N_2199,N_2164);
or U3531 (N_3531,N_2891,N_2115);
nor U3532 (N_3532,N_2446,N_2873);
xor U3533 (N_3533,N_2002,N_2798);
nand U3534 (N_3534,N_2158,N_2828);
and U3535 (N_3535,N_2532,N_2927);
and U3536 (N_3536,N_2564,N_2650);
xor U3537 (N_3537,N_2785,N_2361);
nand U3538 (N_3538,N_2412,N_2614);
or U3539 (N_3539,N_2238,N_2188);
nor U3540 (N_3540,N_2737,N_2524);
nand U3541 (N_3541,N_2491,N_2728);
nand U3542 (N_3542,N_2234,N_2599);
xor U3543 (N_3543,N_2731,N_2011);
nand U3544 (N_3544,N_2809,N_2387);
and U3545 (N_3545,N_2426,N_2554);
or U3546 (N_3546,N_2047,N_2356);
nor U3547 (N_3547,N_2595,N_2527);
nand U3548 (N_3548,N_2937,N_2882);
xnor U3549 (N_3549,N_2152,N_2191);
nand U3550 (N_3550,N_2639,N_2092);
or U3551 (N_3551,N_2130,N_2294);
nor U3552 (N_3552,N_2822,N_2028);
or U3553 (N_3553,N_2242,N_2307);
nor U3554 (N_3554,N_2929,N_2989);
nand U3555 (N_3555,N_2076,N_2884);
nand U3556 (N_3556,N_2722,N_2180);
nand U3557 (N_3557,N_2651,N_2291);
nand U3558 (N_3558,N_2333,N_2872);
nor U3559 (N_3559,N_2190,N_2332);
or U3560 (N_3560,N_2465,N_2466);
xor U3561 (N_3561,N_2196,N_2801);
or U3562 (N_3562,N_2958,N_2126);
and U3563 (N_3563,N_2432,N_2368);
or U3564 (N_3564,N_2674,N_2131);
xnor U3565 (N_3565,N_2239,N_2230);
and U3566 (N_3566,N_2279,N_2206);
or U3567 (N_3567,N_2751,N_2510);
nand U3568 (N_3568,N_2755,N_2568);
xor U3569 (N_3569,N_2106,N_2184);
xor U3570 (N_3570,N_2842,N_2185);
or U3571 (N_3571,N_2386,N_2986);
nor U3572 (N_3572,N_2986,N_2491);
nand U3573 (N_3573,N_2135,N_2802);
xnor U3574 (N_3574,N_2149,N_2847);
nand U3575 (N_3575,N_2174,N_2440);
nor U3576 (N_3576,N_2653,N_2763);
xnor U3577 (N_3577,N_2601,N_2882);
nand U3578 (N_3578,N_2220,N_2392);
xor U3579 (N_3579,N_2431,N_2309);
nand U3580 (N_3580,N_2219,N_2913);
nand U3581 (N_3581,N_2765,N_2540);
nor U3582 (N_3582,N_2423,N_2855);
and U3583 (N_3583,N_2633,N_2385);
or U3584 (N_3584,N_2703,N_2010);
nor U3585 (N_3585,N_2867,N_2897);
or U3586 (N_3586,N_2450,N_2235);
or U3587 (N_3587,N_2206,N_2651);
and U3588 (N_3588,N_2312,N_2209);
nand U3589 (N_3589,N_2398,N_2598);
nand U3590 (N_3590,N_2884,N_2360);
nand U3591 (N_3591,N_2874,N_2154);
and U3592 (N_3592,N_2424,N_2727);
nand U3593 (N_3593,N_2422,N_2543);
and U3594 (N_3594,N_2702,N_2408);
xnor U3595 (N_3595,N_2689,N_2846);
and U3596 (N_3596,N_2204,N_2852);
xnor U3597 (N_3597,N_2789,N_2241);
or U3598 (N_3598,N_2422,N_2934);
xor U3599 (N_3599,N_2943,N_2464);
and U3600 (N_3600,N_2122,N_2948);
xnor U3601 (N_3601,N_2516,N_2586);
and U3602 (N_3602,N_2310,N_2717);
or U3603 (N_3603,N_2153,N_2110);
nor U3604 (N_3604,N_2603,N_2872);
and U3605 (N_3605,N_2968,N_2412);
and U3606 (N_3606,N_2951,N_2517);
or U3607 (N_3607,N_2121,N_2098);
and U3608 (N_3608,N_2555,N_2799);
nand U3609 (N_3609,N_2742,N_2345);
xor U3610 (N_3610,N_2728,N_2059);
and U3611 (N_3611,N_2415,N_2269);
or U3612 (N_3612,N_2913,N_2972);
nor U3613 (N_3613,N_2194,N_2551);
or U3614 (N_3614,N_2420,N_2201);
nand U3615 (N_3615,N_2384,N_2991);
nor U3616 (N_3616,N_2282,N_2818);
or U3617 (N_3617,N_2214,N_2904);
xor U3618 (N_3618,N_2620,N_2798);
and U3619 (N_3619,N_2788,N_2054);
or U3620 (N_3620,N_2442,N_2711);
nor U3621 (N_3621,N_2255,N_2871);
and U3622 (N_3622,N_2514,N_2481);
or U3623 (N_3623,N_2424,N_2200);
or U3624 (N_3624,N_2311,N_2925);
or U3625 (N_3625,N_2904,N_2778);
and U3626 (N_3626,N_2403,N_2369);
or U3627 (N_3627,N_2242,N_2222);
xor U3628 (N_3628,N_2511,N_2294);
and U3629 (N_3629,N_2500,N_2919);
and U3630 (N_3630,N_2585,N_2893);
or U3631 (N_3631,N_2311,N_2916);
nor U3632 (N_3632,N_2199,N_2060);
or U3633 (N_3633,N_2177,N_2662);
nor U3634 (N_3634,N_2278,N_2545);
xor U3635 (N_3635,N_2630,N_2043);
or U3636 (N_3636,N_2792,N_2182);
nor U3637 (N_3637,N_2333,N_2618);
or U3638 (N_3638,N_2921,N_2939);
and U3639 (N_3639,N_2712,N_2620);
nor U3640 (N_3640,N_2599,N_2233);
xnor U3641 (N_3641,N_2229,N_2262);
and U3642 (N_3642,N_2145,N_2325);
xnor U3643 (N_3643,N_2945,N_2953);
or U3644 (N_3644,N_2000,N_2365);
nor U3645 (N_3645,N_2979,N_2192);
or U3646 (N_3646,N_2469,N_2650);
or U3647 (N_3647,N_2477,N_2870);
or U3648 (N_3648,N_2629,N_2871);
or U3649 (N_3649,N_2401,N_2269);
and U3650 (N_3650,N_2108,N_2624);
and U3651 (N_3651,N_2096,N_2406);
xnor U3652 (N_3652,N_2071,N_2871);
or U3653 (N_3653,N_2389,N_2013);
nand U3654 (N_3654,N_2582,N_2045);
nand U3655 (N_3655,N_2612,N_2356);
nor U3656 (N_3656,N_2467,N_2475);
and U3657 (N_3657,N_2795,N_2409);
or U3658 (N_3658,N_2337,N_2673);
xor U3659 (N_3659,N_2126,N_2837);
nand U3660 (N_3660,N_2158,N_2864);
or U3661 (N_3661,N_2506,N_2992);
nor U3662 (N_3662,N_2648,N_2402);
nand U3663 (N_3663,N_2695,N_2983);
or U3664 (N_3664,N_2486,N_2432);
and U3665 (N_3665,N_2674,N_2819);
and U3666 (N_3666,N_2667,N_2391);
xor U3667 (N_3667,N_2868,N_2153);
or U3668 (N_3668,N_2535,N_2131);
and U3669 (N_3669,N_2602,N_2702);
xnor U3670 (N_3670,N_2867,N_2472);
xor U3671 (N_3671,N_2045,N_2147);
xor U3672 (N_3672,N_2716,N_2909);
nor U3673 (N_3673,N_2743,N_2686);
and U3674 (N_3674,N_2869,N_2843);
nand U3675 (N_3675,N_2586,N_2121);
and U3676 (N_3676,N_2596,N_2103);
or U3677 (N_3677,N_2172,N_2022);
and U3678 (N_3678,N_2684,N_2141);
nor U3679 (N_3679,N_2231,N_2932);
nor U3680 (N_3680,N_2762,N_2410);
xnor U3681 (N_3681,N_2163,N_2365);
xnor U3682 (N_3682,N_2795,N_2481);
and U3683 (N_3683,N_2829,N_2562);
or U3684 (N_3684,N_2702,N_2246);
nand U3685 (N_3685,N_2792,N_2602);
nor U3686 (N_3686,N_2696,N_2745);
or U3687 (N_3687,N_2420,N_2004);
nor U3688 (N_3688,N_2744,N_2755);
or U3689 (N_3689,N_2720,N_2989);
xnor U3690 (N_3690,N_2157,N_2232);
nand U3691 (N_3691,N_2246,N_2201);
xnor U3692 (N_3692,N_2546,N_2393);
or U3693 (N_3693,N_2001,N_2787);
nand U3694 (N_3694,N_2157,N_2025);
nor U3695 (N_3695,N_2195,N_2521);
xnor U3696 (N_3696,N_2658,N_2337);
nand U3697 (N_3697,N_2847,N_2512);
and U3698 (N_3698,N_2161,N_2531);
xor U3699 (N_3699,N_2630,N_2718);
xnor U3700 (N_3700,N_2498,N_2585);
nor U3701 (N_3701,N_2310,N_2453);
or U3702 (N_3702,N_2586,N_2874);
or U3703 (N_3703,N_2181,N_2313);
xor U3704 (N_3704,N_2656,N_2742);
nor U3705 (N_3705,N_2798,N_2702);
nand U3706 (N_3706,N_2674,N_2411);
and U3707 (N_3707,N_2853,N_2821);
nor U3708 (N_3708,N_2788,N_2316);
xnor U3709 (N_3709,N_2466,N_2374);
or U3710 (N_3710,N_2043,N_2679);
xor U3711 (N_3711,N_2291,N_2351);
and U3712 (N_3712,N_2654,N_2950);
or U3713 (N_3713,N_2085,N_2568);
xnor U3714 (N_3714,N_2509,N_2003);
or U3715 (N_3715,N_2750,N_2997);
or U3716 (N_3716,N_2392,N_2407);
nand U3717 (N_3717,N_2948,N_2307);
or U3718 (N_3718,N_2515,N_2353);
and U3719 (N_3719,N_2536,N_2493);
nand U3720 (N_3720,N_2825,N_2265);
xor U3721 (N_3721,N_2314,N_2129);
and U3722 (N_3722,N_2848,N_2636);
and U3723 (N_3723,N_2892,N_2560);
or U3724 (N_3724,N_2903,N_2517);
nand U3725 (N_3725,N_2951,N_2528);
or U3726 (N_3726,N_2491,N_2037);
nor U3727 (N_3727,N_2201,N_2581);
or U3728 (N_3728,N_2089,N_2435);
nand U3729 (N_3729,N_2514,N_2128);
and U3730 (N_3730,N_2035,N_2441);
nor U3731 (N_3731,N_2305,N_2964);
nor U3732 (N_3732,N_2234,N_2043);
xor U3733 (N_3733,N_2319,N_2331);
or U3734 (N_3734,N_2626,N_2387);
or U3735 (N_3735,N_2930,N_2826);
or U3736 (N_3736,N_2933,N_2722);
xor U3737 (N_3737,N_2622,N_2784);
xor U3738 (N_3738,N_2289,N_2522);
xor U3739 (N_3739,N_2467,N_2680);
and U3740 (N_3740,N_2916,N_2578);
or U3741 (N_3741,N_2666,N_2830);
xor U3742 (N_3742,N_2409,N_2192);
nor U3743 (N_3743,N_2963,N_2589);
and U3744 (N_3744,N_2948,N_2959);
nand U3745 (N_3745,N_2884,N_2832);
or U3746 (N_3746,N_2325,N_2980);
xnor U3747 (N_3747,N_2573,N_2411);
xor U3748 (N_3748,N_2820,N_2505);
nand U3749 (N_3749,N_2370,N_2834);
or U3750 (N_3750,N_2866,N_2153);
nand U3751 (N_3751,N_2495,N_2219);
nand U3752 (N_3752,N_2800,N_2034);
xor U3753 (N_3753,N_2941,N_2989);
xor U3754 (N_3754,N_2881,N_2437);
or U3755 (N_3755,N_2590,N_2420);
or U3756 (N_3756,N_2135,N_2579);
nand U3757 (N_3757,N_2867,N_2674);
and U3758 (N_3758,N_2227,N_2403);
xnor U3759 (N_3759,N_2873,N_2362);
nand U3760 (N_3760,N_2953,N_2237);
or U3761 (N_3761,N_2379,N_2303);
nand U3762 (N_3762,N_2228,N_2458);
or U3763 (N_3763,N_2765,N_2725);
and U3764 (N_3764,N_2863,N_2029);
xor U3765 (N_3765,N_2458,N_2589);
or U3766 (N_3766,N_2086,N_2113);
xnor U3767 (N_3767,N_2683,N_2491);
nand U3768 (N_3768,N_2451,N_2166);
xnor U3769 (N_3769,N_2873,N_2247);
xor U3770 (N_3770,N_2075,N_2731);
and U3771 (N_3771,N_2763,N_2675);
nor U3772 (N_3772,N_2018,N_2889);
or U3773 (N_3773,N_2020,N_2526);
nor U3774 (N_3774,N_2269,N_2287);
nor U3775 (N_3775,N_2297,N_2909);
nor U3776 (N_3776,N_2947,N_2269);
and U3777 (N_3777,N_2092,N_2948);
or U3778 (N_3778,N_2603,N_2750);
and U3779 (N_3779,N_2785,N_2001);
nor U3780 (N_3780,N_2227,N_2745);
and U3781 (N_3781,N_2888,N_2128);
xor U3782 (N_3782,N_2289,N_2523);
or U3783 (N_3783,N_2717,N_2653);
nor U3784 (N_3784,N_2296,N_2883);
and U3785 (N_3785,N_2645,N_2334);
xnor U3786 (N_3786,N_2457,N_2434);
and U3787 (N_3787,N_2894,N_2845);
nand U3788 (N_3788,N_2173,N_2265);
nand U3789 (N_3789,N_2259,N_2990);
nor U3790 (N_3790,N_2595,N_2137);
and U3791 (N_3791,N_2264,N_2726);
nand U3792 (N_3792,N_2444,N_2003);
xor U3793 (N_3793,N_2488,N_2561);
nand U3794 (N_3794,N_2624,N_2702);
and U3795 (N_3795,N_2804,N_2710);
nand U3796 (N_3796,N_2914,N_2311);
xor U3797 (N_3797,N_2909,N_2074);
nor U3798 (N_3798,N_2618,N_2484);
nand U3799 (N_3799,N_2636,N_2256);
nor U3800 (N_3800,N_2380,N_2024);
nand U3801 (N_3801,N_2428,N_2999);
and U3802 (N_3802,N_2440,N_2965);
and U3803 (N_3803,N_2230,N_2969);
nand U3804 (N_3804,N_2665,N_2989);
nor U3805 (N_3805,N_2164,N_2781);
and U3806 (N_3806,N_2142,N_2686);
xnor U3807 (N_3807,N_2941,N_2690);
nor U3808 (N_3808,N_2715,N_2983);
and U3809 (N_3809,N_2034,N_2180);
xor U3810 (N_3810,N_2529,N_2081);
nor U3811 (N_3811,N_2843,N_2076);
nand U3812 (N_3812,N_2001,N_2852);
or U3813 (N_3813,N_2709,N_2079);
and U3814 (N_3814,N_2267,N_2356);
and U3815 (N_3815,N_2952,N_2639);
or U3816 (N_3816,N_2187,N_2761);
nand U3817 (N_3817,N_2936,N_2637);
or U3818 (N_3818,N_2053,N_2552);
nand U3819 (N_3819,N_2943,N_2072);
and U3820 (N_3820,N_2036,N_2678);
or U3821 (N_3821,N_2136,N_2510);
and U3822 (N_3822,N_2799,N_2166);
xnor U3823 (N_3823,N_2693,N_2649);
nand U3824 (N_3824,N_2019,N_2853);
xor U3825 (N_3825,N_2786,N_2633);
nor U3826 (N_3826,N_2971,N_2326);
xor U3827 (N_3827,N_2010,N_2416);
nor U3828 (N_3828,N_2709,N_2486);
and U3829 (N_3829,N_2125,N_2080);
and U3830 (N_3830,N_2139,N_2178);
and U3831 (N_3831,N_2348,N_2531);
or U3832 (N_3832,N_2505,N_2054);
and U3833 (N_3833,N_2130,N_2487);
and U3834 (N_3834,N_2177,N_2033);
xor U3835 (N_3835,N_2909,N_2994);
nor U3836 (N_3836,N_2821,N_2653);
nand U3837 (N_3837,N_2654,N_2621);
xor U3838 (N_3838,N_2724,N_2617);
and U3839 (N_3839,N_2258,N_2339);
nand U3840 (N_3840,N_2932,N_2042);
and U3841 (N_3841,N_2662,N_2806);
nor U3842 (N_3842,N_2587,N_2136);
nor U3843 (N_3843,N_2902,N_2723);
xor U3844 (N_3844,N_2696,N_2476);
xor U3845 (N_3845,N_2118,N_2437);
and U3846 (N_3846,N_2019,N_2059);
nor U3847 (N_3847,N_2480,N_2395);
nor U3848 (N_3848,N_2018,N_2973);
nand U3849 (N_3849,N_2553,N_2228);
and U3850 (N_3850,N_2184,N_2154);
or U3851 (N_3851,N_2476,N_2202);
nor U3852 (N_3852,N_2742,N_2337);
nand U3853 (N_3853,N_2333,N_2118);
nor U3854 (N_3854,N_2826,N_2555);
or U3855 (N_3855,N_2044,N_2489);
xnor U3856 (N_3856,N_2157,N_2715);
xor U3857 (N_3857,N_2171,N_2080);
nor U3858 (N_3858,N_2632,N_2859);
and U3859 (N_3859,N_2478,N_2535);
nor U3860 (N_3860,N_2149,N_2179);
and U3861 (N_3861,N_2083,N_2421);
xnor U3862 (N_3862,N_2464,N_2553);
nand U3863 (N_3863,N_2697,N_2986);
and U3864 (N_3864,N_2539,N_2994);
nand U3865 (N_3865,N_2453,N_2280);
nand U3866 (N_3866,N_2457,N_2502);
and U3867 (N_3867,N_2250,N_2818);
nor U3868 (N_3868,N_2321,N_2012);
nor U3869 (N_3869,N_2090,N_2340);
or U3870 (N_3870,N_2938,N_2771);
xnor U3871 (N_3871,N_2044,N_2040);
and U3872 (N_3872,N_2605,N_2680);
xnor U3873 (N_3873,N_2048,N_2463);
xnor U3874 (N_3874,N_2593,N_2282);
nor U3875 (N_3875,N_2832,N_2804);
or U3876 (N_3876,N_2971,N_2096);
or U3877 (N_3877,N_2804,N_2822);
xnor U3878 (N_3878,N_2745,N_2087);
and U3879 (N_3879,N_2469,N_2167);
nor U3880 (N_3880,N_2644,N_2211);
nand U3881 (N_3881,N_2669,N_2122);
and U3882 (N_3882,N_2354,N_2480);
nor U3883 (N_3883,N_2501,N_2130);
nand U3884 (N_3884,N_2993,N_2515);
nor U3885 (N_3885,N_2775,N_2414);
and U3886 (N_3886,N_2379,N_2733);
xor U3887 (N_3887,N_2491,N_2643);
or U3888 (N_3888,N_2390,N_2976);
and U3889 (N_3889,N_2520,N_2110);
and U3890 (N_3890,N_2997,N_2651);
or U3891 (N_3891,N_2185,N_2320);
nand U3892 (N_3892,N_2253,N_2882);
or U3893 (N_3893,N_2409,N_2089);
and U3894 (N_3894,N_2840,N_2957);
or U3895 (N_3895,N_2385,N_2306);
xor U3896 (N_3896,N_2717,N_2868);
or U3897 (N_3897,N_2445,N_2220);
or U3898 (N_3898,N_2852,N_2837);
nor U3899 (N_3899,N_2681,N_2018);
xor U3900 (N_3900,N_2223,N_2840);
xnor U3901 (N_3901,N_2207,N_2220);
and U3902 (N_3902,N_2029,N_2150);
nand U3903 (N_3903,N_2459,N_2630);
nor U3904 (N_3904,N_2773,N_2697);
and U3905 (N_3905,N_2091,N_2999);
nor U3906 (N_3906,N_2667,N_2366);
nand U3907 (N_3907,N_2538,N_2912);
nor U3908 (N_3908,N_2689,N_2985);
and U3909 (N_3909,N_2746,N_2421);
nand U3910 (N_3910,N_2627,N_2871);
xnor U3911 (N_3911,N_2028,N_2703);
nand U3912 (N_3912,N_2576,N_2059);
nand U3913 (N_3913,N_2417,N_2390);
and U3914 (N_3914,N_2478,N_2009);
and U3915 (N_3915,N_2934,N_2342);
xnor U3916 (N_3916,N_2912,N_2120);
nand U3917 (N_3917,N_2794,N_2619);
or U3918 (N_3918,N_2994,N_2514);
xor U3919 (N_3919,N_2038,N_2632);
or U3920 (N_3920,N_2091,N_2142);
nand U3921 (N_3921,N_2052,N_2385);
nor U3922 (N_3922,N_2952,N_2065);
nor U3923 (N_3923,N_2395,N_2120);
nand U3924 (N_3924,N_2795,N_2597);
nor U3925 (N_3925,N_2536,N_2909);
or U3926 (N_3926,N_2222,N_2728);
nor U3927 (N_3927,N_2690,N_2843);
xnor U3928 (N_3928,N_2300,N_2492);
or U3929 (N_3929,N_2488,N_2790);
nor U3930 (N_3930,N_2896,N_2169);
nor U3931 (N_3931,N_2867,N_2846);
xnor U3932 (N_3932,N_2898,N_2494);
xnor U3933 (N_3933,N_2380,N_2364);
or U3934 (N_3934,N_2470,N_2525);
nor U3935 (N_3935,N_2120,N_2108);
nor U3936 (N_3936,N_2188,N_2792);
nor U3937 (N_3937,N_2236,N_2092);
or U3938 (N_3938,N_2646,N_2389);
xor U3939 (N_3939,N_2068,N_2184);
xor U3940 (N_3940,N_2127,N_2476);
xnor U3941 (N_3941,N_2058,N_2391);
nand U3942 (N_3942,N_2877,N_2248);
nand U3943 (N_3943,N_2713,N_2394);
xnor U3944 (N_3944,N_2143,N_2349);
or U3945 (N_3945,N_2877,N_2788);
or U3946 (N_3946,N_2832,N_2280);
and U3947 (N_3947,N_2706,N_2025);
nor U3948 (N_3948,N_2248,N_2695);
and U3949 (N_3949,N_2650,N_2676);
nand U3950 (N_3950,N_2195,N_2128);
nand U3951 (N_3951,N_2718,N_2507);
nand U3952 (N_3952,N_2354,N_2481);
nor U3953 (N_3953,N_2853,N_2826);
nor U3954 (N_3954,N_2929,N_2892);
xnor U3955 (N_3955,N_2052,N_2458);
nand U3956 (N_3956,N_2181,N_2936);
xor U3957 (N_3957,N_2418,N_2815);
nand U3958 (N_3958,N_2801,N_2490);
or U3959 (N_3959,N_2425,N_2587);
xnor U3960 (N_3960,N_2404,N_2737);
nor U3961 (N_3961,N_2706,N_2564);
nor U3962 (N_3962,N_2683,N_2035);
or U3963 (N_3963,N_2930,N_2862);
or U3964 (N_3964,N_2830,N_2488);
nor U3965 (N_3965,N_2510,N_2410);
and U3966 (N_3966,N_2731,N_2551);
or U3967 (N_3967,N_2304,N_2677);
or U3968 (N_3968,N_2803,N_2868);
xor U3969 (N_3969,N_2086,N_2731);
xnor U3970 (N_3970,N_2388,N_2210);
or U3971 (N_3971,N_2140,N_2528);
xnor U3972 (N_3972,N_2429,N_2299);
or U3973 (N_3973,N_2802,N_2050);
and U3974 (N_3974,N_2955,N_2289);
nand U3975 (N_3975,N_2317,N_2592);
and U3976 (N_3976,N_2071,N_2236);
nor U3977 (N_3977,N_2237,N_2720);
or U3978 (N_3978,N_2484,N_2711);
and U3979 (N_3979,N_2822,N_2307);
and U3980 (N_3980,N_2568,N_2521);
and U3981 (N_3981,N_2080,N_2027);
nor U3982 (N_3982,N_2146,N_2274);
nor U3983 (N_3983,N_2390,N_2179);
or U3984 (N_3984,N_2756,N_2845);
or U3985 (N_3985,N_2617,N_2532);
and U3986 (N_3986,N_2781,N_2517);
or U3987 (N_3987,N_2539,N_2036);
nor U3988 (N_3988,N_2302,N_2253);
xnor U3989 (N_3989,N_2204,N_2953);
xnor U3990 (N_3990,N_2315,N_2443);
or U3991 (N_3991,N_2963,N_2895);
nor U3992 (N_3992,N_2550,N_2987);
nand U3993 (N_3993,N_2749,N_2867);
nor U3994 (N_3994,N_2926,N_2304);
and U3995 (N_3995,N_2042,N_2396);
nor U3996 (N_3996,N_2733,N_2143);
nand U3997 (N_3997,N_2624,N_2276);
or U3998 (N_3998,N_2976,N_2250);
nand U3999 (N_3999,N_2648,N_2206);
and U4000 (N_4000,N_3912,N_3309);
and U4001 (N_4001,N_3884,N_3272);
or U4002 (N_4002,N_3337,N_3896);
or U4003 (N_4003,N_3778,N_3098);
and U4004 (N_4004,N_3161,N_3878);
or U4005 (N_4005,N_3027,N_3106);
nor U4006 (N_4006,N_3274,N_3495);
xnor U4007 (N_4007,N_3904,N_3548);
xnor U4008 (N_4008,N_3389,N_3002);
xnor U4009 (N_4009,N_3568,N_3544);
xnor U4010 (N_4010,N_3866,N_3244);
and U4011 (N_4011,N_3783,N_3019);
xnor U4012 (N_4012,N_3761,N_3901);
nand U4013 (N_4013,N_3643,N_3746);
and U4014 (N_4014,N_3753,N_3676);
xnor U4015 (N_4015,N_3805,N_3793);
nor U4016 (N_4016,N_3391,N_3048);
or U4017 (N_4017,N_3420,N_3013);
xor U4018 (N_4018,N_3821,N_3807);
xnor U4019 (N_4019,N_3102,N_3942);
nand U4020 (N_4020,N_3026,N_3311);
or U4021 (N_4021,N_3641,N_3701);
and U4022 (N_4022,N_3278,N_3613);
or U4023 (N_4023,N_3677,N_3922);
or U4024 (N_4024,N_3361,N_3642);
or U4025 (N_4025,N_3340,N_3018);
and U4026 (N_4026,N_3044,N_3030);
or U4027 (N_4027,N_3740,N_3808);
nor U4028 (N_4028,N_3686,N_3584);
nor U4029 (N_4029,N_3464,N_3304);
or U4030 (N_4030,N_3656,N_3933);
or U4031 (N_4031,N_3800,N_3806);
xor U4032 (N_4032,N_3528,N_3802);
nor U4033 (N_4033,N_3968,N_3338);
or U4034 (N_4034,N_3149,N_3332);
nand U4035 (N_4035,N_3313,N_3097);
nor U4036 (N_4036,N_3458,N_3981);
nor U4037 (N_4037,N_3356,N_3629);
nand U4038 (N_4038,N_3512,N_3813);
xnor U4039 (N_4039,N_3120,N_3185);
or U4040 (N_4040,N_3339,N_3427);
or U4041 (N_4041,N_3176,N_3985);
or U4042 (N_4042,N_3284,N_3854);
or U4043 (N_4043,N_3024,N_3556);
and U4044 (N_4044,N_3785,N_3654);
nand U4045 (N_4045,N_3868,N_3004);
or U4046 (N_4046,N_3328,N_3890);
nor U4047 (N_4047,N_3152,N_3763);
and U4048 (N_4048,N_3182,N_3877);
nand U4049 (N_4049,N_3704,N_3826);
nand U4050 (N_4050,N_3954,N_3381);
xnor U4051 (N_4051,N_3586,N_3333);
and U4052 (N_4052,N_3660,N_3798);
and U4053 (N_4053,N_3921,N_3727);
xnor U4054 (N_4054,N_3301,N_3545);
xnor U4055 (N_4055,N_3579,N_3809);
and U4056 (N_4056,N_3789,N_3914);
or U4057 (N_4057,N_3071,N_3407);
or U4058 (N_4058,N_3186,N_3526);
xor U4059 (N_4059,N_3036,N_3532);
xor U4060 (N_4060,N_3101,N_3497);
xor U4061 (N_4061,N_3860,N_3399);
nand U4062 (N_4062,N_3134,N_3293);
or U4063 (N_4063,N_3146,N_3855);
nand U4064 (N_4064,N_3370,N_3234);
nor U4065 (N_4065,N_3850,N_3983);
nor U4066 (N_4066,N_3553,N_3580);
nand U4067 (N_4067,N_3531,N_3283);
and U4068 (N_4068,N_3915,N_3111);
xnor U4069 (N_4069,N_3090,N_3961);
xor U4070 (N_4070,N_3198,N_3649);
and U4071 (N_4071,N_3977,N_3235);
xnor U4072 (N_4072,N_3817,N_3771);
xor U4073 (N_4073,N_3907,N_3958);
nand U4074 (N_4074,N_3716,N_3220);
nand U4075 (N_4075,N_3843,N_3379);
xor U4076 (N_4076,N_3687,N_3776);
or U4077 (N_4077,N_3721,N_3374);
xnor U4078 (N_4078,N_3412,N_3562);
nand U4079 (N_4079,N_3023,N_3314);
xnor U4080 (N_4080,N_3009,N_3992);
or U4081 (N_4081,N_3796,N_3558);
nand U4082 (N_4082,N_3836,N_3212);
and U4083 (N_4083,N_3765,N_3247);
xnor U4084 (N_4084,N_3588,N_3706);
nand U4085 (N_4085,N_3608,N_3870);
or U4086 (N_4086,N_3455,N_3975);
and U4087 (N_4087,N_3978,N_3717);
nand U4088 (N_4088,N_3066,N_3797);
xnor U4089 (N_4089,N_3167,N_3243);
xnor U4090 (N_4090,N_3910,N_3277);
nor U4091 (N_4091,N_3054,N_3335);
nand U4092 (N_4092,N_3668,N_3519);
and U4093 (N_4093,N_3856,N_3773);
xnor U4094 (N_4094,N_3296,N_3801);
or U4095 (N_4095,N_3100,N_3445);
xnor U4096 (N_4096,N_3260,N_3892);
nor U4097 (N_4097,N_3351,N_3903);
nand U4098 (N_4098,N_3779,N_3162);
or U4099 (N_4099,N_3061,N_3891);
nor U4100 (N_4100,N_3218,N_3722);
nor U4101 (N_4101,N_3818,N_3148);
xnor U4102 (N_4102,N_3297,N_3058);
nand U4103 (N_4103,N_3128,N_3124);
and U4104 (N_4104,N_3385,N_3893);
xnor U4105 (N_4105,N_3096,N_3040);
nand U4106 (N_4106,N_3122,N_3233);
nand U4107 (N_4107,N_3108,N_3117);
or U4108 (N_4108,N_3083,N_3137);
nand U4109 (N_4109,N_3675,N_3627);
xor U4110 (N_4110,N_3591,N_3095);
nor U4111 (N_4111,N_3460,N_3987);
or U4112 (N_4112,N_3499,N_3334);
nand U4113 (N_4113,N_3032,N_3959);
nand U4114 (N_4114,N_3909,N_3476);
and U4115 (N_4115,N_3368,N_3943);
or U4116 (N_4116,N_3245,N_3489);
xor U4117 (N_4117,N_3572,N_3459);
nand U4118 (N_4118,N_3209,N_3619);
nand U4119 (N_4119,N_3431,N_3841);
nand U4120 (N_4120,N_3863,N_3008);
and U4121 (N_4121,N_3515,N_3275);
and U4122 (N_4122,N_3631,N_3271);
or U4123 (N_4123,N_3190,N_3292);
and U4124 (N_4124,N_3485,N_3352);
or U4125 (N_4125,N_3270,N_3777);
or U4126 (N_4126,N_3127,N_3393);
xor U4127 (N_4127,N_3215,N_3211);
nor U4128 (N_4128,N_3593,N_3700);
and U4129 (N_4129,N_3355,N_3323);
or U4130 (N_4130,N_3669,N_3481);
or U4131 (N_4131,N_3538,N_3590);
xor U4132 (N_4132,N_3522,N_3897);
nor U4133 (N_4133,N_3187,N_3321);
nor U4134 (N_4134,N_3359,N_3782);
xor U4135 (N_4135,N_3599,N_3045);
xor U4136 (N_4136,N_3143,N_3409);
xor U4137 (N_4137,N_3224,N_3116);
xor U4138 (N_4138,N_3831,N_3344);
nor U4139 (N_4139,N_3630,N_3103);
nor U4140 (N_4140,N_3781,N_3421);
nand U4141 (N_4141,N_3307,N_3749);
nand U4142 (N_4142,N_3119,N_3029);
nor U4143 (N_4143,N_3960,N_3154);
or U4144 (N_4144,N_3442,N_3006);
and U4145 (N_4145,N_3788,N_3684);
or U4146 (N_4146,N_3436,N_3611);
and U4147 (N_4147,N_3932,N_3383);
or U4148 (N_4148,N_3074,N_3623);
and U4149 (N_4149,N_3560,N_3653);
xor U4150 (N_4150,N_3078,N_3035);
or U4151 (N_4151,N_3471,N_3620);
or U4152 (N_4152,N_3928,N_3714);
nor U4153 (N_4153,N_3663,N_3400);
nor U4154 (N_4154,N_3659,N_3829);
and U4155 (N_4155,N_3467,N_3624);
nand U4156 (N_4156,N_3741,N_3988);
or U4157 (N_4157,N_3636,N_3769);
nand U4158 (N_4158,N_3726,N_3944);
nand U4159 (N_4159,N_3573,N_3707);
and U4160 (N_4160,N_3839,N_3482);
or U4161 (N_4161,N_3305,N_3377);
or U4162 (N_4162,N_3824,N_3563);
nor U4163 (N_4163,N_3589,N_3709);
nor U4164 (N_4164,N_3658,N_3804);
xnor U4165 (N_4165,N_3888,N_3193);
and U4166 (N_4166,N_3632,N_3229);
nand U4167 (N_4167,N_3937,N_3533);
or U4168 (N_4168,N_3052,N_3894);
and U4169 (N_4169,N_3444,N_3085);
nand U4170 (N_4170,N_3766,N_3419);
and U4171 (N_4171,N_3174,N_3129);
xor U4172 (N_4172,N_3175,N_3979);
xor U4173 (N_4173,N_3595,N_3378);
and U4174 (N_4174,N_3811,N_3472);
xor U4175 (N_4175,N_3133,N_3169);
and U4176 (N_4176,N_3724,N_3037);
nand U4177 (N_4177,N_3557,N_3091);
and U4178 (N_4178,N_3792,N_3849);
nor U4179 (N_4179,N_3582,N_3616);
nor U4180 (N_4180,N_3197,N_3150);
nand U4181 (N_4181,N_3551,N_3496);
nor U4182 (N_4182,N_3994,N_3690);
nand U4183 (N_4183,N_3319,N_3423);
and U4184 (N_4184,N_3131,N_3181);
xnor U4185 (N_4185,N_3474,N_3327);
xnor U4186 (N_4186,N_3331,N_3925);
nand U4187 (N_4187,N_3760,N_3232);
nand U4188 (N_4188,N_3160,N_3547);
nand U4189 (N_4189,N_3565,N_3038);
nand U4190 (N_4190,N_3625,N_3946);
or U4191 (N_4191,N_3844,N_3520);
nand U4192 (N_4192,N_3601,N_3112);
or U4193 (N_4193,N_3947,N_3602);
xor U4194 (N_4194,N_3710,N_3867);
nor U4195 (N_4195,N_3939,N_3068);
and U4196 (N_4196,N_3217,N_3648);
or U4197 (N_4197,N_3158,N_3671);
or U4198 (N_4198,N_3883,N_3934);
xor U4199 (N_4199,N_3222,N_3201);
and U4200 (N_4200,N_3456,N_3432);
xnor U4201 (N_4201,N_3830,N_3810);
nand U4202 (N_4202,N_3437,N_3570);
xor U4203 (N_4203,N_3092,N_3250);
or U4204 (N_4204,N_3479,N_3803);
xor U4205 (N_4205,N_3364,N_3819);
xnor U4206 (N_4206,N_3739,N_3823);
xor U4207 (N_4207,N_3384,N_3329);
nand U4208 (N_4208,N_3758,N_3603);
xnor U4209 (N_4209,N_3923,N_3088);
nand U4210 (N_4210,N_3833,N_3065);
and U4211 (N_4211,N_3967,N_3478);
and U4212 (N_4212,N_3362,N_3498);
nand U4213 (N_4213,N_3372,N_3080);
or U4214 (N_4214,N_3646,N_3057);
xor U4215 (N_4215,N_3737,N_3082);
nand U4216 (N_4216,N_3842,N_3628);
xnor U4217 (N_4217,N_3748,N_3780);
nor U4218 (N_4218,N_3694,N_3125);
nand U4219 (N_4219,N_3592,N_3140);
nand U4220 (N_4220,N_3063,N_3214);
nor U4221 (N_4221,N_3950,N_3564);
and U4222 (N_4222,N_3366,N_3046);
nand U4223 (N_4223,N_3255,N_3055);
xnor U4224 (N_4224,N_3200,N_3104);
nor U4225 (N_4225,N_3527,N_3696);
nand U4226 (N_4226,N_3905,N_3294);
and U4227 (N_4227,N_3952,N_3530);
xor U4228 (N_4228,N_3990,N_3535);
and U4229 (N_4229,N_3864,N_3053);
nor U4230 (N_4230,N_3930,N_3017);
and U4231 (N_4231,N_3415,N_3157);
nand U4232 (N_4232,N_3774,N_3202);
or U4233 (N_4233,N_3493,N_3666);
and U4234 (N_4234,N_3282,N_3230);
or U4235 (N_4235,N_3718,N_3376);
nor U4236 (N_4236,N_3342,N_3099);
or U4237 (N_4237,N_3051,N_3738);
nand U4238 (N_4238,N_3480,N_3486);
nor U4239 (N_4239,N_3069,N_3228);
xnor U4240 (N_4240,N_3205,N_3882);
and U4241 (N_4241,N_3873,N_3510);
xor U4242 (N_4242,N_3791,N_3964);
xnor U4243 (N_4243,N_3031,N_3931);
or U4244 (N_4244,N_3509,N_3240);
xor U4245 (N_4245,N_3135,N_3348);
and U4246 (N_4246,N_3621,N_3600);
nand U4247 (N_4247,N_3501,N_3041);
and U4248 (N_4248,N_3300,N_3237);
xnor U4249 (N_4249,N_3534,N_3448);
nor U4250 (N_4250,N_3768,N_3276);
and U4251 (N_4251,N_3295,N_3574);
nand U4252 (N_4252,N_3492,N_3180);
and U4253 (N_4253,N_3380,N_3587);
or U4254 (N_4254,N_3787,N_3885);
xor U4255 (N_4255,N_3094,N_3859);
or U4256 (N_4256,N_3682,N_3650);
and U4257 (N_4257,N_3397,N_3330);
or U4258 (N_4258,N_3940,N_3281);
or U4259 (N_4259,N_3033,N_3633);
or U4260 (N_4260,N_3916,N_3770);
nand U4261 (N_4261,N_3059,N_3050);
nor U4262 (N_4262,N_3172,N_3517);
nand U4263 (N_4263,N_3439,N_3252);
nor U4264 (N_4264,N_3424,N_3170);
or U4265 (N_4265,N_3750,N_3764);
or U4266 (N_4266,N_3171,N_3132);
nand U4267 (N_4267,N_3264,N_3001);
and U4268 (N_4268,N_3195,N_3734);
xor U4269 (N_4269,N_3425,N_3775);
nand U4270 (N_4270,N_3430,N_3853);
or U4271 (N_4271,N_3196,N_3745);
nor U4272 (N_4272,N_3433,N_3837);
nor U4273 (N_4273,N_3754,N_3070);
nand U4274 (N_4274,N_3609,N_3691);
or U4275 (N_4275,N_3089,N_3536);
nand U4276 (N_4276,N_3109,N_3291);
nand U4277 (N_4277,N_3614,N_3989);
xnor U4278 (N_4278,N_3575,N_3594);
nor U4279 (N_4279,N_3880,N_3213);
and U4280 (N_4280,N_3062,N_3900);
nand U4281 (N_4281,N_3142,N_3279);
nor U4282 (N_4282,N_3207,N_3079);
nand U4283 (N_4283,N_3354,N_3908);
nor U4284 (N_4284,N_3951,N_3917);
xnor U4285 (N_4285,N_3514,N_3151);
nand U4286 (N_4286,N_3010,N_3834);
xor U4287 (N_4287,N_3320,N_3268);
xor U4288 (N_4288,N_3178,N_3258);
and U4289 (N_4289,N_3980,N_3732);
xor U4290 (N_4290,N_3683,N_3454);
nand U4291 (N_4291,N_3503,N_3000);
xnor U4292 (N_4292,N_3452,N_3596);
or U4293 (N_4293,N_3386,N_3487);
and U4294 (N_4294,N_3871,N_3273);
and U4295 (N_4295,N_3845,N_3814);
and U4296 (N_4296,N_3555,N_3657);
nor U4297 (N_4297,N_3612,N_3490);
and U4298 (N_4298,N_3280,N_3123);
xor U4299 (N_4299,N_3508,N_3956);
xor U4300 (N_4300,N_3617,N_3226);
and U4301 (N_4301,N_3879,N_3084);
nor U4302 (N_4302,N_3395,N_3786);
xnor U4303 (N_4303,N_3179,N_3141);
and U4304 (N_4304,N_3513,N_3034);
nor U4305 (N_4305,N_3345,N_3253);
nor U4306 (N_4306,N_3743,N_3540);
or U4307 (N_4307,N_3414,N_3286);
nand U4308 (N_4308,N_3665,N_3681);
and U4309 (N_4309,N_3887,N_3411);
nor U4310 (N_4310,N_3346,N_3177);
or U4311 (N_4311,N_3168,N_3795);
or U4312 (N_4312,N_3488,N_3387);
nand U4313 (N_4313,N_3308,N_3011);
nand U4314 (N_4314,N_3674,N_3685);
nor U4315 (N_4315,N_3477,N_3139);
xor U4316 (N_4316,N_3963,N_3889);
or U4317 (N_4317,N_3126,N_3310);
nand U4318 (N_4318,N_3408,N_3115);
nor U4319 (N_4319,N_3550,N_3049);
or U4320 (N_4320,N_3426,N_3906);
nor U4321 (N_4321,N_3416,N_3056);
or U4322 (N_4322,N_3569,N_3373);
nor U4323 (N_4323,N_3450,N_3715);
or U4324 (N_4324,N_3225,N_3607);
or U4325 (N_4325,N_3166,N_3506);
and U4326 (N_4326,N_3462,N_3610);
xor U4327 (N_4327,N_3326,N_3164);
nor U4328 (N_4328,N_3705,N_3576);
nand U4329 (N_4329,N_3518,N_3266);
and U4330 (N_4330,N_3184,N_3447);
nor U4331 (N_4331,N_3689,N_3434);
xor U4332 (N_4332,N_3413,N_3021);
or U4333 (N_4333,N_3986,N_3578);
or U4334 (N_4334,N_3263,N_3105);
or U4335 (N_4335,N_3438,N_3678);
or U4336 (N_4336,N_3567,N_3406);
xor U4337 (N_4337,N_3075,N_3703);
or U4338 (N_4338,N_3446,N_3812);
or U4339 (N_4339,N_3287,N_3585);
and U4340 (N_4340,N_3651,N_3847);
nand U4341 (N_4341,N_3840,N_3886);
or U4342 (N_4342,N_3929,N_3955);
or U4343 (N_4343,N_3204,N_3862);
and U4344 (N_4344,N_3756,N_3189);
and U4345 (N_4345,N_3144,N_3767);
nand U4346 (N_4346,N_3970,N_3241);
and U4347 (N_4347,N_3820,N_3577);
nand U4348 (N_4348,N_3539,N_3025);
nor U4349 (N_4349,N_3566,N_3832);
nand U4350 (N_4350,N_3554,N_3156);
nand U4351 (N_4351,N_3325,N_3039);
and U4352 (N_4352,N_3957,N_3081);
xnor U4353 (N_4353,N_3679,N_3290);
xnor U4354 (N_4354,N_3846,N_3259);
xnor U4355 (N_4355,N_3524,N_3552);
nand U4356 (N_4356,N_3913,N_3851);
or U4357 (N_4357,N_3265,N_3730);
and U4358 (N_4358,N_3973,N_3073);
or U4359 (N_4359,N_3246,N_3042);
nand U4360 (N_4360,N_3457,N_3639);
nand U4361 (N_4361,N_3113,N_3317);
and U4362 (N_4362,N_3652,N_3662);
or U4363 (N_4363,N_3953,N_3711);
xnor U4364 (N_4364,N_3322,N_3153);
nor U4365 (N_4365,N_3838,N_3945);
or U4366 (N_4366,N_3007,N_3192);
xnor U4367 (N_4367,N_3735,N_3466);
xor U4368 (N_4368,N_3242,N_3731);
or U4369 (N_4369,N_3015,N_3626);
and U4370 (N_4370,N_3751,N_3938);
or U4371 (N_4371,N_3110,N_3667);
or U4372 (N_4372,N_3429,N_3728);
and U4373 (N_4373,N_3504,N_3402);
nor U4374 (N_4374,N_3965,N_3012);
nand U4375 (N_4375,N_3966,N_3350);
nand U4376 (N_4376,N_3637,N_3919);
nor U4377 (N_4377,N_3772,N_3874);
nand U4378 (N_4378,N_3401,N_3483);
xnor U4379 (N_4379,N_3634,N_3147);
and U4380 (N_4380,N_3784,N_3790);
nor U4381 (N_4381,N_3725,N_3145);
xor U4382 (N_4382,N_3561,N_3289);
or U4383 (N_4383,N_3618,N_3227);
nand U4384 (N_4384,N_3759,N_3360);
xnor U4385 (N_4385,N_3163,N_3453);
nor U4386 (N_4386,N_3316,N_3644);
nand U4387 (N_4387,N_3542,N_3606);
nand U4388 (N_4388,N_3249,N_3948);
nand U4389 (N_4389,N_3299,N_3529);
xor U4390 (N_4390,N_3729,N_3712);
xnor U4391 (N_4391,N_3976,N_3405);
and U4392 (N_4392,N_3394,N_3995);
or U4393 (N_4393,N_3604,N_3984);
xor U4394 (N_4394,N_3336,N_3799);
xor U4395 (N_4395,N_3491,N_3615);
nand U4396 (N_4396,N_3872,N_3622);
nand U4397 (N_4397,N_3543,N_3698);
or U4398 (N_4398,N_3390,N_3920);
nor U4399 (N_4399,N_3060,N_3755);
and U4400 (N_4400,N_3206,N_3076);
and U4401 (N_4401,N_3876,N_3303);
or U4402 (N_4402,N_3248,N_3341);
and U4403 (N_4403,N_3918,N_3719);
or U4404 (N_4404,N_3713,N_3869);
or U4405 (N_4405,N_3997,N_3302);
nor U4406 (N_4406,N_3635,N_3645);
xnor U4407 (N_4407,N_3194,N_3417);
or U4408 (N_4408,N_3288,N_3661);
xnor U4409 (N_4409,N_3597,N_3183);
xnor U4410 (N_4410,N_3367,N_3465);
nand U4411 (N_4411,N_3898,N_3136);
xor U4412 (N_4412,N_3216,N_3269);
and U4413 (N_4413,N_3475,N_3312);
nand U4414 (N_4414,N_3525,N_3121);
and U4415 (N_4415,N_3188,N_3461);
xor U4416 (N_4416,N_3638,N_3267);
xnor U4417 (N_4417,N_3469,N_3752);
xor U4418 (N_4418,N_3020,N_3935);
and U4419 (N_4419,N_3523,N_3003);
nand U4420 (N_4420,N_3388,N_3541);
nand U4421 (N_4421,N_3744,N_3583);
and U4422 (N_4422,N_3072,N_3422);
nor U4423 (N_4423,N_3672,N_3165);
or U4424 (N_4424,N_3762,N_3825);
nor U4425 (N_4425,N_3357,N_3256);
nor U4426 (N_4426,N_3982,N_3794);
xnor U4427 (N_4427,N_3511,N_3815);
nand U4428 (N_4428,N_3086,N_3107);
nor U4429 (N_4429,N_3199,N_3902);
nor U4430 (N_4430,N_3191,N_3993);
xor U4431 (N_4431,N_3428,N_3064);
or U4432 (N_4432,N_3521,N_3285);
nor U4433 (N_4433,N_3298,N_3875);
or U4434 (N_4434,N_3014,N_3972);
xor U4435 (N_4435,N_3473,N_3848);
nor U4436 (N_4436,N_3664,N_3353);
xor U4437 (N_4437,N_3358,N_3315);
nor U4438 (N_4438,N_3347,N_3516);
nor U4439 (N_4439,N_3502,N_3559);
and U4440 (N_4440,N_3494,N_3118);
xnor U4441 (N_4441,N_3047,N_3974);
nor U4442 (N_4442,N_3827,N_3911);
xor U4443 (N_4443,N_3404,N_3598);
nor U4444 (N_4444,N_3673,N_3093);
nor U4445 (N_4445,N_3969,N_3403);
xor U4446 (N_4446,N_3443,N_3318);
and U4447 (N_4447,N_3470,N_3221);
or U4448 (N_4448,N_3822,N_3138);
nor U4449 (N_4449,N_3881,N_3835);
and U4450 (N_4450,N_3382,N_3828);
nand U4451 (N_4451,N_3736,N_3996);
xnor U4452 (N_4452,N_3261,N_3369);
and U4453 (N_4453,N_3324,N_3949);
nand U4454 (N_4454,N_3375,N_3449);
nor U4455 (N_4455,N_3605,N_3236);
or U4456 (N_4456,N_3371,N_3219);
nand U4457 (N_4457,N_3971,N_3463);
or U4458 (N_4458,N_3926,N_3418);
nor U4459 (N_4459,N_3043,N_3363);
and U4460 (N_4460,N_3693,N_3927);
xnor U4461 (N_4461,N_3680,N_3130);
nand U4462 (N_4462,N_3349,N_3507);
and U4463 (N_4463,N_3155,N_3251);
or U4464 (N_4464,N_3852,N_3239);
xor U4465 (N_4465,N_3723,N_3546);
or U4466 (N_4466,N_3484,N_3991);
nand U4467 (N_4467,N_3208,N_3865);
nand U4468 (N_4468,N_3757,N_3223);
nor U4469 (N_4469,N_3747,N_3695);
nand U4470 (N_4470,N_3581,N_3699);
or U4471 (N_4471,N_3392,N_3306);
and U4472 (N_4472,N_3396,N_3895);
nor U4473 (N_4473,N_3410,N_3899);
or U4474 (N_4474,N_3742,N_3257);
xor U4475 (N_4475,N_3203,N_3005);
nor U4476 (N_4476,N_3858,N_3720);
or U4477 (N_4477,N_3398,N_3028);
nor U4478 (N_4478,N_3924,N_3500);
and U4479 (N_4479,N_3655,N_3451);
xor U4480 (N_4480,N_3173,N_3861);
nand U4481 (N_4481,N_3262,N_3238);
or U4482 (N_4482,N_3365,N_3733);
or U4483 (N_4483,N_3440,N_3468);
and U4484 (N_4484,N_3999,N_3077);
nand U4485 (N_4485,N_3936,N_3692);
xnor U4486 (N_4486,N_3571,N_3343);
nor U4487 (N_4487,N_3697,N_3016);
nand U4488 (N_4488,N_3087,N_3114);
xor U4489 (N_4489,N_3231,N_3640);
nor U4490 (N_4490,N_3159,N_3435);
nor U4491 (N_4491,N_3254,N_3962);
nand U4492 (N_4492,N_3857,N_3647);
xnor U4493 (N_4493,N_3022,N_3505);
or U4494 (N_4494,N_3688,N_3670);
nor U4495 (N_4495,N_3708,N_3702);
xor U4496 (N_4496,N_3941,N_3816);
xnor U4497 (N_4497,N_3067,N_3441);
and U4498 (N_4498,N_3549,N_3537);
xor U4499 (N_4499,N_3998,N_3210);
or U4500 (N_4500,N_3492,N_3755);
or U4501 (N_4501,N_3271,N_3793);
nand U4502 (N_4502,N_3721,N_3784);
nand U4503 (N_4503,N_3134,N_3817);
xnor U4504 (N_4504,N_3880,N_3692);
nor U4505 (N_4505,N_3565,N_3478);
and U4506 (N_4506,N_3200,N_3792);
xor U4507 (N_4507,N_3400,N_3503);
xnor U4508 (N_4508,N_3957,N_3572);
and U4509 (N_4509,N_3104,N_3440);
or U4510 (N_4510,N_3478,N_3708);
xnor U4511 (N_4511,N_3427,N_3202);
nand U4512 (N_4512,N_3901,N_3538);
nand U4513 (N_4513,N_3088,N_3632);
nor U4514 (N_4514,N_3447,N_3921);
nand U4515 (N_4515,N_3709,N_3036);
and U4516 (N_4516,N_3630,N_3441);
xor U4517 (N_4517,N_3955,N_3648);
nand U4518 (N_4518,N_3526,N_3846);
nor U4519 (N_4519,N_3439,N_3951);
nand U4520 (N_4520,N_3860,N_3916);
nand U4521 (N_4521,N_3039,N_3341);
nand U4522 (N_4522,N_3209,N_3824);
nor U4523 (N_4523,N_3512,N_3777);
or U4524 (N_4524,N_3211,N_3765);
or U4525 (N_4525,N_3941,N_3445);
nand U4526 (N_4526,N_3202,N_3037);
and U4527 (N_4527,N_3607,N_3397);
nor U4528 (N_4528,N_3287,N_3303);
nor U4529 (N_4529,N_3182,N_3206);
nand U4530 (N_4530,N_3522,N_3303);
nor U4531 (N_4531,N_3841,N_3484);
and U4532 (N_4532,N_3732,N_3681);
or U4533 (N_4533,N_3868,N_3468);
nor U4534 (N_4534,N_3974,N_3041);
nor U4535 (N_4535,N_3904,N_3178);
nor U4536 (N_4536,N_3240,N_3366);
and U4537 (N_4537,N_3205,N_3298);
or U4538 (N_4538,N_3329,N_3681);
and U4539 (N_4539,N_3430,N_3595);
or U4540 (N_4540,N_3529,N_3245);
xor U4541 (N_4541,N_3238,N_3782);
xor U4542 (N_4542,N_3141,N_3684);
xnor U4543 (N_4543,N_3461,N_3557);
xor U4544 (N_4544,N_3189,N_3753);
and U4545 (N_4545,N_3824,N_3691);
nand U4546 (N_4546,N_3730,N_3678);
and U4547 (N_4547,N_3384,N_3078);
and U4548 (N_4548,N_3004,N_3183);
nand U4549 (N_4549,N_3294,N_3600);
xor U4550 (N_4550,N_3798,N_3261);
xor U4551 (N_4551,N_3343,N_3611);
nor U4552 (N_4552,N_3054,N_3571);
or U4553 (N_4553,N_3903,N_3977);
nor U4554 (N_4554,N_3620,N_3716);
or U4555 (N_4555,N_3753,N_3122);
and U4556 (N_4556,N_3960,N_3255);
or U4557 (N_4557,N_3890,N_3184);
xnor U4558 (N_4558,N_3807,N_3599);
or U4559 (N_4559,N_3211,N_3337);
nor U4560 (N_4560,N_3925,N_3986);
and U4561 (N_4561,N_3390,N_3348);
nand U4562 (N_4562,N_3138,N_3698);
or U4563 (N_4563,N_3854,N_3594);
xnor U4564 (N_4564,N_3199,N_3728);
or U4565 (N_4565,N_3923,N_3180);
and U4566 (N_4566,N_3859,N_3463);
and U4567 (N_4567,N_3660,N_3739);
and U4568 (N_4568,N_3467,N_3365);
and U4569 (N_4569,N_3077,N_3527);
or U4570 (N_4570,N_3110,N_3012);
nor U4571 (N_4571,N_3324,N_3106);
nor U4572 (N_4572,N_3816,N_3576);
nand U4573 (N_4573,N_3608,N_3617);
xnor U4574 (N_4574,N_3324,N_3904);
nor U4575 (N_4575,N_3992,N_3293);
and U4576 (N_4576,N_3373,N_3097);
nand U4577 (N_4577,N_3282,N_3361);
nor U4578 (N_4578,N_3765,N_3417);
nor U4579 (N_4579,N_3923,N_3400);
nand U4580 (N_4580,N_3083,N_3347);
and U4581 (N_4581,N_3898,N_3818);
nand U4582 (N_4582,N_3936,N_3625);
nor U4583 (N_4583,N_3164,N_3401);
xnor U4584 (N_4584,N_3921,N_3504);
nand U4585 (N_4585,N_3332,N_3916);
xor U4586 (N_4586,N_3700,N_3652);
and U4587 (N_4587,N_3744,N_3577);
nand U4588 (N_4588,N_3996,N_3227);
xnor U4589 (N_4589,N_3672,N_3704);
xor U4590 (N_4590,N_3491,N_3876);
or U4591 (N_4591,N_3554,N_3545);
xor U4592 (N_4592,N_3063,N_3352);
nand U4593 (N_4593,N_3580,N_3680);
nand U4594 (N_4594,N_3703,N_3275);
and U4595 (N_4595,N_3018,N_3946);
xnor U4596 (N_4596,N_3599,N_3565);
and U4597 (N_4597,N_3459,N_3921);
nor U4598 (N_4598,N_3731,N_3817);
nor U4599 (N_4599,N_3953,N_3887);
nand U4600 (N_4600,N_3550,N_3446);
nor U4601 (N_4601,N_3772,N_3136);
xnor U4602 (N_4602,N_3924,N_3147);
nor U4603 (N_4603,N_3655,N_3636);
xnor U4604 (N_4604,N_3010,N_3557);
and U4605 (N_4605,N_3186,N_3027);
xnor U4606 (N_4606,N_3855,N_3956);
and U4607 (N_4607,N_3159,N_3024);
and U4608 (N_4608,N_3490,N_3799);
and U4609 (N_4609,N_3532,N_3542);
nand U4610 (N_4610,N_3656,N_3291);
xnor U4611 (N_4611,N_3424,N_3665);
or U4612 (N_4612,N_3161,N_3014);
xnor U4613 (N_4613,N_3830,N_3015);
nor U4614 (N_4614,N_3507,N_3592);
or U4615 (N_4615,N_3363,N_3293);
xor U4616 (N_4616,N_3121,N_3117);
nand U4617 (N_4617,N_3616,N_3400);
or U4618 (N_4618,N_3536,N_3739);
or U4619 (N_4619,N_3699,N_3509);
nand U4620 (N_4620,N_3460,N_3491);
nand U4621 (N_4621,N_3289,N_3933);
nand U4622 (N_4622,N_3391,N_3485);
or U4623 (N_4623,N_3717,N_3093);
xnor U4624 (N_4624,N_3335,N_3710);
and U4625 (N_4625,N_3545,N_3827);
or U4626 (N_4626,N_3710,N_3080);
nor U4627 (N_4627,N_3915,N_3956);
or U4628 (N_4628,N_3798,N_3538);
and U4629 (N_4629,N_3890,N_3467);
xnor U4630 (N_4630,N_3515,N_3847);
and U4631 (N_4631,N_3254,N_3838);
nor U4632 (N_4632,N_3617,N_3839);
and U4633 (N_4633,N_3229,N_3250);
nor U4634 (N_4634,N_3876,N_3920);
xnor U4635 (N_4635,N_3463,N_3401);
nand U4636 (N_4636,N_3849,N_3067);
or U4637 (N_4637,N_3883,N_3623);
and U4638 (N_4638,N_3629,N_3365);
or U4639 (N_4639,N_3896,N_3591);
xnor U4640 (N_4640,N_3022,N_3288);
or U4641 (N_4641,N_3262,N_3313);
nand U4642 (N_4642,N_3504,N_3960);
and U4643 (N_4643,N_3278,N_3396);
nand U4644 (N_4644,N_3203,N_3263);
and U4645 (N_4645,N_3715,N_3593);
nand U4646 (N_4646,N_3603,N_3466);
nor U4647 (N_4647,N_3845,N_3678);
nor U4648 (N_4648,N_3035,N_3357);
nor U4649 (N_4649,N_3603,N_3923);
and U4650 (N_4650,N_3321,N_3331);
nand U4651 (N_4651,N_3276,N_3924);
nor U4652 (N_4652,N_3389,N_3726);
xor U4653 (N_4653,N_3482,N_3340);
or U4654 (N_4654,N_3773,N_3462);
and U4655 (N_4655,N_3088,N_3915);
or U4656 (N_4656,N_3022,N_3867);
xnor U4657 (N_4657,N_3020,N_3543);
nor U4658 (N_4658,N_3944,N_3076);
and U4659 (N_4659,N_3812,N_3767);
or U4660 (N_4660,N_3121,N_3120);
xor U4661 (N_4661,N_3776,N_3210);
nand U4662 (N_4662,N_3830,N_3791);
or U4663 (N_4663,N_3709,N_3082);
nand U4664 (N_4664,N_3757,N_3852);
or U4665 (N_4665,N_3934,N_3987);
nor U4666 (N_4666,N_3002,N_3384);
nor U4667 (N_4667,N_3107,N_3895);
nor U4668 (N_4668,N_3864,N_3791);
and U4669 (N_4669,N_3489,N_3793);
nand U4670 (N_4670,N_3126,N_3175);
or U4671 (N_4671,N_3421,N_3090);
nand U4672 (N_4672,N_3423,N_3733);
and U4673 (N_4673,N_3836,N_3941);
nor U4674 (N_4674,N_3416,N_3535);
nand U4675 (N_4675,N_3951,N_3934);
nor U4676 (N_4676,N_3929,N_3848);
xor U4677 (N_4677,N_3296,N_3350);
nand U4678 (N_4678,N_3469,N_3536);
xor U4679 (N_4679,N_3865,N_3801);
xor U4680 (N_4680,N_3060,N_3562);
nand U4681 (N_4681,N_3858,N_3871);
or U4682 (N_4682,N_3739,N_3305);
xnor U4683 (N_4683,N_3408,N_3791);
or U4684 (N_4684,N_3914,N_3561);
nor U4685 (N_4685,N_3547,N_3996);
and U4686 (N_4686,N_3209,N_3756);
and U4687 (N_4687,N_3726,N_3516);
nand U4688 (N_4688,N_3226,N_3077);
xnor U4689 (N_4689,N_3506,N_3396);
nor U4690 (N_4690,N_3984,N_3620);
or U4691 (N_4691,N_3367,N_3729);
and U4692 (N_4692,N_3004,N_3363);
xnor U4693 (N_4693,N_3274,N_3203);
nand U4694 (N_4694,N_3268,N_3854);
or U4695 (N_4695,N_3489,N_3756);
nand U4696 (N_4696,N_3723,N_3636);
or U4697 (N_4697,N_3757,N_3038);
nand U4698 (N_4698,N_3575,N_3128);
xnor U4699 (N_4699,N_3681,N_3730);
and U4700 (N_4700,N_3871,N_3006);
xor U4701 (N_4701,N_3306,N_3053);
or U4702 (N_4702,N_3350,N_3072);
nand U4703 (N_4703,N_3746,N_3630);
nand U4704 (N_4704,N_3063,N_3176);
nand U4705 (N_4705,N_3250,N_3028);
nand U4706 (N_4706,N_3928,N_3476);
or U4707 (N_4707,N_3934,N_3002);
and U4708 (N_4708,N_3698,N_3257);
nor U4709 (N_4709,N_3518,N_3405);
nand U4710 (N_4710,N_3077,N_3526);
and U4711 (N_4711,N_3856,N_3780);
and U4712 (N_4712,N_3467,N_3764);
nor U4713 (N_4713,N_3854,N_3428);
and U4714 (N_4714,N_3621,N_3186);
xor U4715 (N_4715,N_3787,N_3959);
nand U4716 (N_4716,N_3609,N_3288);
xor U4717 (N_4717,N_3259,N_3121);
nand U4718 (N_4718,N_3554,N_3322);
xnor U4719 (N_4719,N_3066,N_3214);
nand U4720 (N_4720,N_3631,N_3781);
and U4721 (N_4721,N_3215,N_3795);
nor U4722 (N_4722,N_3330,N_3780);
and U4723 (N_4723,N_3932,N_3179);
or U4724 (N_4724,N_3287,N_3449);
nand U4725 (N_4725,N_3496,N_3047);
xor U4726 (N_4726,N_3770,N_3744);
nor U4727 (N_4727,N_3415,N_3595);
nor U4728 (N_4728,N_3766,N_3668);
xor U4729 (N_4729,N_3356,N_3650);
and U4730 (N_4730,N_3937,N_3812);
nand U4731 (N_4731,N_3164,N_3315);
xor U4732 (N_4732,N_3263,N_3424);
nand U4733 (N_4733,N_3881,N_3312);
nor U4734 (N_4734,N_3751,N_3490);
or U4735 (N_4735,N_3907,N_3607);
nand U4736 (N_4736,N_3918,N_3442);
xor U4737 (N_4737,N_3256,N_3117);
or U4738 (N_4738,N_3110,N_3225);
or U4739 (N_4739,N_3004,N_3563);
and U4740 (N_4740,N_3623,N_3829);
nor U4741 (N_4741,N_3307,N_3352);
xnor U4742 (N_4742,N_3515,N_3375);
nor U4743 (N_4743,N_3676,N_3189);
or U4744 (N_4744,N_3468,N_3476);
or U4745 (N_4745,N_3826,N_3562);
or U4746 (N_4746,N_3573,N_3840);
or U4747 (N_4747,N_3446,N_3825);
xnor U4748 (N_4748,N_3844,N_3029);
and U4749 (N_4749,N_3017,N_3387);
or U4750 (N_4750,N_3764,N_3905);
xor U4751 (N_4751,N_3842,N_3121);
and U4752 (N_4752,N_3146,N_3199);
xnor U4753 (N_4753,N_3144,N_3492);
nor U4754 (N_4754,N_3520,N_3976);
and U4755 (N_4755,N_3962,N_3526);
nand U4756 (N_4756,N_3605,N_3063);
nor U4757 (N_4757,N_3062,N_3040);
nor U4758 (N_4758,N_3771,N_3178);
or U4759 (N_4759,N_3332,N_3492);
nand U4760 (N_4760,N_3204,N_3486);
xor U4761 (N_4761,N_3841,N_3964);
xnor U4762 (N_4762,N_3331,N_3123);
nand U4763 (N_4763,N_3287,N_3357);
nor U4764 (N_4764,N_3060,N_3093);
and U4765 (N_4765,N_3254,N_3762);
or U4766 (N_4766,N_3220,N_3077);
nand U4767 (N_4767,N_3451,N_3633);
and U4768 (N_4768,N_3648,N_3318);
nor U4769 (N_4769,N_3187,N_3903);
and U4770 (N_4770,N_3634,N_3918);
nand U4771 (N_4771,N_3663,N_3850);
nand U4772 (N_4772,N_3039,N_3296);
nand U4773 (N_4773,N_3799,N_3377);
or U4774 (N_4774,N_3453,N_3527);
or U4775 (N_4775,N_3370,N_3757);
xnor U4776 (N_4776,N_3068,N_3153);
and U4777 (N_4777,N_3547,N_3856);
nor U4778 (N_4778,N_3933,N_3086);
nand U4779 (N_4779,N_3630,N_3790);
or U4780 (N_4780,N_3366,N_3165);
or U4781 (N_4781,N_3038,N_3818);
xnor U4782 (N_4782,N_3221,N_3808);
nand U4783 (N_4783,N_3180,N_3838);
and U4784 (N_4784,N_3151,N_3932);
xor U4785 (N_4785,N_3291,N_3653);
nand U4786 (N_4786,N_3643,N_3642);
and U4787 (N_4787,N_3743,N_3296);
or U4788 (N_4788,N_3308,N_3692);
or U4789 (N_4789,N_3371,N_3268);
and U4790 (N_4790,N_3145,N_3455);
nor U4791 (N_4791,N_3932,N_3021);
nand U4792 (N_4792,N_3657,N_3797);
or U4793 (N_4793,N_3017,N_3127);
nand U4794 (N_4794,N_3866,N_3561);
xnor U4795 (N_4795,N_3219,N_3870);
and U4796 (N_4796,N_3385,N_3671);
nor U4797 (N_4797,N_3151,N_3203);
nor U4798 (N_4798,N_3211,N_3979);
xor U4799 (N_4799,N_3553,N_3777);
or U4800 (N_4800,N_3444,N_3750);
xor U4801 (N_4801,N_3312,N_3393);
xor U4802 (N_4802,N_3844,N_3815);
nand U4803 (N_4803,N_3200,N_3666);
nand U4804 (N_4804,N_3495,N_3869);
nor U4805 (N_4805,N_3069,N_3428);
nor U4806 (N_4806,N_3073,N_3944);
xor U4807 (N_4807,N_3579,N_3205);
nor U4808 (N_4808,N_3217,N_3668);
or U4809 (N_4809,N_3233,N_3864);
xor U4810 (N_4810,N_3427,N_3109);
nand U4811 (N_4811,N_3921,N_3924);
nor U4812 (N_4812,N_3562,N_3571);
or U4813 (N_4813,N_3924,N_3696);
or U4814 (N_4814,N_3917,N_3025);
or U4815 (N_4815,N_3213,N_3866);
nand U4816 (N_4816,N_3960,N_3618);
and U4817 (N_4817,N_3951,N_3043);
and U4818 (N_4818,N_3279,N_3845);
or U4819 (N_4819,N_3265,N_3981);
or U4820 (N_4820,N_3141,N_3694);
nand U4821 (N_4821,N_3778,N_3108);
nor U4822 (N_4822,N_3597,N_3760);
nand U4823 (N_4823,N_3629,N_3783);
nor U4824 (N_4824,N_3384,N_3623);
or U4825 (N_4825,N_3880,N_3678);
or U4826 (N_4826,N_3656,N_3198);
or U4827 (N_4827,N_3719,N_3619);
and U4828 (N_4828,N_3260,N_3953);
nand U4829 (N_4829,N_3825,N_3627);
nor U4830 (N_4830,N_3755,N_3959);
nor U4831 (N_4831,N_3643,N_3710);
and U4832 (N_4832,N_3787,N_3556);
xor U4833 (N_4833,N_3523,N_3721);
xor U4834 (N_4834,N_3926,N_3112);
xor U4835 (N_4835,N_3618,N_3946);
nor U4836 (N_4836,N_3929,N_3753);
nand U4837 (N_4837,N_3610,N_3116);
and U4838 (N_4838,N_3394,N_3908);
and U4839 (N_4839,N_3540,N_3848);
xor U4840 (N_4840,N_3806,N_3548);
or U4841 (N_4841,N_3040,N_3389);
xnor U4842 (N_4842,N_3248,N_3653);
xnor U4843 (N_4843,N_3917,N_3670);
or U4844 (N_4844,N_3289,N_3432);
or U4845 (N_4845,N_3730,N_3329);
xor U4846 (N_4846,N_3379,N_3847);
or U4847 (N_4847,N_3874,N_3050);
and U4848 (N_4848,N_3144,N_3358);
nand U4849 (N_4849,N_3970,N_3879);
and U4850 (N_4850,N_3337,N_3571);
or U4851 (N_4851,N_3806,N_3490);
nand U4852 (N_4852,N_3919,N_3162);
and U4853 (N_4853,N_3680,N_3707);
nand U4854 (N_4854,N_3501,N_3653);
nor U4855 (N_4855,N_3528,N_3766);
nor U4856 (N_4856,N_3463,N_3920);
xor U4857 (N_4857,N_3631,N_3390);
or U4858 (N_4858,N_3403,N_3177);
or U4859 (N_4859,N_3303,N_3029);
nor U4860 (N_4860,N_3282,N_3759);
or U4861 (N_4861,N_3166,N_3222);
or U4862 (N_4862,N_3205,N_3363);
and U4863 (N_4863,N_3975,N_3519);
xnor U4864 (N_4864,N_3500,N_3749);
or U4865 (N_4865,N_3191,N_3937);
nor U4866 (N_4866,N_3532,N_3956);
xor U4867 (N_4867,N_3705,N_3085);
and U4868 (N_4868,N_3712,N_3679);
nor U4869 (N_4869,N_3529,N_3835);
and U4870 (N_4870,N_3593,N_3527);
or U4871 (N_4871,N_3699,N_3803);
nand U4872 (N_4872,N_3221,N_3830);
xnor U4873 (N_4873,N_3320,N_3579);
or U4874 (N_4874,N_3037,N_3749);
xor U4875 (N_4875,N_3591,N_3290);
nand U4876 (N_4876,N_3117,N_3837);
or U4877 (N_4877,N_3140,N_3282);
xnor U4878 (N_4878,N_3377,N_3032);
nor U4879 (N_4879,N_3678,N_3394);
or U4880 (N_4880,N_3875,N_3612);
or U4881 (N_4881,N_3928,N_3805);
nor U4882 (N_4882,N_3109,N_3753);
and U4883 (N_4883,N_3582,N_3559);
or U4884 (N_4884,N_3915,N_3597);
nor U4885 (N_4885,N_3320,N_3141);
or U4886 (N_4886,N_3442,N_3250);
or U4887 (N_4887,N_3309,N_3766);
nor U4888 (N_4888,N_3046,N_3356);
or U4889 (N_4889,N_3401,N_3305);
or U4890 (N_4890,N_3874,N_3414);
nand U4891 (N_4891,N_3562,N_3808);
nor U4892 (N_4892,N_3533,N_3864);
nand U4893 (N_4893,N_3933,N_3784);
and U4894 (N_4894,N_3317,N_3782);
nor U4895 (N_4895,N_3882,N_3424);
and U4896 (N_4896,N_3861,N_3429);
nand U4897 (N_4897,N_3779,N_3461);
xnor U4898 (N_4898,N_3236,N_3434);
or U4899 (N_4899,N_3208,N_3122);
nand U4900 (N_4900,N_3240,N_3273);
xnor U4901 (N_4901,N_3560,N_3005);
nand U4902 (N_4902,N_3521,N_3842);
nand U4903 (N_4903,N_3470,N_3578);
nand U4904 (N_4904,N_3665,N_3988);
nor U4905 (N_4905,N_3884,N_3403);
or U4906 (N_4906,N_3865,N_3359);
nor U4907 (N_4907,N_3800,N_3688);
and U4908 (N_4908,N_3112,N_3966);
or U4909 (N_4909,N_3644,N_3822);
and U4910 (N_4910,N_3780,N_3153);
xor U4911 (N_4911,N_3499,N_3188);
nor U4912 (N_4912,N_3193,N_3803);
xnor U4913 (N_4913,N_3624,N_3671);
xor U4914 (N_4914,N_3778,N_3273);
nand U4915 (N_4915,N_3802,N_3114);
or U4916 (N_4916,N_3527,N_3974);
nand U4917 (N_4917,N_3038,N_3228);
and U4918 (N_4918,N_3015,N_3412);
nor U4919 (N_4919,N_3588,N_3277);
xnor U4920 (N_4920,N_3686,N_3016);
nand U4921 (N_4921,N_3870,N_3475);
xor U4922 (N_4922,N_3203,N_3146);
or U4923 (N_4923,N_3618,N_3184);
nor U4924 (N_4924,N_3308,N_3965);
nor U4925 (N_4925,N_3408,N_3844);
or U4926 (N_4926,N_3060,N_3044);
xnor U4927 (N_4927,N_3312,N_3916);
xor U4928 (N_4928,N_3283,N_3656);
or U4929 (N_4929,N_3833,N_3542);
nand U4930 (N_4930,N_3188,N_3290);
nand U4931 (N_4931,N_3474,N_3156);
or U4932 (N_4932,N_3530,N_3905);
nor U4933 (N_4933,N_3332,N_3369);
nor U4934 (N_4934,N_3993,N_3562);
and U4935 (N_4935,N_3383,N_3797);
nand U4936 (N_4936,N_3398,N_3007);
nor U4937 (N_4937,N_3726,N_3522);
or U4938 (N_4938,N_3432,N_3253);
nand U4939 (N_4939,N_3835,N_3507);
nor U4940 (N_4940,N_3562,N_3942);
or U4941 (N_4941,N_3397,N_3855);
xnor U4942 (N_4942,N_3090,N_3833);
nand U4943 (N_4943,N_3262,N_3234);
nand U4944 (N_4944,N_3279,N_3458);
nor U4945 (N_4945,N_3669,N_3120);
nor U4946 (N_4946,N_3157,N_3602);
nor U4947 (N_4947,N_3454,N_3112);
xor U4948 (N_4948,N_3919,N_3787);
nor U4949 (N_4949,N_3979,N_3545);
or U4950 (N_4950,N_3696,N_3224);
xor U4951 (N_4951,N_3882,N_3543);
and U4952 (N_4952,N_3841,N_3134);
nand U4953 (N_4953,N_3117,N_3323);
or U4954 (N_4954,N_3315,N_3097);
xor U4955 (N_4955,N_3028,N_3574);
nand U4956 (N_4956,N_3122,N_3942);
nor U4957 (N_4957,N_3277,N_3237);
nor U4958 (N_4958,N_3463,N_3339);
or U4959 (N_4959,N_3355,N_3448);
nor U4960 (N_4960,N_3023,N_3285);
nor U4961 (N_4961,N_3221,N_3736);
nor U4962 (N_4962,N_3543,N_3042);
nand U4963 (N_4963,N_3155,N_3950);
nor U4964 (N_4964,N_3572,N_3632);
and U4965 (N_4965,N_3949,N_3896);
xnor U4966 (N_4966,N_3330,N_3987);
or U4967 (N_4967,N_3329,N_3505);
nor U4968 (N_4968,N_3848,N_3361);
nor U4969 (N_4969,N_3343,N_3542);
and U4970 (N_4970,N_3076,N_3360);
nand U4971 (N_4971,N_3777,N_3419);
nand U4972 (N_4972,N_3826,N_3451);
nand U4973 (N_4973,N_3308,N_3148);
xor U4974 (N_4974,N_3405,N_3283);
nand U4975 (N_4975,N_3911,N_3691);
xnor U4976 (N_4976,N_3594,N_3622);
xnor U4977 (N_4977,N_3734,N_3955);
or U4978 (N_4978,N_3884,N_3454);
and U4979 (N_4979,N_3521,N_3400);
xor U4980 (N_4980,N_3590,N_3307);
and U4981 (N_4981,N_3115,N_3235);
or U4982 (N_4982,N_3672,N_3880);
nand U4983 (N_4983,N_3507,N_3172);
nor U4984 (N_4984,N_3769,N_3856);
xor U4985 (N_4985,N_3612,N_3286);
nor U4986 (N_4986,N_3889,N_3345);
nand U4987 (N_4987,N_3561,N_3226);
and U4988 (N_4988,N_3293,N_3785);
nor U4989 (N_4989,N_3992,N_3455);
and U4990 (N_4990,N_3372,N_3267);
xor U4991 (N_4991,N_3065,N_3381);
nand U4992 (N_4992,N_3849,N_3615);
nand U4993 (N_4993,N_3593,N_3281);
or U4994 (N_4994,N_3669,N_3219);
nand U4995 (N_4995,N_3265,N_3820);
xnor U4996 (N_4996,N_3979,N_3297);
nand U4997 (N_4997,N_3521,N_3710);
nor U4998 (N_4998,N_3425,N_3373);
nor U4999 (N_4999,N_3079,N_3138);
nor U5000 (N_5000,N_4039,N_4936);
nand U5001 (N_5001,N_4871,N_4033);
and U5002 (N_5002,N_4483,N_4295);
nor U5003 (N_5003,N_4398,N_4649);
nand U5004 (N_5004,N_4457,N_4328);
nand U5005 (N_5005,N_4989,N_4978);
or U5006 (N_5006,N_4016,N_4629);
nand U5007 (N_5007,N_4934,N_4996);
and U5008 (N_5008,N_4838,N_4660);
xnor U5009 (N_5009,N_4741,N_4954);
nor U5010 (N_5010,N_4140,N_4909);
or U5011 (N_5011,N_4368,N_4603);
nor U5012 (N_5012,N_4618,N_4687);
and U5013 (N_5013,N_4121,N_4260);
and U5014 (N_5014,N_4866,N_4758);
and U5015 (N_5015,N_4972,N_4529);
nor U5016 (N_5016,N_4523,N_4502);
or U5017 (N_5017,N_4290,N_4755);
nand U5018 (N_5018,N_4532,N_4263);
xnor U5019 (N_5019,N_4353,N_4462);
xor U5020 (N_5020,N_4329,N_4062);
and U5021 (N_5021,N_4230,N_4746);
and U5022 (N_5022,N_4504,N_4362);
xnor U5023 (N_5023,N_4339,N_4506);
or U5024 (N_5024,N_4992,N_4897);
and U5025 (N_5025,N_4732,N_4659);
nor U5026 (N_5026,N_4586,N_4748);
or U5027 (N_5027,N_4416,N_4813);
nand U5028 (N_5028,N_4227,N_4887);
nor U5029 (N_5029,N_4381,N_4772);
nor U5030 (N_5030,N_4695,N_4827);
xnor U5031 (N_5031,N_4665,N_4805);
or U5032 (N_5032,N_4968,N_4102);
or U5033 (N_5033,N_4366,N_4519);
and U5034 (N_5034,N_4025,N_4355);
nor U5035 (N_5035,N_4760,N_4669);
or U5036 (N_5036,N_4373,N_4509);
xnor U5037 (N_5037,N_4320,N_4393);
and U5038 (N_5038,N_4821,N_4343);
and U5039 (N_5039,N_4734,N_4106);
xnor U5040 (N_5040,N_4820,N_4786);
nor U5041 (N_5041,N_4508,N_4997);
xnor U5042 (N_5042,N_4704,N_4249);
nor U5043 (N_5043,N_4815,N_4971);
and U5044 (N_5044,N_4679,N_4847);
nand U5045 (N_5045,N_4083,N_4712);
or U5046 (N_5046,N_4736,N_4723);
and U5047 (N_5047,N_4044,N_4703);
nand U5048 (N_5048,N_4032,N_4892);
xnor U5049 (N_5049,N_4714,N_4662);
nor U5050 (N_5050,N_4967,N_4409);
or U5051 (N_5051,N_4585,N_4610);
xnor U5052 (N_5052,N_4010,N_4615);
nor U5053 (N_5053,N_4922,N_4981);
and U5054 (N_5054,N_4201,N_4883);
nor U5055 (N_5055,N_4194,N_4783);
nand U5056 (N_5056,N_4440,N_4534);
nand U5057 (N_5057,N_4291,N_4788);
xnor U5058 (N_5058,N_4135,N_4767);
xor U5059 (N_5059,N_4114,N_4361);
or U5060 (N_5060,N_4914,N_4469);
xnor U5061 (N_5061,N_4248,N_4013);
xnor U5062 (N_5062,N_4181,N_4627);
xnor U5063 (N_5063,N_4193,N_4654);
nor U5064 (N_5064,N_4609,N_4715);
xor U5065 (N_5065,N_4738,N_4300);
and U5066 (N_5066,N_4624,N_4728);
xor U5067 (N_5067,N_4397,N_4661);
xor U5068 (N_5068,N_4042,N_4153);
xor U5069 (N_5069,N_4500,N_4672);
nor U5070 (N_5070,N_4594,N_4238);
nor U5071 (N_5071,N_4103,N_4458);
nand U5072 (N_5072,N_4879,N_4943);
or U5073 (N_5073,N_4571,N_4730);
and U5074 (N_5074,N_4801,N_4563);
or U5075 (N_5075,N_4955,N_4432);
and U5076 (N_5076,N_4547,N_4242);
nor U5077 (N_5077,N_4031,N_4975);
nand U5078 (N_5078,N_4485,N_4727);
or U5079 (N_5079,N_4045,N_4894);
or U5080 (N_5080,N_4771,N_4845);
nor U5081 (N_5081,N_4780,N_4619);
or U5082 (N_5082,N_4697,N_4235);
nand U5083 (N_5083,N_4112,N_4258);
or U5084 (N_5084,N_4546,N_4766);
nand U5085 (N_5085,N_4400,N_4512);
and U5086 (N_5086,N_4575,N_4009);
and U5087 (N_5087,N_4977,N_4841);
xnor U5088 (N_5088,N_4239,N_4055);
nand U5089 (N_5089,N_4411,N_4204);
and U5090 (N_5090,N_4860,N_4918);
xnor U5091 (N_5091,N_4360,N_4030);
nand U5092 (N_5092,N_4162,N_4747);
nor U5093 (N_5093,N_4038,N_4941);
nor U5094 (N_5094,N_4979,N_4210);
nand U5095 (N_5095,N_4787,N_4069);
xor U5096 (N_5096,N_4692,N_4449);
xor U5097 (N_5097,N_4602,N_4014);
or U5098 (N_5098,N_4021,N_4399);
xor U5099 (N_5099,N_4154,N_4915);
nand U5100 (N_5100,N_4844,N_4306);
and U5101 (N_5101,N_4183,N_4250);
and U5102 (N_5102,N_4579,N_4643);
and U5103 (N_5103,N_4965,N_4710);
or U5104 (N_5104,N_4430,N_4898);
nand U5105 (N_5105,N_4177,N_4202);
and U5106 (N_5106,N_4445,N_4691);
or U5107 (N_5107,N_4241,N_4716);
and U5108 (N_5108,N_4027,N_4919);
nand U5109 (N_5109,N_4641,N_4208);
nor U5110 (N_5110,N_4735,N_4437);
or U5111 (N_5111,N_4739,N_4453);
nand U5112 (N_5112,N_4549,N_4520);
or U5113 (N_5113,N_4698,N_4463);
or U5114 (N_5114,N_4800,N_4369);
xor U5115 (N_5115,N_4903,N_4294);
and U5116 (N_5116,N_4998,N_4707);
xnor U5117 (N_5117,N_4589,N_4572);
or U5118 (N_5118,N_4964,N_4376);
and U5119 (N_5119,N_4427,N_4782);
nor U5120 (N_5120,N_4465,N_4839);
nand U5121 (N_5121,N_4671,N_4663);
and U5122 (N_5122,N_4528,N_4753);
xnor U5123 (N_5123,N_4060,N_4165);
nor U5124 (N_5124,N_4468,N_4335);
nand U5125 (N_5125,N_4612,N_4085);
and U5126 (N_5126,N_4757,N_4047);
and U5127 (N_5127,N_4680,N_4137);
xor U5128 (N_5128,N_4164,N_4702);
nor U5129 (N_5129,N_4058,N_4002);
xnor U5130 (N_5130,N_4582,N_4994);
nor U5131 (N_5131,N_4299,N_4858);
nor U5132 (N_5132,N_4912,N_4948);
nand U5133 (N_5133,N_4637,N_4598);
and U5134 (N_5134,N_4348,N_4455);
and U5135 (N_5135,N_4775,N_4550);
or U5136 (N_5136,N_4940,N_4065);
nor U5137 (N_5137,N_4507,N_4236);
xnor U5138 (N_5138,N_4479,N_4868);
and U5139 (N_5139,N_4725,N_4960);
nor U5140 (N_5140,N_4726,N_4650);
xnor U5141 (N_5141,N_4478,N_4608);
nor U5142 (N_5142,N_4802,N_4742);
nand U5143 (N_5143,N_4480,N_4623);
or U5144 (N_5144,N_4187,N_4804);
nand U5145 (N_5145,N_4498,N_4438);
nand U5146 (N_5146,N_4341,N_4855);
xnor U5147 (N_5147,N_4818,N_4597);
nor U5148 (N_5148,N_4810,N_4811);
and U5149 (N_5149,N_4491,N_4240);
nand U5150 (N_5150,N_4272,N_4213);
and U5151 (N_5151,N_4321,N_4189);
and U5152 (N_5152,N_4267,N_4426);
nor U5153 (N_5153,N_4560,N_4133);
and U5154 (N_5154,N_4492,N_4079);
or U5155 (N_5155,N_4156,N_4552);
xor U5156 (N_5156,N_4336,N_4277);
and U5157 (N_5157,N_4327,N_4244);
nand U5158 (N_5158,N_4505,N_4770);
or U5159 (N_5159,N_4113,N_4533);
or U5160 (N_5160,N_4929,N_4565);
xor U5161 (N_5161,N_4621,N_4891);
or U5162 (N_5162,N_4385,N_4588);
xnor U5163 (N_5163,N_4987,N_4347);
xor U5164 (N_5164,N_4425,N_4059);
and U5165 (N_5165,N_4819,N_4254);
xor U5166 (N_5166,N_4099,N_4257);
and U5167 (N_5167,N_4326,N_4916);
and U5168 (N_5168,N_4020,N_4041);
and U5169 (N_5169,N_4086,N_4886);
xnor U5170 (N_5170,N_4117,N_4436);
or U5171 (N_5171,N_4447,N_4564);
xor U5172 (N_5172,N_4814,N_4094);
and U5173 (N_5173,N_4640,N_4995);
nand U5174 (N_5174,N_4392,N_4517);
or U5175 (N_5175,N_4461,N_4638);
nor U5176 (N_5176,N_4789,N_4173);
and U5177 (N_5177,N_4273,N_4574);
xnor U5178 (N_5178,N_4614,N_4639);
and U5179 (N_5179,N_4467,N_4799);
xnor U5180 (N_5180,N_4234,N_4876);
nor U5181 (N_5181,N_4731,N_4429);
xnor U5182 (N_5182,N_4902,N_4790);
and U5183 (N_5183,N_4584,N_4356);
nand U5184 (N_5184,N_4690,N_4944);
and U5185 (N_5185,N_4274,N_4881);
nor U5186 (N_5186,N_4620,N_4317);
nor U5187 (N_5187,N_4617,N_4421);
or U5188 (N_5188,N_4297,N_4043);
nand U5189 (N_5189,N_4207,N_4296);
nor U5190 (N_5190,N_4285,N_4825);
and U5191 (N_5191,N_4493,N_4926);
or U5192 (N_5192,N_4313,N_4969);
nor U5193 (N_5193,N_4511,N_4367);
or U5194 (N_5194,N_4974,N_4023);
xor U5195 (N_5195,N_4888,N_4836);
nor U5196 (N_5196,N_4628,N_4885);
xnor U5197 (N_5197,N_4708,N_4951);
and U5198 (N_5198,N_4226,N_4872);
or U5199 (N_5199,N_4939,N_4666);
or U5200 (N_5200,N_4756,N_4322);
xnor U5201 (N_5201,N_4798,N_4068);
and U5202 (N_5202,N_4451,N_4514);
xnor U5203 (N_5203,N_4854,N_4613);
xor U5204 (N_5204,N_4141,N_4759);
or U5205 (N_5205,N_4146,N_4123);
and U5206 (N_5206,N_4082,N_4701);
or U5207 (N_5207,N_4211,N_4937);
or U5208 (N_5208,N_4489,N_4378);
and U5209 (N_5209,N_4066,N_4658);
or U5210 (N_5210,N_4359,N_4157);
and U5211 (N_5211,N_4018,N_4375);
or U5212 (N_5212,N_4214,N_4163);
xor U5213 (N_5213,N_4861,N_4350);
or U5214 (N_5214,N_4000,N_4203);
nand U5215 (N_5215,N_4569,N_4864);
nor U5216 (N_5216,N_4774,N_4152);
xor U5217 (N_5217,N_4778,N_4527);
nor U5218 (N_5218,N_4566,N_4900);
nand U5219 (N_5219,N_4635,N_4548);
nor U5220 (N_5220,N_4721,N_4949);
nor U5221 (N_5221,N_4188,N_4098);
or U5222 (N_5222,N_4587,N_4225);
and U5223 (N_5223,N_4928,N_4158);
xor U5224 (N_5224,N_4829,N_4583);
or U5225 (N_5225,N_4890,N_4407);
and U5226 (N_5226,N_4216,N_4947);
nor U5227 (N_5227,N_4093,N_4011);
xor U5228 (N_5228,N_4521,N_4490);
and U5229 (N_5229,N_4850,N_4344);
and U5230 (N_5230,N_4568,N_4387);
or U5231 (N_5231,N_4870,N_4428);
nor U5232 (N_5232,N_4119,N_4266);
nand U5233 (N_5233,N_4807,N_4749);
nand U5234 (N_5234,N_4873,N_4072);
and U5235 (N_5235,N_4270,N_4848);
nor U5236 (N_5236,N_4388,N_4482);
and U5237 (N_5237,N_4185,N_4365);
nor U5238 (N_5238,N_4842,N_4924);
and U5239 (N_5239,N_4232,N_4452);
and U5240 (N_5240,N_4175,N_4488);
xnor U5241 (N_5241,N_4053,N_4700);
and U5242 (N_5242,N_4791,N_4849);
or U5243 (N_5243,N_4383,N_4166);
xnor U5244 (N_5244,N_4840,N_4435);
nand U5245 (N_5245,N_4503,N_4218);
nand U5246 (N_5246,N_4652,N_4364);
nor U5247 (N_5247,N_4268,N_4785);
xor U5248 (N_5248,N_4139,N_4380);
nor U5249 (N_5249,N_4439,N_4275);
nand U5250 (N_5250,N_4990,N_4808);
nor U5251 (N_5251,N_4554,N_4417);
nor U5252 (N_5252,N_4882,N_4931);
xnor U5253 (N_5253,N_4834,N_4538);
nand U5254 (N_5254,N_4718,N_4953);
and U5255 (N_5255,N_4917,N_4862);
nand U5256 (N_5256,N_4867,N_4875);
or U5257 (N_5257,N_4856,N_4999);
nor U5258 (N_5258,N_4570,N_4389);
or U5259 (N_5259,N_4052,N_4116);
xnor U5260 (N_5260,N_4932,N_4580);
or U5261 (N_5261,N_4980,N_4938);
nor U5262 (N_5262,N_4950,N_4228);
nand U5263 (N_5263,N_4127,N_4282);
or U5264 (N_5264,N_4197,N_4050);
and U5265 (N_5265,N_4180,N_4022);
xnor U5266 (N_5266,N_4831,N_4305);
nand U5267 (N_5267,N_4414,N_4415);
nand U5268 (N_5268,N_4391,N_4957);
nor U5269 (N_5269,N_4309,N_4130);
or U5270 (N_5270,N_4487,N_4418);
and U5271 (N_5271,N_4499,N_4970);
xor U5272 (N_5272,N_4696,N_4184);
nand U5273 (N_5273,N_4644,N_4142);
or U5274 (N_5274,N_4170,N_4051);
xor U5275 (N_5275,N_4255,N_4930);
or U5276 (N_5276,N_4301,N_4984);
nor U5277 (N_5277,N_4160,N_4403);
and U5278 (N_5278,N_4684,N_4822);
or U5279 (N_5279,N_4280,N_4754);
or U5280 (N_5280,N_4973,N_4095);
nor U5281 (N_5281,N_4762,N_4781);
nor U5282 (N_5282,N_4078,N_4105);
and U5283 (N_5283,N_4190,N_4223);
nor U5284 (N_5284,N_4017,N_4431);
and U5285 (N_5285,N_4765,N_4115);
nand U5286 (N_5286,N_4542,N_4222);
and U5287 (N_5287,N_4298,N_4670);
or U5288 (N_5288,N_4963,N_4717);
or U5289 (N_5289,N_4983,N_4460);
or U5290 (N_5290,N_4596,N_4678);
nor U5291 (N_5291,N_4826,N_4828);
xnor U5292 (N_5292,N_4667,N_4656);
or U5293 (N_5293,N_4054,N_4325);
nand U5294 (N_5294,N_4795,N_4904);
nor U5295 (N_5295,N_4131,N_4551);
or U5296 (N_5296,N_4338,N_4982);
and U5297 (N_5297,N_4179,N_4402);
xor U5298 (N_5298,N_4048,N_4486);
nand U5299 (N_5299,N_4709,N_4061);
nand U5300 (N_5300,N_4331,N_4433);
nand U5301 (N_5301,N_4441,N_4634);
nand U5302 (N_5302,N_4256,N_4893);
nor U5303 (N_5303,N_4752,N_4408);
or U5304 (N_5304,N_4231,N_4962);
or U5305 (N_5305,N_4645,N_4019);
and U5306 (N_5306,N_4107,N_4668);
or U5307 (N_5307,N_4633,N_4324);
and U5308 (N_5308,N_4237,N_4713);
nor U5309 (N_5309,N_4776,N_4835);
and U5310 (N_5310,N_4600,N_4101);
nor U5311 (N_5311,N_4186,N_4985);
and U5312 (N_5312,N_4857,N_4518);
nand U5313 (N_5313,N_4281,N_4777);
and U5314 (N_5314,N_4906,N_4074);
and U5315 (N_5315,N_4150,N_4196);
or U5316 (N_5316,N_4056,N_4685);
and U5317 (N_5317,N_4215,N_4007);
nand U5318 (N_5318,N_4719,N_4591);
xor U5319 (N_5319,N_4144,N_4149);
xor U5320 (N_5320,N_4262,N_4959);
xor U5321 (N_5321,N_4357,N_4476);
nand U5322 (N_5322,N_4259,N_4535);
xor U5323 (N_5323,N_4961,N_4859);
nor U5324 (N_5324,N_4443,N_4540);
and U5325 (N_5325,N_4128,N_4221);
and U5326 (N_5326,N_4126,N_4913);
and U5327 (N_5327,N_4159,N_4833);
or U5328 (N_5328,N_4406,N_4952);
nand U5329 (N_5329,N_4145,N_4556);
or U5330 (N_5330,N_4653,N_4803);
xor U5331 (N_5331,N_4539,N_4311);
or U5332 (N_5332,N_4293,N_4288);
or U5333 (N_5333,N_4132,N_4761);
nand U5334 (N_5334,N_4729,N_4993);
and U5335 (N_5335,N_4034,N_4124);
nor U5336 (N_5336,N_4333,N_4657);
nand U5337 (N_5337,N_4648,N_4976);
xnor U5338 (N_5338,N_4351,N_4155);
nor U5339 (N_5339,N_4251,N_4049);
xor U5340 (N_5340,N_4945,N_4269);
xor U5341 (N_5341,N_4377,N_4988);
xnor U5342 (N_5342,N_4806,N_4531);
and U5343 (N_5343,N_4737,N_4136);
nand U5344 (N_5344,N_4349,N_4384);
xnor U5345 (N_5345,N_4664,N_4625);
or U5346 (N_5346,N_4510,N_4674);
nor U5347 (N_5347,N_4420,N_4168);
and U5348 (N_5348,N_4182,N_4530);
and U5349 (N_5349,N_4601,N_4830);
nand U5350 (N_5350,N_4837,N_4573);
or U5351 (N_5351,N_4497,N_4823);
nand U5352 (N_5352,N_4161,N_4394);
xor U5353 (N_5353,N_4524,N_4212);
and U5354 (N_5354,N_4064,N_4442);
xnor U5355 (N_5355,N_4084,N_4006);
or U5356 (N_5356,N_4763,N_4688);
or U5357 (N_5357,N_4318,N_4191);
or U5358 (N_5358,N_4884,N_4075);
xor U5359 (N_5359,N_4129,N_4138);
nand U5360 (N_5360,N_4302,N_4024);
or U5361 (N_5361,N_4475,N_4090);
or U5362 (N_5362,N_4100,N_4581);
nand U5363 (N_5363,N_4779,N_4005);
xnor U5364 (N_5364,N_4076,N_4077);
or U5365 (N_5365,N_4199,N_4846);
and U5366 (N_5366,N_4470,N_4557);
and U5367 (N_5367,N_4046,N_4676);
or U5368 (N_5368,N_4004,N_4401);
xor U5369 (N_5369,N_4632,N_4073);
or U5370 (N_5370,N_4522,N_4865);
nor U5371 (N_5371,N_4063,N_4174);
nand U5372 (N_5372,N_4991,N_4148);
xor U5373 (N_5373,N_4089,N_4330);
nand U5374 (N_5374,N_4382,N_4413);
and U5375 (N_5375,N_4567,N_4410);
and U5376 (N_5376,N_4264,N_4303);
nand U5377 (N_5377,N_4172,N_4942);
nand U5378 (N_5378,N_4108,N_4593);
xnor U5379 (N_5379,N_4604,N_4733);
xor U5380 (N_5380,N_4374,N_4008);
nor U5381 (N_5381,N_4863,N_4553);
nor U5382 (N_5382,N_4292,N_4544);
and U5383 (N_5383,N_4143,N_4686);
or U5384 (N_5384,N_4412,N_4750);
nand U5385 (N_5385,N_4220,N_4271);
and U5386 (N_5386,N_4474,N_4286);
nand U5387 (N_5387,N_4337,N_4080);
and U5388 (N_5388,N_4693,N_4206);
xnor U5389 (N_5389,N_4195,N_4824);
nand U5390 (N_5390,N_4874,N_4395);
xnor U5391 (N_5391,N_4120,N_4740);
xnor U5392 (N_5392,N_4036,N_4927);
nor U5393 (N_5393,N_4908,N_4484);
nor U5394 (N_5394,N_4543,N_4577);
nor U5395 (N_5395,N_4720,N_4422);
xnor U5396 (N_5396,N_4370,N_4342);
nand U5397 (N_5397,N_4466,N_4464);
and U5398 (N_5398,N_4905,N_4711);
and U5399 (N_5399,N_4513,N_4682);
nand U5400 (N_5400,N_4794,N_4946);
xnor U5401 (N_5401,N_4319,N_4880);
or U5402 (N_5402,N_4496,N_4677);
and U5403 (N_5403,N_4310,N_4784);
nor U5404 (N_5404,N_4923,N_4832);
xnor U5405 (N_5405,N_4853,N_4332);
nor U5406 (N_5406,N_4630,N_4109);
nor U5407 (N_5407,N_4261,N_4456);
nand U5408 (N_5408,N_4276,N_4899);
nor U5409 (N_5409,N_4390,N_4590);
and U5410 (N_5410,N_4169,N_4278);
and U5411 (N_5411,N_4473,N_4769);
nand U5412 (N_5412,N_4605,N_4404);
xnor U5413 (N_5413,N_4346,N_4289);
or U5414 (N_5414,N_4792,N_4673);
or U5415 (N_5415,N_4576,N_4386);
or U5416 (N_5416,N_4925,N_4205);
nand U5417 (N_5417,N_4796,N_4448);
nor U5418 (N_5418,N_4015,N_4354);
nor U5419 (N_5419,N_4675,N_4029);
xnor U5420 (N_5420,N_4176,N_4245);
or U5421 (N_5421,N_4631,N_4578);
or U5422 (N_5422,N_4935,N_4423);
nand U5423 (N_5423,N_4444,N_4233);
or U5424 (N_5424,N_4037,N_4012);
and U5425 (N_5425,N_4481,N_4646);
nor U5426 (N_5426,N_4647,N_4209);
or U5427 (N_5427,N_4933,N_4471);
nand U5428 (N_5428,N_4541,N_4764);
nor U5429 (N_5429,N_4151,N_4555);
or U5430 (N_5430,N_4110,N_4642);
and U5431 (N_5431,N_4851,N_4192);
nor U5432 (N_5432,N_4545,N_4745);
and U5433 (N_5433,N_4026,N_4477);
nand U5434 (N_5434,N_4446,N_4334);
xor U5435 (N_5435,N_4681,N_4515);
and U5436 (N_5436,N_4699,N_4224);
and U5437 (N_5437,N_4167,N_4028);
xnor U5438 (N_5438,N_4219,N_4744);
nand U5439 (N_5439,N_4252,N_4537);
or U5440 (N_5440,N_4878,N_4352);
or U5441 (N_5441,N_4340,N_4966);
or U5442 (N_5442,N_4852,N_4622);
and U5443 (N_5443,N_4118,N_4284);
nand U5444 (N_5444,N_4147,N_4877);
xnor U5445 (N_5445,N_4901,N_4751);
xnor U5446 (N_5446,N_4345,N_4869);
or U5447 (N_5447,N_4986,N_4616);
or U5448 (N_5448,N_4817,N_4562);
nor U5449 (N_5449,N_4312,N_4247);
nor U5450 (N_5450,N_4558,N_4459);
or U5451 (N_5451,N_4283,N_4651);
or U5452 (N_5452,N_4405,N_4705);
and U5453 (N_5453,N_4516,N_4253);
and U5454 (N_5454,N_4057,N_4287);
xnor U5455 (N_5455,N_4372,N_4134);
and U5456 (N_5456,N_4200,N_4279);
or U5457 (N_5457,N_4092,N_4889);
nor U5458 (N_5458,N_4472,N_4229);
or U5459 (N_5459,N_4454,N_4314);
nor U5460 (N_5460,N_4307,N_4495);
xnor U5461 (N_5461,N_4316,N_4217);
or U5462 (N_5462,N_4606,N_4525);
and U5463 (N_5463,N_4494,N_4526);
nor U5464 (N_5464,N_4722,N_4363);
nor U5465 (N_5465,N_4070,N_4907);
nand U5466 (N_5466,N_4171,N_4592);
nor U5467 (N_5467,N_4706,N_4626);
nor U5468 (N_5468,N_4122,N_4091);
or U5469 (N_5469,N_4424,N_4071);
and U5470 (N_5470,N_4793,N_4595);
nor U5471 (N_5471,N_4536,N_4920);
nand U5472 (N_5472,N_4561,N_4246);
nand U5473 (N_5473,N_4396,N_4081);
nand U5474 (N_5474,N_4111,N_4607);
nand U5475 (N_5475,N_4896,N_4371);
or U5476 (N_5476,N_4768,N_4087);
or U5477 (N_5477,N_4910,N_4003);
and U5478 (N_5478,N_4096,N_4743);
and U5479 (N_5479,N_4125,N_4694);
or U5480 (N_5480,N_4434,N_4501);
nor U5481 (N_5481,N_4178,N_4911);
or U5482 (N_5482,N_4599,N_4450);
nand U5483 (N_5483,N_4315,N_4689);
nand U5484 (N_5484,N_4797,N_4655);
nand U5485 (N_5485,N_4843,N_4088);
nand U5486 (N_5486,N_4958,N_4308);
xor U5487 (N_5487,N_4358,N_4559);
or U5488 (N_5488,N_4001,N_4773);
or U5489 (N_5489,N_4104,N_4040);
nor U5490 (N_5490,N_4895,N_4611);
nor U5491 (N_5491,N_4683,N_4323);
nand U5492 (N_5492,N_4812,N_4243);
xor U5493 (N_5493,N_4198,N_4809);
and U5494 (N_5494,N_4265,N_4379);
nand U5495 (N_5495,N_4419,N_4816);
nand U5496 (N_5496,N_4724,N_4956);
and U5497 (N_5497,N_4035,N_4097);
nand U5498 (N_5498,N_4304,N_4636);
and U5499 (N_5499,N_4067,N_4921);
xor U5500 (N_5500,N_4305,N_4095);
and U5501 (N_5501,N_4305,N_4390);
nor U5502 (N_5502,N_4570,N_4871);
nand U5503 (N_5503,N_4382,N_4502);
nand U5504 (N_5504,N_4117,N_4669);
xor U5505 (N_5505,N_4296,N_4600);
nor U5506 (N_5506,N_4715,N_4375);
and U5507 (N_5507,N_4040,N_4815);
nor U5508 (N_5508,N_4283,N_4478);
xnor U5509 (N_5509,N_4084,N_4347);
nand U5510 (N_5510,N_4543,N_4523);
or U5511 (N_5511,N_4284,N_4113);
nand U5512 (N_5512,N_4078,N_4711);
nor U5513 (N_5513,N_4310,N_4232);
nand U5514 (N_5514,N_4442,N_4289);
nand U5515 (N_5515,N_4802,N_4921);
or U5516 (N_5516,N_4750,N_4765);
or U5517 (N_5517,N_4690,N_4217);
xor U5518 (N_5518,N_4554,N_4355);
nand U5519 (N_5519,N_4813,N_4231);
and U5520 (N_5520,N_4628,N_4941);
xnor U5521 (N_5521,N_4634,N_4313);
nor U5522 (N_5522,N_4200,N_4787);
nor U5523 (N_5523,N_4759,N_4462);
nor U5524 (N_5524,N_4535,N_4553);
and U5525 (N_5525,N_4007,N_4253);
and U5526 (N_5526,N_4366,N_4250);
xnor U5527 (N_5527,N_4382,N_4895);
xnor U5528 (N_5528,N_4958,N_4457);
and U5529 (N_5529,N_4705,N_4328);
or U5530 (N_5530,N_4693,N_4955);
and U5531 (N_5531,N_4914,N_4383);
nor U5532 (N_5532,N_4639,N_4874);
nand U5533 (N_5533,N_4602,N_4721);
xor U5534 (N_5534,N_4414,N_4015);
and U5535 (N_5535,N_4911,N_4326);
or U5536 (N_5536,N_4973,N_4986);
or U5537 (N_5537,N_4965,N_4942);
and U5538 (N_5538,N_4205,N_4643);
xor U5539 (N_5539,N_4946,N_4348);
or U5540 (N_5540,N_4193,N_4620);
or U5541 (N_5541,N_4723,N_4146);
xnor U5542 (N_5542,N_4614,N_4113);
nand U5543 (N_5543,N_4138,N_4093);
xor U5544 (N_5544,N_4558,N_4987);
nor U5545 (N_5545,N_4661,N_4319);
xor U5546 (N_5546,N_4980,N_4899);
nand U5547 (N_5547,N_4116,N_4879);
and U5548 (N_5548,N_4866,N_4234);
xnor U5549 (N_5549,N_4782,N_4278);
and U5550 (N_5550,N_4811,N_4180);
nand U5551 (N_5551,N_4104,N_4316);
xnor U5552 (N_5552,N_4965,N_4889);
nor U5553 (N_5553,N_4247,N_4012);
nor U5554 (N_5554,N_4382,N_4812);
nand U5555 (N_5555,N_4606,N_4459);
nor U5556 (N_5556,N_4431,N_4478);
xnor U5557 (N_5557,N_4329,N_4476);
nand U5558 (N_5558,N_4869,N_4566);
xnor U5559 (N_5559,N_4162,N_4980);
and U5560 (N_5560,N_4336,N_4157);
xnor U5561 (N_5561,N_4457,N_4769);
nor U5562 (N_5562,N_4653,N_4944);
and U5563 (N_5563,N_4464,N_4096);
nor U5564 (N_5564,N_4311,N_4183);
xor U5565 (N_5565,N_4069,N_4537);
nand U5566 (N_5566,N_4862,N_4281);
or U5567 (N_5567,N_4553,N_4777);
nand U5568 (N_5568,N_4955,N_4488);
nand U5569 (N_5569,N_4757,N_4434);
and U5570 (N_5570,N_4906,N_4028);
and U5571 (N_5571,N_4072,N_4248);
nor U5572 (N_5572,N_4969,N_4105);
nand U5573 (N_5573,N_4760,N_4404);
and U5574 (N_5574,N_4848,N_4914);
and U5575 (N_5575,N_4646,N_4391);
nor U5576 (N_5576,N_4344,N_4668);
nor U5577 (N_5577,N_4980,N_4044);
xor U5578 (N_5578,N_4074,N_4232);
and U5579 (N_5579,N_4346,N_4689);
and U5580 (N_5580,N_4133,N_4096);
and U5581 (N_5581,N_4226,N_4741);
or U5582 (N_5582,N_4871,N_4892);
nor U5583 (N_5583,N_4010,N_4570);
xnor U5584 (N_5584,N_4391,N_4547);
nor U5585 (N_5585,N_4324,N_4275);
or U5586 (N_5586,N_4586,N_4517);
nand U5587 (N_5587,N_4902,N_4114);
or U5588 (N_5588,N_4825,N_4595);
or U5589 (N_5589,N_4415,N_4882);
or U5590 (N_5590,N_4225,N_4643);
nor U5591 (N_5591,N_4479,N_4231);
nor U5592 (N_5592,N_4941,N_4986);
xnor U5593 (N_5593,N_4989,N_4542);
xor U5594 (N_5594,N_4686,N_4641);
nand U5595 (N_5595,N_4452,N_4294);
nand U5596 (N_5596,N_4250,N_4084);
nand U5597 (N_5597,N_4390,N_4995);
nor U5598 (N_5598,N_4480,N_4076);
or U5599 (N_5599,N_4933,N_4045);
xor U5600 (N_5600,N_4175,N_4772);
and U5601 (N_5601,N_4471,N_4379);
xnor U5602 (N_5602,N_4666,N_4265);
nor U5603 (N_5603,N_4445,N_4263);
or U5604 (N_5604,N_4054,N_4785);
nor U5605 (N_5605,N_4863,N_4480);
xnor U5606 (N_5606,N_4701,N_4608);
nor U5607 (N_5607,N_4059,N_4681);
or U5608 (N_5608,N_4895,N_4718);
or U5609 (N_5609,N_4271,N_4593);
nor U5610 (N_5610,N_4636,N_4911);
or U5611 (N_5611,N_4490,N_4334);
nor U5612 (N_5612,N_4290,N_4901);
nor U5613 (N_5613,N_4639,N_4688);
and U5614 (N_5614,N_4984,N_4795);
nor U5615 (N_5615,N_4572,N_4717);
or U5616 (N_5616,N_4610,N_4392);
or U5617 (N_5617,N_4641,N_4827);
or U5618 (N_5618,N_4878,N_4247);
or U5619 (N_5619,N_4851,N_4673);
nor U5620 (N_5620,N_4330,N_4222);
nor U5621 (N_5621,N_4413,N_4732);
nand U5622 (N_5622,N_4320,N_4355);
xnor U5623 (N_5623,N_4402,N_4231);
and U5624 (N_5624,N_4376,N_4691);
nand U5625 (N_5625,N_4065,N_4259);
or U5626 (N_5626,N_4257,N_4402);
and U5627 (N_5627,N_4603,N_4628);
xor U5628 (N_5628,N_4914,N_4085);
xnor U5629 (N_5629,N_4635,N_4169);
nor U5630 (N_5630,N_4827,N_4460);
nand U5631 (N_5631,N_4555,N_4646);
or U5632 (N_5632,N_4093,N_4082);
nand U5633 (N_5633,N_4258,N_4403);
nand U5634 (N_5634,N_4124,N_4304);
or U5635 (N_5635,N_4650,N_4443);
nand U5636 (N_5636,N_4199,N_4054);
nor U5637 (N_5637,N_4632,N_4340);
xnor U5638 (N_5638,N_4868,N_4919);
and U5639 (N_5639,N_4583,N_4497);
and U5640 (N_5640,N_4225,N_4615);
and U5641 (N_5641,N_4396,N_4601);
or U5642 (N_5642,N_4136,N_4093);
or U5643 (N_5643,N_4040,N_4509);
and U5644 (N_5644,N_4221,N_4373);
nor U5645 (N_5645,N_4302,N_4088);
and U5646 (N_5646,N_4911,N_4369);
or U5647 (N_5647,N_4075,N_4520);
xnor U5648 (N_5648,N_4852,N_4917);
or U5649 (N_5649,N_4411,N_4055);
or U5650 (N_5650,N_4155,N_4196);
nor U5651 (N_5651,N_4384,N_4718);
nor U5652 (N_5652,N_4481,N_4230);
and U5653 (N_5653,N_4925,N_4761);
nor U5654 (N_5654,N_4534,N_4624);
xor U5655 (N_5655,N_4675,N_4891);
or U5656 (N_5656,N_4132,N_4215);
nor U5657 (N_5657,N_4595,N_4245);
nand U5658 (N_5658,N_4604,N_4317);
and U5659 (N_5659,N_4327,N_4570);
xnor U5660 (N_5660,N_4644,N_4505);
nor U5661 (N_5661,N_4863,N_4017);
or U5662 (N_5662,N_4653,N_4062);
xnor U5663 (N_5663,N_4566,N_4435);
nand U5664 (N_5664,N_4269,N_4106);
xnor U5665 (N_5665,N_4227,N_4050);
xnor U5666 (N_5666,N_4072,N_4501);
and U5667 (N_5667,N_4488,N_4328);
nor U5668 (N_5668,N_4991,N_4274);
nand U5669 (N_5669,N_4100,N_4670);
and U5670 (N_5670,N_4569,N_4763);
and U5671 (N_5671,N_4815,N_4151);
nand U5672 (N_5672,N_4687,N_4622);
xor U5673 (N_5673,N_4300,N_4372);
or U5674 (N_5674,N_4058,N_4940);
or U5675 (N_5675,N_4424,N_4149);
nor U5676 (N_5676,N_4500,N_4990);
xor U5677 (N_5677,N_4362,N_4230);
or U5678 (N_5678,N_4938,N_4799);
nand U5679 (N_5679,N_4848,N_4173);
or U5680 (N_5680,N_4617,N_4261);
and U5681 (N_5681,N_4229,N_4095);
and U5682 (N_5682,N_4917,N_4842);
xnor U5683 (N_5683,N_4937,N_4281);
xor U5684 (N_5684,N_4358,N_4880);
or U5685 (N_5685,N_4926,N_4190);
and U5686 (N_5686,N_4686,N_4112);
and U5687 (N_5687,N_4281,N_4191);
nor U5688 (N_5688,N_4334,N_4153);
nor U5689 (N_5689,N_4935,N_4562);
nand U5690 (N_5690,N_4106,N_4824);
nor U5691 (N_5691,N_4940,N_4355);
and U5692 (N_5692,N_4330,N_4589);
and U5693 (N_5693,N_4893,N_4335);
xnor U5694 (N_5694,N_4269,N_4176);
xor U5695 (N_5695,N_4196,N_4465);
xnor U5696 (N_5696,N_4755,N_4048);
and U5697 (N_5697,N_4535,N_4866);
nand U5698 (N_5698,N_4829,N_4333);
xnor U5699 (N_5699,N_4681,N_4592);
and U5700 (N_5700,N_4818,N_4520);
and U5701 (N_5701,N_4007,N_4588);
and U5702 (N_5702,N_4608,N_4171);
or U5703 (N_5703,N_4977,N_4902);
nor U5704 (N_5704,N_4586,N_4166);
nor U5705 (N_5705,N_4988,N_4611);
nor U5706 (N_5706,N_4925,N_4585);
nor U5707 (N_5707,N_4477,N_4386);
xor U5708 (N_5708,N_4761,N_4483);
nor U5709 (N_5709,N_4316,N_4056);
nor U5710 (N_5710,N_4826,N_4062);
and U5711 (N_5711,N_4777,N_4965);
nor U5712 (N_5712,N_4388,N_4443);
or U5713 (N_5713,N_4487,N_4819);
nand U5714 (N_5714,N_4872,N_4551);
nand U5715 (N_5715,N_4284,N_4149);
nand U5716 (N_5716,N_4703,N_4684);
and U5717 (N_5717,N_4556,N_4772);
nor U5718 (N_5718,N_4542,N_4851);
nand U5719 (N_5719,N_4322,N_4425);
nor U5720 (N_5720,N_4389,N_4338);
nor U5721 (N_5721,N_4086,N_4526);
or U5722 (N_5722,N_4146,N_4201);
nor U5723 (N_5723,N_4907,N_4383);
nor U5724 (N_5724,N_4271,N_4856);
and U5725 (N_5725,N_4948,N_4438);
nand U5726 (N_5726,N_4098,N_4192);
xnor U5727 (N_5727,N_4320,N_4931);
xor U5728 (N_5728,N_4627,N_4840);
xnor U5729 (N_5729,N_4954,N_4068);
xor U5730 (N_5730,N_4372,N_4891);
and U5731 (N_5731,N_4512,N_4137);
or U5732 (N_5732,N_4309,N_4858);
nor U5733 (N_5733,N_4357,N_4099);
xor U5734 (N_5734,N_4087,N_4120);
nand U5735 (N_5735,N_4685,N_4317);
nor U5736 (N_5736,N_4675,N_4159);
nor U5737 (N_5737,N_4520,N_4606);
nand U5738 (N_5738,N_4288,N_4233);
xnor U5739 (N_5739,N_4383,N_4707);
or U5740 (N_5740,N_4381,N_4883);
and U5741 (N_5741,N_4410,N_4517);
nand U5742 (N_5742,N_4230,N_4467);
and U5743 (N_5743,N_4267,N_4638);
and U5744 (N_5744,N_4576,N_4887);
or U5745 (N_5745,N_4624,N_4617);
nor U5746 (N_5746,N_4790,N_4752);
or U5747 (N_5747,N_4537,N_4511);
and U5748 (N_5748,N_4983,N_4234);
nor U5749 (N_5749,N_4953,N_4240);
nand U5750 (N_5750,N_4223,N_4719);
nand U5751 (N_5751,N_4570,N_4075);
and U5752 (N_5752,N_4570,N_4691);
or U5753 (N_5753,N_4907,N_4984);
nand U5754 (N_5754,N_4548,N_4035);
nand U5755 (N_5755,N_4698,N_4697);
or U5756 (N_5756,N_4127,N_4994);
and U5757 (N_5757,N_4994,N_4789);
or U5758 (N_5758,N_4131,N_4872);
nand U5759 (N_5759,N_4086,N_4339);
xnor U5760 (N_5760,N_4335,N_4156);
nor U5761 (N_5761,N_4753,N_4269);
nand U5762 (N_5762,N_4452,N_4271);
xnor U5763 (N_5763,N_4170,N_4891);
nand U5764 (N_5764,N_4816,N_4677);
nand U5765 (N_5765,N_4847,N_4841);
or U5766 (N_5766,N_4140,N_4153);
or U5767 (N_5767,N_4562,N_4443);
and U5768 (N_5768,N_4131,N_4335);
or U5769 (N_5769,N_4638,N_4259);
and U5770 (N_5770,N_4964,N_4427);
xnor U5771 (N_5771,N_4856,N_4413);
or U5772 (N_5772,N_4239,N_4321);
nor U5773 (N_5773,N_4348,N_4027);
nand U5774 (N_5774,N_4136,N_4243);
nor U5775 (N_5775,N_4081,N_4962);
and U5776 (N_5776,N_4885,N_4784);
and U5777 (N_5777,N_4209,N_4589);
nor U5778 (N_5778,N_4194,N_4526);
nor U5779 (N_5779,N_4612,N_4276);
nor U5780 (N_5780,N_4326,N_4062);
or U5781 (N_5781,N_4460,N_4876);
and U5782 (N_5782,N_4708,N_4434);
nor U5783 (N_5783,N_4679,N_4865);
or U5784 (N_5784,N_4929,N_4287);
or U5785 (N_5785,N_4425,N_4006);
nand U5786 (N_5786,N_4391,N_4220);
nor U5787 (N_5787,N_4068,N_4780);
or U5788 (N_5788,N_4474,N_4960);
and U5789 (N_5789,N_4646,N_4322);
nand U5790 (N_5790,N_4220,N_4198);
nand U5791 (N_5791,N_4325,N_4506);
nor U5792 (N_5792,N_4849,N_4525);
nor U5793 (N_5793,N_4597,N_4501);
or U5794 (N_5794,N_4885,N_4105);
and U5795 (N_5795,N_4802,N_4021);
nor U5796 (N_5796,N_4709,N_4164);
nor U5797 (N_5797,N_4835,N_4955);
or U5798 (N_5798,N_4963,N_4611);
xnor U5799 (N_5799,N_4953,N_4418);
nand U5800 (N_5800,N_4190,N_4226);
nor U5801 (N_5801,N_4611,N_4581);
xor U5802 (N_5802,N_4553,N_4251);
nor U5803 (N_5803,N_4803,N_4494);
or U5804 (N_5804,N_4697,N_4168);
nor U5805 (N_5805,N_4082,N_4192);
or U5806 (N_5806,N_4994,N_4441);
nand U5807 (N_5807,N_4169,N_4747);
nor U5808 (N_5808,N_4058,N_4883);
xnor U5809 (N_5809,N_4189,N_4098);
and U5810 (N_5810,N_4607,N_4543);
and U5811 (N_5811,N_4716,N_4654);
or U5812 (N_5812,N_4304,N_4170);
nand U5813 (N_5813,N_4526,N_4600);
and U5814 (N_5814,N_4165,N_4359);
nand U5815 (N_5815,N_4281,N_4871);
or U5816 (N_5816,N_4664,N_4006);
and U5817 (N_5817,N_4419,N_4378);
or U5818 (N_5818,N_4720,N_4498);
and U5819 (N_5819,N_4204,N_4032);
nor U5820 (N_5820,N_4556,N_4543);
or U5821 (N_5821,N_4795,N_4466);
xor U5822 (N_5822,N_4661,N_4906);
or U5823 (N_5823,N_4743,N_4762);
xor U5824 (N_5824,N_4958,N_4598);
nand U5825 (N_5825,N_4199,N_4642);
or U5826 (N_5826,N_4739,N_4245);
nand U5827 (N_5827,N_4341,N_4340);
and U5828 (N_5828,N_4376,N_4219);
nor U5829 (N_5829,N_4870,N_4140);
and U5830 (N_5830,N_4882,N_4031);
or U5831 (N_5831,N_4934,N_4574);
or U5832 (N_5832,N_4324,N_4197);
xor U5833 (N_5833,N_4057,N_4280);
nand U5834 (N_5834,N_4199,N_4678);
xnor U5835 (N_5835,N_4947,N_4763);
and U5836 (N_5836,N_4562,N_4908);
or U5837 (N_5837,N_4819,N_4508);
and U5838 (N_5838,N_4028,N_4182);
xor U5839 (N_5839,N_4762,N_4146);
nand U5840 (N_5840,N_4441,N_4817);
and U5841 (N_5841,N_4058,N_4202);
and U5842 (N_5842,N_4346,N_4440);
xnor U5843 (N_5843,N_4416,N_4902);
xor U5844 (N_5844,N_4102,N_4725);
or U5845 (N_5845,N_4088,N_4154);
nand U5846 (N_5846,N_4005,N_4587);
xnor U5847 (N_5847,N_4837,N_4105);
nor U5848 (N_5848,N_4973,N_4782);
nand U5849 (N_5849,N_4786,N_4853);
nand U5850 (N_5850,N_4313,N_4427);
or U5851 (N_5851,N_4457,N_4289);
nor U5852 (N_5852,N_4428,N_4275);
nand U5853 (N_5853,N_4274,N_4494);
nand U5854 (N_5854,N_4811,N_4913);
nor U5855 (N_5855,N_4765,N_4502);
and U5856 (N_5856,N_4183,N_4608);
and U5857 (N_5857,N_4383,N_4909);
and U5858 (N_5858,N_4812,N_4395);
xnor U5859 (N_5859,N_4614,N_4540);
nor U5860 (N_5860,N_4518,N_4043);
or U5861 (N_5861,N_4260,N_4640);
nand U5862 (N_5862,N_4983,N_4315);
or U5863 (N_5863,N_4091,N_4167);
xnor U5864 (N_5864,N_4478,N_4905);
nand U5865 (N_5865,N_4325,N_4815);
nor U5866 (N_5866,N_4787,N_4031);
xnor U5867 (N_5867,N_4945,N_4594);
nand U5868 (N_5868,N_4893,N_4157);
and U5869 (N_5869,N_4168,N_4139);
xor U5870 (N_5870,N_4970,N_4058);
nand U5871 (N_5871,N_4971,N_4609);
nand U5872 (N_5872,N_4035,N_4141);
and U5873 (N_5873,N_4150,N_4532);
or U5874 (N_5874,N_4458,N_4932);
nor U5875 (N_5875,N_4997,N_4030);
nor U5876 (N_5876,N_4504,N_4073);
xor U5877 (N_5877,N_4794,N_4078);
nand U5878 (N_5878,N_4999,N_4372);
xor U5879 (N_5879,N_4913,N_4179);
xnor U5880 (N_5880,N_4608,N_4405);
and U5881 (N_5881,N_4434,N_4903);
nand U5882 (N_5882,N_4846,N_4466);
and U5883 (N_5883,N_4100,N_4277);
nor U5884 (N_5884,N_4030,N_4406);
xnor U5885 (N_5885,N_4684,N_4939);
or U5886 (N_5886,N_4087,N_4066);
nor U5887 (N_5887,N_4549,N_4372);
nor U5888 (N_5888,N_4791,N_4356);
nand U5889 (N_5889,N_4019,N_4993);
or U5890 (N_5890,N_4837,N_4129);
xnor U5891 (N_5891,N_4260,N_4271);
and U5892 (N_5892,N_4302,N_4599);
nor U5893 (N_5893,N_4542,N_4667);
or U5894 (N_5894,N_4480,N_4506);
xnor U5895 (N_5895,N_4101,N_4112);
and U5896 (N_5896,N_4959,N_4620);
and U5897 (N_5897,N_4629,N_4800);
xor U5898 (N_5898,N_4454,N_4200);
or U5899 (N_5899,N_4693,N_4101);
and U5900 (N_5900,N_4723,N_4330);
xor U5901 (N_5901,N_4947,N_4716);
xnor U5902 (N_5902,N_4068,N_4384);
nor U5903 (N_5903,N_4289,N_4510);
nor U5904 (N_5904,N_4596,N_4731);
nor U5905 (N_5905,N_4886,N_4741);
and U5906 (N_5906,N_4270,N_4108);
xor U5907 (N_5907,N_4979,N_4311);
nor U5908 (N_5908,N_4678,N_4657);
nor U5909 (N_5909,N_4228,N_4915);
and U5910 (N_5910,N_4156,N_4450);
or U5911 (N_5911,N_4794,N_4369);
or U5912 (N_5912,N_4107,N_4334);
xnor U5913 (N_5913,N_4700,N_4019);
nand U5914 (N_5914,N_4917,N_4691);
xnor U5915 (N_5915,N_4965,N_4978);
xor U5916 (N_5916,N_4142,N_4120);
nand U5917 (N_5917,N_4753,N_4236);
and U5918 (N_5918,N_4789,N_4051);
nor U5919 (N_5919,N_4836,N_4892);
and U5920 (N_5920,N_4765,N_4194);
nand U5921 (N_5921,N_4093,N_4502);
nor U5922 (N_5922,N_4227,N_4085);
nor U5923 (N_5923,N_4593,N_4251);
or U5924 (N_5924,N_4681,N_4284);
nand U5925 (N_5925,N_4528,N_4987);
xor U5926 (N_5926,N_4885,N_4462);
nor U5927 (N_5927,N_4116,N_4838);
or U5928 (N_5928,N_4261,N_4291);
nor U5929 (N_5929,N_4281,N_4044);
nor U5930 (N_5930,N_4582,N_4893);
xor U5931 (N_5931,N_4556,N_4766);
and U5932 (N_5932,N_4828,N_4656);
xor U5933 (N_5933,N_4686,N_4776);
nand U5934 (N_5934,N_4389,N_4406);
xor U5935 (N_5935,N_4127,N_4764);
nor U5936 (N_5936,N_4444,N_4708);
or U5937 (N_5937,N_4942,N_4576);
nor U5938 (N_5938,N_4207,N_4407);
nand U5939 (N_5939,N_4755,N_4578);
nand U5940 (N_5940,N_4634,N_4338);
nor U5941 (N_5941,N_4176,N_4028);
and U5942 (N_5942,N_4622,N_4707);
nor U5943 (N_5943,N_4721,N_4757);
xor U5944 (N_5944,N_4306,N_4126);
nor U5945 (N_5945,N_4499,N_4007);
xor U5946 (N_5946,N_4216,N_4321);
and U5947 (N_5947,N_4178,N_4252);
and U5948 (N_5948,N_4835,N_4893);
and U5949 (N_5949,N_4510,N_4184);
and U5950 (N_5950,N_4053,N_4586);
nor U5951 (N_5951,N_4412,N_4823);
nand U5952 (N_5952,N_4138,N_4618);
and U5953 (N_5953,N_4772,N_4049);
xnor U5954 (N_5954,N_4265,N_4153);
or U5955 (N_5955,N_4366,N_4796);
xor U5956 (N_5956,N_4299,N_4818);
or U5957 (N_5957,N_4331,N_4901);
nor U5958 (N_5958,N_4290,N_4453);
xnor U5959 (N_5959,N_4385,N_4976);
or U5960 (N_5960,N_4872,N_4680);
nand U5961 (N_5961,N_4666,N_4335);
nand U5962 (N_5962,N_4971,N_4221);
and U5963 (N_5963,N_4380,N_4783);
nand U5964 (N_5964,N_4124,N_4816);
or U5965 (N_5965,N_4605,N_4092);
or U5966 (N_5966,N_4227,N_4710);
xor U5967 (N_5967,N_4918,N_4394);
or U5968 (N_5968,N_4529,N_4518);
nor U5969 (N_5969,N_4205,N_4061);
nand U5970 (N_5970,N_4413,N_4040);
nor U5971 (N_5971,N_4500,N_4362);
or U5972 (N_5972,N_4320,N_4647);
nor U5973 (N_5973,N_4913,N_4724);
or U5974 (N_5974,N_4532,N_4590);
or U5975 (N_5975,N_4238,N_4035);
and U5976 (N_5976,N_4299,N_4753);
nand U5977 (N_5977,N_4591,N_4621);
nor U5978 (N_5978,N_4554,N_4639);
nand U5979 (N_5979,N_4659,N_4875);
or U5980 (N_5980,N_4722,N_4313);
or U5981 (N_5981,N_4573,N_4752);
xor U5982 (N_5982,N_4913,N_4798);
or U5983 (N_5983,N_4285,N_4408);
nand U5984 (N_5984,N_4016,N_4871);
or U5985 (N_5985,N_4614,N_4973);
xor U5986 (N_5986,N_4996,N_4061);
and U5987 (N_5987,N_4507,N_4961);
or U5988 (N_5988,N_4649,N_4667);
nand U5989 (N_5989,N_4808,N_4377);
xor U5990 (N_5990,N_4915,N_4747);
xor U5991 (N_5991,N_4923,N_4471);
nand U5992 (N_5992,N_4623,N_4093);
or U5993 (N_5993,N_4595,N_4981);
nor U5994 (N_5994,N_4301,N_4687);
and U5995 (N_5995,N_4709,N_4226);
or U5996 (N_5996,N_4705,N_4458);
and U5997 (N_5997,N_4479,N_4742);
and U5998 (N_5998,N_4813,N_4463);
and U5999 (N_5999,N_4426,N_4329);
nor U6000 (N_6000,N_5771,N_5220);
and U6001 (N_6001,N_5773,N_5879);
and U6002 (N_6002,N_5467,N_5811);
nand U6003 (N_6003,N_5884,N_5036);
nor U6004 (N_6004,N_5170,N_5676);
and U6005 (N_6005,N_5164,N_5473);
xor U6006 (N_6006,N_5753,N_5685);
or U6007 (N_6007,N_5728,N_5695);
xor U6008 (N_6008,N_5292,N_5048);
or U6009 (N_6009,N_5304,N_5149);
or U6010 (N_6010,N_5871,N_5625);
nor U6011 (N_6011,N_5487,N_5984);
nor U6012 (N_6012,N_5863,N_5230);
xnor U6013 (N_6013,N_5612,N_5637);
and U6014 (N_6014,N_5877,N_5723);
and U6015 (N_6015,N_5881,N_5139);
nand U6016 (N_6016,N_5276,N_5092);
or U6017 (N_6017,N_5349,N_5039);
nor U6018 (N_6018,N_5354,N_5835);
nand U6019 (N_6019,N_5511,N_5334);
xor U6020 (N_6020,N_5035,N_5307);
or U6021 (N_6021,N_5576,N_5808);
or U6022 (N_6022,N_5528,N_5980);
nand U6023 (N_6023,N_5687,N_5256);
xor U6024 (N_6024,N_5194,N_5148);
nand U6025 (N_6025,N_5774,N_5804);
or U6026 (N_6026,N_5158,N_5971);
nor U6027 (N_6027,N_5024,N_5937);
nor U6028 (N_6028,N_5477,N_5744);
or U6029 (N_6029,N_5662,N_5490);
nor U6030 (N_6030,N_5111,N_5076);
and U6031 (N_6031,N_5059,N_5905);
nand U6032 (N_6032,N_5225,N_5664);
and U6033 (N_6033,N_5961,N_5845);
nor U6034 (N_6034,N_5031,N_5986);
nor U6035 (N_6035,N_5370,N_5834);
xor U6036 (N_6036,N_5926,N_5671);
xnor U6037 (N_6037,N_5632,N_5814);
nand U6038 (N_6038,N_5901,N_5428);
and U6039 (N_6039,N_5162,N_5897);
or U6040 (N_6040,N_5533,N_5656);
and U6041 (N_6041,N_5185,N_5118);
xor U6042 (N_6042,N_5572,N_5013);
or U6043 (N_6043,N_5481,N_5344);
nor U6044 (N_6044,N_5010,N_5776);
xor U6045 (N_6045,N_5563,N_5817);
nand U6046 (N_6046,N_5618,N_5357);
nand U6047 (N_6047,N_5130,N_5440);
nand U6048 (N_6048,N_5596,N_5343);
nor U6049 (N_6049,N_5271,N_5101);
and U6050 (N_6050,N_5274,N_5942);
nor U6051 (N_6051,N_5963,N_5075);
nor U6052 (N_6052,N_5177,N_5358);
nor U6053 (N_6053,N_5090,N_5785);
xnor U6054 (N_6054,N_5231,N_5923);
and U6055 (N_6055,N_5865,N_5616);
nor U6056 (N_6056,N_5306,N_5453);
or U6057 (N_6057,N_5260,N_5694);
or U6058 (N_6058,N_5526,N_5324);
xnor U6059 (N_6059,N_5506,N_5257);
xnor U6060 (N_6060,N_5883,N_5505);
xnor U6061 (N_6061,N_5957,N_5701);
nor U6062 (N_6062,N_5948,N_5916);
or U6063 (N_6063,N_5810,N_5998);
or U6064 (N_6064,N_5520,N_5837);
xnor U6065 (N_6065,N_5888,N_5109);
nor U6066 (N_6066,N_5770,N_5981);
xnor U6067 (N_6067,N_5407,N_5290);
or U6068 (N_6068,N_5064,N_5764);
or U6069 (N_6069,N_5868,N_5607);
nand U6070 (N_6070,N_5698,N_5012);
or U6071 (N_6071,N_5722,N_5550);
xor U6072 (N_6072,N_5468,N_5248);
and U6073 (N_6073,N_5283,N_5378);
and U6074 (N_6074,N_5931,N_5514);
nor U6075 (N_6075,N_5451,N_5583);
nor U6076 (N_6076,N_5673,N_5310);
nor U6077 (N_6077,N_5187,N_5458);
and U6078 (N_6078,N_5355,N_5930);
nor U6079 (N_6079,N_5706,N_5820);
xnor U6080 (N_6080,N_5859,N_5777);
nand U6081 (N_6081,N_5176,N_5669);
and U6082 (N_6082,N_5245,N_5831);
or U6083 (N_6083,N_5262,N_5345);
and U6084 (N_6084,N_5547,N_5661);
and U6085 (N_6085,N_5329,N_5847);
xor U6086 (N_6086,N_5026,N_5281);
xnor U6087 (N_6087,N_5134,N_5293);
and U6088 (N_6088,N_5207,N_5840);
xor U6089 (N_6089,N_5691,N_5087);
or U6090 (N_6090,N_5083,N_5175);
xor U6091 (N_6091,N_5030,N_5374);
or U6092 (N_6092,N_5760,N_5707);
or U6093 (N_6093,N_5161,N_5296);
xor U6094 (N_6094,N_5584,N_5277);
xor U6095 (N_6095,N_5047,N_5145);
nor U6096 (N_6096,N_5347,N_5014);
xor U6097 (N_6097,N_5392,N_5071);
and U6098 (N_6098,N_5767,N_5802);
and U6099 (N_6099,N_5546,N_5875);
nand U6100 (N_6100,N_5335,N_5366);
or U6101 (N_6101,N_5465,N_5735);
nor U6102 (N_6102,N_5179,N_5166);
or U6103 (N_6103,N_5917,N_5108);
xor U6104 (N_6104,N_5038,N_5094);
nand U6105 (N_6105,N_5002,N_5922);
xnor U6106 (N_6106,N_5388,N_5536);
nand U6107 (N_6107,N_5300,N_5739);
nor U6108 (N_6108,N_5809,N_5791);
or U6109 (N_6109,N_5507,N_5807);
nor U6110 (N_6110,N_5913,N_5023);
or U6111 (N_6111,N_5243,N_5967);
nand U6112 (N_6112,N_5794,N_5210);
xor U6113 (N_6113,N_5123,N_5700);
nand U6114 (N_6114,N_5912,N_5524);
and U6115 (N_6115,N_5822,N_5372);
and U6116 (N_6116,N_5085,N_5990);
nand U6117 (N_6117,N_5270,N_5610);
and U6118 (N_6118,N_5182,N_5034);
or U6119 (N_6119,N_5521,N_5951);
and U6120 (N_6120,N_5713,N_5716);
nor U6121 (N_6121,N_5019,N_5813);
or U6122 (N_6122,N_5525,N_5895);
and U6123 (N_6123,N_5549,N_5932);
or U6124 (N_6124,N_5915,N_5885);
or U6125 (N_6125,N_5833,N_5799);
nor U6126 (N_6126,N_5919,N_5982);
or U6127 (N_6127,N_5497,N_5124);
nor U6128 (N_6128,N_5201,N_5647);
xnor U6129 (N_6129,N_5436,N_5914);
and U6130 (N_6130,N_5630,N_5670);
nand U6131 (N_6131,N_5994,N_5155);
or U6132 (N_6132,N_5627,N_5899);
xor U6133 (N_6133,N_5122,N_5202);
or U6134 (N_6134,N_5054,N_5288);
nor U6135 (N_6135,N_5484,N_5621);
and U6136 (N_6136,N_5940,N_5244);
and U6137 (N_6137,N_5887,N_5353);
and U6138 (N_6138,N_5403,N_5754);
or U6139 (N_6139,N_5812,N_5159);
xnor U6140 (N_6140,N_5070,N_5099);
nor U6141 (N_6141,N_5504,N_5934);
or U6142 (N_6142,N_5255,N_5841);
and U6143 (N_6143,N_5876,N_5455);
nor U6144 (N_6144,N_5551,N_5489);
xor U6145 (N_6145,N_5861,N_5636);
xor U6146 (N_6146,N_5291,N_5638);
nor U6147 (N_6147,N_5667,N_5318);
nand U6148 (N_6148,N_5766,N_5120);
xnor U6149 (N_6149,N_5189,N_5874);
nand U6150 (N_6150,N_5780,N_5975);
nand U6151 (N_6151,N_5678,N_5960);
and U6152 (N_6152,N_5105,N_5554);
xor U6153 (N_6153,N_5703,N_5314);
nor U6154 (N_6154,N_5425,N_5011);
nand U6155 (N_6155,N_5419,N_5223);
and U6156 (N_6156,N_5683,N_5659);
or U6157 (N_6157,N_5828,N_5679);
nor U6158 (N_6158,N_5749,N_5128);
and U6159 (N_6159,N_5096,N_5479);
or U6160 (N_6160,N_5053,N_5169);
xnor U6161 (N_6161,N_5240,N_5401);
nor U6162 (N_6162,N_5502,N_5966);
or U6163 (N_6163,N_5665,N_5394);
xnor U6164 (N_6164,N_5000,N_5269);
xnor U6165 (N_6165,N_5747,N_5725);
and U6166 (N_6166,N_5079,N_5104);
and U6167 (N_6167,N_5266,N_5402);
xnor U6168 (N_6168,N_5389,N_5301);
or U6169 (N_6169,N_5792,N_5309);
and U6170 (N_6170,N_5037,N_5140);
xnor U6171 (N_6171,N_5198,N_5229);
nand U6172 (N_6172,N_5119,N_5340);
xor U6173 (N_6173,N_5606,N_5195);
xor U6174 (N_6174,N_5433,N_5629);
and U6175 (N_6175,N_5686,N_5356);
nand U6176 (N_6176,N_5867,N_5516);
nand U6177 (N_6177,N_5741,N_5411);
xnor U6178 (N_6178,N_5996,N_5545);
nand U6179 (N_6179,N_5815,N_5213);
and U6180 (N_6180,N_5709,N_5228);
and U6181 (N_6181,N_5783,N_5517);
and U6182 (N_6182,N_5247,N_5527);
or U6183 (N_6183,N_5136,N_5480);
xor U6184 (N_6184,N_5363,N_5501);
xnor U6185 (N_6185,N_5945,N_5491);
xnor U6186 (N_6186,N_5761,N_5623);
nor U6187 (N_6187,N_5965,N_5084);
xnor U6188 (N_6188,N_5268,N_5496);
nand U6189 (N_6189,N_5890,N_5611);
nand U6190 (N_6190,N_5369,N_5049);
xor U6191 (N_6191,N_5993,N_5121);
nor U6192 (N_6192,N_5615,N_5880);
and U6193 (N_6193,N_5775,N_5299);
nand U6194 (N_6194,N_5727,N_5066);
and U6195 (N_6195,N_5055,N_5591);
nor U6196 (N_6196,N_5904,N_5331);
or U6197 (N_6197,N_5655,N_5438);
and U6198 (N_6198,N_5574,N_5280);
and U6199 (N_6199,N_5733,N_5658);
xnor U6200 (N_6200,N_5069,N_5180);
or U6201 (N_6201,N_5769,N_5711);
and U6202 (N_6202,N_5829,N_5952);
nand U6203 (N_6203,N_5062,N_5454);
xor U6204 (N_6204,N_5046,N_5232);
xor U6205 (N_6205,N_5843,N_5714);
nand U6206 (N_6206,N_5273,N_5844);
nand U6207 (N_6207,N_5509,N_5386);
and U6208 (N_6208,N_5745,N_5444);
nor U6209 (N_6209,N_5510,N_5652);
and U6210 (N_6210,N_5406,N_5482);
nor U6211 (N_6211,N_5399,N_5925);
and U6212 (N_6212,N_5190,N_5712);
and U6213 (N_6213,N_5962,N_5970);
nand U6214 (N_6214,N_5565,N_5918);
or U6215 (N_6215,N_5405,N_5333);
nand U6216 (N_6216,N_5146,N_5110);
xnor U6217 (N_6217,N_5908,N_5858);
and U6218 (N_6218,N_5864,N_5589);
nor U6219 (N_6219,N_5941,N_5380);
nand U6220 (N_6220,N_5519,N_5224);
nand U6221 (N_6221,N_5854,N_5842);
xor U6222 (N_6222,N_5730,N_5289);
nand U6223 (N_6223,N_5663,N_5924);
nand U6224 (N_6224,N_5560,N_5732);
or U6225 (N_6225,N_5631,N_5464);
nor U6226 (N_6226,N_5226,N_5532);
nand U6227 (N_6227,N_5801,N_5217);
xnor U6228 (N_6228,N_5855,N_5827);
or U6229 (N_6229,N_5173,N_5025);
and U6230 (N_6230,N_5886,N_5499);
and U6231 (N_6231,N_5127,N_5929);
or U6232 (N_6232,N_5736,N_5558);
xor U6233 (N_6233,N_5328,N_5410);
xor U6234 (N_6234,N_5135,N_5423);
and U6235 (N_6235,N_5485,N_5350);
or U6236 (N_6236,N_5786,N_5327);
or U6237 (N_6237,N_5246,N_5535);
and U6238 (N_6238,N_5798,N_5851);
xnor U6239 (N_6239,N_5573,N_5696);
nor U6240 (N_6240,N_5746,N_5595);
and U6241 (N_6241,N_5193,N_5974);
or U6242 (N_6242,N_5088,N_5920);
nor U6243 (N_6243,N_5015,N_5058);
xor U6244 (N_6244,N_5857,N_5992);
xnor U6245 (N_6245,N_5129,N_5098);
xnor U6246 (N_6246,N_5796,N_5103);
and U6247 (N_6247,N_5818,N_5466);
nand U6248 (N_6248,N_5566,N_5461);
xor U6249 (N_6249,N_5494,N_5375);
and U6250 (N_6250,N_5398,N_5206);
xnor U6251 (N_6251,N_5503,N_5530);
and U6252 (N_6252,N_5422,N_5593);
and U6253 (N_6253,N_5654,N_5790);
or U6254 (N_6254,N_5557,N_5977);
nor U6255 (N_6255,N_5515,N_5203);
nor U6256 (N_6256,N_5522,N_5997);
nor U6257 (N_6257,N_5414,N_5462);
or U6258 (N_6258,N_5763,N_5003);
and U6259 (N_6259,N_5889,N_5144);
nor U6260 (N_6260,N_5787,N_5163);
nor U6261 (N_6261,N_5585,N_5635);
nor U6262 (N_6262,N_5027,N_5077);
nand U6263 (N_6263,N_5265,N_5800);
xor U6264 (N_6264,N_5587,N_5167);
and U6265 (N_6265,N_5234,N_5755);
or U6266 (N_6266,N_5445,N_5544);
or U6267 (N_6267,N_5849,N_5385);
xnor U6268 (N_6268,N_5233,N_5690);
nand U6269 (N_6269,N_5191,N_5697);
and U6270 (N_6270,N_5825,N_5236);
nor U6271 (N_6271,N_5021,N_5421);
xor U6272 (N_6272,N_5548,N_5513);
or U6273 (N_6273,N_5717,N_5869);
nor U6274 (N_6274,N_5588,N_5878);
xor U6275 (N_6275,N_5757,N_5330);
or U6276 (N_6276,N_5944,N_5954);
nand U6277 (N_6277,N_5312,N_5253);
nand U6278 (N_6278,N_5586,N_5298);
nand U6279 (N_6279,N_5978,N_5803);
or U6280 (N_6280,N_5337,N_5160);
xnor U6281 (N_6281,N_5097,N_5042);
or U6282 (N_6282,N_5295,N_5379);
or U6283 (N_6283,N_5765,N_5795);
xor U6284 (N_6284,N_5400,N_5117);
or U6285 (N_6285,N_5041,N_5907);
nand U6286 (N_6286,N_5044,N_5056);
or U6287 (N_6287,N_5336,N_5351);
nor U6288 (N_6288,N_5677,N_5626);
nand U6289 (N_6289,N_5750,N_5898);
nor U6290 (N_6290,N_5486,N_5939);
xor U6291 (N_6291,N_5614,N_5321);
and U6292 (N_6292,N_5427,N_5114);
xnor U6293 (N_6293,N_5779,N_5432);
nor U6294 (N_6294,N_5215,N_5577);
nand U6295 (N_6295,N_5107,N_5906);
nand U6296 (N_6296,N_5133,N_5305);
and U6297 (N_6297,N_5640,N_5660);
nand U6298 (N_6298,N_5450,N_5946);
or U6299 (N_6299,N_5238,N_5742);
or U6300 (N_6300,N_5949,N_5692);
or U6301 (N_6301,N_5495,N_5816);
nor U6302 (N_6302,N_5390,N_5726);
nor U6303 (N_6303,N_5032,N_5579);
nor U6304 (N_6304,N_5302,N_5705);
and U6305 (N_6305,N_5483,N_5376);
nor U6306 (N_6306,N_5346,N_5708);
or U6307 (N_6307,N_5208,N_5823);
or U6308 (N_6308,N_5040,N_5052);
and U6309 (N_6309,N_5286,N_5178);
and U6310 (N_6310,N_5418,N_5492);
nor U6311 (N_6311,N_5204,N_5192);
nand U6312 (N_6312,N_5602,N_5838);
or U6313 (N_6313,N_5860,N_5326);
and U6314 (N_6314,N_5737,N_5313);
xnor U6315 (N_6315,N_5430,N_5241);
and U6316 (N_6316,N_5443,N_5424);
nand U6317 (N_6317,N_5218,N_5367);
nor U6318 (N_6318,N_5624,N_5381);
nor U6319 (N_6319,N_5734,N_5921);
xnor U6320 (N_6320,N_5634,N_5580);
or U6321 (N_6321,N_5447,N_5718);
and U6322 (N_6322,N_5074,N_5434);
nand U6323 (N_6323,N_5781,N_5050);
and U6324 (N_6324,N_5500,N_5171);
and U6325 (N_6325,N_5091,N_5200);
and U6326 (N_6326,N_5393,N_5045);
or U6327 (N_6327,N_5836,N_5933);
nor U6328 (N_6328,N_5006,N_5553);
nand U6329 (N_6329,N_5029,N_5995);
nor U6330 (N_6330,N_5682,N_5603);
nor U6331 (N_6331,N_5758,N_5927);
nand U6332 (N_6332,N_5989,N_5891);
or U6333 (N_6333,N_5839,N_5339);
nor U6334 (N_6334,N_5150,N_5784);
or U6335 (N_6335,N_5397,N_5541);
and U6336 (N_6336,N_5151,N_5512);
or U6337 (N_6337,N_5582,N_5368);
nor U6338 (N_6338,N_5721,N_5599);
and U6339 (N_6339,N_5537,N_5352);
nand U6340 (N_6340,N_5209,N_5644);
xnor U6341 (N_6341,N_5227,N_5806);
and U6342 (N_6342,N_5979,N_5057);
and U6343 (N_6343,N_5478,N_5362);
nor U6344 (N_6344,N_5903,N_5360);
xnor U6345 (N_6345,N_5263,N_5242);
and U6346 (N_6346,N_5235,N_5853);
or U6347 (N_6347,N_5910,N_5617);
or U6348 (N_6348,N_5564,N_5555);
and U6349 (N_6349,N_5138,N_5578);
or U6350 (N_6350,N_5862,N_5969);
xor U6351 (N_6351,N_5028,N_5431);
or U6352 (N_6352,N_5604,N_5830);
nor U6353 (N_6353,N_5222,N_5323);
nor U6354 (N_6354,N_5752,N_5928);
xor U6355 (N_6355,N_5633,N_5275);
nor U6356 (N_6356,N_5377,N_5953);
or U6357 (N_6357,N_5646,N_5852);
xor U6358 (N_6358,N_5518,N_5575);
xor U6359 (N_6359,N_5020,N_5793);
xor U6360 (N_6360,N_5259,N_5442);
nand U6361 (N_6361,N_5956,N_5412);
xor U6362 (N_6362,N_5183,N_5063);
and U6363 (N_6363,N_5254,N_5141);
or U6364 (N_6364,N_5866,N_5072);
nor U6365 (N_6365,N_5184,N_5332);
nor U6366 (N_6366,N_5493,N_5470);
and U6367 (N_6367,N_5005,N_5174);
nor U6368 (N_6368,N_5976,N_5987);
xnor U6369 (N_6369,N_5214,N_5341);
nand U6370 (N_6370,N_5724,N_5065);
nand U6371 (N_6371,N_5601,N_5112);
xnor U6372 (N_6372,N_5552,N_5396);
xnor U6373 (N_6373,N_5715,N_5212);
and U6374 (N_6374,N_5832,N_5008);
xnor U6375 (N_6375,N_5297,N_5311);
and U6376 (N_6376,N_5756,N_5870);
and U6377 (N_6377,N_5650,N_5936);
nor U6378 (N_6378,N_5199,N_5142);
xnor U6379 (N_6379,N_5456,N_5605);
nand U6380 (N_6380,N_5279,N_5562);
nor U6381 (N_6381,N_5613,N_5282);
nor U6382 (N_6382,N_5007,N_5873);
nand U6383 (N_6383,N_5082,N_5720);
or U6384 (N_6384,N_5471,N_5017);
nor U6385 (N_6385,N_5556,N_5249);
xor U6386 (N_6386,N_5531,N_5674);
nand U6387 (N_6387,N_5460,N_5294);
and U6388 (N_6388,N_5740,N_5642);
xnor U6389 (N_6389,N_5437,N_5474);
or U6390 (N_6390,N_5619,N_5439);
and U6391 (N_6391,N_5523,N_5080);
nor U6392 (N_6392,N_5395,N_5872);
nor U6393 (N_6393,N_5991,N_5797);
nand U6394 (N_6394,N_5078,N_5022);
or U6395 (N_6395,N_5267,N_5657);
or U6396 (N_6396,N_5985,N_5426);
nand U6397 (N_6397,N_5272,N_5893);
or U6398 (N_6398,N_5081,N_5252);
xnor U6399 (N_6399,N_5384,N_5303);
nand U6400 (N_6400,N_5463,N_5067);
nor U6401 (N_6401,N_5540,N_5089);
and U6402 (N_6402,N_5221,N_5387);
nor U6403 (N_6403,N_5699,N_5219);
xnor U6404 (N_6404,N_5568,N_5016);
nand U6405 (N_6405,N_5570,N_5620);
nor U6406 (N_6406,N_5113,N_5778);
nand U6407 (N_6407,N_5955,N_5534);
nand U6408 (N_6408,N_5689,N_5258);
or U6409 (N_6409,N_5361,N_5846);
and U6410 (N_6410,N_5590,N_5452);
or U6411 (N_6411,N_5762,N_5043);
or U6412 (N_6412,N_5093,N_5639);
nand U6413 (N_6413,N_5968,N_5172);
or U6414 (N_6414,N_5896,N_5782);
xnor U6415 (N_6415,N_5538,N_5529);
xor U6416 (N_6416,N_5475,N_5704);
nand U6417 (N_6417,N_5001,N_5251);
nand U6418 (N_6418,N_5420,N_5947);
or U6419 (N_6419,N_5498,N_5137);
nor U6420 (N_6420,N_5681,N_5719);
xnor U6421 (N_6421,N_5320,N_5628);
nand U6422 (N_6422,N_5364,N_5597);
and U6423 (N_6423,N_5693,N_5116);
nor U6424 (N_6424,N_5571,N_5743);
or U6425 (N_6425,N_5338,N_5789);
or U6426 (N_6426,N_5102,N_5068);
nor U6427 (N_6427,N_5153,N_5147);
and U6428 (N_6428,N_5469,N_5342);
nor U6429 (N_6429,N_5250,N_5018);
and U6430 (N_6430,N_5448,N_5988);
xor U6431 (N_6431,N_5850,N_5567);
xnor U6432 (N_6432,N_5824,N_5156);
nor U6433 (N_6433,N_5666,N_5539);
and U6434 (N_6434,N_5285,N_5100);
xor U6435 (N_6435,N_5805,N_5086);
nand U6436 (N_6436,N_5449,N_5009);
nand U6437 (N_6437,N_5772,N_5413);
nor U6438 (N_6438,N_5581,N_5819);
or U6439 (N_6439,N_5391,N_5609);
nor U6440 (N_6440,N_5278,N_5622);
or U6441 (N_6441,N_5429,N_5417);
and U6442 (N_6442,N_5672,N_5649);
xnor U6443 (N_6443,N_5125,N_5095);
xnor U6444 (N_6444,N_5729,N_5457);
or U6445 (N_6445,N_5973,N_5287);
nor U6446 (N_6446,N_5181,N_5598);
or U6447 (N_6447,N_5592,N_5950);
and U6448 (N_6448,N_5261,N_5909);
nand U6449 (N_6449,N_5959,N_5958);
xor U6450 (N_6450,N_5061,N_5168);
nor U6451 (N_6451,N_5882,N_5131);
nor U6452 (N_6452,N_5702,N_5900);
or U6453 (N_6453,N_5126,N_5165);
xnor U6454 (N_6454,N_5826,N_5365);
nand U6455 (N_6455,N_5416,N_5348);
and U6456 (N_6456,N_5600,N_5073);
or U6457 (N_6457,N_5675,N_5196);
nor U6458 (N_6458,N_5561,N_5308);
and U6459 (N_6459,N_5216,N_5157);
nor U6460 (N_6460,N_5205,N_5115);
nor U6461 (N_6461,N_5731,N_5315);
or U6462 (N_6462,N_5106,N_5476);
or U6463 (N_6463,N_5688,N_5325);
and U6464 (N_6464,N_5768,N_5382);
nand U6465 (N_6465,N_5651,N_5938);
nand U6466 (N_6466,N_5668,N_5542);
and U6467 (N_6467,N_5211,N_5143);
or U6468 (N_6468,N_5154,N_5759);
nand U6469 (N_6469,N_5738,N_5641);
nand U6470 (N_6470,N_5684,N_5237);
or U6471 (N_6471,N_5435,N_5680);
or U6472 (N_6472,N_5911,N_5322);
xnor U6473 (N_6473,N_5999,N_5409);
and U6474 (N_6474,N_5404,N_5441);
and U6475 (N_6475,N_5186,N_5559);
or U6476 (N_6476,N_5371,N_5488);
or U6477 (N_6477,N_5943,N_5415);
nand U6478 (N_6478,N_5788,N_5594);
nor U6479 (N_6479,N_5051,N_5316);
or U6480 (N_6480,N_5935,N_5508);
xnor U6481 (N_6481,N_5964,N_5383);
and U6482 (N_6482,N_5004,N_5848);
nor U6483 (N_6483,N_5060,N_5648);
nor U6484 (N_6484,N_5359,N_5239);
nor U6485 (N_6485,N_5856,N_5902);
nor U6486 (N_6486,N_5132,N_5710);
xnor U6487 (N_6487,N_5317,N_5152);
or U6488 (N_6488,N_5188,N_5197);
nor U6489 (N_6489,N_5608,N_5472);
and U6490 (N_6490,N_5264,N_5821);
nor U6491 (N_6491,N_5373,N_5408);
and U6492 (N_6492,N_5653,N_5319);
and U6493 (N_6493,N_5459,N_5748);
nor U6494 (N_6494,N_5751,N_5643);
or U6495 (N_6495,N_5972,N_5446);
nor U6496 (N_6496,N_5983,N_5894);
nand U6497 (N_6497,N_5645,N_5284);
nand U6498 (N_6498,N_5033,N_5569);
and U6499 (N_6499,N_5892,N_5543);
xnor U6500 (N_6500,N_5611,N_5658);
and U6501 (N_6501,N_5704,N_5724);
and U6502 (N_6502,N_5708,N_5074);
xnor U6503 (N_6503,N_5820,N_5905);
or U6504 (N_6504,N_5967,N_5248);
and U6505 (N_6505,N_5738,N_5834);
and U6506 (N_6506,N_5757,N_5872);
or U6507 (N_6507,N_5803,N_5310);
xnor U6508 (N_6508,N_5543,N_5623);
and U6509 (N_6509,N_5256,N_5906);
nor U6510 (N_6510,N_5087,N_5254);
or U6511 (N_6511,N_5659,N_5158);
or U6512 (N_6512,N_5468,N_5623);
and U6513 (N_6513,N_5410,N_5693);
nor U6514 (N_6514,N_5075,N_5281);
nor U6515 (N_6515,N_5109,N_5199);
nand U6516 (N_6516,N_5060,N_5123);
or U6517 (N_6517,N_5312,N_5895);
or U6518 (N_6518,N_5981,N_5341);
and U6519 (N_6519,N_5366,N_5730);
nand U6520 (N_6520,N_5829,N_5977);
or U6521 (N_6521,N_5686,N_5635);
xor U6522 (N_6522,N_5599,N_5971);
or U6523 (N_6523,N_5929,N_5588);
and U6524 (N_6524,N_5268,N_5980);
xnor U6525 (N_6525,N_5755,N_5473);
nor U6526 (N_6526,N_5094,N_5784);
and U6527 (N_6527,N_5940,N_5062);
or U6528 (N_6528,N_5227,N_5039);
or U6529 (N_6529,N_5858,N_5736);
or U6530 (N_6530,N_5555,N_5096);
or U6531 (N_6531,N_5306,N_5446);
nand U6532 (N_6532,N_5165,N_5946);
or U6533 (N_6533,N_5760,N_5725);
nor U6534 (N_6534,N_5822,N_5552);
or U6535 (N_6535,N_5083,N_5422);
nor U6536 (N_6536,N_5277,N_5170);
nor U6537 (N_6537,N_5864,N_5124);
nor U6538 (N_6538,N_5953,N_5040);
nand U6539 (N_6539,N_5302,N_5915);
and U6540 (N_6540,N_5555,N_5461);
nand U6541 (N_6541,N_5706,N_5838);
nand U6542 (N_6542,N_5716,N_5956);
nor U6543 (N_6543,N_5028,N_5785);
nand U6544 (N_6544,N_5617,N_5122);
nor U6545 (N_6545,N_5997,N_5337);
and U6546 (N_6546,N_5211,N_5214);
xor U6547 (N_6547,N_5797,N_5597);
or U6548 (N_6548,N_5395,N_5280);
and U6549 (N_6549,N_5770,N_5889);
nand U6550 (N_6550,N_5077,N_5061);
or U6551 (N_6551,N_5345,N_5154);
xor U6552 (N_6552,N_5292,N_5012);
nand U6553 (N_6553,N_5858,N_5778);
or U6554 (N_6554,N_5123,N_5473);
nand U6555 (N_6555,N_5836,N_5403);
nand U6556 (N_6556,N_5564,N_5511);
xnor U6557 (N_6557,N_5275,N_5007);
or U6558 (N_6558,N_5535,N_5013);
xnor U6559 (N_6559,N_5289,N_5335);
nand U6560 (N_6560,N_5859,N_5354);
nand U6561 (N_6561,N_5631,N_5341);
nor U6562 (N_6562,N_5778,N_5783);
xnor U6563 (N_6563,N_5325,N_5447);
nor U6564 (N_6564,N_5118,N_5572);
or U6565 (N_6565,N_5468,N_5672);
or U6566 (N_6566,N_5473,N_5994);
and U6567 (N_6567,N_5710,N_5608);
xor U6568 (N_6568,N_5802,N_5382);
and U6569 (N_6569,N_5440,N_5405);
xnor U6570 (N_6570,N_5730,N_5501);
or U6571 (N_6571,N_5955,N_5414);
nor U6572 (N_6572,N_5468,N_5927);
nor U6573 (N_6573,N_5398,N_5999);
xnor U6574 (N_6574,N_5659,N_5569);
nor U6575 (N_6575,N_5576,N_5645);
and U6576 (N_6576,N_5083,N_5596);
nor U6577 (N_6577,N_5489,N_5206);
xnor U6578 (N_6578,N_5705,N_5965);
nand U6579 (N_6579,N_5851,N_5343);
nor U6580 (N_6580,N_5112,N_5252);
xnor U6581 (N_6581,N_5722,N_5965);
and U6582 (N_6582,N_5352,N_5223);
nand U6583 (N_6583,N_5216,N_5899);
xor U6584 (N_6584,N_5372,N_5641);
and U6585 (N_6585,N_5460,N_5928);
nor U6586 (N_6586,N_5127,N_5680);
and U6587 (N_6587,N_5508,N_5007);
nor U6588 (N_6588,N_5152,N_5761);
nand U6589 (N_6589,N_5840,N_5784);
or U6590 (N_6590,N_5136,N_5573);
xor U6591 (N_6591,N_5331,N_5965);
nand U6592 (N_6592,N_5726,N_5324);
or U6593 (N_6593,N_5679,N_5144);
xnor U6594 (N_6594,N_5339,N_5303);
xor U6595 (N_6595,N_5115,N_5128);
or U6596 (N_6596,N_5534,N_5444);
nand U6597 (N_6597,N_5876,N_5912);
xnor U6598 (N_6598,N_5196,N_5752);
or U6599 (N_6599,N_5954,N_5106);
nor U6600 (N_6600,N_5693,N_5090);
nand U6601 (N_6601,N_5788,N_5833);
or U6602 (N_6602,N_5960,N_5614);
and U6603 (N_6603,N_5588,N_5787);
xor U6604 (N_6604,N_5718,N_5670);
or U6605 (N_6605,N_5826,N_5236);
xor U6606 (N_6606,N_5764,N_5367);
and U6607 (N_6607,N_5530,N_5894);
nand U6608 (N_6608,N_5655,N_5723);
and U6609 (N_6609,N_5804,N_5517);
nor U6610 (N_6610,N_5811,N_5560);
nor U6611 (N_6611,N_5880,N_5696);
nor U6612 (N_6612,N_5228,N_5630);
and U6613 (N_6613,N_5548,N_5815);
xnor U6614 (N_6614,N_5704,N_5892);
nand U6615 (N_6615,N_5617,N_5205);
and U6616 (N_6616,N_5937,N_5381);
or U6617 (N_6617,N_5892,N_5410);
or U6618 (N_6618,N_5219,N_5243);
xor U6619 (N_6619,N_5888,N_5108);
xnor U6620 (N_6620,N_5798,N_5452);
nor U6621 (N_6621,N_5724,N_5145);
and U6622 (N_6622,N_5799,N_5875);
nor U6623 (N_6623,N_5067,N_5241);
nor U6624 (N_6624,N_5107,N_5838);
xnor U6625 (N_6625,N_5049,N_5634);
nand U6626 (N_6626,N_5079,N_5754);
nand U6627 (N_6627,N_5240,N_5927);
nand U6628 (N_6628,N_5066,N_5951);
and U6629 (N_6629,N_5585,N_5528);
xnor U6630 (N_6630,N_5270,N_5142);
and U6631 (N_6631,N_5086,N_5328);
or U6632 (N_6632,N_5830,N_5726);
and U6633 (N_6633,N_5149,N_5653);
nor U6634 (N_6634,N_5744,N_5804);
xnor U6635 (N_6635,N_5997,N_5841);
or U6636 (N_6636,N_5550,N_5456);
xnor U6637 (N_6637,N_5000,N_5225);
xor U6638 (N_6638,N_5737,N_5923);
nor U6639 (N_6639,N_5637,N_5243);
or U6640 (N_6640,N_5956,N_5910);
nand U6641 (N_6641,N_5814,N_5343);
nand U6642 (N_6642,N_5726,N_5808);
or U6643 (N_6643,N_5295,N_5885);
xor U6644 (N_6644,N_5984,N_5460);
or U6645 (N_6645,N_5578,N_5694);
and U6646 (N_6646,N_5772,N_5359);
nor U6647 (N_6647,N_5250,N_5193);
xor U6648 (N_6648,N_5891,N_5717);
nor U6649 (N_6649,N_5367,N_5721);
nor U6650 (N_6650,N_5071,N_5656);
nor U6651 (N_6651,N_5801,N_5623);
nor U6652 (N_6652,N_5975,N_5690);
nor U6653 (N_6653,N_5056,N_5502);
or U6654 (N_6654,N_5900,N_5534);
nand U6655 (N_6655,N_5903,N_5320);
nor U6656 (N_6656,N_5508,N_5549);
xor U6657 (N_6657,N_5283,N_5169);
nand U6658 (N_6658,N_5988,N_5042);
or U6659 (N_6659,N_5643,N_5821);
nor U6660 (N_6660,N_5131,N_5831);
nand U6661 (N_6661,N_5099,N_5124);
nor U6662 (N_6662,N_5210,N_5345);
nand U6663 (N_6663,N_5089,N_5098);
xor U6664 (N_6664,N_5757,N_5302);
or U6665 (N_6665,N_5896,N_5841);
nand U6666 (N_6666,N_5865,N_5701);
nand U6667 (N_6667,N_5547,N_5596);
nand U6668 (N_6668,N_5193,N_5388);
xor U6669 (N_6669,N_5654,N_5980);
nand U6670 (N_6670,N_5413,N_5844);
and U6671 (N_6671,N_5112,N_5525);
xnor U6672 (N_6672,N_5841,N_5732);
nand U6673 (N_6673,N_5800,N_5601);
nor U6674 (N_6674,N_5378,N_5171);
or U6675 (N_6675,N_5141,N_5641);
xnor U6676 (N_6676,N_5160,N_5840);
xor U6677 (N_6677,N_5660,N_5646);
xnor U6678 (N_6678,N_5851,N_5996);
nand U6679 (N_6679,N_5080,N_5476);
nor U6680 (N_6680,N_5902,N_5429);
nand U6681 (N_6681,N_5258,N_5502);
or U6682 (N_6682,N_5962,N_5081);
or U6683 (N_6683,N_5229,N_5725);
nor U6684 (N_6684,N_5595,N_5100);
or U6685 (N_6685,N_5899,N_5942);
nand U6686 (N_6686,N_5182,N_5023);
and U6687 (N_6687,N_5207,N_5133);
xnor U6688 (N_6688,N_5431,N_5925);
or U6689 (N_6689,N_5025,N_5019);
or U6690 (N_6690,N_5680,N_5965);
or U6691 (N_6691,N_5175,N_5756);
or U6692 (N_6692,N_5685,N_5673);
and U6693 (N_6693,N_5990,N_5045);
nor U6694 (N_6694,N_5613,N_5255);
or U6695 (N_6695,N_5920,N_5041);
nand U6696 (N_6696,N_5040,N_5354);
nor U6697 (N_6697,N_5325,N_5940);
nor U6698 (N_6698,N_5895,N_5770);
or U6699 (N_6699,N_5015,N_5240);
or U6700 (N_6700,N_5118,N_5848);
and U6701 (N_6701,N_5647,N_5062);
xnor U6702 (N_6702,N_5542,N_5353);
and U6703 (N_6703,N_5654,N_5631);
and U6704 (N_6704,N_5020,N_5346);
and U6705 (N_6705,N_5361,N_5544);
nor U6706 (N_6706,N_5914,N_5245);
xnor U6707 (N_6707,N_5350,N_5102);
nor U6708 (N_6708,N_5019,N_5884);
or U6709 (N_6709,N_5474,N_5941);
or U6710 (N_6710,N_5200,N_5913);
nor U6711 (N_6711,N_5298,N_5303);
and U6712 (N_6712,N_5780,N_5821);
nor U6713 (N_6713,N_5024,N_5084);
or U6714 (N_6714,N_5379,N_5885);
or U6715 (N_6715,N_5638,N_5274);
xor U6716 (N_6716,N_5899,N_5853);
xor U6717 (N_6717,N_5916,N_5517);
or U6718 (N_6718,N_5314,N_5054);
nand U6719 (N_6719,N_5201,N_5303);
xor U6720 (N_6720,N_5216,N_5574);
nor U6721 (N_6721,N_5964,N_5184);
and U6722 (N_6722,N_5392,N_5225);
nand U6723 (N_6723,N_5268,N_5866);
nand U6724 (N_6724,N_5953,N_5193);
and U6725 (N_6725,N_5006,N_5925);
and U6726 (N_6726,N_5566,N_5788);
xnor U6727 (N_6727,N_5652,N_5982);
or U6728 (N_6728,N_5380,N_5706);
xor U6729 (N_6729,N_5512,N_5344);
or U6730 (N_6730,N_5163,N_5599);
or U6731 (N_6731,N_5462,N_5598);
or U6732 (N_6732,N_5685,N_5934);
nor U6733 (N_6733,N_5319,N_5689);
or U6734 (N_6734,N_5057,N_5082);
or U6735 (N_6735,N_5762,N_5354);
xnor U6736 (N_6736,N_5968,N_5351);
and U6737 (N_6737,N_5975,N_5737);
xor U6738 (N_6738,N_5338,N_5971);
xor U6739 (N_6739,N_5405,N_5698);
or U6740 (N_6740,N_5360,N_5480);
or U6741 (N_6741,N_5307,N_5544);
or U6742 (N_6742,N_5627,N_5454);
nor U6743 (N_6743,N_5613,N_5572);
nand U6744 (N_6744,N_5084,N_5863);
nor U6745 (N_6745,N_5604,N_5857);
and U6746 (N_6746,N_5588,N_5185);
and U6747 (N_6747,N_5080,N_5195);
xor U6748 (N_6748,N_5224,N_5991);
xnor U6749 (N_6749,N_5517,N_5682);
or U6750 (N_6750,N_5775,N_5414);
or U6751 (N_6751,N_5298,N_5949);
or U6752 (N_6752,N_5688,N_5982);
nand U6753 (N_6753,N_5853,N_5125);
xor U6754 (N_6754,N_5694,N_5303);
or U6755 (N_6755,N_5441,N_5913);
and U6756 (N_6756,N_5566,N_5798);
and U6757 (N_6757,N_5371,N_5625);
nor U6758 (N_6758,N_5153,N_5716);
or U6759 (N_6759,N_5669,N_5465);
xnor U6760 (N_6760,N_5066,N_5335);
nand U6761 (N_6761,N_5923,N_5160);
and U6762 (N_6762,N_5234,N_5583);
or U6763 (N_6763,N_5433,N_5738);
nor U6764 (N_6764,N_5725,N_5399);
nand U6765 (N_6765,N_5398,N_5605);
and U6766 (N_6766,N_5191,N_5961);
or U6767 (N_6767,N_5573,N_5087);
or U6768 (N_6768,N_5769,N_5780);
nor U6769 (N_6769,N_5165,N_5916);
nand U6770 (N_6770,N_5967,N_5256);
and U6771 (N_6771,N_5913,N_5899);
nor U6772 (N_6772,N_5156,N_5874);
xor U6773 (N_6773,N_5567,N_5004);
and U6774 (N_6774,N_5022,N_5062);
and U6775 (N_6775,N_5034,N_5985);
or U6776 (N_6776,N_5234,N_5719);
nand U6777 (N_6777,N_5148,N_5627);
xor U6778 (N_6778,N_5970,N_5771);
xor U6779 (N_6779,N_5451,N_5570);
xor U6780 (N_6780,N_5654,N_5607);
nand U6781 (N_6781,N_5735,N_5633);
nor U6782 (N_6782,N_5820,N_5720);
and U6783 (N_6783,N_5628,N_5079);
nor U6784 (N_6784,N_5810,N_5713);
and U6785 (N_6785,N_5641,N_5103);
and U6786 (N_6786,N_5932,N_5829);
nor U6787 (N_6787,N_5109,N_5665);
or U6788 (N_6788,N_5534,N_5266);
nor U6789 (N_6789,N_5318,N_5045);
nor U6790 (N_6790,N_5007,N_5299);
nand U6791 (N_6791,N_5407,N_5531);
or U6792 (N_6792,N_5890,N_5080);
or U6793 (N_6793,N_5922,N_5869);
and U6794 (N_6794,N_5602,N_5025);
or U6795 (N_6795,N_5729,N_5532);
or U6796 (N_6796,N_5009,N_5379);
and U6797 (N_6797,N_5352,N_5951);
and U6798 (N_6798,N_5195,N_5197);
nand U6799 (N_6799,N_5900,N_5646);
and U6800 (N_6800,N_5794,N_5914);
nand U6801 (N_6801,N_5661,N_5677);
nand U6802 (N_6802,N_5483,N_5768);
and U6803 (N_6803,N_5602,N_5621);
nor U6804 (N_6804,N_5005,N_5419);
or U6805 (N_6805,N_5949,N_5290);
or U6806 (N_6806,N_5797,N_5888);
or U6807 (N_6807,N_5919,N_5101);
nor U6808 (N_6808,N_5948,N_5713);
nand U6809 (N_6809,N_5500,N_5145);
or U6810 (N_6810,N_5599,N_5458);
xnor U6811 (N_6811,N_5679,N_5550);
nand U6812 (N_6812,N_5817,N_5339);
or U6813 (N_6813,N_5333,N_5930);
xnor U6814 (N_6814,N_5476,N_5641);
xor U6815 (N_6815,N_5022,N_5701);
nor U6816 (N_6816,N_5036,N_5758);
xor U6817 (N_6817,N_5490,N_5626);
and U6818 (N_6818,N_5901,N_5971);
or U6819 (N_6819,N_5271,N_5024);
or U6820 (N_6820,N_5337,N_5183);
and U6821 (N_6821,N_5098,N_5586);
xnor U6822 (N_6822,N_5623,N_5532);
or U6823 (N_6823,N_5053,N_5366);
or U6824 (N_6824,N_5281,N_5386);
nor U6825 (N_6825,N_5706,N_5046);
xor U6826 (N_6826,N_5372,N_5534);
and U6827 (N_6827,N_5811,N_5220);
nand U6828 (N_6828,N_5863,N_5835);
nand U6829 (N_6829,N_5241,N_5591);
xor U6830 (N_6830,N_5783,N_5870);
nand U6831 (N_6831,N_5426,N_5369);
or U6832 (N_6832,N_5396,N_5687);
xor U6833 (N_6833,N_5883,N_5365);
or U6834 (N_6834,N_5328,N_5118);
xnor U6835 (N_6835,N_5149,N_5872);
and U6836 (N_6836,N_5061,N_5473);
or U6837 (N_6837,N_5193,N_5081);
or U6838 (N_6838,N_5337,N_5220);
or U6839 (N_6839,N_5211,N_5849);
xor U6840 (N_6840,N_5230,N_5851);
and U6841 (N_6841,N_5504,N_5458);
or U6842 (N_6842,N_5343,N_5623);
or U6843 (N_6843,N_5388,N_5084);
nor U6844 (N_6844,N_5021,N_5107);
nand U6845 (N_6845,N_5461,N_5086);
or U6846 (N_6846,N_5703,N_5583);
xnor U6847 (N_6847,N_5889,N_5417);
nand U6848 (N_6848,N_5081,N_5024);
nor U6849 (N_6849,N_5364,N_5107);
and U6850 (N_6850,N_5244,N_5966);
or U6851 (N_6851,N_5555,N_5496);
or U6852 (N_6852,N_5532,N_5275);
and U6853 (N_6853,N_5705,N_5042);
or U6854 (N_6854,N_5754,N_5111);
and U6855 (N_6855,N_5211,N_5369);
and U6856 (N_6856,N_5928,N_5465);
nor U6857 (N_6857,N_5008,N_5717);
nand U6858 (N_6858,N_5657,N_5322);
or U6859 (N_6859,N_5625,N_5627);
or U6860 (N_6860,N_5923,N_5462);
or U6861 (N_6861,N_5715,N_5072);
nand U6862 (N_6862,N_5244,N_5453);
nor U6863 (N_6863,N_5306,N_5932);
or U6864 (N_6864,N_5433,N_5573);
xor U6865 (N_6865,N_5309,N_5723);
xnor U6866 (N_6866,N_5655,N_5088);
or U6867 (N_6867,N_5309,N_5670);
nand U6868 (N_6868,N_5696,N_5052);
nor U6869 (N_6869,N_5227,N_5900);
nor U6870 (N_6870,N_5044,N_5628);
nor U6871 (N_6871,N_5835,N_5333);
xnor U6872 (N_6872,N_5051,N_5125);
nor U6873 (N_6873,N_5962,N_5384);
nor U6874 (N_6874,N_5426,N_5335);
or U6875 (N_6875,N_5597,N_5014);
and U6876 (N_6876,N_5672,N_5319);
nand U6877 (N_6877,N_5062,N_5389);
and U6878 (N_6878,N_5645,N_5635);
nand U6879 (N_6879,N_5925,N_5415);
xnor U6880 (N_6880,N_5744,N_5514);
nand U6881 (N_6881,N_5293,N_5455);
xnor U6882 (N_6882,N_5129,N_5584);
nand U6883 (N_6883,N_5826,N_5053);
nor U6884 (N_6884,N_5695,N_5552);
nand U6885 (N_6885,N_5033,N_5825);
nand U6886 (N_6886,N_5804,N_5952);
and U6887 (N_6887,N_5275,N_5946);
nand U6888 (N_6888,N_5531,N_5182);
or U6889 (N_6889,N_5715,N_5172);
or U6890 (N_6890,N_5229,N_5317);
xnor U6891 (N_6891,N_5206,N_5131);
nand U6892 (N_6892,N_5853,N_5942);
or U6893 (N_6893,N_5557,N_5669);
nand U6894 (N_6894,N_5325,N_5545);
and U6895 (N_6895,N_5112,N_5097);
or U6896 (N_6896,N_5652,N_5844);
or U6897 (N_6897,N_5949,N_5426);
nand U6898 (N_6898,N_5896,N_5915);
xnor U6899 (N_6899,N_5061,N_5370);
and U6900 (N_6900,N_5061,N_5971);
and U6901 (N_6901,N_5875,N_5064);
xnor U6902 (N_6902,N_5957,N_5440);
nor U6903 (N_6903,N_5576,N_5485);
xor U6904 (N_6904,N_5323,N_5117);
or U6905 (N_6905,N_5312,N_5257);
and U6906 (N_6906,N_5108,N_5441);
xor U6907 (N_6907,N_5411,N_5442);
and U6908 (N_6908,N_5157,N_5464);
and U6909 (N_6909,N_5155,N_5178);
xnor U6910 (N_6910,N_5860,N_5872);
nand U6911 (N_6911,N_5850,N_5772);
nand U6912 (N_6912,N_5303,N_5199);
nor U6913 (N_6913,N_5488,N_5463);
or U6914 (N_6914,N_5370,N_5634);
nor U6915 (N_6915,N_5713,N_5680);
or U6916 (N_6916,N_5047,N_5151);
nand U6917 (N_6917,N_5816,N_5428);
nand U6918 (N_6918,N_5642,N_5611);
nor U6919 (N_6919,N_5150,N_5999);
xnor U6920 (N_6920,N_5527,N_5689);
nand U6921 (N_6921,N_5993,N_5522);
nor U6922 (N_6922,N_5467,N_5919);
nand U6923 (N_6923,N_5339,N_5793);
or U6924 (N_6924,N_5912,N_5783);
nor U6925 (N_6925,N_5309,N_5020);
or U6926 (N_6926,N_5432,N_5324);
nand U6927 (N_6927,N_5196,N_5521);
xnor U6928 (N_6928,N_5068,N_5854);
nor U6929 (N_6929,N_5477,N_5745);
and U6930 (N_6930,N_5818,N_5031);
and U6931 (N_6931,N_5133,N_5468);
nand U6932 (N_6932,N_5778,N_5061);
xnor U6933 (N_6933,N_5694,N_5038);
or U6934 (N_6934,N_5915,N_5615);
and U6935 (N_6935,N_5294,N_5912);
or U6936 (N_6936,N_5602,N_5940);
or U6937 (N_6937,N_5308,N_5964);
or U6938 (N_6938,N_5013,N_5449);
xnor U6939 (N_6939,N_5780,N_5587);
nor U6940 (N_6940,N_5581,N_5790);
xnor U6941 (N_6941,N_5881,N_5559);
xnor U6942 (N_6942,N_5856,N_5206);
nor U6943 (N_6943,N_5629,N_5565);
nand U6944 (N_6944,N_5539,N_5063);
nor U6945 (N_6945,N_5216,N_5842);
xor U6946 (N_6946,N_5915,N_5708);
xor U6947 (N_6947,N_5360,N_5704);
nor U6948 (N_6948,N_5876,N_5656);
and U6949 (N_6949,N_5482,N_5962);
nand U6950 (N_6950,N_5359,N_5822);
or U6951 (N_6951,N_5564,N_5717);
nor U6952 (N_6952,N_5935,N_5015);
xor U6953 (N_6953,N_5377,N_5213);
and U6954 (N_6954,N_5447,N_5975);
nand U6955 (N_6955,N_5311,N_5993);
or U6956 (N_6956,N_5214,N_5926);
and U6957 (N_6957,N_5366,N_5921);
xor U6958 (N_6958,N_5349,N_5489);
nand U6959 (N_6959,N_5507,N_5180);
and U6960 (N_6960,N_5687,N_5217);
or U6961 (N_6961,N_5954,N_5785);
or U6962 (N_6962,N_5541,N_5848);
xor U6963 (N_6963,N_5838,N_5523);
and U6964 (N_6964,N_5150,N_5554);
nor U6965 (N_6965,N_5664,N_5763);
nor U6966 (N_6966,N_5140,N_5216);
xor U6967 (N_6967,N_5798,N_5772);
nand U6968 (N_6968,N_5884,N_5478);
and U6969 (N_6969,N_5032,N_5008);
xor U6970 (N_6970,N_5929,N_5435);
nand U6971 (N_6971,N_5013,N_5710);
nand U6972 (N_6972,N_5374,N_5573);
or U6973 (N_6973,N_5132,N_5946);
nor U6974 (N_6974,N_5905,N_5555);
and U6975 (N_6975,N_5803,N_5189);
and U6976 (N_6976,N_5783,N_5696);
and U6977 (N_6977,N_5004,N_5559);
nor U6978 (N_6978,N_5100,N_5857);
or U6979 (N_6979,N_5448,N_5737);
nand U6980 (N_6980,N_5097,N_5545);
nand U6981 (N_6981,N_5774,N_5714);
nor U6982 (N_6982,N_5418,N_5143);
xnor U6983 (N_6983,N_5319,N_5863);
and U6984 (N_6984,N_5529,N_5499);
and U6985 (N_6985,N_5483,N_5303);
xor U6986 (N_6986,N_5219,N_5164);
or U6987 (N_6987,N_5522,N_5023);
xnor U6988 (N_6988,N_5278,N_5495);
xor U6989 (N_6989,N_5124,N_5906);
nand U6990 (N_6990,N_5013,N_5060);
or U6991 (N_6991,N_5631,N_5579);
xor U6992 (N_6992,N_5591,N_5221);
and U6993 (N_6993,N_5552,N_5132);
or U6994 (N_6994,N_5712,N_5969);
nor U6995 (N_6995,N_5549,N_5364);
nor U6996 (N_6996,N_5767,N_5835);
xnor U6997 (N_6997,N_5543,N_5650);
nor U6998 (N_6998,N_5645,N_5806);
or U6999 (N_6999,N_5424,N_5975);
nor U7000 (N_7000,N_6734,N_6144);
nand U7001 (N_7001,N_6149,N_6169);
and U7002 (N_7002,N_6581,N_6195);
nor U7003 (N_7003,N_6354,N_6676);
nor U7004 (N_7004,N_6875,N_6163);
xnor U7005 (N_7005,N_6246,N_6740);
nand U7006 (N_7006,N_6468,N_6499);
xnor U7007 (N_7007,N_6827,N_6045);
and U7008 (N_7008,N_6721,N_6567);
nor U7009 (N_7009,N_6935,N_6200);
nand U7010 (N_7010,N_6292,N_6675);
or U7011 (N_7011,N_6456,N_6353);
or U7012 (N_7012,N_6392,N_6320);
and U7013 (N_7013,N_6670,N_6857);
nand U7014 (N_7014,N_6061,N_6267);
and U7015 (N_7015,N_6622,N_6752);
and U7016 (N_7016,N_6583,N_6132);
nand U7017 (N_7017,N_6239,N_6863);
xor U7018 (N_7018,N_6214,N_6650);
nor U7019 (N_7019,N_6559,N_6217);
or U7020 (N_7020,N_6786,N_6791);
nand U7021 (N_7021,N_6991,N_6665);
xor U7022 (N_7022,N_6357,N_6170);
nor U7023 (N_7023,N_6945,N_6871);
xor U7024 (N_7024,N_6589,N_6284);
or U7025 (N_7025,N_6100,N_6775);
nor U7026 (N_7026,N_6031,N_6923);
nand U7027 (N_7027,N_6962,N_6422);
nand U7028 (N_7028,N_6505,N_6606);
nand U7029 (N_7029,N_6829,N_6852);
nand U7030 (N_7030,N_6469,N_6027);
and U7031 (N_7031,N_6057,N_6433);
xor U7032 (N_7032,N_6797,N_6245);
nand U7033 (N_7033,N_6612,N_6271);
nand U7034 (N_7034,N_6849,N_6256);
or U7035 (N_7035,N_6288,N_6196);
nand U7036 (N_7036,N_6794,N_6951);
or U7037 (N_7037,N_6201,N_6632);
or U7038 (N_7038,N_6044,N_6616);
xnor U7039 (N_7039,N_6541,N_6578);
xnor U7040 (N_7040,N_6532,N_6087);
xnor U7041 (N_7041,N_6077,N_6492);
nor U7042 (N_7042,N_6990,N_6550);
nand U7043 (N_7043,N_6926,N_6148);
nor U7044 (N_7044,N_6980,N_6804);
or U7045 (N_7045,N_6411,N_6719);
and U7046 (N_7046,N_6753,N_6687);
nor U7047 (N_7047,N_6723,N_6707);
nor U7048 (N_7048,N_6537,N_6350);
nor U7049 (N_7049,N_6513,N_6437);
and U7050 (N_7050,N_6418,N_6240);
or U7051 (N_7051,N_6983,N_6273);
nand U7052 (N_7052,N_6324,N_6139);
nand U7053 (N_7053,N_6074,N_6472);
and U7054 (N_7054,N_6409,N_6093);
xnor U7055 (N_7055,N_6908,N_6933);
nand U7056 (N_7056,N_6640,N_6075);
xnor U7057 (N_7057,N_6654,N_6968);
nand U7058 (N_7058,N_6175,N_6495);
xnor U7059 (N_7059,N_6026,N_6296);
or U7060 (N_7060,N_6269,N_6035);
or U7061 (N_7061,N_6927,N_6759);
nand U7062 (N_7062,N_6958,N_6717);
nor U7063 (N_7063,N_6358,N_6218);
nor U7064 (N_7064,N_6588,N_6647);
xnor U7065 (N_7065,N_6549,N_6361);
nand U7066 (N_7066,N_6914,N_6446);
nor U7067 (N_7067,N_6376,N_6801);
or U7068 (N_7068,N_6192,N_6224);
and U7069 (N_7069,N_6060,N_6898);
xnor U7070 (N_7070,N_6371,N_6668);
or U7071 (N_7071,N_6498,N_6851);
nand U7072 (N_7072,N_6440,N_6603);
nand U7073 (N_7073,N_6360,N_6826);
nand U7074 (N_7074,N_6839,N_6303);
or U7075 (N_7075,N_6931,N_6773);
nand U7076 (N_7076,N_6483,N_6967);
or U7077 (N_7077,N_6533,N_6973);
or U7078 (N_7078,N_6122,N_6161);
nand U7079 (N_7079,N_6127,N_6414);
and U7080 (N_7080,N_6490,N_6223);
xnor U7081 (N_7081,N_6312,N_6363);
nand U7082 (N_7082,N_6934,N_6020);
or U7083 (N_7083,N_6307,N_6191);
or U7084 (N_7084,N_6452,N_6720);
nand U7085 (N_7085,N_6576,N_6772);
nand U7086 (N_7086,N_6577,N_6098);
and U7087 (N_7087,N_6166,N_6173);
nand U7088 (N_7088,N_6197,N_6325);
nand U7089 (N_7089,N_6294,N_6854);
xnor U7090 (N_7090,N_6940,N_6887);
nand U7091 (N_7091,N_6843,N_6183);
nor U7092 (N_7092,N_6313,N_6838);
xnor U7093 (N_7093,N_6907,N_6090);
or U7094 (N_7094,N_6625,N_6052);
xor U7095 (N_7095,N_6587,N_6339);
xnor U7096 (N_7096,N_6462,N_6870);
or U7097 (N_7097,N_6290,N_6141);
nand U7098 (N_7098,N_6811,N_6517);
nor U7099 (N_7099,N_6008,N_6340);
xor U7100 (N_7100,N_6231,N_6609);
and U7101 (N_7101,N_6971,N_6002);
nand U7102 (N_7102,N_6798,N_6692);
or U7103 (N_7103,N_6477,N_6413);
nor U7104 (N_7104,N_6757,N_6540);
nand U7105 (N_7105,N_6082,N_6886);
nand U7106 (N_7106,N_6874,N_6953);
nand U7107 (N_7107,N_6754,N_6788);
and U7108 (N_7108,N_6880,N_6017);
or U7109 (N_7109,N_6030,N_6561);
nor U7110 (N_7110,N_6145,N_6941);
xor U7111 (N_7111,N_6997,N_6428);
nand U7112 (N_7112,N_6523,N_6251);
and U7113 (N_7113,N_6960,N_6373);
nor U7114 (N_7114,N_6853,N_6512);
nor U7115 (N_7115,N_6084,N_6001);
nand U7116 (N_7116,N_6107,N_6486);
and U7117 (N_7117,N_6733,N_6833);
or U7118 (N_7118,N_6855,N_6432);
and U7119 (N_7119,N_6664,N_6694);
nor U7120 (N_7120,N_6895,N_6203);
and U7121 (N_7121,N_6518,N_6553);
and U7122 (N_7122,N_6234,N_6276);
xor U7123 (N_7123,N_6072,N_6400);
xor U7124 (N_7124,N_6126,N_6321);
and U7125 (N_7125,N_6902,N_6601);
xnor U7126 (N_7126,N_6021,N_6463);
and U7127 (N_7127,N_6386,N_6808);
nor U7128 (N_7128,N_6885,N_6465);
or U7129 (N_7129,N_6153,N_6491);
nor U7130 (N_7130,N_6981,N_6978);
and U7131 (N_7131,N_6097,N_6123);
nor U7132 (N_7132,N_6007,N_6421);
nand U7133 (N_7133,N_6554,N_6441);
nand U7134 (N_7134,N_6894,N_6205);
and U7135 (N_7135,N_6110,N_6538);
and U7136 (N_7136,N_6096,N_6306);
nand U7137 (N_7137,N_6322,N_6388);
nor U7138 (N_7138,N_6326,N_6682);
nor U7139 (N_7139,N_6435,N_6285);
nand U7140 (N_7140,N_6502,N_6129);
nand U7141 (N_7141,N_6627,N_6575);
and U7142 (N_7142,N_6226,N_6447);
or U7143 (N_7143,N_6741,N_6514);
nor U7144 (N_7144,N_6479,N_6207);
nand U7145 (N_7145,N_6936,N_6257);
xor U7146 (N_7146,N_6611,N_6748);
nor U7147 (N_7147,N_6891,N_6423);
nand U7148 (N_7148,N_6275,N_6488);
and U7149 (N_7149,N_6825,N_6824);
or U7150 (N_7150,N_6726,N_6737);
nand U7151 (N_7151,N_6781,N_6248);
or U7152 (N_7152,N_6146,N_6521);
xor U7153 (N_7153,N_6291,N_6000);
xor U7154 (N_7154,N_6293,N_6599);
nand U7155 (N_7155,N_6287,N_6649);
nand U7156 (N_7156,N_6963,N_6982);
and U7157 (N_7157,N_6335,N_6190);
or U7158 (N_7158,N_6069,N_6792);
and U7159 (N_7159,N_6018,N_6316);
nor U7160 (N_7160,N_6023,N_6039);
or U7161 (N_7161,N_6154,N_6579);
and U7162 (N_7162,N_6590,N_6188);
xnor U7163 (N_7163,N_6796,N_6113);
nand U7164 (N_7164,N_6889,N_6375);
nor U7165 (N_7165,N_6487,N_6526);
nor U7166 (N_7166,N_6025,N_6242);
or U7167 (N_7167,N_6939,N_6394);
or U7168 (N_7168,N_6474,N_6716);
or U7169 (N_7169,N_6229,N_6383);
xor U7170 (N_7170,N_6063,N_6950);
nor U7171 (N_7171,N_6172,N_6678);
xnor U7172 (N_7172,N_6047,N_6774);
or U7173 (N_7173,N_6308,N_6262);
or U7174 (N_7174,N_6731,N_6859);
nor U7175 (N_7175,N_6565,N_6673);
xnor U7176 (N_7176,N_6496,N_6571);
xor U7177 (N_7177,N_6543,N_6747);
nor U7178 (N_7178,N_6377,N_6613);
nor U7179 (N_7179,N_6743,N_6124);
nand U7180 (N_7180,N_6661,N_6168);
xor U7181 (N_7181,N_6708,N_6948);
nor U7182 (N_7182,N_6102,N_6238);
or U7183 (N_7183,N_6279,N_6975);
nor U7184 (N_7184,N_6660,N_6648);
or U7185 (N_7185,N_6901,N_6681);
nor U7186 (N_7186,N_6158,N_6142);
xnor U7187 (N_7187,N_6167,N_6473);
nor U7188 (N_7188,N_6602,N_6979);
and U7189 (N_7189,N_6504,N_6445);
nand U7190 (N_7190,N_6497,N_6861);
nand U7191 (N_7191,N_6845,N_6443);
and U7192 (N_7192,N_6888,N_6460);
and U7193 (N_7193,N_6013,N_6766);
nand U7194 (N_7194,N_6823,N_6770);
nand U7195 (N_7195,N_6382,N_6489);
xnor U7196 (N_7196,N_6959,N_6471);
xnor U7197 (N_7197,N_6639,N_6729);
and U7198 (N_7198,N_6568,N_6701);
and U7199 (N_7199,N_6913,N_6209);
and U7200 (N_7200,N_6019,N_6910);
xor U7201 (N_7201,N_6105,N_6187);
nor U7202 (N_7202,N_6091,N_6669);
xnor U7203 (N_7203,N_6448,N_6050);
nand U7204 (N_7204,N_6134,N_6434);
nor U7205 (N_7205,N_6858,N_6955);
and U7206 (N_7206,N_6724,N_6643);
nand U7207 (N_7207,N_6470,N_6131);
nand U7208 (N_7208,N_6011,N_6755);
nor U7209 (N_7209,N_6482,N_6787);
nand U7210 (N_7210,N_6071,N_6679);
nor U7211 (N_7211,N_6580,N_6856);
nand U7212 (N_7212,N_6529,N_6624);
or U7213 (N_7213,N_6403,N_6282);
and U7214 (N_7214,N_6652,N_6921);
nor U7215 (N_7215,N_6943,N_6711);
and U7216 (N_7216,N_6365,N_6278);
nand U7217 (N_7217,N_6546,N_6728);
or U7218 (N_7218,N_6961,N_6356);
or U7219 (N_7219,N_6746,N_6380);
xor U7220 (N_7220,N_6264,N_6806);
or U7221 (N_7221,N_6872,N_6528);
nor U7222 (N_7222,N_6763,N_6993);
xnor U7223 (N_7223,N_6202,N_6867);
or U7224 (N_7224,N_6892,N_6507);
xor U7225 (N_7225,N_6032,N_6138);
xor U7226 (N_7226,N_6212,N_6369);
or U7227 (N_7227,N_6399,N_6244);
or U7228 (N_7228,N_6051,N_6233);
nor U7229 (N_7229,N_6079,N_6884);
xnor U7230 (N_7230,N_6405,N_6947);
nor U7231 (N_7231,N_6516,N_6680);
xor U7232 (N_7232,N_6401,N_6454);
or U7233 (N_7233,N_6835,N_6596);
nand U7234 (N_7234,N_6323,N_6905);
nand U7235 (N_7235,N_6789,N_6222);
xnor U7236 (N_7236,N_6989,N_6566);
and U7237 (N_7237,N_6268,N_6208);
or U7238 (N_7238,N_6150,N_6837);
or U7239 (N_7239,N_6850,N_6607);
and U7240 (N_7240,N_6924,N_6431);
nand U7241 (N_7241,N_6879,N_6174);
nand U7242 (N_7242,N_6416,N_6480);
or U7243 (N_7243,N_6503,N_6584);
or U7244 (N_7244,N_6745,N_6178);
or U7245 (N_7245,N_6310,N_6878);
or U7246 (N_7246,N_6387,N_6524);
nor U7247 (N_7247,N_6976,N_6593);
nand U7248 (N_7248,N_6830,N_6799);
nor U7249 (N_7249,N_6685,N_6557);
and U7250 (N_7250,N_6598,N_6906);
nor U7251 (N_7251,N_6803,N_6918);
and U7252 (N_7252,N_6705,N_6563);
and U7253 (N_7253,N_6646,N_6152);
xor U7254 (N_7254,N_6548,N_6476);
xnor U7255 (N_7255,N_6016,N_6942);
nand U7256 (N_7256,N_6130,N_6569);
or U7257 (N_7257,N_6299,N_6204);
nor U7258 (N_7258,N_6327,N_6143);
nor U7259 (N_7259,N_6121,N_6937);
xor U7260 (N_7260,N_6289,N_6137);
or U7261 (N_7261,N_6620,N_6994);
and U7262 (N_7262,N_6714,N_6427);
or U7263 (N_7263,N_6877,N_6702);
nor U7264 (N_7264,N_6225,N_6847);
xor U7265 (N_7265,N_6128,N_6085);
nor U7266 (N_7266,N_6793,N_6663);
xor U7267 (N_7267,N_6311,N_6272);
and U7268 (N_7268,N_6795,N_6241);
nor U7269 (N_7269,N_6304,N_6033);
or U7270 (N_7270,N_6043,N_6406);
and U7271 (N_7271,N_6227,N_6634);
xnor U7272 (N_7272,N_6184,N_6156);
nor U7273 (N_7273,N_6604,N_6560);
or U7274 (N_7274,N_6623,N_6621);
or U7275 (N_7275,N_6672,N_6281);
xor U7276 (N_7276,N_6253,N_6641);
xnor U7277 (N_7277,N_6535,N_6536);
xor U7278 (N_7278,N_6573,N_6157);
nor U7279 (N_7279,N_6429,N_6783);
or U7280 (N_7280,N_6995,N_6106);
and U7281 (N_7281,N_6352,N_6265);
or U7282 (N_7282,N_6896,N_6366);
nor U7283 (N_7283,N_6710,N_6337);
and U7284 (N_7284,N_6761,N_6062);
and U7285 (N_7285,N_6564,N_6341);
xnor U7286 (N_7286,N_6464,N_6250);
nand U7287 (N_7287,N_6391,N_6351);
nor U7288 (N_7288,N_6812,N_6656);
nand U7289 (N_7289,N_6619,N_6374);
and U7290 (N_7290,N_6562,N_6232);
xor U7291 (N_7291,N_6805,N_6344);
or U7292 (N_7292,N_6667,N_6511);
xor U7293 (N_7293,N_6331,N_6904);
xor U7294 (N_7294,N_6088,N_6539);
nor U7295 (N_7295,N_6461,N_6438);
xnor U7296 (N_7296,N_6005,N_6055);
or U7297 (N_7297,N_6455,N_6645);
or U7298 (N_7298,N_6368,N_6029);
or U7299 (N_7299,N_6508,N_6952);
xnor U7300 (N_7300,N_6735,N_6776);
and U7301 (N_7301,N_6636,N_6343);
or U7302 (N_7302,N_6964,N_6249);
nor U7303 (N_7303,N_6402,N_6751);
xor U7304 (N_7304,N_6220,N_6068);
nand U7305 (N_7305,N_6417,N_6420);
nor U7306 (N_7306,N_6252,N_6844);
nor U7307 (N_7307,N_6099,N_6970);
and U7308 (N_7308,N_6570,N_6920);
nor U7309 (N_7309,N_6618,N_6396);
nor U7310 (N_7310,N_6006,N_6478);
or U7311 (N_7311,N_6444,N_6530);
and U7312 (N_7312,N_6235,N_6592);
and U7313 (N_7313,N_6012,N_6453);
and U7314 (N_7314,N_6458,N_6713);
nand U7315 (N_7315,N_6688,N_6689);
xor U7316 (N_7316,N_6977,N_6346);
nand U7317 (N_7317,N_6355,N_6608);
nand U7318 (N_7318,N_6659,N_6330);
nand U7319 (N_7319,N_6638,N_6022);
and U7320 (N_7320,N_6626,N_6760);
xor U7321 (N_7321,N_6298,N_6500);
nor U7322 (N_7322,N_6348,N_6398);
or U7323 (N_7323,N_6574,N_6078);
and U7324 (N_7324,N_6037,N_6064);
and U7325 (N_7325,N_6738,N_6111);
xor U7326 (N_7326,N_6430,N_6722);
and U7327 (N_7327,N_6984,N_6762);
or U7328 (N_7328,N_6690,N_6800);
nor U7329 (N_7329,N_6545,N_6314);
xor U7330 (N_7330,N_6662,N_6848);
and U7331 (N_7331,N_6695,N_6765);
nand U7332 (N_7332,N_6451,N_6459);
nor U7333 (N_7333,N_6270,N_6467);
nand U7334 (N_7334,N_6415,N_6520);
xnor U7335 (N_7335,N_6116,N_6992);
nand U7336 (N_7336,N_6309,N_6378);
xnor U7337 (N_7337,N_6697,N_6010);
nand U7338 (N_7338,N_6333,N_6860);
nor U7339 (N_7339,N_6785,N_6425);
or U7340 (N_7340,N_6542,N_6778);
xor U7341 (N_7341,N_6115,N_6671);
or U7342 (N_7342,N_6784,N_6181);
and U7343 (N_7343,N_6998,N_6319);
xnor U7344 (N_7344,N_6136,N_6198);
nand U7345 (N_7345,N_6846,N_6868);
or U7346 (N_7346,N_6591,N_6067);
or U7347 (N_7347,N_6744,N_6756);
nor U7348 (N_7348,N_6631,N_6534);
xor U7349 (N_7349,N_6024,N_6318);
nand U7350 (N_7350,N_6089,N_6182);
and U7351 (N_7351,N_6266,N_6666);
xnor U7352 (N_7352,N_6883,N_6015);
xor U7353 (N_7353,N_6258,N_6969);
or U7354 (N_7354,N_6810,N_6911);
and U7355 (N_7355,N_6586,N_6054);
or U7356 (N_7356,N_6243,N_6362);
nor U7357 (N_7357,N_6769,N_6815);
xnor U7358 (N_7358,N_6186,N_6758);
nand U7359 (N_7359,N_6370,N_6436);
nand U7360 (N_7360,N_6882,N_6510);
and U7361 (N_7361,N_6957,N_6114);
or U7362 (N_7362,N_6836,N_6519);
nor U7363 (N_7363,N_6712,N_6164);
and U7364 (N_7364,N_6449,N_6890);
nor U7365 (N_7365,N_6509,N_6112);
xnor U7366 (N_7366,N_6658,N_6556);
and U7367 (N_7367,N_6552,N_6014);
nor U7368 (N_7368,N_6842,N_6653);
nand U7369 (N_7369,N_6206,N_6151);
xnor U7370 (N_7370,N_6210,N_6916);
nor U7371 (N_7371,N_6929,N_6359);
xnor U7372 (N_7372,N_6230,N_6389);
nand U7373 (N_7373,N_6732,N_6442);
and U7374 (N_7374,N_6817,N_6922);
xnor U7375 (N_7375,N_6585,N_6329);
nand U7376 (N_7376,N_6674,N_6261);
xnor U7377 (N_7377,N_6919,N_6347);
xor U7378 (N_7378,N_6259,N_6696);
nand U7379 (N_7379,N_6600,N_6439);
or U7380 (N_7380,N_6730,N_6059);
or U7381 (N_7381,N_6009,N_6683);
nand U7382 (N_7382,N_6677,N_6897);
and U7383 (N_7383,N_6866,N_6424);
xor U7384 (N_7384,N_6159,N_6767);
or U7385 (N_7385,N_6004,N_6295);
nand U7386 (N_7386,N_6221,N_6693);
nor U7387 (N_7387,N_6194,N_6834);
xnor U7388 (N_7388,N_6999,N_6410);
nand U7389 (N_7389,N_6393,N_6108);
or U7390 (N_7390,N_6254,N_6821);
nand U7391 (N_7391,N_6367,N_6986);
nand U7392 (N_7392,N_6832,N_6903);
nor U7393 (N_7393,N_6996,N_6777);
xor U7394 (N_7394,N_6768,N_6555);
xor U7395 (N_7395,N_6614,N_6372);
nand U7396 (N_7396,N_6956,N_6698);
and U7397 (N_7397,N_6237,N_6869);
or U7398 (N_7398,N_6635,N_6450);
or U7399 (N_7399,N_6034,N_6466);
or U7400 (N_7400,N_6255,N_6475);
and U7401 (N_7401,N_6630,N_6816);
nor U7402 (N_7402,N_6819,N_6095);
nand U7403 (N_7403,N_6092,N_6925);
nand U7404 (N_7404,N_6390,N_6501);
and U7405 (N_7405,N_6742,N_6949);
and U7406 (N_7406,N_6109,N_6628);
or U7407 (N_7407,N_6286,N_6135);
and U7408 (N_7408,N_6094,N_6481);
xnor U7409 (N_7409,N_6042,N_6987);
xor U7410 (N_7410,N_6684,N_6617);
nor U7411 (N_7411,N_6899,N_6053);
xnor U7412 (N_7412,N_6040,N_6657);
nand U7413 (N_7413,N_6283,N_6058);
nand U7414 (N_7414,N_6280,N_6219);
xor U7415 (N_7415,N_6699,N_6165);
and U7416 (N_7416,N_6595,N_6828);
xor U7417 (N_7417,N_6300,N_6140);
nor U7418 (N_7418,N_6779,N_6407);
nand U7419 (N_7419,N_6041,N_6820);
nor U7420 (N_7420,N_6814,N_6637);
and U7421 (N_7421,N_6076,N_6893);
and U7422 (N_7422,N_6946,N_6522);
xor U7423 (N_7423,N_6876,N_6066);
or U7424 (N_7424,N_6932,N_6718);
or U7425 (N_7425,N_6809,N_6831);
xnor U7426 (N_7426,N_6484,N_6133);
xor U7427 (N_7427,N_6342,N_6544);
and U7428 (N_7428,N_6048,N_6036);
or U7429 (N_7429,N_6384,N_6912);
xnor U7430 (N_7430,N_6199,N_6715);
or U7431 (N_7431,N_6104,N_6515);
nor U7432 (N_7432,N_6176,N_6119);
nor U7433 (N_7433,N_6764,N_6551);
or U7434 (N_7434,N_6813,N_6065);
xnor U7435 (N_7435,N_6954,N_6909);
and U7436 (N_7436,N_6818,N_6972);
nand U7437 (N_7437,N_6260,N_6080);
nand U7438 (N_7438,N_6691,N_6944);
and U7439 (N_7439,N_6531,N_6610);
xnor U7440 (N_7440,N_6338,N_6385);
and U7441 (N_7441,N_6750,N_6162);
xor U7442 (N_7442,N_6988,N_6873);
or U7443 (N_7443,N_6633,N_6118);
xor U7444 (N_7444,N_6179,N_6247);
nor U7445 (N_7445,N_6651,N_6317);
xor U7446 (N_7446,N_6263,N_6277);
nor U7447 (N_7447,N_6073,N_6228);
or U7448 (N_7448,N_6930,N_6807);
nand U7449 (N_7449,N_6426,N_6103);
nand U7450 (N_7450,N_6525,N_6915);
xor U7451 (N_7451,N_6704,N_6700);
and U7452 (N_7452,N_6302,N_6938);
xor U7453 (N_7453,N_6974,N_6180);
xnor U7454 (N_7454,N_6706,N_6397);
or U7455 (N_7455,N_6336,N_6629);
xnor U7456 (N_7456,N_6594,N_6749);
and U7457 (N_7457,N_6597,N_6185);
nand U7458 (N_7458,N_6642,N_6703);
nor U7459 (N_7459,N_6900,N_6155);
nor U7460 (N_7460,N_6725,N_6822);
nor U7461 (N_7461,N_6081,N_6727);
and U7462 (N_7462,N_6379,N_6419);
xnor U7463 (N_7463,N_6046,N_6038);
nand U7464 (N_7464,N_6686,N_6790);
xor U7465 (N_7465,N_6928,N_6709);
or U7466 (N_7466,N_6494,N_6655);
or U7467 (N_7467,N_6101,N_6003);
xor U7468 (N_7468,N_6615,N_6349);
nand U7469 (N_7469,N_6171,N_6086);
nand U7470 (N_7470,N_6865,N_6404);
nand U7471 (N_7471,N_6274,N_6840);
nor U7472 (N_7472,N_6881,N_6117);
or U7473 (N_7473,N_6802,N_6305);
nand U7474 (N_7474,N_6328,N_6334);
xnor U7475 (N_7475,N_6297,N_6160);
xor U7476 (N_7476,N_6364,N_6049);
nand U7477 (N_7477,N_6527,N_6605);
nor U7478 (N_7478,N_6211,N_6771);
nor U7479 (N_7479,N_6485,N_6193);
or U7480 (N_7480,N_6125,N_6862);
nor U7481 (N_7481,N_6345,N_6147);
xor U7482 (N_7482,N_6985,N_6644);
xnor U7483 (N_7483,N_6736,N_6028);
nor U7484 (N_7484,N_6582,N_6506);
xnor U7485 (N_7485,N_6215,N_6547);
xnor U7486 (N_7486,N_6782,N_6395);
nand U7487 (N_7487,N_6558,N_6189);
and U7488 (N_7488,N_6216,N_6056);
or U7489 (N_7489,N_6332,N_6120);
and U7490 (N_7490,N_6493,N_6408);
and U7491 (N_7491,N_6412,N_6739);
nand U7492 (N_7492,N_6315,N_6457);
xnor U7493 (N_7493,N_6083,N_6965);
or U7494 (N_7494,N_6966,N_6301);
nor U7495 (N_7495,N_6864,N_6213);
nor U7496 (N_7496,N_6236,N_6381);
nor U7497 (N_7497,N_6780,N_6177);
or U7498 (N_7498,N_6841,N_6572);
or U7499 (N_7499,N_6070,N_6917);
nor U7500 (N_7500,N_6136,N_6025);
or U7501 (N_7501,N_6254,N_6468);
nand U7502 (N_7502,N_6631,N_6372);
and U7503 (N_7503,N_6170,N_6278);
nor U7504 (N_7504,N_6426,N_6134);
nand U7505 (N_7505,N_6202,N_6741);
or U7506 (N_7506,N_6154,N_6503);
nand U7507 (N_7507,N_6508,N_6190);
and U7508 (N_7508,N_6702,N_6927);
nand U7509 (N_7509,N_6297,N_6524);
nor U7510 (N_7510,N_6589,N_6329);
nand U7511 (N_7511,N_6568,N_6118);
nor U7512 (N_7512,N_6561,N_6770);
nand U7513 (N_7513,N_6165,N_6049);
xor U7514 (N_7514,N_6295,N_6896);
xor U7515 (N_7515,N_6927,N_6963);
nand U7516 (N_7516,N_6198,N_6962);
or U7517 (N_7517,N_6521,N_6283);
and U7518 (N_7518,N_6479,N_6039);
and U7519 (N_7519,N_6243,N_6648);
or U7520 (N_7520,N_6446,N_6172);
xor U7521 (N_7521,N_6406,N_6678);
xor U7522 (N_7522,N_6902,N_6368);
nor U7523 (N_7523,N_6179,N_6096);
and U7524 (N_7524,N_6245,N_6885);
and U7525 (N_7525,N_6462,N_6233);
nand U7526 (N_7526,N_6322,N_6802);
xor U7527 (N_7527,N_6883,N_6855);
xnor U7528 (N_7528,N_6898,N_6385);
and U7529 (N_7529,N_6017,N_6908);
and U7530 (N_7530,N_6357,N_6299);
xnor U7531 (N_7531,N_6119,N_6397);
or U7532 (N_7532,N_6754,N_6238);
and U7533 (N_7533,N_6278,N_6664);
nand U7534 (N_7534,N_6054,N_6424);
nand U7535 (N_7535,N_6908,N_6388);
nor U7536 (N_7536,N_6413,N_6362);
and U7537 (N_7537,N_6998,N_6324);
or U7538 (N_7538,N_6983,N_6761);
xnor U7539 (N_7539,N_6549,N_6333);
nand U7540 (N_7540,N_6875,N_6551);
and U7541 (N_7541,N_6690,N_6716);
and U7542 (N_7542,N_6964,N_6508);
or U7543 (N_7543,N_6219,N_6946);
and U7544 (N_7544,N_6126,N_6482);
xnor U7545 (N_7545,N_6882,N_6679);
and U7546 (N_7546,N_6520,N_6169);
nand U7547 (N_7547,N_6114,N_6567);
or U7548 (N_7548,N_6985,N_6296);
nor U7549 (N_7549,N_6869,N_6251);
nor U7550 (N_7550,N_6597,N_6662);
xor U7551 (N_7551,N_6795,N_6191);
nor U7552 (N_7552,N_6310,N_6122);
xnor U7553 (N_7553,N_6627,N_6334);
nor U7554 (N_7554,N_6223,N_6033);
or U7555 (N_7555,N_6170,N_6327);
nor U7556 (N_7556,N_6523,N_6269);
xor U7557 (N_7557,N_6519,N_6692);
nor U7558 (N_7558,N_6757,N_6899);
or U7559 (N_7559,N_6008,N_6893);
nand U7560 (N_7560,N_6101,N_6072);
and U7561 (N_7561,N_6736,N_6049);
xnor U7562 (N_7562,N_6513,N_6636);
or U7563 (N_7563,N_6443,N_6127);
xor U7564 (N_7564,N_6122,N_6679);
nor U7565 (N_7565,N_6922,N_6177);
nor U7566 (N_7566,N_6496,N_6386);
nor U7567 (N_7567,N_6862,N_6307);
nand U7568 (N_7568,N_6073,N_6175);
and U7569 (N_7569,N_6941,N_6389);
xnor U7570 (N_7570,N_6293,N_6813);
nor U7571 (N_7571,N_6260,N_6556);
or U7572 (N_7572,N_6147,N_6837);
and U7573 (N_7573,N_6130,N_6231);
and U7574 (N_7574,N_6320,N_6404);
nor U7575 (N_7575,N_6888,N_6874);
xor U7576 (N_7576,N_6092,N_6875);
nor U7577 (N_7577,N_6618,N_6264);
and U7578 (N_7578,N_6003,N_6481);
and U7579 (N_7579,N_6230,N_6703);
or U7580 (N_7580,N_6074,N_6050);
nand U7581 (N_7581,N_6223,N_6848);
and U7582 (N_7582,N_6769,N_6665);
nor U7583 (N_7583,N_6550,N_6109);
xor U7584 (N_7584,N_6826,N_6179);
nand U7585 (N_7585,N_6879,N_6709);
xnor U7586 (N_7586,N_6277,N_6106);
nor U7587 (N_7587,N_6525,N_6660);
or U7588 (N_7588,N_6009,N_6270);
nor U7589 (N_7589,N_6507,N_6731);
and U7590 (N_7590,N_6649,N_6454);
nor U7591 (N_7591,N_6622,N_6063);
and U7592 (N_7592,N_6344,N_6557);
or U7593 (N_7593,N_6913,N_6750);
and U7594 (N_7594,N_6408,N_6314);
nand U7595 (N_7595,N_6027,N_6549);
nor U7596 (N_7596,N_6616,N_6752);
and U7597 (N_7597,N_6640,N_6439);
nand U7598 (N_7598,N_6232,N_6230);
nor U7599 (N_7599,N_6433,N_6585);
nand U7600 (N_7600,N_6262,N_6261);
xnor U7601 (N_7601,N_6289,N_6627);
xnor U7602 (N_7602,N_6501,N_6170);
nor U7603 (N_7603,N_6589,N_6707);
or U7604 (N_7604,N_6783,N_6791);
and U7605 (N_7605,N_6788,N_6575);
and U7606 (N_7606,N_6175,N_6020);
nand U7607 (N_7607,N_6859,N_6010);
xnor U7608 (N_7608,N_6629,N_6845);
or U7609 (N_7609,N_6860,N_6471);
and U7610 (N_7610,N_6807,N_6787);
or U7611 (N_7611,N_6117,N_6303);
and U7612 (N_7612,N_6603,N_6488);
xnor U7613 (N_7613,N_6094,N_6388);
xor U7614 (N_7614,N_6136,N_6038);
and U7615 (N_7615,N_6626,N_6048);
and U7616 (N_7616,N_6657,N_6496);
and U7617 (N_7617,N_6080,N_6945);
and U7618 (N_7618,N_6266,N_6468);
nor U7619 (N_7619,N_6434,N_6991);
nor U7620 (N_7620,N_6835,N_6651);
nor U7621 (N_7621,N_6982,N_6589);
nand U7622 (N_7622,N_6247,N_6228);
and U7623 (N_7623,N_6215,N_6960);
nor U7624 (N_7624,N_6200,N_6823);
and U7625 (N_7625,N_6701,N_6388);
nand U7626 (N_7626,N_6051,N_6303);
or U7627 (N_7627,N_6104,N_6986);
and U7628 (N_7628,N_6998,N_6805);
and U7629 (N_7629,N_6438,N_6963);
or U7630 (N_7630,N_6965,N_6795);
xor U7631 (N_7631,N_6293,N_6593);
nand U7632 (N_7632,N_6595,N_6237);
nand U7633 (N_7633,N_6157,N_6666);
and U7634 (N_7634,N_6632,N_6952);
nand U7635 (N_7635,N_6745,N_6090);
or U7636 (N_7636,N_6723,N_6367);
nor U7637 (N_7637,N_6471,N_6737);
nor U7638 (N_7638,N_6059,N_6944);
xor U7639 (N_7639,N_6574,N_6414);
nand U7640 (N_7640,N_6020,N_6577);
xnor U7641 (N_7641,N_6468,N_6249);
nor U7642 (N_7642,N_6822,N_6051);
nor U7643 (N_7643,N_6396,N_6264);
nand U7644 (N_7644,N_6096,N_6123);
and U7645 (N_7645,N_6271,N_6904);
xnor U7646 (N_7646,N_6714,N_6033);
and U7647 (N_7647,N_6134,N_6310);
xor U7648 (N_7648,N_6287,N_6077);
xor U7649 (N_7649,N_6109,N_6957);
xnor U7650 (N_7650,N_6572,N_6029);
and U7651 (N_7651,N_6499,N_6196);
nor U7652 (N_7652,N_6908,N_6391);
or U7653 (N_7653,N_6333,N_6206);
or U7654 (N_7654,N_6812,N_6654);
xor U7655 (N_7655,N_6914,N_6649);
xnor U7656 (N_7656,N_6558,N_6759);
or U7657 (N_7657,N_6434,N_6287);
nand U7658 (N_7658,N_6799,N_6798);
nor U7659 (N_7659,N_6074,N_6954);
and U7660 (N_7660,N_6293,N_6505);
nand U7661 (N_7661,N_6168,N_6359);
nor U7662 (N_7662,N_6267,N_6421);
nand U7663 (N_7663,N_6400,N_6211);
xor U7664 (N_7664,N_6966,N_6273);
xnor U7665 (N_7665,N_6639,N_6046);
xor U7666 (N_7666,N_6741,N_6985);
nor U7667 (N_7667,N_6052,N_6463);
or U7668 (N_7668,N_6700,N_6052);
nor U7669 (N_7669,N_6473,N_6579);
nor U7670 (N_7670,N_6442,N_6711);
xor U7671 (N_7671,N_6175,N_6889);
nand U7672 (N_7672,N_6531,N_6575);
and U7673 (N_7673,N_6912,N_6284);
nor U7674 (N_7674,N_6013,N_6322);
nor U7675 (N_7675,N_6911,N_6195);
xnor U7676 (N_7676,N_6657,N_6739);
nor U7677 (N_7677,N_6750,N_6275);
and U7678 (N_7678,N_6713,N_6176);
and U7679 (N_7679,N_6968,N_6948);
nor U7680 (N_7680,N_6313,N_6572);
or U7681 (N_7681,N_6132,N_6453);
nor U7682 (N_7682,N_6155,N_6020);
xor U7683 (N_7683,N_6613,N_6087);
and U7684 (N_7684,N_6644,N_6649);
nand U7685 (N_7685,N_6160,N_6335);
xnor U7686 (N_7686,N_6656,N_6777);
nor U7687 (N_7687,N_6202,N_6950);
xnor U7688 (N_7688,N_6737,N_6122);
or U7689 (N_7689,N_6064,N_6766);
or U7690 (N_7690,N_6171,N_6793);
and U7691 (N_7691,N_6081,N_6628);
xor U7692 (N_7692,N_6382,N_6643);
nor U7693 (N_7693,N_6370,N_6512);
nor U7694 (N_7694,N_6434,N_6488);
or U7695 (N_7695,N_6199,N_6505);
xnor U7696 (N_7696,N_6701,N_6127);
xnor U7697 (N_7697,N_6217,N_6633);
and U7698 (N_7698,N_6210,N_6182);
or U7699 (N_7699,N_6721,N_6861);
nand U7700 (N_7700,N_6915,N_6620);
nand U7701 (N_7701,N_6528,N_6896);
and U7702 (N_7702,N_6325,N_6242);
or U7703 (N_7703,N_6020,N_6690);
xnor U7704 (N_7704,N_6498,N_6326);
or U7705 (N_7705,N_6697,N_6272);
nand U7706 (N_7706,N_6793,N_6645);
nand U7707 (N_7707,N_6386,N_6349);
or U7708 (N_7708,N_6442,N_6228);
or U7709 (N_7709,N_6133,N_6440);
nand U7710 (N_7710,N_6139,N_6322);
nor U7711 (N_7711,N_6450,N_6282);
and U7712 (N_7712,N_6288,N_6487);
xnor U7713 (N_7713,N_6254,N_6057);
xor U7714 (N_7714,N_6723,N_6619);
nor U7715 (N_7715,N_6465,N_6264);
and U7716 (N_7716,N_6171,N_6647);
nand U7717 (N_7717,N_6619,N_6266);
and U7718 (N_7718,N_6111,N_6760);
xnor U7719 (N_7719,N_6772,N_6423);
nor U7720 (N_7720,N_6614,N_6545);
and U7721 (N_7721,N_6536,N_6798);
nand U7722 (N_7722,N_6327,N_6895);
nand U7723 (N_7723,N_6350,N_6373);
and U7724 (N_7724,N_6042,N_6307);
and U7725 (N_7725,N_6011,N_6881);
or U7726 (N_7726,N_6874,N_6087);
xor U7727 (N_7727,N_6174,N_6978);
or U7728 (N_7728,N_6796,N_6872);
and U7729 (N_7729,N_6815,N_6280);
xor U7730 (N_7730,N_6322,N_6385);
and U7731 (N_7731,N_6403,N_6414);
xnor U7732 (N_7732,N_6070,N_6998);
xnor U7733 (N_7733,N_6148,N_6772);
and U7734 (N_7734,N_6561,N_6440);
nor U7735 (N_7735,N_6459,N_6211);
nor U7736 (N_7736,N_6802,N_6432);
or U7737 (N_7737,N_6992,N_6673);
xnor U7738 (N_7738,N_6380,N_6226);
xor U7739 (N_7739,N_6855,N_6572);
or U7740 (N_7740,N_6040,N_6332);
nor U7741 (N_7741,N_6328,N_6260);
nand U7742 (N_7742,N_6365,N_6752);
nand U7743 (N_7743,N_6264,N_6411);
xnor U7744 (N_7744,N_6158,N_6702);
xnor U7745 (N_7745,N_6332,N_6813);
or U7746 (N_7746,N_6186,N_6302);
and U7747 (N_7747,N_6909,N_6593);
xor U7748 (N_7748,N_6071,N_6819);
nor U7749 (N_7749,N_6086,N_6127);
and U7750 (N_7750,N_6402,N_6205);
or U7751 (N_7751,N_6372,N_6692);
xnor U7752 (N_7752,N_6870,N_6285);
nor U7753 (N_7753,N_6721,N_6735);
nor U7754 (N_7754,N_6138,N_6589);
xnor U7755 (N_7755,N_6477,N_6144);
or U7756 (N_7756,N_6408,N_6830);
nor U7757 (N_7757,N_6127,N_6159);
and U7758 (N_7758,N_6325,N_6485);
and U7759 (N_7759,N_6244,N_6500);
and U7760 (N_7760,N_6907,N_6270);
nand U7761 (N_7761,N_6096,N_6880);
nand U7762 (N_7762,N_6356,N_6374);
and U7763 (N_7763,N_6487,N_6003);
and U7764 (N_7764,N_6310,N_6354);
nand U7765 (N_7765,N_6882,N_6270);
or U7766 (N_7766,N_6816,N_6081);
or U7767 (N_7767,N_6053,N_6568);
nand U7768 (N_7768,N_6885,N_6077);
and U7769 (N_7769,N_6002,N_6821);
or U7770 (N_7770,N_6056,N_6302);
and U7771 (N_7771,N_6304,N_6249);
or U7772 (N_7772,N_6703,N_6891);
xnor U7773 (N_7773,N_6191,N_6849);
xor U7774 (N_7774,N_6297,N_6284);
nand U7775 (N_7775,N_6626,N_6930);
nor U7776 (N_7776,N_6562,N_6110);
or U7777 (N_7777,N_6647,N_6458);
nor U7778 (N_7778,N_6843,N_6621);
xor U7779 (N_7779,N_6875,N_6087);
or U7780 (N_7780,N_6581,N_6549);
nand U7781 (N_7781,N_6277,N_6081);
xnor U7782 (N_7782,N_6177,N_6691);
nand U7783 (N_7783,N_6763,N_6480);
nand U7784 (N_7784,N_6461,N_6521);
or U7785 (N_7785,N_6954,N_6055);
nor U7786 (N_7786,N_6288,N_6069);
and U7787 (N_7787,N_6405,N_6616);
xor U7788 (N_7788,N_6423,N_6115);
or U7789 (N_7789,N_6955,N_6506);
nand U7790 (N_7790,N_6456,N_6211);
and U7791 (N_7791,N_6689,N_6459);
or U7792 (N_7792,N_6276,N_6662);
and U7793 (N_7793,N_6030,N_6183);
xnor U7794 (N_7794,N_6900,N_6273);
or U7795 (N_7795,N_6667,N_6433);
or U7796 (N_7796,N_6248,N_6098);
and U7797 (N_7797,N_6520,N_6625);
nor U7798 (N_7798,N_6548,N_6899);
xor U7799 (N_7799,N_6693,N_6503);
xor U7800 (N_7800,N_6510,N_6535);
and U7801 (N_7801,N_6635,N_6182);
nor U7802 (N_7802,N_6600,N_6814);
or U7803 (N_7803,N_6522,N_6541);
and U7804 (N_7804,N_6089,N_6062);
xor U7805 (N_7805,N_6720,N_6419);
nor U7806 (N_7806,N_6092,N_6920);
xnor U7807 (N_7807,N_6500,N_6350);
nor U7808 (N_7808,N_6450,N_6515);
and U7809 (N_7809,N_6401,N_6822);
or U7810 (N_7810,N_6931,N_6010);
or U7811 (N_7811,N_6322,N_6691);
nor U7812 (N_7812,N_6727,N_6190);
or U7813 (N_7813,N_6234,N_6204);
xor U7814 (N_7814,N_6843,N_6398);
xor U7815 (N_7815,N_6551,N_6526);
xnor U7816 (N_7816,N_6775,N_6970);
nor U7817 (N_7817,N_6574,N_6102);
or U7818 (N_7818,N_6460,N_6756);
nor U7819 (N_7819,N_6044,N_6082);
or U7820 (N_7820,N_6882,N_6534);
or U7821 (N_7821,N_6706,N_6117);
nor U7822 (N_7822,N_6090,N_6093);
and U7823 (N_7823,N_6911,N_6233);
xnor U7824 (N_7824,N_6732,N_6133);
nand U7825 (N_7825,N_6658,N_6681);
xor U7826 (N_7826,N_6187,N_6089);
nand U7827 (N_7827,N_6498,N_6062);
nand U7828 (N_7828,N_6773,N_6198);
and U7829 (N_7829,N_6787,N_6740);
and U7830 (N_7830,N_6601,N_6718);
nand U7831 (N_7831,N_6603,N_6671);
and U7832 (N_7832,N_6916,N_6637);
and U7833 (N_7833,N_6505,N_6924);
xor U7834 (N_7834,N_6561,N_6656);
nor U7835 (N_7835,N_6104,N_6397);
nand U7836 (N_7836,N_6930,N_6754);
and U7837 (N_7837,N_6871,N_6520);
nor U7838 (N_7838,N_6784,N_6497);
nand U7839 (N_7839,N_6849,N_6938);
nand U7840 (N_7840,N_6358,N_6949);
and U7841 (N_7841,N_6424,N_6462);
xor U7842 (N_7842,N_6948,N_6894);
or U7843 (N_7843,N_6277,N_6921);
or U7844 (N_7844,N_6142,N_6215);
nor U7845 (N_7845,N_6091,N_6034);
or U7846 (N_7846,N_6673,N_6116);
nor U7847 (N_7847,N_6207,N_6632);
or U7848 (N_7848,N_6785,N_6896);
nor U7849 (N_7849,N_6796,N_6185);
and U7850 (N_7850,N_6354,N_6901);
nand U7851 (N_7851,N_6579,N_6349);
and U7852 (N_7852,N_6324,N_6800);
or U7853 (N_7853,N_6989,N_6092);
or U7854 (N_7854,N_6900,N_6140);
and U7855 (N_7855,N_6514,N_6927);
nand U7856 (N_7856,N_6125,N_6151);
nand U7857 (N_7857,N_6089,N_6786);
nand U7858 (N_7858,N_6492,N_6834);
and U7859 (N_7859,N_6417,N_6969);
xor U7860 (N_7860,N_6656,N_6062);
or U7861 (N_7861,N_6605,N_6172);
or U7862 (N_7862,N_6953,N_6066);
xor U7863 (N_7863,N_6073,N_6361);
or U7864 (N_7864,N_6174,N_6627);
or U7865 (N_7865,N_6103,N_6622);
nand U7866 (N_7866,N_6807,N_6396);
nand U7867 (N_7867,N_6033,N_6182);
and U7868 (N_7868,N_6656,N_6522);
xnor U7869 (N_7869,N_6709,N_6299);
and U7870 (N_7870,N_6977,N_6641);
or U7871 (N_7871,N_6862,N_6584);
and U7872 (N_7872,N_6860,N_6127);
or U7873 (N_7873,N_6882,N_6318);
nand U7874 (N_7874,N_6168,N_6546);
and U7875 (N_7875,N_6767,N_6934);
xor U7876 (N_7876,N_6814,N_6475);
nor U7877 (N_7877,N_6347,N_6195);
nor U7878 (N_7878,N_6557,N_6953);
or U7879 (N_7879,N_6945,N_6286);
and U7880 (N_7880,N_6963,N_6608);
nor U7881 (N_7881,N_6545,N_6147);
nand U7882 (N_7882,N_6927,N_6749);
nor U7883 (N_7883,N_6347,N_6800);
and U7884 (N_7884,N_6819,N_6691);
nand U7885 (N_7885,N_6502,N_6006);
nand U7886 (N_7886,N_6065,N_6419);
and U7887 (N_7887,N_6723,N_6613);
or U7888 (N_7888,N_6082,N_6095);
xor U7889 (N_7889,N_6517,N_6832);
nand U7890 (N_7890,N_6199,N_6606);
nor U7891 (N_7891,N_6233,N_6227);
nand U7892 (N_7892,N_6075,N_6743);
nand U7893 (N_7893,N_6247,N_6819);
nand U7894 (N_7894,N_6936,N_6944);
nand U7895 (N_7895,N_6370,N_6344);
or U7896 (N_7896,N_6458,N_6034);
xnor U7897 (N_7897,N_6073,N_6388);
xor U7898 (N_7898,N_6290,N_6960);
or U7899 (N_7899,N_6593,N_6577);
nand U7900 (N_7900,N_6878,N_6942);
and U7901 (N_7901,N_6797,N_6589);
and U7902 (N_7902,N_6249,N_6984);
nand U7903 (N_7903,N_6473,N_6656);
and U7904 (N_7904,N_6100,N_6447);
xnor U7905 (N_7905,N_6591,N_6088);
and U7906 (N_7906,N_6787,N_6489);
nor U7907 (N_7907,N_6762,N_6818);
nand U7908 (N_7908,N_6653,N_6695);
nand U7909 (N_7909,N_6880,N_6786);
xnor U7910 (N_7910,N_6822,N_6538);
or U7911 (N_7911,N_6622,N_6197);
or U7912 (N_7912,N_6905,N_6045);
and U7913 (N_7913,N_6038,N_6137);
and U7914 (N_7914,N_6540,N_6502);
nand U7915 (N_7915,N_6344,N_6284);
nand U7916 (N_7916,N_6290,N_6170);
and U7917 (N_7917,N_6557,N_6358);
nand U7918 (N_7918,N_6499,N_6966);
nor U7919 (N_7919,N_6861,N_6252);
nor U7920 (N_7920,N_6397,N_6650);
nor U7921 (N_7921,N_6182,N_6376);
and U7922 (N_7922,N_6525,N_6316);
nor U7923 (N_7923,N_6542,N_6573);
nor U7924 (N_7924,N_6696,N_6061);
nand U7925 (N_7925,N_6953,N_6231);
nand U7926 (N_7926,N_6124,N_6945);
xnor U7927 (N_7927,N_6336,N_6919);
nand U7928 (N_7928,N_6983,N_6317);
nor U7929 (N_7929,N_6102,N_6812);
xor U7930 (N_7930,N_6281,N_6058);
nand U7931 (N_7931,N_6348,N_6765);
xnor U7932 (N_7932,N_6369,N_6413);
nor U7933 (N_7933,N_6931,N_6441);
and U7934 (N_7934,N_6706,N_6762);
and U7935 (N_7935,N_6940,N_6159);
or U7936 (N_7936,N_6289,N_6328);
or U7937 (N_7937,N_6077,N_6827);
and U7938 (N_7938,N_6518,N_6505);
or U7939 (N_7939,N_6098,N_6756);
and U7940 (N_7940,N_6039,N_6511);
xnor U7941 (N_7941,N_6722,N_6480);
and U7942 (N_7942,N_6045,N_6231);
xnor U7943 (N_7943,N_6524,N_6854);
or U7944 (N_7944,N_6091,N_6966);
xnor U7945 (N_7945,N_6048,N_6375);
and U7946 (N_7946,N_6876,N_6905);
xnor U7947 (N_7947,N_6924,N_6742);
xor U7948 (N_7948,N_6311,N_6722);
nand U7949 (N_7949,N_6431,N_6162);
or U7950 (N_7950,N_6816,N_6625);
or U7951 (N_7951,N_6027,N_6171);
and U7952 (N_7952,N_6516,N_6147);
or U7953 (N_7953,N_6422,N_6913);
and U7954 (N_7954,N_6420,N_6874);
nor U7955 (N_7955,N_6740,N_6562);
xnor U7956 (N_7956,N_6955,N_6757);
nand U7957 (N_7957,N_6272,N_6795);
and U7958 (N_7958,N_6889,N_6082);
and U7959 (N_7959,N_6817,N_6707);
or U7960 (N_7960,N_6231,N_6952);
or U7961 (N_7961,N_6923,N_6083);
nand U7962 (N_7962,N_6492,N_6031);
nor U7963 (N_7963,N_6574,N_6257);
or U7964 (N_7964,N_6141,N_6414);
nand U7965 (N_7965,N_6836,N_6366);
nand U7966 (N_7966,N_6000,N_6323);
nand U7967 (N_7967,N_6998,N_6873);
or U7968 (N_7968,N_6641,N_6479);
and U7969 (N_7969,N_6487,N_6742);
nand U7970 (N_7970,N_6542,N_6472);
and U7971 (N_7971,N_6171,N_6074);
nand U7972 (N_7972,N_6321,N_6101);
xnor U7973 (N_7973,N_6341,N_6457);
and U7974 (N_7974,N_6706,N_6046);
and U7975 (N_7975,N_6631,N_6235);
nand U7976 (N_7976,N_6005,N_6103);
or U7977 (N_7977,N_6197,N_6339);
nand U7978 (N_7978,N_6828,N_6519);
xor U7979 (N_7979,N_6201,N_6673);
nor U7980 (N_7980,N_6063,N_6692);
xnor U7981 (N_7981,N_6836,N_6492);
and U7982 (N_7982,N_6706,N_6512);
and U7983 (N_7983,N_6623,N_6717);
nor U7984 (N_7984,N_6827,N_6916);
or U7985 (N_7985,N_6918,N_6525);
nand U7986 (N_7986,N_6105,N_6867);
nand U7987 (N_7987,N_6378,N_6321);
or U7988 (N_7988,N_6484,N_6524);
and U7989 (N_7989,N_6375,N_6404);
nand U7990 (N_7990,N_6722,N_6747);
xor U7991 (N_7991,N_6353,N_6960);
xnor U7992 (N_7992,N_6186,N_6829);
and U7993 (N_7993,N_6654,N_6344);
nand U7994 (N_7994,N_6386,N_6819);
and U7995 (N_7995,N_6226,N_6422);
or U7996 (N_7996,N_6058,N_6055);
nor U7997 (N_7997,N_6669,N_6532);
nand U7998 (N_7998,N_6039,N_6181);
xnor U7999 (N_7999,N_6886,N_6254);
and U8000 (N_8000,N_7409,N_7546);
nand U8001 (N_8001,N_7202,N_7833);
xor U8002 (N_8002,N_7304,N_7798);
nor U8003 (N_8003,N_7448,N_7857);
xnor U8004 (N_8004,N_7485,N_7818);
nor U8005 (N_8005,N_7559,N_7083);
xnor U8006 (N_8006,N_7901,N_7349);
and U8007 (N_8007,N_7960,N_7249);
nand U8008 (N_8008,N_7987,N_7912);
nand U8009 (N_8009,N_7514,N_7429);
nor U8010 (N_8010,N_7989,N_7804);
and U8011 (N_8011,N_7003,N_7434);
or U8012 (N_8012,N_7056,N_7288);
xor U8013 (N_8013,N_7408,N_7337);
nand U8014 (N_8014,N_7724,N_7879);
nand U8015 (N_8015,N_7175,N_7824);
and U8016 (N_8016,N_7159,N_7185);
or U8017 (N_8017,N_7432,N_7784);
nor U8018 (N_8018,N_7787,N_7872);
and U8019 (N_8019,N_7615,N_7803);
and U8020 (N_8020,N_7402,N_7771);
or U8021 (N_8021,N_7668,N_7186);
xor U8022 (N_8022,N_7767,N_7621);
nor U8023 (N_8023,N_7401,N_7384);
nand U8024 (N_8024,N_7358,N_7971);
and U8025 (N_8025,N_7550,N_7190);
nand U8026 (N_8026,N_7836,N_7555);
nor U8027 (N_8027,N_7160,N_7240);
xnor U8028 (N_8028,N_7831,N_7079);
or U8029 (N_8029,N_7498,N_7835);
xnor U8030 (N_8030,N_7925,N_7568);
nor U8031 (N_8031,N_7375,N_7501);
or U8032 (N_8032,N_7119,N_7379);
or U8033 (N_8033,N_7210,N_7755);
nor U8034 (N_8034,N_7863,N_7254);
nor U8035 (N_8035,N_7522,N_7627);
and U8036 (N_8036,N_7738,N_7947);
xor U8037 (N_8037,N_7101,N_7127);
xnor U8038 (N_8038,N_7759,N_7400);
nor U8039 (N_8039,N_7026,N_7045);
or U8040 (N_8040,N_7881,N_7839);
and U8041 (N_8041,N_7910,N_7195);
nand U8042 (N_8042,N_7601,N_7488);
nor U8043 (N_8043,N_7005,N_7543);
nand U8044 (N_8044,N_7880,N_7981);
nor U8045 (N_8045,N_7727,N_7091);
or U8046 (N_8046,N_7477,N_7343);
or U8047 (N_8047,N_7122,N_7878);
or U8048 (N_8048,N_7914,N_7952);
nand U8049 (N_8049,N_7469,N_7266);
xor U8050 (N_8050,N_7138,N_7310);
xor U8051 (N_8051,N_7636,N_7683);
nand U8052 (N_8052,N_7691,N_7532);
nand U8053 (N_8053,N_7526,N_7296);
or U8054 (N_8054,N_7271,N_7196);
xnor U8055 (N_8055,N_7723,N_7313);
nand U8056 (N_8056,N_7220,N_7499);
or U8057 (N_8057,N_7941,N_7157);
nand U8058 (N_8058,N_7070,N_7285);
nor U8059 (N_8059,N_7467,N_7199);
nand U8060 (N_8060,N_7335,N_7136);
or U8061 (N_8061,N_7184,N_7919);
or U8062 (N_8062,N_7648,N_7675);
nor U8063 (N_8063,N_7143,N_7012);
or U8064 (N_8064,N_7882,N_7242);
or U8065 (N_8065,N_7862,N_7694);
and U8066 (N_8066,N_7244,N_7896);
nor U8067 (N_8067,N_7877,N_7870);
and U8068 (N_8068,N_7782,N_7268);
or U8069 (N_8069,N_7311,N_7867);
nor U8070 (N_8070,N_7284,N_7339);
and U8071 (N_8071,N_7982,N_7654);
and U8072 (N_8072,N_7132,N_7376);
or U8073 (N_8073,N_7397,N_7735);
and U8074 (N_8074,N_7740,N_7355);
nand U8075 (N_8075,N_7347,N_7061);
nand U8076 (N_8076,N_7153,N_7687);
nand U8077 (N_8077,N_7680,N_7642);
or U8078 (N_8078,N_7608,N_7637);
and U8079 (N_8079,N_7262,N_7577);
xnor U8080 (N_8080,N_7991,N_7701);
xor U8081 (N_8081,N_7035,N_7055);
and U8082 (N_8082,N_7366,N_7998);
xnor U8083 (N_8083,N_7997,N_7676);
xor U8084 (N_8084,N_7093,N_7599);
and U8085 (N_8085,N_7293,N_7442);
xnor U8086 (N_8086,N_7886,N_7834);
and U8087 (N_8087,N_7068,N_7438);
nor U8088 (N_8088,N_7380,N_7523);
or U8089 (N_8089,N_7688,N_7123);
and U8090 (N_8090,N_7197,N_7367);
nor U8091 (N_8091,N_7507,N_7785);
nor U8092 (N_8092,N_7255,N_7893);
nor U8093 (N_8093,N_7086,N_7710);
or U8094 (N_8094,N_7425,N_7600);
and U8095 (N_8095,N_7796,N_7411);
nand U8096 (N_8096,N_7113,N_7643);
or U8097 (N_8097,N_7581,N_7351);
or U8098 (N_8098,N_7015,N_7576);
nand U8099 (N_8099,N_7606,N_7780);
nor U8100 (N_8100,N_7842,N_7243);
nor U8101 (N_8101,N_7452,N_7966);
xnor U8102 (N_8102,N_7146,N_7398);
nor U8103 (N_8103,N_7855,N_7126);
xnor U8104 (N_8104,N_7457,N_7161);
nor U8105 (N_8105,N_7923,N_7995);
xor U8106 (N_8106,N_7290,N_7742);
nand U8107 (N_8107,N_7547,N_7830);
nor U8108 (N_8108,N_7224,N_7214);
xnor U8109 (N_8109,N_7903,N_7921);
nor U8110 (N_8110,N_7926,N_7752);
or U8111 (N_8111,N_7010,N_7421);
nor U8112 (N_8112,N_7792,N_7625);
nand U8113 (N_8113,N_7825,N_7120);
xnor U8114 (N_8114,N_7321,N_7336);
nor U8115 (N_8115,N_7228,N_7149);
nor U8116 (N_8116,N_7595,N_7164);
or U8117 (N_8117,N_7038,N_7812);
xor U8118 (N_8118,N_7840,N_7279);
nor U8119 (N_8119,N_7813,N_7873);
nand U8120 (N_8120,N_7217,N_7042);
nor U8121 (N_8121,N_7482,N_7165);
or U8122 (N_8122,N_7890,N_7110);
nor U8123 (N_8123,N_7582,N_7536);
or U8124 (N_8124,N_7605,N_7907);
or U8125 (N_8125,N_7391,N_7588);
xor U8126 (N_8126,N_7297,N_7864);
nand U8127 (N_8127,N_7487,N_7282);
nand U8128 (N_8128,N_7406,N_7837);
or U8129 (N_8129,N_7418,N_7129);
and U8130 (N_8130,N_7585,N_7034);
nand U8131 (N_8131,N_7369,N_7150);
or U8132 (N_8132,N_7416,N_7639);
or U8133 (N_8133,N_7390,N_7117);
nand U8134 (N_8134,N_7078,N_7180);
and U8135 (N_8135,N_7235,N_7757);
nand U8136 (N_8136,N_7189,N_7898);
and U8137 (N_8137,N_7060,N_7081);
and U8138 (N_8138,N_7233,N_7392);
nor U8139 (N_8139,N_7647,N_7541);
xor U8140 (N_8140,N_7399,N_7428);
and U8141 (N_8141,N_7163,N_7763);
xnor U8142 (N_8142,N_7090,N_7631);
and U8143 (N_8143,N_7822,N_7385);
xnor U8144 (N_8144,N_7094,N_7871);
nand U8145 (N_8145,N_7578,N_7678);
and U8146 (N_8146,N_7455,N_7295);
or U8147 (N_8147,N_7371,N_7450);
nand U8148 (N_8148,N_7256,N_7373);
xnor U8149 (N_8149,N_7917,N_7407);
xnor U8150 (N_8150,N_7223,N_7427);
and U8151 (N_8151,N_7116,N_7561);
xnor U8152 (N_8152,N_7789,N_7974);
or U8153 (N_8153,N_7393,N_7460);
nor U8154 (N_8154,N_7325,N_7564);
and U8155 (N_8155,N_7490,N_7483);
nand U8156 (N_8156,N_7975,N_7350);
xor U8157 (N_8157,N_7883,N_7817);
nand U8158 (N_8158,N_7537,N_7622);
xor U8159 (N_8159,N_7732,N_7348);
and U8160 (N_8160,N_7506,N_7986);
and U8161 (N_8161,N_7492,N_7069);
or U8162 (N_8162,N_7875,N_7827);
and U8163 (N_8163,N_7811,N_7970);
xnor U8164 (N_8164,N_7772,N_7741);
and U8165 (N_8165,N_7044,N_7704);
and U8166 (N_8166,N_7207,N_7291);
xor U8167 (N_8167,N_7011,N_7019);
xnor U8168 (N_8168,N_7720,N_7059);
or U8169 (N_8169,N_7014,N_7978);
xnor U8170 (N_8170,N_7441,N_7632);
and U8171 (N_8171,N_7895,N_7505);
or U8172 (N_8172,N_7420,N_7041);
nand U8173 (N_8173,N_7151,N_7236);
or U8174 (N_8174,N_7023,N_7664);
nor U8175 (N_8175,N_7426,N_7072);
and U8176 (N_8176,N_7739,N_7712);
and U8177 (N_8177,N_7852,N_7649);
or U8178 (N_8178,N_7241,N_7865);
xnor U8179 (N_8179,N_7328,N_7264);
nor U8180 (N_8180,N_7777,N_7935);
nor U8181 (N_8181,N_7204,N_7359);
and U8182 (N_8182,N_7230,N_7762);
and U8183 (N_8183,N_7856,N_7203);
xor U8184 (N_8184,N_7048,N_7700);
nand U8185 (N_8185,N_7211,N_7128);
and U8186 (N_8186,N_7502,N_7414);
nand U8187 (N_8187,N_7612,N_7594);
and U8188 (N_8188,N_7580,N_7439);
nor U8189 (N_8189,N_7597,N_7037);
and U8190 (N_8190,N_7692,N_7690);
nor U8191 (N_8191,N_7171,N_7008);
and U8192 (N_8192,N_7449,N_7826);
nor U8193 (N_8193,N_7046,N_7586);
and U8194 (N_8194,N_7111,N_7481);
and U8195 (N_8195,N_7162,N_7112);
nor U8196 (N_8196,N_7212,N_7471);
nor U8197 (N_8197,N_7703,N_7509);
nand U8198 (N_8198,N_7959,N_7731);
nand U8199 (N_8199,N_7039,N_7693);
xnor U8200 (N_8200,N_7570,N_7965);
nor U8201 (N_8201,N_7031,N_7816);
or U8202 (N_8202,N_7948,N_7967);
xnor U8203 (N_8203,N_7334,N_7054);
xor U8204 (N_8204,N_7229,N_7629);
and U8205 (N_8205,N_7861,N_7462);
or U8206 (N_8206,N_7289,N_7372);
nor U8207 (N_8207,N_7567,N_7183);
and U8208 (N_8208,N_7277,N_7250);
and U8209 (N_8209,N_7954,N_7663);
xor U8210 (N_8210,N_7025,N_7064);
and U8211 (N_8211,N_7173,N_7618);
nor U8212 (N_8212,N_7135,N_7084);
and U8213 (N_8213,N_7247,N_7058);
and U8214 (N_8214,N_7307,N_7043);
and U8215 (N_8215,N_7918,N_7503);
xor U8216 (N_8216,N_7109,N_7556);
or U8217 (N_8217,N_7137,N_7049);
xnor U8218 (N_8218,N_7299,N_7177);
xnor U8219 (N_8219,N_7050,N_7098);
xor U8220 (N_8220,N_7144,N_7920);
or U8221 (N_8221,N_7294,N_7187);
nand U8222 (N_8222,N_7887,N_7658);
and U8223 (N_8223,N_7440,N_7188);
or U8224 (N_8224,N_7510,N_7800);
nand U8225 (N_8225,N_7340,N_7227);
and U8226 (N_8226,N_7669,N_7130);
nor U8227 (N_8227,N_7022,N_7644);
nand U8228 (N_8228,N_7333,N_7938);
or U8229 (N_8229,N_7718,N_7319);
and U8230 (N_8230,N_7105,N_7028);
xor U8231 (N_8231,N_7472,N_7215);
xor U8232 (N_8232,N_7200,N_7436);
nor U8233 (N_8233,N_7062,N_7681);
and U8234 (N_8234,N_7451,N_7354);
or U8235 (N_8235,N_7516,N_7844);
and U8236 (N_8236,N_7958,N_7222);
nor U8237 (N_8237,N_7972,N_7794);
and U8238 (N_8238,N_7029,N_7819);
nand U8239 (N_8239,N_7276,N_7733);
or U8240 (N_8240,N_7904,N_7134);
and U8241 (N_8241,N_7610,N_7006);
xor U8242 (N_8242,N_7362,N_7346);
nor U8243 (N_8243,N_7957,N_7040);
and U8244 (N_8244,N_7603,N_7659);
xnor U8245 (N_8245,N_7768,N_7820);
nor U8246 (N_8246,N_7067,N_7549);
nor U8247 (N_8247,N_7590,N_7706);
and U8248 (N_8248,N_7417,N_7237);
nor U8249 (N_8249,N_7773,N_7744);
nand U8250 (N_8250,N_7102,N_7626);
nand U8251 (N_8251,N_7140,N_7684);
nor U8252 (N_8252,N_7765,N_7057);
nor U8253 (N_8253,N_7308,N_7617);
xnor U8254 (N_8254,N_7774,N_7589);
xnor U8255 (N_8255,N_7650,N_7298);
xnor U8256 (N_8256,N_7121,N_7705);
nand U8257 (N_8257,N_7464,N_7540);
and U8258 (N_8258,N_7574,N_7095);
and U8259 (N_8259,N_7758,N_7066);
and U8260 (N_8260,N_7208,N_7182);
nor U8261 (N_8261,N_7990,N_7999);
and U8262 (N_8262,N_7446,N_7922);
nand U8263 (N_8263,N_7437,N_7695);
nor U8264 (N_8264,N_7531,N_7075);
nand U8265 (N_8265,N_7566,N_7345);
xnor U8266 (N_8266,N_7962,N_7232);
nand U8267 (N_8267,N_7623,N_7269);
and U8268 (N_8268,N_7248,N_7115);
xnor U8269 (N_8269,N_7716,N_7667);
and U8270 (N_8270,N_7553,N_7624);
and U8271 (N_8271,N_7021,N_7125);
xnor U8272 (N_8272,N_7992,N_7394);
nand U8273 (N_8273,N_7096,N_7341);
and U8274 (N_8274,N_7697,N_7013);
and U8275 (N_8275,N_7931,N_7107);
xor U8276 (N_8276,N_7360,N_7994);
xnor U8277 (N_8277,N_7497,N_7660);
xor U8278 (N_8278,N_7386,N_7430);
and U8279 (N_8279,N_7709,N_7571);
and U8280 (N_8280,N_7908,N_7943);
and U8281 (N_8281,N_7728,N_7076);
xor U8282 (N_8282,N_7403,N_7300);
nor U8283 (N_8283,N_7786,N_7662);
and U8284 (N_8284,N_7260,N_7641);
nor U8285 (N_8285,N_7218,N_7677);
or U8286 (N_8286,N_7829,N_7000);
or U8287 (N_8287,N_7329,N_7645);
or U8288 (N_8288,N_7737,N_7080);
or U8289 (N_8289,N_7906,N_7287);
or U8290 (N_8290,N_7486,N_7500);
and U8291 (N_8291,N_7572,N_7194);
xnor U8292 (N_8292,N_7719,N_7270);
nor U8293 (N_8293,N_7201,N_7097);
and U8294 (N_8294,N_7722,N_7365);
or U8295 (N_8295,N_7166,N_7356);
and U8296 (N_8296,N_7736,N_7009);
or U8297 (N_8297,N_7885,N_7283);
xnor U8298 (N_8298,N_7565,N_7924);
nor U8299 (N_8299,N_7963,N_7071);
or U8300 (N_8300,N_7979,N_7179);
or U8301 (N_8301,N_7527,N_7533);
or U8302 (N_8302,N_7431,N_7273);
and U8303 (N_8303,N_7281,N_7447);
xnor U8304 (N_8304,N_7213,N_7454);
or U8305 (N_8305,N_7301,N_7192);
nor U8306 (N_8306,N_7381,N_7751);
nor U8307 (N_8307,N_7828,N_7092);
xnor U8308 (N_8308,N_7653,N_7814);
or U8309 (N_8309,N_7776,N_7593);
xor U8310 (N_8310,N_7389,N_7944);
xor U8311 (N_8311,N_7030,N_7156);
and U8312 (N_8312,N_7953,N_7155);
nor U8313 (N_8313,N_7473,N_7051);
nor U8314 (N_8314,N_7239,N_7809);
xnor U8315 (N_8315,N_7916,N_7946);
nor U8316 (N_8316,N_7024,N_7118);
nand U8317 (N_8317,N_7114,N_7303);
nor U8318 (N_8318,N_7415,N_7172);
or U8319 (N_8319,N_7198,N_7387);
nand U8320 (N_8320,N_7754,N_7246);
nor U8321 (N_8321,N_7529,N_7205);
and U8322 (N_8322,N_7476,N_7843);
nand U8323 (N_8323,N_7475,N_7352);
nor U8324 (N_8324,N_7458,N_7638);
nand U8325 (N_8325,N_7193,N_7929);
and U8326 (N_8326,N_7725,N_7309);
xor U8327 (N_8327,N_7085,N_7364);
and U8328 (N_8328,N_7791,N_7563);
nor U8329 (N_8329,N_7750,N_7769);
or U8330 (N_8330,N_7363,N_7779);
or U8331 (N_8331,N_7463,N_7745);
nor U8332 (N_8332,N_7544,N_7849);
or U8333 (N_8333,N_7033,N_7656);
nand U8334 (N_8334,N_7783,N_7259);
nor U8335 (N_8335,N_7583,N_7717);
xnor U8336 (N_8336,N_7027,N_7322);
and U8337 (N_8337,N_7602,N_7592);
and U8338 (N_8338,N_7976,N_7484);
and U8339 (N_8339,N_7404,N_7221);
and U8340 (N_8340,N_7764,N_7479);
xnor U8341 (N_8341,N_7945,N_7884);
or U8342 (N_8342,N_7424,N_7939);
or U8343 (N_8343,N_7630,N_7474);
and U8344 (N_8344,N_7278,N_7145);
and U8345 (N_8345,N_7106,N_7573);
and U8346 (N_8346,N_7419,N_7848);
and U8347 (N_8347,N_7778,N_7410);
nor U8348 (N_8348,N_7614,N_7646);
or U8349 (N_8349,N_7263,N_7815);
or U8350 (N_8350,N_7802,N_7382);
and U8351 (N_8351,N_7805,N_7154);
or U8352 (N_8352,N_7152,N_7489);
and U8353 (N_8353,N_7730,N_7635);
and U8354 (N_8354,N_7951,N_7866);
and U8355 (N_8355,N_7357,N_7845);
nor U8356 (N_8356,N_7234,N_7461);
or U8357 (N_8357,N_7018,N_7673);
or U8358 (N_8358,N_7004,N_7504);
and U8359 (N_8359,N_7715,N_7558);
or U8360 (N_8360,N_7634,N_7374);
xor U8361 (N_8361,N_7591,N_7176);
or U8362 (N_8362,N_7616,N_7832);
or U8363 (N_8363,N_7859,N_7993);
nor U8364 (N_8364,N_7909,N_7074);
xnor U8365 (N_8365,N_7611,N_7928);
xor U8366 (N_8366,N_7726,N_7746);
or U8367 (N_8367,N_7721,N_7312);
or U8368 (N_8368,N_7405,N_7894);
and U8369 (N_8369,N_7219,N_7696);
nor U8370 (N_8370,N_7539,N_7370);
nor U8371 (N_8371,N_7930,N_7619);
or U8372 (N_8372,N_7760,N_7520);
xor U8373 (N_8373,N_7512,N_7496);
or U8374 (N_8374,N_7065,N_7913);
or U8375 (N_8375,N_7860,N_7748);
and U8376 (N_8376,N_7854,N_7983);
and U8377 (N_8377,N_7361,N_7891);
and U8378 (N_8378,N_7036,N_7032);
xor U8379 (N_8379,N_7331,N_7231);
or U8380 (N_8380,N_7324,N_7781);
or U8381 (N_8381,N_7478,N_7053);
and U8382 (N_8382,N_7465,N_7905);
or U8383 (N_8383,N_7554,N_7433);
or U8384 (N_8384,N_7897,N_7089);
nand U8385 (N_8385,N_7584,N_7560);
xor U8386 (N_8386,N_7797,N_7542);
nor U8387 (N_8387,N_7932,N_7142);
nor U8388 (N_8388,N_7342,N_7900);
nor U8389 (N_8389,N_7383,N_7412);
nor U8390 (N_8390,N_7950,N_7874);
nand U8391 (N_8391,N_7806,N_7139);
xor U8392 (N_8392,N_7468,N_7793);
nor U8393 (N_8393,N_7413,N_7655);
or U8394 (N_8394,N_7665,N_7444);
xnor U8395 (N_8395,N_7147,N_7657);
xor U8396 (N_8396,N_7206,N_7020);
nand U8397 (N_8397,N_7052,N_7749);
nand U8398 (N_8398,N_7002,N_7876);
and U8399 (N_8399,N_7823,N_7274);
or U8400 (N_8400,N_7911,N_7557);
xor U8401 (N_8401,N_7973,N_7168);
and U8402 (N_8402,N_7261,N_7521);
or U8403 (N_8403,N_7915,N_7082);
nor U8404 (N_8404,N_7332,N_7548);
xor U8405 (N_8405,N_7511,N_7265);
xnor U8406 (N_8406,N_7851,N_7170);
or U8407 (N_8407,N_7267,N_7853);
or U8408 (N_8408,N_7459,N_7985);
xnor U8409 (N_8409,N_7443,N_7178);
or U8410 (N_8410,N_7984,N_7524);
nand U8411 (N_8411,N_7395,N_7257);
and U8412 (N_8412,N_7988,N_7562);
nand U8413 (N_8413,N_7480,N_7258);
nand U8414 (N_8414,N_7810,N_7252);
or U8415 (N_8415,N_7686,N_7714);
nand U8416 (N_8416,N_7766,N_7315);
nand U8417 (N_8417,N_7934,N_7087);
xnor U8418 (N_8418,N_7933,N_7672);
or U8419 (N_8419,N_7552,N_7821);
and U8420 (N_8420,N_7167,N_7494);
xor U8421 (N_8421,N_7969,N_7850);
nand U8422 (N_8422,N_7841,N_7099);
xnor U8423 (N_8423,N_7598,N_7620);
or U8424 (N_8424,N_7869,N_7305);
nor U8425 (N_8425,N_7517,N_7679);
and U8426 (N_8426,N_7423,N_7302);
or U8427 (N_8427,N_7707,N_7747);
nand U8428 (N_8428,N_7317,N_7949);
nand U8429 (N_8429,N_7807,N_7902);
and U8430 (N_8430,N_7316,N_7569);
nand U8431 (N_8431,N_7661,N_7508);
or U8432 (N_8432,N_7579,N_7801);
and U8433 (N_8433,N_7702,N_7323);
nor U8434 (N_8434,N_7888,N_7330);
nor U8435 (N_8435,N_7513,N_7604);
or U8436 (N_8436,N_7551,N_7326);
nand U8437 (N_8437,N_7073,N_7158);
xor U8438 (N_8438,N_7209,N_7292);
nand U8439 (N_8439,N_7847,N_7734);
nor U8440 (N_8440,N_7396,N_7174);
and U8441 (N_8441,N_7937,N_7245);
and U8442 (N_8442,N_7613,N_7518);
nand U8443 (N_8443,N_7493,N_7216);
nor U8444 (N_8444,N_7596,N_7238);
or U8445 (N_8445,N_7148,N_7956);
nor U8446 (N_8446,N_7682,N_7191);
or U8447 (N_8447,N_7422,N_7977);
xor U8448 (N_8448,N_7689,N_7453);
and U8449 (N_8449,N_7708,N_7275);
nand U8450 (N_8450,N_7670,N_7133);
or U8451 (N_8451,N_7770,N_7108);
and U8452 (N_8452,N_7790,N_7280);
nand U8453 (N_8453,N_7515,N_7756);
xor U8454 (N_8454,N_7327,N_7698);
xor U8455 (N_8455,N_7713,N_7753);
nor U8456 (N_8456,N_7226,N_7955);
and U8457 (N_8457,N_7575,N_7124);
nand U8458 (N_8458,N_7338,N_7017);
and U8459 (N_8459,N_7699,N_7525);
and U8460 (N_8460,N_7927,N_7528);
xnor U8461 (N_8461,N_7251,N_7609);
nor U8462 (N_8462,N_7711,N_7942);
nand U8463 (N_8463,N_7651,N_7535);
xor U8464 (N_8464,N_7306,N_7491);
and U8465 (N_8465,N_7587,N_7470);
nor U8466 (N_8466,N_7799,N_7445);
or U8467 (N_8467,N_7495,N_7466);
and U8468 (N_8468,N_7685,N_7838);
xnor U8469 (N_8469,N_7940,N_7761);
xnor U8470 (N_8470,N_7225,N_7388);
nor U8471 (N_8471,N_7001,N_7980);
and U8472 (N_8472,N_7519,N_7936);
xnor U8473 (N_8473,N_7088,N_7344);
or U8474 (N_8474,N_7007,N_7743);
or U8475 (N_8475,N_7729,N_7253);
nand U8476 (N_8476,N_7545,N_7435);
and U8477 (N_8477,N_7846,N_7775);
nor U8478 (N_8478,N_7104,N_7378);
or U8479 (N_8479,N_7353,N_7534);
or U8480 (N_8480,N_7996,N_7795);
nand U8481 (N_8481,N_7181,N_7131);
nor U8482 (N_8482,N_7286,N_7169);
xor U8483 (N_8483,N_7538,N_7633);
nand U8484 (N_8484,N_7272,N_7666);
or U8485 (N_8485,N_7314,N_7858);
and U8486 (N_8486,N_7674,N_7889);
and U8487 (N_8487,N_7077,N_7964);
or U8488 (N_8488,N_7788,N_7899);
or U8489 (N_8489,N_7063,N_7892);
nor U8490 (N_8490,N_7808,N_7368);
nand U8491 (N_8491,N_7968,N_7016);
xnor U8492 (N_8492,N_7377,N_7607);
or U8493 (N_8493,N_7640,N_7103);
nand U8494 (N_8494,N_7628,N_7318);
or U8495 (N_8495,N_7047,N_7868);
nor U8496 (N_8496,N_7530,N_7671);
or U8497 (N_8497,N_7652,N_7456);
xnor U8498 (N_8498,N_7320,N_7100);
nand U8499 (N_8499,N_7141,N_7961);
and U8500 (N_8500,N_7383,N_7879);
or U8501 (N_8501,N_7755,N_7155);
or U8502 (N_8502,N_7996,N_7389);
or U8503 (N_8503,N_7670,N_7854);
nand U8504 (N_8504,N_7866,N_7949);
or U8505 (N_8505,N_7875,N_7820);
nor U8506 (N_8506,N_7392,N_7780);
xor U8507 (N_8507,N_7516,N_7745);
nand U8508 (N_8508,N_7123,N_7895);
nor U8509 (N_8509,N_7836,N_7887);
nand U8510 (N_8510,N_7315,N_7401);
nor U8511 (N_8511,N_7947,N_7771);
and U8512 (N_8512,N_7978,N_7667);
and U8513 (N_8513,N_7707,N_7526);
xnor U8514 (N_8514,N_7562,N_7376);
or U8515 (N_8515,N_7701,N_7913);
xnor U8516 (N_8516,N_7892,N_7425);
and U8517 (N_8517,N_7574,N_7289);
nor U8518 (N_8518,N_7633,N_7227);
and U8519 (N_8519,N_7932,N_7979);
and U8520 (N_8520,N_7953,N_7651);
nand U8521 (N_8521,N_7621,N_7365);
xor U8522 (N_8522,N_7944,N_7240);
nand U8523 (N_8523,N_7032,N_7548);
or U8524 (N_8524,N_7570,N_7547);
or U8525 (N_8525,N_7297,N_7403);
xnor U8526 (N_8526,N_7666,N_7702);
and U8527 (N_8527,N_7148,N_7321);
nor U8528 (N_8528,N_7320,N_7476);
nand U8529 (N_8529,N_7106,N_7872);
nand U8530 (N_8530,N_7265,N_7547);
xor U8531 (N_8531,N_7480,N_7742);
or U8532 (N_8532,N_7760,N_7883);
nand U8533 (N_8533,N_7384,N_7422);
nor U8534 (N_8534,N_7735,N_7479);
or U8535 (N_8535,N_7225,N_7833);
and U8536 (N_8536,N_7619,N_7586);
nand U8537 (N_8537,N_7895,N_7401);
and U8538 (N_8538,N_7690,N_7786);
nor U8539 (N_8539,N_7923,N_7639);
and U8540 (N_8540,N_7787,N_7251);
nor U8541 (N_8541,N_7111,N_7791);
nand U8542 (N_8542,N_7276,N_7272);
xnor U8543 (N_8543,N_7592,N_7459);
and U8544 (N_8544,N_7105,N_7360);
nand U8545 (N_8545,N_7703,N_7419);
and U8546 (N_8546,N_7900,N_7672);
nand U8547 (N_8547,N_7204,N_7999);
xnor U8548 (N_8548,N_7411,N_7742);
nand U8549 (N_8549,N_7412,N_7719);
and U8550 (N_8550,N_7625,N_7790);
nand U8551 (N_8551,N_7176,N_7815);
nand U8552 (N_8552,N_7141,N_7062);
xnor U8553 (N_8553,N_7877,N_7647);
nor U8554 (N_8554,N_7317,N_7203);
nand U8555 (N_8555,N_7123,N_7387);
nand U8556 (N_8556,N_7386,N_7006);
or U8557 (N_8557,N_7044,N_7670);
and U8558 (N_8558,N_7104,N_7173);
nor U8559 (N_8559,N_7636,N_7510);
xnor U8560 (N_8560,N_7193,N_7524);
or U8561 (N_8561,N_7606,N_7529);
nor U8562 (N_8562,N_7474,N_7987);
xor U8563 (N_8563,N_7834,N_7334);
xor U8564 (N_8564,N_7685,N_7845);
xor U8565 (N_8565,N_7746,N_7336);
and U8566 (N_8566,N_7348,N_7447);
or U8567 (N_8567,N_7253,N_7098);
nand U8568 (N_8568,N_7199,N_7932);
xor U8569 (N_8569,N_7628,N_7319);
nand U8570 (N_8570,N_7088,N_7026);
and U8571 (N_8571,N_7785,N_7970);
nor U8572 (N_8572,N_7657,N_7800);
and U8573 (N_8573,N_7906,N_7237);
nor U8574 (N_8574,N_7346,N_7743);
or U8575 (N_8575,N_7381,N_7561);
nor U8576 (N_8576,N_7226,N_7821);
and U8577 (N_8577,N_7403,N_7028);
xor U8578 (N_8578,N_7287,N_7534);
or U8579 (N_8579,N_7351,N_7830);
nand U8580 (N_8580,N_7864,N_7257);
xor U8581 (N_8581,N_7167,N_7936);
and U8582 (N_8582,N_7033,N_7947);
nor U8583 (N_8583,N_7128,N_7463);
nor U8584 (N_8584,N_7839,N_7549);
xor U8585 (N_8585,N_7838,N_7992);
or U8586 (N_8586,N_7494,N_7767);
and U8587 (N_8587,N_7974,N_7170);
or U8588 (N_8588,N_7527,N_7996);
nor U8589 (N_8589,N_7841,N_7166);
nand U8590 (N_8590,N_7976,N_7800);
or U8591 (N_8591,N_7205,N_7096);
nor U8592 (N_8592,N_7264,N_7061);
xnor U8593 (N_8593,N_7210,N_7731);
or U8594 (N_8594,N_7549,N_7863);
nand U8595 (N_8595,N_7258,N_7816);
nand U8596 (N_8596,N_7275,N_7811);
nor U8597 (N_8597,N_7409,N_7235);
and U8598 (N_8598,N_7596,N_7160);
nor U8599 (N_8599,N_7108,N_7288);
nand U8600 (N_8600,N_7639,N_7174);
nand U8601 (N_8601,N_7138,N_7128);
nor U8602 (N_8602,N_7215,N_7382);
nand U8603 (N_8603,N_7521,N_7440);
or U8604 (N_8604,N_7207,N_7024);
nand U8605 (N_8605,N_7210,N_7666);
xnor U8606 (N_8606,N_7870,N_7145);
or U8607 (N_8607,N_7409,N_7731);
or U8608 (N_8608,N_7562,N_7137);
nand U8609 (N_8609,N_7465,N_7772);
nand U8610 (N_8610,N_7935,N_7547);
nand U8611 (N_8611,N_7931,N_7174);
and U8612 (N_8612,N_7575,N_7063);
nand U8613 (N_8613,N_7046,N_7636);
or U8614 (N_8614,N_7943,N_7456);
or U8615 (N_8615,N_7785,N_7294);
and U8616 (N_8616,N_7072,N_7207);
and U8617 (N_8617,N_7470,N_7758);
nor U8618 (N_8618,N_7721,N_7424);
or U8619 (N_8619,N_7633,N_7961);
or U8620 (N_8620,N_7498,N_7044);
xor U8621 (N_8621,N_7374,N_7194);
or U8622 (N_8622,N_7671,N_7016);
nor U8623 (N_8623,N_7216,N_7691);
nor U8624 (N_8624,N_7893,N_7611);
xor U8625 (N_8625,N_7437,N_7211);
and U8626 (N_8626,N_7563,N_7494);
nand U8627 (N_8627,N_7345,N_7360);
nor U8628 (N_8628,N_7680,N_7794);
nor U8629 (N_8629,N_7941,N_7732);
nor U8630 (N_8630,N_7303,N_7899);
and U8631 (N_8631,N_7125,N_7128);
nand U8632 (N_8632,N_7018,N_7956);
or U8633 (N_8633,N_7354,N_7400);
nand U8634 (N_8634,N_7715,N_7147);
nand U8635 (N_8635,N_7209,N_7848);
and U8636 (N_8636,N_7572,N_7515);
nor U8637 (N_8637,N_7655,N_7103);
or U8638 (N_8638,N_7950,N_7308);
nand U8639 (N_8639,N_7885,N_7278);
nor U8640 (N_8640,N_7882,N_7933);
nand U8641 (N_8641,N_7806,N_7294);
and U8642 (N_8642,N_7425,N_7797);
xor U8643 (N_8643,N_7605,N_7629);
xor U8644 (N_8644,N_7774,N_7255);
nand U8645 (N_8645,N_7138,N_7725);
nand U8646 (N_8646,N_7550,N_7125);
xnor U8647 (N_8647,N_7161,N_7910);
nor U8648 (N_8648,N_7938,N_7608);
nand U8649 (N_8649,N_7412,N_7093);
xnor U8650 (N_8650,N_7575,N_7362);
and U8651 (N_8651,N_7481,N_7367);
nand U8652 (N_8652,N_7921,N_7562);
nand U8653 (N_8653,N_7942,N_7140);
and U8654 (N_8654,N_7132,N_7159);
nor U8655 (N_8655,N_7636,N_7203);
or U8656 (N_8656,N_7627,N_7074);
or U8657 (N_8657,N_7562,N_7608);
nor U8658 (N_8658,N_7141,N_7205);
nor U8659 (N_8659,N_7183,N_7405);
or U8660 (N_8660,N_7085,N_7771);
nand U8661 (N_8661,N_7413,N_7781);
xor U8662 (N_8662,N_7476,N_7705);
or U8663 (N_8663,N_7057,N_7966);
nor U8664 (N_8664,N_7173,N_7331);
nor U8665 (N_8665,N_7799,N_7869);
or U8666 (N_8666,N_7603,N_7703);
or U8667 (N_8667,N_7914,N_7926);
nor U8668 (N_8668,N_7239,N_7435);
or U8669 (N_8669,N_7930,N_7009);
xor U8670 (N_8670,N_7806,N_7697);
nand U8671 (N_8671,N_7828,N_7339);
xnor U8672 (N_8672,N_7677,N_7875);
or U8673 (N_8673,N_7667,N_7736);
nor U8674 (N_8674,N_7584,N_7729);
and U8675 (N_8675,N_7989,N_7348);
or U8676 (N_8676,N_7128,N_7254);
xor U8677 (N_8677,N_7529,N_7293);
and U8678 (N_8678,N_7236,N_7240);
nand U8679 (N_8679,N_7418,N_7833);
and U8680 (N_8680,N_7287,N_7612);
or U8681 (N_8681,N_7863,N_7558);
nor U8682 (N_8682,N_7938,N_7446);
nand U8683 (N_8683,N_7382,N_7148);
and U8684 (N_8684,N_7628,N_7332);
or U8685 (N_8685,N_7346,N_7845);
and U8686 (N_8686,N_7322,N_7456);
xor U8687 (N_8687,N_7149,N_7299);
nor U8688 (N_8688,N_7629,N_7392);
xnor U8689 (N_8689,N_7292,N_7515);
nor U8690 (N_8690,N_7785,N_7164);
or U8691 (N_8691,N_7997,N_7905);
and U8692 (N_8692,N_7921,N_7237);
and U8693 (N_8693,N_7606,N_7750);
nand U8694 (N_8694,N_7748,N_7900);
nor U8695 (N_8695,N_7143,N_7331);
and U8696 (N_8696,N_7118,N_7243);
nor U8697 (N_8697,N_7980,N_7724);
and U8698 (N_8698,N_7120,N_7690);
xnor U8699 (N_8699,N_7506,N_7744);
nand U8700 (N_8700,N_7581,N_7901);
nand U8701 (N_8701,N_7780,N_7706);
or U8702 (N_8702,N_7145,N_7668);
xnor U8703 (N_8703,N_7510,N_7475);
xor U8704 (N_8704,N_7959,N_7580);
or U8705 (N_8705,N_7246,N_7221);
and U8706 (N_8706,N_7046,N_7887);
xor U8707 (N_8707,N_7014,N_7710);
and U8708 (N_8708,N_7611,N_7153);
nand U8709 (N_8709,N_7344,N_7137);
nand U8710 (N_8710,N_7022,N_7451);
nor U8711 (N_8711,N_7391,N_7635);
and U8712 (N_8712,N_7618,N_7297);
nor U8713 (N_8713,N_7279,N_7876);
or U8714 (N_8714,N_7962,N_7359);
and U8715 (N_8715,N_7243,N_7499);
nor U8716 (N_8716,N_7916,N_7864);
or U8717 (N_8717,N_7039,N_7542);
xnor U8718 (N_8718,N_7830,N_7488);
nor U8719 (N_8719,N_7356,N_7129);
nor U8720 (N_8720,N_7136,N_7598);
or U8721 (N_8721,N_7570,N_7382);
xnor U8722 (N_8722,N_7391,N_7459);
xor U8723 (N_8723,N_7100,N_7180);
and U8724 (N_8724,N_7459,N_7231);
nor U8725 (N_8725,N_7074,N_7517);
xor U8726 (N_8726,N_7127,N_7634);
nand U8727 (N_8727,N_7872,N_7040);
or U8728 (N_8728,N_7329,N_7766);
and U8729 (N_8729,N_7978,N_7364);
nor U8730 (N_8730,N_7715,N_7891);
or U8731 (N_8731,N_7279,N_7863);
nor U8732 (N_8732,N_7870,N_7013);
nand U8733 (N_8733,N_7159,N_7484);
nor U8734 (N_8734,N_7361,N_7587);
xor U8735 (N_8735,N_7962,N_7821);
and U8736 (N_8736,N_7450,N_7729);
xnor U8737 (N_8737,N_7387,N_7347);
or U8738 (N_8738,N_7437,N_7639);
nor U8739 (N_8739,N_7706,N_7491);
nor U8740 (N_8740,N_7247,N_7539);
xnor U8741 (N_8741,N_7853,N_7737);
nand U8742 (N_8742,N_7666,N_7662);
or U8743 (N_8743,N_7012,N_7354);
nor U8744 (N_8744,N_7763,N_7498);
xnor U8745 (N_8745,N_7185,N_7740);
xnor U8746 (N_8746,N_7616,N_7146);
xnor U8747 (N_8747,N_7280,N_7699);
and U8748 (N_8748,N_7974,N_7940);
nand U8749 (N_8749,N_7049,N_7028);
nand U8750 (N_8750,N_7661,N_7480);
nand U8751 (N_8751,N_7274,N_7243);
nand U8752 (N_8752,N_7782,N_7925);
nor U8753 (N_8753,N_7778,N_7494);
nand U8754 (N_8754,N_7829,N_7036);
or U8755 (N_8755,N_7328,N_7796);
nor U8756 (N_8756,N_7085,N_7758);
xor U8757 (N_8757,N_7294,N_7515);
or U8758 (N_8758,N_7733,N_7723);
xor U8759 (N_8759,N_7203,N_7676);
xor U8760 (N_8760,N_7894,N_7063);
or U8761 (N_8761,N_7710,N_7885);
or U8762 (N_8762,N_7487,N_7444);
nand U8763 (N_8763,N_7795,N_7381);
nor U8764 (N_8764,N_7705,N_7533);
xnor U8765 (N_8765,N_7550,N_7740);
xor U8766 (N_8766,N_7251,N_7272);
xor U8767 (N_8767,N_7506,N_7951);
or U8768 (N_8768,N_7756,N_7364);
xnor U8769 (N_8769,N_7618,N_7310);
nor U8770 (N_8770,N_7683,N_7290);
xnor U8771 (N_8771,N_7872,N_7955);
and U8772 (N_8772,N_7117,N_7976);
and U8773 (N_8773,N_7046,N_7061);
and U8774 (N_8774,N_7998,N_7231);
nand U8775 (N_8775,N_7582,N_7955);
nor U8776 (N_8776,N_7259,N_7254);
nor U8777 (N_8777,N_7993,N_7503);
or U8778 (N_8778,N_7016,N_7192);
nor U8779 (N_8779,N_7100,N_7240);
or U8780 (N_8780,N_7674,N_7541);
nand U8781 (N_8781,N_7601,N_7706);
nand U8782 (N_8782,N_7414,N_7872);
nor U8783 (N_8783,N_7853,N_7387);
nor U8784 (N_8784,N_7047,N_7467);
nand U8785 (N_8785,N_7227,N_7042);
nor U8786 (N_8786,N_7246,N_7873);
nor U8787 (N_8787,N_7694,N_7132);
and U8788 (N_8788,N_7789,N_7343);
nand U8789 (N_8789,N_7373,N_7448);
nand U8790 (N_8790,N_7595,N_7509);
nor U8791 (N_8791,N_7578,N_7969);
nor U8792 (N_8792,N_7673,N_7437);
and U8793 (N_8793,N_7808,N_7637);
nand U8794 (N_8794,N_7285,N_7843);
and U8795 (N_8795,N_7196,N_7131);
xor U8796 (N_8796,N_7123,N_7304);
or U8797 (N_8797,N_7235,N_7311);
or U8798 (N_8798,N_7383,N_7692);
and U8799 (N_8799,N_7371,N_7850);
nand U8800 (N_8800,N_7772,N_7241);
nor U8801 (N_8801,N_7773,N_7835);
and U8802 (N_8802,N_7302,N_7327);
and U8803 (N_8803,N_7808,N_7018);
nand U8804 (N_8804,N_7262,N_7265);
nand U8805 (N_8805,N_7831,N_7630);
and U8806 (N_8806,N_7164,N_7319);
and U8807 (N_8807,N_7463,N_7490);
and U8808 (N_8808,N_7370,N_7033);
or U8809 (N_8809,N_7379,N_7847);
nand U8810 (N_8810,N_7581,N_7345);
or U8811 (N_8811,N_7413,N_7247);
or U8812 (N_8812,N_7822,N_7749);
nor U8813 (N_8813,N_7529,N_7851);
and U8814 (N_8814,N_7830,N_7226);
or U8815 (N_8815,N_7028,N_7900);
nand U8816 (N_8816,N_7152,N_7170);
and U8817 (N_8817,N_7410,N_7587);
or U8818 (N_8818,N_7209,N_7783);
and U8819 (N_8819,N_7283,N_7098);
or U8820 (N_8820,N_7612,N_7552);
nor U8821 (N_8821,N_7648,N_7708);
xor U8822 (N_8822,N_7081,N_7660);
nand U8823 (N_8823,N_7322,N_7114);
nand U8824 (N_8824,N_7561,N_7388);
and U8825 (N_8825,N_7316,N_7339);
nand U8826 (N_8826,N_7395,N_7595);
nor U8827 (N_8827,N_7821,N_7887);
or U8828 (N_8828,N_7067,N_7317);
nand U8829 (N_8829,N_7531,N_7998);
nand U8830 (N_8830,N_7236,N_7956);
nand U8831 (N_8831,N_7092,N_7338);
or U8832 (N_8832,N_7412,N_7708);
nor U8833 (N_8833,N_7142,N_7217);
xor U8834 (N_8834,N_7785,N_7580);
and U8835 (N_8835,N_7791,N_7306);
nand U8836 (N_8836,N_7162,N_7977);
and U8837 (N_8837,N_7553,N_7876);
or U8838 (N_8838,N_7752,N_7591);
nor U8839 (N_8839,N_7731,N_7765);
or U8840 (N_8840,N_7978,N_7190);
and U8841 (N_8841,N_7917,N_7591);
nand U8842 (N_8842,N_7505,N_7309);
or U8843 (N_8843,N_7776,N_7980);
and U8844 (N_8844,N_7218,N_7095);
nand U8845 (N_8845,N_7239,N_7595);
nor U8846 (N_8846,N_7442,N_7765);
xor U8847 (N_8847,N_7879,N_7910);
nand U8848 (N_8848,N_7715,N_7956);
nand U8849 (N_8849,N_7040,N_7844);
xnor U8850 (N_8850,N_7884,N_7790);
nor U8851 (N_8851,N_7755,N_7814);
xor U8852 (N_8852,N_7201,N_7278);
xor U8853 (N_8853,N_7860,N_7616);
nand U8854 (N_8854,N_7389,N_7777);
nor U8855 (N_8855,N_7392,N_7078);
xor U8856 (N_8856,N_7333,N_7076);
xnor U8857 (N_8857,N_7811,N_7322);
nor U8858 (N_8858,N_7718,N_7703);
nor U8859 (N_8859,N_7270,N_7480);
or U8860 (N_8860,N_7502,N_7785);
or U8861 (N_8861,N_7942,N_7549);
xor U8862 (N_8862,N_7632,N_7823);
nor U8863 (N_8863,N_7033,N_7412);
xor U8864 (N_8864,N_7360,N_7840);
nor U8865 (N_8865,N_7203,N_7073);
xnor U8866 (N_8866,N_7676,N_7613);
nand U8867 (N_8867,N_7392,N_7455);
or U8868 (N_8868,N_7365,N_7201);
xor U8869 (N_8869,N_7462,N_7799);
nor U8870 (N_8870,N_7838,N_7665);
or U8871 (N_8871,N_7262,N_7893);
or U8872 (N_8872,N_7809,N_7281);
and U8873 (N_8873,N_7141,N_7812);
nand U8874 (N_8874,N_7004,N_7424);
nand U8875 (N_8875,N_7446,N_7694);
nor U8876 (N_8876,N_7527,N_7178);
or U8877 (N_8877,N_7350,N_7633);
and U8878 (N_8878,N_7208,N_7334);
xor U8879 (N_8879,N_7459,N_7084);
nor U8880 (N_8880,N_7100,N_7659);
nor U8881 (N_8881,N_7131,N_7925);
and U8882 (N_8882,N_7057,N_7876);
nor U8883 (N_8883,N_7385,N_7007);
nor U8884 (N_8884,N_7101,N_7498);
nand U8885 (N_8885,N_7137,N_7780);
xnor U8886 (N_8886,N_7160,N_7027);
and U8887 (N_8887,N_7860,N_7242);
nand U8888 (N_8888,N_7548,N_7095);
nor U8889 (N_8889,N_7367,N_7831);
nor U8890 (N_8890,N_7275,N_7199);
and U8891 (N_8891,N_7804,N_7004);
or U8892 (N_8892,N_7277,N_7676);
xor U8893 (N_8893,N_7182,N_7025);
xor U8894 (N_8894,N_7753,N_7251);
xnor U8895 (N_8895,N_7855,N_7573);
xnor U8896 (N_8896,N_7473,N_7469);
nand U8897 (N_8897,N_7164,N_7146);
nor U8898 (N_8898,N_7518,N_7094);
and U8899 (N_8899,N_7006,N_7093);
nor U8900 (N_8900,N_7287,N_7711);
nor U8901 (N_8901,N_7512,N_7250);
nor U8902 (N_8902,N_7485,N_7027);
xnor U8903 (N_8903,N_7001,N_7101);
or U8904 (N_8904,N_7748,N_7617);
nand U8905 (N_8905,N_7883,N_7780);
and U8906 (N_8906,N_7538,N_7733);
or U8907 (N_8907,N_7936,N_7029);
or U8908 (N_8908,N_7562,N_7207);
nand U8909 (N_8909,N_7260,N_7658);
and U8910 (N_8910,N_7218,N_7512);
and U8911 (N_8911,N_7356,N_7566);
nor U8912 (N_8912,N_7252,N_7070);
xnor U8913 (N_8913,N_7632,N_7820);
and U8914 (N_8914,N_7176,N_7144);
nor U8915 (N_8915,N_7542,N_7873);
nand U8916 (N_8916,N_7104,N_7000);
nor U8917 (N_8917,N_7321,N_7551);
or U8918 (N_8918,N_7415,N_7942);
nand U8919 (N_8919,N_7856,N_7142);
nand U8920 (N_8920,N_7654,N_7656);
nand U8921 (N_8921,N_7734,N_7125);
nor U8922 (N_8922,N_7522,N_7835);
nor U8923 (N_8923,N_7445,N_7779);
nor U8924 (N_8924,N_7613,N_7358);
xnor U8925 (N_8925,N_7711,N_7069);
nand U8926 (N_8926,N_7247,N_7566);
nand U8927 (N_8927,N_7595,N_7894);
nor U8928 (N_8928,N_7014,N_7350);
or U8929 (N_8929,N_7179,N_7089);
and U8930 (N_8930,N_7769,N_7614);
nand U8931 (N_8931,N_7402,N_7553);
xor U8932 (N_8932,N_7501,N_7031);
or U8933 (N_8933,N_7738,N_7281);
nor U8934 (N_8934,N_7358,N_7742);
and U8935 (N_8935,N_7383,N_7320);
nor U8936 (N_8936,N_7473,N_7617);
xnor U8937 (N_8937,N_7392,N_7901);
nand U8938 (N_8938,N_7296,N_7697);
and U8939 (N_8939,N_7958,N_7304);
xor U8940 (N_8940,N_7237,N_7569);
and U8941 (N_8941,N_7873,N_7520);
nor U8942 (N_8942,N_7879,N_7979);
and U8943 (N_8943,N_7822,N_7184);
and U8944 (N_8944,N_7967,N_7500);
nor U8945 (N_8945,N_7970,N_7003);
nand U8946 (N_8946,N_7226,N_7613);
or U8947 (N_8947,N_7196,N_7146);
nor U8948 (N_8948,N_7185,N_7903);
nor U8949 (N_8949,N_7089,N_7315);
nand U8950 (N_8950,N_7101,N_7035);
nand U8951 (N_8951,N_7596,N_7031);
and U8952 (N_8952,N_7741,N_7845);
and U8953 (N_8953,N_7109,N_7437);
nand U8954 (N_8954,N_7550,N_7404);
or U8955 (N_8955,N_7951,N_7054);
nand U8956 (N_8956,N_7569,N_7046);
nor U8957 (N_8957,N_7848,N_7895);
nand U8958 (N_8958,N_7183,N_7352);
or U8959 (N_8959,N_7250,N_7291);
and U8960 (N_8960,N_7717,N_7542);
and U8961 (N_8961,N_7276,N_7591);
and U8962 (N_8962,N_7141,N_7077);
and U8963 (N_8963,N_7241,N_7265);
xor U8964 (N_8964,N_7887,N_7258);
and U8965 (N_8965,N_7814,N_7409);
or U8966 (N_8966,N_7548,N_7019);
xor U8967 (N_8967,N_7837,N_7997);
nand U8968 (N_8968,N_7741,N_7405);
nor U8969 (N_8969,N_7573,N_7772);
xnor U8970 (N_8970,N_7442,N_7374);
nand U8971 (N_8971,N_7973,N_7443);
nor U8972 (N_8972,N_7082,N_7952);
nand U8973 (N_8973,N_7098,N_7529);
or U8974 (N_8974,N_7606,N_7799);
or U8975 (N_8975,N_7324,N_7978);
nor U8976 (N_8976,N_7858,N_7531);
and U8977 (N_8977,N_7128,N_7835);
or U8978 (N_8978,N_7866,N_7132);
and U8979 (N_8979,N_7932,N_7772);
nor U8980 (N_8980,N_7787,N_7738);
and U8981 (N_8981,N_7393,N_7542);
nand U8982 (N_8982,N_7822,N_7909);
xor U8983 (N_8983,N_7984,N_7278);
and U8984 (N_8984,N_7968,N_7620);
or U8985 (N_8985,N_7528,N_7546);
nand U8986 (N_8986,N_7939,N_7090);
nor U8987 (N_8987,N_7288,N_7721);
xnor U8988 (N_8988,N_7843,N_7542);
nor U8989 (N_8989,N_7487,N_7929);
nor U8990 (N_8990,N_7366,N_7140);
or U8991 (N_8991,N_7106,N_7702);
nand U8992 (N_8992,N_7931,N_7998);
xnor U8993 (N_8993,N_7399,N_7893);
or U8994 (N_8994,N_7808,N_7674);
nor U8995 (N_8995,N_7756,N_7755);
or U8996 (N_8996,N_7165,N_7822);
or U8997 (N_8997,N_7444,N_7049);
and U8998 (N_8998,N_7329,N_7268);
nand U8999 (N_8999,N_7299,N_7368);
or U9000 (N_9000,N_8854,N_8182);
nand U9001 (N_9001,N_8198,N_8493);
nand U9002 (N_9002,N_8266,N_8974);
or U9003 (N_9003,N_8385,N_8552);
xor U9004 (N_9004,N_8861,N_8500);
and U9005 (N_9005,N_8446,N_8807);
nor U9006 (N_9006,N_8509,N_8549);
or U9007 (N_9007,N_8192,N_8325);
nand U9008 (N_9008,N_8047,N_8629);
and U9009 (N_9009,N_8135,N_8515);
xnor U9010 (N_9010,N_8568,N_8508);
nor U9011 (N_9011,N_8819,N_8153);
nor U9012 (N_9012,N_8659,N_8248);
or U9013 (N_9013,N_8028,N_8981);
or U9014 (N_9014,N_8742,N_8187);
or U9015 (N_9015,N_8563,N_8285);
xnor U9016 (N_9016,N_8338,N_8801);
nor U9017 (N_9017,N_8494,N_8214);
xnor U9018 (N_9018,N_8103,N_8776);
nand U9019 (N_9019,N_8816,N_8840);
and U9020 (N_9020,N_8989,N_8298);
nor U9021 (N_9021,N_8792,N_8590);
nor U9022 (N_9022,N_8738,N_8421);
nand U9023 (N_9023,N_8276,N_8995);
and U9024 (N_9024,N_8530,N_8513);
and U9025 (N_9025,N_8420,N_8583);
nand U9026 (N_9026,N_8404,N_8955);
xnor U9027 (N_9027,N_8617,N_8875);
xor U9028 (N_9028,N_8039,N_8966);
nand U9029 (N_9029,N_8473,N_8667);
xor U9030 (N_9030,N_8829,N_8180);
and U9031 (N_9031,N_8706,N_8841);
xnor U9032 (N_9032,N_8979,N_8081);
nand U9033 (N_9033,N_8964,N_8274);
nor U9034 (N_9034,N_8114,N_8394);
xor U9035 (N_9035,N_8315,N_8949);
nand U9036 (N_9036,N_8911,N_8741);
nand U9037 (N_9037,N_8519,N_8167);
nor U9038 (N_9038,N_8049,N_8621);
nand U9039 (N_9039,N_8517,N_8605);
and U9040 (N_9040,N_8104,N_8710);
and U9041 (N_9041,N_8693,N_8270);
and U9042 (N_9042,N_8747,N_8258);
nand U9043 (N_9043,N_8092,N_8306);
or U9044 (N_9044,N_8053,N_8439);
and U9045 (N_9045,N_8123,N_8579);
nand U9046 (N_9046,N_8392,N_8040);
xor U9047 (N_9047,N_8926,N_8284);
xor U9048 (N_9048,N_8928,N_8880);
or U9049 (N_9049,N_8287,N_8072);
nor U9050 (N_9050,N_8891,N_8112);
nor U9051 (N_9051,N_8698,N_8416);
and U9052 (N_9052,N_8189,N_8497);
or U9053 (N_9053,N_8041,N_8814);
or U9054 (N_9054,N_8598,N_8227);
xor U9055 (N_9055,N_8260,N_8254);
or U9056 (N_9056,N_8312,N_8538);
or U9057 (N_9057,N_8600,N_8946);
nor U9058 (N_9058,N_8899,N_8570);
nand U9059 (N_9059,N_8119,N_8753);
xor U9060 (N_9060,N_8060,N_8435);
or U9061 (N_9061,N_8997,N_8217);
xnor U9062 (N_9062,N_8585,N_8384);
or U9063 (N_9063,N_8407,N_8499);
nor U9064 (N_9064,N_8761,N_8272);
nand U9065 (N_9065,N_8280,N_8987);
and U9066 (N_9066,N_8098,N_8766);
xnor U9067 (N_9067,N_8471,N_8190);
and U9068 (N_9068,N_8476,N_8418);
and U9069 (N_9069,N_8111,N_8878);
nand U9070 (N_9070,N_8925,N_8842);
xor U9071 (N_9071,N_8464,N_8457);
nand U9072 (N_9072,N_8614,N_8342);
and U9073 (N_9073,N_8046,N_8283);
nor U9074 (N_9074,N_8310,N_8063);
and U9075 (N_9075,N_8122,N_8799);
or U9076 (N_9076,N_8003,N_8376);
and U9077 (N_9077,N_8129,N_8514);
xnor U9078 (N_9078,N_8662,N_8012);
nand U9079 (N_9079,N_8822,N_8296);
xor U9080 (N_9080,N_8375,N_8004);
xnor U9081 (N_9081,N_8580,N_8474);
xor U9082 (N_9082,N_8690,N_8212);
xor U9083 (N_9083,N_8133,N_8820);
nand U9084 (N_9084,N_8085,N_8870);
or U9085 (N_9085,N_8851,N_8145);
xor U9086 (N_9086,N_8898,N_8152);
or U9087 (N_9087,N_8771,N_8030);
nor U9088 (N_9088,N_8429,N_8055);
nand U9089 (N_9089,N_8548,N_8383);
and U9090 (N_9090,N_8329,N_8764);
and U9091 (N_9091,N_8064,N_8166);
and U9092 (N_9092,N_8239,N_8358);
and U9093 (N_9093,N_8139,N_8466);
nand U9094 (N_9094,N_8666,N_8589);
xor U9095 (N_9095,N_8998,N_8709);
or U9096 (N_9096,N_8909,N_8923);
xnor U9097 (N_9097,N_8467,N_8916);
xnor U9098 (N_9098,N_8451,N_8365);
and U9099 (N_9099,N_8843,N_8594);
xnor U9100 (N_9100,N_8827,N_8089);
and U9101 (N_9101,N_8197,N_8795);
nor U9102 (N_9102,N_8784,N_8551);
nor U9103 (N_9103,N_8014,N_8218);
and U9104 (N_9104,N_8186,N_8951);
nand U9105 (N_9105,N_8204,N_8252);
or U9106 (N_9106,N_8890,N_8953);
and U9107 (N_9107,N_8045,N_8815);
nor U9108 (N_9108,N_8224,N_8381);
nor U9109 (N_9109,N_8729,N_8701);
or U9110 (N_9110,N_8026,N_8165);
nand U9111 (N_9111,N_8007,N_8456);
or U9112 (N_9112,N_8522,N_8846);
nand U9113 (N_9113,N_8199,N_8351);
nand U9114 (N_9114,N_8452,N_8751);
nor U9115 (N_9115,N_8606,N_8770);
nor U9116 (N_9116,N_8582,N_8255);
xor U9117 (N_9117,N_8531,N_8147);
xor U9118 (N_9118,N_8685,N_8632);
and U9119 (N_9119,N_8765,N_8141);
xnor U9120 (N_9120,N_8733,N_8148);
xnor U9121 (N_9121,N_8712,N_8347);
nand U9122 (N_9122,N_8194,N_8249);
xor U9123 (N_9123,N_8626,N_8566);
nand U9124 (N_9124,N_8087,N_8825);
xnor U9125 (N_9125,N_8279,N_8431);
nor U9126 (N_9126,N_8311,N_8893);
nor U9127 (N_9127,N_8286,N_8316);
or U9128 (N_9128,N_8859,N_8554);
and U9129 (N_9129,N_8475,N_8631);
nand U9130 (N_9130,N_8688,N_8382);
and U9131 (N_9131,N_8495,N_8162);
nand U9132 (N_9132,N_8716,N_8798);
xnor U9133 (N_9133,N_8211,N_8427);
and U9134 (N_9134,N_8541,N_8930);
or U9135 (N_9135,N_8806,N_8038);
nor U9136 (N_9136,N_8897,N_8093);
nand U9137 (N_9137,N_8232,N_8663);
and U9138 (N_9138,N_8561,N_8453);
or U9139 (N_9139,N_8426,N_8086);
and U9140 (N_9140,N_8939,N_8067);
and U9141 (N_9141,N_8571,N_8116);
or U9142 (N_9142,N_8529,N_8869);
xnor U9143 (N_9143,N_8425,N_8247);
nor U9144 (N_9144,N_8924,N_8216);
or U9145 (N_9145,N_8313,N_8993);
or U9146 (N_9146,N_8967,N_8892);
and U9147 (N_9147,N_8990,N_8374);
nor U9148 (N_9148,N_8331,N_8683);
and U9149 (N_9149,N_8436,N_8082);
xnor U9150 (N_9150,N_8718,N_8095);
nand U9151 (N_9151,N_8137,N_8231);
nor U9152 (N_9152,N_8428,N_8944);
and U9153 (N_9153,N_8389,N_8681);
or U9154 (N_9154,N_8671,N_8945);
nand U9155 (N_9155,N_8948,N_8547);
nand U9156 (N_9156,N_8482,N_8001);
or U9157 (N_9157,N_8235,N_8936);
xnor U9158 (N_9158,N_8128,N_8678);
nor U9159 (N_9159,N_8088,N_8660);
or U9160 (N_9160,N_8542,N_8059);
xor U9161 (N_9161,N_8206,N_8447);
and U9162 (N_9162,N_8968,N_8615);
or U9163 (N_9163,N_8174,N_8492);
nor U9164 (N_9164,N_8171,N_8895);
or U9165 (N_9165,N_8833,N_8503);
nand U9166 (N_9166,N_8868,N_8469);
or U9167 (N_9167,N_8151,N_8734);
nor U9168 (N_9168,N_8543,N_8303);
nor U9169 (N_9169,N_8346,N_8609);
or U9170 (N_9170,N_8448,N_8483);
nor U9171 (N_9171,N_8886,N_8942);
or U9172 (N_9172,N_8654,N_8149);
nand U9173 (N_9173,N_8648,N_8917);
xor U9174 (N_9174,N_8633,N_8324);
or U9175 (N_9175,N_8022,N_8177);
and U9176 (N_9176,N_8762,N_8835);
and U9177 (N_9177,N_8818,N_8752);
xnor U9178 (N_9178,N_8649,N_8083);
nor U9179 (N_9179,N_8411,N_8188);
nand U9180 (N_9180,N_8226,N_8750);
nor U9181 (N_9181,N_8973,N_8535);
xnor U9182 (N_9182,N_8322,N_8941);
nand U9183 (N_9183,N_8763,N_8512);
nand U9184 (N_9184,N_8146,N_8019);
xor U9185 (N_9185,N_8443,N_8257);
nand U9186 (N_9186,N_8319,N_8159);
nand U9187 (N_9187,N_8777,N_8277);
xnor U9188 (N_9188,N_8700,N_8246);
and U9189 (N_9189,N_8921,N_8341);
nor U9190 (N_9190,N_8075,N_8970);
nor U9191 (N_9191,N_8545,N_8449);
and U9192 (N_9192,N_8574,N_8772);
or U9193 (N_9193,N_8677,N_8321);
nor U9194 (N_9194,N_8963,N_8544);
xor U9195 (N_9195,N_8101,N_8757);
xor U9196 (N_9196,N_8386,N_8525);
nand U9197 (N_9197,N_8785,N_8702);
xor U9198 (N_9198,N_8242,N_8403);
and U9199 (N_9199,N_8077,N_8220);
xnor U9200 (N_9200,N_8913,N_8540);
nand U9201 (N_9201,N_8823,N_8789);
nand U9202 (N_9202,N_8713,N_8359);
nor U9203 (N_9203,N_8269,N_8243);
xnor U9204 (N_9204,N_8048,N_8097);
xor U9205 (N_9205,N_8985,N_8811);
and U9206 (N_9206,N_8790,N_8442);
and U9207 (N_9207,N_8947,N_8644);
nor U9208 (N_9208,N_8971,N_8488);
xor U9209 (N_9209,N_8692,N_8179);
and U9210 (N_9210,N_8185,N_8783);
xnor U9211 (N_9211,N_8694,N_8664);
or U9212 (N_9212,N_8908,N_8641);
or U9213 (N_9213,N_8069,N_8441);
nor U9214 (N_9214,N_8595,N_8665);
and U9215 (N_9215,N_8876,N_8355);
nand U9216 (N_9216,N_8658,N_8202);
nand U9217 (N_9217,N_8016,N_8134);
nand U9218 (N_9218,N_8929,N_8352);
or U9219 (N_9219,N_8309,N_8193);
and U9220 (N_9220,N_8491,N_8651);
nand U9221 (N_9221,N_8465,N_8630);
nor U9222 (N_9222,N_8972,N_8068);
xnor U9223 (N_9223,N_8900,N_8366);
nor U9224 (N_9224,N_8914,N_8977);
nor U9225 (N_9225,N_8035,N_8364);
nor U9226 (N_9226,N_8424,N_8720);
and U9227 (N_9227,N_8136,N_8760);
nor U9228 (N_9228,N_8830,N_8506);
nand U9229 (N_9229,N_8345,N_8219);
or U9230 (N_9230,N_8699,N_8066);
xnor U9231 (N_9231,N_8956,N_8697);
nor U9232 (N_9232,N_8334,N_8959);
xor U9233 (N_9233,N_8797,N_8323);
or U9234 (N_9234,N_8412,N_8740);
xor U9235 (N_9235,N_8078,N_8031);
or U9236 (N_9236,N_8071,N_8826);
nand U9237 (N_9237,N_8935,N_8486);
and U9238 (N_9238,N_8652,N_8691);
or U9239 (N_9239,N_8577,N_8587);
nor U9240 (N_9240,N_8213,N_8100);
nor U9241 (N_9241,N_8050,N_8802);
nor U9242 (N_9242,N_8839,N_8481);
or U9243 (N_9243,N_8578,N_8743);
and U9244 (N_9244,N_8504,N_8268);
xnor U9245 (N_9245,N_8767,N_8521);
xnor U9246 (N_9246,N_8518,N_8236);
and U9247 (N_9247,N_8314,N_8639);
nor U9248 (N_9248,N_8749,N_8222);
and U9249 (N_9249,N_8264,N_8330);
nor U9250 (N_9250,N_8675,N_8592);
nor U9251 (N_9251,N_8455,N_8960);
or U9252 (N_9252,N_8430,N_8943);
nand U9253 (N_9253,N_8724,N_8477);
xor U9254 (N_9254,N_8907,N_8154);
nand U9255 (N_9255,N_8417,N_8808);
and U9256 (N_9256,N_8857,N_8550);
xnor U9257 (N_9257,N_8986,N_8965);
or U9258 (N_9258,N_8882,N_8599);
or U9259 (N_9259,N_8670,N_8295);
nor U9260 (N_9260,N_8335,N_8118);
nor U9261 (N_9261,N_8461,N_8824);
xor U9262 (N_9262,N_8395,N_8327);
xor U9263 (N_9263,N_8237,N_8793);
nor U9264 (N_9264,N_8668,N_8360);
nand U9265 (N_9265,N_8608,N_8132);
nor U9266 (N_9266,N_8127,N_8496);
xor U9267 (N_9267,N_8874,N_8864);
and U9268 (N_9268,N_8920,N_8140);
or U9269 (N_9269,N_8791,N_8391);
nor U9270 (N_9270,N_8234,N_8344);
nand U9271 (N_9271,N_8775,N_8337);
xor U9272 (N_9272,N_8887,N_8037);
nand U9273 (N_9273,N_8402,N_8336);
nor U9274 (N_9274,N_8124,N_8871);
nand U9275 (N_9275,N_8005,N_8487);
nand U9276 (N_9276,N_8090,N_8618);
xnor U9277 (N_9277,N_8051,N_8721);
xor U9278 (N_9278,N_8832,N_8025);
nand U9279 (N_9279,N_8687,N_8291);
or U9280 (N_9280,N_8445,N_8643);
nand U9281 (N_9281,N_8567,N_8203);
nand U9282 (N_9282,N_8009,N_8528);
or U9283 (N_9283,N_8262,N_8021);
xnor U9284 (N_9284,N_8684,N_8719);
xor U9285 (N_9285,N_8302,N_8867);
xnor U9286 (N_9286,N_8036,N_8454);
and U9287 (N_9287,N_8635,N_8155);
and U9288 (N_9288,N_8388,N_8423);
or U9289 (N_9289,N_8156,N_8265);
xnor U9290 (N_9290,N_8230,N_8107);
nand U9291 (N_9291,N_8596,N_8836);
or U9292 (N_9292,N_8183,N_8848);
or U9293 (N_9293,N_8169,N_8866);
or U9294 (N_9294,N_8862,N_8988);
nand U9295 (N_9295,N_8695,N_8273);
or U9296 (N_9296,N_8356,N_8564);
xnor U9297 (N_9297,N_8686,N_8804);
xnor U9298 (N_9298,N_8023,N_8922);
xor U9299 (N_9299,N_8978,N_8511);
or U9300 (N_9300,N_8730,N_8340);
xnor U9301 (N_9301,N_8736,N_8440);
and U9302 (N_9302,N_8507,N_8458);
or U9303 (N_9303,N_8584,N_8079);
or U9304 (N_9304,N_8042,N_8293);
or U9305 (N_9305,N_8387,N_8304);
nor U9306 (N_9306,N_8191,N_8062);
or U9307 (N_9307,N_8301,N_8320);
or U9308 (N_9308,N_8367,N_8433);
and U9309 (N_9309,N_8679,N_8983);
and U9310 (N_9310,N_8195,N_8650);
nor U9311 (N_9311,N_8773,N_8837);
or U9312 (N_9312,N_8844,N_8768);
nand U9313 (N_9313,N_8061,N_8413);
xnor U9314 (N_9314,N_8682,N_8294);
or U9315 (N_9315,N_8396,N_8553);
nand U9316 (N_9316,N_8669,N_8460);
nand U9317 (N_9317,N_8490,N_8940);
and U9318 (N_9318,N_8209,N_8369);
xnor U9319 (N_9319,N_8597,N_8847);
xor U9320 (N_9320,N_8725,N_8353);
or U9321 (N_9321,N_8894,N_8020);
and U9322 (N_9322,N_8468,N_8271);
nand U9323 (N_9323,N_8251,N_8459);
and U9324 (N_9324,N_8976,N_8787);
xor U9325 (N_9325,N_8532,N_8308);
xnor U9326 (N_9326,N_8000,N_8779);
and U9327 (N_9327,N_8073,N_8472);
nor U9328 (N_9328,N_8379,N_8689);
and U9329 (N_9329,N_8646,N_8732);
or U9330 (N_9330,N_8168,N_8070);
nand U9331 (N_9331,N_8558,N_8398);
xnor U9332 (N_9332,N_8786,N_8656);
xor U9333 (N_9333,N_8883,N_8125);
and U9334 (N_9334,N_8906,N_8415);
nand U9335 (N_9335,N_8350,N_8479);
nor U9336 (N_9336,N_8409,N_8094);
or U9337 (N_9337,N_8505,N_8676);
nand U9338 (N_9338,N_8932,N_8708);
and U9339 (N_9339,N_8244,N_8400);
or U9340 (N_9340,N_8520,N_8927);
or U9341 (N_9341,N_8328,N_8307);
nor U9342 (N_9342,N_8860,N_8569);
nor U9343 (N_9343,N_8463,N_8362);
xnor U9344 (N_9344,N_8027,N_8637);
nor U9345 (N_9345,N_8969,N_8339);
xor U9346 (N_9346,N_8253,N_8160);
nand U9347 (N_9347,N_8006,N_8769);
and U9348 (N_9348,N_8628,N_8131);
and U9349 (N_9349,N_8106,N_8813);
xor U9350 (N_9350,N_8640,N_8523);
nor U9351 (N_9351,N_8778,N_8096);
nand U9352 (N_9352,N_8333,N_8809);
or U9353 (N_9353,N_8642,N_8054);
and U9354 (N_9354,N_8225,N_8282);
and U9355 (N_9355,N_8163,N_8432);
xnor U9356 (N_9356,N_8877,N_8625);
and U9357 (N_9357,N_8731,N_8674);
nor U9358 (N_9358,N_8419,N_8673);
nor U9359 (N_9359,N_8378,N_8289);
xor U9360 (N_9360,N_8109,N_8746);
nor U9361 (N_9361,N_8105,N_8343);
and U9362 (N_9362,N_8794,N_8178);
and U9363 (N_9363,N_8902,N_8727);
nor U9364 (N_9364,N_8377,N_8034);
nand U9365 (N_9365,N_8370,N_8657);
nor U9366 (N_9366,N_8011,N_8782);
nor U9367 (N_9367,N_8278,N_8728);
nor U9368 (N_9368,N_8812,N_8414);
nor U9369 (N_9369,N_8560,N_8510);
or U9370 (N_9370,N_8704,N_8390);
or U9371 (N_9371,N_8368,N_8057);
nor U9372 (N_9372,N_8714,N_8437);
nand U9373 (N_9373,N_8410,N_8910);
nor U9374 (N_9374,N_8175,N_8290);
xnor U9375 (N_9375,N_8017,N_8142);
nand U9376 (N_9376,N_8002,N_8828);
and U9377 (N_9377,N_8755,N_8256);
and U9378 (N_9378,N_8241,N_8380);
nand U9379 (N_9379,N_8735,N_8996);
nor U9380 (N_9380,N_8470,N_8354);
or U9381 (N_9381,N_8636,N_8164);
xnor U9382 (N_9382,N_8158,N_8557);
and U9383 (N_9383,N_8572,N_8576);
nor U9384 (N_9384,N_8207,N_8838);
nor U9385 (N_9385,N_8610,N_8008);
and U9386 (N_9386,N_8696,N_8853);
or U9387 (N_9387,N_8317,N_8992);
or U9388 (N_9388,N_8033,N_8991);
nand U9389 (N_9389,N_8121,N_8208);
xnor U9390 (N_9390,N_8601,N_8292);
nor U9391 (N_9391,N_8361,N_8788);
xor U9392 (N_9392,N_8527,N_8903);
or U9393 (N_9393,N_8602,N_8722);
nor U9394 (N_9394,N_8150,N_8371);
nor U9395 (N_9395,N_8305,N_8982);
and U9396 (N_9396,N_8918,N_8221);
nand U9397 (N_9397,N_8707,N_8884);
nor U9398 (N_9398,N_8856,N_8717);
nor U9399 (N_9399,N_8588,N_8524);
nor U9400 (N_9400,N_8076,N_8288);
nand U9401 (N_9401,N_8393,N_8647);
and U9402 (N_9402,N_8397,N_8516);
nor U9403 (N_9403,N_8546,N_8228);
nand U9404 (N_9404,N_8373,N_8612);
nand U9405 (N_9405,N_8817,N_8422);
or U9406 (N_9406,N_8015,N_8739);
and U9407 (N_9407,N_8581,N_8056);
and U9408 (N_9408,N_8952,N_8634);
nor U9409 (N_9409,N_8170,N_8645);
nor U9410 (N_9410,N_8332,N_8950);
nand U9411 (N_9411,N_8904,N_8526);
nand U9412 (N_9412,N_8229,N_8680);
nand U9413 (N_9413,N_8110,N_8120);
xnor U9414 (N_9414,N_8607,N_8958);
nand U9415 (N_9415,N_8052,N_8759);
xnor U9416 (N_9416,N_8478,N_8275);
xor U9417 (N_9417,N_8555,N_8573);
nand U9418 (N_9418,N_8711,N_8613);
xnor U9419 (N_9419,N_8845,N_8603);
nand U9420 (N_9420,N_8896,N_8655);
nand U9421 (N_9421,N_8885,N_8611);
and U9422 (N_9422,N_8401,N_8406);
nand U9423 (N_9423,N_8933,N_8627);
or U9424 (N_9424,N_8593,N_8462);
and U9425 (N_9425,N_8210,N_8043);
xor U9426 (N_9426,N_8800,N_8065);
xor U9427 (N_9427,N_8556,N_8905);
or U9428 (N_9428,N_8623,N_8223);
and U9429 (N_9429,N_8044,N_8803);
xnor U9430 (N_9430,N_8281,N_8653);
nor U9431 (N_9431,N_8534,N_8912);
or U9432 (N_9432,N_8117,N_8852);
and U9433 (N_9433,N_8999,N_8172);
xnor U9434 (N_9434,N_8954,N_8108);
nor U9435 (N_9435,N_8858,N_8024);
xor U9436 (N_9436,N_8937,N_8888);
nor U9437 (N_9437,N_8737,N_8873);
nor U9438 (N_9438,N_8901,N_8173);
xor U9439 (N_9439,N_8215,N_8863);
nand U9440 (N_9440,N_8705,N_8181);
and U9441 (N_9441,N_8539,N_8238);
nand U9442 (N_9442,N_8444,N_8450);
nor U9443 (N_9443,N_8821,N_8502);
nand U9444 (N_9444,N_8919,N_8774);
and U9445 (N_9445,N_8113,N_8091);
nand U9446 (N_9446,N_8715,N_8297);
nor U9447 (N_9447,N_8408,N_8032);
nor U9448 (N_9448,N_8661,N_8620);
or U9449 (N_9449,N_8010,N_8889);
nand U9450 (N_9450,N_8357,N_8261);
xnor U9451 (N_9451,N_8559,N_8962);
xor U9452 (N_9452,N_8604,N_8562);
and U9453 (N_9453,N_8938,N_8879);
and U9454 (N_9454,N_8754,N_8498);
xnor U9455 (N_9455,N_8616,N_8205);
nor U9456 (N_9456,N_8074,N_8849);
and U9457 (N_9457,N_8744,N_8980);
and U9458 (N_9458,N_8931,N_8372);
xnor U9459 (N_9459,N_8591,N_8102);
nand U9460 (N_9460,N_8263,N_8157);
and U9461 (N_9461,N_8018,N_8536);
or U9462 (N_9462,N_8638,N_8196);
nand U9463 (N_9463,N_8915,N_8115);
or U9464 (N_9464,N_8250,N_8143);
xnor U9465 (N_9465,N_8084,N_8934);
nand U9466 (N_9466,N_8200,N_8865);
nand U9467 (N_9467,N_8138,N_8013);
xor U9468 (N_9468,N_8622,N_8703);
or U9469 (N_9469,N_8161,N_8872);
and U9470 (N_9470,N_8961,N_8245);
and U9471 (N_9471,N_8586,N_8850);
nor U9472 (N_9472,N_8624,N_8438);
xnor U9473 (N_9473,N_8300,N_8176);
and U9474 (N_9474,N_8201,N_8348);
xnor U9475 (N_9475,N_8672,N_8099);
nor U9476 (N_9476,N_8748,N_8029);
or U9477 (N_9477,N_8619,N_8126);
xnor U9478 (N_9478,N_8233,N_8855);
xnor U9479 (N_9479,N_8299,N_8537);
nor U9480 (N_9480,N_8745,N_8480);
nand U9481 (N_9481,N_8781,N_8240);
nor U9482 (N_9482,N_8831,N_8575);
nand U9483 (N_9483,N_8810,N_8080);
nand U9484 (N_9484,N_8881,N_8805);
or U9485 (N_9485,N_8758,N_8326);
nand U9486 (N_9486,N_8434,N_8565);
nand U9487 (N_9487,N_8399,N_8485);
or U9488 (N_9488,N_8756,N_8726);
nor U9489 (N_9489,N_8834,N_8349);
xor U9490 (N_9490,N_8489,N_8058);
and U9491 (N_9491,N_8144,N_8533);
nand U9492 (N_9492,N_8405,N_8780);
nor U9493 (N_9493,N_8984,N_8957);
nand U9494 (N_9494,N_8130,N_8267);
or U9495 (N_9495,N_8796,N_8363);
and U9496 (N_9496,N_8994,N_8501);
nand U9497 (N_9497,N_8975,N_8723);
xnor U9498 (N_9498,N_8259,N_8184);
and U9499 (N_9499,N_8318,N_8484);
nand U9500 (N_9500,N_8669,N_8180);
or U9501 (N_9501,N_8566,N_8800);
or U9502 (N_9502,N_8306,N_8705);
and U9503 (N_9503,N_8827,N_8020);
xnor U9504 (N_9504,N_8863,N_8438);
xnor U9505 (N_9505,N_8777,N_8937);
and U9506 (N_9506,N_8104,N_8764);
xnor U9507 (N_9507,N_8999,N_8383);
and U9508 (N_9508,N_8532,N_8619);
xnor U9509 (N_9509,N_8475,N_8826);
nand U9510 (N_9510,N_8717,N_8608);
nand U9511 (N_9511,N_8850,N_8436);
nand U9512 (N_9512,N_8552,N_8093);
xor U9513 (N_9513,N_8976,N_8954);
or U9514 (N_9514,N_8837,N_8377);
or U9515 (N_9515,N_8693,N_8114);
nor U9516 (N_9516,N_8485,N_8331);
xnor U9517 (N_9517,N_8226,N_8859);
xor U9518 (N_9518,N_8396,N_8423);
or U9519 (N_9519,N_8210,N_8600);
nor U9520 (N_9520,N_8379,N_8307);
xnor U9521 (N_9521,N_8118,N_8331);
xnor U9522 (N_9522,N_8848,N_8535);
and U9523 (N_9523,N_8629,N_8926);
or U9524 (N_9524,N_8225,N_8244);
and U9525 (N_9525,N_8210,N_8038);
xor U9526 (N_9526,N_8129,N_8706);
xor U9527 (N_9527,N_8214,N_8321);
xnor U9528 (N_9528,N_8294,N_8589);
nand U9529 (N_9529,N_8316,N_8005);
nor U9530 (N_9530,N_8812,N_8852);
and U9531 (N_9531,N_8237,N_8883);
nand U9532 (N_9532,N_8399,N_8915);
or U9533 (N_9533,N_8724,N_8492);
and U9534 (N_9534,N_8848,N_8700);
and U9535 (N_9535,N_8122,N_8428);
nand U9536 (N_9536,N_8495,N_8870);
nor U9537 (N_9537,N_8851,N_8421);
xnor U9538 (N_9538,N_8092,N_8384);
nor U9539 (N_9539,N_8327,N_8601);
nand U9540 (N_9540,N_8838,N_8150);
and U9541 (N_9541,N_8363,N_8807);
xor U9542 (N_9542,N_8574,N_8682);
xor U9543 (N_9543,N_8598,N_8771);
or U9544 (N_9544,N_8784,N_8923);
xnor U9545 (N_9545,N_8023,N_8634);
nand U9546 (N_9546,N_8886,N_8860);
nor U9547 (N_9547,N_8617,N_8407);
xor U9548 (N_9548,N_8915,N_8301);
xor U9549 (N_9549,N_8972,N_8040);
and U9550 (N_9550,N_8354,N_8809);
or U9551 (N_9551,N_8031,N_8818);
xnor U9552 (N_9552,N_8284,N_8515);
or U9553 (N_9553,N_8746,N_8045);
xor U9554 (N_9554,N_8707,N_8816);
nand U9555 (N_9555,N_8554,N_8988);
nor U9556 (N_9556,N_8309,N_8996);
xor U9557 (N_9557,N_8488,N_8254);
nor U9558 (N_9558,N_8786,N_8836);
and U9559 (N_9559,N_8845,N_8657);
xor U9560 (N_9560,N_8352,N_8760);
nor U9561 (N_9561,N_8541,N_8023);
xor U9562 (N_9562,N_8641,N_8798);
nand U9563 (N_9563,N_8668,N_8535);
xnor U9564 (N_9564,N_8849,N_8025);
nand U9565 (N_9565,N_8052,N_8266);
or U9566 (N_9566,N_8698,N_8671);
nor U9567 (N_9567,N_8085,N_8131);
nand U9568 (N_9568,N_8975,N_8457);
or U9569 (N_9569,N_8294,N_8043);
and U9570 (N_9570,N_8063,N_8746);
xnor U9571 (N_9571,N_8048,N_8315);
and U9572 (N_9572,N_8756,N_8408);
nand U9573 (N_9573,N_8192,N_8594);
nor U9574 (N_9574,N_8709,N_8098);
xor U9575 (N_9575,N_8838,N_8009);
nand U9576 (N_9576,N_8454,N_8207);
nand U9577 (N_9577,N_8235,N_8761);
nand U9578 (N_9578,N_8350,N_8501);
or U9579 (N_9579,N_8498,N_8827);
nor U9580 (N_9580,N_8512,N_8463);
and U9581 (N_9581,N_8735,N_8068);
or U9582 (N_9582,N_8124,N_8870);
nor U9583 (N_9583,N_8366,N_8147);
nor U9584 (N_9584,N_8644,N_8450);
nor U9585 (N_9585,N_8637,N_8930);
nor U9586 (N_9586,N_8421,N_8015);
nor U9587 (N_9587,N_8923,N_8716);
nand U9588 (N_9588,N_8544,N_8007);
nand U9589 (N_9589,N_8275,N_8356);
nor U9590 (N_9590,N_8703,N_8301);
nand U9591 (N_9591,N_8862,N_8351);
or U9592 (N_9592,N_8726,N_8693);
and U9593 (N_9593,N_8918,N_8657);
nand U9594 (N_9594,N_8509,N_8698);
or U9595 (N_9595,N_8439,N_8426);
and U9596 (N_9596,N_8822,N_8061);
xor U9597 (N_9597,N_8366,N_8897);
xnor U9598 (N_9598,N_8794,N_8100);
or U9599 (N_9599,N_8177,N_8730);
nor U9600 (N_9600,N_8461,N_8120);
or U9601 (N_9601,N_8543,N_8404);
or U9602 (N_9602,N_8098,N_8126);
nor U9603 (N_9603,N_8024,N_8293);
nor U9604 (N_9604,N_8096,N_8245);
or U9605 (N_9605,N_8713,N_8033);
nor U9606 (N_9606,N_8014,N_8946);
or U9607 (N_9607,N_8005,N_8150);
nor U9608 (N_9608,N_8471,N_8690);
and U9609 (N_9609,N_8318,N_8445);
or U9610 (N_9610,N_8540,N_8366);
nor U9611 (N_9611,N_8682,N_8472);
xor U9612 (N_9612,N_8045,N_8457);
and U9613 (N_9613,N_8147,N_8331);
nor U9614 (N_9614,N_8760,N_8662);
nor U9615 (N_9615,N_8054,N_8017);
nand U9616 (N_9616,N_8147,N_8854);
and U9617 (N_9617,N_8235,N_8823);
nand U9618 (N_9618,N_8648,N_8554);
nand U9619 (N_9619,N_8008,N_8618);
and U9620 (N_9620,N_8182,N_8801);
nor U9621 (N_9621,N_8277,N_8119);
nor U9622 (N_9622,N_8304,N_8046);
nor U9623 (N_9623,N_8656,N_8073);
nand U9624 (N_9624,N_8003,N_8151);
nor U9625 (N_9625,N_8149,N_8583);
nand U9626 (N_9626,N_8996,N_8601);
and U9627 (N_9627,N_8045,N_8698);
xnor U9628 (N_9628,N_8138,N_8569);
and U9629 (N_9629,N_8689,N_8739);
and U9630 (N_9630,N_8607,N_8507);
xnor U9631 (N_9631,N_8650,N_8335);
nand U9632 (N_9632,N_8969,N_8576);
nor U9633 (N_9633,N_8752,N_8128);
xor U9634 (N_9634,N_8950,N_8707);
and U9635 (N_9635,N_8931,N_8374);
nand U9636 (N_9636,N_8140,N_8881);
nor U9637 (N_9637,N_8516,N_8731);
nand U9638 (N_9638,N_8154,N_8215);
and U9639 (N_9639,N_8199,N_8162);
nor U9640 (N_9640,N_8443,N_8805);
and U9641 (N_9641,N_8132,N_8112);
nor U9642 (N_9642,N_8480,N_8049);
nand U9643 (N_9643,N_8334,N_8368);
or U9644 (N_9644,N_8754,N_8806);
nand U9645 (N_9645,N_8014,N_8258);
nand U9646 (N_9646,N_8572,N_8570);
and U9647 (N_9647,N_8200,N_8996);
nand U9648 (N_9648,N_8886,N_8858);
nor U9649 (N_9649,N_8131,N_8033);
nor U9650 (N_9650,N_8539,N_8462);
and U9651 (N_9651,N_8497,N_8027);
xor U9652 (N_9652,N_8305,N_8995);
nand U9653 (N_9653,N_8672,N_8316);
and U9654 (N_9654,N_8671,N_8245);
xor U9655 (N_9655,N_8039,N_8364);
and U9656 (N_9656,N_8052,N_8558);
xor U9657 (N_9657,N_8243,N_8966);
nor U9658 (N_9658,N_8500,N_8448);
nand U9659 (N_9659,N_8747,N_8456);
xor U9660 (N_9660,N_8347,N_8624);
and U9661 (N_9661,N_8701,N_8938);
and U9662 (N_9662,N_8200,N_8935);
nor U9663 (N_9663,N_8054,N_8783);
xor U9664 (N_9664,N_8919,N_8970);
nor U9665 (N_9665,N_8521,N_8533);
nor U9666 (N_9666,N_8252,N_8814);
or U9667 (N_9667,N_8771,N_8891);
and U9668 (N_9668,N_8742,N_8291);
xnor U9669 (N_9669,N_8268,N_8825);
nand U9670 (N_9670,N_8481,N_8018);
nand U9671 (N_9671,N_8394,N_8354);
and U9672 (N_9672,N_8356,N_8484);
xor U9673 (N_9673,N_8917,N_8004);
nor U9674 (N_9674,N_8929,N_8055);
nand U9675 (N_9675,N_8215,N_8562);
nand U9676 (N_9676,N_8390,N_8970);
nor U9677 (N_9677,N_8277,N_8856);
and U9678 (N_9678,N_8088,N_8082);
or U9679 (N_9679,N_8225,N_8968);
and U9680 (N_9680,N_8695,N_8741);
nor U9681 (N_9681,N_8134,N_8668);
xnor U9682 (N_9682,N_8367,N_8829);
and U9683 (N_9683,N_8464,N_8604);
nor U9684 (N_9684,N_8317,N_8327);
nor U9685 (N_9685,N_8354,N_8841);
nand U9686 (N_9686,N_8551,N_8520);
xor U9687 (N_9687,N_8071,N_8687);
nor U9688 (N_9688,N_8244,N_8983);
nand U9689 (N_9689,N_8869,N_8821);
or U9690 (N_9690,N_8617,N_8187);
nand U9691 (N_9691,N_8789,N_8354);
nand U9692 (N_9692,N_8639,N_8107);
nand U9693 (N_9693,N_8821,N_8324);
nor U9694 (N_9694,N_8271,N_8446);
nand U9695 (N_9695,N_8356,N_8786);
xor U9696 (N_9696,N_8243,N_8920);
nand U9697 (N_9697,N_8037,N_8884);
nand U9698 (N_9698,N_8216,N_8266);
xor U9699 (N_9699,N_8519,N_8157);
or U9700 (N_9700,N_8470,N_8572);
nand U9701 (N_9701,N_8575,N_8926);
nand U9702 (N_9702,N_8999,N_8848);
nor U9703 (N_9703,N_8024,N_8835);
or U9704 (N_9704,N_8028,N_8210);
nor U9705 (N_9705,N_8215,N_8049);
and U9706 (N_9706,N_8667,N_8442);
or U9707 (N_9707,N_8704,N_8168);
nand U9708 (N_9708,N_8319,N_8927);
xor U9709 (N_9709,N_8968,N_8610);
nand U9710 (N_9710,N_8472,N_8730);
nand U9711 (N_9711,N_8965,N_8685);
nor U9712 (N_9712,N_8782,N_8775);
nor U9713 (N_9713,N_8412,N_8279);
nand U9714 (N_9714,N_8506,N_8205);
xor U9715 (N_9715,N_8605,N_8419);
nand U9716 (N_9716,N_8474,N_8935);
and U9717 (N_9717,N_8335,N_8140);
and U9718 (N_9718,N_8319,N_8677);
and U9719 (N_9719,N_8407,N_8658);
nor U9720 (N_9720,N_8108,N_8544);
nand U9721 (N_9721,N_8444,N_8904);
nor U9722 (N_9722,N_8782,N_8913);
and U9723 (N_9723,N_8786,N_8617);
xnor U9724 (N_9724,N_8515,N_8005);
and U9725 (N_9725,N_8026,N_8106);
nor U9726 (N_9726,N_8781,N_8270);
xor U9727 (N_9727,N_8377,N_8490);
xnor U9728 (N_9728,N_8211,N_8498);
and U9729 (N_9729,N_8967,N_8902);
and U9730 (N_9730,N_8090,N_8682);
or U9731 (N_9731,N_8324,N_8851);
nor U9732 (N_9732,N_8847,N_8863);
xnor U9733 (N_9733,N_8915,N_8913);
and U9734 (N_9734,N_8080,N_8765);
and U9735 (N_9735,N_8649,N_8897);
nand U9736 (N_9736,N_8540,N_8008);
nand U9737 (N_9737,N_8610,N_8884);
and U9738 (N_9738,N_8746,N_8187);
or U9739 (N_9739,N_8232,N_8813);
nor U9740 (N_9740,N_8399,N_8252);
nand U9741 (N_9741,N_8824,N_8514);
nand U9742 (N_9742,N_8972,N_8538);
and U9743 (N_9743,N_8573,N_8912);
nand U9744 (N_9744,N_8393,N_8859);
nor U9745 (N_9745,N_8273,N_8206);
and U9746 (N_9746,N_8574,N_8538);
nor U9747 (N_9747,N_8507,N_8814);
nand U9748 (N_9748,N_8058,N_8790);
xnor U9749 (N_9749,N_8109,N_8802);
xor U9750 (N_9750,N_8699,N_8085);
nor U9751 (N_9751,N_8568,N_8394);
and U9752 (N_9752,N_8625,N_8701);
nand U9753 (N_9753,N_8572,N_8483);
or U9754 (N_9754,N_8599,N_8075);
nand U9755 (N_9755,N_8742,N_8239);
xnor U9756 (N_9756,N_8820,N_8284);
nand U9757 (N_9757,N_8519,N_8474);
and U9758 (N_9758,N_8710,N_8630);
or U9759 (N_9759,N_8805,N_8039);
xor U9760 (N_9760,N_8399,N_8686);
nor U9761 (N_9761,N_8022,N_8597);
nand U9762 (N_9762,N_8980,N_8404);
and U9763 (N_9763,N_8769,N_8052);
and U9764 (N_9764,N_8348,N_8160);
nand U9765 (N_9765,N_8624,N_8561);
or U9766 (N_9766,N_8482,N_8388);
or U9767 (N_9767,N_8136,N_8341);
xnor U9768 (N_9768,N_8521,N_8202);
nor U9769 (N_9769,N_8235,N_8833);
nor U9770 (N_9770,N_8917,N_8641);
nor U9771 (N_9771,N_8221,N_8712);
and U9772 (N_9772,N_8179,N_8171);
nand U9773 (N_9773,N_8505,N_8126);
or U9774 (N_9774,N_8732,N_8974);
nor U9775 (N_9775,N_8806,N_8236);
xnor U9776 (N_9776,N_8345,N_8939);
nor U9777 (N_9777,N_8146,N_8906);
and U9778 (N_9778,N_8134,N_8713);
and U9779 (N_9779,N_8611,N_8425);
nor U9780 (N_9780,N_8730,N_8376);
or U9781 (N_9781,N_8207,N_8417);
nor U9782 (N_9782,N_8739,N_8145);
nor U9783 (N_9783,N_8628,N_8359);
nor U9784 (N_9784,N_8947,N_8087);
or U9785 (N_9785,N_8490,N_8362);
xor U9786 (N_9786,N_8344,N_8586);
xor U9787 (N_9787,N_8370,N_8761);
nand U9788 (N_9788,N_8732,N_8016);
nand U9789 (N_9789,N_8230,N_8982);
and U9790 (N_9790,N_8123,N_8211);
or U9791 (N_9791,N_8368,N_8777);
xor U9792 (N_9792,N_8883,N_8502);
or U9793 (N_9793,N_8286,N_8708);
nor U9794 (N_9794,N_8956,N_8844);
nand U9795 (N_9795,N_8437,N_8258);
xnor U9796 (N_9796,N_8579,N_8653);
nor U9797 (N_9797,N_8797,N_8151);
and U9798 (N_9798,N_8629,N_8593);
nand U9799 (N_9799,N_8735,N_8259);
nor U9800 (N_9800,N_8552,N_8424);
xor U9801 (N_9801,N_8283,N_8204);
nor U9802 (N_9802,N_8302,N_8185);
or U9803 (N_9803,N_8065,N_8122);
and U9804 (N_9804,N_8137,N_8305);
or U9805 (N_9805,N_8801,N_8580);
and U9806 (N_9806,N_8049,N_8614);
xor U9807 (N_9807,N_8650,N_8352);
xor U9808 (N_9808,N_8347,N_8757);
or U9809 (N_9809,N_8649,N_8856);
or U9810 (N_9810,N_8491,N_8717);
xnor U9811 (N_9811,N_8152,N_8556);
nor U9812 (N_9812,N_8305,N_8610);
xnor U9813 (N_9813,N_8613,N_8976);
or U9814 (N_9814,N_8624,N_8694);
nand U9815 (N_9815,N_8186,N_8467);
nand U9816 (N_9816,N_8615,N_8321);
nor U9817 (N_9817,N_8971,N_8460);
and U9818 (N_9818,N_8245,N_8639);
xnor U9819 (N_9819,N_8889,N_8703);
and U9820 (N_9820,N_8389,N_8225);
nand U9821 (N_9821,N_8563,N_8755);
or U9822 (N_9822,N_8811,N_8056);
nor U9823 (N_9823,N_8053,N_8939);
and U9824 (N_9824,N_8526,N_8714);
nor U9825 (N_9825,N_8416,N_8268);
or U9826 (N_9826,N_8002,N_8700);
xnor U9827 (N_9827,N_8707,N_8672);
xnor U9828 (N_9828,N_8839,N_8053);
nand U9829 (N_9829,N_8081,N_8514);
nor U9830 (N_9830,N_8423,N_8870);
xnor U9831 (N_9831,N_8376,N_8186);
and U9832 (N_9832,N_8126,N_8802);
nand U9833 (N_9833,N_8131,N_8228);
nand U9834 (N_9834,N_8417,N_8458);
xor U9835 (N_9835,N_8928,N_8954);
nor U9836 (N_9836,N_8756,N_8583);
nor U9837 (N_9837,N_8604,N_8500);
xnor U9838 (N_9838,N_8386,N_8247);
nor U9839 (N_9839,N_8819,N_8914);
xor U9840 (N_9840,N_8453,N_8191);
nor U9841 (N_9841,N_8617,N_8807);
and U9842 (N_9842,N_8841,N_8129);
nor U9843 (N_9843,N_8462,N_8589);
nor U9844 (N_9844,N_8449,N_8752);
xnor U9845 (N_9845,N_8193,N_8655);
nor U9846 (N_9846,N_8135,N_8816);
nor U9847 (N_9847,N_8088,N_8503);
xnor U9848 (N_9848,N_8371,N_8982);
nand U9849 (N_9849,N_8386,N_8448);
nor U9850 (N_9850,N_8810,N_8826);
and U9851 (N_9851,N_8573,N_8584);
and U9852 (N_9852,N_8076,N_8539);
nand U9853 (N_9853,N_8063,N_8071);
nor U9854 (N_9854,N_8393,N_8355);
nand U9855 (N_9855,N_8229,N_8054);
nand U9856 (N_9856,N_8658,N_8971);
or U9857 (N_9857,N_8908,N_8833);
and U9858 (N_9858,N_8141,N_8871);
xnor U9859 (N_9859,N_8404,N_8281);
or U9860 (N_9860,N_8570,N_8108);
xnor U9861 (N_9861,N_8288,N_8567);
nor U9862 (N_9862,N_8690,N_8717);
or U9863 (N_9863,N_8458,N_8155);
xnor U9864 (N_9864,N_8560,N_8620);
nor U9865 (N_9865,N_8924,N_8015);
or U9866 (N_9866,N_8699,N_8662);
xnor U9867 (N_9867,N_8741,N_8318);
and U9868 (N_9868,N_8510,N_8972);
xnor U9869 (N_9869,N_8403,N_8540);
or U9870 (N_9870,N_8880,N_8016);
or U9871 (N_9871,N_8705,N_8803);
or U9872 (N_9872,N_8899,N_8781);
or U9873 (N_9873,N_8598,N_8793);
nor U9874 (N_9874,N_8396,N_8327);
xor U9875 (N_9875,N_8969,N_8807);
and U9876 (N_9876,N_8060,N_8408);
and U9877 (N_9877,N_8951,N_8137);
or U9878 (N_9878,N_8578,N_8495);
and U9879 (N_9879,N_8708,N_8941);
and U9880 (N_9880,N_8835,N_8349);
nor U9881 (N_9881,N_8186,N_8744);
nor U9882 (N_9882,N_8787,N_8108);
or U9883 (N_9883,N_8195,N_8558);
xnor U9884 (N_9884,N_8292,N_8609);
and U9885 (N_9885,N_8664,N_8812);
xnor U9886 (N_9886,N_8625,N_8105);
or U9887 (N_9887,N_8001,N_8659);
and U9888 (N_9888,N_8490,N_8440);
nor U9889 (N_9889,N_8696,N_8139);
nor U9890 (N_9890,N_8600,N_8163);
or U9891 (N_9891,N_8265,N_8660);
or U9892 (N_9892,N_8757,N_8950);
xnor U9893 (N_9893,N_8017,N_8710);
nor U9894 (N_9894,N_8029,N_8475);
nand U9895 (N_9895,N_8428,N_8464);
xor U9896 (N_9896,N_8762,N_8328);
xor U9897 (N_9897,N_8390,N_8421);
nor U9898 (N_9898,N_8176,N_8693);
xnor U9899 (N_9899,N_8659,N_8514);
nor U9900 (N_9900,N_8911,N_8356);
nor U9901 (N_9901,N_8073,N_8735);
or U9902 (N_9902,N_8687,N_8016);
nand U9903 (N_9903,N_8750,N_8401);
xor U9904 (N_9904,N_8821,N_8522);
nor U9905 (N_9905,N_8382,N_8012);
nand U9906 (N_9906,N_8467,N_8436);
xnor U9907 (N_9907,N_8035,N_8853);
nand U9908 (N_9908,N_8308,N_8264);
xnor U9909 (N_9909,N_8610,N_8791);
nand U9910 (N_9910,N_8039,N_8461);
nor U9911 (N_9911,N_8014,N_8289);
xor U9912 (N_9912,N_8795,N_8706);
nor U9913 (N_9913,N_8429,N_8155);
xor U9914 (N_9914,N_8524,N_8122);
nand U9915 (N_9915,N_8102,N_8396);
and U9916 (N_9916,N_8326,N_8820);
nand U9917 (N_9917,N_8809,N_8106);
nor U9918 (N_9918,N_8660,N_8330);
nand U9919 (N_9919,N_8668,N_8946);
or U9920 (N_9920,N_8358,N_8436);
nand U9921 (N_9921,N_8637,N_8061);
nor U9922 (N_9922,N_8122,N_8507);
or U9923 (N_9923,N_8727,N_8285);
or U9924 (N_9924,N_8143,N_8961);
nor U9925 (N_9925,N_8670,N_8805);
nand U9926 (N_9926,N_8482,N_8937);
nand U9927 (N_9927,N_8595,N_8020);
xor U9928 (N_9928,N_8640,N_8317);
nor U9929 (N_9929,N_8214,N_8728);
or U9930 (N_9930,N_8328,N_8516);
nand U9931 (N_9931,N_8349,N_8182);
nand U9932 (N_9932,N_8665,N_8367);
and U9933 (N_9933,N_8796,N_8499);
and U9934 (N_9934,N_8033,N_8104);
nand U9935 (N_9935,N_8902,N_8771);
nor U9936 (N_9936,N_8752,N_8884);
and U9937 (N_9937,N_8386,N_8259);
nor U9938 (N_9938,N_8553,N_8854);
or U9939 (N_9939,N_8583,N_8285);
nor U9940 (N_9940,N_8698,N_8082);
xnor U9941 (N_9941,N_8012,N_8223);
nor U9942 (N_9942,N_8022,N_8116);
nand U9943 (N_9943,N_8438,N_8415);
or U9944 (N_9944,N_8261,N_8386);
and U9945 (N_9945,N_8598,N_8608);
xor U9946 (N_9946,N_8326,N_8912);
and U9947 (N_9947,N_8409,N_8056);
nor U9948 (N_9948,N_8667,N_8429);
and U9949 (N_9949,N_8430,N_8833);
nor U9950 (N_9950,N_8396,N_8550);
or U9951 (N_9951,N_8238,N_8373);
xor U9952 (N_9952,N_8840,N_8417);
xnor U9953 (N_9953,N_8281,N_8609);
and U9954 (N_9954,N_8343,N_8562);
nor U9955 (N_9955,N_8071,N_8089);
and U9956 (N_9956,N_8857,N_8057);
and U9957 (N_9957,N_8406,N_8170);
xnor U9958 (N_9958,N_8647,N_8155);
nand U9959 (N_9959,N_8546,N_8821);
and U9960 (N_9960,N_8001,N_8092);
or U9961 (N_9961,N_8457,N_8925);
and U9962 (N_9962,N_8290,N_8262);
nand U9963 (N_9963,N_8681,N_8457);
xnor U9964 (N_9964,N_8294,N_8144);
nor U9965 (N_9965,N_8995,N_8979);
nand U9966 (N_9966,N_8662,N_8495);
nand U9967 (N_9967,N_8077,N_8423);
or U9968 (N_9968,N_8360,N_8732);
and U9969 (N_9969,N_8632,N_8177);
and U9970 (N_9970,N_8849,N_8402);
and U9971 (N_9971,N_8151,N_8375);
or U9972 (N_9972,N_8190,N_8474);
xnor U9973 (N_9973,N_8040,N_8033);
nand U9974 (N_9974,N_8510,N_8742);
nor U9975 (N_9975,N_8136,N_8840);
xor U9976 (N_9976,N_8367,N_8386);
nor U9977 (N_9977,N_8324,N_8008);
and U9978 (N_9978,N_8046,N_8047);
nor U9979 (N_9979,N_8989,N_8643);
xor U9980 (N_9980,N_8199,N_8725);
or U9981 (N_9981,N_8792,N_8669);
and U9982 (N_9982,N_8850,N_8404);
nand U9983 (N_9983,N_8295,N_8938);
nor U9984 (N_9984,N_8903,N_8343);
and U9985 (N_9985,N_8732,N_8716);
xnor U9986 (N_9986,N_8224,N_8478);
nor U9987 (N_9987,N_8195,N_8875);
nand U9988 (N_9988,N_8161,N_8757);
nand U9989 (N_9989,N_8098,N_8154);
nand U9990 (N_9990,N_8795,N_8422);
or U9991 (N_9991,N_8924,N_8268);
or U9992 (N_9992,N_8018,N_8977);
xor U9993 (N_9993,N_8563,N_8430);
or U9994 (N_9994,N_8380,N_8438);
nand U9995 (N_9995,N_8295,N_8370);
or U9996 (N_9996,N_8832,N_8688);
nor U9997 (N_9997,N_8813,N_8128);
nor U9998 (N_9998,N_8957,N_8685);
and U9999 (N_9999,N_8071,N_8803);
or U10000 (N_10000,N_9603,N_9775);
xor U10001 (N_10001,N_9834,N_9607);
nand U10002 (N_10002,N_9968,N_9242);
or U10003 (N_10003,N_9040,N_9793);
xor U10004 (N_10004,N_9896,N_9489);
xor U10005 (N_10005,N_9759,N_9004);
xor U10006 (N_10006,N_9099,N_9610);
xnor U10007 (N_10007,N_9111,N_9996);
nor U10008 (N_10008,N_9296,N_9168);
and U10009 (N_10009,N_9398,N_9861);
or U10010 (N_10010,N_9782,N_9048);
xor U10011 (N_10011,N_9375,N_9229);
nor U10012 (N_10012,N_9467,N_9729);
and U10013 (N_10013,N_9654,N_9276);
nor U10014 (N_10014,N_9904,N_9611);
or U10015 (N_10015,N_9660,N_9370);
nand U10016 (N_10016,N_9414,N_9681);
and U10017 (N_10017,N_9621,N_9496);
nand U10018 (N_10018,N_9018,N_9689);
and U10019 (N_10019,N_9288,N_9854);
xnor U10020 (N_10020,N_9286,N_9870);
and U10021 (N_10021,N_9228,N_9580);
nor U10022 (N_10022,N_9490,N_9275);
xnor U10023 (N_10023,N_9056,N_9540);
xnor U10024 (N_10024,N_9137,N_9383);
nor U10025 (N_10025,N_9434,N_9876);
nor U10026 (N_10026,N_9149,N_9172);
or U10027 (N_10027,N_9362,N_9957);
xor U10028 (N_10028,N_9795,N_9486);
nor U10029 (N_10029,N_9049,N_9731);
or U10030 (N_10030,N_9444,N_9244);
nand U10031 (N_10031,N_9236,N_9727);
and U10032 (N_10032,N_9059,N_9461);
nand U10033 (N_10033,N_9525,N_9814);
and U10034 (N_10034,N_9800,N_9218);
and U10035 (N_10035,N_9166,N_9928);
nand U10036 (N_10036,N_9431,N_9708);
nand U10037 (N_10037,N_9354,N_9881);
nor U10038 (N_10038,N_9678,N_9754);
nor U10039 (N_10039,N_9969,N_9455);
xor U10040 (N_10040,N_9245,N_9669);
nor U10041 (N_10041,N_9404,N_9034);
nor U10042 (N_10042,N_9052,N_9620);
xnor U10043 (N_10043,N_9790,N_9131);
nand U10044 (N_10044,N_9884,N_9483);
nor U10045 (N_10045,N_9578,N_9779);
xor U10046 (N_10046,N_9157,N_9728);
nor U10047 (N_10047,N_9565,N_9348);
and U10048 (N_10048,N_9984,N_9911);
and U10049 (N_10049,N_9737,N_9602);
or U10050 (N_10050,N_9736,N_9652);
nand U10051 (N_10051,N_9748,N_9614);
nand U10052 (N_10052,N_9688,N_9224);
xnor U10053 (N_10053,N_9591,N_9261);
nand U10054 (N_10054,N_9115,N_9093);
nor U10055 (N_10055,N_9178,N_9910);
and U10056 (N_10056,N_9871,N_9555);
nor U10057 (N_10057,N_9344,N_9371);
or U10058 (N_10058,N_9575,N_9917);
or U10059 (N_10059,N_9703,N_9158);
xor U10060 (N_10060,N_9686,N_9505);
xnor U10061 (N_10061,N_9480,N_9560);
xor U10062 (N_10062,N_9629,N_9290);
nor U10063 (N_10063,N_9246,N_9514);
nor U10064 (N_10064,N_9888,N_9347);
or U10065 (N_10065,N_9476,N_9351);
xor U10066 (N_10066,N_9187,N_9237);
and U10067 (N_10067,N_9940,N_9202);
xnor U10068 (N_10068,N_9912,N_9331);
xor U10069 (N_10069,N_9209,N_9098);
xor U10070 (N_10070,N_9430,N_9134);
and U10071 (N_10071,N_9060,N_9036);
xor U10072 (N_10072,N_9140,N_9777);
and U10073 (N_10073,N_9475,N_9577);
nor U10074 (N_10074,N_9363,N_9494);
or U10075 (N_10075,N_9102,N_9074);
and U10076 (N_10076,N_9420,N_9104);
nor U10077 (N_10077,N_9338,N_9891);
or U10078 (N_10078,N_9898,N_9125);
and U10079 (N_10079,N_9081,N_9346);
nand U10080 (N_10080,N_9023,N_9510);
xnor U10081 (N_10081,N_9674,N_9446);
xor U10082 (N_10082,N_9468,N_9985);
and U10083 (N_10083,N_9887,N_9076);
nor U10084 (N_10084,N_9316,N_9506);
xor U10085 (N_10085,N_9920,N_9132);
and U10086 (N_10086,N_9189,N_9964);
and U10087 (N_10087,N_9762,N_9921);
xor U10088 (N_10088,N_9767,N_9193);
or U10089 (N_10089,N_9963,N_9012);
and U10090 (N_10090,N_9041,N_9367);
nand U10091 (N_10091,N_9027,N_9190);
xnor U10092 (N_10092,N_9211,N_9712);
or U10093 (N_10093,N_9447,N_9450);
or U10094 (N_10094,N_9343,N_9293);
or U10095 (N_10095,N_9504,N_9355);
xor U10096 (N_10096,N_9305,N_9219);
nand U10097 (N_10097,N_9235,N_9820);
and U10098 (N_10098,N_9144,N_9875);
nor U10099 (N_10099,N_9718,N_9271);
nor U10100 (N_10100,N_9417,N_9742);
xor U10101 (N_10101,N_9961,N_9241);
nor U10102 (N_10102,N_9029,N_9666);
nand U10103 (N_10103,N_9693,N_9259);
nor U10104 (N_10104,N_9265,N_9557);
xor U10105 (N_10105,N_9277,N_9208);
xor U10106 (N_10106,N_9735,N_9186);
xor U10107 (N_10107,N_9773,N_9217);
nor U10108 (N_10108,N_9720,N_9069);
or U10109 (N_10109,N_9010,N_9092);
nand U10110 (N_10110,N_9806,N_9582);
or U10111 (N_10111,N_9598,N_9413);
nand U10112 (N_10112,N_9032,N_9634);
nand U10113 (N_10113,N_9571,N_9758);
nor U10114 (N_10114,N_9992,N_9942);
or U10115 (N_10115,N_9195,N_9799);
and U10116 (N_10116,N_9415,N_9472);
xnor U10117 (N_10117,N_9295,N_9661);
nor U10118 (N_10118,N_9792,N_9433);
nor U10119 (N_10119,N_9079,N_9987);
xnor U10120 (N_10120,N_9897,N_9151);
nand U10121 (N_10121,N_9273,N_9118);
xor U10122 (N_10122,N_9618,N_9922);
and U10123 (N_10123,N_9141,N_9308);
nor U10124 (N_10124,N_9667,N_9533);
and U10125 (N_10125,N_9200,N_9460);
or U10126 (N_10126,N_9812,N_9757);
xnor U10127 (N_10127,N_9334,N_9570);
xor U10128 (N_10128,N_9947,N_9873);
nand U10129 (N_10129,N_9329,N_9901);
nor U10130 (N_10130,N_9648,N_9222);
nor U10131 (N_10131,N_9326,N_9791);
or U10132 (N_10132,N_9169,N_9774);
xnor U10133 (N_10133,N_9683,N_9117);
nor U10134 (N_10134,N_9124,N_9590);
nor U10135 (N_10135,N_9154,N_9606);
nor U10136 (N_10136,N_9088,N_9303);
nand U10137 (N_10137,N_9650,N_9000);
xor U10138 (N_10138,N_9630,N_9473);
nand U10139 (N_10139,N_9361,N_9702);
xnor U10140 (N_10140,N_9670,N_9436);
nand U10141 (N_10141,N_9492,N_9238);
nor U10142 (N_10142,N_9958,N_9859);
nand U10143 (N_10143,N_9142,N_9597);
and U10144 (N_10144,N_9082,N_9682);
nand U10145 (N_10145,N_9274,N_9828);
and U10146 (N_10146,N_9804,N_9519);
nand U10147 (N_10147,N_9596,N_9339);
nand U10148 (N_10148,N_9527,N_9579);
nand U10149 (N_10149,N_9651,N_9553);
xor U10150 (N_10150,N_9488,N_9395);
nand U10151 (N_10151,N_9379,N_9127);
nand U10152 (N_10152,N_9412,N_9763);
nor U10153 (N_10153,N_9613,N_9517);
or U10154 (N_10154,N_9826,N_9130);
nand U10155 (N_10155,N_9173,N_9322);
or U10156 (N_10156,N_9498,N_9907);
nor U10157 (N_10157,N_9509,N_9085);
and U10158 (N_10158,N_9396,N_9991);
nor U10159 (N_10159,N_9309,N_9419);
and U10160 (N_10160,N_9556,N_9880);
xnor U10161 (N_10161,N_9179,N_9452);
xor U10162 (N_10162,N_9177,N_9722);
or U10163 (N_10163,N_9824,N_9437);
nand U10164 (N_10164,N_9341,N_9995);
xor U10165 (N_10165,N_9233,N_9442);
nand U10166 (N_10166,N_9655,N_9636);
and U10167 (N_10167,N_9146,N_9045);
or U10168 (N_10168,N_9234,N_9199);
and U10169 (N_10169,N_9979,N_9864);
and U10170 (N_10170,N_9905,N_9285);
nand U10171 (N_10171,N_9687,N_9933);
xor U10172 (N_10172,N_9312,N_9369);
nor U10173 (N_10173,N_9663,N_9647);
and U10174 (N_10174,N_9521,N_9279);
xnor U10175 (N_10175,N_9284,N_9659);
or U10176 (N_10176,N_9213,N_9147);
xnor U10177 (N_10177,N_9156,N_9609);
or U10178 (N_10178,N_9599,N_9402);
nor U10179 (N_10179,N_9340,N_9656);
xor U10180 (N_10180,N_9955,N_9943);
xnor U10181 (N_10181,N_9707,N_9292);
and U10182 (N_10182,N_9903,N_9109);
xnor U10183 (N_10183,N_9332,N_9640);
or U10184 (N_10184,N_9025,N_9256);
and U10185 (N_10185,N_9129,N_9716);
and U10186 (N_10186,N_9809,N_9587);
or U10187 (N_10187,N_9230,N_9106);
or U10188 (N_10188,N_9822,N_9267);
nor U10189 (N_10189,N_9949,N_9105);
and U10190 (N_10190,N_9511,N_9451);
or U10191 (N_10191,N_9251,N_9051);
xnor U10192 (N_10192,N_9207,N_9892);
xor U10193 (N_10193,N_9994,N_9119);
and U10194 (N_10194,N_9091,N_9310);
nor U10195 (N_10195,N_9584,N_9583);
or U10196 (N_10196,N_9948,N_9588);
or U10197 (N_10197,N_9798,N_9950);
and U10198 (N_10198,N_9448,N_9665);
and U10199 (N_10199,N_9679,N_9794);
and U10200 (N_10200,N_9306,N_9358);
nor U10201 (N_10201,N_9047,N_9038);
or U10202 (N_10202,N_9021,N_9198);
nor U10203 (N_10203,N_9740,N_9479);
nor U10204 (N_10204,N_9529,N_9110);
or U10205 (N_10205,N_9877,N_9772);
xnor U10206 (N_10206,N_9150,N_9879);
xnor U10207 (N_10207,N_9171,N_9977);
nor U10208 (N_10208,N_9923,N_9815);
or U10209 (N_10209,N_9366,N_9847);
and U10210 (N_10210,N_9971,N_9014);
xnor U10211 (N_10211,N_9300,N_9990);
nor U10212 (N_10212,N_9321,N_9786);
nand U10213 (N_10213,N_9534,N_9778);
xnor U10214 (N_10214,N_9843,N_9205);
nand U10215 (N_10215,N_9184,N_9170);
and U10216 (N_10216,N_9657,N_9484);
or U10217 (N_10217,N_9280,N_9204);
nand U10218 (N_10218,N_9487,N_9938);
nand U10219 (N_10219,N_9925,N_9960);
or U10220 (N_10220,N_9212,N_9719);
and U10221 (N_10221,N_9016,N_9002);
nor U10222 (N_10222,N_9972,N_9314);
or U10223 (N_10223,N_9311,N_9072);
xnor U10224 (N_10224,N_9668,N_9975);
and U10225 (N_10225,N_9410,N_9680);
and U10226 (N_10226,N_9185,N_9123);
and U10227 (N_10227,N_9988,N_9558);
or U10228 (N_10228,N_9546,N_9068);
and U10229 (N_10229,N_9357,N_9725);
xor U10230 (N_10230,N_9094,N_9073);
or U10231 (N_10231,N_9941,N_9216);
nand U10232 (N_10232,N_9443,N_9999);
and U10233 (N_10233,N_9266,N_9856);
xnor U10234 (N_10234,N_9268,N_9559);
nand U10235 (N_10235,N_9421,N_9684);
nand U10236 (N_10236,N_9262,N_9906);
nor U10237 (N_10237,N_9015,N_9771);
nor U10238 (N_10238,N_9260,N_9739);
nor U10239 (N_10239,N_9075,N_9539);
xnor U10240 (N_10240,N_9165,N_9493);
xor U10241 (N_10241,N_9258,N_9839);
and U10242 (N_10242,N_9645,N_9466);
nor U10243 (N_10243,N_9715,N_9254);
xnor U10244 (N_10244,N_9352,N_9003);
xnor U10245 (N_10245,N_9249,N_9116);
nand U10246 (N_10246,N_9787,N_9019);
and U10247 (N_10247,N_9699,N_9853);
nor U10248 (N_10248,N_9252,N_9840);
or U10249 (N_10249,N_9176,N_9902);
nor U10250 (N_10250,N_9465,N_9627);
nand U10251 (N_10251,N_9829,N_9152);
and U10252 (N_10252,N_9263,N_9574);
nor U10253 (N_10253,N_9225,N_9495);
and U10254 (N_10254,N_9071,N_9913);
nand U10255 (N_10255,N_9457,N_9206);
nor U10256 (N_10256,N_9743,N_9463);
nand U10257 (N_10257,N_9440,N_9783);
nor U10258 (N_10258,N_9653,N_9866);
or U10259 (N_10259,N_9697,N_9622);
xnor U10260 (N_10260,N_9818,N_9924);
and U10261 (N_10261,N_9282,N_9247);
and U10262 (N_10262,N_9210,N_9232);
xnor U10263 (N_10263,N_9320,N_9153);
and U10264 (N_10264,N_9628,N_9882);
and U10265 (N_10265,N_9594,N_9862);
xnor U10266 (N_10266,N_9714,N_9624);
xnor U10267 (N_10267,N_9428,N_9845);
and U10268 (N_10268,N_9087,N_9857);
or U10269 (N_10269,N_9914,N_9313);
nor U10270 (N_10270,N_9530,N_9175);
or U10271 (N_10271,N_9547,N_9641);
xnor U10272 (N_10272,N_9054,N_9044);
and U10273 (N_10273,N_9089,N_9253);
or U10274 (N_10274,N_9980,N_9376);
and U10275 (N_10275,N_9459,N_9808);
or U10276 (N_10276,N_9062,N_9302);
nand U10277 (N_10277,N_9625,N_9781);
or U10278 (N_10278,N_9518,N_9841);
nor U10279 (N_10279,N_9753,N_9600);
nor U10280 (N_10280,N_9512,N_9751);
and U10281 (N_10281,N_9393,N_9899);
nand U10282 (N_10282,N_9848,N_9389);
nand U10283 (N_10283,N_9478,N_9356);
xor U10284 (N_10284,N_9738,N_9989);
or U10285 (N_10285,N_9011,N_9120);
nor U10286 (N_10286,N_9863,N_9272);
or U10287 (N_10287,N_9741,N_9664);
nand U10288 (N_10288,N_9700,N_9020);
nor U10289 (N_10289,N_9935,N_9919);
nor U10290 (N_10290,N_9128,N_9567);
or U10291 (N_10291,N_9974,N_9802);
xor U10292 (N_10292,N_9005,N_9315);
or U10293 (N_10293,N_9294,N_9709);
nand U10294 (N_10294,N_9524,N_9592);
nand U10295 (N_10295,N_9959,N_9978);
or U10296 (N_10296,N_9501,N_9766);
xor U10297 (N_10297,N_9677,N_9477);
xnor U10298 (N_10298,N_9243,N_9837);
xnor U10299 (N_10299,N_9915,N_9255);
xnor U10300 (N_10300,N_9726,N_9585);
nand U10301 (N_10301,N_9456,N_9350);
nand U10302 (N_10302,N_9507,N_9359);
nor U10303 (N_10303,N_9765,N_9564);
nand U10304 (N_10304,N_9746,N_9692);
and U10305 (N_10305,N_9576,N_9058);
nand U10306 (N_10306,N_9033,N_9986);
xnor U10307 (N_10307,N_9240,N_9006);
or U10308 (N_10308,N_9523,N_9724);
nand U10309 (N_10309,N_9471,N_9377);
nor U10310 (N_10310,N_9250,N_9046);
xnor U10311 (N_10311,N_9572,N_9954);
nor U10312 (N_10312,N_9403,N_9333);
xnor U10313 (N_10313,N_9445,N_9874);
xor U10314 (N_10314,N_9387,N_9803);
nand U10315 (N_10315,N_9043,N_9095);
xnor U10316 (N_10316,N_9944,N_9926);
nor U10317 (N_10317,N_9701,N_9878);
and U10318 (N_10318,N_9353,N_9257);
nand U10319 (N_10319,N_9939,N_9161);
nor U10320 (N_10320,N_9723,N_9865);
or U10321 (N_10321,N_9345,N_9976);
xor U10322 (N_10322,N_9932,N_9136);
or U10323 (N_10323,N_9662,N_9744);
nand U10324 (N_10324,N_9439,N_9890);
nand U10325 (N_10325,N_9408,N_9860);
xor U10326 (N_10326,N_9965,N_9164);
nand U10327 (N_10327,N_9077,N_9017);
nor U10328 (N_10328,N_9418,N_9400);
xnor U10329 (N_10329,N_9672,N_9589);
nand U10330 (N_10330,N_9770,N_9318);
nand U10331 (N_10331,N_9894,N_9122);
xnor U10332 (N_10332,N_9562,N_9581);
nand U10333 (N_10333,N_9868,N_9180);
nand U10334 (N_10334,N_9462,N_9126);
nor U10335 (N_10335,N_9385,N_9842);
or U10336 (N_10336,N_9850,N_9223);
xnor U10337 (N_10337,N_9066,N_9671);
xor U10338 (N_10338,N_9830,N_9458);
nand U10339 (N_10339,N_9515,N_9291);
or U10340 (N_10340,N_9438,N_9063);
xor U10341 (N_10341,N_9215,N_9192);
xor U10342 (N_10342,N_9544,N_9227);
nor U10343 (N_10343,N_9858,N_9929);
nor U10344 (N_10344,N_9554,N_9336);
and U10345 (N_10345,N_9807,N_9100);
nand U10346 (N_10346,N_9391,N_9042);
or U10347 (N_10347,N_9900,N_9747);
and U10348 (N_10348,N_9427,N_9080);
nand U10349 (N_10349,N_9704,N_9392);
xor U10350 (N_10350,N_9541,N_9289);
or U10351 (N_10351,N_9373,N_9673);
and U10352 (N_10352,N_9756,N_9776);
nand U10353 (N_10353,N_9372,N_9927);
and U10354 (N_10354,N_9937,N_9601);
or U10355 (N_10355,N_9608,N_9760);
nand U10356 (N_10356,N_9784,N_9852);
nor U10357 (N_10357,N_9733,N_9464);
nand U10358 (N_10358,N_9951,N_9816);
xnor U10359 (N_10359,N_9364,N_9531);
nand U10360 (N_10360,N_9945,N_9849);
nand U10361 (N_10361,N_9573,N_9090);
xor U10362 (N_10362,N_9013,N_9831);
or U10363 (N_10363,N_9103,N_9401);
and U10364 (N_10364,N_9631,N_9998);
nor U10365 (N_10365,N_9752,N_9883);
and U10366 (N_10366,N_9388,N_9500);
nand U10367 (N_10367,N_9694,N_9365);
and U10368 (N_10368,N_9649,N_9827);
or U10369 (N_10369,N_9086,N_9009);
xor U10370 (N_10370,N_9833,N_9623);
and U10371 (N_10371,N_9838,N_9057);
and U10372 (N_10372,N_9821,N_9139);
or U10373 (N_10373,N_9761,N_9167);
and U10374 (N_10374,N_9078,N_9513);
xor U10375 (N_10375,N_9817,N_9307);
and U10376 (N_10376,N_9675,N_9605);
and U10377 (N_10377,N_9819,N_9221);
nor U10378 (N_10378,N_9026,N_9386);
nand U10379 (N_10379,N_9569,N_9851);
nor U10380 (N_10380,N_9297,N_9191);
nand U10381 (N_10381,N_9264,N_9084);
and U10382 (N_10382,N_9616,N_9422);
nor U10383 (N_10383,N_9895,N_9304);
nor U10384 (N_10384,N_9030,N_9532);
or U10385 (N_10385,N_9936,N_9096);
nand U10386 (N_10386,N_9734,N_9639);
nand U10387 (N_10387,N_9327,N_9337);
nor U10388 (N_10388,N_9188,N_9916);
xor U10389 (N_10389,N_9407,N_9001);
nand U10390 (N_10390,N_9368,N_9270);
and U10391 (N_10391,N_9502,N_9441);
or U10392 (N_10392,N_9730,N_9646);
or U10393 (N_10393,N_9552,N_9426);
nand U10394 (N_10394,N_9335,N_9805);
nand U10395 (N_10395,N_9416,N_9226);
and U10396 (N_10396,N_9325,N_9710);
and U10397 (N_10397,N_9070,N_9148);
or U10398 (N_10398,N_9470,N_9114);
nand U10399 (N_10399,N_9846,N_9967);
xor U10400 (N_10400,N_9811,N_9835);
or U10401 (N_10401,N_9526,N_9508);
nor U10402 (N_10402,N_9550,N_9872);
or U10403 (N_10403,N_9566,N_9788);
xor U10404 (N_10404,N_9409,N_9374);
nand U10405 (N_10405,N_9561,N_9381);
nor U10406 (N_10406,N_9330,N_9022);
nor U10407 (N_10407,N_9643,N_9138);
nand U10408 (N_10408,N_9855,N_9966);
nor U10409 (N_10409,N_9503,N_9997);
nor U10410 (N_10410,N_9197,N_9789);
xnor U10411 (N_10411,N_9764,N_9454);
or U10412 (N_10412,N_9121,N_9429);
and U10413 (N_10413,N_9535,N_9520);
nor U10414 (N_10414,N_9112,N_9281);
nor U10415 (N_10415,N_9543,N_9981);
and U10416 (N_10416,N_9008,N_9485);
or U10417 (N_10417,N_9231,N_9453);
or U10418 (N_10418,N_9542,N_9287);
or U10419 (N_10419,N_9360,N_9768);
and U10420 (N_10420,N_9269,N_9182);
or U10421 (N_10421,N_9952,N_9796);
nor U10422 (N_10422,N_9537,N_9705);
xor U10423 (N_10423,N_9918,N_9642);
xnor U10424 (N_10424,N_9844,N_9644);
or U10425 (N_10425,N_9469,N_9203);
or U10426 (N_10426,N_9283,N_9956);
nand U10427 (N_10427,N_9797,N_9946);
or U10428 (N_10428,N_9635,N_9007);
or U10429 (N_10429,N_9239,N_9061);
nor U10430 (N_10430,N_9174,N_9732);
xnor U10431 (N_10431,N_9181,N_9676);
and U10432 (N_10432,N_9324,N_9067);
or U10433 (N_10433,N_9028,N_9711);
nand U10434 (N_10434,N_9886,N_9536);
and U10435 (N_10435,N_9497,N_9491);
and U10436 (N_10436,N_9885,N_9970);
nor U10437 (N_10437,N_9214,N_9721);
and U10438 (N_10438,N_9108,N_9163);
or U10439 (N_10439,N_9449,N_9037);
and U10440 (N_10440,N_9755,N_9399);
nand U10441 (N_10441,N_9113,N_9435);
nor U10442 (N_10442,N_9055,N_9135);
nand U10443 (N_10443,N_9194,N_9397);
xnor U10444 (N_10444,N_9825,N_9548);
xnor U10445 (N_10445,N_9039,N_9384);
and U10446 (N_10446,N_9411,N_9390);
nand U10447 (N_10447,N_9278,N_9973);
nor U10448 (N_10448,N_9035,N_9604);
nand U10449 (N_10449,N_9983,N_9908);
or U10450 (N_10450,N_9319,N_9619);
nand U10451 (N_10451,N_9482,N_9101);
xor U10452 (N_10452,N_9299,N_9638);
xor U10453 (N_10453,N_9380,N_9107);
xor U10454 (N_10454,N_9424,N_9801);
xnor U10455 (N_10455,N_9930,N_9810);
xnor U10456 (N_10456,N_9696,N_9342);
and U10457 (N_10457,N_9159,N_9637);
or U10458 (N_10458,N_9528,N_9425);
nand U10459 (N_10459,N_9617,N_9349);
nand U10460 (N_10460,N_9538,N_9982);
nor U10461 (N_10461,N_9695,N_9909);
nand U10462 (N_10462,N_9934,N_9832);
nand U10463 (N_10463,N_9328,N_9516);
or U10464 (N_10464,N_9220,N_9196);
or U10465 (N_10465,N_9145,N_9551);
or U10466 (N_10466,N_9717,N_9143);
or U10467 (N_10467,N_9658,N_9024);
nand U10468 (N_10468,N_9785,N_9706);
nand U10469 (N_10469,N_9050,N_9083);
xor U10470 (N_10470,N_9615,N_9394);
or U10471 (N_10471,N_9162,N_9522);
nand U10472 (N_10472,N_9889,N_9248);
xor U10473 (N_10473,N_9481,N_9836);
and U10474 (N_10474,N_9612,N_9298);
nand U10475 (N_10475,N_9201,N_9691);
and U10476 (N_10476,N_9595,N_9713);
or U10477 (N_10477,N_9953,N_9780);
nand U10478 (N_10478,N_9155,N_9031);
nor U10479 (N_10479,N_9750,N_9823);
and U10480 (N_10480,N_9893,N_9869);
nor U10481 (N_10481,N_9499,N_9633);
xor U10482 (N_10482,N_9813,N_9690);
and U10483 (N_10483,N_9698,N_9568);
nor U10484 (N_10484,N_9586,N_9317);
nand U10485 (N_10485,N_9301,N_9867);
nand U10486 (N_10486,N_9474,N_9065);
nand U10487 (N_10487,N_9097,N_9549);
and U10488 (N_10488,N_9769,N_9183);
nand U10489 (N_10489,N_9962,N_9406);
and U10490 (N_10490,N_9423,N_9563);
or U10491 (N_10491,N_9053,N_9133);
xnor U10492 (N_10492,N_9685,N_9382);
or U10493 (N_10493,N_9749,N_9064);
xor U10494 (N_10494,N_9593,N_9626);
nor U10495 (N_10495,N_9378,N_9405);
or U10496 (N_10496,N_9545,N_9432);
nand U10497 (N_10497,N_9632,N_9993);
nand U10498 (N_10498,N_9323,N_9931);
or U10499 (N_10499,N_9745,N_9160);
nor U10500 (N_10500,N_9169,N_9274);
nor U10501 (N_10501,N_9445,N_9331);
nor U10502 (N_10502,N_9570,N_9869);
xor U10503 (N_10503,N_9306,N_9695);
or U10504 (N_10504,N_9188,N_9037);
nor U10505 (N_10505,N_9167,N_9432);
nor U10506 (N_10506,N_9393,N_9808);
and U10507 (N_10507,N_9220,N_9569);
nand U10508 (N_10508,N_9404,N_9636);
nor U10509 (N_10509,N_9606,N_9711);
or U10510 (N_10510,N_9370,N_9850);
nor U10511 (N_10511,N_9444,N_9000);
and U10512 (N_10512,N_9182,N_9999);
and U10513 (N_10513,N_9683,N_9194);
and U10514 (N_10514,N_9976,N_9333);
or U10515 (N_10515,N_9922,N_9687);
and U10516 (N_10516,N_9654,N_9902);
nor U10517 (N_10517,N_9461,N_9073);
and U10518 (N_10518,N_9419,N_9116);
or U10519 (N_10519,N_9545,N_9411);
xnor U10520 (N_10520,N_9466,N_9953);
nor U10521 (N_10521,N_9403,N_9694);
and U10522 (N_10522,N_9452,N_9476);
and U10523 (N_10523,N_9532,N_9857);
or U10524 (N_10524,N_9694,N_9417);
or U10525 (N_10525,N_9669,N_9205);
nand U10526 (N_10526,N_9175,N_9981);
nand U10527 (N_10527,N_9786,N_9386);
and U10528 (N_10528,N_9288,N_9986);
and U10529 (N_10529,N_9591,N_9036);
xor U10530 (N_10530,N_9214,N_9994);
xnor U10531 (N_10531,N_9698,N_9152);
nand U10532 (N_10532,N_9600,N_9579);
nor U10533 (N_10533,N_9137,N_9080);
nor U10534 (N_10534,N_9855,N_9568);
xnor U10535 (N_10535,N_9357,N_9407);
nor U10536 (N_10536,N_9359,N_9993);
xor U10537 (N_10537,N_9936,N_9091);
xor U10538 (N_10538,N_9377,N_9018);
and U10539 (N_10539,N_9414,N_9579);
xor U10540 (N_10540,N_9800,N_9555);
xor U10541 (N_10541,N_9486,N_9213);
xnor U10542 (N_10542,N_9266,N_9697);
and U10543 (N_10543,N_9838,N_9476);
xor U10544 (N_10544,N_9134,N_9643);
nor U10545 (N_10545,N_9395,N_9078);
nor U10546 (N_10546,N_9832,N_9528);
and U10547 (N_10547,N_9552,N_9495);
xnor U10548 (N_10548,N_9664,N_9301);
nand U10549 (N_10549,N_9274,N_9509);
and U10550 (N_10550,N_9018,N_9649);
or U10551 (N_10551,N_9152,N_9893);
nand U10552 (N_10552,N_9331,N_9120);
nand U10553 (N_10553,N_9128,N_9530);
nand U10554 (N_10554,N_9013,N_9704);
and U10555 (N_10555,N_9781,N_9002);
nand U10556 (N_10556,N_9992,N_9408);
nor U10557 (N_10557,N_9190,N_9365);
xnor U10558 (N_10558,N_9215,N_9945);
and U10559 (N_10559,N_9942,N_9619);
and U10560 (N_10560,N_9720,N_9334);
nand U10561 (N_10561,N_9786,N_9504);
nand U10562 (N_10562,N_9672,N_9410);
and U10563 (N_10563,N_9813,N_9330);
nor U10564 (N_10564,N_9219,N_9323);
nor U10565 (N_10565,N_9730,N_9215);
nand U10566 (N_10566,N_9255,N_9452);
and U10567 (N_10567,N_9916,N_9119);
and U10568 (N_10568,N_9031,N_9090);
or U10569 (N_10569,N_9301,N_9490);
or U10570 (N_10570,N_9143,N_9608);
xor U10571 (N_10571,N_9237,N_9571);
nor U10572 (N_10572,N_9650,N_9408);
nand U10573 (N_10573,N_9966,N_9941);
or U10574 (N_10574,N_9930,N_9642);
nand U10575 (N_10575,N_9811,N_9980);
and U10576 (N_10576,N_9012,N_9233);
xnor U10577 (N_10577,N_9743,N_9177);
or U10578 (N_10578,N_9494,N_9732);
nand U10579 (N_10579,N_9899,N_9109);
nand U10580 (N_10580,N_9102,N_9049);
xnor U10581 (N_10581,N_9459,N_9660);
nor U10582 (N_10582,N_9774,N_9601);
xor U10583 (N_10583,N_9525,N_9171);
and U10584 (N_10584,N_9739,N_9062);
nor U10585 (N_10585,N_9880,N_9047);
nor U10586 (N_10586,N_9596,N_9406);
xnor U10587 (N_10587,N_9052,N_9558);
xor U10588 (N_10588,N_9631,N_9866);
nand U10589 (N_10589,N_9950,N_9458);
nand U10590 (N_10590,N_9667,N_9518);
xor U10591 (N_10591,N_9215,N_9766);
nand U10592 (N_10592,N_9932,N_9480);
nor U10593 (N_10593,N_9207,N_9640);
xor U10594 (N_10594,N_9709,N_9150);
and U10595 (N_10595,N_9679,N_9917);
and U10596 (N_10596,N_9163,N_9924);
xnor U10597 (N_10597,N_9467,N_9794);
nand U10598 (N_10598,N_9737,N_9628);
and U10599 (N_10599,N_9622,N_9680);
and U10600 (N_10600,N_9894,N_9870);
nor U10601 (N_10601,N_9099,N_9176);
or U10602 (N_10602,N_9591,N_9581);
nand U10603 (N_10603,N_9990,N_9494);
nand U10604 (N_10604,N_9178,N_9050);
or U10605 (N_10605,N_9449,N_9565);
nor U10606 (N_10606,N_9690,N_9190);
nand U10607 (N_10607,N_9051,N_9995);
and U10608 (N_10608,N_9721,N_9532);
and U10609 (N_10609,N_9473,N_9274);
or U10610 (N_10610,N_9903,N_9445);
or U10611 (N_10611,N_9716,N_9588);
or U10612 (N_10612,N_9284,N_9973);
nand U10613 (N_10613,N_9798,N_9278);
nand U10614 (N_10614,N_9090,N_9846);
nor U10615 (N_10615,N_9116,N_9636);
nand U10616 (N_10616,N_9389,N_9584);
nor U10617 (N_10617,N_9371,N_9103);
nor U10618 (N_10618,N_9300,N_9532);
or U10619 (N_10619,N_9927,N_9147);
or U10620 (N_10620,N_9814,N_9642);
xor U10621 (N_10621,N_9784,N_9417);
xor U10622 (N_10622,N_9617,N_9187);
nand U10623 (N_10623,N_9170,N_9717);
nor U10624 (N_10624,N_9897,N_9393);
nand U10625 (N_10625,N_9587,N_9408);
and U10626 (N_10626,N_9569,N_9950);
xnor U10627 (N_10627,N_9956,N_9363);
xor U10628 (N_10628,N_9804,N_9899);
nand U10629 (N_10629,N_9152,N_9106);
xor U10630 (N_10630,N_9523,N_9538);
nor U10631 (N_10631,N_9568,N_9060);
nor U10632 (N_10632,N_9526,N_9738);
nand U10633 (N_10633,N_9790,N_9802);
nand U10634 (N_10634,N_9428,N_9495);
nor U10635 (N_10635,N_9746,N_9900);
and U10636 (N_10636,N_9320,N_9583);
or U10637 (N_10637,N_9960,N_9879);
nor U10638 (N_10638,N_9173,N_9828);
and U10639 (N_10639,N_9744,N_9319);
nor U10640 (N_10640,N_9633,N_9060);
or U10641 (N_10641,N_9741,N_9194);
xor U10642 (N_10642,N_9959,N_9908);
nor U10643 (N_10643,N_9489,N_9116);
or U10644 (N_10644,N_9013,N_9976);
nor U10645 (N_10645,N_9959,N_9583);
nor U10646 (N_10646,N_9241,N_9577);
or U10647 (N_10647,N_9728,N_9151);
nor U10648 (N_10648,N_9615,N_9155);
nand U10649 (N_10649,N_9070,N_9606);
and U10650 (N_10650,N_9685,N_9029);
or U10651 (N_10651,N_9578,N_9310);
nor U10652 (N_10652,N_9954,N_9506);
nor U10653 (N_10653,N_9179,N_9306);
xor U10654 (N_10654,N_9258,N_9765);
nand U10655 (N_10655,N_9414,N_9069);
nand U10656 (N_10656,N_9951,N_9460);
nand U10657 (N_10657,N_9297,N_9861);
xnor U10658 (N_10658,N_9263,N_9016);
nand U10659 (N_10659,N_9747,N_9300);
nand U10660 (N_10660,N_9908,N_9059);
nor U10661 (N_10661,N_9389,N_9159);
xor U10662 (N_10662,N_9789,N_9326);
nand U10663 (N_10663,N_9181,N_9325);
xor U10664 (N_10664,N_9652,N_9202);
or U10665 (N_10665,N_9294,N_9612);
nor U10666 (N_10666,N_9045,N_9319);
nand U10667 (N_10667,N_9617,N_9534);
nor U10668 (N_10668,N_9170,N_9114);
nand U10669 (N_10669,N_9732,N_9353);
xor U10670 (N_10670,N_9573,N_9688);
xnor U10671 (N_10671,N_9699,N_9316);
or U10672 (N_10672,N_9609,N_9123);
and U10673 (N_10673,N_9251,N_9794);
xor U10674 (N_10674,N_9459,N_9007);
and U10675 (N_10675,N_9488,N_9044);
nor U10676 (N_10676,N_9680,N_9985);
nor U10677 (N_10677,N_9802,N_9957);
nand U10678 (N_10678,N_9656,N_9130);
nand U10679 (N_10679,N_9729,N_9367);
or U10680 (N_10680,N_9834,N_9994);
xnor U10681 (N_10681,N_9114,N_9966);
or U10682 (N_10682,N_9963,N_9046);
and U10683 (N_10683,N_9437,N_9844);
nand U10684 (N_10684,N_9476,N_9344);
or U10685 (N_10685,N_9178,N_9051);
nand U10686 (N_10686,N_9696,N_9261);
nor U10687 (N_10687,N_9178,N_9006);
and U10688 (N_10688,N_9522,N_9805);
and U10689 (N_10689,N_9436,N_9664);
xnor U10690 (N_10690,N_9226,N_9453);
and U10691 (N_10691,N_9054,N_9445);
nor U10692 (N_10692,N_9349,N_9452);
nand U10693 (N_10693,N_9847,N_9675);
nor U10694 (N_10694,N_9335,N_9424);
xnor U10695 (N_10695,N_9329,N_9973);
xor U10696 (N_10696,N_9113,N_9534);
nor U10697 (N_10697,N_9700,N_9701);
or U10698 (N_10698,N_9341,N_9946);
nor U10699 (N_10699,N_9207,N_9202);
nand U10700 (N_10700,N_9527,N_9417);
or U10701 (N_10701,N_9598,N_9209);
nor U10702 (N_10702,N_9702,N_9469);
or U10703 (N_10703,N_9354,N_9785);
xnor U10704 (N_10704,N_9709,N_9348);
xor U10705 (N_10705,N_9229,N_9573);
nor U10706 (N_10706,N_9158,N_9423);
xor U10707 (N_10707,N_9081,N_9667);
xnor U10708 (N_10708,N_9175,N_9654);
xor U10709 (N_10709,N_9136,N_9541);
nor U10710 (N_10710,N_9254,N_9482);
nor U10711 (N_10711,N_9538,N_9346);
xnor U10712 (N_10712,N_9947,N_9939);
nor U10713 (N_10713,N_9213,N_9929);
and U10714 (N_10714,N_9475,N_9982);
xnor U10715 (N_10715,N_9481,N_9071);
nand U10716 (N_10716,N_9778,N_9531);
or U10717 (N_10717,N_9653,N_9779);
or U10718 (N_10718,N_9147,N_9224);
xnor U10719 (N_10719,N_9035,N_9181);
nand U10720 (N_10720,N_9153,N_9309);
xor U10721 (N_10721,N_9835,N_9748);
nor U10722 (N_10722,N_9482,N_9243);
nand U10723 (N_10723,N_9553,N_9087);
nor U10724 (N_10724,N_9019,N_9775);
or U10725 (N_10725,N_9757,N_9076);
nand U10726 (N_10726,N_9405,N_9560);
xnor U10727 (N_10727,N_9763,N_9563);
nor U10728 (N_10728,N_9615,N_9661);
xnor U10729 (N_10729,N_9463,N_9872);
and U10730 (N_10730,N_9310,N_9779);
xor U10731 (N_10731,N_9691,N_9501);
or U10732 (N_10732,N_9486,N_9804);
nand U10733 (N_10733,N_9247,N_9245);
or U10734 (N_10734,N_9003,N_9560);
nand U10735 (N_10735,N_9674,N_9336);
nor U10736 (N_10736,N_9361,N_9290);
nor U10737 (N_10737,N_9417,N_9000);
nand U10738 (N_10738,N_9112,N_9352);
nor U10739 (N_10739,N_9751,N_9136);
nor U10740 (N_10740,N_9720,N_9468);
nor U10741 (N_10741,N_9072,N_9690);
and U10742 (N_10742,N_9173,N_9403);
nor U10743 (N_10743,N_9478,N_9548);
xnor U10744 (N_10744,N_9613,N_9708);
xnor U10745 (N_10745,N_9259,N_9907);
or U10746 (N_10746,N_9999,N_9528);
nor U10747 (N_10747,N_9117,N_9809);
xnor U10748 (N_10748,N_9306,N_9208);
and U10749 (N_10749,N_9537,N_9164);
nor U10750 (N_10750,N_9967,N_9297);
xnor U10751 (N_10751,N_9505,N_9445);
and U10752 (N_10752,N_9625,N_9642);
and U10753 (N_10753,N_9614,N_9212);
nor U10754 (N_10754,N_9569,N_9469);
xnor U10755 (N_10755,N_9603,N_9579);
xnor U10756 (N_10756,N_9972,N_9481);
or U10757 (N_10757,N_9967,N_9631);
nor U10758 (N_10758,N_9047,N_9310);
nor U10759 (N_10759,N_9698,N_9335);
and U10760 (N_10760,N_9255,N_9828);
nand U10761 (N_10761,N_9753,N_9710);
and U10762 (N_10762,N_9726,N_9184);
and U10763 (N_10763,N_9583,N_9143);
or U10764 (N_10764,N_9266,N_9449);
nand U10765 (N_10765,N_9975,N_9454);
and U10766 (N_10766,N_9645,N_9261);
nand U10767 (N_10767,N_9209,N_9442);
nor U10768 (N_10768,N_9745,N_9413);
and U10769 (N_10769,N_9138,N_9684);
xnor U10770 (N_10770,N_9875,N_9625);
xnor U10771 (N_10771,N_9273,N_9798);
and U10772 (N_10772,N_9578,N_9378);
nand U10773 (N_10773,N_9044,N_9375);
nor U10774 (N_10774,N_9661,N_9309);
nor U10775 (N_10775,N_9264,N_9618);
nor U10776 (N_10776,N_9463,N_9813);
xnor U10777 (N_10777,N_9756,N_9412);
xnor U10778 (N_10778,N_9001,N_9836);
or U10779 (N_10779,N_9404,N_9641);
nand U10780 (N_10780,N_9510,N_9980);
nand U10781 (N_10781,N_9795,N_9695);
nand U10782 (N_10782,N_9956,N_9991);
nor U10783 (N_10783,N_9083,N_9218);
xnor U10784 (N_10784,N_9623,N_9389);
nor U10785 (N_10785,N_9193,N_9912);
nand U10786 (N_10786,N_9149,N_9568);
and U10787 (N_10787,N_9809,N_9980);
nor U10788 (N_10788,N_9179,N_9996);
nand U10789 (N_10789,N_9955,N_9797);
nand U10790 (N_10790,N_9353,N_9837);
and U10791 (N_10791,N_9027,N_9813);
xor U10792 (N_10792,N_9600,N_9948);
and U10793 (N_10793,N_9208,N_9170);
nor U10794 (N_10794,N_9619,N_9200);
nand U10795 (N_10795,N_9989,N_9006);
nor U10796 (N_10796,N_9076,N_9715);
xnor U10797 (N_10797,N_9050,N_9825);
xnor U10798 (N_10798,N_9665,N_9358);
xor U10799 (N_10799,N_9465,N_9837);
and U10800 (N_10800,N_9390,N_9829);
and U10801 (N_10801,N_9495,N_9259);
xor U10802 (N_10802,N_9098,N_9812);
nand U10803 (N_10803,N_9045,N_9854);
nor U10804 (N_10804,N_9656,N_9881);
xor U10805 (N_10805,N_9265,N_9610);
or U10806 (N_10806,N_9338,N_9892);
xor U10807 (N_10807,N_9401,N_9530);
nand U10808 (N_10808,N_9820,N_9300);
xor U10809 (N_10809,N_9044,N_9176);
or U10810 (N_10810,N_9598,N_9033);
nand U10811 (N_10811,N_9777,N_9480);
and U10812 (N_10812,N_9539,N_9776);
or U10813 (N_10813,N_9716,N_9268);
or U10814 (N_10814,N_9460,N_9270);
nand U10815 (N_10815,N_9994,N_9167);
nor U10816 (N_10816,N_9171,N_9999);
nand U10817 (N_10817,N_9512,N_9696);
nor U10818 (N_10818,N_9030,N_9052);
nand U10819 (N_10819,N_9916,N_9539);
xor U10820 (N_10820,N_9504,N_9247);
or U10821 (N_10821,N_9313,N_9953);
nor U10822 (N_10822,N_9798,N_9928);
or U10823 (N_10823,N_9152,N_9135);
xor U10824 (N_10824,N_9236,N_9962);
and U10825 (N_10825,N_9660,N_9410);
or U10826 (N_10826,N_9931,N_9255);
and U10827 (N_10827,N_9149,N_9895);
nand U10828 (N_10828,N_9098,N_9430);
or U10829 (N_10829,N_9496,N_9747);
and U10830 (N_10830,N_9140,N_9946);
nor U10831 (N_10831,N_9296,N_9519);
xnor U10832 (N_10832,N_9032,N_9391);
nor U10833 (N_10833,N_9725,N_9419);
or U10834 (N_10834,N_9158,N_9966);
nand U10835 (N_10835,N_9224,N_9173);
nor U10836 (N_10836,N_9473,N_9738);
or U10837 (N_10837,N_9420,N_9783);
or U10838 (N_10838,N_9999,N_9816);
nor U10839 (N_10839,N_9779,N_9657);
or U10840 (N_10840,N_9155,N_9000);
nor U10841 (N_10841,N_9584,N_9092);
nand U10842 (N_10842,N_9088,N_9190);
and U10843 (N_10843,N_9325,N_9411);
nand U10844 (N_10844,N_9984,N_9471);
nor U10845 (N_10845,N_9719,N_9094);
and U10846 (N_10846,N_9855,N_9700);
xnor U10847 (N_10847,N_9521,N_9276);
nor U10848 (N_10848,N_9855,N_9179);
nand U10849 (N_10849,N_9619,N_9195);
nand U10850 (N_10850,N_9381,N_9817);
nor U10851 (N_10851,N_9263,N_9965);
or U10852 (N_10852,N_9823,N_9878);
nor U10853 (N_10853,N_9367,N_9214);
and U10854 (N_10854,N_9033,N_9741);
and U10855 (N_10855,N_9274,N_9725);
and U10856 (N_10856,N_9998,N_9851);
nand U10857 (N_10857,N_9479,N_9866);
nand U10858 (N_10858,N_9557,N_9022);
nor U10859 (N_10859,N_9384,N_9314);
nand U10860 (N_10860,N_9415,N_9685);
and U10861 (N_10861,N_9159,N_9320);
and U10862 (N_10862,N_9147,N_9838);
nor U10863 (N_10863,N_9578,N_9730);
xnor U10864 (N_10864,N_9873,N_9147);
nand U10865 (N_10865,N_9858,N_9446);
and U10866 (N_10866,N_9251,N_9642);
or U10867 (N_10867,N_9666,N_9222);
or U10868 (N_10868,N_9682,N_9855);
xnor U10869 (N_10869,N_9648,N_9562);
nand U10870 (N_10870,N_9840,N_9083);
or U10871 (N_10871,N_9748,N_9667);
or U10872 (N_10872,N_9645,N_9753);
xnor U10873 (N_10873,N_9092,N_9629);
and U10874 (N_10874,N_9498,N_9329);
or U10875 (N_10875,N_9939,N_9011);
nor U10876 (N_10876,N_9323,N_9496);
or U10877 (N_10877,N_9137,N_9977);
xor U10878 (N_10878,N_9338,N_9910);
nand U10879 (N_10879,N_9042,N_9483);
nor U10880 (N_10880,N_9013,N_9465);
nand U10881 (N_10881,N_9084,N_9256);
nand U10882 (N_10882,N_9902,N_9850);
or U10883 (N_10883,N_9889,N_9352);
or U10884 (N_10884,N_9475,N_9706);
and U10885 (N_10885,N_9278,N_9046);
xnor U10886 (N_10886,N_9169,N_9245);
nand U10887 (N_10887,N_9099,N_9266);
xnor U10888 (N_10888,N_9542,N_9023);
xor U10889 (N_10889,N_9861,N_9318);
or U10890 (N_10890,N_9413,N_9266);
xor U10891 (N_10891,N_9000,N_9911);
nand U10892 (N_10892,N_9403,N_9599);
and U10893 (N_10893,N_9101,N_9684);
nor U10894 (N_10894,N_9502,N_9081);
nor U10895 (N_10895,N_9252,N_9416);
nand U10896 (N_10896,N_9115,N_9013);
nand U10897 (N_10897,N_9437,N_9352);
and U10898 (N_10898,N_9476,N_9010);
or U10899 (N_10899,N_9246,N_9310);
nor U10900 (N_10900,N_9526,N_9013);
nor U10901 (N_10901,N_9829,N_9837);
and U10902 (N_10902,N_9504,N_9701);
xor U10903 (N_10903,N_9895,N_9052);
and U10904 (N_10904,N_9434,N_9297);
xnor U10905 (N_10905,N_9678,N_9566);
xnor U10906 (N_10906,N_9434,N_9744);
or U10907 (N_10907,N_9562,N_9118);
and U10908 (N_10908,N_9934,N_9514);
xor U10909 (N_10909,N_9248,N_9917);
and U10910 (N_10910,N_9856,N_9744);
nor U10911 (N_10911,N_9642,N_9718);
nor U10912 (N_10912,N_9881,N_9195);
nand U10913 (N_10913,N_9444,N_9449);
and U10914 (N_10914,N_9620,N_9370);
xor U10915 (N_10915,N_9811,N_9867);
xor U10916 (N_10916,N_9555,N_9563);
xor U10917 (N_10917,N_9515,N_9795);
or U10918 (N_10918,N_9313,N_9767);
and U10919 (N_10919,N_9186,N_9279);
nand U10920 (N_10920,N_9712,N_9860);
or U10921 (N_10921,N_9374,N_9881);
or U10922 (N_10922,N_9183,N_9035);
nor U10923 (N_10923,N_9754,N_9659);
nand U10924 (N_10924,N_9881,N_9508);
nor U10925 (N_10925,N_9731,N_9031);
and U10926 (N_10926,N_9118,N_9350);
or U10927 (N_10927,N_9016,N_9854);
and U10928 (N_10928,N_9299,N_9542);
and U10929 (N_10929,N_9383,N_9306);
and U10930 (N_10930,N_9970,N_9897);
or U10931 (N_10931,N_9163,N_9951);
nand U10932 (N_10932,N_9556,N_9258);
nand U10933 (N_10933,N_9046,N_9280);
xor U10934 (N_10934,N_9772,N_9802);
nand U10935 (N_10935,N_9451,N_9228);
xnor U10936 (N_10936,N_9332,N_9930);
xor U10937 (N_10937,N_9120,N_9827);
xor U10938 (N_10938,N_9367,N_9026);
xnor U10939 (N_10939,N_9147,N_9581);
nor U10940 (N_10940,N_9303,N_9576);
nor U10941 (N_10941,N_9064,N_9144);
or U10942 (N_10942,N_9284,N_9232);
and U10943 (N_10943,N_9790,N_9153);
and U10944 (N_10944,N_9413,N_9114);
nor U10945 (N_10945,N_9625,N_9038);
and U10946 (N_10946,N_9669,N_9278);
and U10947 (N_10947,N_9009,N_9333);
and U10948 (N_10948,N_9071,N_9383);
and U10949 (N_10949,N_9785,N_9842);
xnor U10950 (N_10950,N_9683,N_9861);
and U10951 (N_10951,N_9250,N_9814);
or U10952 (N_10952,N_9026,N_9771);
xor U10953 (N_10953,N_9468,N_9505);
nand U10954 (N_10954,N_9152,N_9330);
and U10955 (N_10955,N_9669,N_9241);
and U10956 (N_10956,N_9716,N_9071);
xnor U10957 (N_10957,N_9834,N_9697);
nor U10958 (N_10958,N_9536,N_9949);
nand U10959 (N_10959,N_9052,N_9655);
xnor U10960 (N_10960,N_9115,N_9469);
nor U10961 (N_10961,N_9019,N_9838);
nor U10962 (N_10962,N_9587,N_9754);
or U10963 (N_10963,N_9619,N_9996);
xnor U10964 (N_10964,N_9936,N_9768);
nor U10965 (N_10965,N_9843,N_9262);
nor U10966 (N_10966,N_9890,N_9173);
nor U10967 (N_10967,N_9835,N_9479);
or U10968 (N_10968,N_9336,N_9090);
and U10969 (N_10969,N_9723,N_9235);
xnor U10970 (N_10970,N_9601,N_9371);
and U10971 (N_10971,N_9013,N_9877);
and U10972 (N_10972,N_9872,N_9952);
or U10973 (N_10973,N_9102,N_9982);
xnor U10974 (N_10974,N_9035,N_9362);
or U10975 (N_10975,N_9032,N_9526);
nand U10976 (N_10976,N_9175,N_9005);
nand U10977 (N_10977,N_9333,N_9552);
or U10978 (N_10978,N_9658,N_9091);
or U10979 (N_10979,N_9135,N_9395);
nand U10980 (N_10980,N_9984,N_9580);
and U10981 (N_10981,N_9877,N_9823);
and U10982 (N_10982,N_9708,N_9266);
or U10983 (N_10983,N_9988,N_9446);
and U10984 (N_10984,N_9398,N_9320);
or U10985 (N_10985,N_9104,N_9540);
and U10986 (N_10986,N_9953,N_9479);
xor U10987 (N_10987,N_9353,N_9025);
or U10988 (N_10988,N_9901,N_9309);
xor U10989 (N_10989,N_9487,N_9915);
and U10990 (N_10990,N_9140,N_9227);
or U10991 (N_10991,N_9780,N_9660);
xnor U10992 (N_10992,N_9318,N_9376);
or U10993 (N_10993,N_9598,N_9394);
nand U10994 (N_10994,N_9743,N_9285);
or U10995 (N_10995,N_9706,N_9794);
xnor U10996 (N_10996,N_9032,N_9212);
and U10997 (N_10997,N_9312,N_9845);
or U10998 (N_10998,N_9041,N_9297);
xnor U10999 (N_10999,N_9675,N_9010);
nand U11000 (N_11000,N_10209,N_10776);
or U11001 (N_11001,N_10713,N_10990);
nand U11002 (N_11002,N_10285,N_10965);
and U11003 (N_11003,N_10229,N_10539);
nor U11004 (N_11004,N_10862,N_10097);
or U11005 (N_11005,N_10602,N_10326);
or U11006 (N_11006,N_10944,N_10488);
xnor U11007 (N_11007,N_10305,N_10444);
xnor U11008 (N_11008,N_10096,N_10921);
nor U11009 (N_11009,N_10322,N_10420);
nor U11010 (N_11010,N_10931,N_10119);
nor U11011 (N_11011,N_10727,N_10331);
nor U11012 (N_11012,N_10197,N_10511);
and U11013 (N_11013,N_10695,N_10540);
and U11014 (N_11014,N_10358,N_10378);
or U11015 (N_11015,N_10217,N_10480);
or U11016 (N_11016,N_10479,N_10858);
xor U11017 (N_11017,N_10999,N_10577);
and U11018 (N_11018,N_10430,N_10645);
nor U11019 (N_11019,N_10056,N_10922);
xnor U11020 (N_11020,N_10314,N_10655);
xor U11021 (N_11021,N_10954,N_10110);
xor U11022 (N_11022,N_10049,N_10964);
nand U11023 (N_11023,N_10806,N_10873);
and U11024 (N_11024,N_10886,N_10095);
and U11025 (N_11025,N_10421,N_10158);
or U11026 (N_11026,N_10966,N_10423);
nor U11027 (N_11027,N_10306,N_10971);
and U11028 (N_11028,N_10039,N_10236);
and U11029 (N_11029,N_10061,N_10470);
or U11030 (N_11030,N_10783,N_10477);
xnor U11031 (N_11031,N_10108,N_10203);
nor U11032 (N_11032,N_10397,N_10022);
or U11033 (N_11033,N_10153,N_10215);
xor U11034 (N_11034,N_10652,N_10573);
nand U11035 (N_11035,N_10365,N_10364);
nor U11036 (N_11036,N_10723,N_10431);
nand U11037 (N_11037,N_10004,N_10416);
nor U11038 (N_11038,N_10389,N_10720);
nand U11039 (N_11039,N_10724,N_10002);
nand U11040 (N_11040,N_10237,N_10510);
nor U11041 (N_11041,N_10536,N_10019);
and U11042 (N_11042,N_10796,N_10018);
nand U11043 (N_11043,N_10238,N_10319);
nand U11044 (N_11044,N_10589,N_10294);
xor U11045 (N_11045,N_10026,N_10842);
and U11046 (N_11046,N_10383,N_10140);
xor U11047 (N_11047,N_10731,N_10487);
xnor U11048 (N_11048,N_10504,N_10338);
and U11049 (N_11049,N_10641,N_10586);
or U11050 (N_11050,N_10516,N_10499);
xnor U11051 (N_11051,N_10635,N_10789);
or U11052 (N_11052,N_10846,N_10498);
or U11053 (N_11053,N_10262,N_10376);
nand U11054 (N_11054,N_10975,N_10797);
xnor U11055 (N_11055,N_10054,N_10059);
and U11056 (N_11056,N_10633,N_10067);
nand U11057 (N_11057,N_10979,N_10370);
and U11058 (N_11058,N_10210,N_10472);
nand U11059 (N_11059,N_10085,N_10225);
nand U11060 (N_11060,N_10587,N_10330);
nor U11061 (N_11061,N_10191,N_10801);
and U11062 (N_11062,N_10272,N_10189);
and U11063 (N_11063,N_10742,N_10254);
nor U11064 (N_11064,N_10970,N_10380);
and U11065 (N_11065,N_10277,N_10005);
or U11066 (N_11066,N_10500,N_10893);
nor U11067 (N_11067,N_10768,N_10485);
nor U11068 (N_11068,N_10028,N_10218);
xnor U11069 (N_11069,N_10463,N_10825);
or U11070 (N_11070,N_10164,N_10295);
and U11071 (N_11071,N_10848,N_10875);
nor U11072 (N_11072,N_10402,N_10814);
xor U11073 (N_11073,N_10804,N_10239);
xnor U11074 (N_11074,N_10258,N_10819);
xnor U11075 (N_11075,N_10878,N_10895);
nor U11076 (N_11076,N_10580,N_10696);
nand U11077 (N_11077,N_10055,N_10252);
or U11078 (N_11078,N_10040,N_10943);
or U11079 (N_11079,N_10481,N_10646);
and U11080 (N_11080,N_10777,N_10772);
and U11081 (N_11081,N_10843,N_10601);
nand U11082 (N_11082,N_10951,N_10084);
nand U11083 (N_11083,N_10457,N_10271);
nand U11084 (N_11084,N_10052,N_10057);
and U11085 (N_11085,N_10455,N_10612);
nand U11086 (N_11086,N_10638,N_10029);
nor U11087 (N_11087,N_10839,N_10363);
xor U11088 (N_11088,N_10270,N_10523);
or U11089 (N_11089,N_10637,N_10240);
nor U11090 (N_11090,N_10781,N_10913);
nand U11091 (N_11091,N_10173,N_10766);
or U11092 (N_11092,N_10912,N_10025);
xnor U11093 (N_11093,N_10894,N_10575);
xnor U11094 (N_11094,N_10867,N_10847);
or U11095 (N_11095,N_10991,N_10234);
nor U11096 (N_11096,N_10605,N_10386);
or U11097 (N_11097,N_10442,N_10800);
xor U11098 (N_11098,N_10640,N_10011);
nor U11099 (N_11099,N_10905,N_10930);
nor U11100 (N_11100,N_10593,N_10691);
xnor U11101 (N_11101,N_10547,N_10969);
xnor U11102 (N_11102,N_10856,N_10983);
nand U11103 (N_11103,N_10167,N_10736);
xor U11104 (N_11104,N_10838,N_10245);
xnor U11105 (N_11105,N_10648,N_10268);
and U11106 (N_11106,N_10900,N_10629);
and U11107 (N_11107,N_10687,N_10219);
nand U11108 (N_11108,N_10963,N_10845);
nand U11109 (N_11109,N_10373,N_10161);
and U11110 (N_11110,N_10486,N_10639);
or U11111 (N_11111,N_10413,N_10660);
and U11112 (N_11112,N_10681,N_10279);
nand U11113 (N_11113,N_10955,N_10706);
nor U11114 (N_11114,N_10303,N_10710);
nor U11115 (N_11115,N_10307,N_10206);
and U11116 (N_11116,N_10755,N_10535);
nand U11117 (N_11117,N_10524,N_10497);
xor U11118 (N_11118,N_10773,N_10555);
xnor U11119 (N_11119,N_10574,N_10264);
xnor U11120 (N_11120,N_10348,N_10827);
xor U11121 (N_11121,N_10461,N_10885);
or U11122 (N_11122,N_10948,N_10212);
xnor U11123 (N_11123,N_10630,N_10725);
or U11124 (N_11124,N_10180,N_10143);
or U11125 (N_11125,N_10973,N_10222);
or U11126 (N_11126,N_10447,N_10137);
xor U11127 (N_11127,N_10591,N_10992);
nor U11128 (N_11128,N_10595,N_10767);
nor U11129 (N_11129,N_10419,N_10988);
nor U11130 (N_11130,N_10452,N_10996);
or U11131 (N_11131,N_10293,N_10957);
nand U11132 (N_11132,N_10150,N_10090);
nand U11133 (N_11133,N_10583,N_10074);
or U11134 (N_11134,N_10753,N_10968);
nand U11135 (N_11135,N_10283,N_10065);
nor U11136 (N_11136,N_10513,N_10068);
nand U11137 (N_11137,N_10113,N_10533);
nor U11138 (N_11138,N_10643,N_10906);
nor U11139 (N_11139,N_10947,N_10959);
nor U11140 (N_11140,N_10835,N_10771);
or U11141 (N_11141,N_10897,N_10392);
xor U11142 (N_11142,N_10927,N_10400);
nand U11143 (N_11143,N_10103,N_10746);
nor U11144 (N_11144,N_10989,N_10144);
or U11145 (N_11145,N_10459,N_10501);
nor U11146 (N_11146,N_10749,N_10207);
and U11147 (N_11147,N_10432,N_10571);
or U11148 (N_11148,N_10412,N_10889);
and U11149 (N_11149,N_10024,N_10551);
xnor U11150 (N_11150,N_10344,N_10183);
xnor U11151 (N_11151,N_10978,N_10805);
nand U11152 (N_11152,N_10770,N_10821);
nand U11153 (N_11153,N_10353,N_10266);
and U11154 (N_11154,N_10576,N_10624);
xor U11155 (N_11155,N_10857,N_10558);
nand U11156 (N_11156,N_10142,N_10850);
and U11157 (N_11157,N_10111,N_10122);
nand U11158 (N_11158,N_10661,N_10584);
or U11159 (N_11159,N_10908,N_10078);
xor U11160 (N_11160,N_10154,N_10304);
and U11161 (N_11161,N_10812,N_10786);
or U11162 (N_11162,N_10578,N_10282);
nor U11163 (N_11163,N_10328,N_10077);
nor U11164 (N_11164,N_10977,N_10027);
xor U11165 (N_11165,N_10844,N_10290);
and U11166 (N_11166,N_10828,N_10313);
or U11167 (N_11167,N_10896,N_10355);
xnor U11168 (N_11168,N_10093,N_10087);
or U11169 (N_11169,N_10300,N_10434);
and U11170 (N_11170,N_10393,N_10870);
or U11171 (N_11171,N_10302,N_10834);
or U11172 (N_11172,N_10851,N_10009);
nand U11173 (N_11173,N_10717,N_10903);
and U11174 (N_11174,N_10932,N_10853);
nor U11175 (N_11175,N_10548,N_10426);
nand U11176 (N_11176,N_10615,N_10631);
nor U11177 (N_11177,N_10923,N_10956);
nor U11178 (N_11178,N_10817,N_10179);
nand U11179 (N_11179,N_10483,N_10404);
nand U11180 (N_11180,N_10045,N_10565);
nand U11181 (N_11181,N_10133,N_10686);
xor U11182 (N_11182,N_10634,N_10642);
or U11183 (N_11183,N_10942,N_10650);
and U11184 (N_11184,N_10334,N_10663);
nand U11185 (N_11185,N_10610,N_10337);
and U11186 (N_11186,N_10360,N_10280);
xnor U11187 (N_11187,N_10220,N_10545);
nand U11188 (N_11188,N_10891,N_10403);
nand U11189 (N_11189,N_10157,N_10861);
and U11190 (N_11190,N_10714,N_10803);
or U11191 (N_11191,N_10739,N_10833);
nor U11192 (N_11192,N_10456,N_10445);
or U11193 (N_11193,N_10323,N_10950);
nand U11194 (N_11194,N_10410,N_10566);
xnor U11195 (N_11195,N_10037,N_10744);
or U11196 (N_11196,N_10916,N_10181);
nand U11197 (N_11197,N_10060,N_10134);
nor U11198 (N_11198,N_10721,N_10155);
nor U11199 (N_11199,N_10976,N_10582);
nor U11200 (N_11200,N_10538,N_10118);
and U11201 (N_11201,N_10530,N_10146);
xnor U11202 (N_11202,N_10675,N_10429);
nand U11203 (N_11203,N_10438,N_10176);
nand U11204 (N_11204,N_10993,N_10572);
or U11205 (N_11205,N_10274,N_10518);
and U11206 (N_11206,N_10168,N_10709);
nand U11207 (N_11207,N_10347,N_10756);
nand U11208 (N_11208,N_10604,N_10104);
xor U11209 (N_11209,N_10531,N_10564);
and U11210 (N_11210,N_10126,N_10899);
and U11211 (N_11211,N_10417,N_10299);
nand U11212 (N_11212,N_10815,N_10354);
nand U11213 (N_11213,N_10961,N_10178);
and U11214 (N_11214,N_10329,N_10131);
nand U11215 (N_11215,N_10123,N_10798);
nor U11216 (N_11216,N_10705,N_10737);
or U11217 (N_11217,N_10849,N_10933);
or U11218 (N_11218,N_10936,N_10086);
nand U11219 (N_11219,N_10831,N_10339);
or U11220 (N_11220,N_10958,N_10865);
xor U11221 (N_11221,N_10255,N_10070);
or U11222 (N_11222,N_10351,N_10647);
xor U11223 (N_11223,N_10379,N_10081);
xnor U11224 (N_11224,N_10408,N_10120);
and U11225 (N_11225,N_10046,N_10658);
nor U11226 (N_11226,N_10596,N_10273);
or U11227 (N_11227,N_10139,N_10301);
xnor U11228 (N_11228,N_10945,N_10507);
nor U11229 (N_11229,N_10107,N_10187);
or U11230 (N_11230,N_10361,N_10414);
nor U11231 (N_11231,N_10424,N_10382);
or U11232 (N_11232,N_10678,N_10163);
or U11233 (N_11233,N_10017,N_10008);
nand U11234 (N_11234,N_10779,N_10855);
xor U11235 (N_11235,N_10553,N_10269);
xnor U11236 (N_11236,N_10309,N_10112);
or U11237 (N_11237,N_10000,N_10676);
xnor U11238 (N_11238,N_10882,N_10053);
and U11239 (N_11239,N_10909,N_10907);
nor U11240 (N_11240,N_10275,N_10115);
or U11241 (N_11241,N_10911,N_10474);
nand U11242 (N_11242,N_10836,N_10047);
xor U11243 (N_11243,N_10685,N_10454);
or U11244 (N_11244,N_10101,N_10559);
and U11245 (N_11245,N_10816,N_10719);
nand U11246 (N_11246,N_10117,N_10433);
nand U11247 (N_11247,N_10888,N_10223);
or U11248 (N_11248,N_10038,N_10367);
or U11249 (N_11249,N_10121,N_10341);
and U11250 (N_11250,N_10261,N_10418);
nand U11251 (N_11251,N_10830,N_10509);
nand U11252 (N_11252,N_10297,N_10716);
nor U11253 (N_11253,N_10628,N_10048);
nor U11254 (N_11254,N_10974,N_10561);
nor U11255 (N_11255,N_10464,N_10625);
or U11256 (N_11256,N_10741,N_10473);
nor U11257 (N_11257,N_10763,N_10669);
and U11258 (N_11258,N_10734,N_10357);
nand U11259 (N_11259,N_10792,N_10193);
nor U11260 (N_11260,N_10063,N_10073);
nor U11261 (N_11261,N_10918,N_10259);
nand U11262 (N_11262,N_10491,N_10879);
and U11263 (N_11263,N_10822,N_10984);
xor U11264 (N_11264,N_10995,N_10106);
nand U11265 (N_11265,N_10791,N_10257);
xnor U11266 (N_11266,N_10287,N_10760);
xor U11267 (N_11267,N_10682,N_10529);
nor U11268 (N_11268,N_10042,N_10920);
nand U11269 (N_11269,N_10621,N_10832);
xor U11270 (N_11270,N_10177,N_10315);
xor U11271 (N_11271,N_10672,N_10441);
and U11272 (N_11272,N_10785,N_10190);
and U11273 (N_11273,N_10352,N_10928);
nor U11274 (N_11274,N_10636,N_10369);
nand U11275 (N_11275,N_10415,N_10010);
nand U11276 (N_11276,N_10953,N_10608);
nor U11277 (N_11277,N_10289,N_10493);
nand U11278 (N_11278,N_10693,N_10128);
or U11279 (N_11279,N_10752,N_10651);
nor U11280 (N_11280,N_10409,N_10864);
nor U11281 (N_11281,N_10626,N_10016);
xnor U11282 (N_11282,N_10230,N_10278);
nand U11283 (N_11283,N_10892,N_10708);
xor U11284 (N_11284,N_10506,N_10544);
xor U11285 (N_11285,N_10715,N_10823);
and U11286 (N_11286,N_10689,N_10508);
and U11287 (N_11287,N_10592,N_10915);
and U11288 (N_11288,N_10939,N_10680);
nor U11289 (N_11289,N_10050,N_10435);
nor U11290 (N_11290,N_10649,N_10136);
and U11291 (N_11291,N_10482,N_10324);
and U11292 (N_11292,N_10549,N_10492);
nor U11293 (N_11293,N_10079,N_10664);
nor U11294 (N_11294,N_10703,N_10585);
nand U11295 (N_11295,N_10694,N_10860);
and U11296 (N_11296,N_10526,N_10023);
nand U11297 (N_11297,N_10058,N_10102);
xor U11298 (N_11298,N_10044,N_10759);
or U11299 (N_11299,N_10099,N_10233);
nand U11300 (N_11300,N_10124,N_10151);
and U11301 (N_11301,N_10898,N_10674);
nor U11302 (N_11302,N_10762,N_10632);
xnor U11303 (N_11303,N_10914,N_10072);
nor U11304 (N_11304,N_10250,N_10793);
or U11305 (N_11305,N_10877,N_10901);
nand U11306 (N_11306,N_10904,N_10554);
or U11307 (N_11307,N_10033,N_10406);
or U11308 (N_11308,N_10728,N_10449);
and U11309 (N_11309,N_10671,N_10761);
or U11310 (N_11310,N_10006,N_10618);
nor U11311 (N_11311,N_10296,N_10611);
xnor U11312 (N_11312,N_10665,N_10105);
or U11313 (N_11313,N_10562,N_10982);
nor U11314 (N_11314,N_10623,N_10679);
nor U11315 (N_11315,N_10228,N_10556);
nor U11316 (N_11316,N_10246,N_10702);
or U11317 (N_11317,N_10439,N_10644);
nor U11318 (N_11318,N_10826,N_10350);
nor U11319 (N_11319,N_10949,N_10606);
nor U11320 (N_11320,N_10043,N_10659);
nand U11321 (N_11321,N_10195,N_10778);
nor U11322 (N_11322,N_10541,N_10311);
nand U11323 (N_11323,N_10824,N_10467);
xnor U11324 (N_11324,N_10138,N_10799);
or U11325 (N_11325,N_10820,N_10597);
nor U11326 (N_11326,N_10567,N_10581);
nand U11327 (N_11327,N_10469,N_10780);
xor U11328 (N_11328,N_10325,N_10490);
and U11329 (N_11329,N_10733,N_10654);
nand U11330 (N_11330,N_10747,N_10732);
nand U11331 (N_11331,N_10460,N_10041);
nand U11332 (N_11332,N_10829,N_10598);
or U11333 (N_11333,N_10071,N_10868);
or U11334 (N_11334,N_10080,N_10722);
xnor U11335 (N_11335,N_10711,N_10205);
nor U11336 (N_11336,N_10162,N_10211);
or U11337 (N_11337,N_10251,N_10098);
or U11338 (N_11338,N_10308,N_10349);
nor U11339 (N_11339,N_10557,N_10818);
and U11340 (N_11340,N_10570,N_10613);
xnor U11341 (N_11341,N_10662,N_10869);
xnor U11342 (N_11342,N_10377,N_10226);
nor U11343 (N_11343,N_10863,N_10147);
and U11344 (N_11344,N_10385,N_10148);
nand U11345 (N_11345,N_10787,N_10532);
xor U11346 (N_11346,N_10552,N_10405);
nor U11347 (N_11347,N_10468,N_10462);
or U11348 (N_11348,N_10284,N_10698);
and U11349 (N_11349,N_10465,N_10244);
nand U11350 (N_11350,N_10204,N_10013);
nor U11351 (N_11351,N_10852,N_10960);
nand U11352 (N_11352,N_10866,N_10398);
and U11353 (N_11353,N_10216,N_10336);
nor U11354 (N_11354,N_10346,N_10001);
or U11355 (N_11355,N_10020,N_10619);
nor U11356 (N_11356,N_10871,N_10366);
or U11357 (N_11357,N_10670,N_10627);
and U11358 (N_11358,N_10256,N_10503);
xnor U11359 (N_11359,N_10356,N_10436);
nor U11360 (N_11360,N_10014,N_10345);
xor U11361 (N_11361,N_10840,N_10034);
nor U11362 (N_11362,N_10242,N_10458);
nor U11363 (N_11363,N_10395,N_10224);
and U11364 (N_11364,N_10075,N_10542);
xor U11365 (N_11365,N_10253,N_10129);
xnor U11366 (N_11366,N_10145,N_10740);
nor U11367 (N_11367,N_10902,N_10534);
nand U11368 (N_11368,N_10769,N_10496);
nor U11369 (N_11369,N_10286,N_10750);
and U11370 (N_11370,N_10192,N_10880);
xnor U11371 (N_11371,N_10396,N_10451);
nand U11372 (N_11372,N_10495,N_10288);
nand U11373 (N_11373,N_10962,N_10166);
or U11374 (N_11374,N_10517,N_10765);
nor U11375 (N_11375,N_10281,N_10764);
nand U11376 (N_11376,N_10653,N_10298);
nor U11377 (N_11377,N_10069,N_10340);
xor U11378 (N_11378,N_10657,N_10795);
and U11379 (N_11379,N_10332,N_10489);
and U11380 (N_11380,N_10925,N_10590);
or U11381 (N_11381,N_10094,N_10007);
nor U11382 (N_11382,N_10730,N_10381);
or U11383 (N_11383,N_10872,N_10673);
xor U11384 (N_11384,N_10175,N_10617);
or U11385 (N_11385,N_10446,N_10726);
and U11386 (N_11386,N_10428,N_10335);
xor U11387 (N_11387,N_10550,N_10917);
xor U11388 (N_11388,N_10701,N_10616);
and U11389 (N_11389,N_10291,N_10841);
nor U11390 (N_11390,N_10076,N_10937);
nand U11391 (N_11391,N_10656,N_10876);
or U11392 (N_11392,N_10327,N_10036);
or U11393 (N_11393,N_10267,N_10667);
nand U11394 (N_11394,N_10807,N_10114);
or U11395 (N_11395,N_10362,N_10152);
nand U11396 (N_11396,N_10707,N_10666);
nand U11397 (N_11397,N_10375,N_10994);
nor U11398 (N_11398,N_10172,N_10135);
or U11399 (N_11399,N_10515,N_10374);
xnor U11400 (N_11400,N_10312,N_10609);
or U11401 (N_11401,N_10924,N_10919);
nor U11402 (N_11402,N_10089,N_10031);
and U11403 (N_11403,N_10015,N_10998);
or U11404 (N_11404,N_10184,N_10310);
xnor U11405 (N_11405,N_10321,N_10425);
or U11406 (N_11406,N_10171,N_10697);
xor U11407 (N_11407,N_10132,N_10929);
and U11408 (N_11408,N_10109,N_10884);
nand U11409 (N_11409,N_10088,N_10247);
nand U11410 (N_11410,N_10064,N_10437);
nand U11411 (N_11411,N_10484,N_10494);
nor U11412 (N_11412,N_10668,N_10519);
nor U11413 (N_11413,N_10475,N_10692);
or U11414 (N_11414,N_10704,N_10248);
or U11415 (N_11415,N_10521,N_10188);
xnor U11416 (N_11416,N_10837,N_10359);
xnor U11417 (N_11417,N_10265,N_10520);
and U11418 (N_11418,N_10182,N_10712);
and U11419 (N_11419,N_10387,N_10603);
nand U11420 (N_11420,N_10450,N_10260);
or U11421 (N_11421,N_10677,N_10407);
xor U11422 (N_11422,N_10790,N_10607);
nor U11423 (N_11423,N_10940,N_10802);
and U11424 (N_11424,N_10318,N_10276);
xnor U11425 (N_11425,N_10688,N_10718);
or U11426 (N_11426,N_10091,N_10743);
or U11427 (N_11427,N_10092,N_10141);
nor U11428 (N_11428,N_10537,N_10569);
xnor U11429 (N_11429,N_10985,N_10149);
and U11430 (N_11430,N_10788,N_10967);
nor U11431 (N_11431,N_10810,N_10343);
or U11432 (N_11432,N_10774,N_10185);
nand U11433 (N_11433,N_10476,N_10887);
nor U11434 (N_11434,N_10729,N_10174);
and U11435 (N_11435,N_10232,N_10169);
xnor U11436 (N_11436,N_10754,N_10745);
or U11437 (N_11437,N_10525,N_10030);
nand U11438 (N_11438,N_10201,N_10941);
or U11439 (N_11439,N_10859,N_10411);
and U11440 (N_11440,N_10620,N_10292);
and U11441 (N_11441,N_10987,N_10594);
and U11442 (N_11442,N_10316,N_10116);
and U11443 (N_11443,N_10391,N_10588);
nor U11444 (N_11444,N_10231,N_10599);
nand U11445 (N_11445,N_10125,N_10874);
nor U11446 (N_11446,N_10952,N_10546);
or U11447 (N_11447,N_10758,N_10127);
and U11448 (N_11448,N_10735,N_10478);
or U11449 (N_11449,N_10809,N_10249);
nor U11450 (N_11450,N_10213,N_10563);
or U11451 (N_11451,N_10156,N_10399);
or U11452 (N_11452,N_10981,N_10051);
and U11453 (N_11453,N_10683,N_10471);
or U11454 (N_11454,N_10198,N_10738);
xor U11455 (N_11455,N_10502,N_10986);
nor U11456 (N_11456,N_10946,N_10522);
nor U11457 (N_11457,N_10980,N_10221);
and U11458 (N_11458,N_10782,N_10579);
or U11459 (N_11459,N_10320,N_10775);
or U11460 (N_11460,N_10200,N_10699);
nor U11461 (N_11461,N_10684,N_10700);
and U11462 (N_11462,N_10194,N_10202);
xor U11463 (N_11463,N_10890,N_10243);
nand U11464 (N_11464,N_10186,N_10160);
or U11465 (N_11465,N_10568,N_10165);
nor U11466 (N_11466,N_10935,N_10512);
and U11467 (N_11467,N_10443,N_10066);
nand U11468 (N_11468,N_10241,N_10757);
nand U11469 (N_11469,N_10368,N_10448);
xnor U11470 (N_11470,N_10813,N_10372);
nor U11471 (N_11471,N_10384,N_10938);
nor U11472 (N_11472,N_10159,N_10012);
nor U11473 (N_11473,N_10342,N_10401);
nor U11474 (N_11474,N_10881,N_10371);
or U11475 (N_11475,N_10263,N_10910);
or U11476 (N_11476,N_10748,N_10440);
and U11477 (N_11477,N_10130,N_10527);
nor U11478 (N_11478,N_10543,N_10227);
nand U11479 (N_11479,N_10003,N_10214);
xnor U11480 (N_11480,N_10208,N_10528);
and U11481 (N_11481,N_10062,N_10082);
nand U11482 (N_11482,N_10466,N_10317);
or U11483 (N_11483,N_10196,N_10514);
or U11484 (N_11484,N_10811,N_10751);
xnor U11485 (N_11485,N_10199,N_10035);
xor U11486 (N_11486,N_10333,N_10926);
nand U11487 (N_11487,N_10934,N_10390);
or U11488 (N_11488,N_10784,N_10972);
or U11489 (N_11489,N_10883,N_10808);
or U11490 (N_11490,N_10394,N_10997);
or U11491 (N_11491,N_10505,N_10600);
nand U11492 (N_11492,N_10422,N_10170);
or U11493 (N_11493,N_10622,N_10427);
nand U11494 (N_11494,N_10854,N_10690);
xor U11495 (N_11495,N_10021,N_10100);
xnor U11496 (N_11496,N_10560,N_10083);
nor U11497 (N_11497,N_10453,N_10032);
nand U11498 (N_11498,N_10235,N_10794);
or U11499 (N_11499,N_10614,N_10388);
or U11500 (N_11500,N_10817,N_10018);
and U11501 (N_11501,N_10662,N_10669);
nand U11502 (N_11502,N_10859,N_10935);
xnor U11503 (N_11503,N_10742,N_10895);
or U11504 (N_11504,N_10712,N_10136);
nand U11505 (N_11505,N_10954,N_10647);
nand U11506 (N_11506,N_10798,N_10873);
or U11507 (N_11507,N_10373,N_10095);
and U11508 (N_11508,N_10340,N_10849);
or U11509 (N_11509,N_10693,N_10238);
or U11510 (N_11510,N_10343,N_10591);
xnor U11511 (N_11511,N_10343,N_10242);
or U11512 (N_11512,N_10400,N_10485);
xnor U11513 (N_11513,N_10149,N_10631);
xor U11514 (N_11514,N_10617,N_10180);
nor U11515 (N_11515,N_10727,N_10685);
nor U11516 (N_11516,N_10490,N_10095);
xor U11517 (N_11517,N_10219,N_10077);
or U11518 (N_11518,N_10820,N_10561);
nand U11519 (N_11519,N_10918,N_10291);
xor U11520 (N_11520,N_10889,N_10436);
and U11521 (N_11521,N_10198,N_10629);
and U11522 (N_11522,N_10401,N_10668);
or U11523 (N_11523,N_10526,N_10002);
or U11524 (N_11524,N_10560,N_10749);
nand U11525 (N_11525,N_10404,N_10534);
or U11526 (N_11526,N_10625,N_10499);
nand U11527 (N_11527,N_10743,N_10740);
xor U11528 (N_11528,N_10870,N_10848);
or U11529 (N_11529,N_10999,N_10118);
nand U11530 (N_11530,N_10458,N_10476);
xor U11531 (N_11531,N_10618,N_10743);
nor U11532 (N_11532,N_10882,N_10986);
and U11533 (N_11533,N_10185,N_10405);
xnor U11534 (N_11534,N_10547,N_10630);
or U11535 (N_11535,N_10592,N_10892);
nand U11536 (N_11536,N_10081,N_10896);
and U11537 (N_11537,N_10784,N_10309);
nor U11538 (N_11538,N_10500,N_10256);
or U11539 (N_11539,N_10644,N_10570);
nor U11540 (N_11540,N_10824,N_10735);
and U11541 (N_11541,N_10344,N_10180);
nand U11542 (N_11542,N_10071,N_10495);
nor U11543 (N_11543,N_10178,N_10376);
and U11544 (N_11544,N_10219,N_10514);
and U11545 (N_11545,N_10009,N_10364);
or U11546 (N_11546,N_10715,N_10924);
nand U11547 (N_11547,N_10524,N_10031);
nand U11548 (N_11548,N_10799,N_10363);
xnor U11549 (N_11549,N_10927,N_10243);
nor U11550 (N_11550,N_10538,N_10275);
nor U11551 (N_11551,N_10827,N_10968);
xnor U11552 (N_11552,N_10358,N_10377);
nand U11553 (N_11553,N_10064,N_10457);
or U11554 (N_11554,N_10728,N_10210);
nor U11555 (N_11555,N_10224,N_10351);
nand U11556 (N_11556,N_10717,N_10013);
and U11557 (N_11557,N_10085,N_10787);
nand U11558 (N_11558,N_10375,N_10219);
and U11559 (N_11559,N_10265,N_10377);
xnor U11560 (N_11560,N_10577,N_10296);
nand U11561 (N_11561,N_10209,N_10842);
xor U11562 (N_11562,N_10353,N_10929);
nand U11563 (N_11563,N_10769,N_10497);
nor U11564 (N_11564,N_10100,N_10727);
xnor U11565 (N_11565,N_10661,N_10237);
and U11566 (N_11566,N_10101,N_10425);
and U11567 (N_11567,N_10156,N_10904);
nor U11568 (N_11568,N_10435,N_10644);
or U11569 (N_11569,N_10508,N_10651);
nor U11570 (N_11570,N_10228,N_10438);
nor U11571 (N_11571,N_10434,N_10718);
and U11572 (N_11572,N_10498,N_10838);
and U11573 (N_11573,N_10428,N_10934);
or U11574 (N_11574,N_10980,N_10691);
or U11575 (N_11575,N_10004,N_10531);
nand U11576 (N_11576,N_10100,N_10939);
nand U11577 (N_11577,N_10651,N_10653);
and U11578 (N_11578,N_10749,N_10046);
nand U11579 (N_11579,N_10864,N_10210);
and U11580 (N_11580,N_10891,N_10226);
nor U11581 (N_11581,N_10148,N_10909);
nor U11582 (N_11582,N_10560,N_10677);
nand U11583 (N_11583,N_10104,N_10239);
and U11584 (N_11584,N_10471,N_10925);
and U11585 (N_11585,N_10480,N_10766);
or U11586 (N_11586,N_10973,N_10604);
nor U11587 (N_11587,N_10595,N_10846);
nor U11588 (N_11588,N_10761,N_10301);
and U11589 (N_11589,N_10855,N_10081);
nand U11590 (N_11590,N_10386,N_10097);
xnor U11591 (N_11591,N_10197,N_10085);
xnor U11592 (N_11592,N_10287,N_10993);
nor U11593 (N_11593,N_10694,N_10768);
and U11594 (N_11594,N_10621,N_10268);
and U11595 (N_11595,N_10684,N_10400);
xnor U11596 (N_11596,N_10226,N_10277);
and U11597 (N_11597,N_10371,N_10582);
nor U11598 (N_11598,N_10646,N_10430);
nand U11599 (N_11599,N_10799,N_10559);
or U11600 (N_11600,N_10684,N_10707);
and U11601 (N_11601,N_10954,N_10600);
nand U11602 (N_11602,N_10774,N_10193);
nand U11603 (N_11603,N_10762,N_10214);
nor U11604 (N_11604,N_10061,N_10833);
xor U11605 (N_11605,N_10257,N_10631);
xor U11606 (N_11606,N_10618,N_10315);
nand U11607 (N_11607,N_10591,N_10691);
nor U11608 (N_11608,N_10265,N_10685);
xnor U11609 (N_11609,N_10560,N_10534);
and U11610 (N_11610,N_10577,N_10233);
nand U11611 (N_11611,N_10772,N_10672);
xnor U11612 (N_11612,N_10928,N_10880);
or U11613 (N_11613,N_10013,N_10118);
nor U11614 (N_11614,N_10221,N_10273);
xnor U11615 (N_11615,N_10988,N_10914);
and U11616 (N_11616,N_10009,N_10307);
xnor U11617 (N_11617,N_10954,N_10283);
and U11618 (N_11618,N_10926,N_10653);
and U11619 (N_11619,N_10398,N_10737);
xor U11620 (N_11620,N_10486,N_10389);
nor U11621 (N_11621,N_10491,N_10793);
nand U11622 (N_11622,N_10919,N_10250);
xor U11623 (N_11623,N_10711,N_10226);
and U11624 (N_11624,N_10461,N_10531);
or U11625 (N_11625,N_10617,N_10144);
nand U11626 (N_11626,N_10010,N_10586);
nand U11627 (N_11627,N_10129,N_10542);
nor U11628 (N_11628,N_10900,N_10836);
nand U11629 (N_11629,N_10154,N_10087);
xor U11630 (N_11630,N_10971,N_10035);
xor U11631 (N_11631,N_10692,N_10188);
xnor U11632 (N_11632,N_10003,N_10605);
nand U11633 (N_11633,N_10898,N_10979);
or U11634 (N_11634,N_10534,N_10222);
nor U11635 (N_11635,N_10028,N_10812);
and U11636 (N_11636,N_10138,N_10587);
xor U11637 (N_11637,N_10797,N_10587);
nor U11638 (N_11638,N_10520,N_10910);
or U11639 (N_11639,N_10090,N_10958);
nor U11640 (N_11640,N_10880,N_10131);
xor U11641 (N_11641,N_10165,N_10809);
nor U11642 (N_11642,N_10622,N_10270);
or U11643 (N_11643,N_10499,N_10410);
nor U11644 (N_11644,N_10558,N_10988);
and U11645 (N_11645,N_10507,N_10993);
and U11646 (N_11646,N_10507,N_10654);
nor U11647 (N_11647,N_10053,N_10336);
nor U11648 (N_11648,N_10105,N_10136);
and U11649 (N_11649,N_10612,N_10209);
nor U11650 (N_11650,N_10396,N_10585);
nor U11651 (N_11651,N_10675,N_10621);
nor U11652 (N_11652,N_10365,N_10669);
nor U11653 (N_11653,N_10549,N_10028);
nor U11654 (N_11654,N_10294,N_10817);
or U11655 (N_11655,N_10490,N_10213);
nand U11656 (N_11656,N_10349,N_10740);
or U11657 (N_11657,N_10311,N_10222);
or U11658 (N_11658,N_10249,N_10753);
or U11659 (N_11659,N_10402,N_10311);
xnor U11660 (N_11660,N_10164,N_10356);
or U11661 (N_11661,N_10537,N_10454);
nand U11662 (N_11662,N_10494,N_10956);
nor U11663 (N_11663,N_10329,N_10207);
xnor U11664 (N_11664,N_10942,N_10189);
nor U11665 (N_11665,N_10452,N_10391);
xnor U11666 (N_11666,N_10671,N_10171);
nor U11667 (N_11667,N_10504,N_10466);
xnor U11668 (N_11668,N_10146,N_10603);
nor U11669 (N_11669,N_10356,N_10558);
nand U11670 (N_11670,N_10619,N_10363);
xor U11671 (N_11671,N_10200,N_10123);
nand U11672 (N_11672,N_10775,N_10873);
nand U11673 (N_11673,N_10428,N_10457);
or U11674 (N_11674,N_10250,N_10961);
and U11675 (N_11675,N_10075,N_10288);
and U11676 (N_11676,N_10150,N_10302);
nor U11677 (N_11677,N_10907,N_10781);
nand U11678 (N_11678,N_10870,N_10066);
nor U11679 (N_11679,N_10627,N_10071);
or U11680 (N_11680,N_10084,N_10255);
xnor U11681 (N_11681,N_10506,N_10968);
xor U11682 (N_11682,N_10736,N_10187);
nor U11683 (N_11683,N_10114,N_10366);
nand U11684 (N_11684,N_10351,N_10804);
xnor U11685 (N_11685,N_10139,N_10778);
and U11686 (N_11686,N_10034,N_10943);
nand U11687 (N_11687,N_10950,N_10507);
or U11688 (N_11688,N_10892,N_10625);
nor U11689 (N_11689,N_10249,N_10580);
xor U11690 (N_11690,N_10130,N_10178);
nand U11691 (N_11691,N_10633,N_10652);
and U11692 (N_11692,N_10199,N_10230);
nor U11693 (N_11693,N_10270,N_10228);
and U11694 (N_11694,N_10674,N_10369);
nand U11695 (N_11695,N_10375,N_10831);
xnor U11696 (N_11696,N_10490,N_10530);
nand U11697 (N_11697,N_10049,N_10342);
nand U11698 (N_11698,N_10337,N_10480);
and U11699 (N_11699,N_10142,N_10052);
xor U11700 (N_11700,N_10823,N_10665);
and U11701 (N_11701,N_10985,N_10662);
and U11702 (N_11702,N_10257,N_10307);
nand U11703 (N_11703,N_10693,N_10980);
nand U11704 (N_11704,N_10643,N_10965);
or U11705 (N_11705,N_10596,N_10262);
nor U11706 (N_11706,N_10418,N_10360);
and U11707 (N_11707,N_10532,N_10674);
nor U11708 (N_11708,N_10407,N_10805);
or U11709 (N_11709,N_10378,N_10264);
nand U11710 (N_11710,N_10452,N_10270);
nand U11711 (N_11711,N_10257,N_10822);
xnor U11712 (N_11712,N_10824,N_10701);
nand U11713 (N_11713,N_10965,N_10087);
and U11714 (N_11714,N_10780,N_10579);
nor U11715 (N_11715,N_10483,N_10880);
or U11716 (N_11716,N_10682,N_10432);
or U11717 (N_11717,N_10713,N_10511);
or U11718 (N_11718,N_10925,N_10361);
nand U11719 (N_11719,N_10007,N_10817);
xnor U11720 (N_11720,N_10627,N_10368);
nor U11721 (N_11721,N_10201,N_10546);
or U11722 (N_11722,N_10591,N_10496);
xor U11723 (N_11723,N_10752,N_10446);
xor U11724 (N_11724,N_10698,N_10381);
and U11725 (N_11725,N_10628,N_10475);
xor U11726 (N_11726,N_10106,N_10235);
nor U11727 (N_11727,N_10955,N_10878);
nand U11728 (N_11728,N_10469,N_10905);
nand U11729 (N_11729,N_10671,N_10889);
nor U11730 (N_11730,N_10592,N_10464);
nor U11731 (N_11731,N_10842,N_10862);
and U11732 (N_11732,N_10151,N_10301);
and U11733 (N_11733,N_10153,N_10721);
xnor U11734 (N_11734,N_10435,N_10620);
xor U11735 (N_11735,N_10140,N_10306);
or U11736 (N_11736,N_10325,N_10231);
nand U11737 (N_11737,N_10296,N_10302);
and U11738 (N_11738,N_10557,N_10959);
xnor U11739 (N_11739,N_10190,N_10401);
nor U11740 (N_11740,N_10672,N_10777);
nor U11741 (N_11741,N_10212,N_10234);
or U11742 (N_11742,N_10461,N_10497);
and U11743 (N_11743,N_10260,N_10782);
xnor U11744 (N_11744,N_10164,N_10281);
xor U11745 (N_11745,N_10394,N_10175);
nor U11746 (N_11746,N_10792,N_10485);
nand U11747 (N_11747,N_10128,N_10618);
and U11748 (N_11748,N_10770,N_10328);
nor U11749 (N_11749,N_10466,N_10443);
and U11750 (N_11750,N_10900,N_10534);
or U11751 (N_11751,N_10127,N_10751);
xor U11752 (N_11752,N_10689,N_10132);
and U11753 (N_11753,N_10675,N_10925);
nand U11754 (N_11754,N_10323,N_10481);
and U11755 (N_11755,N_10759,N_10472);
or U11756 (N_11756,N_10395,N_10874);
nor U11757 (N_11757,N_10505,N_10341);
and U11758 (N_11758,N_10017,N_10462);
nor U11759 (N_11759,N_10663,N_10231);
nor U11760 (N_11760,N_10038,N_10175);
or U11761 (N_11761,N_10464,N_10507);
nand U11762 (N_11762,N_10093,N_10316);
nor U11763 (N_11763,N_10308,N_10846);
or U11764 (N_11764,N_10006,N_10234);
nor U11765 (N_11765,N_10520,N_10752);
nor U11766 (N_11766,N_10821,N_10227);
nor U11767 (N_11767,N_10519,N_10183);
xor U11768 (N_11768,N_10338,N_10438);
and U11769 (N_11769,N_10968,N_10632);
xor U11770 (N_11770,N_10495,N_10430);
nand U11771 (N_11771,N_10853,N_10477);
and U11772 (N_11772,N_10412,N_10283);
or U11773 (N_11773,N_10207,N_10613);
or U11774 (N_11774,N_10985,N_10214);
and U11775 (N_11775,N_10186,N_10288);
and U11776 (N_11776,N_10667,N_10689);
or U11777 (N_11777,N_10578,N_10324);
and U11778 (N_11778,N_10095,N_10322);
and U11779 (N_11779,N_10150,N_10239);
nand U11780 (N_11780,N_10439,N_10248);
nor U11781 (N_11781,N_10373,N_10922);
nand U11782 (N_11782,N_10035,N_10991);
and U11783 (N_11783,N_10636,N_10237);
or U11784 (N_11784,N_10351,N_10651);
or U11785 (N_11785,N_10579,N_10824);
nor U11786 (N_11786,N_10508,N_10898);
xor U11787 (N_11787,N_10872,N_10064);
and U11788 (N_11788,N_10675,N_10913);
and U11789 (N_11789,N_10632,N_10998);
nand U11790 (N_11790,N_10629,N_10697);
and U11791 (N_11791,N_10098,N_10707);
nor U11792 (N_11792,N_10726,N_10729);
and U11793 (N_11793,N_10612,N_10373);
xor U11794 (N_11794,N_10647,N_10382);
nor U11795 (N_11795,N_10104,N_10739);
and U11796 (N_11796,N_10325,N_10337);
or U11797 (N_11797,N_10946,N_10641);
xnor U11798 (N_11798,N_10518,N_10311);
nand U11799 (N_11799,N_10184,N_10604);
xnor U11800 (N_11800,N_10369,N_10493);
and U11801 (N_11801,N_10494,N_10008);
nand U11802 (N_11802,N_10872,N_10093);
nand U11803 (N_11803,N_10886,N_10020);
nor U11804 (N_11804,N_10261,N_10960);
and U11805 (N_11805,N_10731,N_10705);
nor U11806 (N_11806,N_10734,N_10850);
and U11807 (N_11807,N_10050,N_10120);
nor U11808 (N_11808,N_10932,N_10831);
nor U11809 (N_11809,N_10139,N_10771);
nand U11810 (N_11810,N_10689,N_10128);
and U11811 (N_11811,N_10023,N_10649);
nand U11812 (N_11812,N_10610,N_10018);
nor U11813 (N_11813,N_10781,N_10694);
nor U11814 (N_11814,N_10074,N_10633);
and U11815 (N_11815,N_10418,N_10442);
xor U11816 (N_11816,N_10121,N_10704);
or U11817 (N_11817,N_10035,N_10567);
xnor U11818 (N_11818,N_10005,N_10211);
nor U11819 (N_11819,N_10565,N_10225);
and U11820 (N_11820,N_10061,N_10667);
or U11821 (N_11821,N_10158,N_10055);
xor U11822 (N_11822,N_10616,N_10294);
xor U11823 (N_11823,N_10642,N_10039);
xnor U11824 (N_11824,N_10581,N_10686);
or U11825 (N_11825,N_10232,N_10989);
nor U11826 (N_11826,N_10201,N_10159);
nand U11827 (N_11827,N_10399,N_10549);
nor U11828 (N_11828,N_10686,N_10142);
xor U11829 (N_11829,N_10425,N_10642);
xor U11830 (N_11830,N_10356,N_10579);
nor U11831 (N_11831,N_10354,N_10730);
and U11832 (N_11832,N_10763,N_10944);
and U11833 (N_11833,N_10286,N_10957);
nand U11834 (N_11834,N_10930,N_10563);
nor U11835 (N_11835,N_10379,N_10866);
nand U11836 (N_11836,N_10914,N_10445);
or U11837 (N_11837,N_10345,N_10887);
xor U11838 (N_11838,N_10050,N_10267);
nor U11839 (N_11839,N_10435,N_10963);
nand U11840 (N_11840,N_10263,N_10577);
nand U11841 (N_11841,N_10167,N_10298);
nor U11842 (N_11842,N_10753,N_10133);
nor U11843 (N_11843,N_10257,N_10997);
xnor U11844 (N_11844,N_10495,N_10587);
or U11845 (N_11845,N_10166,N_10381);
nand U11846 (N_11846,N_10625,N_10151);
nand U11847 (N_11847,N_10969,N_10883);
xnor U11848 (N_11848,N_10941,N_10088);
nand U11849 (N_11849,N_10197,N_10956);
and U11850 (N_11850,N_10207,N_10602);
nand U11851 (N_11851,N_10525,N_10261);
nand U11852 (N_11852,N_10098,N_10629);
or U11853 (N_11853,N_10114,N_10392);
or U11854 (N_11854,N_10551,N_10978);
nor U11855 (N_11855,N_10614,N_10128);
nor U11856 (N_11856,N_10548,N_10961);
nand U11857 (N_11857,N_10760,N_10814);
nor U11858 (N_11858,N_10843,N_10762);
or U11859 (N_11859,N_10834,N_10572);
and U11860 (N_11860,N_10714,N_10134);
and U11861 (N_11861,N_10269,N_10310);
or U11862 (N_11862,N_10486,N_10627);
and U11863 (N_11863,N_10579,N_10251);
nand U11864 (N_11864,N_10223,N_10552);
or U11865 (N_11865,N_10526,N_10165);
or U11866 (N_11866,N_10183,N_10688);
xnor U11867 (N_11867,N_10274,N_10691);
or U11868 (N_11868,N_10059,N_10835);
or U11869 (N_11869,N_10770,N_10576);
or U11870 (N_11870,N_10544,N_10579);
or U11871 (N_11871,N_10947,N_10149);
nor U11872 (N_11872,N_10145,N_10470);
or U11873 (N_11873,N_10738,N_10205);
and U11874 (N_11874,N_10363,N_10000);
nand U11875 (N_11875,N_10051,N_10882);
xor U11876 (N_11876,N_10459,N_10308);
xor U11877 (N_11877,N_10068,N_10903);
or U11878 (N_11878,N_10777,N_10298);
and U11879 (N_11879,N_10830,N_10037);
and U11880 (N_11880,N_10021,N_10268);
or U11881 (N_11881,N_10168,N_10052);
nand U11882 (N_11882,N_10525,N_10859);
xnor U11883 (N_11883,N_10938,N_10926);
xor U11884 (N_11884,N_10344,N_10693);
and U11885 (N_11885,N_10525,N_10884);
and U11886 (N_11886,N_10614,N_10510);
or U11887 (N_11887,N_10427,N_10816);
xnor U11888 (N_11888,N_10982,N_10359);
xnor U11889 (N_11889,N_10590,N_10217);
nor U11890 (N_11890,N_10527,N_10924);
and U11891 (N_11891,N_10460,N_10501);
nor U11892 (N_11892,N_10684,N_10340);
xor U11893 (N_11893,N_10434,N_10227);
or U11894 (N_11894,N_10863,N_10755);
and U11895 (N_11895,N_10285,N_10716);
and U11896 (N_11896,N_10879,N_10831);
nand U11897 (N_11897,N_10014,N_10382);
nand U11898 (N_11898,N_10703,N_10082);
or U11899 (N_11899,N_10542,N_10393);
nor U11900 (N_11900,N_10736,N_10778);
nand U11901 (N_11901,N_10970,N_10666);
nand U11902 (N_11902,N_10116,N_10896);
xor U11903 (N_11903,N_10409,N_10148);
or U11904 (N_11904,N_10244,N_10991);
nor U11905 (N_11905,N_10576,N_10532);
nand U11906 (N_11906,N_10477,N_10114);
and U11907 (N_11907,N_10098,N_10906);
nor U11908 (N_11908,N_10779,N_10751);
and U11909 (N_11909,N_10173,N_10657);
nor U11910 (N_11910,N_10851,N_10195);
nor U11911 (N_11911,N_10747,N_10965);
nand U11912 (N_11912,N_10728,N_10326);
or U11913 (N_11913,N_10427,N_10948);
and U11914 (N_11914,N_10379,N_10567);
nor U11915 (N_11915,N_10021,N_10246);
nand U11916 (N_11916,N_10903,N_10680);
nor U11917 (N_11917,N_10185,N_10017);
nor U11918 (N_11918,N_10694,N_10742);
and U11919 (N_11919,N_10481,N_10992);
and U11920 (N_11920,N_10493,N_10437);
xnor U11921 (N_11921,N_10646,N_10802);
nand U11922 (N_11922,N_10097,N_10408);
or U11923 (N_11923,N_10190,N_10556);
and U11924 (N_11924,N_10132,N_10677);
nand U11925 (N_11925,N_10534,N_10850);
xor U11926 (N_11926,N_10453,N_10512);
or U11927 (N_11927,N_10752,N_10722);
nor U11928 (N_11928,N_10179,N_10488);
and U11929 (N_11929,N_10444,N_10839);
and U11930 (N_11930,N_10135,N_10138);
nor U11931 (N_11931,N_10784,N_10868);
nor U11932 (N_11932,N_10324,N_10665);
xnor U11933 (N_11933,N_10243,N_10234);
and U11934 (N_11934,N_10519,N_10289);
and U11935 (N_11935,N_10308,N_10443);
and U11936 (N_11936,N_10177,N_10054);
and U11937 (N_11937,N_10085,N_10650);
nand U11938 (N_11938,N_10222,N_10684);
and U11939 (N_11939,N_10204,N_10176);
nor U11940 (N_11940,N_10144,N_10686);
xnor U11941 (N_11941,N_10347,N_10696);
and U11942 (N_11942,N_10340,N_10046);
nor U11943 (N_11943,N_10754,N_10059);
nor U11944 (N_11944,N_10857,N_10322);
and U11945 (N_11945,N_10686,N_10990);
or U11946 (N_11946,N_10887,N_10113);
and U11947 (N_11947,N_10190,N_10663);
nor U11948 (N_11948,N_10896,N_10548);
or U11949 (N_11949,N_10570,N_10639);
or U11950 (N_11950,N_10267,N_10840);
xnor U11951 (N_11951,N_10641,N_10444);
nand U11952 (N_11952,N_10898,N_10565);
and U11953 (N_11953,N_10923,N_10435);
or U11954 (N_11954,N_10154,N_10565);
and U11955 (N_11955,N_10140,N_10856);
and U11956 (N_11956,N_10579,N_10785);
nand U11957 (N_11957,N_10068,N_10171);
or U11958 (N_11958,N_10478,N_10886);
xnor U11959 (N_11959,N_10072,N_10910);
or U11960 (N_11960,N_10898,N_10231);
and U11961 (N_11961,N_10581,N_10510);
and U11962 (N_11962,N_10857,N_10984);
or U11963 (N_11963,N_10869,N_10291);
or U11964 (N_11964,N_10735,N_10143);
or U11965 (N_11965,N_10345,N_10989);
or U11966 (N_11966,N_10608,N_10820);
or U11967 (N_11967,N_10556,N_10048);
xor U11968 (N_11968,N_10655,N_10246);
or U11969 (N_11969,N_10641,N_10210);
xnor U11970 (N_11970,N_10205,N_10441);
nand U11971 (N_11971,N_10008,N_10820);
xnor U11972 (N_11972,N_10252,N_10860);
xor U11973 (N_11973,N_10256,N_10599);
and U11974 (N_11974,N_10141,N_10645);
nand U11975 (N_11975,N_10747,N_10120);
nor U11976 (N_11976,N_10212,N_10946);
or U11977 (N_11977,N_10352,N_10706);
and U11978 (N_11978,N_10894,N_10905);
xnor U11979 (N_11979,N_10365,N_10739);
and U11980 (N_11980,N_10880,N_10237);
xor U11981 (N_11981,N_10022,N_10787);
xor U11982 (N_11982,N_10021,N_10929);
nand U11983 (N_11983,N_10217,N_10960);
or U11984 (N_11984,N_10540,N_10004);
or U11985 (N_11985,N_10337,N_10115);
and U11986 (N_11986,N_10425,N_10236);
nor U11987 (N_11987,N_10691,N_10767);
nand U11988 (N_11988,N_10094,N_10950);
xnor U11989 (N_11989,N_10062,N_10244);
nor U11990 (N_11990,N_10861,N_10270);
and U11991 (N_11991,N_10242,N_10214);
or U11992 (N_11992,N_10412,N_10083);
xnor U11993 (N_11993,N_10022,N_10426);
and U11994 (N_11994,N_10757,N_10687);
and U11995 (N_11995,N_10590,N_10580);
nor U11996 (N_11996,N_10127,N_10195);
xnor U11997 (N_11997,N_10150,N_10015);
or U11998 (N_11998,N_10426,N_10563);
or U11999 (N_11999,N_10332,N_10212);
and U12000 (N_12000,N_11520,N_11196);
and U12001 (N_12001,N_11103,N_11840);
and U12002 (N_12002,N_11421,N_11943);
xor U12003 (N_12003,N_11995,N_11937);
or U12004 (N_12004,N_11785,N_11550);
and U12005 (N_12005,N_11330,N_11576);
nor U12006 (N_12006,N_11250,N_11050);
or U12007 (N_12007,N_11644,N_11230);
nand U12008 (N_12008,N_11653,N_11647);
nor U12009 (N_12009,N_11605,N_11185);
and U12010 (N_12010,N_11071,N_11851);
nor U12011 (N_12011,N_11130,N_11542);
xor U12012 (N_12012,N_11583,N_11926);
nand U12013 (N_12013,N_11176,N_11949);
nand U12014 (N_12014,N_11159,N_11489);
xor U12015 (N_12015,N_11763,N_11362);
nand U12016 (N_12016,N_11564,N_11812);
nand U12017 (N_12017,N_11961,N_11596);
nand U12018 (N_12018,N_11641,N_11790);
xnor U12019 (N_12019,N_11157,N_11494);
nand U12020 (N_12020,N_11978,N_11706);
and U12021 (N_12021,N_11984,N_11685);
nand U12022 (N_12022,N_11096,N_11317);
and U12023 (N_12023,N_11166,N_11532);
nor U12024 (N_12024,N_11956,N_11622);
xnor U12025 (N_12025,N_11223,N_11599);
or U12026 (N_12026,N_11424,N_11201);
or U12027 (N_12027,N_11345,N_11575);
and U12028 (N_12028,N_11420,N_11437);
nor U12029 (N_12029,N_11070,N_11303);
and U12030 (N_12030,N_11173,N_11213);
or U12031 (N_12031,N_11615,N_11628);
nand U12032 (N_12032,N_11521,N_11898);
and U12033 (N_12033,N_11434,N_11353);
nor U12034 (N_12034,N_11425,N_11132);
xnor U12035 (N_12035,N_11630,N_11720);
xor U12036 (N_12036,N_11121,N_11052);
xnor U12037 (N_12037,N_11920,N_11650);
nand U12038 (N_12038,N_11057,N_11447);
nand U12039 (N_12039,N_11998,N_11702);
nand U12040 (N_12040,N_11922,N_11453);
xor U12041 (N_12041,N_11301,N_11046);
or U12042 (N_12042,N_11385,N_11939);
or U12043 (N_12043,N_11056,N_11178);
nand U12044 (N_12044,N_11858,N_11661);
nand U12045 (N_12045,N_11125,N_11562);
nand U12046 (N_12046,N_11310,N_11382);
and U12047 (N_12047,N_11439,N_11678);
and U12048 (N_12048,N_11415,N_11264);
and U12049 (N_12049,N_11803,N_11917);
and U12050 (N_12050,N_11624,N_11507);
and U12051 (N_12051,N_11451,N_11901);
xnor U12052 (N_12052,N_11503,N_11681);
or U12053 (N_12053,N_11927,N_11339);
or U12054 (N_12054,N_11783,N_11151);
or U12055 (N_12055,N_11872,N_11934);
nor U12056 (N_12056,N_11545,N_11510);
nor U12057 (N_12057,N_11200,N_11569);
or U12058 (N_12058,N_11587,N_11109);
nor U12059 (N_12059,N_11204,N_11402);
nor U12060 (N_12060,N_11780,N_11667);
or U12061 (N_12061,N_11274,N_11828);
nor U12062 (N_12062,N_11000,N_11391);
nand U12063 (N_12063,N_11859,N_11994);
and U12064 (N_12064,N_11002,N_11277);
or U12065 (N_12065,N_11340,N_11038);
nor U12066 (N_12066,N_11767,N_11919);
and U12067 (N_12067,N_11044,N_11866);
xor U12068 (N_12068,N_11710,N_11383);
xor U12069 (N_12069,N_11006,N_11460);
or U12070 (N_12070,N_11880,N_11065);
xor U12071 (N_12071,N_11062,N_11705);
or U12072 (N_12072,N_11574,N_11017);
nand U12073 (N_12073,N_11184,N_11755);
and U12074 (N_12074,N_11139,N_11895);
nor U12075 (N_12075,N_11222,N_11129);
or U12076 (N_12076,N_11036,N_11386);
nand U12077 (N_12077,N_11498,N_11138);
and U12078 (N_12078,N_11392,N_11633);
and U12079 (N_12079,N_11729,N_11941);
xor U12080 (N_12080,N_11528,N_11850);
nand U12081 (N_12081,N_11808,N_11536);
xnor U12082 (N_12082,N_11761,N_11714);
nor U12083 (N_12083,N_11607,N_11560);
nand U12084 (N_12084,N_11772,N_11098);
nand U12085 (N_12085,N_11465,N_11942);
nor U12086 (N_12086,N_11722,N_11960);
or U12087 (N_12087,N_11068,N_11217);
xor U12088 (N_12088,N_11549,N_11796);
and U12089 (N_12089,N_11619,N_11160);
and U12090 (N_12090,N_11406,N_11401);
nand U12091 (N_12091,N_11302,N_11623);
and U12092 (N_12092,N_11309,N_11945);
nor U12093 (N_12093,N_11189,N_11776);
xnor U12094 (N_12094,N_11271,N_11134);
xnor U12095 (N_12095,N_11110,N_11617);
or U12096 (N_12096,N_11766,N_11579);
or U12097 (N_12097,N_11707,N_11896);
nand U12098 (N_12098,N_11511,N_11290);
nor U12099 (N_12099,N_11873,N_11603);
xor U12100 (N_12100,N_11351,N_11957);
xnor U12101 (N_12101,N_11913,N_11100);
nand U12102 (N_12102,N_11727,N_11304);
nor U12103 (N_12103,N_11212,N_11058);
xor U12104 (N_12104,N_11049,N_11203);
nand U12105 (N_12105,N_11833,N_11344);
or U12106 (N_12106,N_11743,N_11762);
and U12107 (N_12107,N_11053,N_11584);
or U12108 (N_12108,N_11395,N_11933);
or U12109 (N_12109,N_11674,N_11643);
nor U12110 (N_12110,N_11531,N_11343);
nand U12111 (N_12111,N_11249,N_11894);
xor U12112 (N_12112,N_11226,N_11462);
and U12113 (N_12113,N_11903,N_11652);
and U12114 (N_12114,N_11182,N_11556);
or U12115 (N_12115,N_11809,N_11752);
nor U12116 (N_12116,N_11372,N_11951);
and U12117 (N_12117,N_11117,N_11765);
xnor U12118 (N_12118,N_11673,N_11989);
nor U12119 (N_12119,N_11713,N_11580);
or U12120 (N_12120,N_11262,N_11589);
nor U12121 (N_12121,N_11795,N_11443);
xor U12122 (N_12122,N_11384,N_11582);
xnor U12123 (N_12123,N_11375,N_11555);
nand U12124 (N_12124,N_11543,N_11683);
xnor U12125 (N_12125,N_11268,N_11784);
xor U12126 (N_12126,N_11518,N_11063);
nor U12127 (N_12127,N_11320,N_11638);
nand U12128 (N_12128,N_11485,N_11712);
xnor U12129 (N_12129,N_11318,N_11348);
or U12130 (N_12130,N_11064,N_11992);
and U12131 (N_12131,N_11244,N_11448);
and U12132 (N_12132,N_11554,N_11733);
and U12133 (N_12133,N_11608,N_11585);
nor U12134 (N_12134,N_11107,N_11496);
nor U12135 (N_12135,N_11023,N_11430);
or U12136 (N_12136,N_11398,N_11777);
xor U12137 (N_12137,N_11209,N_11037);
or U12138 (N_12138,N_11438,N_11876);
xor U12139 (N_12139,N_11504,N_11466);
or U12140 (N_12140,N_11378,N_11081);
xor U12141 (N_12141,N_11324,N_11971);
or U12142 (N_12142,N_11799,N_11513);
xnor U12143 (N_12143,N_11033,N_11101);
xnor U12144 (N_12144,N_11781,N_11969);
xnor U12145 (N_12145,N_11646,N_11613);
and U12146 (N_12146,N_11088,N_11169);
nand U12147 (N_12147,N_11848,N_11962);
xor U12148 (N_12148,N_11161,N_11745);
nand U12149 (N_12149,N_11404,N_11051);
nor U12150 (N_12150,N_11319,N_11394);
and U12151 (N_12151,N_11573,N_11016);
or U12152 (N_12152,N_11839,N_11306);
and U12153 (N_12153,N_11042,N_11190);
or U12154 (N_12154,N_11538,N_11897);
xor U12155 (N_12155,N_11909,N_11568);
and U12156 (N_12156,N_11136,N_11910);
nand U12157 (N_12157,N_11326,N_11150);
or U12158 (N_12158,N_11860,N_11241);
and U12159 (N_12159,N_11167,N_11061);
nand U12160 (N_12160,N_11486,N_11164);
nand U12161 (N_12161,N_11746,N_11165);
or U12162 (N_12162,N_11516,N_11328);
xor U12163 (N_12163,N_11412,N_11635);
or U12164 (N_12164,N_11233,N_11124);
xor U12165 (N_12165,N_11162,N_11374);
nand U12166 (N_12166,N_11759,N_11311);
xor U12167 (N_12167,N_11907,N_11586);
xor U12168 (N_12168,N_11333,N_11611);
nand U12169 (N_12169,N_11293,N_11551);
and U12170 (N_12170,N_11289,N_11771);
and U12171 (N_12171,N_11476,N_11257);
and U12172 (N_12172,N_11074,N_11719);
nor U12173 (N_12173,N_11208,N_11014);
or U12174 (N_12174,N_11458,N_11915);
and U12175 (N_12175,N_11774,N_11665);
nand U12176 (N_12176,N_11216,N_11120);
or U12177 (N_12177,N_11092,N_11308);
nand U12178 (N_12178,N_11959,N_11626);
nand U12179 (N_12179,N_11400,N_11269);
nor U12180 (N_12180,N_11094,N_11793);
xor U12181 (N_12181,N_11814,N_11990);
xnor U12182 (N_12182,N_11691,N_11155);
xnor U12183 (N_12183,N_11807,N_11664);
nor U12184 (N_12184,N_11001,N_11852);
and U12185 (N_12185,N_11970,N_11679);
or U12186 (N_12186,N_11571,N_11655);
nor U12187 (N_12187,N_11566,N_11887);
nand U12188 (N_12188,N_11688,N_11703);
xnor U12189 (N_12189,N_11905,N_11298);
nor U12190 (N_12190,N_11739,N_11409);
and U12191 (N_12191,N_11530,N_11275);
nand U12192 (N_12192,N_11229,N_11717);
and U12193 (N_12193,N_11742,N_11645);
or U12194 (N_12194,N_11426,N_11354);
nor U12195 (N_12195,N_11168,N_11899);
xor U12196 (N_12196,N_11675,N_11030);
or U12197 (N_12197,N_11794,N_11259);
xor U12198 (N_12198,N_11572,N_11171);
and U12199 (N_12199,N_11371,N_11043);
and U12200 (N_12200,N_11818,N_11299);
xor U12201 (N_12201,N_11238,N_11307);
or U12202 (N_12202,N_11791,N_11716);
nor U12203 (N_12203,N_11844,N_11323);
nor U12204 (N_12204,N_11953,N_11292);
nor U12205 (N_12205,N_11696,N_11735);
nor U12206 (N_12206,N_11728,N_11749);
xor U12207 (N_12207,N_11455,N_11741);
and U12208 (N_12208,N_11916,N_11267);
nand U12209 (N_12209,N_11656,N_11862);
nor U12210 (N_12210,N_11515,N_11258);
nand U12211 (N_12211,N_11379,N_11983);
xnor U12212 (N_12212,N_11699,N_11060);
xor U12213 (N_12213,N_11015,N_11614);
and U12214 (N_12214,N_11272,N_11193);
nand U12215 (N_12215,N_11979,N_11663);
or U12216 (N_12216,N_11886,N_11228);
or U12217 (N_12217,N_11687,N_11867);
xor U12218 (N_12218,N_11529,N_11127);
or U12219 (N_12219,N_11889,N_11751);
nand U12220 (N_12220,N_11593,N_11449);
nor U12221 (N_12221,N_11393,N_11266);
xnor U12222 (N_12222,N_11236,N_11422);
and U12223 (N_12223,N_11283,N_11112);
and U12224 (N_12224,N_11940,N_11747);
and U12225 (N_12225,N_11287,N_11329);
nor U12226 (N_12226,N_11723,N_11879);
nand U12227 (N_12227,N_11158,N_11170);
nand U12228 (N_12228,N_11279,N_11967);
and U12229 (N_12229,N_11836,N_11534);
xnor U12230 (N_12230,N_11789,N_11709);
nand U12231 (N_12231,N_11126,N_11815);
and U12232 (N_12232,N_11715,N_11198);
nand U12233 (N_12233,N_11346,N_11313);
xor U12234 (N_12234,N_11853,N_11616);
or U12235 (N_12235,N_11093,N_11008);
or U12236 (N_12236,N_11801,N_11627);
and U12237 (N_12237,N_11488,N_11788);
and U12238 (N_12238,N_11877,N_11831);
xnor U12239 (N_12239,N_11594,N_11552);
xor U12240 (N_12240,N_11478,N_11718);
or U12241 (N_12241,N_11700,N_11559);
or U12242 (N_12242,N_11740,N_11779);
nor U12243 (N_12243,N_11792,N_11186);
and U12244 (N_12244,N_11314,N_11020);
nor U12245 (N_12245,N_11232,N_11618);
and U12246 (N_12246,N_11407,N_11019);
and U12247 (N_12247,N_11798,N_11822);
nor U12248 (N_12248,N_11141,N_11987);
and U12249 (N_12249,N_11597,N_11454);
or U12250 (N_12250,N_11952,N_11682);
nand U12251 (N_12251,N_11865,N_11570);
or U12252 (N_12252,N_11981,N_11199);
xnor U12253 (N_12253,N_11625,N_11377);
and U12254 (N_12254,N_11535,N_11286);
or U12255 (N_12255,N_11505,N_11900);
xor U12256 (N_12256,N_11502,N_11441);
xnor U12257 (N_12257,N_11756,N_11497);
and U12258 (N_12258,N_11242,N_11546);
nor U12259 (N_12259,N_11077,N_11433);
and U12260 (N_12260,N_11432,N_11929);
nand U12261 (N_12261,N_11370,N_11405);
nand U12262 (N_12262,N_11817,N_11483);
or U12263 (N_12263,N_11890,N_11022);
nand U12264 (N_12264,N_11195,N_11701);
xor U12265 (N_12265,N_11738,N_11211);
nand U12266 (N_12266,N_11857,N_11297);
and U12267 (N_12267,N_11367,N_11854);
xnor U12268 (N_12268,N_11031,N_11659);
nor U12269 (N_12269,N_11474,N_11010);
nor U12270 (N_12270,N_11011,N_11525);
nand U12271 (N_12271,N_11336,N_11111);
nand U12272 (N_12272,N_11035,N_11414);
or U12273 (N_12273,N_11609,N_11446);
nand U12274 (N_12274,N_11565,N_11247);
nand U12275 (N_12275,N_11856,N_11221);
or U12276 (N_12276,N_11855,N_11373);
and U12277 (N_12277,N_11248,N_11380);
xnor U12278 (N_12278,N_11581,N_11331);
xnor U12279 (N_12279,N_11461,N_11684);
nor U12280 (N_12280,N_11428,N_11918);
and U12281 (N_12281,N_11364,N_11731);
nor U12282 (N_12282,N_11018,N_11144);
or U12283 (N_12283,N_11540,N_11089);
nor U12284 (N_12284,N_11143,N_11558);
and U12285 (N_12285,N_11137,N_11032);
nand U12286 (N_12286,N_11177,N_11870);
nand U12287 (N_12287,N_11235,N_11082);
or U12288 (N_12288,N_11084,N_11337);
or U12289 (N_12289,N_11399,N_11519);
xor U12290 (N_12290,N_11726,N_11116);
xor U12291 (N_12291,N_11192,N_11832);
or U12292 (N_12292,N_11194,N_11966);
nor U12293 (N_12293,N_11631,N_11411);
xor U12294 (N_12294,N_11188,N_11285);
nand U12295 (N_12295,N_11086,N_11270);
nand U12296 (N_12296,N_11816,N_11359);
nor U12297 (N_12297,N_11355,N_11369);
xor U12298 (N_12298,N_11163,N_11845);
nand U12299 (N_12299,N_11592,N_11999);
or U12300 (N_12300,N_11930,N_11255);
nand U12301 (N_12301,N_11737,N_11932);
and U12302 (N_12302,N_11245,N_11547);
nand U12303 (N_12303,N_11284,N_11567);
xor U12304 (N_12304,N_11846,N_11725);
nor U12305 (N_12305,N_11768,N_11480);
nor U12306 (N_12306,N_11830,N_11868);
nand U12307 (N_12307,N_11537,N_11207);
nand U12308 (N_12308,N_11914,N_11512);
or U12309 (N_12309,N_11403,N_11459);
xor U12310 (N_12310,N_11252,N_11231);
nand U12311 (N_12311,N_11595,N_11921);
xor U12312 (N_12312,N_11841,N_11179);
xnor U12313 (N_12313,N_11240,N_11327);
and U12314 (N_12314,N_11349,N_11429);
xnor U12315 (N_12315,N_11435,N_11690);
xnor U12316 (N_12316,N_11390,N_11174);
or U12317 (N_12317,N_11588,N_11869);
nor U12318 (N_12318,N_11694,N_11436);
or U12319 (N_12319,N_11076,N_11804);
nand U12320 (N_12320,N_11295,N_11105);
and U12321 (N_12321,N_11396,N_11003);
or U12322 (N_12322,N_11468,N_11153);
nor U12323 (N_12323,N_11823,N_11366);
nand U12324 (N_12324,N_11073,N_11069);
nand U12325 (N_12325,N_11629,N_11358);
xor U12326 (N_12326,N_11689,N_11475);
or U12327 (N_12327,N_11191,N_11368);
xor U12328 (N_12328,N_11491,N_11578);
xnor U12329 (N_12329,N_11102,N_11104);
nor U12330 (N_12330,N_11234,N_11884);
nand U12331 (N_12331,N_11444,N_11256);
and U12332 (N_12332,N_11048,N_11210);
or U12333 (N_12333,N_11753,N_11263);
and U12334 (N_12334,N_11410,N_11864);
or U12335 (N_12335,N_11974,N_11312);
and U12336 (N_12336,N_11183,N_11976);
xor U12337 (N_12337,N_11928,N_11004);
nor U12338 (N_12338,N_11027,N_11591);
nand U12339 (N_12339,N_11007,N_11509);
xor U12340 (N_12340,N_11764,N_11842);
and U12341 (N_12341,N_11938,N_11131);
or U12342 (N_12342,N_11676,N_11265);
and U12343 (N_12343,N_11012,N_11342);
and U12344 (N_12344,N_11600,N_11431);
and U12345 (N_12345,N_11837,N_11985);
nand U12346 (N_12346,N_11332,N_11541);
or U12347 (N_12347,N_11944,N_11782);
xor U12348 (N_12348,N_11135,N_11187);
and U12349 (N_12349,N_11891,N_11055);
nor U12350 (N_12350,N_11500,N_11606);
nand U12351 (N_12351,N_11965,N_11775);
nand U12352 (N_12352,N_11418,N_11246);
nand U12353 (N_12353,N_11632,N_11095);
nor U12354 (N_12354,N_11888,N_11620);
xor U12355 (N_12355,N_11123,N_11072);
xor U12356 (N_12356,N_11175,N_11145);
nor U12357 (N_12357,N_11219,N_11863);
and U12358 (N_12358,N_11300,N_11508);
nor U12359 (N_12359,N_11397,N_11754);
nor U12360 (N_12360,N_11711,N_11322);
or U12361 (N_12361,N_11669,N_11181);
or U12362 (N_12362,N_11469,N_11316);
nand U12363 (N_12363,N_11463,N_11885);
xor U12364 (N_12364,N_11381,N_11610);
nor U12365 (N_12365,N_11612,N_11278);
or U12366 (N_12366,N_11450,N_11834);
xnor U12367 (N_12367,N_11122,N_11553);
nand U12368 (N_12368,N_11954,N_11730);
and U12369 (N_12369,N_11637,N_11251);
or U12370 (N_12370,N_11697,N_11698);
xor U12371 (N_12371,N_11079,N_11254);
nor U12372 (N_12372,N_11524,N_11539);
nor U12373 (N_12373,N_11902,N_11786);
nand U12374 (N_12374,N_11416,N_11097);
and U12375 (N_12375,N_11041,N_11024);
xnor U12376 (N_12376,N_11651,N_11871);
or U12377 (N_12377,N_11215,N_11225);
xor U12378 (N_12378,N_11040,N_11861);
nand U12379 (N_12379,N_11693,N_11334);
xnor U12380 (N_12380,N_11294,N_11677);
xor U12381 (N_12381,N_11442,N_11357);
nor U12382 (N_12382,N_11972,N_11066);
nor U12383 (N_12383,N_11843,N_11973);
nand U12384 (N_12384,N_11800,N_11931);
nand U12385 (N_12385,N_11075,N_11281);
xor U12386 (N_12386,N_11825,N_11660);
xor U12387 (N_12387,N_11090,N_11356);
nor U12388 (N_12388,N_11214,N_11517);
nand U12389 (N_12389,N_11577,N_11769);
and U12390 (N_12390,N_11338,N_11147);
or U12391 (N_12391,N_11108,N_11350);
nor U12392 (N_12392,N_11028,N_11544);
xnor U12393 (N_12393,N_11773,N_11875);
or U12394 (N_12394,N_11993,N_11146);
or U12395 (N_12395,N_11602,N_11522);
nand U12396 (N_12396,N_11039,N_11352);
and U12397 (N_12397,N_11760,N_11601);
nor U12398 (N_12398,N_11946,N_11115);
nor U12399 (N_12399,N_11911,N_11533);
and U12400 (N_12400,N_11963,N_11838);
and U12401 (N_12401,N_11237,N_11315);
and U12402 (N_12402,N_11936,N_11347);
and U12403 (N_12403,N_11413,N_11820);
and U12404 (N_12404,N_11280,N_11388);
nor U12405 (N_12405,N_11452,N_11912);
nor U12406 (N_12406,N_11128,N_11034);
nand U12407 (N_12407,N_11819,N_11205);
or U12408 (N_12408,N_11986,N_11218);
nor U12409 (N_12409,N_11639,N_11479);
nand U12410 (N_12410,N_11363,N_11423);
xnor U12411 (N_12411,N_11149,N_11649);
or U12412 (N_12412,N_11197,N_11239);
or U12413 (N_12413,N_11686,N_11464);
nor U12414 (N_12414,N_11206,N_11964);
or U12415 (N_12415,N_11013,N_11654);
nand U12416 (N_12416,N_11787,N_11490);
or U12417 (N_12417,N_11142,N_11085);
nor U12418 (N_12418,N_11417,N_11335);
or U12419 (N_12419,N_11487,N_11133);
or U12420 (N_12420,N_11757,N_11563);
nor U12421 (N_12421,N_11021,N_11045);
or U12422 (N_12422,N_11982,N_11376);
nand U12423 (N_12423,N_11835,N_11408);
or U12424 (N_12424,N_11980,N_11947);
nand U12425 (N_12425,N_11078,N_11261);
nor U12426 (N_12426,N_11826,N_11672);
xor U12427 (N_12427,N_11878,N_11472);
or U12428 (N_12428,N_11091,N_11227);
nor U12429 (N_12429,N_11827,N_11904);
xor U12430 (N_12430,N_11882,N_11029);
nor U12431 (N_12431,N_11467,N_11924);
or U12432 (N_12432,N_11054,N_11527);
nand U12433 (N_12433,N_11321,N_11389);
nor U12434 (N_12434,N_11724,N_11119);
or U12435 (N_12435,N_11273,N_11906);
or U12436 (N_12436,N_11471,N_11657);
nor U12437 (N_12437,N_11260,N_11810);
xnor U12438 (N_12438,N_11180,N_11477);
xor U12439 (N_12439,N_11708,N_11893);
nor U12440 (N_12440,N_11988,N_11658);
or U12441 (N_12441,N_11883,N_11977);
or U12442 (N_12442,N_11925,N_11670);
xor U12443 (N_12443,N_11276,N_11805);
nor U12444 (N_12444,N_11561,N_11341);
nand U12445 (N_12445,N_11457,N_11470);
nand U12446 (N_12446,N_11958,N_11692);
or U12447 (N_12447,N_11172,N_11634);
nand U12448 (N_12448,N_11590,N_11821);
or U12449 (N_12449,N_11662,N_11671);
and U12450 (N_12450,N_11797,N_11704);
or U12451 (N_12451,N_11695,N_11968);
nand U12452 (N_12452,N_11305,N_11621);
nand U12453 (N_12453,N_11736,N_11948);
and U12454 (N_12454,N_11526,N_11514);
and U12455 (N_12455,N_11080,N_11829);
nand U12456 (N_12456,N_11419,N_11955);
nand U12457 (N_12457,N_11482,N_11824);
or U12458 (N_12458,N_11202,N_11154);
nor U12459 (N_12459,N_11083,N_11440);
or U12460 (N_12460,N_11732,N_11325);
xnor U12461 (N_12461,N_11813,N_11059);
nand U12462 (N_12462,N_11881,N_11365);
xnor U12463 (N_12463,N_11026,N_11758);
or U12464 (N_12464,N_11975,N_11640);
and U12465 (N_12465,N_11288,N_11025);
nor U12466 (N_12466,N_11387,N_11721);
nand U12467 (N_12467,N_11156,N_11636);
nand U12468 (N_12468,N_11047,N_11427);
and U12469 (N_12469,N_11114,N_11243);
and U12470 (N_12470,N_11106,N_11067);
nand U12471 (N_12471,N_11473,N_11806);
xnor U12472 (N_12472,N_11642,N_11481);
nand U12473 (N_12473,N_11009,N_11923);
nand U12474 (N_12474,N_11604,N_11282);
or U12475 (N_12475,N_11557,N_11253);
xor U12476 (N_12476,N_11778,N_11087);
nand U12477 (N_12477,N_11523,N_11291);
or U12478 (N_12478,N_11935,N_11847);
nor U12479 (N_12479,N_11598,N_11680);
or U12480 (N_12480,N_11666,N_11445);
and U12481 (N_12481,N_11148,N_11499);
xnor U12482 (N_12482,N_11744,N_11005);
xor U12483 (N_12483,N_11495,N_11892);
and U12484 (N_12484,N_11748,N_11152);
or U12485 (N_12485,N_11360,N_11849);
or U12486 (N_12486,N_11874,N_11501);
nand U12487 (N_12487,N_11802,N_11492);
xnor U12488 (N_12488,N_11493,N_11734);
xnor U12489 (N_12489,N_11113,N_11668);
and U12490 (N_12490,N_11648,N_11220);
xnor U12491 (N_12491,N_11456,N_11811);
or U12492 (N_12492,N_11361,N_11484);
nand U12493 (N_12493,N_11996,N_11750);
nand U12494 (N_12494,N_11997,N_11991);
and U12495 (N_12495,N_11140,N_11506);
xor U12496 (N_12496,N_11118,N_11296);
nor U12497 (N_12497,N_11770,N_11950);
xnor U12498 (N_12498,N_11099,N_11908);
xnor U12499 (N_12499,N_11548,N_11224);
nand U12500 (N_12500,N_11997,N_11395);
or U12501 (N_12501,N_11874,N_11844);
nor U12502 (N_12502,N_11855,N_11835);
xor U12503 (N_12503,N_11180,N_11985);
xnor U12504 (N_12504,N_11253,N_11602);
or U12505 (N_12505,N_11907,N_11999);
nor U12506 (N_12506,N_11983,N_11691);
nor U12507 (N_12507,N_11801,N_11659);
and U12508 (N_12508,N_11143,N_11468);
and U12509 (N_12509,N_11261,N_11731);
or U12510 (N_12510,N_11680,N_11999);
and U12511 (N_12511,N_11698,N_11380);
and U12512 (N_12512,N_11615,N_11705);
nor U12513 (N_12513,N_11804,N_11422);
nor U12514 (N_12514,N_11744,N_11283);
nor U12515 (N_12515,N_11360,N_11557);
or U12516 (N_12516,N_11274,N_11762);
nand U12517 (N_12517,N_11510,N_11021);
nand U12518 (N_12518,N_11623,N_11427);
nor U12519 (N_12519,N_11936,N_11448);
xnor U12520 (N_12520,N_11500,N_11108);
or U12521 (N_12521,N_11082,N_11215);
nand U12522 (N_12522,N_11975,N_11423);
nand U12523 (N_12523,N_11165,N_11856);
nand U12524 (N_12524,N_11104,N_11020);
nand U12525 (N_12525,N_11432,N_11188);
and U12526 (N_12526,N_11401,N_11913);
nor U12527 (N_12527,N_11794,N_11248);
nor U12528 (N_12528,N_11519,N_11248);
nor U12529 (N_12529,N_11284,N_11073);
nand U12530 (N_12530,N_11949,N_11802);
nor U12531 (N_12531,N_11505,N_11305);
and U12532 (N_12532,N_11058,N_11663);
or U12533 (N_12533,N_11795,N_11878);
nand U12534 (N_12534,N_11938,N_11279);
xnor U12535 (N_12535,N_11411,N_11782);
nand U12536 (N_12536,N_11712,N_11933);
nor U12537 (N_12537,N_11612,N_11299);
nand U12538 (N_12538,N_11089,N_11236);
nand U12539 (N_12539,N_11698,N_11542);
nor U12540 (N_12540,N_11778,N_11643);
nand U12541 (N_12541,N_11552,N_11209);
xor U12542 (N_12542,N_11738,N_11072);
and U12543 (N_12543,N_11806,N_11228);
xor U12544 (N_12544,N_11463,N_11819);
or U12545 (N_12545,N_11692,N_11068);
nand U12546 (N_12546,N_11604,N_11163);
nor U12547 (N_12547,N_11470,N_11841);
nor U12548 (N_12548,N_11940,N_11430);
xor U12549 (N_12549,N_11903,N_11094);
nor U12550 (N_12550,N_11284,N_11752);
xor U12551 (N_12551,N_11861,N_11972);
xnor U12552 (N_12552,N_11897,N_11872);
nor U12553 (N_12553,N_11287,N_11865);
nand U12554 (N_12554,N_11729,N_11761);
nand U12555 (N_12555,N_11373,N_11023);
nor U12556 (N_12556,N_11663,N_11048);
nor U12557 (N_12557,N_11796,N_11108);
or U12558 (N_12558,N_11263,N_11943);
or U12559 (N_12559,N_11117,N_11868);
or U12560 (N_12560,N_11494,N_11501);
or U12561 (N_12561,N_11512,N_11009);
xor U12562 (N_12562,N_11999,N_11346);
nor U12563 (N_12563,N_11196,N_11809);
xnor U12564 (N_12564,N_11666,N_11653);
nor U12565 (N_12565,N_11888,N_11996);
or U12566 (N_12566,N_11318,N_11377);
or U12567 (N_12567,N_11804,N_11041);
or U12568 (N_12568,N_11171,N_11816);
or U12569 (N_12569,N_11629,N_11084);
or U12570 (N_12570,N_11937,N_11266);
xnor U12571 (N_12571,N_11719,N_11797);
or U12572 (N_12572,N_11211,N_11327);
xnor U12573 (N_12573,N_11211,N_11800);
xor U12574 (N_12574,N_11070,N_11987);
nand U12575 (N_12575,N_11591,N_11857);
xor U12576 (N_12576,N_11674,N_11835);
nor U12577 (N_12577,N_11331,N_11252);
nor U12578 (N_12578,N_11270,N_11798);
or U12579 (N_12579,N_11329,N_11123);
or U12580 (N_12580,N_11283,N_11153);
nand U12581 (N_12581,N_11896,N_11868);
nand U12582 (N_12582,N_11965,N_11997);
xor U12583 (N_12583,N_11111,N_11017);
nor U12584 (N_12584,N_11917,N_11646);
xnor U12585 (N_12585,N_11556,N_11412);
or U12586 (N_12586,N_11049,N_11169);
and U12587 (N_12587,N_11762,N_11870);
and U12588 (N_12588,N_11574,N_11026);
nor U12589 (N_12589,N_11565,N_11728);
or U12590 (N_12590,N_11225,N_11313);
nor U12591 (N_12591,N_11226,N_11019);
nor U12592 (N_12592,N_11646,N_11624);
xor U12593 (N_12593,N_11395,N_11441);
xnor U12594 (N_12594,N_11628,N_11805);
or U12595 (N_12595,N_11939,N_11098);
and U12596 (N_12596,N_11389,N_11470);
or U12597 (N_12597,N_11346,N_11573);
nor U12598 (N_12598,N_11101,N_11448);
nand U12599 (N_12599,N_11138,N_11545);
and U12600 (N_12600,N_11125,N_11791);
xor U12601 (N_12601,N_11209,N_11942);
xor U12602 (N_12602,N_11377,N_11520);
or U12603 (N_12603,N_11292,N_11903);
nor U12604 (N_12604,N_11449,N_11890);
and U12605 (N_12605,N_11269,N_11803);
and U12606 (N_12606,N_11058,N_11675);
and U12607 (N_12607,N_11311,N_11729);
and U12608 (N_12608,N_11177,N_11127);
or U12609 (N_12609,N_11140,N_11227);
nand U12610 (N_12610,N_11001,N_11957);
and U12611 (N_12611,N_11640,N_11727);
nor U12612 (N_12612,N_11869,N_11109);
and U12613 (N_12613,N_11946,N_11392);
nor U12614 (N_12614,N_11883,N_11341);
or U12615 (N_12615,N_11654,N_11517);
and U12616 (N_12616,N_11505,N_11590);
nor U12617 (N_12617,N_11844,N_11179);
nor U12618 (N_12618,N_11666,N_11374);
nor U12619 (N_12619,N_11621,N_11339);
or U12620 (N_12620,N_11950,N_11621);
nor U12621 (N_12621,N_11606,N_11507);
xnor U12622 (N_12622,N_11594,N_11982);
and U12623 (N_12623,N_11754,N_11070);
and U12624 (N_12624,N_11648,N_11922);
xor U12625 (N_12625,N_11946,N_11220);
nor U12626 (N_12626,N_11566,N_11298);
or U12627 (N_12627,N_11649,N_11379);
nand U12628 (N_12628,N_11933,N_11730);
xor U12629 (N_12629,N_11965,N_11309);
nor U12630 (N_12630,N_11024,N_11987);
or U12631 (N_12631,N_11615,N_11891);
and U12632 (N_12632,N_11202,N_11625);
nor U12633 (N_12633,N_11102,N_11425);
and U12634 (N_12634,N_11656,N_11741);
or U12635 (N_12635,N_11390,N_11479);
nand U12636 (N_12636,N_11022,N_11381);
xnor U12637 (N_12637,N_11214,N_11396);
nand U12638 (N_12638,N_11628,N_11761);
nor U12639 (N_12639,N_11242,N_11292);
nor U12640 (N_12640,N_11356,N_11233);
and U12641 (N_12641,N_11808,N_11086);
or U12642 (N_12642,N_11817,N_11845);
xnor U12643 (N_12643,N_11752,N_11568);
and U12644 (N_12644,N_11213,N_11638);
nor U12645 (N_12645,N_11705,N_11004);
nor U12646 (N_12646,N_11488,N_11285);
and U12647 (N_12647,N_11678,N_11934);
xnor U12648 (N_12648,N_11888,N_11990);
xnor U12649 (N_12649,N_11318,N_11884);
xnor U12650 (N_12650,N_11077,N_11104);
nor U12651 (N_12651,N_11901,N_11821);
or U12652 (N_12652,N_11348,N_11238);
nor U12653 (N_12653,N_11335,N_11941);
and U12654 (N_12654,N_11069,N_11200);
and U12655 (N_12655,N_11151,N_11034);
nor U12656 (N_12656,N_11175,N_11589);
nand U12657 (N_12657,N_11233,N_11197);
xor U12658 (N_12658,N_11053,N_11863);
nand U12659 (N_12659,N_11035,N_11299);
xnor U12660 (N_12660,N_11313,N_11159);
nor U12661 (N_12661,N_11114,N_11099);
xor U12662 (N_12662,N_11373,N_11277);
xor U12663 (N_12663,N_11612,N_11627);
xor U12664 (N_12664,N_11008,N_11470);
nor U12665 (N_12665,N_11317,N_11517);
xor U12666 (N_12666,N_11039,N_11533);
and U12667 (N_12667,N_11664,N_11157);
nand U12668 (N_12668,N_11537,N_11485);
or U12669 (N_12669,N_11381,N_11704);
or U12670 (N_12670,N_11732,N_11605);
and U12671 (N_12671,N_11161,N_11319);
xor U12672 (N_12672,N_11161,N_11390);
xor U12673 (N_12673,N_11449,N_11355);
and U12674 (N_12674,N_11138,N_11533);
nor U12675 (N_12675,N_11295,N_11656);
nand U12676 (N_12676,N_11869,N_11214);
and U12677 (N_12677,N_11129,N_11058);
or U12678 (N_12678,N_11805,N_11413);
nor U12679 (N_12679,N_11014,N_11454);
or U12680 (N_12680,N_11252,N_11904);
nand U12681 (N_12681,N_11448,N_11289);
nand U12682 (N_12682,N_11723,N_11699);
nor U12683 (N_12683,N_11842,N_11716);
xnor U12684 (N_12684,N_11790,N_11328);
xor U12685 (N_12685,N_11569,N_11533);
nor U12686 (N_12686,N_11897,N_11737);
nand U12687 (N_12687,N_11485,N_11269);
xor U12688 (N_12688,N_11543,N_11281);
xor U12689 (N_12689,N_11552,N_11739);
xor U12690 (N_12690,N_11412,N_11248);
nand U12691 (N_12691,N_11018,N_11201);
nor U12692 (N_12692,N_11415,N_11097);
nand U12693 (N_12693,N_11130,N_11727);
or U12694 (N_12694,N_11644,N_11488);
xor U12695 (N_12695,N_11336,N_11282);
xor U12696 (N_12696,N_11693,N_11083);
nor U12697 (N_12697,N_11380,N_11608);
nand U12698 (N_12698,N_11416,N_11341);
nand U12699 (N_12699,N_11590,N_11056);
nor U12700 (N_12700,N_11728,N_11592);
or U12701 (N_12701,N_11360,N_11706);
and U12702 (N_12702,N_11711,N_11812);
nor U12703 (N_12703,N_11623,N_11584);
nand U12704 (N_12704,N_11857,N_11429);
or U12705 (N_12705,N_11882,N_11989);
and U12706 (N_12706,N_11874,N_11957);
or U12707 (N_12707,N_11855,N_11699);
and U12708 (N_12708,N_11336,N_11067);
and U12709 (N_12709,N_11708,N_11292);
nand U12710 (N_12710,N_11232,N_11403);
nand U12711 (N_12711,N_11602,N_11031);
nand U12712 (N_12712,N_11522,N_11380);
or U12713 (N_12713,N_11602,N_11085);
xnor U12714 (N_12714,N_11176,N_11216);
nand U12715 (N_12715,N_11438,N_11431);
or U12716 (N_12716,N_11516,N_11427);
or U12717 (N_12717,N_11417,N_11466);
or U12718 (N_12718,N_11479,N_11345);
nand U12719 (N_12719,N_11278,N_11614);
and U12720 (N_12720,N_11428,N_11036);
xor U12721 (N_12721,N_11836,N_11321);
nor U12722 (N_12722,N_11302,N_11823);
and U12723 (N_12723,N_11590,N_11449);
or U12724 (N_12724,N_11199,N_11582);
nand U12725 (N_12725,N_11806,N_11513);
xor U12726 (N_12726,N_11927,N_11526);
and U12727 (N_12727,N_11475,N_11850);
and U12728 (N_12728,N_11490,N_11798);
xor U12729 (N_12729,N_11795,N_11628);
xor U12730 (N_12730,N_11231,N_11219);
xnor U12731 (N_12731,N_11325,N_11326);
nand U12732 (N_12732,N_11528,N_11694);
or U12733 (N_12733,N_11417,N_11041);
or U12734 (N_12734,N_11142,N_11070);
xnor U12735 (N_12735,N_11802,N_11868);
and U12736 (N_12736,N_11768,N_11615);
and U12737 (N_12737,N_11543,N_11629);
and U12738 (N_12738,N_11350,N_11200);
or U12739 (N_12739,N_11402,N_11793);
nand U12740 (N_12740,N_11956,N_11034);
and U12741 (N_12741,N_11785,N_11054);
and U12742 (N_12742,N_11647,N_11444);
nor U12743 (N_12743,N_11159,N_11695);
xnor U12744 (N_12744,N_11034,N_11682);
and U12745 (N_12745,N_11902,N_11849);
nor U12746 (N_12746,N_11110,N_11102);
nor U12747 (N_12747,N_11741,N_11154);
nand U12748 (N_12748,N_11446,N_11925);
xnor U12749 (N_12749,N_11408,N_11624);
nor U12750 (N_12750,N_11976,N_11096);
nor U12751 (N_12751,N_11109,N_11511);
nor U12752 (N_12752,N_11018,N_11719);
nor U12753 (N_12753,N_11827,N_11049);
nand U12754 (N_12754,N_11129,N_11115);
nand U12755 (N_12755,N_11660,N_11208);
and U12756 (N_12756,N_11813,N_11812);
nand U12757 (N_12757,N_11060,N_11874);
or U12758 (N_12758,N_11776,N_11456);
or U12759 (N_12759,N_11183,N_11376);
or U12760 (N_12760,N_11772,N_11127);
nand U12761 (N_12761,N_11090,N_11129);
or U12762 (N_12762,N_11292,N_11154);
or U12763 (N_12763,N_11070,N_11174);
and U12764 (N_12764,N_11416,N_11529);
nand U12765 (N_12765,N_11865,N_11707);
nor U12766 (N_12766,N_11227,N_11312);
and U12767 (N_12767,N_11676,N_11027);
nand U12768 (N_12768,N_11818,N_11301);
nand U12769 (N_12769,N_11461,N_11815);
or U12770 (N_12770,N_11917,N_11427);
nand U12771 (N_12771,N_11427,N_11349);
xnor U12772 (N_12772,N_11149,N_11960);
xor U12773 (N_12773,N_11418,N_11235);
nor U12774 (N_12774,N_11408,N_11364);
and U12775 (N_12775,N_11306,N_11960);
or U12776 (N_12776,N_11341,N_11527);
or U12777 (N_12777,N_11396,N_11409);
nor U12778 (N_12778,N_11786,N_11785);
and U12779 (N_12779,N_11813,N_11472);
nor U12780 (N_12780,N_11364,N_11507);
nand U12781 (N_12781,N_11197,N_11542);
or U12782 (N_12782,N_11374,N_11681);
and U12783 (N_12783,N_11736,N_11579);
nor U12784 (N_12784,N_11932,N_11782);
nand U12785 (N_12785,N_11462,N_11993);
and U12786 (N_12786,N_11362,N_11105);
xor U12787 (N_12787,N_11816,N_11167);
nand U12788 (N_12788,N_11045,N_11007);
xnor U12789 (N_12789,N_11631,N_11514);
and U12790 (N_12790,N_11246,N_11350);
nand U12791 (N_12791,N_11720,N_11701);
nand U12792 (N_12792,N_11700,N_11014);
nor U12793 (N_12793,N_11645,N_11269);
and U12794 (N_12794,N_11737,N_11651);
xor U12795 (N_12795,N_11051,N_11036);
nor U12796 (N_12796,N_11096,N_11060);
nor U12797 (N_12797,N_11995,N_11231);
and U12798 (N_12798,N_11568,N_11706);
nor U12799 (N_12799,N_11356,N_11472);
xnor U12800 (N_12800,N_11550,N_11043);
nand U12801 (N_12801,N_11408,N_11010);
or U12802 (N_12802,N_11269,N_11821);
or U12803 (N_12803,N_11485,N_11731);
or U12804 (N_12804,N_11586,N_11638);
or U12805 (N_12805,N_11083,N_11014);
and U12806 (N_12806,N_11000,N_11615);
or U12807 (N_12807,N_11132,N_11060);
and U12808 (N_12808,N_11127,N_11711);
or U12809 (N_12809,N_11441,N_11654);
xor U12810 (N_12810,N_11938,N_11410);
xor U12811 (N_12811,N_11473,N_11081);
or U12812 (N_12812,N_11697,N_11631);
xnor U12813 (N_12813,N_11136,N_11453);
nand U12814 (N_12814,N_11832,N_11689);
nor U12815 (N_12815,N_11037,N_11862);
or U12816 (N_12816,N_11135,N_11592);
xor U12817 (N_12817,N_11210,N_11838);
or U12818 (N_12818,N_11721,N_11777);
nand U12819 (N_12819,N_11880,N_11185);
nor U12820 (N_12820,N_11531,N_11983);
nor U12821 (N_12821,N_11733,N_11395);
nand U12822 (N_12822,N_11248,N_11246);
or U12823 (N_12823,N_11735,N_11123);
or U12824 (N_12824,N_11441,N_11705);
and U12825 (N_12825,N_11502,N_11193);
xnor U12826 (N_12826,N_11117,N_11072);
xnor U12827 (N_12827,N_11424,N_11402);
or U12828 (N_12828,N_11434,N_11595);
xnor U12829 (N_12829,N_11639,N_11087);
and U12830 (N_12830,N_11273,N_11877);
nand U12831 (N_12831,N_11474,N_11051);
nand U12832 (N_12832,N_11241,N_11407);
nor U12833 (N_12833,N_11080,N_11659);
nand U12834 (N_12834,N_11367,N_11520);
nand U12835 (N_12835,N_11067,N_11837);
nor U12836 (N_12836,N_11771,N_11564);
or U12837 (N_12837,N_11368,N_11279);
nor U12838 (N_12838,N_11644,N_11818);
xor U12839 (N_12839,N_11970,N_11250);
nand U12840 (N_12840,N_11551,N_11470);
and U12841 (N_12841,N_11708,N_11139);
nor U12842 (N_12842,N_11563,N_11866);
and U12843 (N_12843,N_11845,N_11557);
or U12844 (N_12844,N_11897,N_11598);
and U12845 (N_12845,N_11306,N_11162);
xor U12846 (N_12846,N_11079,N_11877);
xor U12847 (N_12847,N_11800,N_11090);
nand U12848 (N_12848,N_11866,N_11242);
xor U12849 (N_12849,N_11488,N_11669);
and U12850 (N_12850,N_11435,N_11910);
nor U12851 (N_12851,N_11851,N_11047);
or U12852 (N_12852,N_11737,N_11485);
xnor U12853 (N_12853,N_11119,N_11885);
nand U12854 (N_12854,N_11353,N_11602);
nor U12855 (N_12855,N_11481,N_11764);
nand U12856 (N_12856,N_11802,N_11561);
and U12857 (N_12857,N_11378,N_11738);
nor U12858 (N_12858,N_11741,N_11199);
nand U12859 (N_12859,N_11608,N_11543);
nor U12860 (N_12860,N_11528,N_11253);
nand U12861 (N_12861,N_11505,N_11106);
or U12862 (N_12862,N_11102,N_11628);
and U12863 (N_12863,N_11543,N_11121);
or U12864 (N_12864,N_11945,N_11052);
and U12865 (N_12865,N_11683,N_11239);
and U12866 (N_12866,N_11787,N_11051);
and U12867 (N_12867,N_11383,N_11689);
or U12868 (N_12868,N_11633,N_11172);
xnor U12869 (N_12869,N_11700,N_11967);
nor U12870 (N_12870,N_11381,N_11689);
xnor U12871 (N_12871,N_11482,N_11720);
nand U12872 (N_12872,N_11350,N_11094);
or U12873 (N_12873,N_11455,N_11268);
xor U12874 (N_12874,N_11596,N_11517);
nand U12875 (N_12875,N_11190,N_11549);
nor U12876 (N_12876,N_11809,N_11955);
nor U12877 (N_12877,N_11095,N_11692);
nor U12878 (N_12878,N_11102,N_11446);
and U12879 (N_12879,N_11065,N_11422);
or U12880 (N_12880,N_11682,N_11233);
or U12881 (N_12881,N_11011,N_11980);
nand U12882 (N_12882,N_11424,N_11011);
or U12883 (N_12883,N_11797,N_11382);
nor U12884 (N_12884,N_11756,N_11804);
and U12885 (N_12885,N_11748,N_11639);
nor U12886 (N_12886,N_11359,N_11160);
nand U12887 (N_12887,N_11803,N_11492);
nand U12888 (N_12888,N_11368,N_11223);
nor U12889 (N_12889,N_11497,N_11580);
or U12890 (N_12890,N_11901,N_11486);
or U12891 (N_12891,N_11157,N_11368);
or U12892 (N_12892,N_11258,N_11566);
or U12893 (N_12893,N_11997,N_11844);
xnor U12894 (N_12894,N_11346,N_11338);
nor U12895 (N_12895,N_11939,N_11050);
xnor U12896 (N_12896,N_11462,N_11301);
and U12897 (N_12897,N_11660,N_11032);
nand U12898 (N_12898,N_11134,N_11106);
nand U12899 (N_12899,N_11973,N_11430);
xnor U12900 (N_12900,N_11147,N_11214);
or U12901 (N_12901,N_11369,N_11783);
nor U12902 (N_12902,N_11582,N_11630);
xor U12903 (N_12903,N_11632,N_11809);
nand U12904 (N_12904,N_11795,N_11479);
nor U12905 (N_12905,N_11219,N_11342);
xor U12906 (N_12906,N_11240,N_11264);
and U12907 (N_12907,N_11754,N_11445);
nor U12908 (N_12908,N_11867,N_11104);
xor U12909 (N_12909,N_11687,N_11670);
and U12910 (N_12910,N_11797,N_11537);
or U12911 (N_12911,N_11924,N_11665);
nand U12912 (N_12912,N_11242,N_11692);
nor U12913 (N_12913,N_11940,N_11627);
xnor U12914 (N_12914,N_11490,N_11203);
and U12915 (N_12915,N_11054,N_11007);
and U12916 (N_12916,N_11238,N_11701);
and U12917 (N_12917,N_11806,N_11191);
nand U12918 (N_12918,N_11532,N_11306);
and U12919 (N_12919,N_11675,N_11374);
or U12920 (N_12920,N_11521,N_11687);
nand U12921 (N_12921,N_11866,N_11597);
or U12922 (N_12922,N_11256,N_11447);
xor U12923 (N_12923,N_11759,N_11303);
nor U12924 (N_12924,N_11992,N_11274);
xor U12925 (N_12925,N_11431,N_11921);
and U12926 (N_12926,N_11095,N_11577);
and U12927 (N_12927,N_11560,N_11844);
and U12928 (N_12928,N_11163,N_11449);
nand U12929 (N_12929,N_11532,N_11197);
and U12930 (N_12930,N_11052,N_11130);
and U12931 (N_12931,N_11728,N_11776);
or U12932 (N_12932,N_11846,N_11188);
nor U12933 (N_12933,N_11541,N_11935);
or U12934 (N_12934,N_11178,N_11011);
xnor U12935 (N_12935,N_11786,N_11156);
nor U12936 (N_12936,N_11766,N_11364);
and U12937 (N_12937,N_11181,N_11375);
or U12938 (N_12938,N_11618,N_11425);
and U12939 (N_12939,N_11220,N_11362);
and U12940 (N_12940,N_11976,N_11791);
nand U12941 (N_12941,N_11481,N_11004);
nor U12942 (N_12942,N_11849,N_11424);
xnor U12943 (N_12943,N_11863,N_11275);
or U12944 (N_12944,N_11804,N_11236);
and U12945 (N_12945,N_11450,N_11218);
nand U12946 (N_12946,N_11438,N_11762);
and U12947 (N_12947,N_11405,N_11123);
or U12948 (N_12948,N_11882,N_11302);
or U12949 (N_12949,N_11656,N_11118);
xor U12950 (N_12950,N_11877,N_11771);
xnor U12951 (N_12951,N_11279,N_11009);
nor U12952 (N_12952,N_11770,N_11720);
or U12953 (N_12953,N_11478,N_11601);
xnor U12954 (N_12954,N_11887,N_11291);
xnor U12955 (N_12955,N_11416,N_11418);
nor U12956 (N_12956,N_11579,N_11340);
nand U12957 (N_12957,N_11141,N_11836);
and U12958 (N_12958,N_11932,N_11390);
nor U12959 (N_12959,N_11683,N_11565);
nand U12960 (N_12960,N_11451,N_11263);
xnor U12961 (N_12961,N_11674,N_11465);
nor U12962 (N_12962,N_11977,N_11304);
nor U12963 (N_12963,N_11264,N_11729);
nand U12964 (N_12964,N_11951,N_11619);
nor U12965 (N_12965,N_11790,N_11754);
or U12966 (N_12966,N_11392,N_11847);
nor U12967 (N_12967,N_11733,N_11816);
nand U12968 (N_12968,N_11298,N_11194);
xnor U12969 (N_12969,N_11538,N_11426);
nor U12970 (N_12970,N_11148,N_11412);
and U12971 (N_12971,N_11949,N_11506);
or U12972 (N_12972,N_11730,N_11269);
nand U12973 (N_12973,N_11055,N_11803);
and U12974 (N_12974,N_11074,N_11952);
nand U12975 (N_12975,N_11721,N_11216);
or U12976 (N_12976,N_11865,N_11261);
and U12977 (N_12977,N_11409,N_11806);
nor U12978 (N_12978,N_11819,N_11745);
nand U12979 (N_12979,N_11633,N_11409);
and U12980 (N_12980,N_11425,N_11581);
and U12981 (N_12981,N_11756,N_11817);
nand U12982 (N_12982,N_11193,N_11165);
nand U12983 (N_12983,N_11902,N_11104);
nand U12984 (N_12984,N_11780,N_11525);
xor U12985 (N_12985,N_11974,N_11404);
nor U12986 (N_12986,N_11011,N_11806);
and U12987 (N_12987,N_11941,N_11878);
and U12988 (N_12988,N_11295,N_11437);
nand U12989 (N_12989,N_11192,N_11910);
nand U12990 (N_12990,N_11453,N_11053);
or U12991 (N_12991,N_11301,N_11327);
nand U12992 (N_12992,N_11163,N_11345);
nor U12993 (N_12993,N_11805,N_11581);
xnor U12994 (N_12994,N_11462,N_11688);
and U12995 (N_12995,N_11650,N_11539);
and U12996 (N_12996,N_11588,N_11804);
xor U12997 (N_12997,N_11842,N_11637);
nor U12998 (N_12998,N_11894,N_11938);
xor U12999 (N_12999,N_11736,N_11134);
nor U13000 (N_13000,N_12542,N_12297);
or U13001 (N_13001,N_12829,N_12757);
xor U13002 (N_13002,N_12903,N_12392);
xor U13003 (N_13003,N_12989,N_12747);
and U13004 (N_13004,N_12375,N_12415);
and U13005 (N_13005,N_12028,N_12045);
nor U13006 (N_13006,N_12697,N_12178);
xor U13007 (N_13007,N_12300,N_12058);
or U13008 (N_13008,N_12044,N_12263);
and U13009 (N_13009,N_12991,N_12020);
xor U13010 (N_13010,N_12167,N_12124);
or U13011 (N_13011,N_12533,N_12384);
nand U13012 (N_13012,N_12377,N_12061);
nor U13013 (N_13013,N_12270,N_12064);
nand U13014 (N_13014,N_12987,N_12002);
or U13015 (N_13015,N_12670,N_12496);
nand U13016 (N_13016,N_12210,N_12379);
nand U13017 (N_13017,N_12161,N_12198);
xor U13018 (N_13018,N_12705,N_12333);
and U13019 (N_13019,N_12878,N_12145);
xnor U13020 (N_13020,N_12181,N_12628);
nor U13021 (N_13021,N_12049,N_12784);
xor U13022 (N_13022,N_12823,N_12822);
xor U13023 (N_13023,N_12015,N_12717);
or U13024 (N_13024,N_12732,N_12071);
or U13025 (N_13025,N_12977,N_12998);
or U13026 (N_13026,N_12662,N_12909);
nor U13027 (N_13027,N_12986,N_12069);
or U13028 (N_13028,N_12520,N_12046);
nand U13029 (N_13029,N_12597,N_12952);
and U13030 (N_13030,N_12033,N_12357);
or U13031 (N_13031,N_12828,N_12367);
or U13032 (N_13032,N_12479,N_12984);
nand U13033 (N_13033,N_12087,N_12125);
and U13034 (N_13034,N_12268,N_12723);
and U13035 (N_13035,N_12889,N_12431);
nand U13036 (N_13036,N_12816,N_12738);
nand U13037 (N_13037,N_12113,N_12502);
nand U13038 (N_13038,N_12638,N_12907);
and U13039 (N_13039,N_12218,N_12538);
xor U13040 (N_13040,N_12805,N_12331);
and U13041 (N_13041,N_12912,N_12311);
and U13042 (N_13042,N_12819,N_12872);
xnor U13043 (N_13043,N_12525,N_12604);
or U13044 (N_13044,N_12323,N_12477);
and U13045 (N_13045,N_12294,N_12922);
and U13046 (N_13046,N_12899,N_12447);
xor U13047 (N_13047,N_12933,N_12378);
nor U13048 (N_13048,N_12056,N_12134);
and U13049 (N_13049,N_12778,N_12004);
and U13050 (N_13050,N_12966,N_12097);
xor U13051 (N_13051,N_12650,N_12754);
nor U13052 (N_13052,N_12963,N_12352);
nand U13053 (N_13053,N_12132,N_12715);
xor U13054 (N_13054,N_12651,N_12656);
xor U13055 (N_13055,N_12718,N_12328);
xnor U13056 (N_13056,N_12234,N_12424);
xnor U13057 (N_13057,N_12469,N_12136);
or U13058 (N_13058,N_12141,N_12835);
nor U13059 (N_13059,N_12193,N_12343);
nand U13060 (N_13060,N_12327,N_12126);
xor U13061 (N_13061,N_12402,N_12882);
xnor U13062 (N_13062,N_12517,N_12495);
nand U13063 (N_13063,N_12122,N_12674);
and U13064 (N_13064,N_12555,N_12285);
and U13065 (N_13065,N_12936,N_12873);
nor U13066 (N_13066,N_12528,N_12272);
nor U13067 (N_13067,N_12649,N_12036);
nor U13068 (N_13068,N_12802,N_12950);
nand U13069 (N_13069,N_12480,N_12523);
nand U13070 (N_13070,N_12295,N_12971);
and U13071 (N_13071,N_12475,N_12632);
xor U13072 (N_13072,N_12164,N_12283);
nand U13073 (N_13073,N_12111,N_12332);
xnor U13074 (N_13074,N_12432,N_12789);
xnor U13075 (N_13075,N_12260,N_12478);
nor U13076 (N_13076,N_12485,N_12934);
xnor U13077 (N_13077,N_12782,N_12834);
xor U13078 (N_13078,N_12644,N_12760);
and U13079 (N_13079,N_12448,N_12460);
xor U13080 (N_13080,N_12329,N_12054);
and U13081 (N_13081,N_12494,N_12959);
nand U13082 (N_13082,N_12668,N_12930);
nor U13083 (N_13083,N_12314,N_12844);
and U13084 (N_13084,N_12923,N_12369);
xnor U13085 (N_13085,N_12557,N_12890);
xor U13086 (N_13086,N_12550,N_12146);
and U13087 (N_13087,N_12077,N_12827);
or U13088 (N_13088,N_12277,N_12673);
or U13089 (N_13089,N_12059,N_12669);
nor U13090 (N_13090,N_12356,N_12306);
nand U13091 (N_13091,N_12565,N_12355);
xor U13092 (N_13092,N_12464,N_12364);
nor U13093 (N_13093,N_12007,N_12645);
or U13094 (N_13094,N_12060,N_12012);
or U13095 (N_13095,N_12967,N_12707);
nand U13096 (N_13096,N_12252,N_12716);
nor U13097 (N_13097,N_12762,N_12014);
xor U13098 (N_13098,N_12736,N_12596);
xnor U13099 (N_13099,N_12980,N_12326);
xnor U13100 (N_13100,N_12999,N_12545);
and U13101 (N_13101,N_12220,N_12353);
and U13102 (N_13102,N_12699,N_12454);
xnor U13103 (N_13103,N_12826,N_12261);
nand U13104 (N_13104,N_12595,N_12793);
xor U13105 (N_13105,N_12691,N_12927);
nor U13106 (N_13106,N_12667,N_12773);
nand U13107 (N_13107,N_12990,N_12947);
nor U13108 (N_13108,N_12640,N_12706);
nor U13109 (N_13109,N_12157,N_12886);
nor U13110 (N_13110,N_12450,N_12586);
or U13111 (N_13111,N_12531,N_12063);
nor U13112 (N_13112,N_12606,N_12488);
or U13113 (N_13113,N_12030,N_12983);
nor U13114 (N_13114,N_12229,N_12547);
nand U13115 (N_13115,N_12993,N_12339);
and U13116 (N_13116,N_12133,N_12841);
xnor U13117 (N_13117,N_12901,N_12374);
or U13118 (N_13118,N_12582,N_12455);
nor U13119 (N_13119,N_12150,N_12753);
nand U13120 (N_13120,N_12420,N_12221);
nor U13121 (N_13121,N_12937,N_12387);
nor U13122 (N_13122,N_12072,N_12965);
nand U13123 (N_13123,N_12729,N_12010);
nor U13124 (N_13124,N_12226,N_12245);
and U13125 (N_13125,N_12804,N_12838);
nand U13126 (N_13126,N_12183,N_12724);
or U13127 (N_13127,N_12682,N_12380);
xor U13128 (N_13128,N_12401,N_12344);
and U13129 (N_13129,N_12140,N_12879);
xnor U13130 (N_13130,N_12009,N_12803);
or U13131 (N_13131,N_12155,N_12259);
and U13132 (N_13132,N_12227,N_12516);
nand U13133 (N_13133,N_12439,N_12437);
or U13134 (N_13134,N_12385,N_12438);
or U13135 (N_13135,N_12184,N_12043);
and U13136 (N_13136,N_12591,N_12486);
nand U13137 (N_13137,N_12027,N_12601);
and U13138 (N_13138,N_12771,N_12588);
and U13139 (N_13139,N_12708,N_12700);
xor U13140 (N_13140,N_12679,N_12476);
or U13141 (N_13141,N_12888,N_12530);
nor U13142 (N_13142,N_12880,N_12660);
and U13143 (N_13143,N_12642,N_12928);
nand U13144 (N_13144,N_12951,N_12631);
nand U13145 (N_13145,N_12726,N_12837);
or U13146 (N_13146,N_12511,N_12877);
or U13147 (N_13147,N_12501,N_12042);
nand U13148 (N_13148,N_12085,N_12625);
and U13149 (N_13149,N_12571,N_12047);
nor U13150 (N_13150,N_12116,N_12053);
nor U13151 (N_13151,N_12500,N_12428);
nand U13152 (N_13152,N_12840,N_12080);
nor U13153 (N_13153,N_12713,N_12037);
nand U13154 (N_13154,N_12953,N_12459);
nor U13155 (N_13155,N_12932,N_12281);
xor U13156 (N_13156,N_12924,N_12858);
and U13157 (N_13157,N_12780,N_12659);
nor U13158 (N_13158,N_12792,N_12949);
nand U13159 (N_13159,N_12179,N_12162);
and U13160 (N_13160,N_12925,N_12630);
nor U13161 (N_13161,N_12745,N_12749);
nor U13162 (N_13162,N_12766,N_12246);
nor U13163 (N_13163,N_12103,N_12107);
or U13164 (N_13164,N_12169,N_12529);
nor U13165 (N_13165,N_12605,N_12068);
or U13166 (N_13166,N_12000,N_12764);
nand U13167 (N_13167,N_12076,N_12358);
and U13168 (N_13168,N_12962,N_12251);
or U13169 (N_13169,N_12634,N_12399);
nand U13170 (N_13170,N_12472,N_12710);
nor U13171 (N_13171,N_12284,N_12238);
or U13172 (N_13172,N_12919,N_12563);
or U13173 (N_13173,N_12482,N_12614);
nand U13174 (N_13174,N_12173,N_12958);
nand U13175 (N_13175,N_12973,N_12170);
nand U13176 (N_13176,N_12016,N_12405);
xor U13177 (N_13177,N_12677,N_12808);
and U13178 (N_13178,N_12131,N_12203);
xor U13179 (N_13179,N_12532,N_12964);
nand U13180 (N_13180,N_12845,N_12940);
xnor U13181 (N_13181,N_12629,N_12381);
or U13182 (N_13182,N_12553,N_12807);
xnor U13183 (N_13183,N_12939,N_12201);
xnor U13184 (N_13184,N_12239,N_12893);
nand U13185 (N_13185,N_12487,N_12118);
nand U13186 (N_13186,N_12023,N_12585);
and U13187 (N_13187,N_12204,N_12862);
nor U13188 (N_13188,N_12641,N_12894);
nand U13189 (N_13189,N_12335,N_12470);
nor U13190 (N_13190,N_12457,N_12904);
xor U13191 (N_13191,N_12313,N_12172);
or U13192 (N_13192,N_12598,N_12534);
or U13193 (N_13193,N_12573,N_12154);
and U13194 (N_13194,N_12296,N_12138);
nand U13195 (N_13195,N_12618,N_12086);
and U13196 (N_13196,N_12190,N_12489);
nand U13197 (N_13197,N_12159,N_12094);
or U13198 (N_13198,N_12775,N_12073);
and U13199 (N_13199,N_12446,N_12096);
nor U13200 (N_13200,N_12216,N_12338);
or U13201 (N_13201,N_12915,N_12633);
xor U13202 (N_13202,N_12413,N_12391);
nor U13203 (N_13203,N_12276,N_12404);
and U13204 (N_13204,N_12115,N_12746);
or U13205 (N_13205,N_12365,N_12196);
nor U13206 (N_13206,N_12315,N_12847);
or U13207 (N_13207,N_12900,N_12207);
xor U13208 (N_13208,N_12978,N_12280);
or U13209 (N_13209,N_12084,N_12818);
xnor U13210 (N_13210,N_12689,N_12104);
or U13211 (N_13211,N_12067,N_12288);
and U13212 (N_13212,N_12083,N_12627);
nand U13213 (N_13213,N_12617,N_12175);
and U13214 (N_13214,N_12011,N_12194);
xnor U13215 (N_13215,N_12318,N_12740);
and U13216 (N_13216,N_12386,N_12896);
and U13217 (N_13217,N_12982,N_12995);
xnor U13218 (N_13218,N_12102,N_12619);
xnor U13219 (N_13219,N_12798,N_12916);
and U13220 (N_13220,N_12021,N_12974);
xor U13221 (N_13221,N_12564,N_12636);
and U13222 (N_13222,N_12892,N_12935);
or U13223 (N_13223,N_12735,N_12709);
nand U13224 (N_13224,N_12174,N_12350);
or U13225 (N_13225,N_12442,N_12539);
and U13226 (N_13226,N_12988,N_12088);
nand U13227 (N_13227,N_12739,N_12055);
and U13228 (N_13228,N_12751,N_12763);
and U13229 (N_13229,N_12224,N_12451);
xnor U13230 (N_13230,N_12490,N_12461);
nor U13231 (N_13231,N_12694,N_12695);
and U13232 (N_13232,N_12954,N_12748);
xor U13233 (N_13233,N_12264,N_12149);
or U13234 (N_13234,N_12870,N_12655);
nor U13235 (N_13235,N_12594,N_12209);
and U13236 (N_13236,N_12497,N_12254);
and U13237 (N_13237,N_12981,N_12910);
nor U13238 (N_13238,N_12859,N_12307);
and U13239 (N_13239,N_12456,N_12540);
nor U13240 (N_13240,N_12292,N_12257);
nor U13241 (N_13241,N_12051,N_12733);
xor U13242 (N_13242,N_12544,N_12503);
and U13243 (N_13243,N_12092,N_12883);
nand U13244 (N_13244,N_12473,N_12574);
xnor U13245 (N_13245,N_12678,N_12696);
nand U13246 (N_13246,N_12309,N_12985);
and U13247 (N_13247,N_12906,N_12139);
and U13248 (N_13248,N_12039,N_12558);
and U13249 (N_13249,N_12787,N_12852);
nand U13250 (N_13250,N_12017,N_12824);
nor U13251 (N_13251,N_12767,N_12452);
nor U13252 (N_13252,N_12219,N_12024);
xnor U13253 (N_13253,N_12722,N_12742);
and U13254 (N_13254,N_12171,N_12814);
nand U13255 (N_13255,N_12120,N_12079);
and U13256 (N_13256,N_12110,N_12022);
or U13257 (N_13257,N_12945,N_12199);
and U13258 (N_13258,N_12508,N_12316);
and U13259 (N_13259,N_12383,N_12731);
or U13260 (N_13260,N_12885,N_12177);
xnor U13261 (N_13261,N_12714,N_12869);
and U13262 (N_13262,N_12918,N_12799);
or U13263 (N_13263,N_12917,N_12408);
and U13264 (N_13264,N_12626,N_12683);
xnor U13265 (N_13265,N_12554,N_12266);
and U13266 (N_13266,N_12248,N_12361);
nor U13267 (N_13267,N_12941,N_12692);
and U13268 (N_13268,N_12992,N_12240);
xor U13269 (N_13269,N_12166,N_12944);
nor U13270 (N_13270,N_12290,N_12895);
xor U13271 (N_13271,N_12664,N_12400);
xnor U13272 (N_13272,N_12622,N_12008);
and U13273 (N_13273,N_12688,N_12524);
and U13274 (N_13274,N_12492,N_12427);
or U13275 (N_13275,N_12801,N_12498);
xnor U13276 (N_13276,N_12752,N_12395);
xor U13277 (N_13277,N_12815,N_12693);
and U13278 (N_13278,N_12646,N_12790);
nor U13279 (N_13279,N_12599,N_12567);
nand U13280 (N_13280,N_12881,N_12412);
nor U13281 (N_13281,N_12310,N_12647);
and U13282 (N_13282,N_12756,N_12225);
or U13283 (N_13283,N_12509,N_12794);
nor U13284 (N_13284,N_12189,N_12855);
xnor U13285 (N_13285,N_12863,N_12394);
and U13286 (N_13286,N_12806,N_12652);
and U13287 (N_13287,N_12481,N_12969);
nor U13288 (N_13288,N_12275,N_12279);
nor U13289 (N_13289,N_12127,N_12579);
and U13290 (N_13290,N_12854,N_12610);
nor U13291 (N_13291,N_12330,N_12018);
xnor U13292 (N_13292,N_12360,N_12293);
or U13293 (N_13293,N_12825,N_12301);
or U13294 (N_13294,N_12961,N_12050);
or U13295 (N_13295,N_12351,N_12144);
nand U13296 (N_13296,N_12362,N_12434);
xor U13297 (N_13297,N_12772,N_12968);
nand U13298 (N_13298,N_12876,N_12850);
nor U13299 (N_13299,N_12552,N_12317);
or U13300 (N_13300,N_12129,N_12830);
nor U13301 (N_13301,N_12419,N_12908);
and U13302 (N_13302,N_12615,N_12271);
nand U13303 (N_13303,N_12556,N_12119);
or U13304 (N_13304,N_12425,N_12602);
and U13305 (N_13305,N_12666,N_12026);
nor U13306 (N_13306,N_12108,N_12099);
nand U13307 (N_13307,N_12758,N_12302);
nor U13308 (N_13308,N_12341,N_12730);
nor U13309 (N_13309,N_12551,N_12874);
nor U13310 (N_13310,N_12635,N_12836);
xor U13311 (N_13311,N_12608,N_12440);
or U13312 (N_13312,N_12624,N_12675);
and U13313 (N_13313,N_12593,N_12583);
or U13314 (N_13314,N_12324,N_12491);
and U13315 (N_13315,N_12156,N_12403);
and U13316 (N_13316,N_12676,N_12712);
xnor U13317 (N_13317,N_12643,N_12654);
nand U13318 (N_13318,N_12371,N_12781);
nand U13319 (N_13319,N_12512,N_12005);
nor U13320 (N_13320,N_12397,N_12443);
and U13321 (N_13321,N_12561,N_12422);
xor U13322 (N_13322,N_12833,N_12960);
and U13323 (N_13323,N_12414,N_12421);
xor U13324 (N_13324,N_12319,N_12884);
xnor U13325 (N_13325,N_12543,N_12861);
nand U13326 (N_13326,N_12518,N_12286);
and U13327 (N_13327,N_12527,N_12267);
nand U13328 (N_13328,N_12979,N_12291);
nor U13329 (N_13329,N_12029,N_12349);
and U13330 (N_13330,N_12737,N_12359);
nor U13331 (N_13331,N_12347,N_12727);
xor U13332 (N_13332,N_12074,N_12537);
or U13333 (N_13333,N_12112,N_12920);
xnor U13334 (N_13334,N_12613,N_12938);
or U13335 (N_13335,N_12151,N_12168);
nand U13336 (N_13336,N_12776,N_12957);
and U13337 (N_13337,N_12955,N_12911);
nand U13338 (N_13338,N_12857,N_12719);
nand U13339 (N_13339,N_12897,N_12811);
or U13340 (N_13340,N_12163,N_12759);
and U13341 (N_13341,N_12548,N_12325);
and U13342 (N_13342,N_12831,N_12657);
or U13343 (N_13343,N_12721,N_12546);
xor U13344 (N_13344,N_12100,N_12188);
or U13345 (N_13345,N_12779,N_12137);
xnor U13346 (N_13346,N_12734,N_12621);
nand U13347 (N_13347,N_12505,N_12340);
and U13348 (N_13348,N_12817,N_12230);
nor U13349 (N_13349,N_12744,N_12942);
and U13350 (N_13350,N_12926,N_12215);
nand U13351 (N_13351,N_12943,N_12493);
nor U13352 (N_13352,N_12994,N_12269);
or U13353 (N_13353,N_12462,N_12444);
nand U13354 (N_13354,N_12609,N_12466);
or U13355 (N_13355,N_12703,N_12777);
xnor U13356 (N_13356,N_12453,N_12856);
nand U13357 (N_13357,N_12867,N_12253);
and U13358 (N_13358,N_12101,N_12580);
nand U13359 (N_13359,N_12006,N_12148);
or U13360 (N_13360,N_12914,N_12001);
xnor U13361 (N_13361,N_12449,N_12013);
nand U13362 (N_13362,N_12303,N_12728);
or U13363 (N_13363,N_12346,N_12468);
nand U13364 (N_13364,N_12376,N_12684);
nor U13365 (N_13365,N_12282,N_12681);
nor U13366 (N_13366,N_12791,N_12244);
nor U13367 (N_13367,N_12192,N_12813);
nand U13368 (N_13368,N_12887,N_12458);
nand U13369 (N_13369,N_12577,N_12143);
and U13370 (N_13370,N_12623,N_12312);
and U13371 (N_13371,N_12255,N_12373);
nand U13372 (N_13372,N_12471,N_12334);
xor U13373 (N_13373,N_12406,N_12299);
or U13374 (N_13374,N_12003,N_12465);
or U13375 (N_13375,N_12569,N_12320);
and U13376 (N_13376,N_12091,N_12510);
xor U13377 (N_13377,N_12342,N_12905);
or U13378 (N_13378,N_12584,N_12515);
nor U13379 (N_13379,N_12972,N_12435);
xor U13380 (N_13380,N_12182,N_12363);
xor U13381 (N_13381,N_12337,N_12956);
nand U13382 (N_13382,N_12158,N_12114);
and U13383 (N_13383,N_12687,N_12568);
xnor U13384 (N_13384,N_12783,N_12536);
or U13385 (N_13385,N_12411,N_12235);
or U13386 (N_13386,N_12250,N_12066);
nand U13387 (N_13387,N_12770,N_12637);
or U13388 (N_13388,N_12418,N_12186);
nor U13389 (N_13389,N_12052,N_12081);
or U13390 (N_13390,N_12680,N_12416);
xor U13391 (N_13391,N_12590,N_12843);
or U13392 (N_13392,N_12430,N_12562);
nand U13393 (N_13393,N_12720,N_12875);
xor U13394 (N_13394,N_12663,N_12019);
xnor U13395 (N_13395,N_12535,N_12612);
xor U13396 (N_13396,N_12600,N_12786);
nor U13397 (N_13397,N_12589,N_12390);
xor U13398 (N_13398,N_12274,N_12304);
or U13399 (N_13399,N_12519,N_12389);
nand U13400 (N_13400,N_12587,N_12997);
and U13401 (N_13401,N_12195,N_12851);
nor U13402 (N_13402,N_12109,N_12262);
or U13403 (N_13403,N_12025,N_12152);
and U13404 (N_13404,N_12233,N_12040);
and U13405 (N_13405,N_12768,N_12948);
nor U13406 (N_13406,N_12526,N_12970);
xor U13407 (N_13407,N_12130,N_12785);
nor U13408 (N_13408,N_12153,N_12575);
xor U13409 (N_13409,N_12871,N_12217);
or U13410 (N_13410,N_12581,N_12348);
xnor U13411 (N_13411,N_12034,N_12445);
or U13412 (N_13412,N_12795,N_12812);
xor U13413 (N_13413,N_12241,N_12846);
and U13414 (N_13414,N_12407,N_12228);
nand U13415 (N_13415,N_12370,N_12278);
xor U13416 (N_13416,N_12231,N_12820);
and U13417 (N_13417,N_12147,N_12032);
or U13418 (N_13418,N_12976,N_12160);
xor U13419 (N_13419,N_12265,N_12499);
or U13420 (N_13420,N_12409,N_12522);
or U13421 (N_13421,N_12105,N_12075);
or U13422 (N_13422,N_12410,N_12506);
nor U13423 (N_13423,N_12237,N_12396);
xnor U13424 (N_13424,N_12648,N_12214);
xnor U13425 (N_13425,N_12821,N_12197);
and U13426 (N_13426,N_12603,N_12514);
xnor U13427 (N_13427,N_12504,N_12607);
and U13428 (N_13428,N_12913,N_12572);
and U13429 (N_13429,N_12321,N_12433);
xor U13430 (N_13430,N_12142,N_12866);
xnor U13431 (N_13431,N_12839,N_12661);
nor U13432 (N_13432,N_12298,N_12236);
or U13433 (N_13433,N_12429,N_12180);
nor U13434 (N_13434,N_12665,N_12741);
xnor U13435 (N_13435,N_12135,N_12592);
and U13436 (N_13436,N_12128,N_12672);
xor U13437 (N_13437,N_12576,N_12322);
nor U13438 (N_13438,N_12921,N_12521);
nand U13439 (N_13439,N_12711,N_12243);
nand U13440 (N_13440,N_12273,N_12223);
or U13441 (N_13441,N_12382,N_12653);
nand U13442 (N_13442,N_12256,N_12832);
nand U13443 (N_13443,N_12366,N_12769);
nand U13444 (N_13444,N_12176,N_12702);
xnor U13445 (N_13445,N_12810,N_12078);
nor U13446 (N_13446,N_12975,N_12388);
or U13447 (N_13447,N_12860,N_12743);
or U13448 (N_13448,N_12788,N_12725);
nand U13449 (N_13449,N_12774,N_12089);
and U13450 (N_13450,N_12185,N_12507);
or U13451 (N_13451,N_12368,N_12848);
or U13452 (N_13452,N_12658,N_12698);
nor U13453 (N_13453,N_12853,N_12616);
or U13454 (N_13454,N_12849,N_12242);
xor U13455 (N_13455,N_12200,N_12123);
and U13456 (N_13456,N_12308,N_12797);
and U13457 (N_13457,N_12423,N_12249);
nand U13458 (N_13458,N_12578,N_12426);
or U13459 (N_13459,N_12620,N_12931);
nor U13460 (N_13460,N_12093,N_12765);
or U13461 (N_13461,N_12098,N_12570);
and U13462 (N_13462,N_12121,N_12441);
and U13463 (N_13463,N_12639,N_12398);
nor U13464 (N_13464,N_12187,N_12095);
nand U13465 (N_13465,N_12483,N_12041);
and U13466 (N_13466,N_12842,N_12513);
or U13467 (N_13467,N_12305,N_12070);
or U13468 (N_13468,N_12467,N_12704);
and U13469 (N_13469,N_12484,N_12165);
xnor U13470 (N_13470,N_12474,N_12232);
nand U13471 (N_13471,N_12864,N_12549);
xnor U13472 (N_13472,N_12289,N_12031);
nor U13473 (N_13473,N_12996,N_12809);
xnor U13474 (N_13474,N_12206,N_12761);
nor U13475 (N_13475,N_12048,N_12701);
and U13476 (N_13476,N_12685,N_12417);
nor U13477 (N_13477,N_12566,N_12258);
nor U13478 (N_13478,N_12212,N_12560);
nand U13479 (N_13479,N_12065,N_12208);
nor U13480 (N_13480,N_12062,N_12898);
xnor U13481 (N_13481,N_12463,N_12611);
nand U13482 (N_13482,N_12671,N_12800);
nand U13483 (N_13483,N_12090,N_12436);
or U13484 (N_13484,N_12117,N_12211);
nor U13485 (N_13485,N_12559,N_12082);
xor U13486 (N_13486,N_12750,N_12336);
nand U13487 (N_13487,N_12891,N_12287);
nor U13488 (N_13488,N_12038,N_12372);
and U13489 (N_13489,N_12222,N_12106);
and U13490 (N_13490,N_12902,N_12929);
nor U13491 (N_13491,N_12755,N_12946);
xnor U13492 (N_13492,N_12796,N_12205);
nand U13493 (N_13493,N_12191,N_12686);
and U13494 (N_13494,N_12690,N_12213);
nor U13495 (N_13495,N_12202,N_12035);
nand U13496 (N_13496,N_12868,N_12057);
nor U13497 (N_13497,N_12393,N_12865);
nand U13498 (N_13498,N_12345,N_12541);
and U13499 (N_13499,N_12354,N_12247);
nand U13500 (N_13500,N_12463,N_12747);
nand U13501 (N_13501,N_12245,N_12636);
or U13502 (N_13502,N_12715,N_12316);
nor U13503 (N_13503,N_12946,N_12667);
and U13504 (N_13504,N_12857,N_12741);
or U13505 (N_13505,N_12409,N_12379);
or U13506 (N_13506,N_12039,N_12505);
or U13507 (N_13507,N_12061,N_12135);
or U13508 (N_13508,N_12354,N_12052);
and U13509 (N_13509,N_12750,N_12849);
nor U13510 (N_13510,N_12699,N_12981);
or U13511 (N_13511,N_12934,N_12713);
or U13512 (N_13512,N_12114,N_12227);
or U13513 (N_13513,N_12945,N_12428);
or U13514 (N_13514,N_12408,N_12071);
xnor U13515 (N_13515,N_12154,N_12065);
nand U13516 (N_13516,N_12872,N_12740);
xnor U13517 (N_13517,N_12222,N_12879);
or U13518 (N_13518,N_12143,N_12136);
and U13519 (N_13519,N_12260,N_12445);
xor U13520 (N_13520,N_12920,N_12092);
nand U13521 (N_13521,N_12276,N_12647);
nor U13522 (N_13522,N_12362,N_12353);
xor U13523 (N_13523,N_12957,N_12097);
or U13524 (N_13524,N_12402,N_12679);
nor U13525 (N_13525,N_12716,N_12564);
or U13526 (N_13526,N_12918,N_12575);
nand U13527 (N_13527,N_12087,N_12176);
nand U13528 (N_13528,N_12455,N_12971);
and U13529 (N_13529,N_12462,N_12003);
xor U13530 (N_13530,N_12712,N_12324);
or U13531 (N_13531,N_12913,N_12352);
and U13532 (N_13532,N_12332,N_12393);
or U13533 (N_13533,N_12961,N_12323);
or U13534 (N_13534,N_12346,N_12897);
and U13535 (N_13535,N_12373,N_12937);
nand U13536 (N_13536,N_12401,N_12162);
xor U13537 (N_13537,N_12336,N_12505);
nand U13538 (N_13538,N_12944,N_12249);
nor U13539 (N_13539,N_12219,N_12092);
xor U13540 (N_13540,N_12387,N_12850);
nor U13541 (N_13541,N_12172,N_12995);
nor U13542 (N_13542,N_12665,N_12552);
and U13543 (N_13543,N_12733,N_12594);
xor U13544 (N_13544,N_12136,N_12833);
nand U13545 (N_13545,N_12403,N_12397);
nand U13546 (N_13546,N_12071,N_12672);
xor U13547 (N_13547,N_12196,N_12096);
nor U13548 (N_13548,N_12140,N_12664);
nor U13549 (N_13549,N_12578,N_12118);
and U13550 (N_13550,N_12571,N_12905);
xor U13551 (N_13551,N_12139,N_12106);
or U13552 (N_13552,N_12053,N_12134);
nor U13553 (N_13553,N_12971,N_12814);
and U13554 (N_13554,N_12249,N_12456);
or U13555 (N_13555,N_12858,N_12897);
nor U13556 (N_13556,N_12512,N_12306);
nand U13557 (N_13557,N_12764,N_12363);
or U13558 (N_13558,N_12914,N_12071);
xor U13559 (N_13559,N_12225,N_12137);
nor U13560 (N_13560,N_12707,N_12462);
nor U13561 (N_13561,N_12144,N_12054);
and U13562 (N_13562,N_12838,N_12380);
or U13563 (N_13563,N_12355,N_12181);
or U13564 (N_13564,N_12357,N_12276);
xnor U13565 (N_13565,N_12631,N_12896);
xor U13566 (N_13566,N_12213,N_12684);
nand U13567 (N_13567,N_12123,N_12386);
nor U13568 (N_13568,N_12295,N_12707);
xnor U13569 (N_13569,N_12093,N_12797);
nor U13570 (N_13570,N_12490,N_12886);
nor U13571 (N_13571,N_12751,N_12351);
xnor U13572 (N_13572,N_12558,N_12669);
nand U13573 (N_13573,N_12630,N_12339);
or U13574 (N_13574,N_12630,N_12841);
xor U13575 (N_13575,N_12791,N_12794);
and U13576 (N_13576,N_12463,N_12977);
and U13577 (N_13577,N_12034,N_12177);
and U13578 (N_13578,N_12074,N_12767);
or U13579 (N_13579,N_12034,N_12409);
or U13580 (N_13580,N_12427,N_12668);
or U13581 (N_13581,N_12521,N_12540);
and U13582 (N_13582,N_12937,N_12057);
nand U13583 (N_13583,N_12302,N_12548);
nand U13584 (N_13584,N_12081,N_12203);
or U13585 (N_13585,N_12608,N_12362);
and U13586 (N_13586,N_12288,N_12565);
nor U13587 (N_13587,N_12311,N_12613);
xnor U13588 (N_13588,N_12676,N_12091);
nand U13589 (N_13589,N_12355,N_12804);
xnor U13590 (N_13590,N_12015,N_12269);
nand U13591 (N_13591,N_12981,N_12410);
or U13592 (N_13592,N_12668,N_12821);
and U13593 (N_13593,N_12363,N_12807);
nor U13594 (N_13594,N_12597,N_12642);
or U13595 (N_13595,N_12933,N_12471);
or U13596 (N_13596,N_12721,N_12932);
xnor U13597 (N_13597,N_12007,N_12384);
and U13598 (N_13598,N_12664,N_12766);
nor U13599 (N_13599,N_12357,N_12121);
nor U13600 (N_13600,N_12967,N_12277);
xnor U13601 (N_13601,N_12160,N_12503);
and U13602 (N_13602,N_12310,N_12255);
nand U13603 (N_13603,N_12137,N_12845);
nand U13604 (N_13604,N_12714,N_12293);
or U13605 (N_13605,N_12275,N_12431);
or U13606 (N_13606,N_12321,N_12334);
and U13607 (N_13607,N_12995,N_12675);
or U13608 (N_13608,N_12845,N_12193);
or U13609 (N_13609,N_12696,N_12375);
nand U13610 (N_13610,N_12055,N_12566);
xor U13611 (N_13611,N_12973,N_12924);
xnor U13612 (N_13612,N_12723,N_12356);
xor U13613 (N_13613,N_12033,N_12896);
nand U13614 (N_13614,N_12145,N_12164);
or U13615 (N_13615,N_12499,N_12657);
xnor U13616 (N_13616,N_12573,N_12685);
nor U13617 (N_13617,N_12936,N_12495);
nor U13618 (N_13618,N_12541,N_12899);
and U13619 (N_13619,N_12694,N_12387);
nor U13620 (N_13620,N_12691,N_12511);
or U13621 (N_13621,N_12203,N_12059);
or U13622 (N_13622,N_12536,N_12873);
nor U13623 (N_13623,N_12596,N_12125);
and U13624 (N_13624,N_12238,N_12392);
nand U13625 (N_13625,N_12630,N_12247);
nor U13626 (N_13626,N_12177,N_12281);
nor U13627 (N_13627,N_12245,N_12193);
xnor U13628 (N_13628,N_12540,N_12696);
or U13629 (N_13629,N_12400,N_12960);
nand U13630 (N_13630,N_12783,N_12278);
or U13631 (N_13631,N_12169,N_12094);
nand U13632 (N_13632,N_12833,N_12231);
nor U13633 (N_13633,N_12791,N_12138);
nand U13634 (N_13634,N_12085,N_12437);
nand U13635 (N_13635,N_12255,N_12401);
xnor U13636 (N_13636,N_12917,N_12150);
nand U13637 (N_13637,N_12753,N_12123);
or U13638 (N_13638,N_12535,N_12116);
and U13639 (N_13639,N_12328,N_12614);
and U13640 (N_13640,N_12431,N_12876);
nor U13641 (N_13641,N_12043,N_12961);
or U13642 (N_13642,N_12730,N_12589);
or U13643 (N_13643,N_12836,N_12169);
nand U13644 (N_13644,N_12552,N_12319);
nand U13645 (N_13645,N_12558,N_12814);
xnor U13646 (N_13646,N_12163,N_12867);
or U13647 (N_13647,N_12605,N_12780);
or U13648 (N_13648,N_12890,N_12780);
xnor U13649 (N_13649,N_12450,N_12534);
and U13650 (N_13650,N_12342,N_12501);
xor U13651 (N_13651,N_12773,N_12420);
or U13652 (N_13652,N_12636,N_12689);
xnor U13653 (N_13653,N_12036,N_12659);
or U13654 (N_13654,N_12791,N_12964);
nor U13655 (N_13655,N_12596,N_12715);
or U13656 (N_13656,N_12706,N_12165);
nand U13657 (N_13657,N_12732,N_12859);
nand U13658 (N_13658,N_12576,N_12299);
xnor U13659 (N_13659,N_12818,N_12814);
xor U13660 (N_13660,N_12443,N_12951);
nor U13661 (N_13661,N_12789,N_12680);
xor U13662 (N_13662,N_12301,N_12927);
nand U13663 (N_13663,N_12947,N_12794);
nand U13664 (N_13664,N_12111,N_12287);
and U13665 (N_13665,N_12526,N_12283);
and U13666 (N_13666,N_12054,N_12830);
and U13667 (N_13667,N_12593,N_12213);
and U13668 (N_13668,N_12305,N_12580);
and U13669 (N_13669,N_12816,N_12600);
xnor U13670 (N_13670,N_12323,N_12660);
and U13671 (N_13671,N_12011,N_12569);
and U13672 (N_13672,N_12093,N_12376);
or U13673 (N_13673,N_12131,N_12048);
nor U13674 (N_13674,N_12721,N_12925);
and U13675 (N_13675,N_12356,N_12429);
and U13676 (N_13676,N_12188,N_12507);
nand U13677 (N_13677,N_12386,N_12221);
nand U13678 (N_13678,N_12262,N_12937);
xor U13679 (N_13679,N_12837,N_12083);
nand U13680 (N_13680,N_12693,N_12804);
xor U13681 (N_13681,N_12150,N_12732);
or U13682 (N_13682,N_12376,N_12327);
nand U13683 (N_13683,N_12132,N_12502);
nor U13684 (N_13684,N_12550,N_12430);
and U13685 (N_13685,N_12973,N_12030);
nor U13686 (N_13686,N_12329,N_12142);
and U13687 (N_13687,N_12456,N_12316);
nand U13688 (N_13688,N_12624,N_12808);
or U13689 (N_13689,N_12454,N_12466);
nor U13690 (N_13690,N_12974,N_12725);
nand U13691 (N_13691,N_12404,N_12311);
and U13692 (N_13692,N_12481,N_12639);
or U13693 (N_13693,N_12133,N_12783);
or U13694 (N_13694,N_12327,N_12366);
or U13695 (N_13695,N_12514,N_12246);
and U13696 (N_13696,N_12243,N_12365);
nor U13697 (N_13697,N_12707,N_12499);
and U13698 (N_13698,N_12478,N_12416);
nor U13699 (N_13699,N_12131,N_12416);
and U13700 (N_13700,N_12180,N_12106);
and U13701 (N_13701,N_12100,N_12592);
xnor U13702 (N_13702,N_12135,N_12861);
nor U13703 (N_13703,N_12726,N_12361);
xor U13704 (N_13704,N_12133,N_12486);
nor U13705 (N_13705,N_12940,N_12973);
and U13706 (N_13706,N_12016,N_12187);
nor U13707 (N_13707,N_12428,N_12338);
nor U13708 (N_13708,N_12393,N_12158);
and U13709 (N_13709,N_12964,N_12263);
xor U13710 (N_13710,N_12534,N_12932);
and U13711 (N_13711,N_12417,N_12376);
nor U13712 (N_13712,N_12900,N_12984);
nand U13713 (N_13713,N_12969,N_12359);
or U13714 (N_13714,N_12169,N_12894);
nand U13715 (N_13715,N_12222,N_12863);
nor U13716 (N_13716,N_12581,N_12381);
or U13717 (N_13717,N_12638,N_12494);
and U13718 (N_13718,N_12793,N_12556);
or U13719 (N_13719,N_12009,N_12750);
and U13720 (N_13720,N_12178,N_12382);
nand U13721 (N_13721,N_12142,N_12659);
nand U13722 (N_13722,N_12777,N_12074);
nor U13723 (N_13723,N_12739,N_12605);
and U13724 (N_13724,N_12687,N_12086);
xnor U13725 (N_13725,N_12658,N_12887);
nand U13726 (N_13726,N_12585,N_12162);
or U13727 (N_13727,N_12380,N_12684);
nand U13728 (N_13728,N_12232,N_12258);
and U13729 (N_13729,N_12500,N_12557);
nor U13730 (N_13730,N_12127,N_12996);
or U13731 (N_13731,N_12833,N_12534);
nand U13732 (N_13732,N_12199,N_12543);
and U13733 (N_13733,N_12386,N_12659);
or U13734 (N_13734,N_12537,N_12640);
nor U13735 (N_13735,N_12361,N_12039);
and U13736 (N_13736,N_12492,N_12825);
and U13737 (N_13737,N_12881,N_12379);
xnor U13738 (N_13738,N_12782,N_12090);
xor U13739 (N_13739,N_12778,N_12882);
and U13740 (N_13740,N_12949,N_12519);
or U13741 (N_13741,N_12338,N_12471);
and U13742 (N_13742,N_12075,N_12989);
nand U13743 (N_13743,N_12566,N_12703);
nor U13744 (N_13744,N_12404,N_12649);
and U13745 (N_13745,N_12395,N_12011);
xor U13746 (N_13746,N_12739,N_12951);
xor U13747 (N_13747,N_12221,N_12260);
and U13748 (N_13748,N_12763,N_12521);
xor U13749 (N_13749,N_12527,N_12136);
xor U13750 (N_13750,N_12010,N_12691);
and U13751 (N_13751,N_12641,N_12420);
or U13752 (N_13752,N_12280,N_12818);
nand U13753 (N_13753,N_12617,N_12647);
nand U13754 (N_13754,N_12416,N_12047);
nor U13755 (N_13755,N_12633,N_12980);
nand U13756 (N_13756,N_12605,N_12853);
nand U13757 (N_13757,N_12281,N_12274);
xor U13758 (N_13758,N_12342,N_12968);
and U13759 (N_13759,N_12326,N_12758);
nor U13760 (N_13760,N_12066,N_12302);
nor U13761 (N_13761,N_12301,N_12355);
or U13762 (N_13762,N_12981,N_12718);
and U13763 (N_13763,N_12958,N_12883);
and U13764 (N_13764,N_12522,N_12285);
or U13765 (N_13765,N_12955,N_12223);
xnor U13766 (N_13766,N_12181,N_12208);
or U13767 (N_13767,N_12450,N_12147);
and U13768 (N_13768,N_12267,N_12526);
nor U13769 (N_13769,N_12554,N_12940);
and U13770 (N_13770,N_12656,N_12596);
xnor U13771 (N_13771,N_12580,N_12016);
or U13772 (N_13772,N_12777,N_12648);
nand U13773 (N_13773,N_12429,N_12980);
xor U13774 (N_13774,N_12653,N_12500);
nand U13775 (N_13775,N_12326,N_12316);
nand U13776 (N_13776,N_12930,N_12538);
and U13777 (N_13777,N_12927,N_12480);
nor U13778 (N_13778,N_12206,N_12381);
nand U13779 (N_13779,N_12151,N_12331);
nand U13780 (N_13780,N_12898,N_12428);
nor U13781 (N_13781,N_12255,N_12092);
or U13782 (N_13782,N_12197,N_12605);
nand U13783 (N_13783,N_12371,N_12971);
xnor U13784 (N_13784,N_12745,N_12357);
nand U13785 (N_13785,N_12567,N_12712);
xnor U13786 (N_13786,N_12617,N_12109);
nand U13787 (N_13787,N_12846,N_12901);
nand U13788 (N_13788,N_12979,N_12834);
xor U13789 (N_13789,N_12844,N_12698);
nor U13790 (N_13790,N_12351,N_12505);
nand U13791 (N_13791,N_12138,N_12487);
nor U13792 (N_13792,N_12661,N_12208);
xor U13793 (N_13793,N_12623,N_12439);
nand U13794 (N_13794,N_12751,N_12842);
nand U13795 (N_13795,N_12947,N_12291);
or U13796 (N_13796,N_12423,N_12345);
and U13797 (N_13797,N_12674,N_12340);
nor U13798 (N_13798,N_12912,N_12328);
nor U13799 (N_13799,N_12333,N_12755);
xor U13800 (N_13800,N_12006,N_12328);
or U13801 (N_13801,N_12290,N_12227);
and U13802 (N_13802,N_12002,N_12991);
nand U13803 (N_13803,N_12050,N_12901);
nand U13804 (N_13804,N_12308,N_12211);
nand U13805 (N_13805,N_12673,N_12185);
nand U13806 (N_13806,N_12143,N_12513);
nand U13807 (N_13807,N_12012,N_12970);
and U13808 (N_13808,N_12245,N_12433);
nand U13809 (N_13809,N_12990,N_12858);
and U13810 (N_13810,N_12943,N_12853);
xor U13811 (N_13811,N_12269,N_12303);
and U13812 (N_13812,N_12538,N_12096);
and U13813 (N_13813,N_12136,N_12067);
and U13814 (N_13814,N_12480,N_12984);
nand U13815 (N_13815,N_12961,N_12731);
nor U13816 (N_13816,N_12362,N_12551);
xor U13817 (N_13817,N_12599,N_12419);
nand U13818 (N_13818,N_12752,N_12365);
nor U13819 (N_13819,N_12874,N_12244);
or U13820 (N_13820,N_12161,N_12685);
xnor U13821 (N_13821,N_12956,N_12464);
nand U13822 (N_13822,N_12437,N_12308);
xnor U13823 (N_13823,N_12320,N_12146);
nand U13824 (N_13824,N_12421,N_12649);
xnor U13825 (N_13825,N_12010,N_12630);
xnor U13826 (N_13826,N_12976,N_12079);
or U13827 (N_13827,N_12908,N_12663);
nand U13828 (N_13828,N_12234,N_12370);
and U13829 (N_13829,N_12849,N_12745);
nand U13830 (N_13830,N_12975,N_12211);
nand U13831 (N_13831,N_12932,N_12636);
nand U13832 (N_13832,N_12317,N_12691);
xnor U13833 (N_13833,N_12941,N_12861);
nor U13834 (N_13834,N_12933,N_12805);
xnor U13835 (N_13835,N_12133,N_12614);
xor U13836 (N_13836,N_12168,N_12066);
xor U13837 (N_13837,N_12092,N_12733);
xor U13838 (N_13838,N_12689,N_12407);
nor U13839 (N_13839,N_12307,N_12388);
xor U13840 (N_13840,N_12687,N_12278);
xnor U13841 (N_13841,N_12824,N_12799);
and U13842 (N_13842,N_12373,N_12083);
xnor U13843 (N_13843,N_12927,N_12232);
nand U13844 (N_13844,N_12191,N_12937);
nand U13845 (N_13845,N_12572,N_12218);
nor U13846 (N_13846,N_12920,N_12412);
and U13847 (N_13847,N_12377,N_12593);
and U13848 (N_13848,N_12340,N_12605);
nor U13849 (N_13849,N_12854,N_12753);
or U13850 (N_13850,N_12333,N_12768);
nor U13851 (N_13851,N_12348,N_12607);
xnor U13852 (N_13852,N_12094,N_12091);
xnor U13853 (N_13853,N_12083,N_12385);
or U13854 (N_13854,N_12765,N_12191);
or U13855 (N_13855,N_12980,N_12761);
nor U13856 (N_13856,N_12389,N_12441);
xnor U13857 (N_13857,N_12808,N_12671);
and U13858 (N_13858,N_12347,N_12748);
nor U13859 (N_13859,N_12782,N_12152);
and U13860 (N_13860,N_12965,N_12535);
xor U13861 (N_13861,N_12277,N_12144);
or U13862 (N_13862,N_12743,N_12531);
nand U13863 (N_13863,N_12271,N_12668);
nor U13864 (N_13864,N_12230,N_12758);
nand U13865 (N_13865,N_12417,N_12644);
or U13866 (N_13866,N_12153,N_12157);
nand U13867 (N_13867,N_12762,N_12195);
xor U13868 (N_13868,N_12946,N_12125);
xor U13869 (N_13869,N_12574,N_12504);
nor U13870 (N_13870,N_12686,N_12946);
and U13871 (N_13871,N_12436,N_12409);
nor U13872 (N_13872,N_12505,N_12738);
xor U13873 (N_13873,N_12229,N_12536);
xor U13874 (N_13874,N_12497,N_12993);
xor U13875 (N_13875,N_12300,N_12368);
nor U13876 (N_13876,N_12179,N_12123);
nand U13877 (N_13877,N_12449,N_12576);
xnor U13878 (N_13878,N_12176,N_12528);
and U13879 (N_13879,N_12332,N_12035);
or U13880 (N_13880,N_12442,N_12544);
and U13881 (N_13881,N_12450,N_12442);
nor U13882 (N_13882,N_12710,N_12604);
and U13883 (N_13883,N_12655,N_12387);
nand U13884 (N_13884,N_12112,N_12092);
xnor U13885 (N_13885,N_12444,N_12088);
xnor U13886 (N_13886,N_12734,N_12619);
and U13887 (N_13887,N_12290,N_12313);
or U13888 (N_13888,N_12331,N_12731);
xor U13889 (N_13889,N_12741,N_12656);
or U13890 (N_13890,N_12284,N_12721);
nor U13891 (N_13891,N_12037,N_12232);
nand U13892 (N_13892,N_12634,N_12357);
nor U13893 (N_13893,N_12547,N_12760);
xnor U13894 (N_13894,N_12673,N_12870);
or U13895 (N_13895,N_12689,N_12511);
xor U13896 (N_13896,N_12819,N_12444);
and U13897 (N_13897,N_12701,N_12107);
xnor U13898 (N_13898,N_12061,N_12758);
or U13899 (N_13899,N_12696,N_12310);
and U13900 (N_13900,N_12606,N_12845);
and U13901 (N_13901,N_12269,N_12102);
or U13902 (N_13902,N_12071,N_12872);
nand U13903 (N_13903,N_12794,N_12732);
and U13904 (N_13904,N_12765,N_12315);
nand U13905 (N_13905,N_12139,N_12233);
or U13906 (N_13906,N_12011,N_12100);
and U13907 (N_13907,N_12006,N_12628);
xor U13908 (N_13908,N_12420,N_12594);
and U13909 (N_13909,N_12233,N_12729);
nand U13910 (N_13910,N_12135,N_12129);
nor U13911 (N_13911,N_12062,N_12336);
nor U13912 (N_13912,N_12315,N_12175);
xor U13913 (N_13913,N_12610,N_12768);
nor U13914 (N_13914,N_12328,N_12945);
nand U13915 (N_13915,N_12367,N_12559);
nand U13916 (N_13916,N_12714,N_12228);
or U13917 (N_13917,N_12115,N_12185);
and U13918 (N_13918,N_12272,N_12709);
xnor U13919 (N_13919,N_12867,N_12943);
nand U13920 (N_13920,N_12971,N_12924);
nor U13921 (N_13921,N_12143,N_12989);
nand U13922 (N_13922,N_12068,N_12420);
nor U13923 (N_13923,N_12749,N_12282);
xor U13924 (N_13924,N_12374,N_12124);
nand U13925 (N_13925,N_12548,N_12480);
and U13926 (N_13926,N_12525,N_12167);
xnor U13927 (N_13927,N_12142,N_12978);
xnor U13928 (N_13928,N_12922,N_12835);
xor U13929 (N_13929,N_12995,N_12289);
nand U13930 (N_13930,N_12192,N_12304);
and U13931 (N_13931,N_12496,N_12669);
and U13932 (N_13932,N_12439,N_12756);
or U13933 (N_13933,N_12216,N_12745);
nor U13934 (N_13934,N_12480,N_12350);
and U13935 (N_13935,N_12797,N_12376);
xor U13936 (N_13936,N_12918,N_12354);
xor U13937 (N_13937,N_12493,N_12039);
nand U13938 (N_13938,N_12446,N_12003);
or U13939 (N_13939,N_12610,N_12892);
nor U13940 (N_13940,N_12260,N_12684);
nand U13941 (N_13941,N_12148,N_12851);
or U13942 (N_13942,N_12865,N_12611);
xnor U13943 (N_13943,N_12881,N_12597);
nor U13944 (N_13944,N_12076,N_12426);
xnor U13945 (N_13945,N_12360,N_12539);
nor U13946 (N_13946,N_12871,N_12453);
xor U13947 (N_13947,N_12601,N_12015);
xnor U13948 (N_13948,N_12435,N_12893);
nor U13949 (N_13949,N_12726,N_12523);
nor U13950 (N_13950,N_12330,N_12422);
nand U13951 (N_13951,N_12960,N_12353);
xor U13952 (N_13952,N_12612,N_12058);
and U13953 (N_13953,N_12792,N_12636);
nor U13954 (N_13954,N_12071,N_12156);
nor U13955 (N_13955,N_12658,N_12001);
nor U13956 (N_13956,N_12956,N_12232);
xor U13957 (N_13957,N_12046,N_12282);
nand U13958 (N_13958,N_12645,N_12008);
or U13959 (N_13959,N_12511,N_12699);
nor U13960 (N_13960,N_12022,N_12134);
nor U13961 (N_13961,N_12594,N_12977);
xnor U13962 (N_13962,N_12533,N_12195);
and U13963 (N_13963,N_12093,N_12543);
or U13964 (N_13964,N_12251,N_12862);
nand U13965 (N_13965,N_12757,N_12578);
or U13966 (N_13966,N_12531,N_12236);
xnor U13967 (N_13967,N_12699,N_12363);
xnor U13968 (N_13968,N_12427,N_12442);
nor U13969 (N_13969,N_12294,N_12160);
nand U13970 (N_13970,N_12962,N_12420);
and U13971 (N_13971,N_12075,N_12484);
nand U13972 (N_13972,N_12380,N_12468);
and U13973 (N_13973,N_12753,N_12452);
nor U13974 (N_13974,N_12803,N_12858);
nor U13975 (N_13975,N_12713,N_12940);
nand U13976 (N_13976,N_12308,N_12745);
nand U13977 (N_13977,N_12438,N_12149);
and U13978 (N_13978,N_12407,N_12851);
and U13979 (N_13979,N_12436,N_12170);
xnor U13980 (N_13980,N_12850,N_12397);
and U13981 (N_13981,N_12935,N_12660);
and U13982 (N_13982,N_12501,N_12068);
nor U13983 (N_13983,N_12829,N_12520);
xor U13984 (N_13984,N_12928,N_12673);
or U13985 (N_13985,N_12998,N_12193);
xor U13986 (N_13986,N_12411,N_12874);
and U13987 (N_13987,N_12053,N_12216);
and U13988 (N_13988,N_12395,N_12052);
xor U13989 (N_13989,N_12540,N_12949);
nand U13990 (N_13990,N_12238,N_12224);
and U13991 (N_13991,N_12527,N_12550);
or U13992 (N_13992,N_12602,N_12467);
or U13993 (N_13993,N_12344,N_12466);
nor U13994 (N_13994,N_12137,N_12042);
and U13995 (N_13995,N_12638,N_12354);
nor U13996 (N_13996,N_12806,N_12139);
and U13997 (N_13997,N_12669,N_12715);
or U13998 (N_13998,N_12079,N_12333);
or U13999 (N_13999,N_12140,N_12219);
nor U14000 (N_14000,N_13398,N_13653);
nor U14001 (N_14001,N_13149,N_13699);
xor U14002 (N_14002,N_13172,N_13162);
xnor U14003 (N_14003,N_13374,N_13052);
xnor U14004 (N_14004,N_13008,N_13990);
and U14005 (N_14005,N_13808,N_13764);
and U14006 (N_14006,N_13747,N_13570);
and U14007 (N_14007,N_13914,N_13640);
and U14008 (N_14008,N_13622,N_13606);
xnor U14009 (N_14009,N_13238,N_13658);
nor U14010 (N_14010,N_13341,N_13303);
nor U14011 (N_14011,N_13415,N_13116);
nor U14012 (N_14012,N_13582,N_13426);
nand U14013 (N_14013,N_13020,N_13531);
xor U14014 (N_14014,N_13359,N_13174);
nor U14015 (N_14015,N_13815,N_13437);
xor U14016 (N_14016,N_13140,N_13476);
xor U14017 (N_14017,N_13504,N_13920);
xor U14018 (N_14018,N_13707,N_13631);
nand U14019 (N_14019,N_13790,N_13089);
xnor U14020 (N_14020,N_13480,N_13642);
nor U14021 (N_14021,N_13235,N_13186);
or U14022 (N_14022,N_13798,N_13313);
nand U14023 (N_14023,N_13510,N_13938);
nor U14024 (N_14024,N_13922,N_13716);
or U14025 (N_14025,N_13961,N_13445);
or U14026 (N_14026,N_13527,N_13381);
and U14027 (N_14027,N_13100,N_13943);
xor U14028 (N_14028,N_13626,N_13109);
nor U14029 (N_14029,N_13175,N_13344);
or U14030 (N_14030,N_13421,N_13461);
xor U14031 (N_14031,N_13268,N_13214);
xor U14032 (N_14032,N_13442,N_13971);
nor U14033 (N_14033,N_13255,N_13645);
nand U14034 (N_14034,N_13927,N_13820);
and U14035 (N_14035,N_13728,N_13240);
and U14036 (N_14036,N_13368,N_13743);
or U14037 (N_14037,N_13017,N_13698);
and U14038 (N_14038,N_13842,N_13173);
nand U14039 (N_14039,N_13039,N_13505);
or U14040 (N_14040,N_13540,N_13541);
and U14041 (N_14041,N_13915,N_13835);
and U14042 (N_14042,N_13388,N_13691);
nand U14043 (N_14043,N_13278,N_13515);
xnor U14044 (N_14044,N_13661,N_13521);
nor U14045 (N_14045,N_13804,N_13280);
or U14046 (N_14046,N_13126,N_13809);
or U14047 (N_14047,N_13573,N_13945);
and U14048 (N_14048,N_13205,N_13551);
nand U14049 (N_14049,N_13482,N_13674);
or U14050 (N_14050,N_13550,N_13111);
and U14051 (N_14051,N_13057,N_13935);
or U14052 (N_14052,N_13704,N_13206);
nand U14053 (N_14053,N_13178,N_13928);
and U14054 (N_14054,N_13256,N_13384);
or U14055 (N_14055,N_13377,N_13748);
and U14056 (N_14056,N_13035,N_13107);
or U14057 (N_14057,N_13428,N_13431);
nand U14058 (N_14058,N_13625,N_13117);
nor U14059 (N_14059,N_13060,N_13718);
and U14060 (N_14060,N_13731,N_13309);
nor U14061 (N_14061,N_13609,N_13357);
and U14062 (N_14062,N_13131,N_13106);
nand U14063 (N_14063,N_13023,N_13318);
nor U14064 (N_14064,N_13055,N_13182);
nand U14065 (N_14065,N_13019,N_13319);
nand U14066 (N_14066,N_13221,N_13564);
xnor U14067 (N_14067,N_13746,N_13877);
xor U14068 (N_14068,N_13477,N_13752);
and U14069 (N_14069,N_13132,N_13618);
and U14070 (N_14070,N_13483,N_13392);
nand U14071 (N_14071,N_13233,N_13115);
nor U14072 (N_14072,N_13033,N_13993);
and U14073 (N_14073,N_13336,N_13678);
and U14074 (N_14074,N_13497,N_13941);
and U14075 (N_14075,N_13837,N_13843);
or U14076 (N_14076,N_13955,N_13644);
nor U14077 (N_14077,N_13378,N_13904);
and U14078 (N_14078,N_13185,N_13158);
nand U14079 (N_14079,N_13857,N_13859);
xor U14080 (N_14080,N_13129,N_13879);
nand U14081 (N_14081,N_13119,N_13204);
and U14082 (N_14082,N_13416,N_13036);
xnor U14083 (N_14083,N_13267,N_13293);
and U14084 (N_14084,N_13247,N_13623);
nand U14085 (N_14085,N_13688,N_13676);
nand U14086 (N_14086,N_13213,N_13352);
or U14087 (N_14087,N_13466,N_13296);
or U14088 (N_14088,N_13127,N_13545);
and U14089 (N_14089,N_13321,N_13519);
xor U14090 (N_14090,N_13340,N_13702);
nand U14091 (N_14091,N_13639,N_13565);
and U14092 (N_14092,N_13844,N_13074);
nor U14093 (N_14093,N_13011,N_13712);
nor U14094 (N_14094,N_13390,N_13272);
nor U14095 (N_14095,N_13153,N_13435);
nor U14096 (N_14096,N_13291,N_13059);
nor U14097 (N_14097,N_13067,N_13758);
and U14098 (N_14098,N_13710,N_13138);
and U14099 (N_14099,N_13867,N_13113);
nor U14100 (N_14100,N_13382,N_13741);
nor U14101 (N_14101,N_13725,N_13327);
xor U14102 (N_14102,N_13995,N_13749);
xor U14103 (N_14103,N_13056,N_13845);
nor U14104 (N_14104,N_13950,N_13686);
and U14105 (N_14105,N_13054,N_13283);
and U14106 (N_14106,N_13148,N_13443);
nand U14107 (N_14107,N_13836,N_13763);
and U14108 (N_14108,N_13043,N_13222);
xor U14109 (N_14109,N_13219,N_13974);
nand U14110 (N_14110,N_13456,N_13422);
xor U14111 (N_14111,N_13157,N_13875);
and U14112 (N_14112,N_13306,N_13114);
and U14113 (N_14113,N_13916,N_13734);
and U14114 (N_14114,N_13290,N_13241);
or U14115 (N_14115,N_13643,N_13769);
nor U14116 (N_14116,N_13629,N_13690);
and U14117 (N_14117,N_13951,N_13264);
or U14118 (N_14118,N_13579,N_13137);
and U14119 (N_14119,N_13890,N_13617);
nor U14120 (N_14120,N_13458,N_13553);
nand U14121 (N_14121,N_13199,N_13635);
xnor U14122 (N_14122,N_13896,N_13365);
nand U14123 (N_14123,N_13464,N_13776);
nand U14124 (N_14124,N_13998,N_13533);
nor U14125 (N_14125,N_13713,N_13438);
nand U14126 (N_14126,N_13536,N_13874);
and U14127 (N_14127,N_13670,N_13898);
nand U14128 (N_14128,N_13795,N_13886);
xor U14129 (N_14129,N_13633,N_13791);
nor U14130 (N_14130,N_13288,N_13072);
nand U14131 (N_14131,N_13616,N_13701);
or U14132 (N_14132,N_13355,N_13555);
xnor U14133 (N_14133,N_13093,N_13248);
or U14134 (N_14134,N_13893,N_13848);
nand U14135 (N_14135,N_13604,N_13169);
nand U14136 (N_14136,N_13332,N_13677);
xor U14137 (N_14137,N_13239,N_13963);
xor U14138 (N_14138,N_13964,N_13261);
and U14139 (N_14139,N_13451,N_13312);
nor U14140 (N_14140,N_13673,N_13145);
xnor U14141 (N_14141,N_13962,N_13449);
xor U14142 (N_14142,N_13002,N_13038);
xnor U14143 (N_14143,N_13793,N_13194);
or U14144 (N_14144,N_13782,N_13584);
nand U14145 (N_14145,N_13663,N_13460);
nand U14146 (N_14146,N_13311,N_13349);
and U14147 (N_14147,N_13393,N_13130);
nand U14148 (N_14148,N_13574,N_13929);
xnor U14149 (N_14149,N_13491,N_13825);
or U14150 (N_14150,N_13755,N_13598);
nor U14151 (N_14151,N_13887,N_13164);
nor U14152 (N_14152,N_13554,N_13258);
xnor U14153 (N_14153,N_13528,N_13170);
nor U14154 (N_14154,N_13833,N_13975);
nor U14155 (N_14155,N_13537,N_13823);
nor U14156 (N_14156,N_13197,N_13930);
xnor U14157 (N_14157,N_13076,N_13988);
or U14158 (N_14158,N_13097,N_13168);
and U14159 (N_14159,N_13919,N_13361);
or U14160 (N_14160,N_13607,N_13738);
xnor U14161 (N_14161,N_13784,N_13511);
or U14162 (N_14162,N_13888,N_13362);
and U14163 (N_14163,N_13750,N_13289);
xor U14164 (N_14164,N_13696,N_13918);
nand U14165 (N_14165,N_13910,N_13517);
xnor U14166 (N_14166,N_13274,N_13212);
and U14167 (N_14167,N_13736,N_13839);
and U14168 (N_14168,N_13789,N_13908);
nand U14169 (N_14169,N_13367,N_13356);
nor U14170 (N_14170,N_13439,N_13489);
nor U14171 (N_14171,N_13577,N_13905);
or U14172 (N_14172,N_13754,N_13939);
nor U14173 (N_14173,N_13369,N_13473);
xnor U14174 (N_14174,N_13447,N_13231);
nand U14175 (N_14175,N_13925,N_13891);
and U14176 (N_14176,N_13029,N_13408);
or U14177 (N_14177,N_13123,N_13147);
nand U14178 (N_14178,N_13246,N_13207);
and U14179 (N_14179,N_13648,N_13657);
nand U14180 (N_14180,N_13529,N_13134);
or U14181 (N_14181,N_13650,N_13487);
xor U14182 (N_14182,N_13014,N_13018);
nand U14183 (N_14183,N_13665,N_13819);
and U14184 (N_14184,N_13612,N_13351);
nor U14185 (N_14185,N_13952,N_13826);
xor U14186 (N_14186,N_13649,N_13371);
or U14187 (N_14187,N_13889,N_13066);
or U14188 (N_14188,N_13335,N_13088);
or U14189 (N_14189,N_13675,N_13615);
nand U14190 (N_14190,N_13781,N_13596);
nand U14191 (N_14191,N_13403,N_13853);
xor U14192 (N_14192,N_13987,N_13370);
nand U14193 (N_14193,N_13244,N_13227);
and U14194 (N_14194,N_13711,N_13389);
nand U14195 (N_14195,N_13811,N_13454);
and U14196 (N_14196,N_13779,N_13721);
nor U14197 (N_14197,N_13202,N_13404);
xor U14198 (N_14198,N_13933,N_13253);
or U14199 (N_14199,N_13757,N_13346);
nor U14200 (N_14200,N_13772,N_13042);
nand U14201 (N_14201,N_13180,N_13501);
and U14202 (N_14202,N_13237,N_13986);
xor U14203 (N_14203,N_13210,N_13250);
or U14204 (N_14204,N_13307,N_13632);
and U14205 (N_14205,N_13103,N_13006);
xor U14206 (N_14206,N_13603,N_13948);
xor U14207 (N_14207,N_13785,N_13331);
xor U14208 (N_14208,N_13139,N_13523);
and U14209 (N_14209,N_13997,N_13401);
xnor U14210 (N_14210,N_13957,N_13440);
nand U14211 (N_14211,N_13176,N_13801);
xnor U14212 (N_14212,N_13308,N_13259);
or U14213 (N_14213,N_13330,N_13216);
and U14214 (N_14214,N_13496,N_13756);
nand U14215 (N_14215,N_13960,N_13478);
xor U14216 (N_14216,N_13128,N_13071);
or U14217 (N_14217,N_13864,N_13709);
and U14218 (N_14218,N_13298,N_13156);
or U14219 (N_14219,N_13223,N_13587);
nor U14220 (N_14220,N_13166,N_13695);
xor U14221 (N_14221,N_13446,N_13485);
nor U14222 (N_14222,N_13965,N_13683);
xor U14223 (N_14223,N_13979,N_13028);
xor U14224 (N_14224,N_13234,N_13061);
xor U14225 (N_14225,N_13708,N_13856);
nand U14226 (N_14226,N_13050,N_13942);
xor U14227 (N_14227,N_13144,N_13585);
xor U14228 (N_14228,N_13479,N_13009);
and U14229 (N_14229,N_13868,N_13581);
or U14230 (N_14230,N_13735,N_13552);
or U14231 (N_14231,N_13342,N_13567);
xnor U14232 (N_14232,N_13124,N_13405);
nor U14233 (N_14233,N_13003,N_13046);
and U14234 (N_14234,N_13242,N_13507);
xnor U14235 (N_14235,N_13705,N_13099);
or U14236 (N_14236,N_13034,N_13871);
xnor U14237 (N_14237,N_13096,N_13339);
nand U14238 (N_14238,N_13771,N_13027);
nor U14239 (N_14239,N_13885,N_13159);
xor U14240 (N_14240,N_13851,N_13984);
or U14241 (N_14241,N_13761,N_13410);
nor U14242 (N_14242,N_13154,N_13522);
nand U14243 (N_14243,N_13467,N_13681);
nand U14244 (N_14244,N_13614,N_13337);
nand U14245 (N_14245,N_13282,N_13829);
or U14246 (N_14246,N_13266,N_13729);
or U14247 (N_14247,N_13098,N_13778);
and U14248 (N_14248,N_13917,N_13816);
or U14249 (N_14249,N_13849,N_13899);
and U14250 (N_14250,N_13338,N_13160);
nand U14251 (N_14251,N_13733,N_13142);
or U14252 (N_14252,N_13465,N_13292);
xor U14253 (N_14253,N_13193,N_13973);
nor U14254 (N_14254,N_13576,N_13559);
xor U14255 (N_14255,N_13506,N_13353);
nor U14256 (N_14256,N_13902,N_13909);
and U14257 (N_14257,N_13730,N_13400);
nand U14258 (N_14258,N_13693,N_13599);
nand U14259 (N_14259,N_13469,N_13641);
or U14260 (N_14260,N_13095,N_13051);
or U14261 (N_14261,N_13862,N_13016);
nand U14262 (N_14262,N_13135,N_13189);
xor U14263 (N_14263,N_13386,N_13269);
xnor U14264 (N_14264,N_13004,N_13832);
xnor U14265 (N_14265,N_13834,N_13668);
and U14266 (N_14266,N_13672,N_13287);
or U14267 (N_14267,N_13907,N_13830);
xnor U14268 (N_14268,N_13740,N_13083);
nor U14269 (N_14269,N_13230,N_13627);
nand U14270 (N_14270,N_13817,N_13660);
nand U14271 (N_14271,N_13094,N_13595);
nor U14272 (N_14272,N_13860,N_13276);
and U14273 (N_14273,N_13068,N_13812);
and U14274 (N_14274,N_13538,N_13444);
or U14275 (N_14275,N_13429,N_13406);
xor U14276 (N_14276,N_13620,N_13275);
and U14277 (N_14277,N_13947,N_13989);
nor U14278 (N_14278,N_13759,N_13053);
xnor U14279 (N_14279,N_13912,N_13310);
and U14280 (N_14280,N_13802,N_13383);
nand U14281 (N_14281,N_13179,N_13122);
or U14282 (N_14282,N_13396,N_13294);
xnor U14283 (N_14283,N_13608,N_13766);
nand U14284 (N_14284,N_13080,N_13031);
nand U14285 (N_14285,N_13846,N_13201);
nand U14286 (N_14286,N_13807,N_13827);
xnor U14287 (N_14287,N_13262,N_13171);
nor U14288 (N_14288,N_13831,N_13092);
nor U14289 (N_14289,N_13884,N_13305);
or U14290 (N_14290,N_13525,N_13358);
xnor U14291 (N_14291,N_13613,N_13569);
xnor U14292 (N_14292,N_13502,N_13744);
and U14293 (N_14293,N_13873,N_13316);
or U14294 (N_14294,N_13881,N_13363);
or U14295 (N_14295,N_13105,N_13121);
nor U14296 (N_14296,N_13425,N_13077);
xnor U14297 (N_14297,N_13513,N_13315);
xor U14298 (N_14298,N_13897,N_13423);
nand U14299 (N_14299,N_13968,N_13911);
nand U14300 (N_14300,N_13064,N_13300);
and U14301 (N_14301,N_13548,N_13719);
and U14302 (N_14302,N_13659,N_13045);
and U14303 (N_14303,N_13638,N_13463);
xor U14304 (N_14304,N_13783,N_13254);
xnor U14305 (N_14305,N_13796,N_13767);
and U14306 (N_14306,N_13325,N_13328);
or U14307 (N_14307,N_13838,N_13697);
and U14308 (N_14308,N_13903,N_13803);
xor U14309 (N_14309,N_13547,N_13568);
and U14310 (N_14310,N_13391,N_13112);
nand U14311 (N_14311,N_13012,N_13544);
or U14312 (N_14312,N_13414,N_13081);
and U14313 (N_14313,N_13208,N_13788);
xnor U14314 (N_14314,N_13087,N_13813);
nand U14315 (N_14315,N_13015,N_13263);
nand U14316 (N_14316,N_13739,N_13110);
nor U14317 (N_14317,N_13196,N_13379);
nor U14318 (N_14318,N_13430,N_13026);
and U14319 (N_14319,N_13492,N_13590);
xnor U14320 (N_14320,N_13571,N_13800);
nor U14321 (N_14321,N_13184,N_13854);
xnor U14322 (N_14322,N_13656,N_13503);
or U14323 (N_14323,N_13366,N_13666);
nor U14324 (N_14324,N_13586,N_13575);
nand U14325 (N_14325,N_13322,N_13556);
nand U14326 (N_14326,N_13058,N_13892);
nor U14327 (N_14327,N_13768,N_13152);
xnor U14328 (N_14328,N_13524,N_13580);
nor U14329 (N_14329,N_13286,N_13500);
and U14330 (N_14330,N_13628,N_13498);
and U14331 (N_14331,N_13424,N_13700);
and U14332 (N_14332,N_13224,N_13745);
nand U14333 (N_14333,N_13413,N_13013);
nand U14334 (N_14334,N_13490,N_13946);
nand U14335 (N_14335,N_13218,N_13163);
or U14336 (N_14336,N_13514,N_13084);
and U14337 (N_14337,N_13985,N_13679);
and U14338 (N_14338,N_13495,N_13277);
nand U14339 (N_14339,N_13714,N_13876);
or U14340 (N_14340,N_13407,N_13777);
xnor U14341 (N_14341,N_13090,N_13921);
and U14342 (N_14342,N_13726,N_13376);
nand U14343 (N_14343,N_13079,N_13694);
and U14344 (N_14344,N_13970,N_13509);
xnor U14345 (N_14345,N_13822,N_13217);
nand U14346 (N_14346,N_13932,N_13484);
and U14347 (N_14347,N_13775,N_13592);
or U14348 (N_14348,N_13563,N_13474);
nand U14349 (N_14349,N_13448,N_13865);
nor U14350 (N_14350,N_13047,N_13324);
xnor U14351 (N_14351,N_13048,N_13343);
nor U14352 (N_14352,N_13901,N_13872);
nor U14353 (N_14353,N_13078,N_13380);
nand U14354 (N_14354,N_13462,N_13601);
and U14355 (N_14355,N_13387,N_13652);
nor U14356 (N_14356,N_13317,N_13198);
nand U14357 (N_14357,N_13419,N_13323);
and U14358 (N_14358,N_13770,N_13546);
xor U14359 (N_14359,N_13302,N_13953);
and U14360 (N_14360,N_13200,N_13432);
xnor U14361 (N_14361,N_13395,N_13345);
nand U14362 (N_14362,N_13040,N_13488);
nand U14363 (N_14363,N_13285,N_13228);
nand U14364 (N_14364,N_13284,N_13441);
or U14365 (N_14365,N_13146,N_13773);
xor U14366 (N_14366,N_13797,N_13118);
nand U14367 (N_14367,N_13411,N_13455);
and U14368 (N_14368,N_13279,N_13883);
xnor U14369 (N_14369,N_13150,N_13976);
nand U14370 (N_14370,N_13102,N_13805);
and U14371 (N_14371,N_13229,N_13958);
xor U14372 (N_14372,N_13999,N_13591);
xnor U14373 (N_14373,N_13966,N_13457);
nor U14374 (N_14374,N_13468,N_13314);
xnor U14375 (N_14375,N_13453,N_13372);
and U14376 (N_14376,N_13774,N_13913);
nand U14377 (N_14377,N_13792,N_13022);
xnor U14378 (N_14378,N_13646,N_13923);
nor U14379 (N_14379,N_13543,N_13824);
and U14380 (N_14380,N_13732,N_13954);
xor U14381 (N_14381,N_13526,N_13669);
and U14382 (N_14382,N_13481,N_13737);
nand U14383 (N_14383,N_13265,N_13720);
xnor U14384 (N_14384,N_13924,N_13433);
xnor U14385 (N_14385,N_13000,N_13715);
nor U14386 (N_14386,N_13252,N_13086);
or U14387 (N_14387,N_13073,N_13271);
or U14388 (N_14388,N_13760,N_13530);
xor U14389 (N_14389,N_13520,N_13840);
xor U14390 (N_14390,N_13155,N_13977);
and U14391 (N_14391,N_13062,N_13956);
nor U14392 (N_14392,N_13814,N_13049);
nor U14393 (N_14393,N_13188,N_13295);
nand U14394 (N_14394,N_13594,N_13177);
xor U14395 (N_14395,N_13895,N_13597);
and U14396 (N_14396,N_13181,N_13753);
nand U14397 (N_14397,N_13991,N_13667);
or U14398 (N_14398,N_13085,N_13794);
xnor U14399 (N_14399,N_13882,N_13810);
and U14400 (N_14400,N_13535,N_13818);
or U14401 (N_14401,N_13420,N_13687);
xor U14402 (N_14402,N_13717,N_13499);
nor U14403 (N_14403,N_13486,N_13136);
or U14404 (N_14404,N_13301,N_13021);
or U14405 (N_14405,N_13001,N_13082);
and U14406 (N_14406,N_13191,N_13742);
and U14407 (N_14407,N_13373,N_13894);
and U14408 (N_14408,N_13024,N_13692);
or U14409 (N_14409,N_13647,N_13931);
nand U14410 (N_14410,N_13044,N_13727);
nand U14411 (N_14411,N_13637,N_13578);
or U14412 (N_14412,N_13347,N_13981);
xor U14413 (N_14413,N_13630,N_13141);
nand U14414 (N_14414,N_13065,N_13187);
and U14415 (N_14415,N_13589,N_13249);
nor U14416 (N_14416,N_13621,N_13211);
or U14417 (N_14417,N_13906,N_13260);
and U14418 (N_14418,N_13671,N_13010);
and U14419 (N_14419,N_13558,N_13326);
and U14420 (N_14420,N_13101,N_13183);
and U14421 (N_14421,N_13075,N_13703);
and U14422 (N_14422,N_13516,N_13151);
or U14423 (N_14423,N_13588,N_13394);
xnor U14424 (N_14424,N_13333,N_13226);
nor U14425 (N_14425,N_13518,N_13969);
nor U14426 (N_14426,N_13494,N_13232);
or U14427 (N_14427,N_13662,N_13475);
xor U14428 (N_14428,N_13192,N_13780);
or U14429 (N_14429,N_13828,N_13593);
and U14430 (N_14430,N_13190,N_13348);
and U14431 (N_14431,N_13220,N_13320);
or U14432 (N_14432,N_13940,N_13664);
xor U14433 (N_14433,N_13399,N_13450);
xor U14434 (N_14434,N_13651,N_13858);
or U14435 (N_14435,N_13270,N_13304);
nor U14436 (N_14436,N_13852,N_13070);
and U14437 (N_14437,N_13821,N_13354);
or U14438 (N_14438,N_13689,N_13165);
xnor U14439 (N_14439,N_13944,N_13245);
nor U14440 (N_14440,N_13243,N_13215);
nand U14441 (N_14441,N_13980,N_13091);
or U14442 (N_14442,N_13751,N_13926);
nand U14443 (N_14443,N_13032,N_13459);
nor U14444 (N_14444,N_13257,N_13562);
xor U14445 (N_14445,N_13967,N_13610);
xor U14446 (N_14446,N_13417,N_13120);
or U14447 (N_14447,N_13005,N_13557);
nor U14448 (N_14448,N_13007,N_13472);
nand U14449 (N_14449,N_13360,N_13655);
and U14450 (N_14450,N_13209,N_13602);
xor U14451 (N_14451,N_13682,N_13996);
and U14452 (N_14452,N_13937,N_13680);
nor U14453 (N_14453,N_13195,N_13037);
nand U14454 (N_14454,N_13900,N_13685);
and U14455 (N_14455,N_13108,N_13041);
or U14456 (N_14456,N_13787,N_13436);
nor U14457 (N_14457,N_13161,N_13619);
and U14458 (N_14458,N_13063,N_13611);
xor U14459 (N_14459,N_13104,N_13549);
nor U14460 (N_14460,N_13225,N_13847);
nor U14461 (N_14461,N_13841,N_13203);
nand U14462 (N_14462,N_13855,N_13402);
nand U14463 (N_14463,N_13978,N_13654);
and U14464 (N_14464,N_13470,N_13936);
xnor U14465 (N_14465,N_13512,N_13982);
nand U14466 (N_14466,N_13125,N_13364);
nor U14467 (N_14467,N_13959,N_13030);
nand U14468 (N_14468,N_13297,N_13133);
or U14469 (N_14469,N_13493,N_13375);
nand U14470 (N_14470,N_13329,N_13532);
or U14471 (N_14471,N_13273,N_13299);
nand U14472 (N_14472,N_13850,N_13869);
nor U14473 (N_14473,N_13870,N_13878);
nand U14474 (N_14474,N_13534,N_13236);
nand U14475 (N_14475,N_13572,N_13281);
or U14476 (N_14476,N_13983,N_13724);
and U14477 (N_14477,N_13799,N_13806);
nand U14478 (N_14478,N_13605,N_13452);
nand U14479 (N_14479,N_13624,N_13706);
xnor U14480 (N_14480,N_13251,N_13069);
xor U14481 (N_14481,N_13723,N_13397);
nand U14482 (N_14482,N_13542,N_13434);
nand U14483 (N_14483,N_13418,N_13722);
nand U14484 (N_14484,N_13427,N_13866);
or U14485 (N_14485,N_13167,N_13143);
nand U14486 (N_14486,N_13409,N_13566);
nor U14487 (N_14487,N_13861,N_13994);
nand U14488 (N_14488,N_13350,N_13583);
xor U14489 (N_14489,N_13385,N_13471);
and U14490 (N_14490,N_13786,N_13334);
or U14491 (N_14491,N_13636,N_13634);
nand U14492 (N_14492,N_13684,N_13560);
or U14493 (N_14493,N_13992,N_13949);
nand U14494 (N_14494,N_13600,N_13025);
and U14495 (N_14495,N_13765,N_13880);
and U14496 (N_14496,N_13508,N_13561);
nor U14497 (N_14497,N_13863,N_13539);
and U14498 (N_14498,N_13762,N_13972);
or U14499 (N_14499,N_13934,N_13412);
or U14500 (N_14500,N_13188,N_13340);
or U14501 (N_14501,N_13096,N_13982);
nand U14502 (N_14502,N_13015,N_13813);
and U14503 (N_14503,N_13101,N_13987);
or U14504 (N_14504,N_13620,N_13358);
and U14505 (N_14505,N_13635,N_13853);
nor U14506 (N_14506,N_13629,N_13048);
nand U14507 (N_14507,N_13970,N_13284);
or U14508 (N_14508,N_13889,N_13014);
xnor U14509 (N_14509,N_13592,N_13954);
nor U14510 (N_14510,N_13673,N_13321);
nand U14511 (N_14511,N_13679,N_13520);
xor U14512 (N_14512,N_13913,N_13063);
or U14513 (N_14513,N_13493,N_13757);
nor U14514 (N_14514,N_13134,N_13180);
xnor U14515 (N_14515,N_13432,N_13546);
xor U14516 (N_14516,N_13769,N_13341);
and U14517 (N_14517,N_13626,N_13024);
nor U14518 (N_14518,N_13838,N_13730);
nand U14519 (N_14519,N_13563,N_13582);
xor U14520 (N_14520,N_13205,N_13641);
nand U14521 (N_14521,N_13777,N_13469);
nor U14522 (N_14522,N_13133,N_13571);
xnor U14523 (N_14523,N_13980,N_13240);
nor U14524 (N_14524,N_13453,N_13748);
or U14525 (N_14525,N_13812,N_13372);
nor U14526 (N_14526,N_13100,N_13390);
or U14527 (N_14527,N_13775,N_13416);
or U14528 (N_14528,N_13523,N_13414);
or U14529 (N_14529,N_13543,N_13574);
xor U14530 (N_14530,N_13376,N_13856);
and U14531 (N_14531,N_13526,N_13273);
and U14532 (N_14532,N_13201,N_13978);
or U14533 (N_14533,N_13642,N_13130);
nand U14534 (N_14534,N_13134,N_13112);
or U14535 (N_14535,N_13485,N_13341);
xnor U14536 (N_14536,N_13506,N_13577);
nor U14537 (N_14537,N_13788,N_13198);
xnor U14538 (N_14538,N_13775,N_13158);
xor U14539 (N_14539,N_13045,N_13576);
nand U14540 (N_14540,N_13273,N_13744);
nand U14541 (N_14541,N_13423,N_13603);
or U14542 (N_14542,N_13424,N_13411);
nor U14543 (N_14543,N_13875,N_13296);
nand U14544 (N_14544,N_13846,N_13056);
nor U14545 (N_14545,N_13667,N_13843);
xnor U14546 (N_14546,N_13412,N_13661);
or U14547 (N_14547,N_13274,N_13667);
and U14548 (N_14548,N_13976,N_13459);
nor U14549 (N_14549,N_13965,N_13929);
and U14550 (N_14550,N_13155,N_13474);
xnor U14551 (N_14551,N_13205,N_13138);
and U14552 (N_14552,N_13201,N_13919);
xnor U14553 (N_14553,N_13268,N_13755);
or U14554 (N_14554,N_13968,N_13553);
and U14555 (N_14555,N_13597,N_13349);
nor U14556 (N_14556,N_13146,N_13242);
or U14557 (N_14557,N_13887,N_13806);
nand U14558 (N_14558,N_13524,N_13725);
xor U14559 (N_14559,N_13313,N_13975);
nand U14560 (N_14560,N_13907,N_13996);
and U14561 (N_14561,N_13875,N_13248);
nor U14562 (N_14562,N_13557,N_13977);
and U14563 (N_14563,N_13358,N_13319);
xnor U14564 (N_14564,N_13266,N_13131);
or U14565 (N_14565,N_13952,N_13548);
xnor U14566 (N_14566,N_13631,N_13279);
and U14567 (N_14567,N_13879,N_13676);
nor U14568 (N_14568,N_13590,N_13398);
nor U14569 (N_14569,N_13909,N_13641);
and U14570 (N_14570,N_13014,N_13218);
nand U14571 (N_14571,N_13713,N_13614);
nor U14572 (N_14572,N_13384,N_13332);
nand U14573 (N_14573,N_13631,N_13452);
nor U14574 (N_14574,N_13286,N_13367);
or U14575 (N_14575,N_13868,N_13635);
nor U14576 (N_14576,N_13483,N_13927);
nor U14577 (N_14577,N_13765,N_13830);
or U14578 (N_14578,N_13703,N_13224);
xor U14579 (N_14579,N_13693,N_13454);
nand U14580 (N_14580,N_13560,N_13545);
nor U14581 (N_14581,N_13627,N_13259);
nand U14582 (N_14582,N_13249,N_13138);
or U14583 (N_14583,N_13151,N_13644);
or U14584 (N_14584,N_13384,N_13804);
and U14585 (N_14585,N_13323,N_13172);
or U14586 (N_14586,N_13488,N_13473);
or U14587 (N_14587,N_13312,N_13959);
xor U14588 (N_14588,N_13568,N_13879);
and U14589 (N_14589,N_13532,N_13701);
and U14590 (N_14590,N_13866,N_13592);
nor U14591 (N_14591,N_13852,N_13243);
xnor U14592 (N_14592,N_13535,N_13831);
nor U14593 (N_14593,N_13843,N_13656);
nor U14594 (N_14594,N_13380,N_13160);
or U14595 (N_14595,N_13568,N_13297);
xor U14596 (N_14596,N_13037,N_13859);
nand U14597 (N_14597,N_13720,N_13747);
nand U14598 (N_14598,N_13790,N_13655);
xor U14599 (N_14599,N_13110,N_13730);
or U14600 (N_14600,N_13136,N_13579);
nor U14601 (N_14601,N_13590,N_13312);
nor U14602 (N_14602,N_13238,N_13353);
and U14603 (N_14603,N_13557,N_13716);
nor U14604 (N_14604,N_13181,N_13091);
nand U14605 (N_14605,N_13230,N_13200);
xnor U14606 (N_14606,N_13873,N_13604);
nor U14607 (N_14607,N_13364,N_13706);
or U14608 (N_14608,N_13493,N_13957);
or U14609 (N_14609,N_13367,N_13728);
nand U14610 (N_14610,N_13197,N_13625);
or U14611 (N_14611,N_13393,N_13534);
and U14612 (N_14612,N_13364,N_13508);
nor U14613 (N_14613,N_13000,N_13425);
and U14614 (N_14614,N_13726,N_13802);
nor U14615 (N_14615,N_13727,N_13364);
and U14616 (N_14616,N_13088,N_13374);
nand U14617 (N_14617,N_13318,N_13992);
and U14618 (N_14618,N_13484,N_13365);
or U14619 (N_14619,N_13884,N_13910);
nor U14620 (N_14620,N_13674,N_13364);
or U14621 (N_14621,N_13764,N_13844);
and U14622 (N_14622,N_13527,N_13437);
or U14623 (N_14623,N_13955,N_13280);
and U14624 (N_14624,N_13886,N_13572);
and U14625 (N_14625,N_13602,N_13498);
xor U14626 (N_14626,N_13483,N_13802);
xnor U14627 (N_14627,N_13502,N_13046);
nand U14628 (N_14628,N_13245,N_13179);
or U14629 (N_14629,N_13519,N_13095);
or U14630 (N_14630,N_13360,N_13453);
or U14631 (N_14631,N_13764,N_13101);
or U14632 (N_14632,N_13994,N_13010);
xor U14633 (N_14633,N_13793,N_13880);
or U14634 (N_14634,N_13415,N_13102);
nor U14635 (N_14635,N_13713,N_13401);
or U14636 (N_14636,N_13777,N_13577);
or U14637 (N_14637,N_13835,N_13576);
nand U14638 (N_14638,N_13124,N_13760);
and U14639 (N_14639,N_13576,N_13292);
nor U14640 (N_14640,N_13233,N_13079);
nand U14641 (N_14641,N_13058,N_13396);
xnor U14642 (N_14642,N_13220,N_13350);
nor U14643 (N_14643,N_13438,N_13649);
or U14644 (N_14644,N_13876,N_13471);
or U14645 (N_14645,N_13830,N_13703);
nand U14646 (N_14646,N_13826,N_13563);
nand U14647 (N_14647,N_13663,N_13120);
nor U14648 (N_14648,N_13805,N_13560);
nor U14649 (N_14649,N_13560,N_13349);
nand U14650 (N_14650,N_13083,N_13295);
or U14651 (N_14651,N_13391,N_13728);
and U14652 (N_14652,N_13293,N_13378);
nand U14653 (N_14653,N_13847,N_13921);
nand U14654 (N_14654,N_13223,N_13733);
or U14655 (N_14655,N_13896,N_13421);
and U14656 (N_14656,N_13180,N_13050);
nand U14657 (N_14657,N_13266,N_13098);
or U14658 (N_14658,N_13100,N_13744);
nor U14659 (N_14659,N_13873,N_13815);
nand U14660 (N_14660,N_13499,N_13238);
nor U14661 (N_14661,N_13339,N_13843);
xnor U14662 (N_14662,N_13735,N_13590);
and U14663 (N_14663,N_13980,N_13028);
nand U14664 (N_14664,N_13711,N_13317);
xnor U14665 (N_14665,N_13338,N_13334);
nor U14666 (N_14666,N_13644,N_13714);
xor U14667 (N_14667,N_13601,N_13276);
nor U14668 (N_14668,N_13062,N_13270);
nand U14669 (N_14669,N_13680,N_13084);
and U14670 (N_14670,N_13163,N_13792);
nand U14671 (N_14671,N_13731,N_13779);
and U14672 (N_14672,N_13933,N_13791);
nand U14673 (N_14673,N_13278,N_13634);
nor U14674 (N_14674,N_13263,N_13904);
nand U14675 (N_14675,N_13092,N_13948);
nor U14676 (N_14676,N_13115,N_13985);
nor U14677 (N_14677,N_13064,N_13138);
xnor U14678 (N_14678,N_13967,N_13422);
nand U14679 (N_14679,N_13979,N_13564);
nor U14680 (N_14680,N_13846,N_13038);
nand U14681 (N_14681,N_13965,N_13175);
and U14682 (N_14682,N_13197,N_13824);
or U14683 (N_14683,N_13011,N_13384);
xnor U14684 (N_14684,N_13900,N_13858);
and U14685 (N_14685,N_13554,N_13653);
or U14686 (N_14686,N_13830,N_13808);
or U14687 (N_14687,N_13384,N_13947);
xnor U14688 (N_14688,N_13223,N_13175);
xnor U14689 (N_14689,N_13834,N_13279);
xnor U14690 (N_14690,N_13657,N_13579);
nand U14691 (N_14691,N_13168,N_13200);
xnor U14692 (N_14692,N_13314,N_13677);
nand U14693 (N_14693,N_13451,N_13743);
and U14694 (N_14694,N_13505,N_13005);
nor U14695 (N_14695,N_13782,N_13179);
nor U14696 (N_14696,N_13667,N_13737);
xnor U14697 (N_14697,N_13345,N_13950);
xnor U14698 (N_14698,N_13842,N_13495);
nand U14699 (N_14699,N_13936,N_13069);
nor U14700 (N_14700,N_13235,N_13067);
xnor U14701 (N_14701,N_13089,N_13592);
nand U14702 (N_14702,N_13302,N_13678);
or U14703 (N_14703,N_13316,N_13495);
and U14704 (N_14704,N_13810,N_13939);
xnor U14705 (N_14705,N_13094,N_13991);
or U14706 (N_14706,N_13402,N_13592);
nand U14707 (N_14707,N_13103,N_13606);
xor U14708 (N_14708,N_13901,N_13791);
and U14709 (N_14709,N_13550,N_13644);
or U14710 (N_14710,N_13957,N_13893);
xnor U14711 (N_14711,N_13461,N_13125);
xnor U14712 (N_14712,N_13898,N_13593);
nand U14713 (N_14713,N_13512,N_13242);
and U14714 (N_14714,N_13036,N_13850);
nor U14715 (N_14715,N_13875,N_13257);
xor U14716 (N_14716,N_13902,N_13311);
or U14717 (N_14717,N_13181,N_13624);
nor U14718 (N_14718,N_13189,N_13975);
and U14719 (N_14719,N_13752,N_13873);
xor U14720 (N_14720,N_13836,N_13841);
and U14721 (N_14721,N_13967,N_13688);
and U14722 (N_14722,N_13317,N_13226);
xnor U14723 (N_14723,N_13274,N_13477);
and U14724 (N_14724,N_13139,N_13744);
and U14725 (N_14725,N_13472,N_13351);
and U14726 (N_14726,N_13186,N_13839);
and U14727 (N_14727,N_13254,N_13128);
or U14728 (N_14728,N_13695,N_13855);
or U14729 (N_14729,N_13382,N_13875);
xor U14730 (N_14730,N_13830,N_13078);
xor U14731 (N_14731,N_13255,N_13977);
or U14732 (N_14732,N_13589,N_13580);
and U14733 (N_14733,N_13403,N_13977);
nand U14734 (N_14734,N_13239,N_13819);
nor U14735 (N_14735,N_13044,N_13167);
or U14736 (N_14736,N_13029,N_13380);
or U14737 (N_14737,N_13373,N_13082);
xnor U14738 (N_14738,N_13588,N_13673);
xor U14739 (N_14739,N_13426,N_13560);
xnor U14740 (N_14740,N_13077,N_13629);
nand U14741 (N_14741,N_13915,N_13513);
nand U14742 (N_14742,N_13171,N_13866);
nand U14743 (N_14743,N_13806,N_13601);
xnor U14744 (N_14744,N_13010,N_13674);
and U14745 (N_14745,N_13213,N_13388);
or U14746 (N_14746,N_13436,N_13475);
nand U14747 (N_14747,N_13037,N_13803);
nand U14748 (N_14748,N_13453,N_13257);
xnor U14749 (N_14749,N_13108,N_13106);
and U14750 (N_14750,N_13194,N_13243);
nor U14751 (N_14751,N_13337,N_13528);
nand U14752 (N_14752,N_13560,N_13043);
nor U14753 (N_14753,N_13770,N_13847);
and U14754 (N_14754,N_13466,N_13414);
nor U14755 (N_14755,N_13914,N_13862);
or U14756 (N_14756,N_13876,N_13254);
nor U14757 (N_14757,N_13295,N_13057);
nand U14758 (N_14758,N_13556,N_13795);
nor U14759 (N_14759,N_13766,N_13273);
nor U14760 (N_14760,N_13009,N_13374);
and U14761 (N_14761,N_13070,N_13242);
nand U14762 (N_14762,N_13231,N_13842);
xnor U14763 (N_14763,N_13266,N_13635);
xnor U14764 (N_14764,N_13111,N_13816);
nand U14765 (N_14765,N_13877,N_13282);
nor U14766 (N_14766,N_13518,N_13009);
nand U14767 (N_14767,N_13198,N_13229);
and U14768 (N_14768,N_13167,N_13041);
nor U14769 (N_14769,N_13140,N_13077);
nand U14770 (N_14770,N_13003,N_13851);
xor U14771 (N_14771,N_13014,N_13892);
nor U14772 (N_14772,N_13830,N_13709);
nor U14773 (N_14773,N_13394,N_13501);
and U14774 (N_14774,N_13903,N_13132);
nand U14775 (N_14775,N_13007,N_13519);
and U14776 (N_14776,N_13600,N_13527);
and U14777 (N_14777,N_13836,N_13151);
xor U14778 (N_14778,N_13660,N_13008);
xor U14779 (N_14779,N_13852,N_13744);
nor U14780 (N_14780,N_13557,N_13850);
nand U14781 (N_14781,N_13020,N_13967);
nor U14782 (N_14782,N_13077,N_13167);
xnor U14783 (N_14783,N_13650,N_13274);
or U14784 (N_14784,N_13547,N_13452);
xnor U14785 (N_14785,N_13933,N_13116);
nor U14786 (N_14786,N_13548,N_13141);
and U14787 (N_14787,N_13636,N_13035);
or U14788 (N_14788,N_13205,N_13396);
nand U14789 (N_14789,N_13234,N_13409);
nor U14790 (N_14790,N_13137,N_13507);
nand U14791 (N_14791,N_13835,N_13665);
nand U14792 (N_14792,N_13454,N_13133);
nor U14793 (N_14793,N_13595,N_13106);
xor U14794 (N_14794,N_13563,N_13321);
or U14795 (N_14795,N_13484,N_13556);
or U14796 (N_14796,N_13752,N_13937);
and U14797 (N_14797,N_13633,N_13050);
or U14798 (N_14798,N_13953,N_13139);
xor U14799 (N_14799,N_13325,N_13840);
nand U14800 (N_14800,N_13020,N_13515);
xor U14801 (N_14801,N_13454,N_13559);
nand U14802 (N_14802,N_13780,N_13727);
and U14803 (N_14803,N_13370,N_13419);
and U14804 (N_14804,N_13592,N_13393);
or U14805 (N_14805,N_13009,N_13305);
xor U14806 (N_14806,N_13600,N_13383);
xnor U14807 (N_14807,N_13331,N_13492);
nor U14808 (N_14808,N_13072,N_13743);
nor U14809 (N_14809,N_13794,N_13186);
and U14810 (N_14810,N_13670,N_13527);
xnor U14811 (N_14811,N_13399,N_13716);
nand U14812 (N_14812,N_13882,N_13776);
or U14813 (N_14813,N_13629,N_13509);
nand U14814 (N_14814,N_13849,N_13991);
and U14815 (N_14815,N_13214,N_13998);
nand U14816 (N_14816,N_13510,N_13411);
and U14817 (N_14817,N_13111,N_13383);
and U14818 (N_14818,N_13847,N_13198);
nor U14819 (N_14819,N_13168,N_13846);
nand U14820 (N_14820,N_13107,N_13559);
xnor U14821 (N_14821,N_13321,N_13733);
or U14822 (N_14822,N_13929,N_13164);
or U14823 (N_14823,N_13491,N_13537);
nand U14824 (N_14824,N_13835,N_13432);
and U14825 (N_14825,N_13515,N_13259);
and U14826 (N_14826,N_13357,N_13956);
nor U14827 (N_14827,N_13108,N_13738);
or U14828 (N_14828,N_13527,N_13928);
nor U14829 (N_14829,N_13691,N_13269);
nand U14830 (N_14830,N_13115,N_13703);
nand U14831 (N_14831,N_13959,N_13996);
nor U14832 (N_14832,N_13777,N_13410);
nor U14833 (N_14833,N_13201,N_13273);
nand U14834 (N_14834,N_13792,N_13253);
xor U14835 (N_14835,N_13337,N_13836);
and U14836 (N_14836,N_13291,N_13063);
or U14837 (N_14837,N_13716,N_13407);
nand U14838 (N_14838,N_13238,N_13051);
or U14839 (N_14839,N_13382,N_13842);
and U14840 (N_14840,N_13133,N_13746);
and U14841 (N_14841,N_13894,N_13039);
nand U14842 (N_14842,N_13677,N_13654);
xnor U14843 (N_14843,N_13929,N_13737);
and U14844 (N_14844,N_13106,N_13911);
and U14845 (N_14845,N_13811,N_13772);
nand U14846 (N_14846,N_13242,N_13561);
nand U14847 (N_14847,N_13371,N_13389);
or U14848 (N_14848,N_13662,N_13146);
nand U14849 (N_14849,N_13044,N_13123);
xnor U14850 (N_14850,N_13166,N_13710);
and U14851 (N_14851,N_13814,N_13240);
or U14852 (N_14852,N_13299,N_13238);
and U14853 (N_14853,N_13642,N_13557);
or U14854 (N_14854,N_13126,N_13154);
nor U14855 (N_14855,N_13449,N_13007);
nand U14856 (N_14856,N_13336,N_13649);
nand U14857 (N_14857,N_13242,N_13191);
nand U14858 (N_14858,N_13197,N_13342);
nor U14859 (N_14859,N_13673,N_13899);
and U14860 (N_14860,N_13948,N_13753);
and U14861 (N_14861,N_13550,N_13421);
xor U14862 (N_14862,N_13315,N_13010);
nand U14863 (N_14863,N_13907,N_13316);
xnor U14864 (N_14864,N_13233,N_13287);
and U14865 (N_14865,N_13701,N_13065);
nand U14866 (N_14866,N_13935,N_13670);
nand U14867 (N_14867,N_13012,N_13816);
or U14868 (N_14868,N_13516,N_13745);
nor U14869 (N_14869,N_13039,N_13047);
and U14870 (N_14870,N_13972,N_13669);
or U14871 (N_14871,N_13967,N_13403);
xnor U14872 (N_14872,N_13554,N_13692);
and U14873 (N_14873,N_13944,N_13361);
or U14874 (N_14874,N_13836,N_13319);
nor U14875 (N_14875,N_13745,N_13474);
nand U14876 (N_14876,N_13850,N_13501);
nor U14877 (N_14877,N_13268,N_13431);
nand U14878 (N_14878,N_13276,N_13730);
nand U14879 (N_14879,N_13696,N_13045);
nand U14880 (N_14880,N_13634,N_13341);
nor U14881 (N_14881,N_13931,N_13269);
xor U14882 (N_14882,N_13500,N_13205);
or U14883 (N_14883,N_13891,N_13264);
xor U14884 (N_14884,N_13921,N_13924);
and U14885 (N_14885,N_13132,N_13491);
xnor U14886 (N_14886,N_13270,N_13442);
nor U14887 (N_14887,N_13472,N_13230);
xor U14888 (N_14888,N_13334,N_13607);
nor U14889 (N_14889,N_13596,N_13162);
and U14890 (N_14890,N_13079,N_13427);
xnor U14891 (N_14891,N_13366,N_13352);
xnor U14892 (N_14892,N_13510,N_13079);
or U14893 (N_14893,N_13641,N_13689);
nor U14894 (N_14894,N_13476,N_13314);
nand U14895 (N_14895,N_13750,N_13071);
or U14896 (N_14896,N_13161,N_13170);
and U14897 (N_14897,N_13520,N_13403);
nor U14898 (N_14898,N_13389,N_13387);
nand U14899 (N_14899,N_13073,N_13006);
nor U14900 (N_14900,N_13833,N_13420);
or U14901 (N_14901,N_13616,N_13628);
nor U14902 (N_14902,N_13759,N_13831);
nor U14903 (N_14903,N_13683,N_13098);
nor U14904 (N_14904,N_13844,N_13742);
nand U14905 (N_14905,N_13821,N_13981);
nor U14906 (N_14906,N_13595,N_13140);
xnor U14907 (N_14907,N_13253,N_13164);
nand U14908 (N_14908,N_13129,N_13620);
or U14909 (N_14909,N_13252,N_13677);
and U14910 (N_14910,N_13101,N_13124);
and U14911 (N_14911,N_13725,N_13479);
xnor U14912 (N_14912,N_13332,N_13186);
xnor U14913 (N_14913,N_13876,N_13724);
nand U14914 (N_14914,N_13502,N_13774);
and U14915 (N_14915,N_13960,N_13373);
and U14916 (N_14916,N_13998,N_13791);
and U14917 (N_14917,N_13430,N_13376);
xor U14918 (N_14918,N_13551,N_13471);
or U14919 (N_14919,N_13408,N_13825);
xor U14920 (N_14920,N_13969,N_13508);
xnor U14921 (N_14921,N_13452,N_13953);
or U14922 (N_14922,N_13638,N_13454);
or U14923 (N_14923,N_13098,N_13578);
xnor U14924 (N_14924,N_13296,N_13089);
and U14925 (N_14925,N_13319,N_13250);
and U14926 (N_14926,N_13995,N_13709);
nor U14927 (N_14927,N_13530,N_13416);
nand U14928 (N_14928,N_13319,N_13737);
and U14929 (N_14929,N_13067,N_13403);
nand U14930 (N_14930,N_13398,N_13069);
nor U14931 (N_14931,N_13004,N_13049);
nor U14932 (N_14932,N_13841,N_13482);
and U14933 (N_14933,N_13708,N_13422);
xor U14934 (N_14934,N_13583,N_13242);
and U14935 (N_14935,N_13205,N_13425);
xnor U14936 (N_14936,N_13728,N_13086);
xnor U14937 (N_14937,N_13970,N_13122);
or U14938 (N_14938,N_13474,N_13725);
nor U14939 (N_14939,N_13093,N_13374);
nand U14940 (N_14940,N_13425,N_13541);
and U14941 (N_14941,N_13995,N_13994);
nand U14942 (N_14942,N_13533,N_13722);
nand U14943 (N_14943,N_13584,N_13362);
or U14944 (N_14944,N_13162,N_13735);
and U14945 (N_14945,N_13388,N_13841);
nand U14946 (N_14946,N_13206,N_13516);
and U14947 (N_14947,N_13987,N_13554);
nor U14948 (N_14948,N_13624,N_13478);
xor U14949 (N_14949,N_13470,N_13685);
or U14950 (N_14950,N_13353,N_13225);
nor U14951 (N_14951,N_13438,N_13221);
xor U14952 (N_14952,N_13889,N_13754);
or U14953 (N_14953,N_13285,N_13151);
or U14954 (N_14954,N_13002,N_13552);
nand U14955 (N_14955,N_13099,N_13020);
xnor U14956 (N_14956,N_13123,N_13370);
and U14957 (N_14957,N_13530,N_13161);
nand U14958 (N_14958,N_13216,N_13496);
xor U14959 (N_14959,N_13320,N_13820);
xor U14960 (N_14960,N_13180,N_13283);
xnor U14961 (N_14961,N_13882,N_13994);
and U14962 (N_14962,N_13986,N_13568);
nor U14963 (N_14963,N_13546,N_13398);
and U14964 (N_14964,N_13199,N_13655);
or U14965 (N_14965,N_13757,N_13826);
or U14966 (N_14966,N_13344,N_13836);
and U14967 (N_14967,N_13537,N_13091);
or U14968 (N_14968,N_13049,N_13383);
nor U14969 (N_14969,N_13894,N_13349);
and U14970 (N_14970,N_13909,N_13453);
nand U14971 (N_14971,N_13413,N_13316);
nand U14972 (N_14972,N_13760,N_13248);
or U14973 (N_14973,N_13051,N_13624);
nand U14974 (N_14974,N_13103,N_13043);
nand U14975 (N_14975,N_13870,N_13865);
xor U14976 (N_14976,N_13670,N_13737);
nand U14977 (N_14977,N_13490,N_13760);
and U14978 (N_14978,N_13910,N_13113);
xor U14979 (N_14979,N_13234,N_13844);
xor U14980 (N_14980,N_13993,N_13303);
xnor U14981 (N_14981,N_13860,N_13381);
or U14982 (N_14982,N_13225,N_13817);
and U14983 (N_14983,N_13631,N_13803);
or U14984 (N_14984,N_13441,N_13400);
xnor U14985 (N_14985,N_13915,N_13639);
nor U14986 (N_14986,N_13845,N_13450);
nand U14987 (N_14987,N_13156,N_13381);
nand U14988 (N_14988,N_13911,N_13772);
nor U14989 (N_14989,N_13941,N_13598);
nand U14990 (N_14990,N_13663,N_13611);
nor U14991 (N_14991,N_13735,N_13723);
xor U14992 (N_14992,N_13221,N_13812);
or U14993 (N_14993,N_13808,N_13190);
nand U14994 (N_14994,N_13348,N_13850);
nor U14995 (N_14995,N_13052,N_13714);
nand U14996 (N_14996,N_13967,N_13549);
or U14997 (N_14997,N_13429,N_13197);
and U14998 (N_14998,N_13282,N_13725);
xor U14999 (N_14999,N_13916,N_13784);
and U15000 (N_15000,N_14819,N_14991);
nand U15001 (N_15001,N_14737,N_14671);
or U15002 (N_15002,N_14237,N_14486);
and U15003 (N_15003,N_14846,N_14868);
xor U15004 (N_15004,N_14653,N_14851);
nand U15005 (N_15005,N_14973,N_14919);
and U15006 (N_15006,N_14173,N_14692);
nand U15007 (N_15007,N_14383,N_14764);
xnor U15008 (N_15008,N_14338,N_14368);
xor U15009 (N_15009,N_14392,N_14298);
xnor U15010 (N_15010,N_14801,N_14594);
nor U15011 (N_15011,N_14472,N_14260);
or U15012 (N_15012,N_14906,N_14204);
xnor U15013 (N_15013,N_14591,N_14966);
nand U15014 (N_15014,N_14954,N_14208);
nand U15015 (N_15015,N_14573,N_14342);
nand U15016 (N_15016,N_14274,N_14353);
and U15017 (N_15017,N_14960,N_14610);
and U15018 (N_15018,N_14092,N_14993);
nand U15019 (N_15019,N_14125,N_14878);
xnor U15020 (N_15020,N_14654,N_14159);
or U15021 (N_15021,N_14041,N_14038);
nor U15022 (N_15022,N_14155,N_14069);
nor U15023 (N_15023,N_14563,N_14174);
nor U15024 (N_15024,N_14992,N_14169);
xnor U15025 (N_15025,N_14347,N_14782);
or U15026 (N_15026,N_14139,N_14218);
or U15027 (N_15027,N_14776,N_14238);
and U15028 (N_15028,N_14754,N_14874);
or U15029 (N_15029,N_14912,N_14437);
nor U15030 (N_15030,N_14939,N_14430);
nand U15031 (N_15031,N_14224,N_14048);
nand U15032 (N_15032,N_14194,N_14081);
nor U15033 (N_15033,N_14447,N_14718);
or U15034 (N_15034,N_14351,N_14371);
and U15035 (N_15035,N_14134,N_14748);
nor U15036 (N_15036,N_14757,N_14297);
and U15037 (N_15037,N_14651,N_14883);
xor U15038 (N_15038,N_14561,N_14207);
and U15039 (N_15039,N_14168,N_14617);
nand U15040 (N_15040,N_14699,N_14181);
xnor U15041 (N_15041,N_14427,N_14147);
nor U15042 (N_15042,N_14149,N_14106);
and U15043 (N_15043,N_14549,N_14229);
or U15044 (N_15044,N_14952,N_14049);
nor U15045 (N_15045,N_14201,N_14997);
nor U15046 (N_15046,N_14643,N_14900);
and U15047 (N_15047,N_14683,N_14184);
xor U15048 (N_15048,N_14557,N_14070);
xor U15049 (N_15049,N_14312,N_14836);
nor U15050 (N_15050,N_14290,N_14166);
or U15051 (N_15051,N_14924,N_14894);
and U15052 (N_15052,N_14859,N_14235);
xnor U15053 (N_15053,N_14161,N_14592);
nand U15054 (N_15054,N_14625,N_14632);
xnor U15055 (N_15055,N_14619,N_14817);
or U15056 (N_15056,N_14690,N_14119);
or U15057 (N_15057,N_14828,N_14571);
nand U15058 (N_15058,N_14216,N_14225);
or U15059 (N_15059,N_14132,N_14334);
and U15060 (N_15060,N_14087,N_14405);
nor U15061 (N_15061,N_14027,N_14256);
nand U15062 (N_15062,N_14964,N_14475);
nor U15063 (N_15063,N_14882,N_14620);
and U15064 (N_15064,N_14996,N_14967);
xnor U15065 (N_15065,N_14163,N_14156);
and U15066 (N_15066,N_14527,N_14525);
or U15067 (N_15067,N_14073,N_14465);
xnor U15068 (N_15068,N_14463,N_14792);
and U15069 (N_15069,N_14877,N_14955);
nand U15070 (N_15070,N_14300,N_14953);
nand U15071 (N_15071,N_14917,N_14309);
or U15072 (N_15072,N_14470,N_14120);
xnor U15073 (N_15073,N_14506,N_14323);
or U15074 (N_15074,N_14822,N_14382);
nand U15075 (N_15075,N_14986,N_14228);
xnor U15076 (N_15076,N_14698,N_14056);
and U15077 (N_15077,N_14408,N_14213);
nand U15078 (N_15078,N_14553,N_14321);
xor U15079 (N_15079,N_14700,N_14179);
and U15080 (N_15080,N_14037,N_14773);
or U15081 (N_15081,N_14865,N_14372);
and U15082 (N_15082,N_14708,N_14880);
nand U15083 (N_15083,N_14262,N_14394);
nor U15084 (N_15084,N_14978,N_14626);
xnor U15085 (N_15085,N_14729,N_14043);
or U15086 (N_15086,N_14790,N_14283);
nor U15087 (N_15087,N_14121,N_14640);
nor U15088 (N_15088,N_14258,N_14257);
and U15089 (N_15089,N_14249,N_14143);
nand U15090 (N_15090,N_14407,N_14903);
or U15091 (N_15091,N_14328,N_14602);
nand U15092 (N_15092,N_14449,N_14908);
nand U15093 (N_15093,N_14493,N_14325);
and U15094 (N_15094,N_14936,N_14870);
and U15095 (N_15095,N_14058,N_14129);
nand U15096 (N_15096,N_14809,N_14433);
and U15097 (N_15097,N_14178,N_14646);
nor U15098 (N_15098,N_14293,N_14462);
nor U15099 (N_15099,N_14971,N_14974);
nor U15100 (N_15100,N_14086,N_14999);
and U15101 (N_15101,N_14886,N_14580);
nand U15102 (N_15102,N_14963,N_14341);
nand U15103 (N_15103,N_14855,N_14582);
or U15104 (N_15104,N_14720,N_14250);
xor U15105 (N_15105,N_14652,N_14417);
xnor U15106 (N_15106,N_14768,N_14703);
and U15107 (N_15107,N_14907,N_14306);
nand U15108 (N_15108,N_14196,N_14667);
nor U15109 (N_15109,N_14375,N_14324);
and U15110 (N_15110,N_14876,N_14487);
and U15111 (N_15111,N_14236,N_14827);
xnor U15112 (N_15112,N_14858,N_14649);
and U15113 (N_15113,N_14932,N_14872);
and U15114 (N_15114,N_14969,N_14558);
and U15115 (N_15115,N_14674,N_14977);
and U15116 (N_15116,N_14047,N_14336);
and U15117 (N_15117,N_14248,N_14590);
xor U15118 (N_15118,N_14404,N_14403);
or U15119 (N_15119,N_14024,N_14148);
nand U15120 (N_15120,N_14255,N_14787);
or U15121 (N_15121,N_14473,N_14210);
nor U15122 (N_15122,N_14630,N_14477);
nor U15123 (N_15123,N_14280,N_14252);
or U15124 (N_15124,N_14150,N_14152);
nand U15125 (N_15125,N_14655,N_14818);
nor U15126 (N_15126,N_14076,N_14844);
nor U15127 (N_15127,N_14937,N_14440);
xor U15128 (N_15128,N_14537,N_14541);
and U15129 (N_15129,N_14175,N_14975);
xnor U15130 (N_15130,N_14396,N_14253);
nor U15131 (N_15131,N_14740,N_14095);
nor U15132 (N_15132,N_14489,N_14352);
nor U15133 (N_15133,N_14555,N_14284);
xor U15134 (N_15134,N_14164,N_14562);
nor U15135 (N_15135,N_14744,N_14534);
and U15136 (N_15136,N_14837,N_14616);
and U15137 (N_15137,N_14202,N_14856);
and U15138 (N_15138,N_14581,N_14866);
nand U15139 (N_15139,N_14222,N_14522);
nor U15140 (N_15140,N_14116,N_14722);
xor U15141 (N_15141,N_14415,N_14310);
xor U15142 (N_15142,N_14084,N_14554);
xor U15143 (N_15143,N_14063,N_14188);
or U15144 (N_15144,N_14521,N_14454);
nor U15145 (N_15145,N_14854,N_14520);
or U15146 (N_15146,N_14266,N_14777);
or U15147 (N_15147,N_14881,N_14285);
and U15148 (N_15148,N_14459,N_14244);
xnor U15149 (N_15149,N_14714,N_14313);
nor U15150 (N_15150,N_14998,N_14045);
nand U15151 (N_15151,N_14367,N_14711);
and U15152 (N_15152,N_14781,N_14439);
and U15153 (N_15153,N_14055,N_14545);
and U15154 (N_15154,N_14614,N_14395);
nand U15155 (N_15155,N_14171,N_14526);
and U15156 (N_15156,N_14438,N_14896);
and U15157 (N_15157,N_14778,N_14765);
nand U15158 (N_15158,N_14685,N_14798);
or U15159 (N_15159,N_14186,N_14034);
or U15160 (N_15160,N_14593,N_14431);
nor U15161 (N_15161,N_14731,N_14595);
nand U15162 (N_15162,N_14420,N_14990);
nand U15163 (N_15163,N_14374,N_14752);
and U15164 (N_15164,N_14017,N_14004);
xnor U15165 (N_15165,N_14314,N_14468);
and U15166 (N_15166,N_14810,N_14915);
xnor U15167 (N_15167,N_14606,N_14206);
xnor U15168 (N_15168,N_14968,N_14343);
or U15169 (N_15169,N_14108,N_14390);
xnor U15170 (N_15170,N_14267,N_14833);
and U15171 (N_15171,N_14605,N_14240);
nor U15172 (N_15172,N_14904,N_14769);
and U15173 (N_15173,N_14763,N_14679);
and U15174 (N_15174,N_14887,N_14215);
and U15175 (N_15175,N_14421,N_14035);
nor U15176 (N_15176,N_14745,N_14838);
xnor U15177 (N_15177,N_14816,N_14586);
nor U15178 (N_15178,N_14361,N_14780);
or U15179 (N_15179,N_14976,N_14232);
and U15180 (N_15180,N_14388,N_14067);
xnor U15181 (N_15181,N_14721,N_14344);
or U15182 (N_15182,N_14962,N_14185);
xor U15183 (N_15183,N_14425,N_14085);
nand U15184 (N_15184,N_14712,N_14270);
nor U15185 (N_15185,N_14281,N_14268);
nand U15186 (N_15186,N_14369,N_14613);
and U15187 (N_15187,N_14277,N_14009);
nand U15188 (N_15188,N_14766,N_14197);
or U15189 (N_15189,N_14808,N_14137);
or U15190 (N_15190,N_14423,N_14584);
xnor U15191 (N_15191,N_14016,N_14516);
xnor U15192 (N_15192,N_14519,N_14317);
or U15193 (N_15193,N_14219,N_14189);
xnor U15194 (N_15194,N_14354,N_14355);
nor U15195 (N_15195,N_14448,N_14302);
nor U15196 (N_15196,N_14066,N_14378);
nand U15197 (N_15197,N_14287,N_14012);
nor U15198 (N_15198,N_14538,N_14669);
nor U15199 (N_15199,N_14981,N_14141);
nand U15200 (N_15200,N_14788,N_14406);
and U15201 (N_15201,N_14029,N_14938);
and U15202 (N_15202,N_14071,N_14124);
and U15203 (N_15203,N_14411,N_14949);
xor U15204 (N_15204,N_14400,N_14303);
xor U15205 (N_15205,N_14741,N_14536);
nor U15206 (N_15206,N_14020,N_14205);
or U15207 (N_15207,N_14743,N_14001);
nor U15208 (N_15208,N_14589,N_14869);
nor U15209 (N_15209,N_14501,N_14133);
xor U15210 (N_15210,N_14771,N_14820);
xnor U15211 (N_15211,N_14840,N_14693);
xnor U15212 (N_15212,N_14456,N_14180);
nor U15213 (N_15213,N_14040,N_14126);
nor U15214 (N_15214,N_14299,N_14362);
nand U15215 (N_15215,N_14412,N_14665);
nor U15216 (N_15216,N_14760,N_14504);
and U15217 (N_15217,N_14621,N_14793);
or U15218 (N_15218,N_14660,N_14663);
or U15219 (N_15219,N_14103,N_14572);
nand U15220 (N_15220,N_14985,N_14755);
or U15221 (N_15221,N_14018,N_14770);
and U15222 (N_15222,N_14366,N_14570);
and U15223 (N_15223,N_14989,N_14596);
nand U15224 (N_15224,N_14730,N_14146);
or U15225 (N_15225,N_14025,N_14631);
or U15226 (N_15226,N_14933,N_14127);
or U15227 (N_15227,N_14370,N_14011);
nand U15228 (N_15228,N_14987,N_14320);
xor U15229 (N_15229,N_14107,N_14686);
nand U15230 (N_15230,N_14588,N_14226);
or U15231 (N_15231,N_14072,N_14661);
nand U15232 (N_15232,N_14233,N_14387);
or U15233 (N_15233,N_14359,N_14023);
or U15234 (N_15234,N_14995,N_14575);
and U15235 (N_15235,N_14873,N_14241);
nand U15236 (N_15236,N_14805,N_14062);
nor U15237 (N_15237,N_14007,N_14672);
xor U15238 (N_15238,N_14598,N_14191);
xor U15239 (N_15239,N_14791,N_14416);
nor U15240 (N_15240,N_14746,N_14158);
and U15241 (N_15241,N_14641,N_14847);
xor U15242 (N_15242,N_14078,N_14157);
xnor U15243 (N_15243,N_14532,N_14920);
nor U15244 (N_15244,N_14079,N_14867);
nand U15245 (N_15245,N_14142,N_14322);
nand U15246 (N_15246,N_14719,N_14734);
nand U15247 (N_15247,N_14559,N_14576);
nand U15248 (N_15248,N_14909,N_14892);
and U15249 (N_15249,N_14102,N_14587);
nand U15250 (N_15250,N_14825,N_14348);
and U15251 (N_15251,N_14871,N_14494);
nor U15252 (N_15252,N_14203,N_14318);
xnor U15253 (N_15253,N_14065,N_14453);
xor U15254 (N_15254,N_14294,N_14128);
and U15255 (N_15255,N_14162,N_14929);
xor U15256 (N_15256,N_14508,N_14360);
and U15257 (N_15257,N_14008,N_14272);
xnor U15258 (N_15258,N_14524,N_14888);
nand U15259 (N_15259,N_14019,N_14650);
nand U15260 (N_15260,N_14339,N_14357);
or U15261 (N_15261,N_14376,N_14167);
or U15262 (N_15262,N_14824,N_14583);
nand U15263 (N_15263,N_14381,N_14409);
xnor U15264 (N_15264,N_14402,N_14261);
nor U15265 (N_15265,N_14002,N_14443);
nor U15266 (N_15266,N_14807,N_14481);
or U15267 (N_15267,N_14511,N_14796);
or U15268 (N_15268,N_14279,N_14278);
or U15269 (N_15269,N_14850,N_14227);
nor U15270 (N_15270,N_14217,N_14221);
xor U15271 (N_15271,N_14623,N_14467);
or U15272 (N_15272,N_14544,N_14944);
nor U15273 (N_15273,N_14308,N_14889);
and U15274 (N_15274,N_14057,N_14391);
and U15275 (N_15275,N_14350,N_14926);
xnor U15276 (N_15276,N_14502,N_14492);
xor U15277 (N_15277,N_14988,N_14678);
xor U15278 (N_15278,N_14797,N_14327);
or U15279 (N_15279,N_14356,N_14223);
nor U15280 (N_15280,N_14109,N_14957);
nand U15281 (N_15281,N_14922,N_14145);
xor U15282 (N_15282,N_14895,N_14499);
and U15283 (N_15283,N_14728,N_14947);
xor U15284 (N_15284,N_14154,N_14435);
or U15285 (N_15285,N_14961,N_14483);
nor U15286 (N_15286,N_14529,N_14951);
xnor U15287 (N_15287,N_14635,N_14172);
and U15288 (N_15288,N_14068,N_14265);
xnor U15289 (N_15289,N_14612,N_14136);
or U15290 (N_15290,N_14577,N_14014);
xnor U15291 (N_15291,N_14775,N_14264);
nand U15292 (N_15292,N_14662,N_14751);
xor U15293 (N_15293,N_14445,N_14688);
xor U15294 (N_15294,N_14422,N_14015);
or U15295 (N_15295,N_14694,N_14050);
and U15296 (N_15296,N_14622,N_14239);
nor U15297 (N_15297,N_14916,N_14160);
xnor U15298 (N_15298,N_14668,N_14940);
and U15299 (N_15299,N_14498,N_14419);
or U15300 (N_15300,N_14080,N_14677);
nand U15301 (N_15301,N_14315,N_14736);
nand U15302 (N_15302,N_14935,N_14607);
nor U15303 (N_15303,N_14377,N_14384);
and U15304 (N_15304,N_14330,N_14785);
nor U15305 (N_15305,N_14316,N_14113);
xor U15306 (N_15306,N_14512,N_14902);
nand U15307 (N_15307,N_14091,N_14311);
nand U15308 (N_15308,N_14738,N_14097);
xnor U15309 (N_15309,N_14689,N_14183);
nor U15310 (N_15310,N_14064,N_14861);
nand U15311 (N_15311,N_14636,N_14259);
or U15312 (N_15312,N_14893,N_14531);
or U15313 (N_15313,N_14604,N_14681);
nor U15314 (N_15314,N_14735,N_14611);
nor U15315 (N_15315,N_14021,N_14638);
nand U15316 (N_15316,N_14211,N_14182);
or U15317 (N_15317,N_14444,N_14032);
nor U15318 (N_15318,N_14263,N_14138);
nor U15319 (N_15319,N_14082,N_14042);
xnor U15320 (N_15320,N_14251,N_14424);
nor U15321 (N_15321,N_14931,N_14495);
nand U15322 (N_15322,N_14905,N_14918);
xor U15323 (N_15323,N_14601,N_14083);
and U15324 (N_15324,N_14634,N_14701);
and U15325 (N_15325,N_14784,N_14476);
xor U15326 (N_15326,N_14845,N_14254);
nor U15327 (N_15327,N_14296,N_14212);
xor U15328 (N_15328,N_14418,N_14676);
and U15329 (N_15329,N_14659,N_14835);
and U15330 (N_15330,N_14863,N_14565);
and U15331 (N_15331,N_14715,N_14637);
and U15332 (N_15332,N_14972,N_14105);
xnor U15333 (N_15333,N_14560,N_14564);
nor U15334 (N_15334,N_14648,N_14276);
xor U15335 (N_15335,N_14984,N_14839);
xor U15336 (N_15336,N_14717,N_14513);
xor U15337 (N_15337,N_14460,N_14923);
and U15338 (N_15338,N_14994,N_14795);
nand U15339 (N_15339,N_14135,N_14273);
or U15340 (N_15340,N_14786,N_14115);
xor U15341 (N_15341,N_14275,N_14709);
xnor U15342 (N_15342,N_14812,N_14026);
nand U15343 (N_15343,N_14505,N_14089);
xor U15344 (N_15344,N_14242,N_14941);
and U15345 (N_15345,N_14547,N_14518);
and U15346 (N_15346,N_14800,N_14710);
xnor U15347 (N_15347,N_14428,N_14666);
and U15348 (N_15348,N_14245,N_14144);
or U15349 (N_15349,N_14772,N_14639);
nand U15350 (N_15350,N_14096,N_14195);
nand U15351 (N_15351,N_14053,N_14429);
nand U15352 (N_15352,N_14762,N_14603);
nand U15353 (N_15353,N_14482,N_14691);
nand U15354 (N_15354,N_14958,N_14200);
or U15355 (N_15355,N_14434,N_14829);
xor U15356 (N_15356,N_14455,N_14331);
nor U15357 (N_15357,N_14140,N_14335);
nor U15358 (N_15358,N_14658,N_14288);
nand U15359 (N_15359,N_14177,N_14899);
or U15360 (N_15360,N_14852,N_14891);
xnor U15361 (N_15361,N_14804,N_14304);
nand U15362 (N_15362,N_14857,N_14118);
and U15363 (N_15363,N_14705,N_14243);
and U15364 (N_15364,N_14644,N_14684);
nand U15365 (N_15365,N_14401,N_14077);
xor U15366 (N_15366,N_14811,N_14380);
nor U15367 (N_15367,N_14530,N_14497);
or U15368 (N_15368,N_14373,N_14340);
or U15369 (N_15369,N_14843,N_14758);
or U15370 (N_15370,N_14507,N_14059);
xnor U15371 (N_15371,N_14286,N_14704);
and U15372 (N_15372,N_14488,N_14231);
xnor U15373 (N_15373,N_14333,N_14442);
or U15374 (N_15374,N_14815,N_14618);
nor U15375 (N_15375,N_14830,N_14187);
and U15376 (N_15376,N_14193,N_14673);
or U15377 (N_15377,N_14696,N_14170);
and U15378 (N_15378,N_14291,N_14664);
nand U15379 (N_15379,N_14597,N_14033);
nor U15380 (N_15380,N_14123,N_14329);
nor U15381 (N_15381,N_14724,N_14979);
and U15382 (N_15382,N_14198,N_14849);
xnor U15383 (N_15383,N_14911,N_14122);
and U15384 (N_15384,N_14295,N_14948);
and U15385 (N_15385,N_14432,N_14413);
or U15386 (N_15386,N_14337,N_14956);
nor U15387 (N_15387,N_14946,N_14379);
xor U15388 (N_15388,N_14733,N_14950);
and U15389 (N_15389,N_14457,N_14036);
and U15390 (N_15390,N_14345,N_14551);
or U15391 (N_15391,N_14358,N_14864);
and U15392 (N_15392,N_14365,N_14980);
xnor U15393 (N_15393,N_14490,N_14841);
nand U15394 (N_15394,N_14750,N_14441);
nand U15395 (N_15395,N_14398,N_14307);
and U15396 (N_15396,N_14474,N_14389);
and U15397 (N_15397,N_14052,N_14742);
nor U15398 (N_15398,N_14542,N_14890);
nor U15399 (N_15399,N_14051,N_14657);
nand U15400 (N_15400,N_14970,N_14624);
xnor U15401 (N_15401,N_14176,N_14680);
nor U15402 (N_15402,N_14028,N_14509);
nor U15403 (N_15403,N_14633,N_14647);
nand U15404 (N_15404,N_14117,N_14292);
nand U15405 (N_15405,N_14656,N_14496);
nand U15406 (N_15406,N_14615,N_14451);
or U15407 (N_15407,N_14569,N_14627);
nor U15408 (N_15408,N_14349,N_14723);
xor U15409 (N_15409,N_14479,N_14747);
and U15410 (N_15410,N_14727,N_14151);
xor U15411 (N_15411,N_14774,N_14713);
xor U15412 (N_15412,N_14862,N_14585);
or U15413 (N_15413,N_14675,N_14707);
nor U15414 (N_15414,N_14914,N_14943);
or U15415 (N_15415,N_14461,N_14190);
nand U15416 (N_15416,N_14271,N_14875);
or U15417 (N_15417,N_14094,N_14523);
nand U15418 (N_15418,N_14061,N_14884);
nand U15419 (N_15419,N_14925,N_14165);
or U15420 (N_15420,N_14716,N_14921);
nand U15421 (N_15421,N_14739,N_14054);
and U15422 (N_15422,N_14199,N_14111);
and U15423 (N_15423,N_14214,N_14848);
xor U15424 (N_15424,N_14060,N_14568);
xor U15425 (N_15425,N_14897,N_14075);
xnor U15426 (N_15426,N_14006,N_14927);
xnor U15427 (N_15427,N_14794,N_14399);
nor U15428 (N_15428,N_14130,N_14697);
or U15429 (N_15429,N_14753,N_14885);
or U15430 (N_15430,N_14806,N_14942);
and U15431 (N_15431,N_14528,N_14393);
or U15432 (N_15432,N_14574,N_14458);
nor U15433 (N_15433,N_14789,N_14823);
nor U15434 (N_15434,N_14983,N_14834);
nand U15435 (N_15435,N_14514,N_14234);
xor U15436 (N_15436,N_14725,N_14687);
or U15437 (N_15437,N_14552,N_14030);
or U15438 (N_15438,N_14799,N_14093);
xnor U15439 (N_15439,N_14044,N_14230);
xnor U15440 (N_15440,N_14578,N_14670);
nor U15441 (N_15441,N_14192,N_14548);
xor U15442 (N_15442,N_14879,N_14289);
and U15443 (N_15443,N_14515,N_14599);
nand U15444 (N_15444,N_14579,N_14114);
nand U15445 (N_15445,N_14860,N_14543);
or U15446 (N_15446,N_14510,N_14756);
and U15447 (N_15447,N_14556,N_14101);
or U15448 (N_15448,N_14682,N_14550);
nor U15449 (N_15449,N_14491,N_14153);
xor U15450 (N_15450,N_14484,N_14100);
xnor U15451 (N_15451,N_14842,N_14803);
xor U15452 (N_15452,N_14464,N_14046);
or U15453 (N_15453,N_14645,N_14098);
or U15454 (N_15454,N_14003,N_14022);
or U15455 (N_15455,N_14832,N_14783);
nand U15456 (N_15456,N_14246,N_14749);
or U15457 (N_15457,N_14090,N_14301);
and U15458 (N_15458,N_14831,N_14385);
and U15459 (N_15459,N_14898,N_14517);
nand U15460 (N_15460,N_14629,N_14959);
xnor U15461 (N_15461,N_14364,N_14104);
nand U15462 (N_15462,N_14546,N_14220);
xor U15463 (N_15463,N_14363,N_14500);
and U15464 (N_15464,N_14540,N_14934);
and U15465 (N_15465,N_14600,N_14013);
xor U15466 (N_15466,N_14131,N_14469);
xor U15467 (N_15467,N_14539,N_14965);
nor U15468 (N_15468,N_14695,N_14319);
or U15469 (N_15469,N_14779,N_14928);
or U15470 (N_15470,N_14269,N_14000);
and U15471 (N_15471,N_14567,N_14346);
or U15472 (N_15472,N_14426,N_14913);
nor U15473 (N_15473,N_14628,N_14031);
and U15474 (N_15474,N_14566,N_14386);
and U15475 (N_15475,N_14282,N_14110);
nor U15476 (N_15476,N_14397,N_14326);
and U15477 (N_15477,N_14450,N_14813);
nor U15478 (N_15478,N_14074,N_14247);
xor U15479 (N_15479,N_14802,N_14010);
or U15480 (N_15480,N_14732,N_14332);
xor U15481 (N_15481,N_14466,N_14814);
xor U15482 (N_15482,N_14726,N_14471);
xor U15483 (N_15483,N_14702,N_14112);
and U15484 (N_15484,N_14099,N_14005);
xor U15485 (N_15485,N_14452,N_14767);
nand U15486 (N_15486,N_14901,N_14414);
and U15487 (N_15487,N_14826,N_14821);
xnor U15488 (N_15488,N_14088,N_14039);
xnor U15489 (N_15489,N_14642,N_14945);
nor U15490 (N_15490,N_14485,N_14608);
xor U15491 (N_15491,N_14478,N_14982);
nand U15492 (N_15492,N_14853,N_14761);
nand U15493 (N_15493,N_14503,N_14209);
xnor U15494 (N_15494,N_14706,N_14305);
xnor U15495 (N_15495,N_14609,N_14910);
and U15496 (N_15496,N_14436,N_14410);
nand U15497 (N_15497,N_14759,N_14535);
and U15498 (N_15498,N_14446,N_14480);
and U15499 (N_15499,N_14930,N_14533);
or U15500 (N_15500,N_14971,N_14631);
and U15501 (N_15501,N_14138,N_14241);
and U15502 (N_15502,N_14399,N_14205);
or U15503 (N_15503,N_14765,N_14148);
and U15504 (N_15504,N_14577,N_14496);
nor U15505 (N_15505,N_14301,N_14371);
or U15506 (N_15506,N_14643,N_14349);
nand U15507 (N_15507,N_14959,N_14194);
and U15508 (N_15508,N_14678,N_14278);
xnor U15509 (N_15509,N_14129,N_14424);
nor U15510 (N_15510,N_14861,N_14234);
and U15511 (N_15511,N_14152,N_14828);
and U15512 (N_15512,N_14504,N_14090);
nand U15513 (N_15513,N_14507,N_14197);
or U15514 (N_15514,N_14756,N_14196);
nand U15515 (N_15515,N_14900,N_14394);
and U15516 (N_15516,N_14111,N_14420);
nand U15517 (N_15517,N_14238,N_14581);
or U15518 (N_15518,N_14733,N_14931);
nand U15519 (N_15519,N_14863,N_14173);
or U15520 (N_15520,N_14138,N_14770);
xnor U15521 (N_15521,N_14429,N_14769);
nor U15522 (N_15522,N_14745,N_14207);
and U15523 (N_15523,N_14876,N_14189);
xor U15524 (N_15524,N_14168,N_14680);
or U15525 (N_15525,N_14403,N_14925);
xnor U15526 (N_15526,N_14050,N_14775);
and U15527 (N_15527,N_14618,N_14164);
or U15528 (N_15528,N_14884,N_14832);
nand U15529 (N_15529,N_14597,N_14528);
or U15530 (N_15530,N_14062,N_14754);
or U15531 (N_15531,N_14354,N_14845);
and U15532 (N_15532,N_14207,N_14377);
and U15533 (N_15533,N_14596,N_14390);
and U15534 (N_15534,N_14634,N_14508);
nor U15535 (N_15535,N_14226,N_14554);
nor U15536 (N_15536,N_14731,N_14097);
and U15537 (N_15537,N_14968,N_14576);
and U15538 (N_15538,N_14237,N_14751);
xor U15539 (N_15539,N_14288,N_14316);
nor U15540 (N_15540,N_14020,N_14235);
and U15541 (N_15541,N_14083,N_14079);
xnor U15542 (N_15542,N_14232,N_14873);
and U15543 (N_15543,N_14004,N_14432);
xnor U15544 (N_15544,N_14339,N_14221);
nor U15545 (N_15545,N_14705,N_14953);
nor U15546 (N_15546,N_14838,N_14897);
nand U15547 (N_15547,N_14120,N_14726);
nand U15548 (N_15548,N_14224,N_14256);
or U15549 (N_15549,N_14915,N_14179);
xor U15550 (N_15550,N_14282,N_14874);
nand U15551 (N_15551,N_14970,N_14944);
and U15552 (N_15552,N_14859,N_14064);
nor U15553 (N_15553,N_14633,N_14941);
nor U15554 (N_15554,N_14942,N_14871);
or U15555 (N_15555,N_14691,N_14289);
and U15556 (N_15556,N_14869,N_14249);
nor U15557 (N_15557,N_14015,N_14750);
xor U15558 (N_15558,N_14249,N_14451);
or U15559 (N_15559,N_14925,N_14220);
xnor U15560 (N_15560,N_14598,N_14414);
or U15561 (N_15561,N_14375,N_14653);
xnor U15562 (N_15562,N_14346,N_14884);
nand U15563 (N_15563,N_14537,N_14785);
nor U15564 (N_15564,N_14540,N_14606);
xor U15565 (N_15565,N_14530,N_14672);
xor U15566 (N_15566,N_14787,N_14174);
nor U15567 (N_15567,N_14078,N_14238);
and U15568 (N_15568,N_14640,N_14983);
xnor U15569 (N_15569,N_14251,N_14817);
and U15570 (N_15570,N_14359,N_14342);
and U15571 (N_15571,N_14868,N_14496);
nor U15572 (N_15572,N_14344,N_14048);
nor U15573 (N_15573,N_14642,N_14903);
xnor U15574 (N_15574,N_14255,N_14933);
xnor U15575 (N_15575,N_14436,N_14552);
or U15576 (N_15576,N_14327,N_14860);
nor U15577 (N_15577,N_14700,N_14247);
nand U15578 (N_15578,N_14112,N_14732);
and U15579 (N_15579,N_14602,N_14054);
and U15580 (N_15580,N_14091,N_14940);
and U15581 (N_15581,N_14551,N_14676);
nor U15582 (N_15582,N_14934,N_14617);
or U15583 (N_15583,N_14729,N_14265);
xor U15584 (N_15584,N_14133,N_14002);
or U15585 (N_15585,N_14950,N_14354);
or U15586 (N_15586,N_14371,N_14014);
xnor U15587 (N_15587,N_14190,N_14145);
nand U15588 (N_15588,N_14617,N_14214);
nand U15589 (N_15589,N_14079,N_14828);
or U15590 (N_15590,N_14128,N_14251);
or U15591 (N_15591,N_14837,N_14994);
nor U15592 (N_15592,N_14394,N_14803);
nor U15593 (N_15593,N_14789,N_14357);
nand U15594 (N_15594,N_14677,N_14721);
nor U15595 (N_15595,N_14423,N_14133);
nand U15596 (N_15596,N_14774,N_14000);
xor U15597 (N_15597,N_14325,N_14951);
or U15598 (N_15598,N_14536,N_14663);
xor U15599 (N_15599,N_14052,N_14496);
or U15600 (N_15600,N_14334,N_14852);
xnor U15601 (N_15601,N_14606,N_14554);
and U15602 (N_15602,N_14955,N_14884);
nor U15603 (N_15603,N_14005,N_14508);
or U15604 (N_15604,N_14337,N_14033);
xor U15605 (N_15605,N_14734,N_14128);
nand U15606 (N_15606,N_14686,N_14499);
xor U15607 (N_15607,N_14944,N_14266);
and U15608 (N_15608,N_14872,N_14915);
nor U15609 (N_15609,N_14952,N_14934);
nand U15610 (N_15610,N_14155,N_14249);
nand U15611 (N_15611,N_14000,N_14956);
and U15612 (N_15612,N_14837,N_14146);
and U15613 (N_15613,N_14881,N_14737);
nor U15614 (N_15614,N_14686,N_14415);
xnor U15615 (N_15615,N_14848,N_14580);
xor U15616 (N_15616,N_14946,N_14503);
or U15617 (N_15617,N_14393,N_14159);
nand U15618 (N_15618,N_14444,N_14522);
nand U15619 (N_15619,N_14388,N_14400);
and U15620 (N_15620,N_14641,N_14305);
nand U15621 (N_15621,N_14207,N_14868);
xnor U15622 (N_15622,N_14722,N_14062);
and U15623 (N_15623,N_14438,N_14155);
nor U15624 (N_15624,N_14780,N_14981);
and U15625 (N_15625,N_14680,N_14815);
or U15626 (N_15626,N_14178,N_14773);
and U15627 (N_15627,N_14470,N_14258);
nor U15628 (N_15628,N_14872,N_14876);
and U15629 (N_15629,N_14529,N_14715);
nand U15630 (N_15630,N_14927,N_14086);
and U15631 (N_15631,N_14944,N_14309);
and U15632 (N_15632,N_14385,N_14300);
and U15633 (N_15633,N_14585,N_14379);
or U15634 (N_15634,N_14057,N_14684);
xnor U15635 (N_15635,N_14574,N_14651);
or U15636 (N_15636,N_14300,N_14313);
and U15637 (N_15637,N_14711,N_14539);
nor U15638 (N_15638,N_14288,N_14387);
nand U15639 (N_15639,N_14462,N_14003);
or U15640 (N_15640,N_14645,N_14972);
nand U15641 (N_15641,N_14531,N_14135);
and U15642 (N_15642,N_14562,N_14137);
and U15643 (N_15643,N_14159,N_14617);
nand U15644 (N_15644,N_14121,N_14034);
xor U15645 (N_15645,N_14177,N_14684);
nor U15646 (N_15646,N_14451,N_14469);
or U15647 (N_15647,N_14379,N_14858);
nor U15648 (N_15648,N_14999,N_14119);
and U15649 (N_15649,N_14740,N_14893);
nor U15650 (N_15650,N_14317,N_14240);
or U15651 (N_15651,N_14031,N_14105);
or U15652 (N_15652,N_14576,N_14241);
and U15653 (N_15653,N_14338,N_14162);
or U15654 (N_15654,N_14082,N_14808);
or U15655 (N_15655,N_14352,N_14479);
and U15656 (N_15656,N_14302,N_14977);
nor U15657 (N_15657,N_14322,N_14390);
xnor U15658 (N_15658,N_14750,N_14880);
nor U15659 (N_15659,N_14968,N_14842);
xnor U15660 (N_15660,N_14034,N_14443);
or U15661 (N_15661,N_14881,N_14167);
and U15662 (N_15662,N_14480,N_14563);
nand U15663 (N_15663,N_14229,N_14028);
or U15664 (N_15664,N_14824,N_14856);
or U15665 (N_15665,N_14351,N_14839);
and U15666 (N_15666,N_14627,N_14550);
nor U15667 (N_15667,N_14675,N_14421);
or U15668 (N_15668,N_14909,N_14654);
nand U15669 (N_15669,N_14563,N_14048);
xor U15670 (N_15670,N_14433,N_14191);
and U15671 (N_15671,N_14207,N_14293);
nand U15672 (N_15672,N_14585,N_14558);
xnor U15673 (N_15673,N_14111,N_14870);
nand U15674 (N_15674,N_14747,N_14712);
and U15675 (N_15675,N_14205,N_14076);
and U15676 (N_15676,N_14700,N_14403);
or U15677 (N_15677,N_14542,N_14419);
xnor U15678 (N_15678,N_14462,N_14260);
nand U15679 (N_15679,N_14427,N_14582);
or U15680 (N_15680,N_14496,N_14838);
nand U15681 (N_15681,N_14890,N_14446);
nand U15682 (N_15682,N_14517,N_14587);
nor U15683 (N_15683,N_14570,N_14799);
nand U15684 (N_15684,N_14595,N_14039);
and U15685 (N_15685,N_14524,N_14463);
and U15686 (N_15686,N_14156,N_14853);
and U15687 (N_15687,N_14127,N_14810);
nor U15688 (N_15688,N_14993,N_14586);
or U15689 (N_15689,N_14396,N_14398);
xor U15690 (N_15690,N_14731,N_14037);
and U15691 (N_15691,N_14724,N_14179);
or U15692 (N_15692,N_14584,N_14107);
and U15693 (N_15693,N_14310,N_14265);
xnor U15694 (N_15694,N_14805,N_14545);
nor U15695 (N_15695,N_14155,N_14990);
xnor U15696 (N_15696,N_14751,N_14315);
xnor U15697 (N_15697,N_14380,N_14992);
nor U15698 (N_15698,N_14543,N_14512);
nor U15699 (N_15699,N_14255,N_14292);
nor U15700 (N_15700,N_14508,N_14659);
xor U15701 (N_15701,N_14379,N_14813);
xor U15702 (N_15702,N_14140,N_14249);
xnor U15703 (N_15703,N_14904,N_14298);
nor U15704 (N_15704,N_14483,N_14266);
or U15705 (N_15705,N_14420,N_14164);
or U15706 (N_15706,N_14571,N_14181);
xor U15707 (N_15707,N_14242,N_14040);
and U15708 (N_15708,N_14081,N_14342);
and U15709 (N_15709,N_14934,N_14197);
and U15710 (N_15710,N_14705,N_14905);
nor U15711 (N_15711,N_14528,N_14509);
or U15712 (N_15712,N_14647,N_14550);
nor U15713 (N_15713,N_14481,N_14199);
nor U15714 (N_15714,N_14378,N_14573);
nor U15715 (N_15715,N_14869,N_14947);
nand U15716 (N_15716,N_14274,N_14142);
nand U15717 (N_15717,N_14510,N_14121);
nand U15718 (N_15718,N_14977,N_14931);
nor U15719 (N_15719,N_14486,N_14946);
nand U15720 (N_15720,N_14913,N_14390);
nand U15721 (N_15721,N_14450,N_14323);
nand U15722 (N_15722,N_14473,N_14213);
nand U15723 (N_15723,N_14872,N_14387);
xor U15724 (N_15724,N_14433,N_14975);
nor U15725 (N_15725,N_14976,N_14271);
nand U15726 (N_15726,N_14481,N_14874);
xor U15727 (N_15727,N_14717,N_14160);
or U15728 (N_15728,N_14225,N_14030);
or U15729 (N_15729,N_14754,N_14929);
xor U15730 (N_15730,N_14083,N_14033);
nor U15731 (N_15731,N_14048,N_14696);
and U15732 (N_15732,N_14533,N_14817);
or U15733 (N_15733,N_14610,N_14637);
and U15734 (N_15734,N_14763,N_14748);
or U15735 (N_15735,N_14330,N_14797);
or U15736 (N_15736,N_14403,N_14237);
xnor U15737 (N_15737,N_14357,N_14320);
xor U15738 (N_15738,N_14549,N_14396);
and U15739 (N_15739,N_14382,N_14655);
nor U15740 (N_15740,N_14268,N_14066);
and U15741 (N_15741,N_14158,N_14574);
nor U15742 (N_15742,N_14454,N_14039);
or U15743 (N_15743,N_14793,N_14020);
xor U15744 (N_15744,N_14096,N_14615);
and U15745 (N_15745,N_14918,N_14924);
or U15746 (N_15746,N_14713,N_14740);
xnor U15747 (N_15747,N_14207,N_14220);
nor U15748 (N_15748,N_14621,N_14274);
or U15749 (N_15749,N_14288,N_14652);
or U15750 (N_15750,N_14011,N_14521);
nor U15751 (N_15751,N_14489,N_14134);
nor U15752 (N_15752,N_14450,N_14886);
nor U15753 (N_15753,N_14893,N_14804);
nand U15754 (N_15754,N_14498,N_14912);
nor U15755 (N_15755,N_14983,N_14811);
nor U15756 (N_15756,N_14876,N_14464);
and U15757 (N_15757,N_14897,N_14981);
or U15758 (N_15758,N_14254,N_14410);
nand U15759 (N_15759,N_14985,N_14343);
nand U15760 (N_15760,N_14085,N_14334);
and U15761 (N_15761,N_14626,N_14419);
nand U15762 (N_15762,N_14859,N_14181);
and U15763 (N_15763,N_14880,N_14557);
and U15764 (N_15764,N_14665,N_14852);
nor U15765 (N_15765,N_14217,N_14570);
or U15766 (N_15766,N_14749,N_14912);
and U15767 (N_15767,N_14400,N_14743);
xnor U15768 (N_15768,N_14329,N_14642);
xnor U15769 (N_15769,N_14175,N_14259);
nor U15770 (N_15770,N_14593,N_14166);
xor U15771 (N_15771,N_14442,N_14978);
or U15772 (N_15772,N_14522,N_14281);
xnor U15773 (N_15773,N_14006,N_14899);
and U15774 (N_15774,N_14538,N_14310);
or U15775 (N_15775,N_14178,N_14409);
and U15776 (N_15776,N_14810,N_14513);
and U15777 (N_15777,N_14079,N_14964);
and U15778 (N_15778,N_14144,N_14347);
nand U15779 (N_15779,N_14232,N_14868);
nor U15780 (N_15780,N_14562,N_14859);
nor U15781 (N_15781,N_14224,N_14818);
or U15782 (N_15782,N_14693,N_14189);
nand U15783 (N_15783,N_14760,N_14331);
or U15784 (N_15784,N_14046,N_14936);
or U15785 (N_15785,N_14545,N_14592);
nor U15786 (N_15786,N_14971,N_14935);
nand U15787 (N_15787,N_14428,N_14361);
nand U15788 (N_15788,N_14356,N_14149);
nor U15789 (N_15789,N_14936,N_14639);
nor U15790 (N_15790,N_14067,N_14926);
nor U15791 (N_15791,N_14944,N_14429);
nand U15792 (N_15792,N_14000,N_14977);
and U15793 (N_15793,N_14772,N_14561);
xnor U15794 (N_15794,N_14837,N_14510);
or U15795 (N_15795,N_14658,N_14463);
and U15796 (N_15796,N_14246,N_14680);
xor U15797 (N_15797,N_14147,N_14395);
nor U15798 (N_15798,N_14157,N_14311);
or U15799 (N_15799,N_14753,N_14546);
xnor U15800 (N_15800,N_14750,N_14074);
and U15801 (N_15801,N_14436,N_14818);
nand U15802 (N_15802,N_14891,N_14381);
xor U15803 (N_15803,N_14493,N_14712);
xor U15804 (N_15804,N_14967,N_14702);
and U15805 (N_15805,N_14505,N_14473);
nand U15806 (N_15806,N_14666,N_14273);
nand U15807 (N_15807,N_14356,N_14912);
and U15808 (N_15808,N_14935,N_14380);
and U15809 (N_15809,N_14723,N_14418);
nor U15810 (N_15810,N_14115,N_14127);
and U15811 (N_15811,N_14377,N_14687);
and U15812 (N_15812,N_14753,N_14999);
or U15813 (N_15813,N_14170,N_14085);
nor U15814 (N_15814,N_14974,N_14408);
xor U15815 (N_15815,N_14545,N_14664);
nand U15816 (N_15816,N_14355,N_14477);
and U15817 (N_15817,N_14336,N_14951);
nor U15818 (N_15818,N_14338,N_14437);
nand U15819 (N_15819,N_14356,N_14675);
and U15820 (N_15820,N_14040,N_14042);
nand U15821 (N_15821,N_14363,N_14820);
nand U15822 (N_15822,N_14812,N_14244);
xnor U15823 (N_15823,N_14981,N_14797);
xor U15824 (N_15824,N_14158,N_14915);
nand U15825 (N_15825,N_14054,N_14052);
xor U15826 (N_15826,N_14783,N_14927);
nor U15827 (N_15827,N_14928,N_14100);
xor U15828 (N_15828,N_14893,N_14640);
nor U15829 (N_15829,N_14310,N_14300);
xor U15830 (N_15830,N_14995,N_14703);
or U15831 (N_15831,N_14184,N_14089);
nor U15832 (N_15832,N_14530,N_14777);
nor U15833 (N_15833,N_14958,N_14717);
nand U15834 (N_15834,N_14568,N_14464);
or U15835 (N_15835,N_14952,N_14732);
nor U15836 (N_15836,N_14826,N_14096);
nor U15837 (N_15837,N_14642,N_14259);
or U15838 (N_15838,N_14173,N_14630);
xnor U15839 (N_15839,N_14352,N_14257);
nor U15840 (N_15840,N_14226,N_14132);
nand U15841 (N_15841,N_14496,N_14606);
xnor U15842 (N_15842,N_14699,N_14465);
and U15843 (N_15843,N_14262,N_14806);
nand U15844 (N_15844,N_14127,N_14654);
nand U15845 (N_15845,N_14896,N_14684);
or U15846 (N_15846,N_14271,N_14747);
nor U15847 (N_15847,N_14644,N_14466);
or U15848 (N_15848,N_14467,N_14063);
xnor U15849 (N_15849,N_14862,N_14708);
xnor U15850 (N_15850,N_14218,N_14840);
and U15851 (N_15851,N_14545,N_14709);
nand U15852 (N_15852,N_14090,N_14159);
nand U15853 (N_15853,N_14362,N_14283);
nor U15854 (N_15854,N_14577,N_14344);
xnor U15855 (N_15855,N_14977,N_14482);
or U15856 (N_15856,N_14308,N_14960);
nand U15857 (N_15857,N_14877,N_14299);
nor U15858 (N_15858,N_14336,N_14177);
and U15859 (N_15859,N_14439,N_14269);
and U15860 (N_15860,N_14491,N_14443);
or U15861 (N_15861,N_14646,N_14700);
or U15862 (N_15862,N_14312,N_14662);
or U15863 (N_15863,N_14222,N_14302);
nor U15864 (N_15864,N_14880,N_14546);
or U15865 (N_15865,N_14007,N_14291);
nor U15866 (N_15866,N_14240,N_14976);
and U15867 (N_15867,N_14575,N_14738);
nand U15868 (N_15868,N_14113,N_14053);
and U15869 (N_15869,N_14686,N_14249);
and U15870 (N_15870,N_14678,N_14566);
nor U15871 (N_15871,N_14678,N_14627);
nor U15872 (N_15872,N_14163,N_14168);
xnor U15873 (N_15873,N_14774,N_14071);
nand U15874 (N_15874,N_14886,N_14856);
nor U15875 (N_15875,N_14830,N_14159);
nand U15876 (N_15876,N_14845,N_14509);
nand U15877 (N_15877,N_14439,N_14466);
and U15878 (N_15878,N_14763,N_14437);
and U15879 (N_15879,N_14204,N_14379);
and U15880 (N_15880,N_14560,N_14149);
and U15881 (N_15881,N_14274,N_14437);
nand U15882 (N_15882,N_14056,N_14378);
xor U15883 (N_15883,N_14860,N_14233);
nand U15884 (N_15884,N_14693,N_14134);
and U15885 (N_15885,N_14102,N_14754);
and U15886 (N_15886,N_14787,N_14979);
and U15887 (N_15887,N_14576,N_14990);
xnor U15888 (N_15888,N_14015,N_14442);
nor U15889 (N_15889,N_14697,N_14224);
or U15890 (N_15890,N_14423,N_14496);
xnor U15891 (N_15891,N_14783,N_14382);
or U15892 (N_15892,N_14068,N_14624);
xor U15893 (N_15893,N_14978,N_14844);
nand U15894 (N_15894,N_14952,N_14043);
or U15895 (N_15895,N_14107,N_14479);
nor U15896 (N_15896,N_14857,N_14485);
or U15897 (N_15897,N_14328,N_14961);
nand U15898 (N_15898,N_14381,N_14054);
nand U15899 (N_15899,N_14316,N_14531);
nor U15900 (N_15900,N_14512,N_14805);
xor U15901 (N_15901,N_14301,N_14785);
and U15902 (N_15902,N_14313,N_14256);
nor U15903 (N_15903,N_14518,N_14324);
and U15904 (N_15904,N_14636,N_14984);
nor U15905 (N_15905,N_14979,N_14341);
nor U15906 (N_15906,N_14323,N_14847);
xor U15907 (N_15907,N_14113,N_14157);
or U15908 (N_15908,N_14118,N_14545);
or U15909 (N_15909,N_14931,N_14757);
nor U15910 (N_15910,N_14195,N_14757);
nand U15911 (N_15911,N_14391,N_14561);
nor U15912 (N_15912,N_14461,N_14390);
nor U15913 (N_15913,N_14050,N_14403);
or U15914 (N_15914,N_14272,N_14876);
xnor U15915 (N_15915,N_14684,N_14116);
and U15916 (N_15916,N_14116,N_14310);
nand U15917 (N_15917,N_14139,N_14209);
nor U15918 (N_15918,N_14742,N_14094);
or U15919 (N_15919,N_14242,N_14541);
and U15920 (N_15920,N_14071,N_14390);
or U15921 (N_15921,N_14704,N_14788);
or U15922 (N_15922,N_14331,N_14627);
or U15923 (N_15923,N_14580,N_14667);
or U15924 (N_15924,N_14426,N_14110);
nor U15925 (N_15925,N_14160,N_14013);
xor U15926 (N_15926,N_14230,N_14812);
nor U15927 (N_15927,N_14413,N_14073);
and U15928 (N_15928,N_14381,N_14477);
xor U15929 (N_15929,N_14011,N_14978);
nand U15930 (N_15930,N_14944,N_14177);
nand U15931 (N_15931,N_14078,N_14965);
nor U15932 (N_15932,N_14573,N_14011);
xnor U15933 (N_15933,N_14593,N_14836);
nor U15934 (N_15934,N_14914,N_14912);
nand U15935 (N_15935,N_14365,N_14083);
nand U15936 (N_15936,N_14407,N_14808);
or U15937 (N_15937,N_14339,N_14386);
or U15938 (N_15938,N_14342,N_14476);
and U15939 (N_15939,N_14288,N_14472);
nor U15940 (N_15940,N_14888,N_14351);
xnor U15941 (N_15941,N_14667,N_14996);
nand U15942 (N_15942,N_14175,N_14009);
and U15943 (N_15943,N_14051,N_14383);
and U15944 (N_15944,N_14892,N_14466);
nor U15945 (N_15945,N_14122,N_14715);
and U15946 (N_15946,N_14983,N_14961);
or U15947 (N_15947,N_14281,N_14116);
nor U15948 (N_15948,N_14990,N_14407);
or U15949 (N_15949,N_14434,N_14219);
or U15950 (N_15950,N_14068,N_14192);
nor U15951 (N_15951,N_14305,N_14491);
nand U15952 (N_15952,N_14802,N_14579);
xor U15953 (N_15953,N_14439,N_14131);
xor U15954 (N_15954,N_14983,N_14549);
nor U15955 (N_15955,N_14983,N_14654);
nor U15956 (N_15956,N_14112,N_14989);
and U15957 (N_15957,N_14214,N_14180);
nor U15958 (N_15958,N_14403,N_14177);
nand U15959 (N_15959,N_14222,N_14012);
or U15960 (N_15960,N_14347,N_14119);
and U15961 (N_15961,N_14770,N_14569);
nand U15962 (N_15962,N_14892,N_14131);
nor U15963 (N_15963,N_14515,N_14677);
xor U15964 (N_15964,N_14768,N_14801);
xor U15965 (N_15965,N_14808,N_14966);
nor U15966 (N_15966,N_14016,N_14331);
and U15967 (N_15967,N_14953,N_14447);
and U15968 (N_15968,N_14337,N_14490);
or U15969 (N_15969,N_14245,N_14397);
and U15970 (N_15970,N_14099,N_14411);
or U15971 (N_15971,N_14719,N_14729);
and U15972 (N_15972,N_14218,N_14779);
xnor U15973 (N_15973,N_14794,N_14866);
nand U15974 (N_15974,N_14872,N_14814);
or U15975 (N_15975,N_14651,N_14554);
or U15976 (N_15976,N_14705,N_14416);
or U15977 (N_15977,N_14670,N_14879);
and U15978 (N_15978,N_14128,N_14572);
nor U15979 (N_15979,N_14601,N_14388);
and U15980 (N_15980,N_14990,N_14766);
and U15981 (N_15981,N_14089,N_14156);
nor U15982 (N_15982,N_14274,N_14186);
xnor U15983 (N_15983,N_14616,N_14940);
nand U15984 (N_15984,N_14495,N_14892);
nand U15985 (N_15985,N_14389,N_14663);
xor U15986 (N_15986,N_14342,N_14271);
nor U15987 (N_15987,N_14658,N_14483);
xor U15988 (N_15988,N_14287,N_14343);
nor U15989 (N_15989,N_14807,N_14583);
nor U15990 (N_15990,N_14536,N_14042);
and U15991 (N_15991,N_14657,N_14625);
and U15992 (N_15992,N_14414,N_14137);
and U15993 (N_15993,N_14897,N_14032);
or U15994 (N_15994,N_14823,N_14816);
or U15995 (N_15995,N_14798,N_14781);
or U15996 (N_15996,N_14908,N_14057);
nor U15997 (N_15997,N_14296,N_14277);
nor U15998 (N_15998,N_14082,N_14286);
and U15999 (N_15999,N_14689,N_14144);
xor U16000 (N_16000,N_15707,N_15696);
xnor U16001 (N_16001,N_15799,N_15263);
xor U16002 (N_16002,N_15964,N_15672);
and U16003 (N_16003,N_15265,N_15302);
and U16004 (N_16004,N_15908,N_15213);
nand U16005 (N_16005,N_15088,N_15418);
xnor U16006 (N_16006,N_15045,N_15516);
and U16007 (N_16007,N_15085,N_15327);
nand U16008 (N_16008,N_15087,N_15862);
or U16009 (N_16009,N_15639,N_15453);
xnor U16010 (N_16010,N_15595,N_15950);
and U16011 (N_16011,N_15977,N_15976);
nand U16012 (N_16012,N_15973,N_15369);
nand U16013 (N_16013,N_15670,N_15214);
xor U16014 (N_16014,N_15103,N_15067);
nor U16015 (N_16015,N_15482,N_15511);
xnor U16016 (N_16016,N_15250,N_15972);
nor U16017 (N_16017,N_15996,N_15926);
nor U16018 (N_16018,N_15613,N_15424);
nor U16019 (N_16019,N_15824,N_15141);
xor U16020 (N_16020,N_15392,N_15134);
and U16021 (N_16021,N_15106,N_15589);
or U16022 (N_16022,N_15512,N_15069);
nand U16023 (N_16023,N_15929,N_15682);
nand U16024 (N_16024,N_15312,N_15017);
or U16025 (N_16025,N_15710,N_15115);
xor U16026 (N_16026,N_15391,N_15281);
nor U16027 (N_16027,N_15959,N_15660);
or U16028 (N_16028,N_15695,N_15366);
nand U16029 (N_16029,N_15025,N_15947);
xor U16030 (N_16030,N_15162,N_15731);
and U16031 (N_16031,N_15374,N_15687);
xor U16032 (N_16032,N_15494,N_15782);
xnor U16033 (N_16033,N_15989,N_15870);
and U16034 (N_16034,N_15669,N_15264);
nor U16035 (N_16035,N_15365,N_15328);
nor U16036 (N_16036,N_15411,N_15320);
or U16037 (N_16037,N_15933,N_15384);
or U16038 (N_16038,N_15757,N_15754);
xor U16039 (N_16039,N_15838,N_15075);
or U16040 (N_16040,N_15130,N_15771);
nand U16041 (N_16041,N_15598,N_15079);
nand U16042 (N_16042,N_15431,N_15561);
or U16043 (N_16043,N_15258,N_15129);
xor U16044 (N_16044,N_15186,N_15225);
or U16045 (N_16045,N_15305,N_15153);
xnor U16046 (N_16046,N_15139,N_15237);
xor U16047 (N_16047,N_15458,N_15316);
xnor U16048 (N_16048,N_15904,N_15405);
and U16049 (N_16049,N_15415,N_15789);
and U16050 (N_16050,N_15448,N_15556);
nor U16051 (N_16051,N_15519,N_15994);
nor U16052 (N_16052,N_15887,N_15545);
xor U16053 (N_16053,N_15402,N_15636);
and U16054 (N_16054,N_15676,N_15109);
nor U16055 (N_16055,N_15168,N_15289);
nor U16056 (N_16056,N_15603,N_15260);
or U16057 (N_16057,N_15196,N_15205);
xor U16058 (N_16058,N_15954,N_15428);
nand U16059 (N_16059,N_15201,N_15946);
xor U16060 (N_16060,N_15536,N_15801);
xor U16061 (N_16061,N_15764,N_15744);
nand U16062 (N_16062,N_15648,N_15591);
nand U16063 (N_16063,N_15299,N_15429);
xor U16064 (N_16064,N_15247,N_15403);
nand U16065 (N_16065,N_15357,N_15283);
or U16066 (N_16066,N_15863,N_15037);
nand U16067 (N_16067,N_15203,N_15664);
nor U16068 (N_16068,N_15271,N_15578);
xor U16069 (N_16069,N_15029,N_15066);
xnor U16070 (N_16070,N_15057,N_15112);
xor U16071 (N_16071,N_15319,N_15766);
nor U16072 (N_16072,N_15637,N_15301);
nor U16073 (N_16073,N_15315,N_15163);
xor U16074 (N_16074,N_15416,N_15108);
and U16075 (N_16075,N_15097,N_15035);
and U16076 (N_16076,N_15845,N_15548);
or U16077 (N_16077,N_15261,N_15704);
and U16078 (N_16078,N_15308,N_15174);
nand U16079 (N_16079,N_15387,N_15086);
nand U16080 (N_16080,N_15834,N_15177);
nor U16081 (N_16081,N_15490,N_15126);
nand U16082 (N_16082,N_15787,N_15767);
xor U16083 (N_16083,N_15313,N_15449);
nand U16084 (N_16084,N_15122,N_15630);
nand U16085 (N_16085,N_15641,N_15846);
xnor U16086 (N_16086,N_15331,N_15063);
nor U16087 (N_16087,N_15812,N_15893);
nand U16088 (N_16088,N_15456,N_15004);
nand U16089 (N_16089,N_15988,N_15509);
or U16090 (N_16090,N_15282,N_15667);
nor U16091 (N_16091,N_15781,N_15323);
nor U16092 (N_16092,N_15071,N_15951);
nand U16093 (N_16093,N_15111,N_15379);
or U16094 (N_16094,N_15161,N_15350);
xnor U16095 (N_16095,N_15635,N_15593);
and U16096 (N_16096,N_15124,N_15249);
and U16097 (N_16097,N_15193,N_15318);
nand U16098 (N_16098,N_15625,N_15277);
or U16099 (N_16099,N_15464,N_15851);
nor U16100 (N_16100,N_15463,N_15276);
and U16101 (N_16101,N_15525,N_15987);
and U16102 (N_16102,N_15114,N_15955);
nand U16103 (N_16103,N_15551,N_15394);
or U16104 (N_16104,N_15995,N_15375);
xnor U16105 (N_16105,N_15446,N_15944);
and U16106 (N_16106,N_15738,N_15986);
and U16107 (N_16107,N_15270,N_15390);
nor U16108 (N_16108,N_15686,N_15792);
or U16109 (N_16109,N_15259,N_15907);
or U16110 (N_16110,N_15604,N_15455);
or U16111 (N_16111,N_15256,N_15520);
nor U16112 (N_16112,N_15585,N_15212);
and U16113 (N_16113,N_15244,N_15860);
nor U16114 (N_16114,N_15303,N_15880);
or U16115 (N_16115,N_15985,N_15257);
or U16116 (N_16116,N_15466,N_15889);
nand U16117 (N_16117,N_15068,N_15024);
nand U16118 (N_16118,N_15278,N_15385);
nand U16119 (N_16119,N_15090,N_15022);
and U16120 (N_16120,N_15138,N_15871);
or U16121 (N_16121,N_15373,N_15432);
nor U16122 (N_16122,N_15412,N_15714);
xor U16123 (N_16123,N_15430,N_15900);
and U16124 (N_16124,N_15940,N_15688);
nand U16125 (N_16125,N_15340,N_15252);
nor U16126 (N_16126,N_15467,N_15049);
nand U16127 (N_16127,N_15083,N_15306);
or U16128 (N_16128,N_15184,N_15673);
and U16129 (N_16129,N_15531,N_15700);
nand U16130 (N_16130,N_15822,N_15052);
nand U16131 (N_16131,N_15421,N_15471);
and U16132 (N_16132,N_15496,N_15921);
nor U16133 (N_16133,N_15050,N_15070);
nor U16134 (N_16134,N_15517,N_15012);
or U16135 (N_16135,N_15107,N_15590);
nand U16136 (N_16136,N_15961,N_15560);
and U16137 (N_16137,N_15844,N_15169);
and U16138 (N_16138,N_15849,N_15843);
xor U16139 (N_16139,N_15565,N_15209);
xor U16140 (N_16140,N_15145,N_15788);
nand U16141 (N_16141,N_15178,N_15727);
and U16142 (N_16142,N_15267,N_15662);
xor U16143 (N_16143,N_15233,N_15170);
xor U16144 (N_16144,N_15349,N_15489);
and U16145 (N_16145,N_15003,N_15745);
or U16146 (N_16146,N_15747,N_15222);
xor U16147 (N_16147,N_15776,N_15440);
nand U16148 (N_16148,N_15847,N_15073);
nor U16149 (N_16149,N_15563,N_15854);
or U16150 (N_16150,N_15798,N_15619);
and U16151 (N_16151,N_15901,N_15216);
nor U16152 (N_16152,N_15371,N_15000);
xor U16153 (N_16153,N_15291,N_15609);
nand U16154 (N_16154,N_15869,N_15758);
xor U16155 (N_16155,N_15800,N_15229);
xor U16156 (N_16156,N_15397,N_15797);
or U16157 (N_16157,N_15884,N_15314);
nor U16158 (N_16158,N_15383,N_15182);
xnor U16159 (N_16159,N_15028,N_15633);
and U16160 (N_16160,N_15875,N_15930);
and U16161 (N_16161,N_15890,N_15981);
nor U16162 (N_16162,N_15649,N_15891);
and U16163 (N_16163,N_15469,N_15396);
nor U16164 (N_16164,N_15147,N_15909);
xnor U16165 (N_16165,N_15650,N_15290);
or U16166 (N_16166,N_15634,N_15828);
nand U16167 (N_16167,N_15555,N_15861);
nand U16168 (N_16168,N_15393,N_15239);
nand U16169 (N_16169,N_15803,N_15321);
nand U16170 (N_16170,N_15805,N_15832);
and U16171 (N_16171,N_15559,N_15666);
nand U16172 (N_16172,N_15238,N_15338);
and U16173 (N_16173,N_15220,N_15279);
xnor U16174 (N_16174,N_15942,N_15841);
and U16175 (N_16175,N_15487,N_15451);
and U16176 (N_16176,N_15151,N_15928);
and U16177 (N_16177,N_15401,N_15643);
nand U16178 (N_16178,N_15499,N_15542);
nand U16179 (N_16179,N_15567,N_15039);
and U16180 (N_16180,N_15804,N_15872);
and U16181 (N_16181,N_15808,N_15576);
nor U16182 (N_16182,N_15718,N_15699);
xor U16183 (N_16183,N_15910,N_15164);
or U16184 (N_16184,N_15952,N_15288);
and U16185 (N_16185,N_15839,N_15179);
xor U16186 (N_16186,N_15165,N_15647);
and U16187 (N_16187,N_15475,N_15888);
and U16188 (N_16188,N_15286,N_15535);
and U16189 (N_16189,N_15484,N_15608);
or U16190 (N_16190,N_15297,N_15992);
nor U16191 (N_16191,N_15816,N_15998);
and U16192 (N_16192,N_15053,N_15631);
xnor U16193 (N_16193,N_15046,N_15825);
and U16194 (N_16194,N_15354,N_15262);
xnor U16195 (N_16195,N_15389,N_15304);
xor U16196 (N_16196,N_15645,N_15091);
and U16197 (N_16197,N_15809,N_15150);
and U16198 (N_16198,N_15284,N_15077);
nand U16199 (N_16199,N_15915,N_15336);
and U16200 (N_16200,N_15739,N_15020);
or U16201 (N_16201,N_15245,N_15902);
or U16202 (N_16202,N_15510,N_15006);
nor U16203 (N_16203,N_15051,N_15167);
nand U16204 (N_16204,N_15195,N_15675);
or U16205 (N_16205,N_15452,N_15410);
or U16206 (N_16206,N_15518,N_15971);
and U16207 (N_16207,N_15231,N_15348);
xnor U16208 (N_16208,N_15160,N_15364);
nand U16209 (N_16209,N_15065,N_15859);
or U16210 (N_16210,N_15476,N_15626);
nand U16211 (N_16211,N_15166,N_15681);
nor U16212 (N_16212,N_15557,N_15076);
xor U16213 (N_16213,N_15334,N_15918);
nor U16214 (N_16214,N_15554,N_15969);
and U16215 (N_16215,N_15523,N_15811);
nand U16216 (N_16216,N_15400,N_15128);
nor U16217 (N_16217,N_15269,N_15558);
nor U16218 (N_16218,N_15345,N_15180);
or U16219 (N_16219,N_15979,N_15795);
xnor U16220 (N_16220,N_15137,N_15356);
or U16221 (N_16221,N_15735,N_15602);
or U16222 (N_16222,N_15765,N_15703);
nand U16223 (N_16223,N_15204,N_15656);
nand U16224 (N_16224,N_15713,N_15759);
nand U16225 (N_16225,N_15337,N_15529);
and U16226 (N_16226,N_15949,N_15600);
nand U16227 (N_16227,N_15454,N_15913);
xor U16228 (N_16228,N_15524,N_15016);
xor U16229 (N_16229,N_15341,N_15857);
and U16230 (N_16230,N_15208,N_15034);
and U16231 (N_16231,N_15136,N_15246);
nand U16232 (N_16232,N_15584,N_15419);
or U16233 (N_16233,N_15895,N_15980);
nand U16234 (N_16234,N_15459,N_15434);
xor U16235 (N_16235,N_15597,N_15780);
nor U16236 (N_16236,N_15149,N_15358);
nand U16237 (N_16237,N_15866,N_15948);
nand U16238 (N_16238,N_15274,N_15021);
or U16239 (N_16239,N_15101,N_15506);
or U16240 (N_16240,N_15224,N_15105);
nand U16241 (N_16241,N_15723,N_15175);
and U16242 (N_16242,N_15155,N_15359);
nor U16243 (N_16243,N_15970,N_15785);
nand U16244 (N_16244,N_15102,N_15532);
or U16245 (N_16245,N_15990,N_15912);
xnor U16246 (N_16246,N_15386,N_15852);
nor U16247 (N_16247,N_15708,N_15855);
and U16248 (N_16248,N_15381,N_15351);
or U16249 (N_16249,N_15993,N_15539);
or U16250 (N_16250,N_15268,N_15646);
and U16251 (N_16251,N_15310,N_15867);
nand U16252 (N_16252,N_15118,N_15937);
and U16253 (N_16253,N_15541,N_15878);
and U16254 (N_16254,N_15058,N_15644);
or U16255 (N_16255,N_15943,N_15848);
nor U16256 (N_16256,N_15599,N_15579);
nand U16257 (N_16257,N_15094,N_15956);
and U16258 (N_16258,N_15292,N_15295);
or U16259 (N_16259,N_15573,N_15019);
nand U16260 (N_16260,N_15367,N_15716);
and U16261 (N_16261,N_15014,N_15574);
nand U16262 (N_16262,N_15740,N_15010);
or U16263 (N_16263,N_15527,N_15048);
xor U16264 (N_16264,N_15922,N_15468);
and U16265 (N_16265,N_15719,N_15362);
nand U16266 (N_16266,N_15936,N_15836);
xnor U16267 (N_16267,N_15181,N_15678);
or U16268 (N_16268,N_15479,N_15837);
nor U16269 (N_16269,N_15702,N_15734);
or U16270 (N_16270,N_15885,N_15380);
xor U16271 (N_16271,N_15997,N_15978);
xnor U16272 (N_16272,N_15187,N_15814);
or U16273 (N_16273,N_15472,N_15829);
or U16274 (N_16274,N_15422,N_15243);
nor U16275 (N_16275,N_15533,N_15865);
xor U16276 (N_16276,N_15121,N_15013);
nand U16277 (N_16277,N_15616,N_15553);
and U16278 (N_16278,N_15705,N_15540);
and U16279 (N_16279,N_15363,N_15655);
nor U16280 (N_16280,N_15113,N_15706);
or U16281 (N_16281,N_15858,N_15123);
and U16282 (N_16282,N_15342,N_15856);
or U16283 (N_16283,N_15508,N_15720);
and U16284 (N_16284,N_15406,N_15711);
nor U16285 (N_16285,N_15596,N_15728);
or U16286 (N_16286,N_15343,N_15679);
or U16287 (N_16287,N_15498,N_15810);
and U16288 (N_16288,N_15623,N_15173);
or U16289 (N_16289,N_15218,N_15934);
or U16290 (N_16290,N_15298,N_15690);
or U16291 (N_16291,N_15691,N_15654);
nor U16292 (N_16292,N_15924,N_15685);
and U16293 (N_16293,N_15762,N_15158);
nor U16294 (N_16294,N_15743,N_15975);
xnor U16295 (N_16295,N_15194,N_15486);
xor U16296 (N_16296,N_15462,N_15493);
and U16297 (N_16297,N_15125,N_15564);
nand U16298 (N_16298,N_15730,N_15032);
or U16299 (N_16299,N_15436,N_15089);
xnor U16300 (N_16300,N_15242,N_15437);
nand U16301 (N_16301,N_15618,N_15960);
and U16302 (N_16302,N_15941,N_15156);
and U16303 (N_16303,N_15546,N_15569);
nand U16304 (N_16304,N_15041,N_15823);
and U16305 (N_16305,N_15382,N_15793);
or U16306 (N_16306,N_15749,N_15606);
nand U16307 (N_16307,N_15287,N_15709);
nor U16308 (N_16308,N_15119,N_15333);
or U16309 (N_16309,N_15587,N_15272);
or U16310 (N_16310,N_15409,N_15568);
xor U16311 (N_16311,N_15729,N_15399);
and U16312 (N_16312,N_15697,N_15157);
nand U16313 (N_16313,N_15368,N_15096);
or U16314 (N_16314,N_15296,N_15586);
nor U16315 (N_16315,N_15931,N_15481);
xor U16316 (N_16316,N_15724,N_15172);
or U16317 (N_16317,N_15737,N_15752);
nor U16318 (N_16318,N_15495,N_15802);
nor U16319 (N_16319,N_15221,N_15098);
xnor U16320 (N_16320,N_15092,N_15898);
xor U16321 (N_16321,N_15612,N_15248);
xor U16322 (N_16322,N_15876,N_15513);
xor U16323 (N_16323,N_15974,N_15742);
nand U16324 (N_16324,N_15404,N_15084);
or U16325 (N_16325,N_15671,N_15117);
xnor U16326 (N_16326,N_15146,N_15171);
or U16327 (N_16327,N_15492,N_15522);
nand U16328 (N_16328,N_15899,N_15355);
nor U16329 (N_16329,N_15007,N_15370);
and U16330 (N_16330,N_15202,N_15544);
nand U16331 (N_16331,N_15701,N_15223);
xor U16332 (N_16332,N_15461,N_15733);
or U16333 (N_16333,N_15991,N_15120);
or U16334 (N_16334,N_15966,N_15778);
nand U16335 (N_16335,N_15460,N_15309);
or U16336 (N_16336,N_15769,N_15774);
nor U16337 (N_16337,N_15601,N_15651);
or U16338 (N_16338,N_15783,N_15879);
or U16339 (N_16339,N_15426,N_15457);
or U16340 (N_16340,N_15031,N_15441);
and U16341 (N_16341,N_15030,N_15632);
xor U16342 (N_16342,N_15503,N_15427);
xor U16343 (N_16343,N_15033,N_15131);
xnor U16344 (N_16344,N_15684,N_15906);
nand U16345 (N_16345,N_15372,N_15059);
and U16346 (N_16346,N_15330,N_15502);
nor U16347 (N_16347,N_15190,N_15080);
nor U16348 (N_16348,N_15622,N_15215);
nor U16349 (N_16349,N_15773,N_15116);
nand U16350 (N_16350,N_15689,N_15605);
nor U16351 (N_16351,N_15199,N_15721);
nand U16352 (N_16352,N_15444,N_15465);
nor U16353 (N_16353,N_15549,N_15148);
or U16354 (N_16354,N_15488,N_15192);
nor U16355 (N_16355,N_15617,N_15905);
nand U16356 (N_16356,N_15234,N_15001);
nor U16357 (N_16357,N_15777,N_15477);
xor U16358 (N_16358,N_15074,N_15945);
and U16359 (N_16359,N_15110,N_15483);
or U16360 (N_16360,N_15300,N_15505);
nor U16361 (N_16361,N_15850,N_15853);
nor U16362 (N_16362,N_15868,N_15935);
nor U16363 (N_16363,N_15807,N_15712);
or U16364 (N_16364,N_15273,N_15806);
and U16365 (N_16365,N_15515,N_15683);
xnor U16366 (N_16366,N_15361,N_15135);
and U16367 (N_16367,N_15968,N_15817);
xnor U16368 (N_16368,N_15307,N_15347);
xor U16369 (N_16369,N_15226,N_15717);
nand U16370 (N_16370,N_15582,N_15093);
nor U16371 (N_16371,N_15322,N_15255);
xor U16372 (N_16372,N_15607,N_15668);
nor U16373 (N_16373,N_15755,N_15919);
and U16374 (N_16374,N_15413,N_15235);
and U16375 (N_16375,N_15819,N_15999);
xor U16376 (N_16376,N_15023,N_15026);
and U16377 (N_16377,N_15897,N_15528);
nand U16378 (N_16378,N_15514,N_15615);
xnor U16379 (N_16379,N_15217,N_15610);
or U16380 (N_16380,N_15732,N_15060);
nor U16381 (N_16381,N_15562,N_15638);
nand U16382 (N_16382,N_15435,N_15693);
nand U16383 (N_16383,N_15159,N_15530);
nand U16384 (N_16384,N_15911,N_15056);
xor U16385 (N_16385,N_15133,N_15659);
xor U16386 (N_16386,N_15750,N_15967);
xnor U16387 (N_16387,N_15620,N_15251);
xor U16388 (N_16388,N_15236,N_15715);
nor U16389 (N_16389,N_15763,N_15726);
nand U16390 (N_16390,N_15550,N_15478);
nor U16391 (N_16391,N_15230,N_15751);
and U16392 (N_16392,N_15920,N_15042);
xor U16393 (N_16393,N_15501,N_15054);
and U16394 (N_16394,N_15965,N_15826);
or U16395 (N_16395,N_15015,N_15674);
xor U16396 (N_16396,N_15253,N_15219);
xnor U16397 (N_16397,N_15140,N_15197);
and U16398 (N_16398,N_15748,N_15772);
or U16399 (N_16399,N_15142,N_15200);
nor U16400 (N_16400,N_15830,N_15725);
and U16401 (N_16401,N_15640,N_15534);
or U16402 (N_16402,N_15002,N_15916);
or U16403 (N_16403,N_15627,N_15285);
and U16404 (N_16404,N_15661,N_15198);
nand U16405 (N_16405,N_15538,N_15443);
xor U16406 (N_16406,N_15005,N_15417);
xor U16407 (N_16407,N_15537,N_15439);
nand U16408 (N_16408,N_15815,N_15873);
xnor U16409 (N_16409,N_15081,N_15784);
xor U16410 (N_16410,N_15588,N_15746);
xnor U16411 (N_16411,N_15566,N_15144);
or U16412 (N_16412,N_15211,N_15188);
xor U16413 (N_16413,N_15621,N_15473);
xor U16414 (N_16414,N_15692,N_15570);
nor U16415 (N_16415,N_15317,N_15191);
nand U16416 (N_16416,N_15500,N_15326);
nand U16417 (N_16417,N_15339,N_15572);
nor U16418 (N_16418,N_15329,N_15917);
nor U16419 (N_16419,N_15504,N_15183);
nor U16420 (N_16420,N_15594,N_15526);
and U16421 (N_16421,N_15127,N_15925);
xor U16422 (N_16422,N_15293,N_15378);
xnor U16423 (N_16423,N_15680,N_15629);
xor U16424 (N_16424,N_15521,N_15958);
xor U16425 (N_16425,N_15982,N_15894);
nor U16426 (N_16426,N_15794,N_15474);
nor U16427 (N_16427,N_15414,N_15027);
and U16428 (N_16428,N_15770,N_15407);
or U16429 (N_16429,N_15877,N_15756);
nor U16430 (N_16430,N_15818,N_15741);
xor U16431 (N_16431,N_15485,N_15240);
xor U16432 (N_16432,N_15938,N_15099);
xor U16433 (N_16433,N_15442,N_15152);
and U16434 (N_16434,N_15983,N_15280);
nor U16435 (N_16435,N_15753,N_15332);
nor U16436 (N_16436,N_15497,N_15927);
or U16437 (N_16437,N_15658,N_15408);
or U16438 (N_16438,N_15831,N_15423);
xnor U16439 (N_16439,N_15360,N_15210);
or U16440 (N_16440,N_15663,N_15132);
and U16441 (N_16441,N_15571,N_15575);
nand U16442 (N_16442,N_15018,N_15491);
or U16443 (N_16443,N_15353,N_15324);
nand U16444 (N_16444,N_15078,N_15722);
xor U16445 (N_16445,N_15470,N_15064);
nand U16446 (N_16446,N_15984,N_15227);
nor U16447 (N_16447,N_15425,N_15547);
or U16448 (N_16448,N_15311,N_15939);
xnor U16449 (N_16449,N_15796,N_15398);
or U16450 (N_16450,N_15864,N_15543);
and U16451 (N_16451,N_15228,N_15953);
xnor U16452 (N_16452,N_15827,N_15963);
or U16453 (N_16453,N_15881,N_15698);
xnor U16454 (N_16454,N_15914,N_15040);
nor U16455 (N_16455,N_15813,N_15624);
nand U16456 (N_16456,N_15694,N_15294);
or U16457 (N_16457,N_15896,N_15011);
or U16458 (N_16458,N_15335,N_15447);
and U16459 (N_16459,N_15377,N_15833);
or U16460 (N_16460,N_15821,N_15266);
nand U16461 (N_16461,N_15450,N_15395);
or U16462 (N_16462,N_15592,N_15047);
nor U16463 (N_16463,N_15008,N_15665);
xnor U16464 (N_16464,N_15642,N_15189);
nor U16465 (N_16465,N_15154,N_15962);
xnor U16466 (N_16466,N_15736,N_15892);
nand U16467 (N_16467,N_15062,N_15611);
or U16468 (N_16468,N_15344,N_15036);
xor U16469 (N_16469,N_15761,N_15652);
nor U16470 (N_16470,N_15275,N_15043);
or U16471 (N_16471,N_15628,N_15820);
or U16472 (N_16472,N_15874,N_15438);
nor U16473 (N_16473,N_15653,N_15352);
nand U16474 (N_16474,N_15957,N_15614);
nand U16475 (N_16475,N_15420,N_15176);
and U16476 (N_16476,N_15082,N_15786);
and U16477 (N_16477,N_15581,N_15842);
nor U16478 (N_16478,N_15388,N_15480);
nand U16479 (N_16479,N_15768,N_15886);
nor U16480 (N_16480,N_15445,N_15241);
nand U16481 (N_16481,N_15791,N_15932);
xnor U16482 (N_16482,N_15882,N_15044);
nand U16483 (N_16483,N_15790,N_15552);
nor U16484 (N_16484,N_15325,N_15206);
or U16485 (N_16485,N_15760,N_15254);
or U16486 (N_16486,N_15104,N_15580);
nor U16487 (N_16487,N_15577,N_15346);
nand U16488 (N_16488,N_15657,N_15095);
xor U16489 (N_16489,N_15583,N_15507);
xor U16490 (N_16490,N_15232,N_15185);
nand U16491 (N_16491,N_15009,N_15779);
nand U16492 (N_16492,N_15376,N_15923);
and U16493 (N_16493,N_15840,N_15433);
xnor U16494 (N_16494,N_15100,N_15061);
and U16495 (N_16495,N_15207,N_15072);
xnor U16496 (N_16496,N_15883,N_15835);
or U16497 (N_16497,N_15677,N_15143);
or U16498 (N_16498,N_15055,N_15038);
nor U16499 (N_16499,N_15903,N_15775);
xor U16500 (N_16500,N_15076,N_15294);
or U16501 (N_16501,N_15577,N_15006);
or U16502 (N_16502,N_15560,N_15780);
and U16503 (N_16503,N_15509,N_15080);
or U16504 (N_16504,N_15865,N_15919);
nand U16505 (N_16505,N_15309,N_15199);
xnor U16506 (N_16506,N_15067,N_15755);
or U16507 (N_16507,N_15639,N_15626);
xor U16508 (N_16508,N_15192,N_15117);
nand U16509 (N_16509,N_15220,N_15243);
or U16510 (N_16510,N_15088,N_15799);
nor U16511 (N_16511,N_15084,N_15758);
xnor U16512 (N_16512,N_15364,N_15833);
or U16513 (N_16513,N_15115,N_15310);
xor U16514 (N_16514,N_15448,N_15462);
or U16515 (N_16515,N_15524,N_15896);
xor U16516 (N_16516,N_15203,N_15051);
xnor U16517 (N_16517,N_15061,N_15024);
nand U16518 (N_16518,N_15761,N_15534);
and U16519 (N_16519,N_15516,N_15940);
nand U16520 (N_16520,N_15055,N_15962);
nor U16521 (N_16521,N_15143,N_15303);
nor U16522 (N_16522,N_15827,N_15941);
nand U16523 (N_16523,N_15436,N_15327);
or U16524 (N_16524,N_15475,N_15351);
nand U16525 (N_16525,N_15803,N_15566);
and U16526 (N_16526,N_15590,N_15885);
nand U16527 (N_16527,N_15276,N_15531);
xor U16528 (N_16528,N_15320,N_15202);
and U16529 (N_16529,N_15567,N_15468);
xor U16530 (N_16530,N_15846,N_15732);
or U16531 (N_16531,N_15075,N_15114);
and U16532 (N_16532,N_15374,N_15808);
nor U16533 (N_16533,N_15634,N_15618);
and U16534 (N_16534,N_15295,N_15652);
nor U16535 (N_16535,N_15027,N_15403);
xor U16536 (N_16536,N_15252,N_15139);
nor U16537 (N_16537,N_15366,N_15485);
or U16538 (N_16538,N_15214,N_15292);
nor U16539 (N_16539,N_15172,N_15573);
and U16540 (N_16540,N_15423,N_15364);
nor U16541 (N_16541,N_15901,N_15700);
and U16542 (N_16542,N_15236,N_15530);
and U16543 (N_16543,N_15168,N_15206);
nor U16544 (N_16544,N_15691,N_15299);
nand U16545 (N_16545,N_15550,N_15646);
xnor U16546 (N_16546,N_15319,N_15523);
nor U16547 (N_16547,N_15742,N_15795);
nor U16548 (N_16548,N_15108,N_15322);
nand U16549 (N_16549,N_15536,N_15035);
and U16550 (N_16550,N_15286,N_15563);
xnor U16551 (N_16551,N_15317,N_15646);
nand U16552 (N_16552,N_15423,N_15001);
and U16553 (N_16553,N_15813,N_15896);
or U16554 (N_16554,N_15164,N_15669);
nor U16555 (N_16555,N_15392,N_15399);
nand U16556 (N_16556,N_15368,N_15753);
nor U16557 (N_16557,N_15363,N_15108);
xor U16558 (N_16558,N_15389,N_15615);
and U16559 (N_16559,N_15216,N_15855);
xor U16560 (N_16560,N_15110,N_15541);
xnor U16561 (N_16561,N_15404,N_15164);
nand U16562 (N_16562,N_15061,N_15481);
nand U16563 (N_16563,N_15119,N_15011);
xnor U16564 (N_16564,N_15984,N_15423);
xor U16565 (N_16565,N_15734,N_15784);
nor U16566 (N_16566,N_15594,N_15404);
nand U16567 (N_16567,N_15518,N_15881);
nand U16568 (N_16568,N_15533,N_15171);
nor U16569 (N_16569,N_15760,N_15580);
and U16570 (N_16570,N_15894,N_15200);
nand U16571 (N_16571,N_15297,N_15399);
nor U16572 (N_16572,N_15036,N_15177);
nor U16573 (N_16573,N_15359,N_15067);
nand U16574 (N_16574,N_15627,N_15976);
nor U16575 (N_16575,N_15791,N_15250);
or U16576 (N_16576,N_15098,N_15366);
xnor U16577 (N_16577,N_15039,N_15696);
nand U16578 (N_16578,N_15194,N_15401);
or U16579 (N_16579,N_15754,N_15272);
and U16580 (N_16580,N_15563,N_15500);
nor U16581 (N_16581,N_15267,N_15551);
and U16582 (N_16582,N_15695,N_15431);
and U16583 (N_16583,N_15659,N_15739);
and U16584 (N_16584,N_15844,N_15032);
nand U16585 (N_16585,N_15343,N_15233);
nor U16586 (N_16586,N_15264,N_15710);
xor U16587 (N_16587,N_15126,N_15879);
xnor U16588 (N_16588,N_15919,N_15720);
or U16589 (N_16589,N_15743,N_15418);
nand U16590 (N_16590,N_15983,N_15706);
nor U16591 (N_16591,N_15383,N_15308);
nor U16592 (N_16592,N_15391,N_15170);
or U16593 (N_16593,N_15309,N_15202);
or U16594 (N_16594,N_15820,N_15640);
xor U16595 (N_16595,N_15479,N_15310);
nor U16596 (N_16596,N_15581,N_15963);
nor U16597 (N_16597,N_15362,N_15136);
and U16598 (N_16598,N_15124,N_15847);
nor U16599 (N_16599,N_15915,N_15306);
nor U16600 (N_16600,N_15567,N_15398);
xnor U16601 (N_16601,N_15522,N_15239);
or U16602 (N_16602,N_15770,N_15506);
or U16603 (N_16603,N_15619,N_15014);
or U16604 (N_16604,N_15918,N_15902);
and U16605 (N_16605,N_15312,N_15240);
or U16606 (N_16606,N_15386,N_15612);
nand U16607 (N_16607,N_15449,N_15018);
and U16608 (N_16608,N_15849,N_15285);
xor U16609 (N_16609,N_15282,N_15921);
nor U16610 (N_16610,N_15439,N_15675);
xnor U16611 (N_16611,N_15773,N_15506);
or U16612 (N_16612,N_15015,N_15478);
and U16613 (N_16613,N_15092,N_15957);
nor U16614 (N_16614,N_15816,N_15474);
or U16615 (N_16615,N_15398,N_15562);
nand U16616 (N_16616,N_15863,N_15455);
and U16617 (N_16617,N_15846,N_15539);
xnor U16618 (N_16618,N_15620,N_15500);
xor U16619 (N_16619,N_15474,N_15434);
and U16620 (N_16620,N_15705,N_15299);
nor U16621 (N_16621,N_15541,N_15473);
or U16622 (N_16622,N_15539,N_15494);
or U16623 (N_16623,N_15446,N_15565);
or U16624 (N_16624,N_15707,N_15799);
and U16625 (N_16625,N_15043,N_15185);
or U16626 (N_16626,N_15688,N_15564);
nor U16627 (N_16627,N_15183,N_15676);
xnor U16628 (N_16628,N_15288,N_15354);
and U16629 (N_16629,N_15578,N_15609);
nand U16630 (N_16630,N_15556,N_15116);
and U16631 (N_16631,N_15058,N_15118);
nand U16632 (N_16632,N_15331,N_15696);
nor U16633 (N_16633,N_15047,N_15254);
or U16634 (N_16634,N_15635,N_15907);
xor U16635 (N_16635,N_15201,N_15841);
or U16636 (N_16636,N_15242,N_15557);
nand U16637 (N_16637,N_15690,N_15753);
xnor U16638 (N_16638,N_15297,N_15777);
nor U16639 (N_16639,N_15860,N_15686);
nor U16640 (N_16640,N_15033,N_15970);
nand U16641 (N_16641,N_15997,N_15550);
xor U16642 (N_16642,N_15890,N_15191);
xnor U16643 (N_16643,N_15584,N_15155);
or U16644 (N_16644,N_15659,N_15629);
and U16645 (N_16645,N_15132,N_15231);
xor U16646 (N_16646,N_15650,N_15407);
nand U16647 (N_16647,N_15009,N_15474);
nor U16648 (N_16648,N_15251,N_15501);
or U16649 (N_16649,N_15609,N_15614);
xor U16650 (N_16650,N_15301,N_15437);
or U16651 (N_16651,N_15130,N_15485);
and U16652 (N_16652,N_15768,N_15795);
nor U16653 (N_16653,N_15705,N_15290);
or U16654 (N_16654,N_15780,N_15156);
xor U16655 (N_16655,N_15023,N_15471);
nand U16656 (N_16656,N_15234,N_15566);
and U16657 (N_16657,N_15994,N_15159);
nand U16658 (N_16658,N_15609,N_15606);
nor U16659 (N_16659,N_15812,N_15889);
xnor U16660 (N_16660,N_15323,N_15906);
xor U16661 (N_16661,N_15345,N_15428);
or U16662 (N_16662,N_15232,N_15680);
xor U16663 (N_16663,N_15683,N_15843);
xor U16664 (N_16664,N_15730,N_15333);
xor U16665 (N_16665,N_15472,N_15657);
and U16666 (N_16666,N_15660,N_15059);
xnor U16667 (N_16667,N_15883,N_15230);
xnor U16668 (N_16668,N_15928,N_15118);
nand U16669 (N_16669,N_15668,N_15985);
and U16670 (N_16670,N_15621,N_15845);
xnor U16671 (N_16671,N_15217,N_15178);
xor U16672 (N_16672,N_15924,N_15848);
nor U16673 (N_16673,N_15526,N_15697);
nor U16674 (N_16674,N_15520,N_15684);
xnor U16675 (N_16675,N_15040,N_15362);
nand U16676 (N_16676,N_15981,N_15993);
xnor U16677 (N_16677,N_15173,N_15066);
and U16678 (N_16678,N_15163,N_15107);
xor U16679 (N_16679,N_15552,N_15855);
or U16680 (N_16680,N_15413,N_15988);
nand U16681 (N_16681,N_15071,N_15634);
or U16682 (N_16682,N_15556,N_15457);
nand U16683 (N_16683,N_15019,N_15580);
nor U16684 (N_16684,N_15319,N_15055);
or U16685 (N_16685,N_15504,N_15367);
nor U16686 (N_16686,N_15659,N_15380);
and U16687 (N_16687,N_15612,N_15814);
and U16688 (N_16688,N_15857,N_15521);
xor U16689 (N_16689,N_15492,N_15796);
xor U16690 (N_16690,N_15586,N_15891);
nand U16691 (N_16691,N_15795,N_15864);
xor U16692 (N_16692,N_15187,N_15951);
or U16693 (N_16693,N_15856,N_15023);
nand U16694 (N_16694,N_15581,N_15914);
nor U16695 (N_16695,N_15949,N_15314);
nand U16696 (N_16696,N_15147,N_15385);
nor U16697 (N_16697,N_15210,N_15743);
nand U16698 (N_16698,N_15579,N_15231);
nor U16699 (N_16699,N_15483,N_15695);
and U16700 (N_16700,N_15816,N_15250);
nand U16701 (N_16701,N_15220,N_15842);
nor U16702 (N_16702,N_15949,N_15531);
xnor U16703 (N_16703,N_15079,N_15065);
or U16704 (N_16704,N_15657,N_15806);
nand U16705 (N_16705,N_15573,N_15239);
or U16706 (N_16706,N_15952,N_15292);
xnor U16707 (N_16707,N_15016,N_15876);
nor U16708 (N_16708,N_15467,N_15041);
or U16709 (N_16709,N_15173,N_15465);
and U16710 (N_16710,N_15485,N_15076);
nand U16711 (N_16711,N_15454,N_15250);
nand U16712 (N_16712,N_15666,N_15121);
and U16713 (N_16713,N_15887,N_15162);
and U16714 (N_16714,N_15286,N_15192);
or U16715 (N_16715,N_15334,N_15633);
nor U16716 (N_16716,N_15399,N_15548);
and U16717 (N_16717,N_15871,N_15592);
xnor U16718 (N_16718,N_15634,N_15970);
nand U16719 (N_16719,N_15953,N_15281);
nor U16720 (N_16720,N_15932,N_15216);
and U16721 (N_16721,N_15513,N_15763);
and U16722 (N_16722,N_15848,N_15979);
xnor U16723 (N_16723,N_15438,N_15887);
nor U16724 (N_16724,N_15628,N_15294);
or U16725 (N_16725,N_15643,N_15601);
nor U16726 (N_16726,N_15517,N_15472);
or U16727 (N_16727,N_15746,N_15743);
or U16728 (N_16728,N_15598,N_15456);
nand U16729 (N_16729,N_15515,N_15579);
nor U16730 (N_16730,N_15317,N_15909);
nand U16731 (N_16731,N_15093,N_15308);
or U16732 (N_16732,N_15876,N_15624);
nand U16733 (N_16733,N_15843,N_15466);
or U16734 (N_16734,N_15719,N_15777);
and U16735 (N_16735,N_15742,N_15233);
or U16736 (N_16736,N_15660,N_15263);
xor U16737 (N_16737,N_15373,N_15151);
or U16738 (N_16738,N_15571,N_15357);
and U16739 (N_16739,N_15758,N_15766);
and U16740 (N_16740,N_15050,N_15584);
nor U16741 (N_16741,N_15699,N_15126);
or U16742 (N_16742,N_15745,N_15877);
nor U16743 (N_16743,N_15317,N_15648);
and U16744 (N_16744,N_15026,N_15899);
nor U16745 (N_16745,N_15545,N_15664);
and U16746 (N_16746,N_15541,N_15332);
nand U16747 (N_16747,N_15143,N_15500);
xor U16748 (N_16748,N_15565,N_15004);
xor U16749 (N_16749,N_15941,N_15678);
nand U16750 (N_16750,N_15240,N_15430);
or U16751 (N_16751,N_15278,N_15395);
or U16752 (N_16752,N_15306,N_15226);
nand U16753 (N_16753,N_15530,N_15770);
xnor U16754 (N_16754,N_15104,N_15678);
nand U16755 (N_16755,N_15297,N_15778);
nor U16756 (N_16756,N_15436,N_15354);
nor U16757 (N_16757,N_15910,N_15833);
xor U16758 (N_16758,N_15961,N_15297);
xor U16759 (N_16759,N_15320,N_15570);
or U16760 (N_16760,N_15476,N_15733);
xor U16761 (N_16761,N_15846,N_15026);
nor U16762 (N_16762,N_15501,N_15326);
or U16763 (N_16763,N_15271,N_15369);
nand U16764 (N_16764,N_15373,N_15559);
nor U16765 (N_16765,N_15085,N_15052);
and U16766 (N_16766,N_15625,N_15985);
and U16767 (N_16767,N_15870,N_15445);
nand U16768 (N_16768,N_15680,N_15697);
xor U16769 (N_16769,N_15450,N_15754);
and U16770 (N_16770,N_15613,N_15907);
nand U16771 (N_16771,N_15843,N_15829);
nor U16772 (N_16772,N_15808,N_15326);
or U16773 (N_16773,N_15045,N_15552);
or U16774 (N_16774,N_15352,N_15211);
nor U16775 (N_16775,N_15515,N_15932);
nor U16776 (N_16776,N_15397,N_15284);
and U16777 (N_16777,N_15247,N_15604);
and U16778 (N_16778,N_15051,N_15665);
nor U16779 (N_16779,N_15066,N_15156);
and U16780 (N_16780,N_15171,N_15697);
nor U16781 (N_16781,N_15927,N_15590);
xnor U16782 (N_16782,N_15544,N_15473);
and U16783 (N_16783,N_15431,N_15261);
nor U16784 (N_16784,N_15581,N_15009);
and U16785 (N_16785,N_15906,N_15282);
and U16786 (N_16786,N_15762,N_15498);
xnor U16787 (N_16787,N_15153,N_15606);
or U16788 (N_16788,N_15317,N_15717);
or U16789 (N_16789,N_15660,N_15443);
xnor U16790 (N_16790,N_15788,N_15797);
nor U16791 (N_16791,N_15264,N_15385);
xnor U16792 (N_16792,N_15322,N_15623);
or U16793 (N_16793,N_15918,N_15372);
nor U16794 (N_16794,N_15732,N_15811);
nor U16795 (N_16795,N_15967,N_15056);
nor U16796 (N_16796,N_15081,N_15496);
nor U16797 (N_16797,N_15545,N_15059);
or U16798 (N_16798,N_15917,N_15029);
and U16799 (N_16799,N_15660,N_15296);
and U16800 (N_16800,N_15575,N_15417);
and U16801 (N_16801,N_15633,N_15394);
nor U16802 (N_16802,N_15106,N_15267);
and U16803 (N_16803,N_15743,N_15569);
xor U16804 (N_16804,N_15262,N_15050);
or U16805 (N_16805,N_15570,N_15554);
nor U16806 (N_16806,N_15357,N_15781);
or U16807 (N_16807,N_15043,N_15755);
and U16808 (N_16808,N_15173,N_15120);
or U16809 (N_16809,N_15939,N_15199);
or U16810 (N_16810,N_15952,N_15302);
or U16811 (N_16811,N_15783,N_15420);
nor U16812 (N_16812,N_15852,N_15128);
and U16813 (N_16813,N_15621,N_15671);
nand U16814 (N_16814,N_15295,N_15659);
and U16815 (N_16815,N_15093,N_15432);
nor U16816 (N_16816,N_15210,N_15145);
xor U16817 (N_16817,N_15548,N_15231);
xnor U16818 (N_16818,N_15473,N_15894);
xnor U16819 (N_16819,N_15457,N_15327);
and U16820 (N_16820,N_15173,N_15477);
or U16821 (N_16821,N_15398,N_15054);
or U16822 (N_16822,N_15108,N_15686);
nor U16823 (N_16823,N_15772,N_15684);
nor U16824 (N_16824,N_15458,N_15965);
xor U16825 (N_16825,N_15559,N_15633);
nand U16826 (N_16826,N_15295,N_15343);
and U16827 (N_16827,N_15614,N_15753);
or U16828 (N_16828,N_15652,N_15518);
or U16829 (N_16829,N_15307,N_15495);
nand U16830 (N_16830,N_15608,N_15923);
and U16831 (N_16831,N_15173,N_15621);
and U16832 (N_16832,N_15183,N_15895);
or U16833 (N_16833,N_15519,N_15723);
nor U16834 (N_16834,N_15405,N_15841);
nor U16835 (N_16835,N_15291,N_15522);
xnor U16836 (N_16836,N_15005,N_15625);
and U16837 (N_16837,N_15469,N_15058);
xnor U16838 (N_16838,N_15715,N_15810);
nor U16839 (N_16839,N_15652,N_15204);
and U16840 (N_16840,N_15975,N_15733);
or U16841 (N_16841,N_15963,N_15762);
xor U16842 (N_16842,N_15660,N_15389);
or U16843 (N_16843,N_15215,N_15558);
or U16844 (N_16844,N_15715,N_15107);
xor U16845 (N_16845,N_15491,N_15926);
nand U16846 (N_16846,N_15656,N_15894);
nand U16847 (N_16847,N_15712,N_15197);
and U16848 (N_16848,N_15652,N_15777);
or U16849 (N_16849,N_15191,N_15257);
xnor U16850 (N_16850,N_15202,N_15847);
or U16851 (N_16851,N_15100,N_15908);
xor U16852 (N_16852,N_15318,N_15502);
nor U16853 (N_16853,N_15938,N_15717);
xor U16854 (N_16854,N_15460,N_15663);
nor U16855 (N_16855,N_15257,N_15045);
xor U16856 (N_16856,N_15559,N_15813);
and U16857 (N_16857,N_15833,N_15231);
or U16858 (N_16858,N_15810,N_15448);
xnor U16859 (N_16859,N_15983,N_15772);
xnor U16860 (N_16860,N_15121,N_15863);
and U16861 (N_16861,N_15857,N_15692);
or U16862 (N_16862,N_15443,N_15220);
nor U16863 (N_16863,N_15645,N_15014);
nor U16864 (N_16864,N_15643,N_15388);
nand U16865 (N_16865,N_15419,N_15224);
and U16866 (N_16866,N_15998,N_15358);
xnor U16867 (N_16867,N_15403,N_15656);
or U16868 (N_16868,N_15052,N_15634);
xor U16869 (N_16869,N_15032,N_15153);
nand U16870 (N_16870,N_15512,N_15441);
or U16871 (N_16871,N_15987,N_15973);
and U16872 (N_16872,N_15711,N_15996);
xor U16873 (N_16873,N_15150,N_15671);
and U16874 (N_16874,N_15944,N_15074);
or U16875 (N_16875,N_15464,N_15813);
nand U16876 (N_16876,N_15215,N_15098);
nor U16877 (N_16877,N_15965,N_15753);
or U16878 (N_16878,N_15178,N_15002);
or U16879 (N_16879,N_15888,N_15436);
nand U16880 (N_16880,N_15766,N_15010);
or U16881 (N_16881,N_15854,N_15574);
nor U16882 (N_16882,N_15045,N_15927);
and U16883 (N_16883,N_15947,N_15663);
nor U16884 (N_16884,N_15711,N_15623);
xnor U16885 (N_16885,N_15536,N_15838);
xnor U16886 (N_16886,N_15786,N_15460);
nand U16887 (N_16887,N_15377,N_15463);
or U16888 (N_16888,N_15637,N_15769);
nand U16889 (N_16889,N_15082,N_15566);
or U16890 (N_16890,N_15842,N_15469);
nand U16891 (N_16891,N_15664,N_15266);
xnor U16892 (N_16892,N_15543,N_15897);
xnor U16893 (N_16893,N_15659,N_15837);
nor U16894 (N_16894,N_15737,N_15720);
xnor U16895 (N_16895,N_15408,N_15381);
nor U16896 (N_16896,N_15921,N_15393);
xor U16897 (N_16897,N_15260,N_15233);
xnor U16898 (N_16898,N_15042,N_15417);
nand U16899 (N_16899,N_15453,N_15602);
or U16900 (N_16900,N_15939,N_15913);
or U16901 (N_16901,N_15302,N_15282);
and U16902 (N_16902,N_15025,N_15423);
or U16903 (N_16903,N_15830,N_15912);
and U16904 (N_16904,N_15665,N_15502);
nand U16905 (N_16905,N_15128,N_15058);
or U16906 (N_16906,N_15109,N_15294);
nor U16907 (N_16907,N_15569,N_15852);
and U16908 (N_16908,N_15338,N_15168);
nand U16909 (N_16909,N_15065,N_15087);
nand U16910 (N_16910,N_15360,N_15803);
and U16911 (N_16911,N_15866,N_15830);
or U16912 (N_16912,N_15105,N_15823);
nor U16913 (N_16913,N_15732,N_15441);
xor U16914 (N_16914,N_15510,N_15644);
and U16915 (N_16915,N_15296,N_15939);
nand U16916 (N_16916,N_15622,N_15913);
or U16917 (N_16917,N_15214,N_15007);
nand U16918 (N_16918,N_15114,N_15673);
or U16919 (N_16919,N_15914,N_15686);
nand U16920 (N_16920,N_15835,N_15804);
and U16921 (N_16921,N_15769,N_15827);
nand U16922 (N_16922,N_15328,N_15428);
or U16923 (N_16923,N_15032,N_15192);
or U16924 (N_16924,N_15060,N_15441);
xnor U16925 (N_16925,N_15495,N_15102);
nand U16926 (N_16926,N_15889,N_15926);
nor U16927 (N_16927,N_15752,N_15642);
nand U16928 (N_16928,N_15824,N_15557);
and U16929 (N_16929,N_15907,N_15244);
or U16930 (N_16930,N_15599,N_15656);
nand U16931 (N_16931,N_15728,N_15003);
nor U16932 (N_16932,N_15289,N_15321);
or U16933 (N_16933,N_15502,N_15873);
nor U16934 (N_16934,N_15643,N_15605);
or U16935 (N_16935,N_15838,N_15687);
or U16936 (N_16936,N_15838,N_15591);
xnor U16937 (N_16937,N_15922,N_15039);
nand U16938 (N_16938,N_15433,N_15273);
nand U16939 (N_16939,N_15604,N_15605);
xor U16940 (N_16940,N_15129,N_15983);
nand U16941 (N_16941,N_15323,N_15183);
nand U16942 (N_16942,N_15491,N_15185);
nor U16943 (N_16943,N_15924,N_15306);
xnor U16944 (N_16944,N_15021,N_15369);
nor U16945 (N_16945,N_15478,N_15928);
nand U16946 (N_16946,N_15676,N_15941);
nor U16947 (N_16947,N_15113,N_15606);
nand U16948 (N_16948,N_15978,N_15444);
nor U16949 (N_16949,N_15379,N_15812);
nor U16950 (N_16950,N_15307,N_15841);
nor U16951 (N_16951,N_15019,N_15017);
xor U16952 (N_16952,N_15463,N_15734);
or U16953 (N_16953,N_15467,N_15934);
and U16954 (N_16954,N_15093,N_15821);
or U16955 (N_16955,N_15035,N_15849);
nand U16956 (N_16956,N_15322,N_15366);
and U16957 (N_16957,N_15635,N_15570);
xor U16958 (N_16958,N_15861,N_15248);
and U16959 (N_16959,N_15212,N_15491);
nor U16960 (N_16960,N_15799,N_15514);
nor U16961 (N_16961,N_15616,N_15379);
nor U16962 (N_16962,N_15959,N_15831);
nor U16963 (N_16963,N_15267,N_15243);
nand U16964 (N_16964,N_15648,N_15362);
or U16965 (N_16965,N_15866,N_15664);
nand U16966 (N_16966,N_15307,N_15989);
nor U16967 (N_16967,N_15231,N_15519);
and U16968 (N_16968,N_15536,N_15948);
or U16969 (N_16969,N_15664,N_15239);
nand U16970 (N_16970,N_15955,N_15532);
nor U16971 (N_16971,N_15109,N_15805);
xnor U16972 (N_16972,N_15780,N_15988);
or U16973 (N_16973,N_15483,N_15894);
nor U16974 (N_16974,N_15568,N_15167);
nand U16975 (N_16975,N_15378,N_15905);
nor U16976 (N_16976,N_15821,N_15984);
nor U16977 (N_16977,N_15264,N_15261);
or U16978 (N_16978,N_15460,N_15502);
or U16979 (N_16979,N_15186,N_15132);
xor U16980 (N_16980,N_15191,N_15561);
xor U16981 (N_16981,N_15676,N_15665);
and U16982 (N_16982,N_15491,N_15213);
nor U16983 (N_16983,N_15256,N_15472);
and U16984 (N_16984,N_15694,N_15258);
and U16985 (N_16985,N_15153,N_15449);
and U16986 (N_16986,N_15195,N_15667);
or U16987 (N_16987,N_15614,N_15701);
nand U16988 (N_16988,N_15022,N_15360);
nor U16989 (N_16989,N_15416,N_15768);
or U16990 (N_16990,N_15815,N_15345);
or U16991 (N_16991,N_15082,N_15681);
or U16992 (N_16992,N_15367,N_15021);
and U16993 (N_16993,N_15455,N_15066);
xnor U16994 (N_16994,N_15162,N_15454);
nand U16995 (N_16995,N_15200,N_15306);
or U16996 (N_16996,N_15010,N_15909);
nor U16997 (N_16997,N_15911,N_15860);
or U16998 (N_16998,N_15733,N_15272);
and U16999 (N_16999,N_15859,N_15262);
nor U17000 (N_17000,N_16072,N_16595);
nor U17001 (N_17001,N_16321,N_16652);
nand U17002 (N_17002,N_16323,N_16913);
or U17003 (N_17003,N_16331,N_16443);
xnor U17004 (N_17004,N_16371,N_16144);
nand U17005 (N_17005,N_16713,N_16274);
or U17006 (N_17006,N_16971,N_16455);
nand U17007 (N_17007,N_16977,N_16644);
nor U17008 (N_17008,N_16044,N_16200);
or U17009 (N_17009,N_16918,N_16536);
nand U17010 (N_17010,N_16648,N_16880);
and U17011 (N_17011,N_16499,N_16119);
nor U17012 (N_17012,N_16877,N_16653);
nand U17013 (N_17013,N_16475,N_16764);
and U17014 (N_17014,N_16597,N_16706);
and U17015 (N_17015,N_16296,N_16839);
xnor U17016 (N_17016,N_16273,N_16821);
xnor U17017 (N_17017,N_16987,N_16288);
or U17018 (N_17018,N_16898,N_16926);
or U17019 (N_17019,N_16818,N_16613);
or U17020 (N_17020,N_16509,N_16389);
xnor U17021 (N_17021,N_16844,N_16832);
nand U17022 (N_17022,N_16013,N_16654);
and U17023 (N_17023,N_16493,N_16699);
and U17024 (N_17024,N_16248,N_16922);
xnor U17025 (N_17025,N_16451,N_16137);
or U17026 (N_17026,N_16481,N_16092);
nand U17027 (N_17027,N_16776,N_16978);
nor U17028 (N_17028,N_16082,N_16400);
nor U17029 (N_17029,N_16416,N_16546);
and U17030 (N_17030,N_16610,N_16523);
xor U17031 (N_17031,N_16322,N_16645);
nor U17032 (N_17032,N_16851,N_16552);
xor U17033 (N_17033,N_16736,N_16385);
nand U17034 (N_17034,N_16696,N_16008);
xnor U17035 (N_17035,N_16688,N_16808);
and U17036 (N_17036,N_16684,N_16030);
nand U17037 (N_17037,N_16533,N_16335);
and U17038 (N_17038,N_16143,N_16373);
nor U17039 (N_17039,N_16333,N_16437);
nand U17040 (N_17040,N_16570,N_16290);
xnor U17041 (N_17041,N_16716,N_16365);
or U17042 (N_17042,N_16332,N_16282);
or U17043 (N_17043,N_16802,N_16780);
or U17044 (N_17044,N_16297,N_16845);
xnor U17045 (N_17045,N_16559,N_16658);
nand U17046 (N_17046,N_16895,N_16228);
nor U17047 (N_17047,N_16305,N_16381);
nand U17048 (N_17048,N_16635,N_16853);
or U17049 (N_17049,N_16720,N_16916);
xor U17050 (N_17050,N_16584,N_16754);
nor U17051 (N_17051,N_16992,N_16530);
or U17052 (N_17052,N_16039,N_16002);
nor U17053 (N_17053,N_16842,N_16714);
or U17054 (N_17054,N_16370,N_16792);
nand U17055 (N_17055,N_16167,N_16677);
xor U17056 (N_17056,N_16545,N_16899);
nand U17057 (N_17057,N_16140,N_16760);
nand U17058 (N_17058,N_16099,N_16395);
nor U17059 (N_17059,N_16589,N_16594);
nand U17060 (N_17060,N_16567,N_16734);
xor U17061 (N_17061,N_16314,N_16446);
nor U17062 (N_17062,N_16420,N_16948);
xnor U17063 (N_17063,N_16958,N_16284);
nor U17064 (N_17064,N_16096,N_16988);
or U17065 (N_17065,N_16979,N_16620);
nor U17066 (N_17066,N_16689,N_16006);
and U17067 (N_17067,N_16937,N_16957);
xnor U17068 (N_17068,N_16369,N_16883);
and U17069 (N_17069,N_16797,N_16568);
xor U17070 (N_17070,N_16257,N_16266);
xnor U17071 (N_17071,N_16120,N_16291);
nor U17072 (N_17072,N_16307,N_16587);
nand U17073 (N_17073,N_16026,N_16772);
and U17074 (N_17074,N_16544,N_16703);
or U17075 (N_17075,N_16472,N_16383);
nand U17076 (N_17076,N_16474,N_16016);
or U17077 (N_17077,N_16878,N_16153);
xor U17078 (N_17078,N_16789,N_16555);
xnor U17079 (N_17079,N_16510,N_16516);
or U17080 (N_17080,N_16670,N_16833);
xor U17081 (N_17081,N_16168,N_16742);
and U17082 (N_17082,N_16207,N_16885);
nor U17083 (N_17083,N_16537,N_16040);
xor U17084 (N_17084,N_16513,N_16460);
xor U17085 (N_17085,N_16372,N_16521);
and U17086 (N_17086,N_16377,N_16005);
or U17087 (N_17087,N_16285,N_16969);
or U17088 (N_17088,N_16840,N_16114);
nand U17089 (N_17089,N_16019,N_16055);
xor U17090 (N_17090,N_16301,N_16686);
or U17091 (N_17091,N_16669,N_16512);
nand U17092 (N_17092,N_16866,N_16729);
xor U17093 (N_17093,N_16308,N_16449);
nand U17094 (N_17094,N_16339,N_16945);
and U17095 (N_17095,N_16286,N_16538);
or U17096 (N_17096,N_16352,N_16267);
or U17097 (N_17097,N_16965,N_16073);
and U17098 (N_17098,N_16439,N_16432);
xor U17099 (N_17099,N_16626,N_16127);
and U17100 (N_17100,N_16817,N_16132);
nor U17101 (N_17101,N_16747,N_16960);
or U17102 (N_17102,N_16912,N_16309);
and U17103 (N_17103,N_16972,N_16730);
or U17104 (N_17104,N_16025,N_16794);
xnor U17105 (N_17105,N_16611,N_16763);
xnor U17106 (N_17106,N_16588,N_16751);
or U17107 (N_17107,N_16678,N_16048);
nand U17108 (N_17108,N_16846,N_16075);
xor U17109 (N_17109,N_16453,N_16507);
nor U17110 (N_17110,N_16310,N_16262);
and U17111 (N_17111,N_16150,N_16094);
nor U17112 (N_17112,N_16024,N_16231);
nor U17113 (N_17113,N_16185,N_16638);
nor U17114 (N_17114,N_16955,N_16164);
nor U17115 (N_17115,N_16614,N_16906);
xnor U17116 (N_17116,N_16836,N_16175);
nor U17117 (N_17117,N_16116,N_16964);
xnor U17118 (N_17118,N_16664,N_16494);
nor U17119 (N_17119,N_16469,N_16596);
or U17120 (N_17120,N_16289,N_16236);
xor U17121 (N_17121,N_16190,N_16078);
nor U17122 (N_17122,N_16705,N_16911);
xor U17123 (N_17123,N_16542,N_16362);
xnor U17124 (N_17124,N_16483,N_16875);
nand U17125 (N_17125,N_16174,N_16146);
and U17126 (N_17126,N_16857,N_16725);
and U17127 (N_17127,N_16386,N_16962);
xnor U17128 (N_17128,N_16206,N_16525);
xnor U17129 (N_17129,N_16800,N_16612);
nor U17130 (N_17130,N_16023,N_16709);
nand U17131 (N_17131,N_16738,N_16882);
and U17132 (N_17132,N_16179,N_16886);
and U17133 (N_17133,N_16995,N_16276);
nand U17134 (N_17134,N_16178,N_16388);
nand U17135 (N_17135,N_16884,N_16104);
nand U17136 (N_17136,N_16828,N_16038);
nor U17137 (N_17137,N_16065,N_16947);
nand U17138 (N_17138,N_16363,N_16246);
nand U17139 (N_17139,N_16300,N_16219);
or U17140 (N_17140,N_16887,N_16717);
and U17141 (N_17141,N_16452,N_16259);
and U17142 (N_17142,N_16348,N_16409);
and U17143 (N_17143,N_16001,N_16152);
nand U17144 (N_17144,N_16811,N_16741);
or U17145 (N_17145,N_16448,N_16484);
xnor U17146 (N_17146,N_16057,N_16616);
and U17147 (N_17147,N_16701,N_16914);
or U17148 (N_17148,N_16180,N_16526);
xnor U17149 (N_17149,N_16757,N_16010);
nor U17150 (N_17150,N_16495,N_16674);
nand U17151 (N_17151,N_16889,N_16275);
or U17152 (N_17152,N_16089,N_16498);
or U17153 (N_17153,N_16492,N_16222);
and U17154 (N_17154,N_16047,N_16744);
nand U17155 (N_17155,N_16902,N_16569);
or U17156 (N_17156,N_16302,N_16756);
or U17157 (N_17157,N_16227,N_16938);
xnor U17158 (N_17158,N_16681,N_16470);
or U17159 (N_17159,N_16551,N_16874);
nand U17160 (N_17160,N_16984,N_16848);
nand U17161 (N_17161,N_16360,N_16924);
or U17162 (N_17162,N_16873,N_16214);
nand U17163 (N_17163,N_16535,N_16553);
nor U17164 (N_17164,N_16819,N_16769);
xor U17165 (N_17165,N_16069,N_16733);
nor U17166 (N_17166,N_16000,N_16087);
nand U17167 (N_17167,N_16656,N_16356);
xnor U17168 (N_17168,N_16325,N_16903);
and U17169 (N_17169,N_16518,N_16864);
and U17170 (N_17170,N_16514,N_16162);
nor U17171 (N_17171,N_16932,N_16447);
xnor U17172 (N_17172,N_16735,N_16342);
nor U17173 (N_17173,N_16752,N_16404);
nand U17174 (N_17174,N_16511,N_16487);
nand U17175 (N_17175,N_16459,N_16215);
and U17176 (N_17176,N_16033,N_16031);
xor U17177 (N_17177,N_16963,N_16317);
and U17178 (N_17178,N_16501,N_16692);
or U17179 (N_17179,N_16436,N_16240);
or U17180 (N_17180,N_16576,N_16824);
and U17181 (N_17181,N_16672,N_16251);
xnor U17182 (N_17182,N_16944,N_16118);
or U17183 (N_17183,N_16489,N_16123);
and U17184 (N_17184,N_16950,N_16354);
or U17185 (N_17185,N_16990,N_16812);
nor U17186 (N_17186,N_16849,N_16032);
or U17187 (N_17187,N_16066,N_16376);
xor U17188 (N_17188,N_16939,N_16758);
nand U17189 (N_17189,N_16136,N_16476);
nor U17190 (N_17190,N_16575,N_16904);
xnor U17191 (N_17191,N_16585,N_16181);
and U17192 (N_17192,N_16640,N_16519);
or U17193 (N_17193,N_16091,N_16350);
xnor U17194 (N_17194,N_16975,N_16009);
nand U17195 (N_17195,N_16052,N_16766);
or U17196 (N_17196,N_16238,N_16531);
xor U17197 (N_17197,N_16163,N_16117);
and U17198 (N_17198,N_16156,N_16177);
xnor U17199 (N_17199,N_16602,N_16014);
xnor U17200 (N_17200,N_16349,N_16625);
or U17201 (N_17201,N_16172,N_16619);
and U17202 (N_17202,N_16471,N_16265);
or U17203 (N_17203,N_16485,N_16900);
or U17204 (N_17204,N_16609,N_16869);
nand U17205 (N_17205,N_16249,N_16337);
nor U17206 (N_17206,N_16233,N_16834);
nor U17207 (N_17207,N_16011,N_16423);
nor U17208 (N_17208,N_16534,N_16115);
xnor U17209 (N_17209,N_16169,N_16632);
or U17210 (N_17210,N_16433,N_16490);
or U17211 (N_17211,N_16745,N_16319);
nand U17212 (N_17212,N_16486,N_16891);
or U17213 (N_17213,N_16201,N_16051);
or U17214 (N_17214,N_16659,N_16934);
or U17215 (N_17215,N_16410,N_16943);
and U17216 (N_17216,N_16788,N_16893);
xor U17217 (N_17217,N_16151,N_16973);
nand U17218 (N_17218,N_16415,N_16724);
xor U17219 (N_17219,N_16936,N_16401);
or U17220 (N_17220,N_16384,N_16829);
nor U17221 (N_17221,N_16107,N_16917);
and U17222 (N_17222,N_16564,N_16879);
or U17223 (N_17223,N_16761,N_16359);
or U17224 (N_17224,N_16131,N_16442);
or U17225 (N_17225,N_16358,N_16908);
nand U17226 (N_17226,N_16128,N_16791);
nor U17227 (N_17227,N_16850,N_16599);
or U17228 (N_17228,N_16141,N_16762);
nor U17229 (N_17229,N_16650,N_16807);
xor U17230 (N_17230,N_16574,N_16054);
nor U17231 (N_17231,N_16550,N_16601);
nor U17232 (N_17232,N_16160,N_16790);
and U17233 (N_17233,N_16515,N_16814);
and U17234 (N_17234,N_16852,N_16081);
and U17235 (N_17235,N_16028,N_16643);
or U17236 (N_17236,N_16872,N_16456);
nand U17237 (N_17237,N_16434,N_16759);
xnor U17238 (N_17238,N_16974,N_16399);
nor U17239 (N_17239,N_16197,N_16184);
or U17240 (N_17240,N_16621,N_16665);
or U17241 (N_17241,N_16774,N_16581);
and U17242 (N_17242,N_16843,N_16649);
or U17243 (N_17243,N_16134,N_16578);
xnor U17244 (N_17244,N_16722,N_16517);
xnor U17245 (N_17245,N_16135,N_16586);
nand U17246 (N_17246,N_16707,N_16755);
nor U17247 (N_17247,N_16847,N_16631);
nor U17248 (N_17248,N_16213,N_16017);
or U17249 (N_17249,N_16211,N_16929);
nor U17250 (N_17250,N_16690,N_16749);
nor U17251 (N_17251,N_16269,N_16029);
xnor U17252 (N_17252,N_16666,N_16870);
and U17253 (N_17253,N_16204,N_16086);
xnor U17254 (N_17254,N_16264,N_16881);
nor U17255 (N_17255,N_16225,N_16928);
or U17256 (N_17256,N_16813,N_16272);
nand U17257 (N_17257,N_16124,N_16042);
nor U17258 (N_17258,N_16208,N_16743);
nand U17259 (N_17259,N_16629,N_16252);
or U17260 (N_17260,N_16226,N_16217);
or U17261 (N_17261,N_16778,N_16303);
and U17262 (N_17262,N_16380,N_16826);
nand U17263 (N_17263,N_16205,N_16637);
nor U17264 (N_17264,N_16727,N_16986);
xnor U17265 (N_17265,N_16241,N_16083);
or U17266 (N_17266,N_16557,N_16667);
xnor U17267 (N_17267,N_16892,N_16700);
nor U17268 (N_17268,N_16060,N_16771);
nand U17269 (N_17269,N_16837,N_16897);
nor U17270 (N_17270,N_16953,N_16867);
nand U17271 (N_17271,N_16425,N_16781);
and U17272 (N_17272,N_16478,N_16464);
and U17273 (N_17273,N_16565,N_16283);
nor U17274 (N_17274,N_16951,N_16675);
or U17275 (N_17275,N_16737,N_16462);
nor U17276 (N_17276,N_16035,N_16607);
xnor U17277 (N_17277,N_16159,N_16740);
nor U17278 (N_17278,N_16046,N_16015);
nand U17279 (N_17279,N_16655,N_16704);
nand U17280 (N_17280,N_16693,N_16003);
nor U17281 (N_17281,N_16413,N_16138);
nand U17282 (N_17282,N_16147,N_16697);
nand U17283 (N_17283,N_16925,N_16676);
and U17284 (N_17284,N_16428,N_16268);
nand U17285 (N_17285,N_16503,N_16242);
nor U17286 (N_17286,N_16406,N_16858);
nor U17287 (N_17287,N_16261,N_16835);
nor U17288 (N_17288,N_16004,N_16113);
and U17289 (N_17289,N_16393,N_16823);
xor U17290 (N_17290,N_16901,N_16554);
nand U17291 (N_17291,N_16194,N_16295);
nand U17292 (N_17292,N_16894,N_16304);
nor U17293 (N_17293,N_16458,N_16045);
xor U17294 (N_17294,N_16255,N_16798);
and U17295 (N_17295,N_16170,N_16027);
xnor U17296 (N_17296,N_16815,N_16970);
or U17297 (N_17297,N_16299,N_16862);
nand U17298 (N_17298,N_16876,N_16748);
and U17299 (N_17299,N_16088,N_16253);
nor U17300 (N_17300,N_16775,N_16392);
xnor U17301 (N_17301,N_16281,N_16804);
nor U17302 (N_17302,N_16598,N_16106);
nand U17303 (N_17303,N_16549,N_16058);
or U17304 (N_17304,N_16216,N_16329);
nor U17305 (N_17305,N_16547,N_16440);
or U17306 (N_17306,N_16129,N_16830);
or U17307 (N_17307,N_16822,N_16695);
nand U17308 (N_17308,N_16571,N_16430);
xnor U17309 (N_17309,N_16340,N_16673);
or U17310 (N_17310,N_16959,N_16109);
nand U17311 (N_17311,N_16427,N_16603);
and U17312 (N_17312,N_16419,N_16165);
or U17313 (N_17313,N_16173,N_16841);
and U17314 (N_17314,N_16050,N_16020);
nor U17315 (N_17315,N_16983,N_16825);
and U17316 (N_17316,N_16346,N_16863);
nor U17317 (N_17317,N_16624,N_16454);
nor U17318 (N_17318,N_16909,N_16394);
xnor U17319 (N_17319,N_16777,N_16161);
xor U17320 (N_17320,N_16101,N_16431);
and U17321 (N_17321,N_16647,N_16803);
xor U17322 (N_17322,N_16491,N_16018);
xor U17323 (N_17323,N_16053,N_16338);
and U17324 (N_17324,N_16539,N_16468);
nand U17325 (N_17325,N_16328,N_16563);
xor U17326 (N_17326,N_16508,N_16418);
or U17327 (N_17327,N_16708,N_16865);
xor U17328 (N_17328,N_16949,N_16520);
xor U17329 (N_17329,N_16441,N_16682);
xor U17330 (N_17330,N_16074,N_16068);
xor U17331 (N_17331,N_16254,N_16529);
or U17332 (N_17332,N_16782,N_16558);
xor U17333 (N_17333,N_16787,N_16770);
nand U17334 (N_17334,N_16580,N_16732);
nand U17335 (N_17335,N_16506,N_16411);
nor U17336 (N_17336,N_16671,N_16378);
xnor U17337 (N_17337,N_16157,N_16361);
and U17338 (N_17338,N_16919,N_16479);
or U17339 (N_17339,N_16502,N_16036);
or U17340 (N_17340,N_16634,N_16998);
and U17341 (N_17341,N_16292,N_16258);
xor U17342 (N_17342,N_16799,N_16382);
nor U17343 (N_17343,N_16930,N_16311);
nand U17344 (N_17344,N_16606,N_16076);
nor U17345 (N_17345,N_16999,N_16473);
nand U17346 (N_17346,N_16271,N_16723);
and U17347 (N_17347,N_16855,N_16633);
nor U17348 (N_17348,N_16202,N_16345);
nor U17349 (N_17349,N_16910,N_16968);
and U17350 (N_17350,N_16059,N_16111);
xnor U17351 (N_17351,N_16605,N_16312);
xnor U17352 (N_17352,N_16773,N_16711);
and U17353 (N_17353,N_16560,N_16646);
xnor U17354 (N_17354,N_16408,N_16691);
xnor U17355 (N_17355,N_16237,N_16920);
nor U17356 (N_17356,N_16239,N_16330);
nand U17357 (N_17357,N_16316,N_16355);
nand U17358 (N_17358,N_16989,N_16218);
or U17359 (N_17359,N_16095,N_16145);
and U17360 (N_17360,N_16617,N_16927);
nor U17361 (N_17361,N_16426,N_16067);
xor U17362 (N_17362,N_16270,N_16366);
or U17363 (N_17363,N_16592,N_16718);
nand U17364 (N_17364,N_16593,N_16698);
xor U17365 (N_17365,N_16931,N_16294);
or U17366 (N_17366,N_16942,N_16445);
xor U17367 (N_17367,N_16859,N_16133);
nand U17368 (N_17368,N_16199,N_16196);
or U17369 (N_17369,N_16188,N_16341);
nor U17370 (N_17370,N_16056,N_16022);
nor U17371 (N_17371,N_16315,N_16712);
nand U17372 (N_17372,N_16353,N_16923);
nand U17373 (N_17373,N_16187,N_16336);
or U17374 (N_17374,N_16753,N_16422);
and U17375 (N_17375,N_16043,N_16793);
xor U17376 (N_17376,N_16868,N_16591);
and U17377 (N_17377,N_16779,N_16896);
or U17378 (N_17378,N_16726,N_16946);
nor U17379 (N_17379,N_16125,N_16838);
nor U17380 (N_17380,N_16278,N_16412);
xnor U17381 (N_17381,N_16583,N_16077);
xnor U17382 (N_17382,N_16993,N_16561);
nor U17383 (N_17383,N_16049,N_16579);
nor U17384 (N_17384,N_16831,N_16933);
nor U17385 (N_17385,N_16126,N_16347);
nor U17386 (N_17386,N_16604,N_16505);
or U17387 (N_17387,N_16334,N_16182);
nand U17388 (N_17388,N_16192,N_16405);
or U17389 (N_17389,N_16244,N_16379);
or U17390 (N_17390,N_16064,N_16063);
nor U17391 (N_17391,N_16710,N_16457);
or U17392 (N_17392,N_16750,N_16662);
and U17393 (N_17393,N_16176,N_16728);
nand U17394 (N_17394,N_16041,N_16577);
nand U17395 (N_17395,N_16450,N_16391);
nand U17396 (N_17396,N_16820,N_16622);
nand U17397 (N_17397,N_16260,N_16084);
and U17398 (N_17398,N_16191,N_16854);
xnor U17399 (N_17399,N_16203,N_16739);
xor U17400 (N_17400,N_16907,N_16071);
nor U17401 (N_17401,N_16209,N_16466);
and U17402 (N_17402,N_16528,N_16277);
and U17403 (N_17403,N_16805,N_16888);
nand U17404 (N_17404,N_16980,N_16566);
nand U17405 (N_17405,N_16608,N_16871);
nand U17406 (N_17406,N_16232,N_16496);
nor U17407 (N_17407,N_16250,N_16098);
or U17408 (N_17408,N_16500,N_16952);
and U17409 (N_17409,N_16364,N_16367);
xnor U17410 (N_17410,N_16618,N_16424);
nor U17411 (N_17411,N_16785,N_16375);
nand U17412 (N_17412,N_16421,N_16573);
xor U17413 (N_17413,N_16210,N_16719);
or U17414 (N_17414,N_16221,N_16097);
xnor U17415 (N_17415,N_16856,N_16324);
and U17416 (N_17416,N_16085,N_16540);
xor U17417 (N_17417,N_16861,N_16139);
and U17418 (N_17418,N_16108,N_16809);
xnor U17419 (N_17419,N_16186,N_16996);
nand U17420 (N_17420,N_16628,N_16198);
nand U17421 (N_17421,N_16235,N_16212);
nor U17422 (N_17422,N_16796,N_16224);
xor U17423 (N_17423,N_16940,N_16827);
and U17424 (N_17424,N_16784,N_16070);
nand U17425 (N_17425,N_16630,N_16243);
xor U17426 (N_17426,N_16981,N_16543);
xnor U17427 (N_17427,N_16414,N_16661);
and U17428 (N_17428,N_16343,N_16021);
nor U17429 (N_17429,N_16615,N_16149);
or U17430 (N_17430,N_16407,N_16522);
xnor U17431 (N_17431,N_16398,N_16403);
xor U17432 (N_17432,N_16247,N_16482);
nand U17433 (N_17433,N_16721,N_16320);
or U17434 (N_17434,N_16890,N_16627);
nor U17435 (N_17435,N_16444,N_16477);
or U17436 (N_17436,N_16193,N_16480);
and U17437 (N_17437,N_16102,N_16155);
nand U17438 (N_17438,N_16112,N_16397);
and U17439 (N_17439,N_16387,N_16158);
xnor U17440 (N_17440,N_16687,N_16171);
or U17441 (N_17441,N_16189,N_16183);
xor U17442 (N_17442,N_16642,N_16702);
xnor U17443 (N_17443,N_16079,N_16110);
xnor U17444 (N_17444,N_16467,N_16142);
nor U17445 (N_17445,N_16582,N_16765);
and U17446 (N_17446,N_16062,N_16103);
nor U17447 (N_17447,N_16982,N_16746);
and U17448 (N_17448,N_16600,N_16154);
or U17449 (N_17449,N_16357,N_16636);
or U17450 (N_17450,N_16572,N_16548);
nand U17451 (N_17451,N_16795,N_16954);
or U17452 (N_17452,N_16438,N_16037);
or U17453 (N_17453,N_16080,N_16463);
xor U17454 (N_17454,N_16012,N_16562);
nand U17455 (N_17455,N_16280,N_16234);
xnor U17456 (N_17456,N_16223,N_16121);
and U17457 (N_17457,N_16351,N_16967);
xor U17458 (N_17458,N_16679,N_16166);
or U17459 (N_17459,N_16651,N_16994);
or U17460 (N_17460,N_16786,N_16093);
and U17461 (N_17461,N_16402,N_16293);
nor U17462 (N_17462,N_16417,N_16504);
xnor U17463 (N_17463,N_16801,N_16090);
nor U17464 (N_17464,N_16298,N_16767);
nand U17465 (N_17465,N_16195,N_16396);
and U17466 (N_17466,N_16461,N_16263);
nor U17467 (N_17467,N_16245,N_16623);
and U17468 (N_17468,N_16905,N_16344);
nor U17469 (N_17469,N_16488,N_16694);
nand U17470 (N_17470,N_16768,N_16663);
nor U17471 (N_17471,N_16668,N_16368);
and U17472 (N_17472,N_16921,N_16122);
nand U17473 (N_17473,N_16390,N_16007);
xor U17474 (N_17474,N_16497,N_16061);
nand U17475 (N_17475,N_16783,N_16527);
or U17476 (N_17476,N_16230,N_16326);
nand U17477 (N_17477,N_16683,N_16465);
nor U17478 (N_17478,N_16148,N_16327);
nand U17479 (N_17479,N_16806,N_16034);
or U17480 (N_17480,N_16306,N_16976);
nor U17481 (N_17481,N_16524,N_16590);
and U17482 (N_17482,N_16313,N_16130);
and U17483 (N_17483,N_16429,N_16810);
and U17484 (N_17484,N_16287,N_16941);
xnor U17485 (N_17485,N_16991,N_16956);
nand U17486 (N_17486,N_16860,N_16279);
nor U17487 (N_17487,N_16435,N_16318);
nor U17488 (N_17488,N_16966,N_16935);
xor U17489 (N_17489,N_16105,N_16715);
xnor U17490 (N_17490,N_16657,N_16985);
xor U17491 (N_17491,N_16541,N_16816);
and U17492 (N_17492,N_16374,N_16532);
nor U17493 (N_17493,N_16639,N_16229);
xnor U17494 (N_17494,N_16997,N_16731);
xnor U17495 (N_17495,N_16220,N_16556);
nor U17496 (N_17496,N_16685,N_16961);
and U17497 (N_17497,N_16915,N_16680);
and U17498 (N_17498,N_16660,N_16256);
nor U17499 (N_17499,N_16100,N_16641);
nor U17500 (N_17500,N_16648,N_16468);
or U17501 (N_17501,N_16580,N_16029);
or U17502 (N_17502,N_16494,N_16688);
and U17503 (N_17503,N_16669,N_16107);
nand U17504 (N_17504,N_16396,N_16857);
and U17505 (N_17505,N_16854,N_16512);
and U17506 (N_17506,N_16736,N_16630);
nor U17507 (N_17507,N_16754,N_16808);
nor U17508 (N_17508,N_16471,N_16665);
nand U17509 (N_17509,N_16733,N_16346);
nand U17510 (N_17510,N_16090,N_16310);
nor U17511 (N_17511,N_16075,N_16234);
or U17512 (N_17512,N_16509,N_16392);
or U17513 (N_17513,N_16765,N_16647);
nor U17514 (N_17514,N_16068,N_16780);
nand U17515 (N_17515,N_16265,N_16511);
or U17516 (N_17516,N_16066,N_16139);
or U17517 (N_17517,N_16203,N_16663);
xnor U17518 (N_17518,N_16201,N_16803);
or U17519 (N_17519,N_16704,N_16439);
or U17520 (N_17520,N_16326,N_16969);
nor U17521 (N_17521,N_16259,N_16583);
nand U17522 (N_17522,N_16825,N_16552);
xnor U17523 (N_17523,N_16645,N_16105);
or U17524 (N_17524,N_16872,N_16027);
or U17525 (N_17525,N_16441,N_16238);
nand U17526 (N_17526,N_16518,N_16739);
nand U17527 (N_17527,N_16615,N_16523);
nand U17528 (N_17528,N_16294,N_16875);
xor U17529 (N_17529,N_16839,N_16506);
nand U17530 (N_17530,N_16907,N_16544);
xor U17531 (N_17531,N_16128,N_16184);
nor U17532 (N_17532,N_16781,N_16079);
xor U17533 (N_17533,N_16490,N_16538);
xor U17534 (N_17534,N_16917,N_16392);
nor U17535 (N_17535,N_16015,N_16343);
or U17536 (N_17536,N_16193,N_16172);
xnor U17537 (N_17537,N_16798,N_16912);
nand U17538 (N_17538,N_16389,N_16291);
or U17539 (N_17539,N_16774,N_16747);
or U17540 (N_17540,N_16414,N_16111);
and U17541 (N_17541,N_16399,N_16256);
or U17542 (N_17542,N_16918,N_16493);
or U17543 (N_17543,N_16994,N_16597);
or U17544 (N_17544,N_16812,N_16407);
and U17545 (N_17545,N_16462,N_16915);
xnor U17546 (N_17546,N_16066,N_16920);
nand U17547 (N_17547,N_16777,N_16273);
or U17548 (N_17548,N_16026,N_16269);
nand U17549 (N_17549,N_16347,N_16419);
or U17550 (N_17550,N_16450,N_16841);
xor U17551 (N_17551,N_16439,N_16517);
xnor U17552 (N_17552,N_16136,N_16191);
xor U17553 (N_17553,N_16298,N_16986);
xnor U17554 (N_17554,N_16151,N_16889);
nand U17555 (N_17555,N_16405,N_16672);
and U17556 (N_17556,N_16623,N_16445);
nor U17557 (N_17557,N_16957,N_16848);
or U17558 (N_17558,N_16357,N_16593);
and U17559 (N_17559,N_16381,N_16583);
nand U17560 (N_17560,N_16057,N_16825);
or U17561 (N_17561,N_16702,N_16999);
and U17562 (N_17562,N_16018,N_16666);
nor U17563 (N_17563,N_16044,N_16132);
or U17564 (N_17564,N_16444,N_16980);
nand U17565 (N_17565,N_16887,N_16479);
or U17566 (N_17566,N_16295,N_16296);
nand U17567 (N_17567,N_16972,N_16670);
or U17568 (N_17568,N_16302,N_16763);
or U17569 (N_17569,N_16298,N_16799);
xor U17570 (N_17570,N_16471,N_16020);
or U17571 (N_17571,N_16789,N_16347);
or U17572 (N_17572,N_16240,N_16187);
nor U17573 (N_17573,N_16781,N_16598);
or U17574 (N_17574,N_16251,N_16569);
nor U17575 (N_17575,N_16177,N_16834);
nand U17576 (N_17576,N_16790,N_16037);
and U17577 (N_17577,N_16923,N_16132);
xor U17578 (N_17578,N_16320,N_16637);
and U17579 (N_17579,N_16665,N_16206);
and U17580 (N_17580,N_16872,N_16471);
xor U17581 (N_17581,N_16906,N_16590);
nor U17582 (N_17582,N_16924,N_16702);
nor U17583 (N_17583,N_16523,N_16201);
xnor U17584 (N_17584,N_16266,N_16359);
xnor U17585 (N_17585,N_16652,N_16951);
or U17586 (N_17586,N_16542,N_16239);
nand U17587 (N_17587,N_16019,N_16855);
and U17588 (N_17588,N_16338,N_16477);
nand U17589 (N_17589,N_16975,N_16016);
or U17590 (N_17590,N_16884,N_16705);
nand U17591 (N_17591,N_16567,N_16020);
nand U17592 (N_17592,N_16166,N_16803);
nor U17593 (N_17593,N_16134,N_16143);
nand U17594 (N_17594,N_16763,N_16205);
nand U17595 (N_17595,N_16410,N_16992);
nor U17596 (N_17596,N_16838,N_16158);
xnor U17597 (N_17597,N_16065,N_16429);
nor U17598 (N_17598,N_16974,N_16882);
or U17599 (N_17599,N_16022,N_16917);
xor U17600 (N_17600,N_16224,N_16897);
nor U17601 (N_17601,N_16626,N_16686);
and U17602 (N_17602,N_16875,N_16045);
nor U17603 (N_17603,N_16808,N_16450);
nor U17604 (N_17604,N_16271,N_16468);
nor U17605 (N_17605,N_16139,N_16753);
or U17606 (N_17606,N_16593,N_16834);
nor U17607 (N_17607,N_16618,N_16612);
or U17608 (N_17608,N_16293,N_16917);
nor U17609 (N_17609,N_16967,N_16723);
or U17610 (N_17610,N_16371,N_16681);
xor U17611 (N_17611,N_16107,N_16867);
xnor U17612 (N_17612,N_16116,N_16546);
and U17613 (N_17613,N_16751,N_16131);
or U17614 (N_17614,N_16367,N_16100);
nor U17615 (N_17615,N_16695,N_16220);
nand U17616 (N_17616,N_16842,N_16504);
or U17617 (N_17617,N_16627,N_16714);
and U17618 (N_17618,N_16832,N_16190);
xnor U17619 (N_17619,N_16991,N_16022);
or U17620 (N_17620,N_16165,N_16055);
nor U17621 (N_17621,N_16787,N_16876);
xnor U17622 (N_17622,N_16837,N_16068);
or U17623 (N_17623,N_16208,N_16092);
or U17624 (N_17624,N_16669,N_16783);
nand U17625 (N_17625,N_16533,N_16757);
nor U17626 (N_17626,N_16866,N_16918);
or U17627 (N_17627,N_16283,N_16722);
and U17628 (N_17628,N_16837,N_16109);
nand U17629 (N_17629,N_16555,N_16948);
nand U17630 (N_17630,N_16211,N_16823);
nand U17631 (N_17631,N_16399,N_16727);
nand U17632 (N_17632,N_16505,N_16241);
or U17633 (N_17633,N_16314,N_16569);
nand U17634 (N_17634,N_16743,N_16041);
or U17635 (N_17635,N_16164,N_16851);
nor U17636 (N_17636,N_16321,N_16992);
and U17637 (N_17637,N_16167,N_16333);
or U17638 (N_17638,N_16049,N_16931);
nand U17639 (N_17639,N_16513,N_16227);
or U17640 (N_17640,N_16185,N_16616);
and U17641 (N_17641,N_16706,N_16205);
nand U17642 (N_17642,N_16082,N_16967);
and U17643 (N_17643,N_16844,N_16550);
and U17644 (N_17644,N_16139,N_16677);
xnor U17645 (N_17645,N_16943,N_16382);
or U17646 (N_17646,N_16595,N_16454);
xnor U17647 (N_17647,N_16146,N_16881);
nor U17648 (N_17648,N_16836,N_16621);
xnor U17649 (N_17649,N_16775,N_16378);
or U17650 (N_17650,N_16659,N_16387);
and U17651 (N_17651,N_16468,N_16381);
or U17652 (N_17652,N_16163,N_16807);
xnor U17653 (N_17653,N_16395,N_16365);
nor U17654 (N_17654,N_16679,N_16002);
nor U17655 (N_17655,N_16928,N_16076);
and U17656 (N_17656,N_16947,N_16287);
and U17657 (N_17657,N_16871,N_16420);
xor U17658 (N_17658,N_16123,N_16991);
nand U17659 (N_17659,N_16968,N_16531);
nand U17660 (N_17660,N_16283,N_16603);
nand U17661 (N_17661,N_16962,N_16667);
and U17662 (N_17662,N_16027,N_16625);
nand U17663 (N_17663,N_16845,N_16092);
nand U17664 (N_17664,N_16358,N_16152);
nor U17665 (N_17665,N_16096,N_16979);
nor U17666 (N_17666,N_16158,N_16622);
or U17667 (N_17667,N_16500,N_16049);
nor U17668 (N_17668,N_16030,N_16707);
and U17669 (N_17669,N_16806,N_16153);
nor U17670 (N_17670,N_16176,N_16921);
or U17671 (N_17671,N_16148,N_16764);
and U17672 (N_17672,N_16409,N_16316);
xor U17673 (N_17673,N_16051,N_16427);
or U17674 (N_17674,N_16286,N_16650);
nand U17675 (N_17675,N_16689,N_16305);
nand U17676 (N_17676,N_16203,N_16340);
nor U17677 (N_17677,N_16023,N_16323);
xnor U17678 (N_17678,N_16087,N_16918);
nor U17679 (N_17679,N_16090,N_16103);
xnor U17680 (N_17680,N_16779,N_16607);
nor U17681 (N_17681,N_16833,N_16534);
and U17682 (N_17682,N_16111,N_16564);
xnor U17683 (N_17683,N_16200,N_16046);
xnor U17684 (N_17684,N_16749,N_16378);
xnor U17685 (N_17685,N_16300,N_16705);
xor U17686 (N_17686,N_16664,N_16252);
xnor U17687 (N_17687,N_16309,N_16947);
nor U17688 (N_17688,N_16239,N_16590);
and U17689 (N_17689,N_16538,N_16877);
and U17690 (N_17690,N_16297,N_16613);
or U17691 (N_17691,N_16217,N_16609);
or U17692 (N_17692,N_16397,N_16303);
and U17693 (N_17693,N_16604,N_16542);
nand U17694 (N_17694,N_16413,N_16187);
or U17695 (N_17695,N_16031,N_16622);
xnor U17696 (N_17696,N_16049,N_16733);
xor U17697 (N_17697,N_16804,N_16303);
or U17698 (N_17698,N_16981,N_16915);
nand U17699 (N_17699,N_16712,N_16054);
nor U17700 (N_17700,N_16686,N_16783);
nor U17701 (N_17701,N_16227,N_16068);
nor U17702 (N_17702,N_16033,N_16825);
nand U17703 (N_17703,N_16022,N_16151);
and U17704 (N_17704,N_16339,N_16564);
xnor U17705 (N_17705,N_16484,N_16427);
or U17706 (N_17706,N_16183,N_16350);
or U17707 (N_17707,N_16198,N_16558);
nand U17708 (N_17708,N_16388,N_16883);
nand U17709 (N_17709,N_16461,N_16424);
nand U17710 (N_17710,N_16842,N_16752);
nand U17711 (N_17711,N_16649,N_16346);
and U17712 (N_17712,N_16302,N_16370);
xnor U17713 (N_17713,N_16591,N_16051);
nand U17714 (N_17714,N_16063,N_16233);
and U17715 (N_17715,N_16508,N_16296);
nand U17716 (N_17716,N_16449,N_16434);
xor U17717 (N_17717,N_16925,N_16162);
and U17718 (N_17718,N_16321,N_16561);
or U17719 (N_17719,N_16736,N_16421);
and U17720 (N_17720,N_16686,N_16905);
or U17721 (N_17721,N_16071,N_16142);
nor U17722 (N_17722,N_16176,N_16877);
and U17723 (N_17723,N_16799,N_16636);
or U17724 (N_17724,N_16591,N_16353);
and U17725 (N_17725,N_16287,N_16361);
or U17726 (N_17726,N_16593,N_16973);
nand U17727 (N_17727,N_16699,N_16411);
nor U17728 (N_17728,N_16298,N_16821);
xnor U17729 (N_17729,N_16017,N_16783);
and U17730 (N_17730,N_16631,N_16422);
and U17731 (N_17731,N_16091,N_16173);
nor U17732 (N_17732,N_16171,N_16263);
xor U17733 (N_17733,N_16324,N_16435);
and U17734 (N_17734,N_16519,N_16391);
nor U17735 (N_17735,N_16089,N_16190);
and U17736 (N_17736,N_16557,N_16852);
or U17737 (N_17737,N_16512,N_16954);
and U17738 (N_17738,N_16520,N_16443);
or U17739 (N_17739,N_16836,N_16269);
or U17740 (N_17740,N_16966,N_16237);
xor U17741 (N_17741,N_16465,N_16643);
nand U17742 (N_17742,N_16116,N_16967);
nor U17743 (N_17743,N_16162,N_16848);
nand U17744 (N_17744,N_16645,N_16135);
nor U17745 (N_17745,N_16924,N_16434);
and U17746 (N_17746,N_16458,N_16876);
xnor U17747 (N_17747,N_16753,N_16269);
nor U17748 (N_17748,N_16837,N_16522);
and U17749 (N_17749,N_16739,N_16102);
nor U17750 (N_17750,N_16804,N_16030);
nand U17751 (N_17751,N_16307,N_16513);
xnor U17752 (N_17752,N_16631,N_16763);
nand U17753 (N_17753,N_16121,N_16964);
or U17754 (N_17754,N_16842,N_16452);
or U17755 (N_17755,N_16551,N_16074);
xnor U17756 (N_17756,N_16402,N_16092);
and U17757 (N_17757,N_16934,N_16163);
or U17758 (N_17758,N_16298,N_16819);
nand U17759 (N_17759,N_16190,N_16931);
and U17760 (N_17760,N_16088,N_16967);
and U17761 (N_17761,N_16416,N_16665);
nand U17762 (N_17762,N_16000,N_16953);
xor U17763 (N_17763,N_16107,N_16714);
and U17764 (N_17764,N_16156,N_16696);
nand U17765 (N_17765,N_16698,N_16993);
xnor U17766 (N_17766,N_16114,N_16132);
xnor U17767 (N_17767,N_16122,N_16271);
nand U17768 (N_17768,N_16382,N_16913);
or U17769 (N_17769,N_16302,N_16807);
nor U17770 (N_17770,N_16368,N_16117);
xnor U17771 (N_17771,N_16582,N_16538);
nand U17772 (N_17772,N_16770,N_16568);
or U17773 (N_17773,N_16157,N_16468);
and U17774 (N_17774,N_16165,N_16531);
and U17775 (N_17775,N_16366,N_16032);
and U17776 (N_17776,N_16547,N_16704);
or U17777 (N_17777,N_16509,N_16965);
and U17778 (N_17778,N_16063,N_16690);
nor U17779 (N_17779,N_16669,N_16641);
and U17780 (N_17780,N_16038,N_16627);
or U17781 (N_17781,N_16367,N_16514);
nand U17782 (N_17782,N_16320,N_16329);
or U17783 (N_17783,N_16741,N_16695);
and U17784 (N_17784,N_16825,N_16805);
and U17785 (N_17785,N_16080,N_16148);
or U17786 (N_17786,N_16086,N_16083);
nand U17787 (N_17787,N_16867,N_16575);
nand U17788 (N_17788,N_16373,N_16717);
and U17789 (N_17789,N_16390,N_16835);
and U17790 (N_17790,N_16175,N_16923);
nand U17791 (N_17791,N_16772,N_16306);
nand U17792 (N_17792,N_16771,N_16625);
and U17793 (N_17793,N_16248,N_16848);
nand U17794 (N_17794,N_16295,N_16907);
xnor U17795 (N_17795,N_16670,N_16155);
or U17796 (N_17796,N_16982,N_16080);
and U17797 (N_17797,N_16428,N_16083);
or U17798 (N_17798,N_16268,N_16237);
xnor U17799 (N_17799,N_16836,N_16389);
nand U17800 (N_17800,N_16989,N_16098);
and U17801 (N_17801,N_16779,N_16586);
xnor U17802 (N_17802,N_16695,N_16940);
nand U17803 (N_17803,N_16110,N_16471);
nand U17804 (N_17804,N_16880,N_16608);
nand U17805 (N_17805,N_16300,N_16418);
nor U17806 (N_17806,N_16026,N_16604);
nor U17807 (N_17807,N_16878,N_16819);
xnor U17808 (N_17808,N_16406,N_16673);
nand U17809 (N_17809,N_16794,N_16371);
and U17810 (N_17810,N_16218,N_16684);
xnor U17811 (N_17811,N_16235,N_16738);
nand U17812 (N_17812,N_16494,N_16041);
xor U17813 (N_17813,N_16664,N_16870);
nor U17814 (N_17814,N_16384,N_16339);
or U17815 (N_17815,N_16914,N_16695);
or U17816 (N_17816,N_16883,N_16269);
and U17817 (N_17817,N_16360,N_16423);
xnor U17818 (N_17818,N_16342,N_16496);
nor U17819 (N_17819,N_16583,N_16123);
or U17820 (N_17820,N_16968,N_16032);
nand U17821 (N_17821,N_16448,N_16575);
xor U17822 (N_17822,N_16678,N_16009);
xnor U17823 (N_17823,N_16073,N_16781);
and U17824 (N_17824,N_16444,N_16903);
xor U17825 (N_17825,N_16102,N_16261);
nand U17826 (N_17826,N_16787,N_16641);
nor U17827 (N_17827,N_16630,N_16110);
xor U17828 (N_17828,N_16226,N_16719);
nand U17829 (N_17829,N_16355,N_16534);
or U17830 (N_17830,N_16467,N_16319);
xor U17831 (N_17831,N_16642,N_16818);
or U17832 (N_17832,N_16937,N_16259);
and U17833 (N_17833,N_16916,N_16604);
or U17834 (N_17834,N_16022,N_16359);
or U17835 (N_17835,N_16346,N_16008);
nor U17836 (N_17836,N_16693,N_16508);
or U17837 (N_17837,N_16714,N_16648);
and U17838 (N_17838,N_16405,N_16411);
nand U17839 (N_17839,N_16693,N_16922);
nand U17840 (N_17840,N_16413,N_16077);
nand U17841 (N_17841,N_16288,N_16647);
nand U17842 (N_17842,N_16265,N_16140);
nand U17843 (N_17843,N_16598,N_16335);
xnor U17844 (N_17844,N_16226,N_16167);
xor U17845 (N_17845,N_16985,N_16233);
xor U17846 (N_17846,N_16224,N_16740);
and U17847 (N_17847,N_16834,N_16613);
nor U17848 (N_17848,N_16149,N_16294);
or U17849 (N_17849,N_16125,N_16380);
or U17850 (N_17850,N_16807,N_16474);
nor U17851 (N_17851,N_16948,N_16527);
and U17852 (N_17852,N_16348,N_16671);
nand U17853 (N_17853,N_16819,N_16806);
xor U17854 (N_17854,N_16516,N_16434);
nor U17855 (N_17855,N_16998,N_16132);
nor U17856 (N_17856,N_16236,N_16464);
and U17857 (N_17857,N_16183,N_16563);
nand U17858 (N_17858,N_16662,N_16268);
or U17859 (N_17859,N_16495,N_16657);
and U17860 (N_17860,N_16159,N_16906);
or U17861 (N_17861,N_16417,N_16166);
nor U17862 (N_17862,N_16487,N_16783);
nand U17863 (N_17863,N_16551,N_16244);
xor U17864 (N_17864,N_16928,N_16405);
nor U17865 (N_17865,N_16567,N_16142);
nor U17866 (N_17866,N_16362,N_16888);
nand U17867 (N_17867,N_16660,N_16939);
or U17868 (N_17868,N_16575,N_16346);
and U17869 (N_17869,N_16432,N_16508);
nor U17870 (N_17870,N_16194,N_16856);
and U17871 (N_17871,N_16514,N_16973);
nand U17872 (N_17872,N_16331,N_16677);
nand U17873 (N_17873,N_16124,N_16790);
or U17874 (N_17874,N_16789,N_16868);
or U17875 (N_17875,N_16435,N_16028);
nand U17876 (N_17876,N_16246,N_16521);
or U17877 (N_17877,N_16226,N_16907);
xnor U17878 (N_17878,N_16928,N_16408);
and U17879 (N_17879,N_16087,N_16101);
nand U17880 (N_17880,N_16583,N_16879);
or U17881 (N_17881,N_16997,N_16112);
or U17882 (N_17882,N_16708,N_16899);
nor U17883 (N_17883,N_16017,N_16852);
nand U17884 (N_17884,N_16304,N_16831);
and U17885 (N_17885,N_16681,N_16725);
and U17886 (N_17886,N_16066,N_16389);
and U17887 (N_17887,N_16601,N_16019);
xor U17888 (N_17888,N_16436,N_16174);
nor U17889 (N_17889,N_16996,N_16224);
and U17890 (N_17890,N_16355,N_16715);
and U17891 (N_17891,N_16123,N_16649);
nor U17892 (N_17892,N_16128,N_16091);
or U17893 (N_17893,N_16095,N_16399);
and U17894 (N_17894,N_16912,N_16212);
nor U17895 (N_17895,N_16860,N_16611);
or U17896 (N_17896,N_16200,N_16518);
and U17897 (N_17897,N_16210,N_16055);
and U17898 (N_17898,N_16700,N_16576);
and U17899 (N_17899,N_16079,N_16136);
or U17900 (N_17900,N_16201,N_16196);
and U17901 (N_17901,N_16903,N_16836);
nor U17902 (N_17902,N_16736,N_16732);
nand U17903 (N_17903,N_16654,N_16420);
or U17904 (N_17904,N_16415,N_16328);
xor U17905 (N_17905,N_16553,N_16222);
xor U17906 (N_17906,N_16762,N_16885);
or U17907 (N_17907,N_16423,N_16825);
nand U17908 (N_17908,N_16741,N_16074);
nor U17909 (N_17909,N_16386,N_16401);
nand U17910 (N_17910,N_16893,N_16374);
xnor U17911 (N_17911,N_16750,N_16017);
and U17912 (N_17912,N_16516,N_16006);
or U17913 (N_17913,N_16797,N_16934);
nand U17914 (N_17914,N_16275,N_16571);
or U17915 (N_17915,N_16256,N_16410);
xnor U17916 (N_17916,N_16802,N_16050);
nand U17917 (N_17917,N_16032,N_16022);
nor U17918 (N_17918,N_16404,N_16992);
and U17919 (N_17919,N_16227,N_16285);
or U17920 (N_17920,N_16430,N_16518);
or U17921 (N_17921,N_16373,N_16885);
and U17922 (N_17922,N_16523,N_16796);
or U17923 (N_17923,N_16451,N_16136);
or U17924 (N_17924,N_16489,N_16496);
xnor U17925 (N_17925,N_16261,N_16990);
or U17926 (N_17926,N_16670,N_16576);
nor U17927 (N_17927,N_16063,N_16904);
nand U17928 (N_17928,N_16645,N_16727);
and U17929 (N_17929,N_16996,N_16208);
nand U17930 (N_17930,N_16705,N_16054);
nor U17931 (N_17931,N_16965,N_16200);
and U17932 (N_17932,N_16182,N_16233);
or U17933 (N_17933,N_16796,N_16792);
nand U17934 (N_17934,N_16136,N_16008);
nor U17935 (N_17935,N_16454,N_16243);
or U17936 (N_17936,N_16830,N_16668);
xnor U17937 (N_17937,N_16382,N_16297);
nand U17938 (N_17938,N_16541,N_16576);
or U17939 (N_17939,N_16911,N_16417);
and U17940 (N_17940,N_16764,N_16994);
nor U17941 (N_17941,N_16487,N_16029);
and U17942 (N_17942,N_16441,N_16415);
or U17943 (N_17943,N_16032,N_16514);
and U17944 (N_17944,N_16488,N_16979);
nor U17945 (N_17945,N_16076,N_16132);
or U17946 (N_17946,N_16094,N_16095);
nand U17947 (N_17947,N_16023,N_16745);
nand U17948 (N_17948,N_16017,N_16994);
and U17949 (N_17949,N_16933,N_16132);
nand U17950 (N_17950,N_16574,N_16102);
and U17951 (N_17951,N_16670,N_16642);
xnor U17952 (N_17952,N_16712,N_16410);
xnor U17953 (N_17953,N_16178,N_16916);
xnor U17954 (N_17954,N_16739,N_16770);
or U17955 (N_17955,N_16969,N_16127);
and U17956 (N_17956,N_16945,N_16229);
xnor U17957 (N_17957,N_16002,N_16537);
xor U17958 (N_17958,N_16116,N_16095);
and U17959 (N_17959,N_16134,N_16329);
and U17960 (N_17960,N_16617,N_16930);
or U17961 (N_17961,N_16516,N_16368);
and U17962 (N_17962,N_16892,N_16587);
nand U17963 (N_17963,N_16100,N_16103);
and U17964 (N_17964,N_16527,N_16242);
xor U17965 (N_17965,N_16946,N_16413);
nor U17966 (N_17966,N_16693,N_16455);
nor U17967 (N_17967,N_16164,N_16623);
or U17968 (N_17968,N_16683,N_16617);
nor U17969 (N_17969,N_16550,N_16283);
or U17970 (N_17970,N_16770,N_16260);
and U17971 (N_17971,N_16966,N_16161);
and U17972 (N_17972,N_16277,N_16519);
xnor U17973 (N_17973,N_16022,N_16244);
xor U17974 (N_17974,N_16949,N_16765);
nor U17975 (N_17975,N_16768,N_16740);
xor U17976 (N_17976,N_16923,N_16029);
and U17977 (N_17977,N_16267,N_16900);
nor U17978 (N_17978,N_16720,N_16267);
or U17979 (N_17979,N_16219,N_16217);
nor U17980 (N_17980,N_16352,N_16988);
nand U17981 (N_17981,N_16917,N_16370);
nand U17982 (N_17982,N_16961,N_16073);
nand U17983 (N_17983,N_16296,N_16430);
nand U17984 (N_17984,N_16395,N_16387);
nor U17985 (N_17985,N_16390,N_16060);
nor U17986 (N_17986,N_16051,N_16648);
xor U17987 (N_17987,N_16094,N_16433);
nand U17988 (N_17988,N_16443,N_16555);
or U17989 (N_17989,N_16639,N_16134);
xnor U17990 (N_17990,N_16188,N_16171);
xor U17991 (N_17991,N_16256,N_16456);
nand U17992 (N_17992,N_16373,N_16646);
or U17993 (N_17993,N_16120,N_16340);
nor U17994 (N_17994,N_16644,N_16264);
nand U17995 (N_17995,N_16979,N_16655);
nor U17996 (N_17996,N_16128,N_16929);
nor U17997 (N_17997,N_16192,N_16734);
and U17998 (N_17998,N_16873,N_16198);
nand U17999 (N_17999,N_16598,N_16934);
and U18000 (N_18000,N_17282,N_17361);
nand U18001 (N_18001,N_17280,N_17024);
or U18002 (N_18002,N_17208,N_17342);
nor U18003 (N_18003,N_17083,N_17314);
nor U18004 (N_18004,N_17009,N_17265);
nand U18005 (N_18005,N_17848,N_17476);
nand U18006 (N_18006,N_17446,N_17750);
or U18007 (N_18007,N_17878,N_17398);
nor U18008 (N_18008,N_17684,N_17195);
and U18009 (N_18009,N_17906,N_17251);
and U18010 (N_18010,N_17775,N_17281);
xnor U18011 (N_18011,N_17839,N_17834);
and U18012 (N_18012,N_17113,N_17308);
xor U18013 (N_18013,N_17223,N_17135);
nand U18014 (N_18014,N_17094,N_17924);
nand U18015 (N_18015,N_17136,N_17787);
xnor U18016 (N_18016,N_17564,N_17007);
xor U18017 (N_18017,N_17451,N_17663);
xnor U18018 (N_18018,N_17077,N_17606);
nand U18019 (N_18019,N_17743,N_17440);
and U18020 (N_18020,N_17394,N_17101);
xnor U18021 (N_18021,N_17941,N_17719);
or U18022 (N_18022,N_17213,N_17233);
xnor U18023 (N_18023,N_17329,N_17250);
nor U18024 (N_18024,N_17738,N_17594);
xor U18025 (N_18025,N_17469,N_17279);
nor U18026 (N_18026,N_17784,N_17563);
nor U18027 (N_18027,N_17006,N_17244);
and U18028 (N_18028,N_17060,N_17598);
and U18029 (N_18029,N_17286,N_17146);
nand U18030 (N_18030,N_17069,N_17845);
xor U18031 (N_18031,N_17708,N_17652);
xnor U18032 (N_18032,N_17876,N_17133);
or U18033 (N_18033,N_17152,N_17484);
and U18034 (N_18034,N_17013,N_17438);
and U18035 (N_18035,N_17258,N_17592);
nand U18036 (N_18036,N_17796,N_17953);
nand U18037 (N_18037,N_17826,N_17224);
and U18038 (N_18038,N_17338,N_17502);
nor U18039 (N_18039,N_17819,N_17657);
or U18040 (N_18040,N_17068,N_17951);
nand U18041 (N_18041,N_17707,N_17190);
nor U18042 (N_18042,N_17119,N_17519);
or U18043 (N_18043,N_17752,N_17940);
nor U18044 (N_18044,N_17745,N_17794);
or U18045 (N_18045,N_17340,N_17534);
xnor U18046 (N_18046,N_17595,N_17716);
xor U18047 (N_18047,N_17769,N_17260);
or U18048 (N_18048,N_17210,N_17615);
nand U18049 (N_18049,N_17602,N_17669);
nor U18050 (N_18050,N_17710,N_17942);
xor U18051 (N_18051,N_17215,N_17943);
nand U18052 (N_18052,N_17473,N_17551);
nand U18053 (N_18053,N_17331,N_17447);
xnor U18054 (N_18054,N_17552,N_17423);
and U18055 (N_18055,N_17161,N_17678);
nor U18056 (N_18056,N_17601,N_17801);
or U18057 (N_18057,N_17366,N_17809);
and U18058 (N_18058,N_17604,N_17759);
nand U18059 (N_18059,N_17566,N_17687);
or U18060 (N_18060,N_17610,N_17505);
xor U18061 (N_18061,N_17689,N_17677);
xor U18062 (N_18062,N_17075,N_17957);
or U18063 (N_18063,N_17702,N_17170);
nor U18064 (N_18064,N_17246,N_17421);
nor U18065 (N_18065,N_17693,N_17490);
nor U18066 (N_18066,N_17033,N_17929);
nand U18067 (N_18067,N_17402,N_17907);
and U18068 (N_18068,N_17503,N_17354);
xnor U18069 (N_18069,N_17115,N_17003);
nand U18070 (N_18070,N_17525,N_17729);
nor U18071 (N_18071,N_17150,N_17914);
or U18072 (N_18072,N_17934,N_17818);
nor U18073 (N_18073,N_17675,N_17144);
and U18074 (N_18074,N_17475,N_17046);
and U18075 (N_18075,N_17961,N_17828);
and U18076 (N_18076,N_17206,N_17108);
nand U18077 (N_18077,N_17509,N_17103);
nand U18078 (N_18078,N_17999,N_17890);
xnor U18079 (N_18079,N_17200,N_17699);
nand U18080 (N_18080,N_17931,N_17294);
nor U18081 (N_18081,N_17691,N_17293);
and U18082 (N_18082,N_17531,N_17084);
nand U18083 (N_18083,N_17291,N_17718);
or U18084 (N_18084,N_17893,N_17586);
nand U18085 (N_18085,N_17825,N_17134);
nand U18086 (N_18086,N_17695,N_17635);
nor U18087 (N_18087,N_17792,N_17982);
and U18088 (N_18088,N_17029,N_17494);
xnor U18089 (N_18089,N_17268,N_17079);
nor U18090 (N_18090,N_17905,N_17499);
or U18091 (N_18091,N_17761,N_17676);
nor U18092 (N_18092,N_17372,N_17863);
nand U18093 (N_18093,N_17478,N_17032);
nor U18094 (N_18094,N_17590,N_17406);
nand U18095 (N_18095,N_17043,N_17674);
nand U18096 (N_18096,N_17751,N_17212);
and U18097 (N_18097,N_17576,N_17577);
or U18098 (N_18098,N_17508,N_17178);
and U18099 (N_18099,N_17168,N_17411);
or U18100 (N_18100,N_17724,N_17516);
and U18101 (N_18101,N_17884,N_17741);
nand U18102 (N_18102,N_17472,N_17328);
xor U18103 (N_18103,N_17017,N_17336);
nor U18104 (N_18104,N_17063,N_17995);
xnor U18105 (N_18105,N_17603,N_17870);
xor U18106 (N_18106,N_17238,N_17468);
nand U18107 (N_18107,N_17522,N_17706);
nand U18108 (N_18108,N_17569,N_17984);
nand U18109 (N_18109,N_17944,N_17764);
nand U18110 (N_18110,N_17184,N_17380);
nand U18111 (N_18111,N_17424,N_17073);
or U18112 (N_18112,N_17644,N_17098);
nand U18113 (N_18113,N_17524,N_17933);
xnor U18114 (N_18114,N_17393,N_17580);
nor U18115 (N_18115,N_17530,N_17437);
nor U18116 (N_18116,N_17371,N_17172);
nand U18117 (N_18117,N_17449,N_17128);
and U18118 (N_18118,N_17790,N_17864);
nor U18119 (N_18119,N_17422,N_17085);
nor U18120 (N_18120,N_17105,N_17429);
nor U18121 (N_18121,N_17182,N_17810);
nand U18122 (N_18122,N_17344,N_17841);
and U18123 (N_18123,N_17688,N_17175);
nand U18124 (N_18124,N_17425,N_17097);
xnor U18125 (N_18125,N_17658,N_17129);
nand U18126 (N_18126,N_17117,N_17978);
nor U18127 (N_18127,N_17089,N_17339);
or U18128 (N_18128,N_17474,N_17747);
xnor U18129 (N_18129,N_17131,N_17302);
nand U18130 (N_18130,N_17964,N_17805);
nor U18131 (N_18131,N_17510,N_17395);
nor U18132 (N_18132,N_17428,N_17697);
nand U18133 (N_18133,N_17323,N_17091);
and U18134 (N_18134,N_17655,N_17002);
or U18135 (N_18135,N_17426,N_17376);
xor U18136 (N_18136,N_17186,N_17616);
nand U18137 (N_18137,N_17039,N_17920);
xnor U18138 (N_18138,N_17231,N_17740);
nor U18139 (N_18139,N_17058,N_17278);
nor U18140 (N_18140,N_17885,N_17081);
nor U18141 (N_18141,N_17628,N_17584);
nor U18142 (N_18142,N_17936,N_17082);
nand U18143 (N_18143,N_17501,N_17322);
xnor U18144 (N_18144,N_17883,N_17318);
or U18145 (N_18145,N_17972,N_17317);
nor U18146 (N_18146,N_17194,N_17201);
or U18147 (N_18147,N_17433,N_17773);
xnor U18148 (N_18148,N_17756,N_17630);
nand U18149 (N_18149,N_17027,N_17660);
or U18150 (N_18150,N_17403,N_17946);
and U18151 (N_18151,N_17381,N_17162);
nor U18152 (N_18152,N_17815,N_17517);
nand U18153 (N_18153,N_17557,N_17151);
xor U18154 (N_18154,N_17225,N_17641);
or U18155 (N_18155,N_17672,N_17263);
xnor U18156 (N_18156,N_17913,N_17319);
and U18157 (N_18157,N_17585,N_17698);
nand U18158 (N_18158,N_17176,N_17589);
xnor U18159 (N_18159,N_17917,N_17645);
nand U18160 (N_18160,N_17703,N_17252);
or U18161 (N_18161,N_17374,N_17550);
and U18162 (N_18162,N_17044,N_17442);
nor U18163 (N_18163,N_17080,N_17975);
nand U18164 (N_18164,N_17992,N_17014);
nand U18165 (N_18165,N_17141,N_17363);
nand U18166 (N_18166,N_17991,N_17351);
xor U18167 (N_18167,N_17617,N_17096);
or U18168 (N_18168,N_17872,N_17357);
nor U18169 (N_18169,N_17048,N_17036);
and U18170 (N_18170,N_17731,N_17812);
xnor U18171 (N_18171,N_17065,N_17904);
xnor U18172 (N_18172,N_17989,N_17770);
or U18173 (N_18173,N_17078,N_17056);
or U18174 (N_18174,N_17420,N_17732);
xor U18175 (N_18175,N_17835,N_17070);
or U18176 (N_18176,N_17345,N_17607);
or U18177 (N_18177,N_17664,N_17343);
nand U18178 (N_18178,N_17611,N_17918);
nand U18179 (N_18179,N_17409,N_17249);
and U18180 (N_18180,N_17859,N_17389);
and U18181 (N_18181,N_17754,N_17774);
nor U18182 (N_18182,N_17137,N_17633);
and U18183 (N_18183,N_17763,N_17988);
and U18184 (N_18184,N_17071,N_17247);
and U18185 (N_18185,N_17391,N_17035);
or U18186 (N_18186,N_17894,N_17205);
and U18187 (N_18187,N_17460,N_17518);
or U18188 (N_18188,N_17515,N_17000);
nor U18189 (N_18189,N_17945,N_17998);
xor U18190 (N_18190,N_17836,N_17434);
xor U18191 (N_18191,N_17020,N_17368);
and U18192 (N_18192,N_17537,N_17970);
nor U18193 (N_18193,N_17412,N_17234);
nand U18194 (N_18194,N_17207,N_17237);
and U18195 (N_18195,N_17459,N_17310);
xnor U18196 (N_18196,N_17148,N_17275);
or U18197 (N_18197,N_17983,N_17634);
and U18198 (N_18198,N_17004,N_17692);
nor U18199 (N_18199,N_17288,N_17649);
and U18200 (N_18200,N_17221,N_17383);
or U18201 (N_18201,N_17867,N_17514);
or U18202 (N_18202,N_17414,N_17780);
nand U18203 (N_18203,N_17396,N_17193);
nor U18204 (N_18204,N_17730,N_17683);
and U18205 (N_18205,N_17037,N_17903);
and U18206 (N_18206,N_17049,N_17976);
xnor U18207 (N_18207,N_17297,N_17558);
and U18208 (N_18208,N_17820,N_17852);
nand U18209 (N_18209,N_17100,N_17259);
and U18210 (N_18210,N_17582,N_17857);
nand U18211 (N_18211,N_17267,N_17019);
nor U18212 (N_18212,N_17637,N_17847);
xor U18213 (N_18213,N_17378,N_17869);
or U18214 (N_18214,N_17753,N_17532);
nor U18215 (N_18215,N_17315,N_17572);
xnor U18216 (N_18216,N_17189,N_17654);
or U18217 (N_18217,N_17722,N_17120);
nor U18218 (N_18218,N_17147,N_17132);
nand U18219 (N_18219,N_17799,N_17018);
or U18220 (N_18220,N_17296,N_17384);
xnor U18221 (N_18221,N_17568,N_17821);
and U18222 (N_18222,N_17778,N_17456);
nand U18223 (N_18223,N_17123,N_17928);
nor U18224 (N_18224,N_17229,N_17896);
and U18225 (N_18225,N_17717,N_17307);
nor U18226 (N_18226,N_17882,N_17276);
nor U18227 (N_18227,N_17900,N_17118);
nor U18228 (N_18228,N_17031,N_17122);
or U18229 (N_18229,N_17377,N_17632);
nand U18230 (N_18230,N_17696,N_17335);
and U18231 (N_18231,N_17057,N_17289);
and U18232 (N_18232,N_17846,N_17614);
nor U18233 (N_18233,N_17832,N_17042);
xor U18234 (N_18234,N_17199,N_17090);
nor U18235 (N_18235,N_17140,N_17179);
or U18236 (N_18236,N_17369,N_17316);
xor U18237 (N_18237,N_17578,N_17909);
and U18238 (N_18238,N_17116,N_17155);
or U18239 (N_18239,N_17274,N_17880);
or U18240 (N_18240,N_17666,N_17496);
and U18241 (N_18241,N_17492,N_17748);
xnor U18242 (N_18242,N_17230,N_17668);
nor U18243 (N_18243,N_17016,N_17145);
and U18244 (N_18244,N_17862,N_17837);
xnor U18245 (N_18245,N_17023,N_17538);
xnor U18246 (N_18246,N_17670,N_17375);
nor U18247 (N_18247,N_17489,N_17171);
nand U18248 (N_18248,N_17618,N_17605);
nand U18249 (N_18249,N_17777,N_17979);
and U18250 (N_18250,N_17427,N_17413);
or U18251 (N_18251,N_17401,N_17854);
or U18252 (N_18252,N_17111,N_17648);
nor U18253 (N_18253,N_17416,N_17897);
xnor U18254 (N_18254,N_17977,N_17776);
nor U18255 (N_18255,N_17255,N_17910);
xnor U18256 (N_18256,N_17269,N_17581);
nand U18257 (N_18257,N_17143,N_17797);
and U18258 (N_18258,N_17352,N_17966);
or U18259 (N_18259,N_17481,N_17311);
or U18260 (N_18260,N_17919,N_17888);
nand U18261 (N_18261,N_17153,N_17453);
xor U18262 (N_18262,N_17823,N_17922);
or U18263 (N_18263,N_17507,N_17653);
and U18264 (N_18264,N_17925,N_17962);
nand U18265 (N_18265,N_17824,N_17520);
or U18266 (N_18266,N_17831,N_17270);
and U18267 (N_18267,N_17665,N_17448);
and U18268 (N_18268,N_17497,N_17930);
nand U18269 (N_18269,N_17723,N_17198);
xor U18270 (N_18270,N_17713,N_17295);
xnor U18271 (N_18271,N_17298,N_17892);
nand U18272 (N_18272,N_17768,N_17177);
or U18273 (N_18273,N_17842,N_17921);
xnor U18274 (N_18274,N_17785,N_17871);
xor U18275 (N_18275,N_17860,N_17591);
xnor U18276 (N_18276,N_17593,N_17483);
nor U18277 (N_18277,N_17849,N_17012);
nor U18278 (N_18278,N_17054,N_17087);
xor U18279 (N_18279,N_17196,N_17993);
or U18280 (N_18280,N_17938,N_17370);
or U18281 (N_18281,N_17498,N_17734);
nor U18282 (N_18282,N_17454,N_17300);
xor U18283 (N_18283,N_17908,N_17673);
nand U18284 (N_18284,N_17347,N_17158);
nor U18285 (N_18285,N_17619,N_17099);
and U18286 (N_18286,N_17542,N_17963);
xor U18287 (N_18287,N_17721,N_17226);
and U18288 (N_18288,N_17804,N_17535);
xnor U18289 (N_18289,N_17387,N_17450);
nor U18290 (N_18290,N_17061,N_17671);
xnor U18291 (N_18291,N_17681,N_17802);
xor U18292 (N_18292,N_17996,N_17588);
nand U18293 (N_18293,N_17879,N_17047);
and U18294 (N_18294,N_17359,N_17325);
or U18295 (N_18295,N_17495,N_17320);
nor U18296 (N_18296,N_17239,N_17114);
nand U18297 (N_18297,N_17292,N_17465);
nand U18298 (N_18298,N_17102,N_17109);
or U18299 (N_18299,N_17877,N_17651);
and U18300 (N_18300,N_17545,N_17197);
or U18301 (N_18301,N_17912,N_17562);
nor U18302 (N_18302,N_17088,N_17822);
xnor U18303 (N_18303,N_17445,N_17573);
and U18304 (N_18304,N_17874,N_17388);
or U18305 (N_18305,N_17549,N_17482);
nand U18306 (N_18306,N_17959,N_17981);
xor U18307 (N_18307,N_17858,N_17216);
and U18308 (N_18308,N_17733,N_17891);
and U18309 (N_18309,N_17001,N_17139);
or U18310 (N_18310,N_17807,N_17640);
nor U18311 (N_18311,N_17887,N_17844);
or U18312 (N_18312,N_17939,N_17500);
nand U18313 (N_18313,N_17701,N_17303);
nand U18314 (N_18314,N_17220,N_17783);
nor U18315 (N_18315,N_17800,N_17597);
nand U18316 (N_18316,N_17365,N_17985);
xor U18317 (N_18317,N_17694,N_17620);
and U18318 (N_18318,N_17142,N_17861);
and U18319 (N_18319,N_17690,N_17742);
and U18320 (N_18320,N_17779,N_17355);
or U18321 (N_18321,N_17159,N_17462);
nand U18322 (N_18322,N_17901,N_17332);
nor U18323 (N_18323,N_17192,N_17219);
nand U18324 (N_18324,N_17881,N_17301);
or U18325 (N_18325,N_17166,N_17390);
xnor U18326 (N_18326,N_17028,N_17621);
nor U18327 (N_18327,N_17609,N_17362);
and U18328 (N_18328,N_17541,N_17299);
xor U18329 (N_18329,N_17261,N_17488);
and U18330 (N_18330,N_17808,N_17364);
xnor U18331 (N_18331,N_17138,N_17766);
and U18332 (N_18332,N_17803,N_17479);
and U18333 (N_18333,N_17127,N_17232);
nand U18334 (N_18334,N_17485,N_17556);
and U18335 (N_18335,N_17181,N_17560);
or U18336 (N_18336,N_17030,N_17160);
nand U18337 (N_18337,N_17010,N_17283);
xor U18338 (N_18338,N_17466,N_17548);
xnor U18339 (N_18339,N_17650,N_17272);
nand U18340 (N_18340,N_17539,N_17521);
nor U18341 (N_18341,N_17873,N_17284);
and U18342 (N_18342,N_17180,N_17106);
nand U18343 (N_18343,N_17682,N_17266);
nor U18344 (N_18344,N_17379,N_17072);
nor U18345 (N_18345,N_17021,N_17817);
nand U18346 (N_18346,N_17540,N_17714);
nand U18347 (N_18347,N_17157,N_17022);
and U18348 (N_18348,N_17868,N_17257);
and U18349 (N_18349,N_17165,N_17191);
nand U18350 (N_18350,N_17636,N_17720);
xor U18351 (N_18351,N_17506,N_17523);
xor U18352 (N_18352,N_17949,N_17646);
nand U18353 (N_18353,N_17045,N_17543);
nor U18354 (N_18354,N_17313,N_17187);
or U18355 (N_18355,N_17055,N_17185);
nand U18356 (N_18356,N_17736,N_17994);
nor U18357 (N_18357,N_17241,N_17712);
nor U18358 (N_18358,N_17726,N_17725);
nor U18359 (N_18359,N_17680,N_17008);
and U18360 (N_18360,N_17074,N_17765);
and U18361 (N_18361,N_17631,N_17217);
nand U18362 (N_18362,N_17789,N_17554);
nor U18363 (N_18363,N_17243,N_17575);
xor U18364 (N_18364,N_17290,N_17544);
and U18365 (N_18365,N_17419,N_17309);
nor U18366 (N_18366,N_17086,N_17813);
and U18367 (N_18367,N_17130,N_17348);
and U18368 (N_18368,N_17271,N_17728);
or U18369 (N_18369,N_17613,N_17277);
or U18370 (N_18370,N_17125,N_17647);
xor U18371 (N_18371,N_17608,N_17798);
nor U18372 (N_18372,N_17895,N_17470);
or U18373 (N_18373,N_17059,N_17850);
xor U18374 (N_18374,N_17504,N_17005);
or U18375 (N_18375,N_17337,N_17902);
and U18376 (N_18376,N_17571,N_17679);
or U18377 (N_18377,N_17772,N_17211);
or U18378 (N_18378,N_17561,N_17547);
nand U18379 (N_18379,N_17104,N_17969);
nand U18380 (N_18380,N_17092,N_17856);
and U18381 (N_18381,N_17321,N_17947);
or U18382 (N_18382,N_17285,N_17464);
nand U18383 (N_18383,N_17987,N_17218);
or U18384 (N_18384,N_17242,N_17853);
nor U18385 (N_18385,N_17974,N_17526);
nor U18386 (N_18386,N_17851,N_17408);
xor U18387 (N_18387,N_17559,N_17173);
or U18388 (N_18388,N_17816,N_17353);
and U18389 (N_18389,N_17306,N_17980);
or U18390 (N_18390,N_17711,N_17038);
xnor U18391 (N_18391,N_17952,N_17112);
xnor U18392 (N_18392,N_17349,N_17625);
nor U18393 (N_18393,N_17843,N_17898);
and U18394 (N_18394,N_17791,N_17051);
or U18395 (N_18395,N_17567,N_17458);
xnor U18396 (N_18396,N_17467,N_17040);
xor U18397 (N_18397,N_17762,N_17746);
xnor U18398 (N_18398,N_17596,N_17360);
and U18399 (N_18399,N_17262,N_17062);
and U18400 (N_18400,N_17164,N_17067);
and U18401 (N_18401,N_17960,N_17064);
and U18402 (N_18402,N_17052,N_17011);
xor U18403 (N_18403,N_17154,N_17967);
or U18404 (N_18404,N_17382,N_17916);
or U18405 (N_18405,N_17417,N_17471);
and U18406 (N_18406,N_17410,N_17405);
and U18407 (N_18407,N_17188,N_17553);
nand U18408 (N_18408,N_17441,N_17958);
nor U18409 (N_18409,N_17415,N_17167);
and U18410 (N_18410,N_17737,N_17889);
and U18411 (N_18411,N_17076,N_17829);
xnor U18412 (N_18412,N_17627,N_17397);
nand U18413 (N_18413,N_17386,N_17656);
nor U18414 (N_18414,N_17926,N_17662);
nor U18415 (N_18415,N_17124,N_17997);
nand U18416 (N_18416,N_17156,N_17487);
nand U18417 (N_18417,N_17767,N_17624);
or U18418 (N_18418,N_17418,N_17511);
xor U18419 (N_18419,N_17899,N_17626);
xnor U18420 (N_18420,N_17659,N_17838);
nor U18421 (N_18421,N_17202,N_17121);
nand U18422 (N_18422,N_17579,N_17050);
nand U18423 (N_18423,N_17830,N_17373);
and U18424 (N_18424,N_17436,N_17053);
or U18425 (N_18425,N_17399,N_17404);
nand U18426 (N_18426,N_17806,N_17760);
xnor U18427 (N_18427,N_17749,N_17583);
xnor U18428 (N_18428,N_17227,N_17755);
or U18429 (N_18429,N_17093,N_17923);
nor U18430 (N_18430,N_17305,N_17439);
and U18431 (N_18431,N_17533,N_17430);
and U18432 (N_18432,N_17358,N_17623);
nor U18433 (N_18433,N_17811,N_17932);
and U18434 (N_18434,N_17287,N_17529);
or U18435 (N_18435,N_17444,N_17705);
nor U18436 (N_18436,N_17457,N_17350);
nor U18437 (N_18437,N_17330,N_17709);
or U18438 (N_18438,N_17565,N_17110);
or U18439 (N_18439,N_17204,N_17727);
or U18440 (N_18440,N_17574,N_17512);
or U18441 (N_18441,N_17025,N_17245);
and U18442 (N_18442,N_17095,N_17528);
xnor U18443 (N_18443,N_17435,N_17781);
or U18444 (N_18444,N_17240,N_17312);
and U18445 (N_18445,N_17840,N_17570);
or U18446 (N_18446,N_17346,N_17385);
nor U18447 (N_18447,N_17786,N_17066);
and U18448 (N_18448,N_17214,N_17341);
or U18449 (N_18449,N_17744,N_17264);
xor U18450 (N_18450,N_17327,N_17367);
and U18451 (N_18451,N_17174,N_17954);
nor U18452 (N_18452,N_17715,N_17638);
xnor U18453 (N_18453,N_17041,N_17235);
nor U18454 (N_18454,N_17911,N_17392);
nand U18455 (N_18455,N_17782,N_17950);
or U18456 (N_18456,N_17431,N_17203);
and U18457 (N_18457,N_17855,N_17356);
nand U18458 (N_18458,N_17757,N_17814);
xor U18459 (N_18459,N_17333,N_17927);
xor U18460 (N_18460,N_17513,N_17795);
nor U18461 (N_18461,N_17700,N_17407);
or U18462 (N_18462,N_17493,N_17827);
xor U18463 (N_18463,N_17491,N_17948);
or U18464 (N_18464,N_17248,N_17486);
xor U18465 (N_18465,N_17739,N_17771);
or U18466 (N_18466,N_17990,N_17704);
or U18467 (N_18467,N_17622,N_17236);
nor U18468 (N_18468,N_17477,N_17788);
nor U18469 (N_18469,N_17163,N_17965);
nor U18470 (N_18470,N_17546,N_17273);
or U18471 (N_18471,N_17527,N_17735);
and U18472 (N_18472,N_17443,N_17661);
nand U18473 (N_18473,N_17955,N_17937);
or U18474 (N_18474,N_17400,N_17865);
nand U18475 (N_18475,N_17209,N_17452);
nor U18476 (N_18476,N_17222,N_17639);
or U18477 (N_18477,N_17793,N_17973);
or U18478 (N_18478,N_17643,N_17685);
xor U18479 (N_18479,N_17326,N_17107);
and U18480 (N_18480,N_17968,N_17758);
and U18481 (N_18481,N_17642,N_17228);
xor U18482 (N_18482,N_17555,N_17026);
xnor U18483 (N_18483,N_17956,N_17536);
and U18484 (N_18484,N_17015,N_17480);
nand U18485 (N_18485,N_17629,N_17304);
nand U18486 (N_18486,N_17612,N_17886);
or U18487 (N_18487,N_17455,N_17599);
or U18488 (N_18488,N_17971,N_17986);
nor U18489 (N_18489,N_17667,N_17256);
nor U18490 (N_18490,N_17833,N_17334);
nor U18491 (N_18491,N_17463,N_17432);
nand U18492 (N_18492,N_17253,N_17686);
nand U18493 (N_18493,N_17324,N_17169);
and U18494 (N_18494,N_17461,N_17866);
and U18495 (N_18495,N_17935,N_17915);
nand U18496 (N_18496,N_17600,N_17875);
and U18497 (N_18497,N_17034,N_17126);
xnor U18498 (N_18498,N_17587,N_17149);
and U18499 (N_18499,N_17254,N_17183);
nor U18500 (N_18500,N_17198,N_17185);
xnor U18501 (N_18501,N_17564,N_17189);
or U18502 (N_18502,N_17344,N_17937);
and U18503 (N_18503,N_17815,N_17198);
xnor U18504 (N_18504,N_17540,N_17465);
or U18505 (N_18505,N_17307,N_17950);
or U18506 (N_18506,N_17338,N_17243);
nand U18507 (N_18507,N_17716,N_17718);
xor U18508 (N_18508,N_17448,N_17161);
xnor U18509 (N_18509,N_17273,N_17625);
nor U18510 (N_18510,N_17006,N_17069);
xor U18511 (N_18511,N_17778,N_17328);
and U18512 (N_18512,N_17908,N_17487);
and U18513 (N_18513,N_17156,N_17832);
nor U18514 (N_18514,N_17891,N_17600);
or U18515 (N_18515,N_17831,N_17743);
nor U18516 (N_18516,N_17871,N_17930);
and U18517 (N_18517,N_17043,N_17225);
or U18518 (N_18518,N_17904,N_17175);
xor U18519 (N_18519,N_17938,N_17726);
nand U18520 (N_18520,N_17099,N_17193);
xnor U18521 (N_18521,N_17858,N_17342);
nand U18522 (N_18522,N_17315,N_17333);
or U18523 (N_18523,N_17131,N_17498);
xor U18524 (N_18524,N_17166,N_17629);
xnor U18525 (N_18525,N_17110,N_17134);
and U18526 (N_18526,N_17118,N_17933);
or U18527 (N_18527,N_17018,N_17838);
nor U18528 (N_18528,N_17592,N_17598);
or U18529 (N_18529,N_17382,N_17667);
nand U18530 (N_18530,N_17877,N_17464);
nor U18531 (N_18531,N_17754,N_17122);
xnor U18532 (N_18532,N_17875,N_17683);
xor U18533 (N_18533,N_17502,N_17442);
xor U18534 (N_18534,N_17789,N_17639);
xor U18535 (N_18535,N_17577,N_17813);
xnor U18536 (N_18536,N_17631,N_17763);
nand U18537 (N_18537,N_17495,N_17908);
or U18538 (N_18538,N_17092,N_17812);
nand U18539 (N_18539,N_17011,N_17049);
nand U18540 (N_18540,N_17670,N_17459);
or U18541 (N_18541,N_17517,N_17244);
or U18542 (N_18542,N_17458,N_17885);
nand U18543 (N_18543,N_17003,N_17767);
xnor U18544 (N_18544,N_17626,N_17736);
or U18545 (N_18545,N_17616,N_17629);
or U18546 (N_18546,N_17810,N_17369);
and U18547 (N_18547,N_17789,N_17934);
xnor U18548 (N_18548,N_17320,N_17209);
xor U18549 (N_18549,N_17861,N_17338);
xor U18550 (N_18550,N_17196,N_17902);
and U18551 (N_18551,N_17377,N_17586);
or U18552 (N_18552,N_17434,N_17764);
xnor U18553 (N_18553,N_17747,N_17139);
nand U18554 (N_18554,N_17626,N_17723);
nor U18555 (N_18555,N_17596,N_17299);
xnor U18556 (N_18556,N_17668,N_17761);
nand U18557 (N_18557,N_17376,N_17614);
or U18558 (N_18558,N_17757,N_17340);
and U18559 (N_18559,N_17581,N_17965);
nor U18560 (N_18560,N_17649,N_17324);
and U18561 (N_18561,N_17714,N_17375);
nor U18562 (N_18562,N_17809,N_17348);
nand U18563 (N_18563,N_17371,N_17288);
nor U18564 (N_18564,N_17601,N_17190);
nand U18565 (N_18565,N_17520,N_17587);
xnor U18566 (N_18566,N_17178,N_17477);
and U18567 (N_18567,N_17494,N_17505);
nand U18568 (N_18568,N_17736,N_17577);
xnor U18569 (N_18569,N_17301,N_17970);
and U18570 (N_18570,N_17078,N_17556);
and U18571 (N_18571,N_17564,N_17639);
xnor U18572 (N_18572,N_17898,N_17005);
or U18573 (N_18573,N_17004,N_17848);
and U18574 (N_18574,N_17034,N_17209);
nand U18575 (N_18575,N_17496,N_17485);
and U18576 (N_18576,N_17646,N_17049);
or U18577 (N_18577,N_17455,N_17030);
and U18578 (N_18578,N_17597,N_17383);
nor U18579 (N_18579,N_17685,N_17547);
xnor U18580 (N_18580,N_17589,N_17362);
xnor U18581 (N_18581,N_17252,N_17174);
xor U18582 (N_18582,N_17206,N_17032);
or U18583 (N_18583,N_17360,N_17507);
nor U18584 (N_18584,N_17905,N_17410);
nor U18585 (N_18585,N_17722,N_17845);
xor U18586 (N_18586,N_17433,N_17317);
xor U18587 (N_18587,N_17507,N_17325);
and U18588 (N_18588,N_17860,N_17500);
xnor U18589 (N_18589,N_17644,N_17802);
and U18590 (N_18590,N_17562,N_17168);
or U18591 (N_18591,N_17313,N_17375);
xor U18592 (N_18592,N_17169,N_17775);
xnor U18593 (N_18593,N_17986,N_17267);
nand U18594 (N_18594,N_17805,N_17920);
nand U18595 (N_18595,N_17211,N_17215);
nand U18596 (N_18596,N_17793,N_17397);
nor U18597 (N_18597,N_17388,N_17093);
nor U18598 (N_18598,N_17630,N_17313);
or U18599 (N_18599,N_17457,N_17065);
nor U18600 (N_18600,N_17066,N_17903);
nor U18601 (N_18601,N_17561,N_17509);
nand U18602 (N_18602,N_17524,N_17002);
and U18603 (N_18603,N_17396,N_17203);
and U18604 (N_18604,N_17941,N_17561);
xnor U18605 (N_18605,N_17353,N_17439);
nand U18606 (N_18606,N_17689,N_17230);
nand U18607 (N_18607,N_17778,N_17047);
nor U18608 (N_18608,N_17612,N_17544);
and U18609 (N_18609,N_17399,N_17427);
xnor U18610 (N_18610,N_17669,N_17453);
xor U18611 (N_18611,N_17079,N_17531);
nor U18612 (N_18612,N_17485,N_17471);
xor U18613 (N_18613,N_17694,N_17036);
xnor U18614 (N_18614,N_17794,N_17112);
nor U18615 (N_18615,N_17817,N_17959);
nor U18616 (N_18616,N_17058,N_17110);
nand U18617 (N_18617,N_17881,N_17718);
and U18618 (N_18618,N_17560,N_17766);
nor U18619 (N_18619,N_17748,N_17375);
or U18620 (N_18620,N_17299,N_17654);
or U18621 (N_18621,N_17155,N_17745);
nand U18622 (N_18622,N_17291,N_17676);
nand U18623 (N_18623,N_17714,N_17217);
and U18624 (N_18624,N_17003,N_17328);
xor U18625 (N_18625,N_17761,N_17601);
nor U18626 (N_18626,N_17633,N_17038);
nand U18627 (N_18627,N_17240,N_17681);
and U18628 (N_18628,N_17505,N_17947);
and U18629 (N_18629,N_17045,N_17424);
nor U18630 (N_18630,N_17893,N_17037);
or U18631 (N_18631,N_17078,N_17234);
or U18632 (N_18632,N_17445,N_17766);
xnor U18633 (N_18633,N_17657,N_17036);
and U18634 (N_18634,N_17390,N_17966);
nor U18635 (N_18635,N_17840,N_17165);
and U18636 (N_18636,N_17471,N_17966);
nor U18637 (N_18637,N_17541,N_17295);
or U18638 (N_18638,N_17945,N_17588);
xor U18639 (N_18639,N_17943,N_17395);
xor U18640 (N_18640,N_17661,N_17919);
nor U18641 (N_18641,N_17212,N_17487);
nand U18642 (N_18642,N_17950,N_17989);
xnor U18643 (N_18643,N_17583,N_17986);
xor U18644 (N_18644,N_17332,N_17217);
nand U18645 (N_18645,N_17038,N_17708);
or U18646 (N_18646,N_17022,N_17016);
nand U18647 (N_18647,N_17207,N_17141);
or U18648 (N_18648,N_17672,N_17164);
nor U18649 (N_18649,N_17665,N_17428);
or U18650 (N_18650,N_17507,N_17246);
xnor U18651 (N_18651,N_17779,N_17530);
or U18652 (N_18652,N_17907,N_17231);
and U18653 (N_18653,N_17548,N_17777);
nor U18654 (N_18654,N_17721,N_17926);
and U18655 (N_18655,N_17400,N_17090);
and U18656 (N_18656,N_17908,N_17951);
nand U18657 (N_18657,N_17455,N_17546);
nand U18658 (N_18658,N_17367,N_17582);
or U18659 (N_18659,N_17690,N_17803);
and U18660 (N_18660,N_17459,N_17339);
xnor U18661 (N_18661,N_17213,N_17767);
nand U18662 (N_18662,N_17815,N_17200);
and U18663 (N_18663,N_17674,N_17999);
nor U18664 (N_18664,N_17289,N_17969);
nor U18665 (N_18665,N_17600,N_17394);
or U18666 (N_18666,N_17439,N_17328);
or U18667 (N_18667,N_17537,N_17289);
nand U18668 (N_18668,N_17915,N_17652);
or U18669 (N_18669,N_17213,N_17873);
nor U18670 (N_18670,N_17874,N_17967);
xor U18671 (N_18671,N_17593,N_17061);
nor U18672 (N_18672,N_17282,N_17824);
xnor U18673 (N_18673,N_17756,N_17738);
nand U18674 (N_18674,N_17087,N_17197);
or U18675 (N_18675,N_17152,N_17415);
or U18676 (N_18676,N_17749,N_17967);
xnor U18677 (N_18677,N_17115,N_17903);
nand U18678 (N_18678,N_17216,N_17407);
nand U18679 (N_18679,N_17613,N_17902);
or U18680 (N_18680,N_17648,N_17972);
and U18681 (N_18681,N_17579,N_17862);
and U18682 (N_18682,N_17702,N_17371);
nor U18683 (N_18683,N_17243,N_17099);
xnor U18684 (N_18684,N_17949,N_17682);
or U18685 (N_18685,N_17123,N_17143);
nand U18686 (N_18686,N_17201,N_17603);
and U18687 (N_18687,N_17409,N_17086);
xnor U18688 (N_18688,N_17792,N_17679);
nand U18689 (N_18689,N_17562,N_17272);
or U18690 (N_18690,N_17581,N_17229);
xor U18691 (N_18691,N_17980,N_17694);
xnor U18692 (N_18692,N_17693,N_17178);
nand U18693 (N_18693,N_17422,N_17430);
and U18694 (N_18694,N_17610,N_17111);
nor U18695 (N_18695,N_17068,N_17748);
nand U18696 (N_18696,N_17290,N_17942);
nand U18697 (N_18697,N_17903,N_17751);
nand U18698 (N_18698,N_17907,N_17734);
and U18699 (N_18699,N_17484,N_17305);
xor U18700 (N_18700,N_17141,N_17619);
nor U18701 (N_18701,N_17757,N_17813);
nand U18702 (N_18702,N_17678,N_17961);
xnor U18703 (N_18703,N_17813,N_17835);
nand U18704 (N_18704,N_17487,N_17939);
or U18705 (N_18705,N_17721,N_17013);
xor U18706 (N_18706,N_17336,N_17722);
or U18707 (N_18707,N_17352,N_17464);
nand U18708 (N_18708,N_17353,N_17967);
nand U18709 (N_18709,N_17926,N_17421);
and U18710 (N_18710,N_17000,N_17984);
and U18711 (N_18711,N_17305,N_17281);
nand U18712 (N_18712,N_17246,N_17745);
nand U18713 (N_18713,N_17682,N_17852);
nand U18714 (N_18714,N_17193,N_17599);
and U18715 (N_18715,N_17927,N_17432);
xor U18716 (N_18716,N_17102,N_17475);
and U18717 (N_18717,N_17833,N_17016);
nor U18718 (N_18718,N_17382,N_17645);
nand U18719 (N_18719,N_17135,N_17763);
and U18720 (N_18720,N_17435,N_17128);
nand U18721 (N_18721,N_17472,N_17771);
xnor U18722 (N_18722,N_17356,N_17447);
xor U18723 (N_18723,N_17399,N_17209);
and U18724 (N_18724,N_17995,N_17390);
xor U18725 (N_18725,N_17076,N_17889);
nand U18726 (N_18726,N_17037,N_17481);
and U18727 (N_18727,N_17189,N_17355);
nand U18728 (N_18728,N_17654,N_17886);
xnor U18729 (N_18729,N_17444,N_17037);
nor U18730 (N_18730,N_17227,N_17152);
nand U18731 (N_18731,N_17827,N_17155);
and U18732 (N_18732,N_17541,N_17347);
or U18733 (N_18733,N_17583,N_17152);
nor U18734 (N_18734,N_17906,N_17553);
nor U18735 (N_18735,N_17977,N_17992);
nor U18736 (N_18736,N_17596,N_17129);
and U18737 (N_18737,N_17738,N_17542);
and U18738 (N_18738,N_17791,N_17851);
nand U18739 (N_18739,N_17147,N_17714);
nor U18740 (N_18740,N_17495,N_17818);
nor U18741 (N_18741,N_17502,N_17788);
and U18742 (N_18742,N_17173,N_17839);
nand U18743 (N_18743,N_17543,N_17598);
or U18744 (N_18744,N_17780,N_17247);
nor U18745 (N_18745,N_17071,N_17229);
or U18746 (N_18746,N_17732,N_17906);
xnor U18747 (N_18747,N_17742,N_17628);
and U18748 (N_18748,N_17644,N_17873);
or U18749 (N_18749,N_17870,N_17326);
or U18750 (N_18750,N_17000,N_17996);
or U18751 (N_18751,N_17854,N_17348);
nor U18752 (N_18752,N_17497,N_17241);
xor U18753 (N_18753,N_17212,N_17035);
xnor U18754 (N_18754,N_17077,N_17275);
xor U18755 (N_18755,N_17692,N_17643);
nor U18756 (N_18756,N_17930,N_17588);
nor U18757 (N_18757,N_17815,N_17896);
or U18758 (N_18758,N_17464,N_17330);
nand U18759 (N_18759,N_17463,N_17118);
nor U18760 (N_18760,N_17619,N_17130);
and U18761 (N_18761,N_17996,N_17648);
xor U18762 (N_18762,N_17862,N_17113);
nor U18763 (N_18763,N_17307,N_17687);
or U18764 (N_18764,N_17636,N_17911);
and U18765 (N_18765,N_17921,N_17806);
xor U18766 (N_18766,N_17892,N_17838);
nor U18767 (N_18767,N_17724,N_17939);
nor U18768 (N_18768,N_17599,N_17658);
nand U18769 (N_18769,N_17087,N_17479);
xnor U18770 (N_18770,N_17947,N_17197);
nor U18771 (N_18771,N_17549,N_17548);
nand U18772 (N_18772,N_17657,N_17221);
or U18773 (N_18773,N_17540,N_17546);
and U18774 (N_18774,N_17814,N_17013);
nor U18775 (N_18775,N_17825,N_17489);
xnor U18776 (N_18776,N_17423,N_17647);
nand U18777 (N_18777,N_17828,N_17113);
nand U18778 (N_18778,N_17613,N_17164);
nor U18779 (N_18779,N_17606,N_17291);
and U18780 (N_18780,N_17822,N_17612);
nand U18781 (N_18781,N_17503,N_17250);
and U18782 (N_18782,N_17203,N_17397);
xnor U18783 (N_18783,N_17159,N_17567);
nand U18784 (N_18784,N_17388,N_17345);
nand U18785 (N_18785,N_17829,N_17648);
or U18786 (N_18786,N_17801,N_17404);
and U18787 (N_18787,N_17256,N_17721);
xnor U18788 (N_18788,N_17355,N_17455);
or U18789 (N_18789,N_17573,N_17688);
xor U18790 (N_18790,N_17975,N_17310);
or U18791 (N_18791,N_17321,N_17801);
xor U18792 (N_18792,N_17098,N_17824);
nand U18793 (N_18793,N_17049,N_17896);
nor U18794 (N_18794,N_17468,N_17576);
or U18795 (N_18795,N_17665,N_17376);
nor U18796 (N_18796,N_17095,N_17954);
and U18797 (N_18797,N_17046,N_17985);
and U18798 (N_18798,N_17625,N_17466);
nand U18799 (N_18799,N_17323,N_17623);
or U18800 (N_18800,N_17645,N_17566);
xor U18801 (N_18801,N_17261,N_17166);
nand U18802 (N_18802,N_17922,N_17047);
nand U18803 (N_18803,N_17381,N_17729);
or U18804 (N_18804,N_17592,N_17350);
nand U18805 (N_18805,N_17218,N_17444);
nand U18806 (N_18806,N_17409,N_17666);
nor U18807 (N_18807,N_17351,N_17283);
nor U18808 (N_18808,N_17972,N_17337);
nand U18809 (N_18809,N_17255,N_17989);
or U18810 (N_18810,N_17817,N_17621);
and U18811 (N_18811,N_17390,N_17564);
nor U18812 (N_18812,N_17682,N_17887);
nor U18813 (N_18813,N_17893,N_17142);
and U18814 (N_18814,N_17005,N_17553);
or U18815 (N_18815,N_17383,N_17136);
and U18816 (N_18816,N_17675,N_17156);
or U18817 (N_18817,N_17427,N_17501);
or U18818 (N_18818,N_17790,N_17686);
or U18819 (N_18819,N_17328,N_17845);
or U18820 (N_18820,N_17546,N_17439);
or U18821 (N_18821,N_17608,N_17563);
or U18822 (N_18822,N_17124,N_17840);
nor U18823 (N_18823,N_17667,N_17109);
nand U18824 (N_18824,N_17099,N_17800);
xnor U18825 (N_18825,N_17945,N_17025);
nor U18826 (N_18826,N_17078,N_17620);
and U18827 (N_18827,N_17582,N_17314);
nand U18828 (N_18828,N_17397,N_17894);
xnor U18829 (N_18829,N_17279,N_17327);
nand U18830 (N_18830,N_17626,N_17944);
and U18831 (N_18831,N_17129,N_17506);
or U18832 (N_18832,N_17579,N_17612);
or U18833 (N_18833,N_17392,N_17967);
and U18834 (N_18834,N_17817,N_17274);
xor U18835 (N_18835,N_17485,N_17559);
or U18836 (N_18836,N_17532,N_17349);
and U18837 (N_18837,N_17453,N_17511);
and U18838 (N_18838,N_17483,N_17896);
nor U18839 (N_18839,N_17607,N_17744);
nor U18840 (N_18840,N_17715,N_17595);
and U18841 (N_18841,N_17427,N_17715);
and U18842 (N_18842,N_17120,N_17744);
nand U18843 (N_18843,N_17663,N_17631);
and U18844 (N_18844,N_17503,N_17797);
nor U18845 (N_18845,N_17100,N_17880);
nor U18846 (N_18846,N_17239,N_17042);
or U18847 (N_18847,N_17683,N_17743);
nand U18848 (N_18848,N_17338,N_17092);
xor U18849 (N_18849,N_17906,N_17247);
and U18850 (N_18850,N_17645,N_17780);
nand U18851 (N_18851,N_17785,N_17545);
and U18852 (N_18852,N_17370,N_17311);
or U18853 (N_18853,N_17691,N_17879);
nand U18854 (N_18854,N_17280,N_17625);
and U18855 (N_18855,N_17214,N_17547);
and U18856 (N_18856,N_17330,N_17166);
and U18857 (N_18857,N_17292,N_17551);
nand U18858 (N_18858,N_17929,N_17712);
and U18859 (N_18859,N_17913,N_17968);
xor U18860 (N_18860,N_17109,N_17411);
xnor U18861 (N_18861,N_17990,N_17477);
or U18862 (N_18862,N_17570,N_17770);
nand U18863 (N_18863,N_17548,N_17858);
nor U18864 (N_18864,N_17382,N_17346);
or U18865 (N_18865,N_17923,N_17655);
nand U18866 (N_18866,N_17663,N_17328);
or U18867 (N_18867,N_17747,N_17896);
nor U18868 (N_18868,N_17291,N_17158);
nor U18869 (N_18869,N_17647,N_17434);
xor U18870 (N_18870,N_17924,N_17063);
or U18871 (N_18871,N_17875,N_17571);
and U18872 (N_18872,N_17829,N_17263);
nor U18873 (N_18873,N_17965,N_17967);
or U18874 (N_18874,N_17057,N_17074);
nor U18875 (N_18875,N_17730,N_17675);
nand U18876 (N_18876,N_17316,N_17023);
and U18877 (N_18877,N_17039,N_17788);
or U18878 (N_18878,N_17938,N_17828);
xor U18879 (N_18879,N_17698,N_17442);
and U18880 (N_18880,N_17229,N_17262);
or U18881 (N_18881,N_17137,N_17523);
and U18882 (N_18882,N_17664,N_17468);
nand U18883 (N_18883,N_17675,N_17386);
and U18884 (N_18884,N_17172,N_17636);
nand U18885 (N_18885,N_17463,N_17483);
xnor U18886 (N_18886,N_17570,N_17278);
nand U18887 (N_18887,N_17069,N_17879);
nand U18888 (N_18888,N_17140,N_17490);
xnor U18889 (N_18889,N_17797,N_17401);
nor U18890 (N_18890,N_17374,N_17198);
nand U18891 (N_18891,N_17532,N_17281);
nand U18892 (N_18892,N_17799,N_17518);
and U18893 (N_18893,N_17690,N_17205);
nor U18894 (N_18894,N_17369,N_17541);
nor U18895 (N_18895,N_17543,N_17307);
and U18896 (N_18896,N_17770,N_17162);
and U18897 (N_18897,N_17396,N_17455);
and U18898 (N_18898,N_17174,N_17349);
or U18899 (N_18899,N_17216,N_17567);
xor U18900 (N_18900,N_17552,N_17417);
and U18901 (N_18901,N_17006,N_17561);
nor U18902 (N_18902,N_17658,N_17483);
xnor U18903 (N_18903,N_17705,N_17992);
xor U18904 (N_18904,N_17413,N_17142);
and U18905 (N_18905,N_17333,N_17928);
xor U18906 (N_18906,N_17979,N_17292);
xor U18907 (N_18907,N_17158,N_17900);
and U18908 (N_18908,N_17497,N_17898);
xnor U18909 (N_18909,N_17631,N_17230);
and U18910 (N_18910,N_17142,N_17286);
nor U18911 (N_18911,N_17479,N_17156);
nand U18912 (N_18912,N_17072,N_17946);
xnor U18913 (N_18913,N_17655,N_17009);
and U18914 (N_18914,N_17682,N_17826);
nor U18915 (N_18915,N_17938,N_17650);
or U18916 (N_18916,N_17739,N_17221);
or U18917 (N_18917,N_17479,N_17987);
nor U18918 (N_18918,N_17060,N_17959);
and U18919 (N_18919,N_17828,N_17140);
or U18920 (N_18920,N_17997,N_17117);
or U18921 (N_18921,N_17823,N_17153);
nand U18922 (N_18922,N_17193,N_17192);
or U18923 (N_18923,N_17665,N_17141);
or U18924 (N_18924,N_17948,N_17289);
nand U18925 (N_18925,N_17049,N_17110);
nand U18926 (N_18926,N_17591,N_17742);
and U18927 (N_18927,N_17653,N_17096);
nand U18928 (N_18928,N_17226,N_17349);
or U18929 (N_18929,N_17581,N_17752);
nor U18930 (N_18930,N_17409,N_17904);
xor U18931 (N_18931,N_17972,N_17900);
and U18932 (N_18932,N_17504,N_17865);
nor U18933 (N_18933,N_17500,N_17941);
nor U18934 (N_18934,N_17935,N_17913);
and U18935 (N_18935,N_17211,N_17937);
xor U18936 (N_18936,N_17838,N_17259);
nand U18937 (N_18937,N_17243,N_17361);
xor U18938 (N_18938,N_17690,N_17170);
nor U18939 (N_18939,N_17257,N_17063);
nor U18940 (N_18940,N_17394,N_17619);
and U18941 (N_18941,N_17789,N_17577);
xnor U18942 (N_18942,N_17492,N_17818);
and U18943 (N_18943,N_17984,N_17818);
or U18944 (N_18944,N_17153,N_17902);
and U18945 (N_18945,N_17980,N_17191);
nor U18946 (N_18946,N_17943,N_17504);
xor U18947 (N_18947,N_17520,N_17127);
or U18948 (N_18948,N_17830,N_17249);
or U18949 (N_18949,N_17204,N_17935);
xor U18950 (N_18950,N_17201,N_17003);
or U18951 (N_18951,N_17177,N_17143);
nor U18952 (N_18952,N_17088,N_17096);
or U18953 (N_18953,N_17201,N_17620);
nand U18954 (N_18954,N_17030,N_17741);
nand U18955 (N_18955,N_17270,N_17925);
or U18956 (N_18956,N_17767,N_17838);
xnor U18957 (N_18957,N_17926,N_17747);
xor U18958 (N_18958,N_17927,N_17261);
and U18959 (N_18959,N_17334,N_17809);
and U18960 (N_18960,N_17603,N_17339);
and U18961 (N_18961,N_17579,N_17501);
or U18962 (N_18962,N_17605,N_17620);
or U18963 (N_18963,N_17305,N_17912);
nor U18964 (N_18964,N_17530,N_17937);
or U18965 (N_18965,N_17518,N_17635);
xnor U18966 (N_18966,N_17627,N_17975);
nand U18967 (N_18967,N_17259,N_17756);
or U18968 (N_18968,N_17781,N_17459);
or U18969 (N_18969,N_17454,N_17271);
xor U18970 (N_18970,N_17091,N_17771);
or U18971 (N_18971,N_17850,N_17353);
or U18972 (N_18972,N_17246,N_17784);
or U18973 (N_18973,N_17267,N_17549);
xnor U18974 (N_18974,N_17698,N_17906);
and U18975 (N_18975,N_17042,N_17924);
nor U18976 (N_18976,N_17387,N_17349);
nand U18977 (N_18977,N_17534,N_17658);
nor U18978 (N_18978,N_17702,N_17427);
nor U18979 (N_18979,N_17252,N_17477);
nor U18980 (N_18980,N_17643,N_17874);
nand U18981 (N_18981,N_17567,N_17729);
and U18982 (N_18982,N_17093,N_17942);
or U18983 (N_18983,N_17157,N_17190);
xor U18984 (N_18984,N_17037,N_17614);
nand U18985 (N_18985,N_17356,N_17044);
nor U18986 (N_18986,N_17238,N_17702);
or U18987 (N_18987,N_17634,N_17576);
or U18988 (N_18988,N_17629,N_17855);
and U18989 (N_18989,N_17474,N_17961);
xnor U18990 (N_18990,N_17797,N_17999);
and U18991 (N_18991,N_17592,N_17030);
nand U18992 (N_18992,N_17521,N_17449);
xnor U18993 (N_18993,N_17295,N_17279);
or U18994 (N_18994,N_17263,N_17687);
nor U18995 (N_18995,N_17599,N_17043);
nor U18996 (N_18996,N_17989,N_17160);
or U18997 (N_18997,N_17506,N_17854);
nand U18998 (N_18998,N_17223,N_17248);
nand U18999 (N_18999,N_17745,N_17683);
nor U19000 (N_19000,N_18521,N_18164);
xnor U19001 (N_19001,N_18782,N_18530);
nor U19002 (N_19002,N_18195,N_18386);
or U19003 (N_19003,N_18991,N_18414);
nor U19004 (N_19004,N_18206,N_18799);
xor U19005 (N_19005,N_18999,N_18268);
or U19006 (N_19006,N_18748,N_18681);
and U19007 (N_19007,N_18775,N_18265);
or U19008 (N_19008,N_18026,N_18417);
nor U19009 (N_19009,N_18781,N_18547);
xnor U19010 (N_19010,N_18773,N_18944);
nand U19011 (N_19011,N_18533,N_18849);
and U19012 (N_19012,N_18976,N_18526);
xor U19013 (N_19013,N_18177,N_18093);
nand U19014 (N_19014,N_18495,N_18353);
xnor U19015 (N_19015,N_18829,N_18313);
and U19016 (N_19016,N_18755,N_18559);
nor U19017 (N_19017,N_18408,N_18046);
nor U19018 (N_19018,N_18585,N_18742);
nand U19019 (N_19019,N_18772,N_18867);
nor U19020 (N_19020,N_18270,N_18831);
nor U19021 (N_19021,N_18394,N_18440);
nand U19022 (N_19022,N_18760,N_18610);
and U19023 (N_19023,N_18184,N_18611);
nor U19024 (N_19024,N_18818,N_18591);
or U19025 (N_19025,N_18697,N_18438);
and U19026 (N_19026,N_18683,N_18628);
nand U19027 (N_19027,N_18938,N_18930);
and U19028 (N_19028,N_18152,N_18161);
or U19029 (N_19029,N_18001,N_18666);
or U19030 (N_19030,N_18920,N_18701);
xor U19031 (N_19031,N_18513,N_18665);
xor U19032 (N_19032,N_18817,N_18463);
and U19033 (N_19033,N_18291,N_18770);
nand U19034 (N_19034,N_18565,N_18214);
xor U19035 (N_19035,N_18955,N_18556);
or U19036 (N_19036,N_18859,N_18128);
xor U19037 (N_19037,N_18101,N_18658);
xor U19038 (N_19038,N_18235,N_18435);
xnor U19039 (N_19039,N_18471,N_18809);
or U19040 (N_19040,N_18765,N_18832);
or U19041 (N_19041,N_18323,N_18549);
and U19042 (N_19042,N_18346,N_18006);
xnor U19043 (N_19043,N_18605,N_18857);
nor U19044 (N_19044,N_18534,N_18956);
and U19045 (N_19045,N_18117,N_18641);
xor U19046 (N_19046,N_18788,N_18081);
xnor U19047 (N_19047,N_18361,N_18669);
nor U19048 (N_19048,N_18300,N_18858);
xor U19049 (N_19049,N_18227,N_18306);
nand U19050 (N_19050,N_18953,N_18318);
xnor U19051 (N_19051,N_18162,N_18183);
xnor U19052 (N_19052,N_18627,N_18529);
and U19053 (N_19053,N_18058,N_18151);
and U19054 (N_19054,N_18025,N_18899);
nand U19055 (N_19055,N_18631,N_18430);
nand U19056 (N_19056,N_18708,N_18888);
and U19057 (N_19057,N_18780,N_18543);
nor U19058 (N_19058,N_18222,N_18057);
or U19059 (N_19059,N_18497,N_18219);
or U19060 (N_19060,N_18454,N_18401);
xor U19061 (N_19061,N_18808,N_18089);
nor U19062 (N_19062,N_18267,N_18802);
nand U19063 (N_19063,N_18558,N_18800);
nand U19064 (N_19064,N_18961,N_18672);
and U19065 (N_19065,N_18277,N_18531);
nand U19066 (N_19066,N_18078,N_18874);
nor U19067 (N_19067,N_18236,N_18049);
or U19068 (N_19068,N_18727,N_18718);
and U19069 (N_19069,N_18916,N_18994);
nand U19070 (N_19070,N_18040,N_18600);
xor U19071 (N_19071,N_18871,N_18295);
or U19072 (N_19072,N_18753,N_18243);
and U19073 (N_19073,N_18848,N_18349);
xnor U19074 (N_19074,N_18992,N_18480);
or U19075 (N_19075,N_18877,N_18338);
xnor U19076 (N_19076,N_18751,N_18998);
and U19077 (N_19077,N_18493,N_18758);
nand U19078 (N_19078,N_18217,N_18569);
xor U19079 (N_19079,N_18729,N_18134);
xnor U19080 (N_19080,N_18553,N_18292);
xor U19081 (N_19081,N_18122,N_18798);
and U19082 (N_19082,N_18473,N_18429);
nand U19083 (N_19083,N_18275,N_18392);
or U19084 (N_19084,N_18891,N_18157);
nor U19085 (N_19085,N_18575,N_18482);
or U19086 (N_19086,N_18316,N_18145);
xor U19087 (N_19087,N_18964,N_18837);
nor U19088 (N_19088,N_18839,N_18873);
nor U19089 (N_19089,N_18237,N_18474);
xnor U19090 (N_19090,N_18540,N_18951);
nand U19091 (N_19091,N_18189,N_18357);
nor U19092 (N_19092,N_18741,N_18035);
nand U19093 (N_19093,N_18902,N_18036);
nor U19094 (N_19094,N_18375,N_18745);
or U19095 (N_19095,N_18198,N_18312);
nor U19096 (N_19096,N_18393,N_18550);
nor U19097 (N_19097,N_18649,N_18965);
nor U19098 (N_19098,N_18546,N_18351);
nand U19099 (N_19099,N_18031,N_18703);
or U19100 (N_19100,N_18862,N_18284);
and U19101 (N_19101,N_18000,N_18608);
or U19102 (N_19102,N_18475,N_18717);
and U19103 (N_19103,N_18344,N_18112);
nor U19104 (N_19104,N_18586,N_18050);
nand U19105 (N_19105,N_18983,N_18617);
nor U19106 (N_19106,N_18459,N_18042);
nand U19107 (N_19107,N_18372,N_18340);
nor U19108 (N_19108,N_18055,N_18861);
nand U19109 (N_19109,N_18982,N_18619);
nand U19110 (N_19110,N_18988,N_18716);
xor U19111 (N_19111,N_18460,N_18133);
xnor U19112 (N_19112,N_18850,N_18095);
xnor U19113 (N_19113,N_18045,N_18579);
xor U19114 (N_19114,N_18905,N_18041);
nor U19115 (N_19115,N_18362,N_18015);
and U19116 (N_19116,N_18067,N_18111);
or U19117 (N_19117,N_18694,N_18621);
or U19118 (N_19118,N_18505,N_18677);
and U19119 (N_19119,N_18803,N_18088);
or U19120 (N_19120,N_18166,N_18943);
and U19121 (N_19121,N_18257,N_18187);
nor U19122 (N_19122,N_18171,N_18406);
and U19123 (N_19123,N_18806,N_18130);
nand U19124 (N_19124,N_18519,N_18931);
and U19125 (N_19125,N_18739,N_18653);
or U19126 (N_19126,N_18525,N_18894);
xnor U19127 (N_19127,N_18977,N_18342);
nor U19128 (N_19128,N_18704,N_18216);
nor U19129 (N_19129,N_18733,N_18470);
nand U19130 (N_19130,N_18181,N_18626);
and U19131 (N_19131,N_18796,N_18185);
and U19132 (N_19132,N_18256,N_18172);
or U19133 (N_19133,N_18528,N_18539);
nand U19134 (N_19134,N_18768,N_18702);
or U19135 (N_19135,N_18110,N_18103);
nor U19136 (N_19136,N_18437,N_18979);
nand U19137 (N_19137,N_18978,N_18288);
nor U19138 (N_19138,N_18347,N_18826);
or U19139 (N_19139,N_18228,N_18940);
and U19140 (N_19140,N_18197,N_18464);
nor U19141 (N_19141,N_18064,N_18129);
nand U19142 (N_19142,N_18106,N_18352);
nand U19143 (N_19143,N_18461,N_18835);
and U19144 (N_19144,N_18247,N_18391);
xnor U19145 (N_19145,N_18146,N_18335);
and U19146 (N_19146,N_18434,N_18008);
and U19147 (N_19147,N_18893,N_18638);
or U19148 (N_19148,N_18934,N_18179);
nor U19149 (N_19149,N_18696,N_18834);
and U19150 (N_19150,N_18618,N_18620);
and U19151 (N_19151,N_18757,N_18512);
nand U19152 (N_19152,N_18625,N_18900);
nand U19153 (N_19153,N_18245,N_18465);
nand U19154 (N_19154,N_18327,N_18801);
and U19155 (N_19155,N_18141,N_18113);
nor U19156 (N_19156,N_18845,N_18178);
nand U19157 (N_19157,N_18333,N_18136);
or U19158 (N_19158,N_18661,N_18334);
nand U19159 (N_19159,N_18397,N_18173);
or U19160 (N_19160,N_18767,N_18950);
nand U19161 (N_19161,N_18815,N_18224);
nand U19162 (N_19162,N_18844,N_18494);
and U19163 (N_19163,N_18840,N_18079);
and U19164 (N_19164,N_18825,N_18730);
xor U19165 (N_19165,N_18853,N_18090);
nand U19166 (N_19166,N_18407,N_18623);
xnor U19167 (N_19167,N_18148,N_18663);
or U19168 (N_19168,N_18545,N_18211);
nand U19169 (N_19169,N_18980,N_18252);
nor U19170 (N_19170,N_18912,N_18032);
nand U19171 (N_19171,N_18131,N_18984);
xor U19172 (N_19172,N_18885,N_18761);
xor U19173 (N_19173,N_18005,N_18795);
or U19174 (N_19174,N_18012,N_18642);
xor U19175 (N_19175,N_18144,N_18186);
or U19176 (N_19176,N_18538,N_18897);
and U19177 (N_19177,N_18180,N_18478);
or U19178 (N_19178,N_18385,N_18643);
nor U19179 (N_19179,N_18142,N_18380);
nand U19180 (N_19180,N_18400,N_18226);
nor U19181 (N_19181,N_18154,N_18132);
xnor U19182 (N_19182,N_18294,N_18830);
nor U19183 (N_19183,N_18926,N_18710);
nand U19184 (N_19184,N_18432,N_18039);
xor U19185 (N_19185,N_18975,N_18820);
or U19186 (N_19186,N_18827,N_18678);
and U19187 (N_19187,N_18426,N_18963);
nor U19188 (N_19188,N_18439,N_18213);
and U19189 (N_19189,N_18937,N_18573);
and U19190 (N_19190,N_18254,N_18399);
nor U19191 (N_19191,N_18870,N_18193);
and U19192 (N_19192,N_18952,N_18996);
or U19193 (N_19193,N_18396,N_18149);
xor U19194 (N_19194,N_18107,N_18909);
or U19195 (N_19195,N_18700,N_18421);
or U19196 (N_19196,N_18210,N_18508);
or U19197 (N_19197,N_18080,N_18379);
xnor U19198 (N_19198,N_18604,N_18690);
xor U19199 (N_19199,N_18687,N_18315);
nand U19200 (N_19200,N_18776,N_18972);
and U19201 (N_19201,N_18726,N_18358);
or U19202 (N_19202,N_18833,N_18572);
nand U19203 (N_19203,N_18234,N_18192);
nor U19204 (N_19204,N_18632,N_18410);
and U19205 (N_19205,N_18285,N_18652);
nand U19206 (N_19206,N_18680,N_18232);
xnor U19207 (N_19207,N_18489,N_18960);
and U19208 (N_19208,N_18679,N_18566);
xnor U19209 (N_19209,N_18427,N_18024);
and U19210 (N_19210,N_18875,N_18403);
or U19211 (N_19211,N_18260,N_18962);
nand U19212 (N_19212,N_18092,N_18348);
xor U19213 (N_19213,N_18728,N_18087);
nor U19214 (N_19214,N_18374,N_18203);
nand U19215 (N_19215,N_18370,N_18967);
nand U19216 (N_19216,N_18371,N_18928);
nand U19217 (N_19217,N_18664,N_18455);
and U19218 (N_19218,N_18249,N_18423);
and U19219 (N_19219,N_18202,N_18121);
nor U19220 (N_19220,N_18878,N_18174);
or U19221 (N_19221,N_18248,N_18948);
nor U19222 (N_19222,N_18021,N_18947);
and U19223 (N_19223,N_18648,N_18303);
or U19224 (N_19224,N_18066,N_18156);
nor U19225 (N_19225,N_18766,N_18492);
nand U19226 (N_19226,N_18030,N_18231);
or U19227 (N_19227,N_18317,N_18954);
nand U19228 (N_19228,N_18935,N_18901);
nor U19229 (N_19229,N_18376,N_18259);
and U19230 (N_19230,N_18517,N_18774);
or U19231 (N_19231,N_18524,N_18242);
or U19232 (N_19232,N_18932,N_18028);
and U19233 (N_19233,N_18744,N_18220);
xor U19234 (N_19234,N_18139,N_18446);
nor U19235 (N_19235,N_18555,N_18673);
nor U19236 (N_19236,N_18711,N_18458);
nor U19237 (N_19237,N_18230,N_18903);
nand U19238 (N_19238,N_18881,N_18548);
nor U19239 (N_19239,N_18309,N_18887);
or U19240 (N_19240,N_18176,N_18662);
or U19241 (N_19241,N_18233,N_18215);
nand U19242 (N_19242,N_18207,N_18002);
xor U19243 (N_19243,N_18759,N_18108);
or U19244 (N_19244,N_18476,N_18823);
and U19245 (N_19245,N_18229,N_18511);
and U19246 (N_19246,N_18056,N_18957);
nor U19247 (N_19247,N_18890,N_18749);
and U19248 (N_19248,N_18650,N_18160);
and U19249 (N_19249,N_18424,N_18044);
or U19250 (N_19250,N_18686,N_18262);
nand U19251 (N_19251,N_18995,N_18264);
and U19252 (N_19252,N_18712,N_18034);
xor U19253 (N_19253,N_18986,N_18851);
and U19254 (N_19254,N_18514,N_18587);
xnor U19255 (N_19255,N_18194,N_18743);
xor U19256 (N_19256,N_18367,N_18822);
nand U19257 (N_19257,N_18856,N_18280);
xnor U19258 (N_19258,N_18790,N_18168);
and U19259 (N_19259,N_18593,N_18824);
nor U19260 (N_19260,N_18283,N_18736);
nor U19261 (N_19261,N_18813,N_18286);
or U19262 (N_19262,N_18289,N_18395);
and U19263 (N_19263,N_18135,N_18420);
xor U19264 (N_19264,N_18488,N_18506);
xor U19265 (N_19265,N_18125,N_18239);
nor U19266 (N_19266,N_18048,N_18910);
nand U19267 (N_19267,N_18022,N_18936);
xor U19268 (N_19268,N_18898,N_18792);
or U19269 (N_19269,N_18281,N_18656);
nand U19270 (N_19270,N_18787,N_18724);
nand U19271 (N_19271,N_18671,N_18409);
nor U19272 (N_19272,N_18051,N_18115);
and U19273 (N_19273,N_18865,N_18784);
xor U19274 (N_19274,N_18725,N_18287);
or U19275 (N_19275,N_18322,N_18273);
xor U19276 (N_19276,N_18915,N_18794);
nor U19277 (N_19277,N_18918,N_18276);
and U19278 (N_19278,N_18301,N_18968);
nand U19279 (N_19279,N_18043,N_18373);
nor U19280 (N_19280,N_18923,N_18140);
nor U19281 (N_19281,N_18904,N_18942);
xnor U19282 (N_19282,N_18246,N_18007);
or U19283 (N_19283,N_18250,N_18483);
nor U19284 (N_19284,N_18634,N_18116);
nor U19285 (N_19285,N_18053,N_18989);
nand U19286 (N_19286,N_18448,N_18381);
or U19287 (N_19287,N_18445,N_18453);
xor U19288 (N_19288,N_18630,N_18272);
and U19289 (N_19289,N_18499,N_18378);
or U19290 (N_19290,N_18212,N_18554);
nor U19291 (N_19291,N_18959,N_18114);
nor U19292 (N_19292,N_18484,N_18563);
and U19293 (N_19293,N_18033,N_18155);
xnor U19294 (N_19294,N_18769,N_18094);
nand U19295 (N_19295,N_18576,N_18271);
xor U19296 (N_19296,N_18298,N_18412);
xor U19297 (N_19297,N_18864,N_18688);
or U19298 (N_19298,N_18692,N_18188);
nor U19299 (N_19299,N_18501,N_18723);
nor U19300 (N_19300,N_18685,N_18158);
nor U19301 (N_19301,N_18970,N_18100);
or U19302 (N_19302,N_18072,N_18544);
nor U19303 (N_19303,N_18330,N_18945);
nor U19304 (N_19304,N_18191,N_18536);
nand U19305 (N_19305,N_18302,N_18869);
and U19306 (N_19306,N_18812,N_18675);
xor U19307 (N_19307,N_18324,N_18595);
xnor U19308 (N_19308,N_18906,N_18456);
nand U19309 (N_19309,N_18974,N_18908);
xor U19310 (N_19310,N_18752,N_18355);
xor U19311 (N_19311,N_18054,N_18805);
or U19312 (N_19312,N_18969,N_18472);
nand U19313 (N_19313,N_18023,N_18382);
nand U19314 (N_19314,N_18365,N_18466);
nand U19315 (N_19315,N_18615,N_18364);
xnor U19316 (N_19316,N_18383,N_18523);
or U19317 (N_19317,N_18535,N_18428);
nor U19318 (N_19318,N_18366,N_18336);
nor U19319 (N_19319,N_18077,N_18771);
xnor U19320 (N_19320,N_18542,N_18667);
nor U19321 (N_19321,N_18709,N_18527);
xnor U19322 (N_19322,N_18496,N_18075);
and U19323 (N_19323,N_18791,N_18913);
nor U19324 (N_19324,N_18098,N_18705);
or U19325 (N_19325,N_18571,N_18655);
nand U19326 (N_19326,N_18209,N_18124);
or U19327 (N_19327,N_18838,N_18126);
nand U19328 (N_19328,N_18640,N_18221);
nor U19329 (N_19329,N_18096,N_18084);
xor U19330 (N_19330,N_18811,N_18360);
or U19331 (N_19331,N_18413,N_18481);
nor U19332 (N_19332,N_18722,N_18907);
nor U19333 (N_19333,N_18895,N_18612);
or U19334 (N_19334,N_18987,N_18314);
or U19335 (N_19335,N_18764,N_18855);
and U19336 (N_19336,N_18433,N_18783);
and U19337 (N_19337,N_18919,N_18516);
nor U19338 (N_19338,N_18949,N_18841);
nand U19339 (N_19339,N_18583,N_18010);
or U19340 (N_19340,N_18356,N_18889);
and U19341 (N_19341,N_18924,N_18404);
xnor U19342 (N_19342,N_18085,N_18981);
nor U19343 (N_19343,N_18946,N_18328);
or U19344 (N_19344,N_18581,N_18606);
nand U19345 (N_19345,N_18785,N_18468);
and U19346 (N_19346,N_18485,N_18778);
nand U19347 (N_19347,N_18104,N_18200);
and U19348 (N_19348,N_18442,N_18509);
nor U19349 (N_19349,N_18359,N_18598);
or U19350 (N_19350,N_18170,N_18063);
and U19351 (N_19351,N_18646,N_18308);
xor U19352 (N_19352,N_18819,N_18502);
nor U19353 (N_19353,N_18914,N_18190);
and U19354 (N_19354,N_18027,N_18486);
nor U19355 (N_19355,N_18293,N_18105);
nor U19356 (N_19356,N_18074,N_18389);
xor U19357 (N_19357,N_18601,N_18062);
or U19358 (N_19358,N_18343,N_18756);
nand U19359 (N_19359,N_18592,N_18966);
nor U19360 (N_19360,N_18828,N_18789);
nand U19361 (N_19361,N_18065,N_18016);
or U19362 (N_19362,N_18290,N_18750);
xor U19363 (N_19363,N_18925,N_18674);
nor U19364 (N_19364,N_18415,N_18880);
nand U19365 (N_19365,N_18561,N_18447);
nor U19366 (N_19366,N_18196,N_18003);
xor U19367 (N_19367,N_18614,N_18911);
nor U19368 (N_19368,N_18603,N_18941);
nand U19369 (N_19369,N_18059,N_18052);
or U19370 (N_19370,N_18296,N_18487);
nor U19371 (N_19371,N_18274,N_18804);
nor U19372 (N_19372,N_18584,N_18354);
nor U19373 (N_19373,N_18629,N_18076);
xnor U19374 (N_19374,N_18255,N_18325);
xnor U19375 (N_19375,N_18821,N_18670);
nand U19376 (N_19376,N_18444,N_18917);
and U19377 (N_19377,N_18279,N_18807);
nand U19378 (N_19378,N_18208,N_18150);
nor U19379 (N_19379,N_18251,N_18167);
nor U19380 (N_19380,N_18163,N_18320);
nand U19381 (N_19381,N_18402,N_18238);
and U19382 (N_19382,N_18311,N_18594);
nand U19383 (N_19383,N_18071,N_18574);
nand U19384 (N_19384,N_18069,N_18326);
nand U19385 (N_19385,N_18416,N_18754);
nor U19386 (N_19386,N_18720,N_18588);
or U19387 (N_19387,N_18706,N_18261);
xnor U19388 (N_19388,N_18011,N_18589);
nor U19389 (N_19389,N_18896,N_18863);
or U19390 (N_19390,N_18120,N_18738);
nor U19391 (N_19391,N_18985,N_18387);
or U19392 (N_19392,N_18816,N_18633);
nand U19393 (N_19393,N_18580,N_18143);
or U19394 (N_19394,N_18278,N_18304);
nand U19395 (N_19395,N_18398,N_18266);
nand U19396 (N_19396,N_18047,N_18363);
xnor U19397 (N_19397,N_18282,N_18479);
or U19398 (N_19398,N_18689,N_18345);
or U19399 (N_19399,N_18939,N_18137);
nand U19400 (N_19400,N_18518,N_18390);
nor U19401 (N_19401,N_18038,N_18609);
nand U19402 (N_19402,N_18868,N_18225);
nand U19403 (N_19403,N_18639,N_18321);
nand U19404 (N_19404,N_18099,N_18847);
and U19405 (N_19405,N_18223,N_18973);
xor U19406 (N_19406,N_18568,N_18684);
or U19407 (N_19407,N_18814,N_18477);
nor U19408 (N_19408,N_18425,N_18651);
nor U19409 (N_19409,N_18882,N_18127);
and U19410 (N_19410,N_18119,N_18169);
nor U19411 (N_19411,N_18451,N_18017);
and U19412 (N_19412,N_18377,N_18929);
or U19413 (N_19413,N_18922,N_18810);
nand U19414 (N_19414,N_18138,N_18436);
xnor U19415 (N_19415,N_18083,N_18469);
nor U19416 (N_19416,N_18731,N_18746);
and U19417 (N_19417,N_18721,N_18872);
and U19418 (N_19418,N_18654,N_18199);
xor U19419 (N_19419,N_18297,N_18596);
nand U19420 (N_19420,N_18457,N_18061);
nand U19421 (N_19421,N_18734,N_18644);
nand U19422 (N_19422,N_18507,N_18740);
nand U19423 (N_19423,N_18793,N_18244);
or U19424 (N_19424,N_18892,N_18452);
and U19425 (N_19425,N_18645,N_18777);
nand U19426 (N_19426,N_18258,N_18013);
nand U19427 (N_19427,N_18153,N_18577);
nor U19428 (N_19428,N_18564,N_18510);
xnor U19429 (N_19429,N_18602,N_18560);
or U19430 (N_19430,N_18990,N_18682);
nand U19431 (N_19431,N_18599,N_18541);
xnor U19432 (N_19432,N_18443,N_18405);
or U19433 (N_19433,N_18737,N_18004);
xor U19434 (N_19434,N_18691,N_18886);
nand U19435 (N_19435,N_18073,N_18159);
nand U19436 (N_19436,N_18498,N_18567);
nand U19437 (N_19437,N_18018,N_18009);
and U19438 (N_19438,N_18332,N_18341);
or U19439 (N_19439,N_18747,N_18616);
nand U19440 (N_19440,N_18622,N_18797);
xor U19441 (N_19441,N_18866,N_18263);
and U19442 (N_19442,N_18933,N_18102);
xor U19443 (N_19443,N_18422,N_18411);
nand U19444 (N_19444,N_18713,N_18647);
and U19445 (N_19445,N_18578,N_18503);
xnor U19446 (N_19446,N_18388,N_18319);
and U19447 (N_19447,N_18462,N_18520);
and U19448 (N_19448,N_18676,N_18091);
and U19449 (N_19449,N_18491,N_18082);
nor U19450 (N_19450,N_18883,N_18431);
or U19451 (N_19451,N_18971,N_18331);
nor U19452 (N_19452,N_18876,N_18993);
or U19453 (N_19453,N_18927,N_18201);
and U19454 (N_19454,N_18597,N_18182);
or U19455 (N_19455,N_18515,N_18860);
and U19456 (N_19456,N_18842,N_18714);
xnor U19457 (N_19457,N_18607,N_18384);
xor U19458 (N_19458,N_18532,N_18350);
or U19459 (N_19459,N_18779,N_18337);
or U19460 (N_19460,N_18732,N_18707);
or U19461 (N_19461,N_18060,N_18582);
or U19462 (N_19462,N_18836,N_18118);
and U19463 (N_19463,N_18715,N_18086);
or U19464 (N_19464,N_18636,N_18241);
xor U19465 (N_19465,N_18562,N_18537);
xor U19466 (N_19466,N_18299,N_18668);
and U19467 (N_19467,N_18624,N_18014);
nand U19468 (N_19468,N_18368,N_18490);
nor U19469 (N_19469,N_18635,N_18109);
xnor U19470 (N_19470,N_18418,N_18762);
nor U19471 (N_19471,N_18659,N_18467);
nand U19472 (N_19472,N_18068,N_18253);
nand U19473 (N_19473,N_18029,N_18570);
and U19474 (N_19474,N_18419,N_18165);
or U19475 (N_19475,N_18852,N_18997);
xor U19476 (N_19476,N_18846,N_18329);
and U19477 (N_19477,N_18305,N_18339);
nand U19478 (N_19478,N_18637,N_18522);
nor U19479 (N_19479,N_18205,N_18551);
or U19480 (N_19480,N_18719,N_18450);
or U19481 (N_19481,N_18097,N_18699);
xnor U19482 (N_19482,N_18763,N_18879);
xor U19483 (N_19483,N_18657,N_18449);
xor U19484 (N_19484,N_18884,N_18369);
or U19485 (N_19485,N_18958,N_18070);
nand U19486 (N_19486,N_18786,N_18552);
xnor U19487 (N_19487,N_18204,N_18175);
or U19488 (N_19488,N_18019,N_18590);
nor U19489 (N_19489,N_18854,N_18123);
and U19490 (N_19490,N_18613,N_18441);
xnor U19491 (N_19491,N_18557,N_18307);
nand U19492 (N_19492,N_18269,N_18310);
or U19493 (N_19493,N_18504,N_18037);
nand U19494 (N_19494,N_18500,N_18020);
xnor U19495 (N_19495,N_18843,N_18147);
nor U19496 (N_19496,N_18693,N_18218);
and U19497 (N_19497,N_18240,N_18735);
and U19498 (N_19498,N_18695,N_18921);
xnor U19499 (N_19499,N_18698,N_18660);
or U19500 (N_19500,N_18391,N_18093);
nand U19501 (N_19501,N_18165,N_18535);
nor U19502 (N_19502,N_18114,N_18011);
and U19503 (N_19503,N_18252,N_18513);
nand U19504 (N_19504,N_18450,N_18866);
or U19505 (N_19505,N_18232,N_18331);
and U19506 (N_19506,N_18002,N_18973);
nor U19507 (N_19507,N_18277,N_18293);
nor U19508 (N_19508,N_18185,N_18961);
nand U19509 (N_19509,N_18436,N_18864);
and U19510 (N_19510,N_18679,N_18938);
or U19511 (N_19511,N_18570,N_18786);
xor U19512 (N_19512,N_18036,N_18444);
xnor U19513 (N_19513,N_18509,N_18368);
or U19514 (N_19514,N_18967,N_18630);
nand U19515 (N_19515,N_18607,N_18466);
nand U19516 (N_19516,N_18538,N_18631);
nand U19517 (N_19517,N_18194,N_18013);
xor U19518 (N_19518,N_18646,N_18544);
nand U19519 (N_19519,N_18258,N_18137);
nand U19520 (N_19520,N_18676,N_18499);
or U19521 (N_19521,N_18570,N_18944);
nor U19522 (N_19522,N_18488,N_18268);
nor U19523 (N_19523,N_18997,N_18095);
nand U19524 (N_19524,N_18649,N_18493);
nand U19525 (N_19525,N_18300,N_18206);
or U19526 (N_19526,N_18585,N_18527);
nand U19527 (N_19527,N_18440,N_18182);
xnor U19528 (N_19528,N_18899,N_18006);
or U19529 (N_19529,N_18924,N_18477);
nor U19530 (N_19530,N_18821,N_18044);
and U19531 (N_19531,N_18613,N_18432);
nor U19532 (N_19532,N_18321,N_18068);
xnor U19533 (N_19533,N_18657,N_18545);
and U19534 (N_19534,N_18100,N_18016);
nor U19535 (N_19535,N_18890,N_18861);
nand U19536 (N_19536,N_18844,N_18595);
and U19537 (N_19537,N_18041,N_18196);
xnor U19538 (N_19538,N_18272,N_18889);
and U19539 (N_19539,N_18690,N_18558);
or U19540 (N_19540,N_18595,N_18934);
nand U19541 (N_19541,N_18015,N_18701);
nor U19542 (N_19542,N_18463,N_18751);
xnor U19543 (N_19543,N_18433,N_18208);
xor U19544 (N_19544,N_18766,N_18557);
xnor U19545 (N_19545,N_18043,N_18325);
nor U19546 (N_19546,N_18554,N_18399);
nor U19547 (N_19547,N_18622,N_18697);
and U19548 (N_19548,N_18559,N_18265);
nand U19549 (N_19549,N_18800,N_18567);
nor U19550 (N_19550,N_18835,N_18988);
nand U19551 (N_19551,N_18357,N_18102);
xnor U19552 (N_19552,N_18468,N_18368);
xnor U19553 (N_19553,N_18314,N_18422);
or U19554 (N_19554,N_18085,N_18487);
nand U19555 (N_19555,N_18178,N_18800);
nand U19556 (N_19556,N_18182,N_18721);
and U19557 (N_19557,N_18508,N_18736);
xnor U19558 (N_19558,N_18760,N_18756);
nand U19559 (N_19559,N_18256,N_18769);
nor U19560 (N_19560,N_18512,N_18279);
nor U19561 (N_19561,N_18609,N_18238);
nand U19562 (N_19562,N_18927,N_18018);
and U19563 (N_19563,N_18951,N_18409);
xnor U19564 (N_19564,N_18811,N_18579);
xnor U19565 (N_19565,N_18784,N_18535);
or U19566 (N_19566,N_18204,N_18623);
xnor U19567 (N_19567,N_18123,N_18011);
xnor U19568 (N_19568,N_18791,N_18085);
nand U19569 (N_19569,N_18072,N_18221);
nor U19570 (N_19570,N_18820,N_18214);
or U19571 (N_19571,N_18054,N_18014);
nor U19572 (N_19572,N_18158,N_18357);
nor U19573 (N_19573,N_18298,N_18972);
or U19574 (N_19574,N_18839,N_18048);
nand U19575 (N_19575,N_18663,N_18485);
nand U19576 (N_19576,N_18063,N_18204);
xnor U19577 (N_19577,N_18819,N_18823);
nor U19578 (N_19578,N_18289,N_18103);
nand U19579 (N_19579,N_18207,N_18117);
and U19580 (N_19580,N_18537,N_18549);
or U19581 (N_19581,N_18657,N_18525);
and U19582 (N_19582,N_18851,N_18974);
nand U19583 (N_19583,N_18569,N_18643);
xnor U19584 (N_19584,N_18052,N_18131);
xnor U19585 (N_19585,N_18785,N_18305);
or U19586 (N_19586,N_18298,N_18114);
or U19587 (N_19587,N_18541,N_18555);
nor U19588 (N_19588,N_18196,N_18452);
or U19589 (N_19589,N_18302,N_18885);
or U19590 (N_19590,N_18864,N_18952);
or U19591 (N_19591,N_18138,N_18646);
xor U19592 (N_19592,N_18324,N_18597);
xnor U19593 (N_19593,N_18867,N_18161);
nor U19594 (N_19594,N_18066,N_18589);
nor U19595 (N_19595,N_18007,N_18611);
or U19596 (N_19596,N_18169,N_18922);
nor U19597 (N_19597,N_18302,N_18520);
nand U19598 (N_19598,N_18023,N_18936);
nor U19599 (N_19599,N_18214,N_18578);
xor U19600 (N_19600,N_18994,N_18669);
or U19601 (N_19601,N_18837,N_18303);
nand U19602 (N_19602,N_18865,N_18958);
nor U19603 (N_19603,N_18416,N_18649);
or U19604 (N_19604,N_18028,N_18260);
nand U19605 (N_19605,N_18934,N_18111);
or U19606 (N_19606,N_18040,N_18048);
and U19607 (N_19607,N_18117,N_18790);
nand U19608 (N_19608,N_18839,N_18029);
nor U19609 (N_19609,N_18750,N_18858);
nor U19610 (N_19610,N_18217,N_18937);
xnor U19611 (N_19611,N_18421,N_18092);
nor U19612 (N_19612,N_18745,N_18651);
and U19613 (N_19613,N_18555,N_18094);
xor U19614 (N_19614,N_18999,N_18148);
nand U19615 (N_19615,N_18955,N_18662);
xnor U19616 (N_19616,N_18727,N_18118);
xor U19617 (N_19617,N_18451,N_18166);
and U19618 (N_19618,N_18476,N_18835);
xnor U19619 (N_19619,N_18679,N_18386);
nor U19620 (N_19620,N_18499,N_18769);
or U19621 (N_19621,N_18806,N_18473);
nand U19622 (N_19622,N_18932,N_18234);
nor U19623 (N_19623,N_18527,N_18813);
and U19624 (N_19624,N_18580,N_18188);
xnor U19625 (N_19625,N_18204,N_18874);
or U19626 (N_19626,N_18513,N_18265);
xor U19627 (N_19627,N_18549,N_18621);
nand U19628 (N_19628,N_18410,N_18826);
and U19629 (N_19629,N_18293,N_18977);
nand U19630 (N_19630,N_18553,N_18075);
or U19631 (N_19631,N_18007,N_18070);
or U19632 (N_19632,N_18143,N_18514);
nor U19633 (N_19633,N_18122,N_18406);
nor U19634 (N_19634,N_18886,N_18962);
xor U19635 (N_19635,N_18521,N_18487);
or U19636 (N_19636,N_18727,N_18590);
and U19637 (N_19637,N_18550,N_18294);
or U19638 (N_19638,N_18666,N_18818);
and U19639 (N_19639,N_18079,N_18054);
nand U19640 (N_19640,N_18991,N_18889);
or U19641 (N_19641,N_18949,N_18513);
or U19642 (N_19642,N_18893,N_18461);
or U19643 (N_19643,N_18367,N_18240);
and U19644 (N_19644,N_18128,N_18335);
nor U19645 (N_19645,N_18487,N_18436);
xor U19646 (N_19646,N_18580,N_18899);
and U19647 (N_19647,N_18858,N_18214);
nand U19648 (N_19648,N_18854,N_18785);
and U19649 (N_19649,N_18399,N_18073);
xnor U19650 (N_19650,N_18236,N_18007);
nor U19651 (N_19651,N_18155,N_18976);
or U19652 (N_19652,N_18234,N_18204);
nand U19653 (N_19653,N_18315,N_18575);
xor U19654 (N_19654,N_18689,N_18392);
or U19655 (N_19655,N_18816,N_18246);
or U19656 (N_19656,N_18868,N_18700);
or U19657 (N_19657,N_18955,N_18563);
or U19658 (N_19658,N_18767,N_18884);
nand U19659 (N_19659,N_18806,N_18167);
and U19660 (N_19660,N_18093,N_18094);
and U19661 (N_19661,N_18131,N_18282);
nor U19662 (N_19662,N_18281,N_18610);
xor U19663 (N_19663,N_18512,N_18477);
nor U19664 (N_19664,N_18884,N_18082);
nand U19665 (N_19665,N_18528,N_18731);
nor U19666 (N_19666,N_18101,N_18035);
or U19667 (N_19667,N_18808,N_18257);
or U19668 (N_19668,N_18450,N_18518);
nand U19669 (N_19669,N_18409,N_18089);
nand U19670 (N_19670,N_18256,N_18559);
and U19671 (N_19671,N_18157,N_18093);
or U19672 (N_19672,N_18928,N_18452);
or U19673 (N_19673,N_18192,N_18386);
nand U19674 (N_19674,N_18708,N_18761);
xnor U19675 (N_19675,N_18501,N_18994);
nor U19676 (N_19676,N_18972,N_18166);
or U19677 (N_19677,N_18809,N_18950);
or U19678 (N_19678,N_18078,N_18912);
or U19679 (N_19679,N_18982,N_18091);
and U19680 (N_19680,N_18280,N_18542);
or U19681 (N_19681,N_18027,N_18256);
nand U19682 (N_19682,N_18079,N_18092);
nand U19683 (N_19683,N_18870,N_18832);
xnor U19684 (N_19684,N_18145,N_18564);
xnor U19685 (N_19685,N_18386,N_18572);
xnor U19686 (N_19686,N_18706,N_18100);
nand U19687 (N_19687,N_18630,N_18425);
and U19688 (N_19688,N_18474,N_18325);
and U19689 (N_19689,N_18626,N_18044);
and U19690 (N_19690,N_18122,N_18071);
nand U19691 (N_19691,N_18405,N_18537);
nor U19692 (N_19692,N_18479,N_18108);
nand U19693 (N_19693,N_18496,N_18130);
nor U19694 (N_19694,N_18368,N_18276);
nand U19695 (N_19695,N_18166,N_18544);
xnor U19696 (N_19696,N_18076,N_18025);
xor U19697 (N_19697,N_18788,N_18348);
nor U19698 (N_19698,N_18456,N_18736);
xnor U19699 (N_19699,N_18202,N_18742);
or U19700 (N_19700,N_18379,N_18507);
xnor U19701 (N_19701,N_18962,N_18147);
xnor U19702 (N_19702,N_18577,N_18092);
and U19703 (N_19703,N_18758,N_18121);
and U19704 (N_19704,N_18366,N_18437);
and U19705 (N_19705,N_18272,N_18491);
nor U19706 (N_19706,N_18724,N_18798);
xnor U19707 (N_19707,N_18247,N_18314);
nor U19708 (N_19708,N_18960,N_18997);
nor U19709 (N_19709,N_18272,N_18006);
or U19710 (N_19710,N_18257,N_18966);
xnor U19711 (N_19711,N_18432,N_18103);
or U19712 (N_19712,N_18197,N_18547);
and U19713 (N_19713,N_18628,N_18793);
xor U19714 (N_19714,N_18633,N_18496);
or U19715 (N_19715,N_18666,N_18362);
xnor U19716 (N_19716,N_18041,N_18342);
or U19717 (N_19717,N_18262,N_18372);
nand U19718 (N_19718,N_18416,N_18404);
nand U19719 (N_19719,N_18391,N_18003);
or U19720 (N_19720,N_18144,N_18845);
nand U19721 (N_19721,N_18276,N_18347);
xnor U19722 (N_19722,N_18441,N_18416);
nor U19723 (N_19723,N_18545,N_18194);
and U19724 (N_19724,N_18628,N_18737);
and U19725 (N_19725,N_18455,N_18334);
and U19726 (N_19726,N_18323,N_18182);
or U19727 (N_19727,N_18377,N_18951);
or U19728 (N_19728,N_18465,N_18638);
nand U19729 (N_19729,N_18180,N_18533);
xnor U19730 (N_19730,N_18160,N_18163);
and U19731 (N_19731,N_18305,N_18935);
xnor U19732 (N_19732,N_18056,N_18010);
and U19733 (N_19733,N_18276,N_18184);
or U19734 (N_19734,N_18430,N_18898);
and U19735 (N_19735,N_18358,N_18950);
nand U19736 (N_19736,N_18602,N_18442);
or U19737 (N_19737,N_18162,N_18909);
or U19738 (N_19738,N_18795,N_18651);
nand U19739 (N_19739,N_18212,N_18408);
xnor U19740 (N_19740,N_18244,N_18375);
or U19741 (N_19741,N_18461,N_18542);
xor U19742 (N_19742,N_18338,N_18453);
xor U19743 (N_19743,N_18145,N_18017);
or U19744 (N_19744,N_18393,N_18676);
xnor U19745 (N_19745,N_18794,N_18708);
nor U19746 (N_19746,N_18925,N_18508);
nand U19747 (N_19747,N_18528,N_18616);
and U19748 (N_19748,N_18595,N_18365);
or U19749 (N_19749,N_18210,N_18063);
nand U19750 (N_19750,N_18649,N_18936);
and U19751 (N_19751,N_18422,N_18924);
or U19752 (N_19752,N_18192,N_18723);
or U19753 (N_19753,N_18818,N_18302);
nand U19754 (N_19754,N_18421,N_18624);
nand U19755 (N_19755,N_18502,N_18271);
or U19756 (N_19756,N_18732,N_18181);
and U19757 (N_19757,N_18125,N_18343);
or U19758 (N_19758,N_18286,N_18635);
or U19759 (N_19759,N_18623,N_18768);
nand U19760 (N_19760,N_18284,N_18603);
xor U19761 (N_19761,N_18997,N_18034);
xor U19762 (N_19762,N_18055,N_18493);
xor U19763 (N_19763,N_18455,N_18679);
or U19764 (N_19764,N_18757,N_18499);
xor U19765 (N_19765,N_18447,N_18107);
xnor U19766 (N_19766,N_18872,N_18464);
nor U19767 (N_19767,N_18682,N_18564);
nand U19768 (N_19768,N_18146,N_18159);
nor U19769 (N_19769,N_18634,N_18915);
nor U19770 (N_19770,N_18683,N_18318);
nand U19771 (N_19771,N_18040,N_18191);
or U19772 (N_19772,N_18874,N_18794);
or U19773 (N_19773,N_18986,N_18271);
nor U19774 (N_19774,N_18782,N_18337);
xnor U19775 (N_19775,N_18920,N_18338);
nand U19776 (N_19776,N_18912,N_18110);
or U19777 (N_19777,N_18148,N_18442);
or U19778 (N_19778,N_18132,N_18979);
nor U19779 (N_19779,N_18397,N_18399);
or U19780 (N_19780,N_18106,N_18525);
nor U19781 (N_19781,N_18105,N_18979);
xor U19782 (N_19782,N_18043,N_18552);
or U19783 (N_19783,N_18588,N_18504);
nand U19784 (N_19784,N_18687,N_18955);
nor U19785 (N_19785,N_18433,N_18960);
nand U19786 (N_19786,N_18028,N_18591);
xor U19787 (N_19787,N_18270,N_18676);
nor U19788 (N_19788,N_18604,N_18945);
xor U19789 (N_19789,N_18977,N_18444);
xor U19790 (N_19790,N_18980,N_18937);
nor U19791 (N_19791,N_18409,N_18999);
nor U19792 (N_19792,N_18236,N_18311);
and U19793 (N_19793,N_18342,N_18401);
and U19794 (N_19794,N_18414,N_18394);
or U19795 (N_19795,N_18648,N_18618);
and U19796 (N_19796,N_18148,N_18323);
or U19797 (N_19797,N_18095,N_18725);
nand U19798 (N_19798,N_18458,N_18049);
xor U19799 (N_19799,N_18121,N_18131);
xnor U19800 (N_19800,N_18117,N_18414);
and U19801 (N_19801,N_18771,N_18141);
nand U19802 (N_19802,N_18521,N_18246);
nand U19803 (N_19803,N_18649,N_18295);
nor U19804 (N_19804,N_18889,N_18345);
and U19805 (N_19805,N_18448,N_18795);
and U19806 (N_19806,N_18484,N_18577);
and U19807 (N_19807,N_18277,N_18539);
and U19808 (N_19808,N_18029,N_18203);
and U19809 (N_19809,N_18868,N_18572);
nor U19810 (N_19810,N_18677,N_18027);
and U19811 (N_19811,N_18088,N_18620);
xor U19812 (N_19812,N_18832,N_18332);
or U19813 (N_19813,N_18130,N_18109);
or U19814 (N_19814,N_18218,N_18726);
xor U19815 (N_19815,N_18103,N_18097);
or U19816 (N_19816,N_18020,N_18818);
xnor U19817 (N_19817,N_18781,N_18383);
nor U19818 (N_19818,N_18364,N_18468);
or U19819 (N_19819,N_18346,N_18557);
and U19820 (N_19820,N_18366,N_18838);
and U19821 (N_19821,N_18271,N_18694);
nor U19822 (N_19822,N_18714,N_18117);
nor U19823 (N_19823,N_18962,N_18972);
nand U19824 (N_19824,N_18739,N_18084);
nand U19825 (N_19825,N_18615,N_18196);
xor U19826 (N_19826,N_18022,N_18104);
and U19827 (N_19827,N_18843,N_18432);
nor U19828 (N_19828,N_18450,N_18629);
xnor U19829 (N_19829,N_18352,N_18192);
nor U19830 (N_19830,N_18029,N_18036);
nor U19831 (N_19831,N_18915,N_18507);
nand U19832 (N_19832,N_18527,N_18662);
nor U19833 (N_19833,N_18972,N_18898);
nand U19834 (N_19834,N_18274,N_18601);
and U19835 (N_19835,N_18447,N_18175);
and U19836 (N_19836,N_18894,N_18527);
nand U19837 (N_19837,N_18794,N_18643);
nand U19838 (N_19838,N_18651,N_18399);
xnor U19839 (N_19839,N_18350,N_18858);
xor U19840 (N_19840,N_18218,N_18521);
xnor U19841 (N_19841,N_18002,N_18623);
xor U19842 (N_19842,N_18392,N_18591);
and U19843 (N_19843,N_18791,N_18690);
or U19844 (N_19844,N_18627,N_18428);
xnor U19845 (N_19845,N_18323,N_18125);
nor U19846 (N_19846,N_18157,N_18736);
xor U19847 (N_19847,N_18997,N_18672);
or U19848 (N_19848,N_18594,N_18836);
or U19849 (N_19849,N_18671,N_18338);
nor U19850 (N_19850,N_18055,N_18620);
xnor U19851 (N_19851,N_18349,N_18053);
nand U19852 (N_19852,N_18270,N_18914);
or U19853 (N_19853,N_18574,N_18814);
nor U19854 (N_19854,N_18377,N_18823);
nand U19855 (N_19855,N_18445,N_18452);
or U19856 (N_19856,N_18977,N_18612);
nor U19857 (N_19857,N_18113,N_18743);
nor U19858 (N_19858,N_18229,N_18546);
xor U19859 (N_19859,N_18970,N_18494);
nor U19860 (N_19860,N_18242,N_18236);
and U19861 (N_19861,N_18862,N_18003);
or U19862 (N_19862,N_18721,N_18854);
xnor U19863 (N_19863,N_18999,N_18871);
or U19864 (N_19864,N_18480,N_18321);
xor U19865 (N_19865,N_18592,N_18396);
or U19866 (N_19866,N_18176,N_18040);
xor U19867 (N_19867,N_18582,N_18967);
nor U19868 (N_19868,N_18906,N_18260);
and U19869 (N_19869,N_18087,N_18209);
and U19870 (N_19870,N_18720,N_18549);
and U19871 (N_19871,N_18388,N_18672);
xnor U19872 (N_19872,N_18659,N_18317);
nor U19873 (N_19873,N_18504,N_18602);
xnor U19874 (N_19874,N_18627,N_18009);
or U19875 (N_19875,N_18296,N_18481);
xnor U19876 (N_19876,N_18919,N_18179);
nand U19877 (N_19877,N_18508,N_18884);
nor U19878 (N_19878,N_18844,N_18427);
or U19879 (N_19879,N_18221,N_18048);
nand U19880 (N_19880,N_18268,N_18876);
nand U19881 (N_19881,N_18416,N_18503);
or U19882 (N_19882,N_18669,N_18744);
nor U19883 (N_19883,N_18541,N_18894);
nand U19884 (N_19884,N_18844,N_18305);
xnor U19885 (N_19885,N_18541,N_18994);
xnor U19886 (N_19886,N_18110,N_18288);
and U19887 (N_19887,N_18839,N_18127);
nor U19888 (N_19888,N_18843,N_18823);
nor U19889 (N_19889,N_18644,N_18731);
and U19890 (N_19890,N_18262,N_18227);
and U19891 (N_19891,N_18255,N_18858);
or U19892 (N_19892,N_18398,N_18340);
or U19893 (N_19893,N_18784,N_18156);
xor U19894 (N_19894,N_18824,N_18966);
nor U19895 (N_19895,N_18952,N_18594);
xnor U19896 (N_19896,N_18155,N_18553);
nor U19897 (N_19897,N_18275,N_18872);
nor U19898 (N_19898,N_18666,N_18592);
and U19899 (N_19899,N_18367,N_18691);
and U19900 (N_19900,N_18606,N_18938);
nor U19901 (N_19901,N_18729,N_18925);
or U19902 (N_19902,N_18337,N_18507);
and U19903 (N_19903,N_18657,N_18024);
xnor U19904 (N_19904,N_18477,N_18037);
nand U19905 (N_19905,N_18158,N_18555);
xor U19906 (N_19906,N_18697,N_18037);
and U19907 (N_19907,N_18045,N_18680);
and U19908 (N_19908,N_18135,N_18924);
nand U19909 (N_19909,N_18511,N_18930);
nor U19910 (N_19910,N_18786,N_18906);
nor U19911 (N_19911,N_18198,N_18979);
nor U19912 (N_19912,N_18180,N_18590);
xnor U19913 (N_19913,N_18950,N_18670);
nand U19914 (N_19914,N_18407,N_18311);
xor U19915 (N_19915,N_18280,N_18001);
nor U19916 (N_19916,N_18828,N_18946);
xor U19917 (N_19917,N_18611,N_18265);
xnor U19918 (N_19918,N_18085,N_18956);
nor U19919 (N_19919,N_18419,N_18186);
xnor U19920 (N_19920,N_18227,N_18378);
nor U19921 (N_19921,N_18947,N_18994);
xnor U19922 (N_19922,N_18289,N_18765);
xnor U19923 (N_19923,N_18469,N_18660);
and U19924 (N_19924,N_18020,N_18094);
and U19925 (N_19925,N_18843,N_18287);
nand U19926 (N_19926,N_18528,N_18764);
xor U19927 (N_19927,N_18325,N_18484);
and U19928 (N_19928,N_18921,N_18575);
nor U19929 (N_19929,N_18349,N_18304);
nor U19930 (N_19930,N_18185,N_18306);
xor U19931 (N_19931,N_18492,N_18505);
and U19932 (N_19932,N_18436,N_18687);
and U19933 (N_19933,N_18990,N_18335);
and U19934 (N_19934,N_18979,N_18815);
xnor U19935 (N_19935,N_18900,N_18436);
nor U19936 (N_19936,N_18102,N_18004);
nor U19937 (N_19937,N_18498,N_18600);
nand U19938 (N_19938,N_18718,N_18522);
and U19939 (N_19939,N_18443,N_18026);
or U19940 (N_19940,N_18387,N_18249);
nor U19941 (N_19941,N_18007,N_18091);
nand U19942 (N_19942,N_18416,N_18913);
and U19943 (N_19943,N_18526,N_18269);
nand U19944 (N_19944,N_18558,N_18130);
or U19945 (N_19945,N_18621,N_18118);
or U19946 (N_19946,N_18375,N_18514);
xor U19947 (N_19947,N_18819,N_18714);
and U19948 (N_19948,N_18308,N_18899);
nand U19949 (N_19949,N_18466,N_18911);
nor U19950 (N_19950,N_18734,N_18190);
xor U19951 (N_19951,N_18338,N_18711);
xor U19952 (N_19952,N_18768,N_18290);
or U19953 (N_19953,N_18949,N_18404);
nor U19954 (N_19954,N_18259,N_18336);
nor U19955 (N_19955,N_18430,N_18091);
nor U19956 (N_19956,N_18596,N_18240);
xor U19957 (N_19957,N_18140,N_18101);
nand U19958 (N_19958,N_18782,N_18409);
nor U19959 (N_19959,N_18206,N_18966);
and U19960 (N_19960,N_18004,N_18439);
and U19961 (N_19961,N_18028,N_18423);
or U19962 (N_19962,N_18167,N_18000);
and U19963 (N_19963,N_18628,N_18935);
xor U19964 (N_19964,N_18874,N_18093);
and U19965 (N_19965,N_18796,N_18103);
xor U19966 (N_19966,N_18390,N_18524);
and U19967 (N_19967,N_18894,N_18778);
or U19968 (N_19968,N_18207,N_18219);
or U19969 (N_19969,N_18570,N_18139);
and U19970 (N_19970,N_18992,N_18153);
nand U19971 (N_19971,N_18809,N_18257);
or U19972 (N_19972,N_18012,N_18198);
xnor U19973 (N_19973,N_18827,N_18519);
xor U19974 (N_19974,N_18405,N_18944);
and U19975 (N_19975,N_18631,N_18875);
nand U19976 (N_19976,N_18047,N_18910);
xnor U19977 (N_19977,N_18562,N_18718);
nand U19978 (N_19978,N_18891,N_18503);
nand U19979 (N_19979,N_18845,N_18490);
nor U19980 (N_19980,N_18679,N_18570);
xnor U19981 (N_19981,N_18720,N_18616);
xor U19982 (N_19982,N_18606,N_18838);
nor U19983 (N_19983,N_18527,N_18938);
and U19984 (N_19984,N_18543,N_18372);
or U19985 (N_19985,N_18468,N_18049);
nand U19986 (N_19986,N_18141,N_18630);
nor U19987 (N_19987,N_18164,N_18446);
nand U19988 (N_19988,N_18092,N_18579);
nor U19989 (N_19989,N_18030,N_18062);
nand U19990 (N_19990,N_18519,N_18026);
xnor U19991 (N_19991,N_18097,N_18193);
or U19992 (N_19992,N_18223,N_18581);
xnor U19993 (N_19993,N_18942,N_18237);
nor U19994 (N_19994,N_18425,N_18077);
nor U19995 (N_19995,N_18847,N_18897);
xnor U19996 (N_19996,N_18743,N_18888);
nand U19997 (N_19997,N_18132,N_18085);
nand U19998 (N_19998,N_18494,N_18827);
and U19999 (N_19999,N_18216,N_18166);
nand UO_0 (O_0,N_19273,N_19852);
and UO_1 (O_1,N_19744,N_19821);
or UO_2 (O_2,N_19669,N_19574);
xor UO_3 (O_3,N_19392,N_19867);
or UO_4 (O_4,N_19056,N_19366);
and UO_5 (O_5,N_19992,N_19742);
or UO_6 (O_6,N_19594,N_19402);
nor UO_7 (O_7,N_19009,N_19229);
nand UO_8 (O_8,N_19072,N_19370);
or UO_9 (O_9,N_19558,N_19639);
and UO_10 (O_10,N_19678,N_19160);
and UO_11 (O_11,N_19423,N_19339);
nand UO_12 (O_12,N_19422,N_19874);
or UO_13 (O_13,N_19491,N_19705);
or UO_14 (O_14,N_19687,N_19391);
and UO_15 (O_15,N_19762,N_19085);
xnor UO_16 (O_16,N_19469,N_19136);
xor UO_17 (O_17,N_19913,N_19731);
or UO_18 (O_18,N_19832,N_19692);
xor UO_19 (O_19,N_19472,N_19825);
or UO_20 (O_20,N_19512,N_19355);
nor UO_21 (O_21,N_19965,N_19327);
nor UO_22 (O_22,N_19066,N_19257);
nand UO_23 (O_23,N_19433,N_19971);
xnor UO_24 (O_24,N_19771,N_19441);
nor UO_25 (O_25,N_19973,N_19814);
xnor UO_26 (O_26,N_19408,N_19443);
nor UO_27 (O_27,N_19298,N_19984);
nor UO_28 (O_28,N_19276,N_19727);
nand UO_29 (O_29,N_19959,N_19995);
or UO_30 (O_30,N_19537,N_19330);
and UO_31 (O_31,N_19754,N_19407);
nor UO_32 (O_32,N_19732,N_19958);
and UO_33 (O_33,N_19487,N_19395);
nor UO_34 (O_34,N_19680,N_19657);
or UO_35 (O_35,N_19474,N_19204);
or UO_36 (O_36,N_19962,N_19007);
nand UO_37 (O_37,N_19131,N_19698);
xnor UO_38 (O_38,N_19910,N_19592);
nand UO_39 (O_39,N_19767,N_19784);
or UO_40 (O_40,N_19760,N_19865);
and UO_41 (O_41,N_19079,N_19262);
nor UO_42 (O_42,N_19340,N_19166);
nand UO_43 (O_43,N_19719,N_19180);
nor UO_44 (O_44,N_19288,N_19244);
xor UO_45 (O_45,N_19075,N_19186);
and UO_46 (O_46,N_19764,N_19159);
nand UO_47 (O_47,N_19134,N_19815);
nand UO_48 (O_48,N_19893,N_19505);
and UO_49 (O_49,N_19745,N_19854);
xnor UO_50 (O_50,N_19647,N_19923);
xnor UO_51 (O_51,N_19855,N_19289);
nand UO_52 (O_52,N_19444,N_19036);
nand UO_53 (O_53,N_19686,N_19055);
nor UO_54 (O_54,N_19064,N_19779);
and UO_55 (O_55,N_19634,N_19305);
xor UO_56 (O_56,N_19429,N_19254);
nor UO_57 (O_57,N_19994,N_19871);
nor UO_58 (O_58,N_19718,N_19615);
xor UO_59 (O_59,N_19747,N_19570);
or UO_60 (O_60,N_19794,N_19556);
xnor UO_61 (O_61,N_19112,N_19979);
nor UO_62 (O_62,N_19479,N_19403);
xnor UO_63 (O_63,N_19697,N_19337);
xor UO_64 (O_64,N_19541,N_19387);
nand UO_65 (O_65,N_19290,N_19781);
xnor UO_66 (O_66,N_19125,N_19384);
nand UO_67 (O_67,N_19675,N_19077);
or UO_68 (O_68,N_19383,N_19349);
nand UO_69 (O_69,N_19437,N_19324);
xor UO_70 (O_70,N_19957,N_19926);
and UO_71 (O_71,N_19086,N_19532);
nand UO_72 (O_72,N_19242,N_19191);
nand UO_73 (O_73,N_19184,N_19380);
nor UO_74 (O_74,N_19507,N_19665);
or UO_75 (O_75,N_19533,N_19695);
nand UO_76 (O_76,N_19252,N_19357);
and UO_77 (O_77,N_19772,N_19827);
nand UO_78 (O_78,N_19361,N_19153);
nor UO_79 (O_79,N_19224,N_19037);
and UO_80 (O_80,N_19757,N_19202);
and UO_81 (O_81,N_19530,N_19683);
nor UO_82 (O_82,N_19911,N_19809);
and UO_83 (O_83,N_19409,N_19644);
or UO_84 (O_84,N_19411,N_19081);
xor UO_85 (O_85,N_19619,N_19377);
nand UO_86 (O_86,N_19005,N_19097);
xnor UO_87 (O_87,N_19713,N_19988);
and UO_88 (O_88,N_19144,N_19044);
nor UO_89 (O_89,N_19999,N_19516);
or UO_90 (O_90,N_19301,N_19483);
nand UO_91 (O_91,N_19451,N_19351);
and UO_92 (O_92,N_19199,N_19869);
xnor UO_93 (O_93,N_19755,N_19328);
and UO_94 (O_94,N_19930,N_19632);
nor UO_95 (O_95,N_19167,N_19808);
xnor UO_96 (O_96,N_19246,N_19297);
nor UO_97 (O_97,N_19266,N_19836);
nor UO_98 (O_98,N_19130,N_19780);
nor UO_99 (O_99,N_19816,N_19714);
and UO_100 (O_100,N_19459,N_19864);
or UO_101 (O_101,N_19287,N_19927);
nor UO_102 (O_102,N_19972,N_19169);
and UO_103 (O_103,N_19255,N_19398);
and UO_104 (O_104,N_19104,N_19114);
nor UO_105 (O_105,N_19019,N_19741);
nor UO_106 (O_106,N_19148,N_19905);
and UO_107 (O_107,N_19465,N_19672);
or UO_108 (O_108,N_19799,N_19138);
or UO_109 (O_109,N_19903,N_19782);
xnor UO_110 (O_110,N_19553,N_19660);
or UO_111 (O_111,N_19579,N_19376);
nand UO_112 (O_112,N_19597,N_19162);
nand UO_113 (O_113,N_19623,N_19209);
and UO_114 (O_114,N_19861,N_19121);
xnor UO_115 (O_115,N_19758,N_19993);
nand UO_116 (O_116,N_19006,N_19664);
and UO_117 (O_117,N_19928,N_19371);
xnor UO_118 (O_118,N_19944,N_19618);
nor UO_119 (O_119,N_19043,N_19385);
or UO_120 (O_120,N_19790,N_19899);
nand UO_121 (O_121,N_19318,N_19083);
or UO_122 (O_122,N_19050,N_19550);
nand UO_123 (O_123,N_19178,N_19179);
and UO_124 (O_124,N_19481,N_19207);
or UO_125 (O_125,N_19116,N_19460);
nor UO_126 (O_126,N_19902,N_19651);
xor UO_127 (O_127,N_19195,N_19974);
xor UO_128 (O_128,N_19292,N_19878);
nand UO_129 (O_129,N_19040,N_19524);
and UO_130 (O_130,N_19613,N_19908);
or UO_131 (O_131,N_19452,N_19545);
xnor UO_132 (O_132,N_19251,N_19822);
nand UO_133 (O_133,N_19534,N_19461);
xor UO_134 (O_134,N_19563,N_19175);
and UO_135 (O_135,N_19835,N_19201);
xor UO_136 (O_136,N_19271,N_19838);
and UO_137 (O_137,N_19844,N_19120);
or UO_138 (O_138,N_19765,N_19074);
xor UO_139 (O_139,N_19113,N_19051);
nor UO_140 (O_140,N_19653,N_19087);
or UO_141 (O_141,N_19614,N_19866);
and UO_142 (O_142,N_19791,N_19593);
nand UO_143 (O_143,N_19666,N_19062);
and UO_144 (O_144,N_19933,N_19981);
nor UO_145 (O_145,N_19197,N_19830);
nor UO_146 (O_146,N_19875,N_19900);
or UO_147 (O_147,N_19863,N_19624);
nor UO_148 (O_148,N_19343,N_19227);
nand UO_149 (O_149,N_19949,N_19659);
and UO_150 (O_150,N_19796,N_19859);
and UO_151 (O_151,N_19599,N_19560);
nor UO_152 (O_152,N_19544,N_19369);
nand UO_153 (O_153,N_19696,N_19945);
nand UO_154 (O_154,N_19372,N_19468);
nand UO_155 (O_155,N_19308,N_19420);
xor UO_156 (O_156,N_19098,N_19803);
xnor UO_157 (O_157,N_19275,N_19840);
and UO_158 (O_158,N_19270,N_19707);
nor UO_159 (O_159,N_19219,N_19956);
nor UO_160 (O_160,N_19071,N_19506);
nor UO_161 (O_161,N_19884,N_19342);
nand UO_162 (O_162,N_19806,N_19497);
xor UO_163 (O_163,N_19249,N_19011);
nor UO_164 (O_164,N_19636,N_19906);
or UO_165 (O_165,N_19662,N_19724);
xnor UO_166 (O_166,N_19117,N_19737);
xnor UO_167 (O_167,N_19777,N_19982);
and UO_168 (O_168,N_19548,N_19968);
nor UO_169 (O_169,N_19735,N_19538);
or UO_170 (O_170,N_19084,N_19552);
or UO_171 (O_171,N_19950,N_19922);
nand UO_172 (O_172,N_19496,N_19853);
nand UO_173 (O_173,N_19730,N_19492);
xor UO_174 (O_174,N_19291,N_19650);
and UO_175 (O_175,N_19953,N_19453);
nor UO_176 (O_176,N_19736,N_19596);
or UO_177 (O_177,N_19888,N_19183);
nand UO_178 (O_178,N_19536,N_19786);
nand UO_179 (O_179,N_19137,N_19334);
and UO_180 (O_180,N_19058,N_19756);
and UO_181 (O_181,N_19316,N_19447);
nand UO_182 (O_182,N_19582,N_19753);
xnor UO_183 (O_183,N_19454,N_19263);
xor UO_184 (O_184,N_19157,N_19699);
xnor UO_185 (O_185,N_19435,N_19709);
nor UO_186 (O_186,N_19752,N_19093);
and UO_187 (O_187,N_19450,N_19419);
nand UO_188 (O_188,N_19256,N_19823);
xnor UO_189 (O_189,N_19400,N_19522);
xor UO_190 (O_190,N_19528,N_19679);
xor UO_191 (O_191,N_19245,N_19099);
xnor UO_192 (O_192,N_19529,N_19549);
and UO_193 (O_193,N_19174,N_19480);
and UO_194 (O_194,N_19417,N_19627);
xor UO_195 (O_195,N_19152,N_19939);
xor UO_196 (O_196,N_19439,N_19012);
nor UO_197 (O_197,N_19033,N_19525);
and UO_198 (O_198,N_19129,N_19498);
nor UO_199 (O_199,N_19527,N_19605);
nand UO_200 (O_200,N_19029,N_19161);
and UO_201 (O_201,N_19094,N_19111);
nand UO_202 (O_202,N_19321,N_19502);
xor UO_203 (O_203,N_19942,N_19243);
nor UO_204 (O_204,N_19685,N_19426);
xnor UO_205 (O_205,N_19022,N_19941);
and UO_206 (O_206,N_19586,N_19035);
nand UO_207 (O_207,N_19891,N_19213);
and UO_208 (O_208,N_19135,N_19917);
or UO_209 (O_209,N_19237,N_19018);
nand UO_210 (O_210,N_19590,N_19860);
nand UO_211 (O_211,N_19168,N_19580);
nor UO_212 (O_212,N_19551,N_19555);
nor UO_213 (O_213,N_19132,N_19115);
xnor UO_214 (O_214,N_19931,N_19151);
and UO_215 (O_215,N_19936,N_19015);
nor UO_216 (O_216,N_19438,N_19314);
and UO_217 (O_217,N_19065,N_19028);
nor UO_218 (O_218,N_19014,N_19716);
xnor UO_219 (O_219,N_19748,N_19572);
xnor UO_220 (O_220,N_19609,N_19427);
nor UO_221 (O_221,N_19837,N_19518);
nand UO_222 (O_222,N_19769,N_19681);
nand UO_223 (O_223,N_19708,N_19969);
and UO_224 (O_224,N_19236,N_19940);
xor UO_225 (O_225,N_19610,N_19870);
nor UO_226 (O_226,N_19476,N_19785);
nand UO_227 (O_227,N_19310,N_19034);
or UO_228 (O_228,N_19268,N_19918);
xor UO_229 (O_229,N_19879,N_19892);
xnor UO_230 (O_230,N_19482,N_19535);
and UO_231 (O_231,N_19598,N_19671);
or UO_232 (O_232,N_19225,N_19985);
nor UO_233 (O_233,N_19848,N_19010);
or UO_234 (O_234,N_19766,N_19206);
nor UO_235 (O_235,N_19353,N_19004);
or UO_236 (O_236,N_19947,N_19734);
or UO_237 (O_237,N_19456,N_19198);
xnor UO_238 (O_238,N_19171,N_19172);
nand UO_239 (O_239,N_19743,N_19412);
nand UO_240 (O_240,N_19631,N_19581);
xnor UO_241 (O_241,N_19336,N_19915);
xor UO_242 (O_242,N_19788,N_19073);
and UO_243 (O_243,N_19858,N_19248);
nand UO_244 (O_244,N_19514,N_19163);
xor UO_245 (O_245,N_19303,N_19575);
nand UO_246 (O_246,N_19063,N_19519);
xor UO_247 (O_247,N_19595,N_19494);
nor UO_248 (O_248,N_19819,N_19526);
or UO_249 (O_249,N_19674,N_19712);
and UO_250 (O_250,N_19967,N_19102);
and UO_251 (O_251,N_19280,N_19108);
nor UO_252 (O_252,N_19325,N_19721);
nor UO_253 (O_253,N_19381,N_19946);
xnor UO_254 (O_254,N_19872,N_19216);
nand UO_255 (O_255,N_19868,N_19850);
and UO_256 (O_256,N_19269,N_19682);
nand UO_257 (O_257,N_19846,N_19466);
or UO_258 (O_258,N_19642,N_19834);
or UO_259 (O_259,N_19265,N_19080);
nor UO_260 (O_260,N_19226,N_19188);
and UO_261 (O_261,N_19127,N_19440);
xor UO_262 (O_262,N_19296,N_19475);
nand UO_263 (O_263,N_19652,N_19897);
nand UO_264 (O_264,N_19069,N_19676);
nand UO_265 (O_265,N_19640,N_19641);
nand UO_266 (O_266,N_19591,N_19568);
and UO_267 (O_267,N_19739,N_19284);
and UO_268 (O_268,N_19285,N_19635);
nor UO_269 (O_269,N_19364,N_19404);
or UO_270 (O_270,N_19561,N_19701);
nor UO_271 (O_271,N_19805,N_19042);
nand UO_272 (O_272,N_19215,N_19811);
xnor UO_273 (O_273,N_19416,N_19733);
and UO_274 (O_274,N_19410,N_19078);
xnor UO_275 (O_275,N_19873,N_19820);
nor UO_276 (O_276,N_19002,N_19934);
or UO_277 (O_277,N_19626,N_19775);
xnor UO_278 (O_278,N_19311,N_19637);
xor UO_279 (O_279,N_19883,N_19513);
xor UO_280 (O_280,N_19667,N_19123);
nor UO_281 (O_281,N_19307,N_19761);
nor UO_282 (O_282,N_19470,N_19106);
xor UO_283 (O_283,N_19194,N_19890);
or UO_284 (O_284,N_19829,N_19393);
xnor UO_285 (O_285,N_19049,N_19889);
xnor UO_286 (O_286,N_19170,N_19193);
xor UO_287 (O_287,N_19625,N_19576);
nand UO_288 (O_288,N_19231,N_19208);
or UO_289 (O_289,N_19156,N_19881);
nand UO_290 (O_290,N_19319,N_19954);
nor UO_291 (O_291,N_19501,N_19442);
xor UO_292 (O_292,N_19149,N_19960);
and UO_293 (O_293,N_19176,N_19976);
xnor UO_294 (O_294,N_19673,N_19463);
and UO_295 (O_295,N_19260,N_19789);
nor UO_296 (O_296,N_19750,N_19185);
or UO_297 (O_297,N_19432,N_19354);
nand UO_298 (O_298,N_19158,N_19842);
or UO_299 (O_299,N_19831,N_19633);
or UO_300 (O_300,N_19038,N_19360);
or UO_301 (O_301,N_19247,N_19068);
nor UO_302 (O_302,N_19768,N_19021);
and UO_303 (O_303,N_19052,N_19203);
nor UO_304 (O_304,N_19912,N_19800);
xor UO_305 (O_305,N_19620,N_19783);
and UO_306 (O_306,N_19932,N_19141);
xor UO_307 (O_307,N_19181,N_19684);
xnor UO_308 (O_308,N_19955,N_19374);
nor UO_309 (O_309,N_19668,N_19489);
nor UO_310 (O_310,N_19663,N_19047);
xor UO_311 (O_311,N_19143,N_19546);
or UO_312 (O_312,N_19046,N_19150);
or UO_313 (O_313,N_19510,N_19001);
or UO_314 (O_314,N_19100,N_19192);
xnor UO_315 (O_315,N_19801,N_19856);
or UO_316 (O_316,N_19414,N_19629);
xor UO_317 (O_317,N_19986,N_19896);
xnor UO_318 (O_318,N_19214,N_19421);
xor UO_319 (O_319,N_19948,N_19196);
nand UO_320 (O_320,N_19253,N_19415);
or UO_321 (O_321,N_19622,N_19026);
nand UO_322 (O_322,N_19951,N_19857);
nand UO_323 (O_323,N_19961,N_19147);
nor UO_324 (O_324,N_19189,N_19312);
xnor UO_325 (O_325,N_19616,N_19924);
nor UO_326 (O_326,N_19278,N_19817);
nand UO_327 (O_327,N_19573,N_19013);
and UO_328 (O_328,N_19406,N_19880);
nand UO_329 (O_329,N_19320,N_19096);
nor UO_330 (O_330,N_19740,N_19023);
and UO_331 (O_331,N_19362,N_19164);
nand UO_332 (O_332,N_19375,N_19401);
or UO_333 (O_333,N_19987,N_19045);
and UO_334 (O_334,N_19751,N_19966);
xnor UO_335 (O_335,N_19723,N_19390);
or UO_336 (O_336,N_19710,N_19562);
or UO_337 (O_337,N_19567,N_19016);
nor UO_338 (O_338,N_19359,N_19515);
nand UO_339 (O_339,N_19998,N_19826);
and UO_340 (O_340,N_19523,N_19057);
or UO_341 (O_341,N_19797,N_19397);
or UO_342 (O_342,N_19140,N_19477);
or UO_343 (O_343,N_19557,N_19331);
nand UO_344 (O_344,N_19101,N_19282);
nand UO_345 (O_345,N_19606,N_19338);
xnor UO_346 (O_346,N_19833,N_19024);
xor UO_347 (O_347,N_19983,N_19763);
and UO_348 (O_348,N_19554,N_19943);
xnor UO_349 (O_349,N_19520,N_19177);
or UO_350 (O_350,N_19504,N_19082);
or UO_351 (O_351,N_19818,N_19017);
nor UO_352 (O_352,N_19658,N_19455);
nor UO_353 (O_353,N_19975,N_19105);
nand UO_354 (O_354,N_19793,N_19352);
or UO_355 (O_355,N_19937,N_19919);
and UO_356 (O_356,N_19600,N_19980);
nand UO_357 (O_357,N_19645,N_19405);
nor UO_358 (O_358,N_19259,N_19485);
or UO_359 (O_359,N_19715,N_19128);
xor UO_360 (O_360,N_19493,N_19604);
xnor UO_361 (O_361,N_19322,N_19810);
or UO_362 (O_362,N_19088,N_19607);
xnor UO_363 (O_363,N_19720,N_19388);
nand UO_364 (O_364,N_19274,N_19076);
and UO_365 (O_365,N_19495,N_19847);
nand UO_366 (O_366,N_19500,N_19368);
nand UO_367 (O_367,N_19585,N_19446);
or UO_368 (O_368,N_19335,N_19521);
or UO_369 (O_369,N_19222,N_19990);
and UO_370 (O_370,N_19603,N_19283);
nor UO_371 (O_371,N_19656,N_19584);
or UO_372 (O_372,N_19473,N_19299);
xor UO_373 (O_373,N_19155,N_19851);
nor UO_374 (O_374,N_19670,N_19508);
or UO_375 (O_375,N_19306,N_19503);
and UO_376 (O_376,N_19139,N_19389);
nand UO_377 (O_377,N_19531,N_19458);
and UO_378 (O_378,N_19119,N_19677);
xor UO_379 (O_379,N_19587,N_19240);
xnor UO_380 (O_380,N_19694,N_19540);
and UO_381 (O_381,N_19935,N_19457);
nand UO_382 (O_382,N_19802,N_19261);
nor UO_383 (O_383,N_19471,N_19221);
or UO_384 (O_384,N_19382,N_19738);
or UO_385 (O_385,N_19228,N_19795);
and UO_386 (O_386,N_19997,N_19323);
and UO_387 (O_387,N_19118,N_19304);
nor UO_388 (O_388,N_19938,N_19027);
and UO_389 (O_389,N_19000,N_19386);
xnor UO_390 (O_390,N_19281,N_19054);
nor UO_391 (O_391,N_19726,N_19272);
nor UO_392 (O_392,N_19577,N_19326);
nand UO_393 (O_393,N_19346,N_19929);
or UO_394 (O_394,N_19431,N_19812);
or UO_395 (O_395,N_19190,N_19728);
nor UO_396 (O_396,N_19689,N_19329);
xnor UO_397 (O_397,N_19601,N_19145);
or UO_398 (O_398,N_19341,N_19895);
nor UO_399 (O_399,N_19060,N_19230);
nor UO_400 (O_400,N_19428,N_19053);
or UO_401 (O_401,N_19630,N_19649);
and UO_402 (O_402,N_19711,N_19031);
nand UO_403 (O_403,N_19876,N_19841);
or UO_404 (O_404,N_19569,N_19424);
or UO_405 (O_405,N_19898,N_19302);
xor UO_406 (O_406,N_19090,N_19749);
and UO_407 (O_407,N_19565,N_19286);
xor UO_408 (O_408,N_19356,N_19977);
nor UO_409 (O_409,N_19773,N_19571);
xor UO_410 (O_410,N_19617,N_19588);
xnor UO_411 (O_411,N_19061,N_19578);
nand UO_412 (O_412,N_19277,N_19210);
or UO_413 (O_413,N_19436,N_19107);
xnor UO_414 (O_414,N_19041,N_19729);
and UO_415 (O_415,N_19916,N_19638);
nand UO_416 (O_416,N_19882,N_19020);
and UO_417 (O_417,N_19792,N_19464);
or UO_418 (O_418,N_19234,N_19843);
and UO_419 (O_419,N_19347,N_19646);
nand UO_420 (O_420,N_19235,N_19543);
nand UO_421 (O_421,N_19365,N_19103);
nand UO_422 (O_422,N_19434,N_19413);
xor UO_423 (O_423,N_19564,N_19511);
nand UO_424 (O_424,N_19688,N_19539);
nor UO_425 (O_425,N_19925,N_19309);
or UO_426 (O_426,N_19849,N_19358);
xnor UO_427 (O_427,N_19367,N_19970);
or UO_428 (O_428,N_19643,N_19217);
and UO_429 (O_429,N_19462,N_19070);
nand UO_430 (O_430,N_19887,N_19776);
or UO_431 (O_431,N_19654,N_19396);
xnor UO_432 (O_432,N_19399,N_19091);
or UO_433 (O_433,N_19904,N_19770);
nand UO_434 (O_434,N_19067,N_19279);
nor UO_435 (O_435,N_19547,N_19449);
xnor UO_436 (O_436,N_19661,N_19488);
nand UO_437 (O_437,N_19725,N_19963);
nand UO_438 (O_438,N_19220,N_19059);
and UO_439 (O_439,N_19717,N_19300);
nor UO_440 (O_440,N_19690,N_19182);
nor UO_441 (O_441,N_19146,N_19122);
xor UO_442 (O_442,N_19238,N_19722);
xnor UO_443 (O_443,N_19828,N_19109);
nor UO_444 (O_444,N_19813,N_19212);
or UO_445 (O_445,N_19704,N_19430);
nor UO_446 (O_446,N_19909,N_19089);
nor UO_447 (O_447,N_19648,N_19223);
nor UO_448 (O_448,N_19907,N_19914);
and UO_449 (O_449,N_19845,N_19348);
or UO_450 (O_450,N_19700,N_19608);
xor UO_451 (O_451,N_19862,N_19894);
nand UO_452 (O_452,N_19378,N_19706);
nor UO_453 (O_453,N_19778,N_19294);
xor UO_454 (O_454,N_19394,N_19486);
nor UO_455 (O_455,N_19205,N_19315);
nor UO_456 (O_456,N_19759,N_19509);
and UO_457 (O_457,N_19232,N_19142);
xnor UO_458 (O_458,N_19542,N_19964);
and UO_459 (O_459,N_19048,N_19425);
or UO_460 (O_460,N_19313,N_19373);
nor UO_461 (O_461,N_19559,N_19345);
nand UO_462 (O_462,N_19239,N_19187);
and UO_463 (O_463,N_19165,N_19517);
nor UO_464 (O_464,N_19901,N_19258);
nand UO_465 (O_465,N_19008,N_19092);
or UO_466 (O_466,N_19798,N_19173);
and UO_467 (O_467,N_19332,N_19703);
and UO_468 (O_468,N_19611,N_19241);
and UO_469 (O_469,N_19877,N_19133);
xnor UO_470 (O_470,N_19110,N_19126);
or UO_471 (O_471,N_19003,N_19612);
and UO_472 (O_472,N_19317,N_19774);
nor UO_473 (O_473,N_19996,N_19589);
or UO_474 (O_474,N_19499,N_19267);
xnor UO_475 (O_475,N_19628,N_19200);
nor UO_476 (O_476,N_19746,N_19920);
nor UO_477 (O_477,N_19921,N_19154);
nand UO_478 (O_478,N_19333,N_19566);
nand UO_479 (O_479,N_19583,N_19095);
and UO_480 (O_480,N_19702,N_19293);
nor UO_481 (O_481,N_19363,N_19787);
xor UO_482 (O_482,N_19218,N_19804);
xor UO_483 (O_483,N_19693,N_19602);
or UO_484 (O_484,N_19991,N_19621);
nor UO_485 (O_485,N_19989,N_19025);
and UO_486 (O_486,N_19839,N_19490);
xnor UO_487 (O_487,N_19484,N_19350);
xor UO_488 (O_488,N_19379,N_19952);
xor UO_489 (O_489,N_19418,N_19824);
nand UO_490 (O_490,N_19264,N_19295);
or UO_491 (O_491,N_19467,N_19250);
or UO_492 (O_492,N_19448,N_19478);
and UO_493 (O_493,N_19978,N_19030);
nand UO_494 (O_494,N_19885,N_19691);
nand UO_495 (O_495,N_19039,N_19211);
nor UO_496 (O_496,N_19445,N_19655);
and UO_497 (O_497,N_19344,N_19233);
nand UO_498 (O_498,N_19807,N_19886);
and UO_499 (O_499,N_19124,N_19032);
and UO_500 (O_500,N_19782,N_19961);
xor UO_501 (O_501,N_19960,N_19338);
nand UO_502 (O_502,N_19940,N_19838);
or UO_503 (O_503,N_19685,N_19903);
or UO_504 (O_504,N_19884,N_19668);
or UO_505 (O_505,N_19272,N_19243);
nor UO_506 (O_506,N_19707,N_19745);
nor UO_507 (O_507,N_19669,N_19329);
nor UO_508 (O_508,N_19637,N_19706);
xnor UO_509 (O_509,N_19413,N_19411);
xor UO_510 (O_510,N_19574,N_19799);
nor UO_511 (O_511,N_19939,N_19393);
or UO_512 (O_512,N_19573,N_19808);
nand UO_513 (O_513,N_19212,N_19020);
and UO_514 (O_514,N_19525,N_19078);
and UO_515 (O_515,N_19661,N_19643);
nand UO_516 (O_516,N_19688,N_19698);
xor UO_517 (O_517,N_19949,N_19053);
nor UO_518 (O_518,N_19965,N_19672);
and UO_519 (O_519,N_19294,N_19331);
or UO_520 (O_520,N_19108,N_19246);
or UO_521 (O_521,N_19858,N_19095);
or UO_522 (O_522,N_19899,N_19666);
nand UO_523 (O_523,N_19049,N_19104);
nand UO_524 (O_524,N_19455,N_19652);
or UO_525 (O_525,N_19334,N_19302);
nand UO_526 (O_526,N_19483,N_19723);
or UO_527 (O_527,N_19226,N_19988);
nor UO_528 (O_528,N_19524,N_19380);
nor UO_529 (O_529,N_19640,N_19556);
nand UO_530 (O_530,N_19057,N_19185);
and UO_531 (O_531,N_19834,N_19891);
xor UO_532 (O_532,N_19106,N_19803);
and UO_533 (O_533,N_19154,N_19212);
xnor UO_534 (O_534,N_19553,N_19499);
and UO_535 (O_535,N_19662,N_19142);
xor UO_536 (O_536,N_19834,N_19283);
nand UO_537 (O_537,N_19309,N_19217);
and UO_538 (O_538,N_19095,N_19480);
nor UO_539 (O_539,N_19420,N_19312);
and UO_540 (O_540,N_19539,N_19400);
and UO_541 (O_541,N_19857,N_19343);
nor UO_542 (O_542,N_19521,N_19635);
and UO_543 (O_543,N_19542,N_19359);
or UO_544 (O_544,N_19317,N_19984);
nor UO_545 (O_545,N_19583,N_19063);
nand UO_546 (O_546,N_19590,N_19066);
xnor UO_547 (O_547,N_19190,N_19451);
and UO_548 (O_548,N_19404,N_19424);
xor UO_549 (O_549,N_19005,N_19156);
nand UO_550 (O_550,N_19835,N_19468);
nand UO_551 (O_551,N_19989,N_19843);
nor UO_552 (O_552,N_19736,N_19789);
xnor UO_553 (O_553,N_19464,N_19279);
xnor UO_554 (O_554,N_19354,N_19385);
or UO_555 (O_555,N_19858,N_19107);
or UO_556 (O_556,N_19025,N_19098);
xnor UO_557 (O_557,N_19951,N_19077);
and UO_558 (O_558,N_19725,N_19529);
nand UO_559 (O_559,N_19751,N_19984);
and UO_560 (O_560,N_19776,N_19162);
and UO_561 (O_561,N_19425,N_19771);
nor UO_562 (O_562,N_19362,N_19064);
and UO_563 (O_563,N_19438,N_19580);
or UO_564 (O_564,N_19460,N_19625);
or UO_565 (O_565,N_19592,N_19400);
xor UO_566 (O_566,N_19057,N_19333);
xor UO_567 (O_567,N_19310,N_19779);
nor UO_568 (O_568,N_19232,N_19851);
nand UO_569 (O_569,N_19868,N_19212);
or UO_570 (O_570,N_19559,N_19856);
or UO_571 (O_571,N_19125,N_19174);
xnor UO_572 (O_572,N_19178,N_19967);
nand UO_573 (O_573,N_19130,N_19358);
xnor UO_574 (O_574,N_19734,N_19922);
nand UO_575 (O_575,N_19820,N_19328);
and UO_576 (O_576,N_19846,N_19728);
nand UO_577 (O_577,N_19062,N_19817);
nand UO_578 (O_578,N_19145,N_19418);
nand UO_579 (O_579,N_19590,N_19551);
or UO_580 (O_580,N_19205,N_19183);
or UO_581 (O_581,N_19899,N_19364);
nand UO_582 (O_582,N_19745,N_19086);
and UO_583 (O_583,N_19779,N_19816);
xor UO_584 (O_584,N_19299,N_19079);
xnor UO_585 (O_585,N_19932,N_19824);
xor UO_586 (O_586,N_19368,N_19590);
or UO_587 (O_587,N_19087,N_19816);
and UO_588 (O_588,N_19749,N_19682);
or UO_589 (O_589,N_19997,N_19448);
and UO_590 (O_590,N_19691,N_19663);
nand UO_591 (O_591,N_19969,N_19008);
or UO_592 (O_592,N_19657,N_19859);
and UO_593 (O_593,N_19170,N_19006);
and UO_594 (O_594,N_19791,N_19403);
xnor UO_595 (O_595,N_19977,N_19769);
nor UO_596 (O_596,N_19328,N_19787);
or UO_597 (O_597,N_19511,N_19050);
nand UO_598 (O_598,N_19862,N_19498);
nor UO_599 (O_599,N_19629,N_19219);
and UO_600 (O_600,N_19131,N_19982);
or UO_601 (O_601,N_19305,N_19299);
nand UO_602 (O_602,N_19843,N_19465);
nand UO_603 (O_603,N_19281,N_19078);
xnor UO_604 (O_604,N_19547,N_19111);
and UO_605 (O_605,N_19383,N_19256);
or UO_606 (O_606,N_19446,N_19540);
and UO_607 (O_607,N_19539,N_19403);
xnor UO_608 (O_608,N_19867,N_19494);
or UO_609 (O_609,N_19363,N_19390);
or UO_610 (O_610,N_19407,N_19610);
nor UO_611 (O_611,N_19140,N_19302);
xnor UO_612 (O_612,N_19239,N_19967);
and UO_613 (O_613,N_19057,N_19539);
and UO_614 (O_614,N_19553,N_19159);
nor UO_615 (O_615,N_19635,N_19889);
and UO_616 (O_616,N_19765,N_19461);
nand UO_617 (O_617,N_19083,N_19231);
or UO_618 (O_618,N_19240,N_19970);
xor UO_619 (O_619,N_19842,N_19476);
or UO_620 (O_620,N_19388,N_19742);
xor UO_621 (O_621,N_19980,N_19799);
nor UO_622 (O_622,N_19250,N_19016);
xor UO_623 (O_623,N_19253,N_19586);
nand UO_624 (O_624,N_19599,N_19985);
and UO_625 (O_625,N_19657,N_19145);
and UO_626 (O_626,N_19364,N_19897);
and UO_627 (O_627,N_19188,N_19143);
or UO_628 (O_628,N_19216,N_19557);
or UO_629 (O_629,N_19932,N_19804);
nand UO_630 (O_630,N_19993,N_19542);
xor UO_631 (O_631,N_19809,N_19598);
or UO_632 (O_632,N_19263,N_19162);
or UO_633 (O_633,N_19436,N_19926);
nor UO_634 (O_634,N_19136,N_19137);
nand UO_635 (O_635,N_19109,N_19863);
and UO_636 (O_636,N_19169,N_19838);
nand UO_637 (O_637,N_19910,N_19687);
nor UO_638 (O_638,N_19572,N_19194);
xor UO_639 (O_639,N_19403,N_19230);
xor UO_640 (O_640,N_19164,N_19535);
or UO_641 (O_641,N_19039,N_19894);
nor UO_642 (O_642,N_19991,N_19172);
or UO_643 (O_643,N_19211,N_19818);
xnor UO_644 (O_644,N_19444,N_19412);
or UO_645 (O_645,N_19852,N_19563);
xor UO_646 (O_646,N_19635,N_19605);
or UO_647 (O_647,N_19834,N_19552);
and UO_648 (O_648,N_19785,N_19548);
nor UO_649 (O_649,N_19551,N_19018);
or UO_650 (O_650,N_19160,N_19701);
or UO_651 (O_651,N_19833,N_19352);
or UO_652 (O_652,N_19269,N_19011);
xnor UO_653 (O_653,N_19837,N_19367);
nand UO_654 (O_654,N_19997,N_19009);
and UO_655 (O_655,N_19527,N_19606);
or UO_656 (O_656,N_19387,N_19381);
nand UO_657 (O_657,N_19167,N_19540);
and UO_658 (O_658,N_19357,N_19388);
nand UO_659 (O_659,N_19465,N_19906);
and UO_660 (O_660,N_19623,N_19571);
xnor UO_661 (O_661,N_19318,N_19984);
xnor UO_662 (O_662,N_19663,N_19153);
and UO_663 (O_663,N_19382,N_19180);
xor UO_664 (O_664,N_19795,N_19747);
and UO_665 (O_665,N_19088,N_19781);
and UO_666 (O_666,N_19255,N_19946);
and UO_667 (O_667,N_19893,N_19000);
and UO_668 (O_668,N_19646,N_19092);
or UO_669 (O_669,N_19110,N_19509);
nand UO_670 (O_670,N_19107,N_19757);
nor UO_671 (O_671,N_19363,N_19921);
nand UO_672 (O_672,N_19231,N_19644);
or UO_673 (O_673,N_19845,N_19855);
nand UO_674 (O_674,N_19551,N_19331);
xnor UO_675 (O_675,N_19217,N_19001);
and UO_676 (O_676,N_19057,N_19566);
xor UO_677 (O_677,N_19261,N_19102);
or UO_678 (O_678,N_19937,N_19450);
and UO_679 (O_679,N_19804,N_19518);
or UO_680 (O_680,N_19848,N_19273);
nor UO_681 (O_681,N_19267,N_19153);
nand UO_682 (O_682,N_19391,N_19412);
nor UO_683 (O_683,N_19432,N_19312);
or UO_684 (O_684,N_19868,N_19956);
nand UO_685 (O_685,N_19519,N_19757);
or UO_686 (O_686,N_19777,N_19710);
nor UO_687 (O_687,N_19263,N_19663);
or UO_688 (O_688,N_19349,N_19875);
xnor UO_689 (O_689,N_19381,N_19834);
nor UO_690 (O_690,N_19089,N_19611);
or UO_691 (O_691,N_19697,N_19461);
or UO_692 (O_692,N_19506,N_19955);
or UO_693 (O_693,N_19096,N_19938);
or UO_694 (O_694,N_19282,N_19458);
nor UO_695 (O_695,N_19330,N_19742);
and UO_696 (O_696,N_19673,N_19942);
and UO_697 (O_697,N_19466,N_19998);
nor UO_698 (O_698,N_19923,N_19498);
nor UO_699 (O_699,N_19393,N_19858);
nand UO_700 (O_700,N_19121,N_19203);
or UO_701 (O_701,N_19406,N_19263);
and UO_702 (O_702,N_19710,N_19635);
xnor UO_703 (O_703,N_19090,N_19696);
xor UO_704 (O_704,N_19166,N_19631);
or UO_705 (O_705,N_19140,N_19115);
xnor UO_706 (O_706,N_19129,N_19883);
and UO_707 (O_707,N_19400,N_19726);
xor UO_708 (O_708,N_19787,N_19345);
or UO_709 (O_709,N_19934,N_19140);
xnor UO_710 (O_710,N_19635,N_19807);
and UO_711 (O_711,N_19371,N_19063);
or UO_712 (O_712,N_19465,N_19938);
nand UO_713 (O_713,N_19804,N_19860);
or UO_714 (O_714,N_19145,N_19474);
xnor UO_715 (O_715,N_19275,N_19169);
xor UO_716 (O_716,N_19055,N_19713);
and UO_717 (O_717,N_19887,N_19726);
and UO_718 (O_718,N_19806,N_19319);
and UO_719 (O_719,N_19341,N_19206);
nor UO_720 (O_720,N_19856,N_19402);
and UO_721 (O_721,N_19837,N_19400);
and UO_722 (O_722,N_19181,N_19220);
or UO_723 (O_723,N_19444,N_19144);
xor UO_724 (O_724,N_19434,N_19809);
xnor UO_725 (O_725,N_19847,N_19433);
or UO_726 (O_726,N_19417,N_19366);
nand UO_727 (O_727,N_19783,N_19152);
and UO_728 (O_728,N_19413,N_19585);
nor UO_729 (O_729,N_19408,N_19979);
or UO_730 (O_730,N_19251,N_19188);
nand UO_731 (O_731,N_19749,N_19196);
or UO_732 (O_732,N_19230,N_19914);
and UO_733 (O_733,N_19505,N_19328);
nor UO_734 (O_734,N_19379,N_19355);
or UO_735 (O_735,N_19273,N_19350);
or UO_736 (O_736,N_19666,N_19898);
nand UO_737 (O_737,N_19332,N_19899);
or UO_738 (O_738,N_19234,N_19109);
or UO_739 (O_739,N_19184,N_19638);
nor UO_740 (O_740,N_19893,N_19844);
nand UO_741 (O_741,N_19292,N_19537);
xor UO_742 (O_742,N_19552,N_19872);
nand UO_743 (O_743,N_19915,N_19085);
or UO_744 (O_744,N_19675,N_19847);
xor UO_745 (O_745,N_19915,N_19643);
nor UO_746 (O_746,N_19896,N_19081);
nand UO_747 (O_747,N_19119,N_19998);
nor UO_748 (O_748,N_19547,N_19454);
nand UO_749 (O_749,N_19373,N_19273);
xnor UO_750 (O_750,N_19193,N_19157);
nand UO_751 (O_751,N_19079,N_19130);
xor UO_752 (O_752,N_19905,N_19762);
nor UO_753 (O_753,N_19142,N_19031);
or UO_754 (O_754,N_19483,N_19040);
nor UO_755 (O_755,N_19892,N_19760);
and UO_756 (O_756,N_19415,N_19685);
xor UO_757 (O_757,N_19272,N_19382);
or UO_758 (O_758,N_19905,N_19182);
xnor UO_759 (O_759,N_19222,N_19660);
or UO_760 (O_760,N_19144,N_19177);
nand UO_761 (O_761,N_19356,N_19885);
nor UO_762 (O_762,N_19646,N_19381);
xnor UO_763 (O_763,N_19907,N_19129);
or UO_764 (O_764,N_19604,N_19223);
nor UO_765 (O_765,N_19907,N_19112);
and UO_766 (O_766,N_19390,N_19121);
xnor UO_767 (O_767,N_19797,N_19200);
or UO_768 (O_768,N_19825,N_19696);
or UO_769 (O_769,N_19007,N_19540);
and UO_770 (O_770,N_19716,N_19250);
and UO_771 (O_771,N_19969,N_19678);
xor UO_772 (O_772,N_19370,N_19947);
nand UO_773 (O_773,N_19076,N_19158);
nand UO_774 (O_774,N_19404,N_19250);
xnor UO_775 (O_775,N_19600,N_19569);
and UO_776 (O_776,N_19288,N_19709);
or UO_777 (O_777,N_19252,N_19575);
nor UO_778 (O_778,N_19251,N_19374);
or UO_779 (O_779,N_19263,N_19008);
nor UO_780 (O_780,N_19502,N_19631);
xnor UO_781 (O_781,N_19734,N_19774);
nand UO_782 (O_782,N_19484,N_19964);
and UO_783 (O_783,N_19586,N_19800);
nor UO_784 (O_784,N_19290,N_19542);
nand UO_785 (O_785,N_19703,N_19179);
xnor UO_786 (O_786,N_19532,N_19745);
or UO_787 (O_787,N_19677,N_19649);
and UO_788 (O_788,N_19215,N_19499);
and UO_789 (O_789,N_19531,N_19774);
or UO_790 (O_790,N_19051,N_19986);
and UO_791 (O_791,N_19626,N_19228);
xnor UO_792 (O_792,N_19890,N_19616);
nand UO_793 (O_793,N_19699,N_19138);
or UO_794 (O_794,N_19183,N_19696);
nand UO_795 (O_795,N_19732,N_19443);
nor UO_796 (O_796,N_19438,N_19666);
and UO_797 (O_797,N_19215,N_19626);
and UO_798 (O_798,N_19277,N_19826);
and UO_799 (O_799,N_19522,N_19272);
and UO_800 (O_800,N_19547,N_19438);
nor UO_801 (O_801,N_19688,N_19770);
nor UO_802 (O_802,N_19120,N_19881);
xnor UO_803 (O_803,N_19398,N_19751);
or UO_804 (O_804,N_19373,N_19386);
xnor UO_805 (O_805,N_19593,N_19797);
and UO_806 (O_806,N_19083,N_19618);
nor UO_807 (O_807,N_19887,N_19184);
nand UO_808 (O_808,N_19542,N_19270);
or UO_809 (O_809,N_19563,N_19288);
nor UO_810 (O_810,N_19876,N_19474);
xnor UO_811 (O_811,N_19112,N_19714);
nor UO_812 (O_812,N_19617,N_19740);
nor UO_813 (O_813,N_19778,N_19459);
nor UO_814 (O_814,N_19383,N_19974);
xor UO_815 (O_815,N_19563,N_19602);
xnor UO_816 (O_816,N_19179,N_19607);
nand UO_817 (O_817,N_19094,N_19564);
xor UO_818 (O_818,N_19212,N_19254);
or UO_819 (O_819,N_19133,N_19495);
nor UO_820 (O_820,N_19133,N_19935);
nand UO_821 (O_821,N_19416,N_19961);
and UO_822 (O_822,N_19501,N_19627);
xor UO_823 (O_823,N_19853,N_19409);
nor UO_824 (O_824,N_19442,N_19015);
or UO_825 (O_825,N_19576,N_19154);
or UO_826 (O_826,N_19094,N_19776);
and UO_827 (O_827,N_19365,N_19083);
or UO_828 (O_828,N_19342,N_19360);
nor UO_829 (O_829,N_19093,N_19444);
xnor UO_830 (O_830,N_19350,N_19440);
nand UO_831 (O_831,N_19127,N_19182);
nor UO_832 (O_832,N_19190,N_19347);
or UO_833 (O_833,N_19114,N_19751);
nor UO_834 (O_834,N_19173,N_19399);
or UO_835 (O_835,N_19955,N_19534);
nor UO_836 (O_836,N_19185,N_19573);
xnor UO_837 (O_837,N_19142,N_19069);
xnor UO_838 (O_838,N_19838,N_19369);
xor UO_839 (O_839,N_19564,N_19768);
and UO_840 (O_840,N_19378,N_19570);
xnor UO_841 (O_841,N_19651,N_19366);
nand UO_842 (O_842,N_19383,N_19586);
and UO_843 (O_843,N_19176,N_19356);
and UO_844 (O_844,N_19280,N_19272);
or UO_845 (O_845,N_19398,N_19381);
and UO_846 (O_846,N_19029,N_19212);
or UO_847 (O_847,N_19475,N_19347);
nand UO_848 (O_848,N_19133,N_19872);
xor UO_849 (O_849,N_19804,N_19411);
and UO_850 (O_850,N_19150,N_19273);
and UO_851 (O_851,N_19107,N_19985);
nand UO_852 (O_852,N_19823,N_19293);
nand UO_853 (O_853,N_19169,N_19329);
nor UO_854 (O_854,N_19268,N_19181);
or UO_855 (O_855,N_19737,N_19646);
nor UO_856 (O_856,N_19446,N_19943);
xor UO_857 (O_857,N_19126,N_19243);
nand UO_858 (O_858,N_19999,N_19956);
xnor UO_859 (O_859,N_19713,N_19146);
nand UO_860 (O_860,N_19385,N_19841);
or UO_861 (O_861,N_19453,N_19675);
nor UO_862 (O_862,N_19310,N_19624);
nand UO_863 (O_863,N_19879,N_19802);
or UO_864 (O_864,N_19655,N_19035);
nor UO_865 (O_865,N_19180,N_19591);
nand UO_866 (O_866,N_19448,N_19422);
nor UO_867 (O_867,N_19984,N_19989);
nand UO_868 (O_868,N_19633,N_19716);
and UO_869 (O_869,N_19550,N_19123);
nand UO_870 (O_870,N_19111,N_19181);
or UO_871 (O_871,N_19407,N_19139);
or UO_872 (O_872,N_19133,N_19200);
and UO_873 (O_873,N_19889,N_19059);
nor UO_874 (O_874,N_19061,N_19261);
and UO_875 (O_875,N_19709,N_19096);
xnor UO_876 (O_876,N_19743,N_19539);
and UO_877 (O_877,N_19717,N_19633);
xor UO_878 (O_878,N_19243,N_19283);
nor UO_879 (O_879,N_19009,N_19593);
nor UO_880 (O_880,N_19337,N_19489);
and UO_881 (O_881,N_19088,N_19574);
nand UO_882 (O_882,N_19537,N_19769);
nand UO_883 (O_883,N_19719,N_19379);
nor UO_884 (O_884,N_19536,N_19856);
xnor UO_885 (O_885,N_19347,N_19296);
nor UO_886 (O_886,N_19206,N_19443);
and UO_887 (O_887,N_19396,N_19126);
xnor UO_888 (O_888,N_19198,N_19741);
and UO_889 (O_889,N_19666,N_19089);
xnor UO_890 (O_890,N_19099,N_19572);
nor UO_891 (O_891,N_19530,N_19779);
xor UO_892 (O_892,N_19952,N_19720);
xnor UO_893 (O_893,N_19194,N_19948);
and UO_894 (O_894,N_19818,N_19347);
xor UO_895 (O_895,N_19437,N_19775);
or UO_896 (O_896,N_19285,N_19752);
nor UO_897 (O_897,N_19475,N_19495);
or UO_898 (O_898,N_19226,N_19903);
or UO_899 (O_899,N_19608,N_19928);
nand UO_900 (O_900,N_19633,N_19871);
nand UO_901 (O_901,N_19782,N_19275);
xnor UO_902 (O_902,N_19694,N_19464);
and UO_903 (O_903,N_19919,N_19655);
nor UO_904 (O_904,N_19068,N_19412);
or UO_905 (O_905,N_19118,N_19363);
nor UO_906 (O_906,N_19430,N_19988);
and UO_907 (O_907,N_19254,N_19240);
nand UO_908 (O_908,N_19462,N_19917);
nor UO_909 (O_909,N_19525,N_19775);
xor UO_910 (O_910,N_19674,N_19321);
nand UO_911 (O_911,N_19054,N_19824);
and UO_912 (O_912,N_19490,N_19703);
and UO_913 (O_913,N_19106,N_19709);
nand UO_914 (O_914,N_19035,N_19396);
nand UO_915 (O_915,N_19703,N_19187);
nor UO_916 (O_916,N_19096,N_19318);
or UO_917 (O_917,N_19335,N_19505);
xor UO_918 (O_918,N_19078,N_19602);
xor UO_919 (O_919,N_19152,N_19916);
xnor UO_920 (O_920,N_19041,N_19597);
and UO_921 (O_921,N_19279,N_19498);
nand UO_922 (O_922,N_19146,N_19123);
xor UO_923 (O_923,N_19386,N_19586);
nand UO_924 (O_924,N_19592,N_19165);
and UO_925 (O_925,N_19105,N_19595);
or UO_926 (O_926,N_19226,N_19339);
and UO_927 (O_927,N_19556,N_19695);
or UO_928 (O_928,N_19026,N_19762);
nand UO_929 (O_929,N_19428,N_19484);
or UO_930 (O_930,N_19315,N_19730);
and UO_931 (O_931,N_19612,N_19518);
nor UO_932 (O_932,N_19516,N_19931);
nand UO_933 (O_933,N_19575,N_19184);
or UO_934 (O_934,N_19949,N_19080);
or UO_935 (O_935,N_19383,N_19993);
nand UO_936 (O_936,N_19823,N_19981);
and UO_937 (O_937,N_19545,N_19268);
xnor UO_938 (O_938,N_19708,N_19831);
and UO_939 (O_939,N_19734,N_19458);
nor UO_940 (O_940,N_19801,N_19011);
nand UO_941 (O_941,N_19630,N_19205);
and UO_942 (O_942,N_19277,N_19624);
and UO_943 (O_943,N_19044,N_19325);
or UO_944 (O_944,N_19268,N_19358);
nor UO_945 (O_945,N_19254,N_19674);
nand UO_946 (O_946,N_19835,N_19488);
or UO_947 (O_947,N_19718,N_19964);
and UO_948 (O_948,N_19135,N_19423);
nand UO_949 (O_949,N_19047,N_19501);
nor UO_950 (O_950,N_19262,N_19010);
or UO_951 (O_951,N_19208,N_19159);
or UO_952 (O_952,N_19739,N_19797);
nand UO_953 (O_953,N_19559,N_19597);
nor UO_954 (O_954,N_19430,N_19414);
nand UO_955 (O_955,N_19063,N_19192);
nand UO_956 (O_956,N_19761,N_19265);
xor UO_957 (O_957,N_19902,N_19683);
nand UO_958 (O_958,N_19875,N_19964);
xnor UO_959 (O_959,N_19940,N_19929);
nor UO_960 (O_960,N_19120,N_19964);
nor UO_961 (O_961,N_19538,N_19584);
and UO_962 (O_962,N_19386,N_19516);
or UO_963 (O_963,N_19325,N_19939);
xnor UO_964 (O_964,N_19334,N_19784);
or UO_965 (O_965,N_19224,N_19338);
nor UO_966 (O_966,N_19008,N_19244);
and UO_967 (O_967,N_19669,N_19241);
nand UO_968 (O_968,N_19322,N_19527);
nand UO_969 (O_969,N_19059,N_19645);
and UO_970 (O_970,N_19644,N_19037);
and UO_971 (O_971,N_19339,N_19002);
xnor UO_972 (O_972,N_19306,N_19478);
nand UO_973 (O_973,N_19755,N_19788);
xor UO_974 (O_974,N_19632,N_19201);
nand UO_975 (O_975,N_19854,N_19897);
nand UO_976 (O_976,N_19494,N_19739);
and UO_977 (O_977,N_19491,N_19013);
xor UO_978 (O_978,N_19074,N_19830);
nand UO_979 (O_979,N_19492,N_19958);
xnor UO_980 (O_980,N_19109,N_19684);
and UO_981 (O_981,N_19280,N_19513);
xnor UO_982 (O_982,N_19479,N_19297);
nor UO_983 (O_983,N_19502,N_19785);
and UO_984 (O_984,N_19485,N_19652);
nand UO_985 (O_985,N_19067,N_19241);
and UO_986 (O_986,N_19396,N_19762);
nand UO_987 (O_987,N_19726,N_19751);
and UO_988 (O_988,N_19758,N_19665);
or UO_989 (O_989,N_19647,N_19382);
nor UO_990 (O_990,N_19992,N_19570);
and UO_991 (O_991,N_19635,N_19062);
nor UO_992 (O_992,N_19009,N_19018);
nand UO_993 (O_993,N_19291,N_19607);
nor UO_994 (O_994,N_19326,N_19823);
or UO_995 (O_995,N_19145,N_19955);
nor UO_996 (O_996,N_19756,N_19884);
nand UO_997 (O_997,N_19913,N_19162);
xnor UO_998 (O_998,N_19252,N_19309);
xor UO_999 (O_999,N_19396,N_19920);
nand UO_1000 (O_1000,N_19077,N_19821);
nand UO_1001 (O_1001,N_19501,N_19207);
or UO_1002 (O_1002,N_19423,N_19603);
nor UO_1003 (O_1003,N_19204,N_19393);
nor UO_1004 (O_1004,N_19532,N_19130);
and UO_1005 (O_1005,N_19696,N_19952);
xnor UO_1006 (O_1006,N_19841,N_19695);
nand UO_1007 (O_1007,N_19920,N_19382);
or UO_1008 (O_1008,N_19803,N_19797);
nand UO_1009 (O_1009,N_19807,N_19853);
xor UO_1010 (O_1010,N_19848,N_19604);
xor UO_1011 (O_1011,N_19688,N_19933);
or UO_1012 (O_1012,N_19876,N_19330);
nand UO_1013 (O_1013,N_19209,N_19728);
and UO_1014 (O_1014,N_19406,N_19155);
nand UO_1015 (O_1015,N_19221,N_19661);
or UO_1016 (O_1016,N_19444,N_19197);
xnor UO_1017 (O_1017,N_19081,N_19524);
nand UO_1018 (O_1018,N_19592,N_19229);
xnor UO_1019 (O_1019,N_19151,N_19056);
and UO_1020 (O_1020,N_19817,N_19241);
or UO_1021 (O_1021,N_19501,N_19947);
or UO_1022 (O_1022,N_19110,N_19899);
xor UO_1023 (O_1023,N_19488,N_19347);
nor UO_1024 (O_1024,N_19111,N_19053);
nor UO_1025 (O_1025,N_19902,N_19328);
nand UO_1026 (O_1026,N_19209,N_19163);
nand UO_1027 (O_1027,N_19974,N_19178);
and UO_1028 (O_1028,N_19768,N_19363);
nand UO_1029 (O_1029,N_19122,N_19108);
xnor UO_1030 (O_1030,N_19203,N_19782);
and UO_1031 (O_1031,N_19383,N_19151);
nor UO_1032 (O_1032,N_19939,N_19899);
xnor UO_1033 (O_1033,N_19732,N_19005);
nor UO_1034 (O_1034,N_19926,N_19388);
or UO_1035 (O_1035,N_19753,N_19940);
nor UO_1036 (O_1036,N_19286,N_19361);
xnor UO_1037 (O_1037,N_19359,N_19475);
or UO_1038 (O_1038,N_19715,N_19619);
or UO_1039 (O_1039,N_19175,N_19167);
or UO_1040 (O_1040,N_19076,N_19749);
xnor UO_1041 (O_1041,N_19033,N_19409);
and UO_1042 (O_1042,N_19702,N_19548);
or UO_1043 (O_1043,N_19938,N_19450);
nand UO_1044 (O_1044,N_19053,N_19010);
xnor UO_1045 (O_1045,N_19358,N_19438);
xor UO_1046 (O_1046,N_19345,N_19940);
xnor UO_1047 (O_1047,N_19056,N_19977);
nand UO_1048 (O_1048,N_19593,N_19467);
xnor UO_1049 (O_1049,N_19872,N_19305);
or UO_1050 (O_1050,N_19486,N_19206);
and UO_1051 (O_1051,N_19345,N_19041);
or UO_1052 (O_1052,N_19816,N_19387);
nor UO_1053 (O_1053,N_19117,N_19534);
nand UO_1054 (O_1054,N_19267,N_19511);
xnor UO_1055 (O_1055,N_19189,N_19725);
and UO_1056 (O_1056,N_19954,N_19786);
and UO_1057 (O_1057,N_19712,N_19786);
or UO_1058 (O_1058,N_19208,N_19063);
nand UO_1059 (O_1059,N_19161,N_19866);
or UO_1060 (O_1060,N_19502,N_19582);
xnor UO_1061 (O_1061,N_19596,N_19803);
nand UO_1062 (O_1062,N_19894,N_19916);
and UO_1063 (O_1063,N_19357,N_19118);
nand UO_1064 (O_1064,N_19677,N_19208);
or UO_1065 (O_1065,N_19745,N_19873);
or UO_1066 (O_1066,N_19480,N_19241);
nor UO_1067 (O_1067,N_19952,N_19924);
nand UO_1068 (O_1068,N_19985,N_19694);
and UO_1069 (O_1069,N_19549,N_19308);
xor UO_1070 (O_1070,N_19132,N_19967);
xor UO_1071 (O_1071,N_19292,N_19441);
xor UO_1072 (O_1072,N_19975,N_19908);
or UO_1073 (O_1073,N_19961,N_19505);
nand UO_1074 (O_1074,N_19383,N_19918);
nand UO_1075 (O_1075,N_19898,N_19405);
nor UO_1076 (O_1076,N_19109,N_19604);
and UO_1077 (O_1077,N_19763,N_19273);
nor UO_1078 (O_1078,N_19913,N_19165);
or UO_1079 (O_1079,N_19156,N_19832);
nor UO_1080 (O_1080,N_19285,N_19521);
nor UO_1081 (O_1081,N_19714,N_19015);
nor UO_1082 (O_1082,N_19494,N_19639);
and UO_1083 (O_1083,N_19378,N_19163);
nand UO_1084 (O_1084,N_19510,N_19595);
nand UO_1085 (O_1085,N_19271,N_19529);
nor UO_1086 (O_1086,N_19461,N_19134);
nand UO_1087 (O_1087,N_19591,N_19814);
xnor UO_1088 (O_1088,N_19317,N_19641);
xnor UO_1089 (O_1089,N_19845,N_19442);
or UO_1090 (O_1090,N_19401,N_19753);
nor UO_1091 (O_1091,N_19379,N_19171);
xnor UO_1092 (O_1092,N_19276,N_19430);
nor UO_1093 (O_1093,N_19478,N_19626);
or UO_1094 (O_1094,N_19759,N_19394);
nor UO_1095 (O_1095,N_19574,N_19508);
and UO_1096 (O_1096,N_19134,N_19109);
xor UO_1097 (O_1097,N_19888,N_19384);
and UO_1098 (O_1098,N_19564,N_19636);
or UO_1099 (O_1099,N_19651,N_19448);
nor UO_1100 (O_1100,N_19246,N_19882);
xor UO_1101 (O_1101,N_19084,N_19303);
xor UO_1102 (O_1102,N_19531,N_19208);
nand UO_1103 (O_1103,N_19208,N_19218);
nand UO_1104 (O_1104,N_19935,N_19025);
and UO_1105 (O_1105,N_19840,N_19664);
nand UO_1106 (O_1106,N_19718,N_19025);
or UO_1107 (O_1107,N_19055,N_19962);
and UO_1108 (O_1108,N_19643,N_19052);
nand UO_1109 (O_1109,N_19857,N_19048);
or UO_1110 (O_1110,N_19234,N_19974);
and UO_1111 (O_1111,N_19876,N_19324);
or UO_1112 (O_1112,N_19758,N_19754);
nor UO_1113 (O_1113,N_19816,N_19072);
and UO_1114 (O_1114,N_19963,N_19743);
xor UO_1115 (O_1115,N_19248,N_19514);
and UO_1116 (O_1116,N_19840,N_19100);
nor UO_1117 (O_1117,N_19653,N_19846);
or UO_1118 (O_1118,N_19668,N_19555);
or UO_1119 (O_1119,N_19770,N_19067);
and UO_1120 (O_1120,N_19927,N_19840);
and UO_1121 (O_1121,N_19368,N_19473);
or UO_1122 (O_1122,N_19856,N_19115);
nor UO_1123 (O_1123,N_19639,N_19343);
and UO_1124 (O_1124,N_19741,N_19582);
nand UO_1125 (O_1125,N_19709,N_19195);
xnor UO_1126 (O_1126,N_19126,N_19020);
nand UO_1127 (O_1127,N_19818,N_19509);
nand UO_1128 (O_1128,N_19617,N_19871);
nor UO_1129 (O_1129,N_19053,N_19558);
nor UO_1130 (O_1130,N_19570,N_19175);
nand UO_1131 (O_1131,N_19267,N_19658);
xnor UO_1132 (O_1132,N_19942,N_19094);
and UO_1133 (O_1133,N_19699,N_19295);
and UO_1134 (O_1134,N_19982,N_19586);
nor UO_1135 (O_1135,N_19263,N_19748);
or UO_1136 (O_1136,N_19519,N_19319);
and UO_1137 (O_1137,N_19525,N_19147);
nor UO_1138 (O_1138,N_19467,N_19473);
and UO_1139 (O_1139,N_19187,N_19382);
nor UO_1140 (O_1140,N_19616,N_19797);
xnor UO_1141 (O_1141,N_19535,N_19430);
or UO_1142 (O_1142,N_19386,N_19914);
and UO_1143 (O_1143,N_19476,N_19494);
nand UO_1144 (O_1144,N_19801,N_19205);
or UO_1145 (O_1145,N_19279,N_19410);
nand UO_1146 (O_1146,N_19058,N_19596);
nand UO_1147 (O_1147,N_19596,N_19096);
or UO_1148 (O_1148,N_19446,N_19853);
or UO_1149 (O_1149,N_19066,N_19026);
nand UO_1150 (O_1150,N_19158,N_19401);
and UO_1151 (O_1151,N_19268,N_19154);
nand UO_1152 (O_1152,N_19567,N_19568);
and UO_1153 (O_1153,N_19800,N_19836);
and UO_1154 (O_1154,N_19169,N_19189);
nand UO_1155 (O_1155,N_19453,N_19932);
or UO_1156 (O_1156,N_19009,N_19494);
xor UO_1157 (O_1157,N_19469,N_19354);
xor UO_1158 (O_1158,N_19470,N_19974);
nand UO_1159 (O_1159,N_19317,N_19888);
and UO_1160 (O_1160,N_19686,N_19762);
nor UO_1161 (O_1161,N_19353,N_19468);
or UO_1162 (O_1162,N_19705,N_19368);
nor UO_1163 (O_1163,N_19259,N_19793);
xnor UO_1164 (O_1164,N_19430,N_19954);
or UO_1165 (O_1165,N_19295,N_19895);
and UO_1166 (O_1166,N_19953,N_19209);
xor UO_1167 (O_1167,N_19873,N_19728);
or UO_1168 (O_1168,N_19072,N_19022);
or UO_1169 (O_1169,N_19595,N_19965);
or UO_1170 (O_1170,N_19147,N_19677);
nor UO_1171 (O_1171,N_19258,N_19900);
nand UO_1172 (O_1172,N_19468,N_19344);
xnor UO_1173 (O_1173,N_19164,N_19337);
nand UO_1174 (O_1174,N_19253,N_19649);
xor UO_1175 (O_1175,N_19756,N_19390);
or UO_1176 (O_1176,N_19013,N_19538);
xnor UO_1177 (O_1177,N_19539,N_19052);
and UO_1178 (O_1178,N_19391,N_19765);
nor UO_1179 (O_1179,N_19305,N_19814);
and UO_1180 (O_1180,N_19504,N_19041);
nor UO_1181 (O_1181,N_19093,N_19479);
xnor UO_1182 (O_1182,N_19598,N_19303);
xor UO_1183 (O_1183,N_19248,N_19998);
and UO_1184 (O_1184,N_19314,N_19109);
xor UO_1185 (O_1185,N_19499,N_19199);
and UO_1186 (O_1186,N_19002,N_19869);
or UO_1187 (O_1187,N_19046,N_19603);
nand UO_1188 (O_1188,N_19224,N_19359);
xnor UO_1189 (O_1189,N_19153,N_19555);
xnor UO_1190 (O_1190,N_19630,N_19437);
and UO_1191 (O_1191,N_19599,N_19009);
xnor UO_1192 (O_1192,N_19391,N_19310);
and UO_1193 (O_1193,N_19713,N_19965);
xor UO_1194 (O_1194,N_19623,N_19287);
or UO_1195 (O_1195,N_19359,N_19560);
and UO_1196 (O_1196,N_19857,N_19684);
or UO_1197 (O_1197,N_19422,N_19341);
xor UO_1198 (O_1198,N_19111,N_19827);
and UO_1199 (O_1199,N_19415,N_19798);
or UO_1200 (O_1200,N_19704,N_19047);
nor UO_1201 (O_1201,N_19089,N_19912);
nor UO_1202 (O_1202,N_19443,N_19028);
nor UO_1203 (O_1203,N_19690,N_19831);
or UO_1204 (O_1204,N_19092,N_19376);
and UO_1205 (O_1205,N_19778,N_19550);
nor UO_1206 (O_1206,N_19103,N_19565);
nor UO_1207 (O_1207,N_19555,N_19276);
and UO_1208 (O_1208,N_19896,N_19259);
nor UO_1209 (O_1209,N_19511,N_19256);
and UO_1210 (O_1210,N_19572,N_19228);
and UO_1211 (O_1211,N_19296,N_19476);
nand UO_1212 (O_1212,N_19454,N_19104);
nand UO_1213 (O_1213,N_19678,N_19631);
xor UO_1214 (O_1214,N_19887,N_19947);
nor UO_1215 (O_1215,N_19471,N_19131);
nor UO_1216 (O_1216,N_19929,N_19711);
or UO_1217 (O_1217,N_19645,N_19119);
nand UO_1218 (O_1218,N_19647,N_19735);
nand UO_1219 (O_1219,N_19424,N_19521);
nand UO_1220 (O_1220,N_19513,N_19414);
or UO_1221 (O_1221,N_19094,N_19957);
nor UO_1222 (O_1222,N_19026,N_19330);
or UO_1223 (O_1223,N_19715,N_19130);
or UO_1224 (O_1224,N_19421,N_19677);
or UO_1225 (O_1225,N_19972,N_19201);
nand UO_1226 (O_1226,N_19770,N_19778);
nand UO_1227 (O_1227,N_19996,N_19455);
nand UO_1228 (O_1228,N_19186,N_19429);
nor UO_1229 (O_1229,N_19159,N_19525);
and UO_1230 (O_1230,N_19781,N_19147);
or UO_1231 (O_1231,N_19222,N_19703);
or UO_1232 (O_1232,N_19585,N_19952);
xor UO_1233 (O_1233,N_19330,N_19601);
and UO_1234 (O_1234,N_19544,N_19596);
xnor UO_1235 (O_1235,N_19076,N_19110);
and UO_1236 (O_1236,N_19850,N_19799);
or UO_1237 (O_1237,N_19647,N_19989);
or UO_1238 (O_1238,N_19774,N_19432);
xor UO_1239 (O_1239,N_19319,N_19223);
or UO_1240 (O_1240,N_19945,N_19280);
nand UO_1241 (O_1241,N_19749,N_19093);
nor UO_1242 (O_1242,N_19960,N_19113);
or UO_1243 (O_1243,N_19058,N_19952);
or UO_1244 (O_1244,N_19098,N_19609);
or UO_1245 (O_1245,N_19575,N_19860);
and UO_1246 (O_1246,N_19647,N_19046);
nor UO_1247 (O_1247,N_19124,N_19722);
and UO_1248 (O_1248,N_19776,N_19133);
xor UO_1249 (O_1249,N_19545,N_19832);
xor UO_1250 (O_1250,N_19059,N_19199);
or UO_1251 (O_1251,N_19798,N_19698);
nand UO_1252 (O_1252,N_19545,N_19161);
and UO_1253 (O_1253,N_19318,N_19408);
xnor UO_1254 (O_1254,N_19290,N_19620);
nand UO_1255 (O_1255,N_19529,N_19853);
or UO_1256 (O_1256,N_19149,N_19865);
nor UO_1257 (O_1257,N_19392,N_19339);
xor UO_1258 (O_1258,N_19980,N_19885);
or UO_1259 (O_1259,N_19644,N_19213);
xnor UO_1260 (O_1260,N_19958,N_19060);
and UO_1261 (O_1261,N_19492,N_19277);
xnor UO_1262 (O_1262,N_19312,N_19647);
or UO_1263 (O_1263,N_19416,N_19660);
or UO_1264 (O_1264,N_19854,N_19693);
or UO_1265 (O_1265,N_19259,N_19868);
nand UO_1266 (O_1266,N_19007,N_19695);
nand UO_1267 (O_1267,N_19219,N_19578);
nand UO_1268 (O_1268,N_19242,N_19813);
xor UO_1269 (O_1269,N_19778,N_19178);
xnor UO_1270 (O_1270,N_19292,N_19598);
or UO_1271 (O_1271,N_19211,N_19036);
or UO_1272 (O_1272,N_19141,N_19534);
and UO_1273 (O_1273,N_19253,N_19905);
or UO_1274 (O_1274,N_19095,N_19654);
nor UO_1275 (O_1275,N_19514,N_19431);
nor UO_1276 (O_1276,N_19993,N_19130);
nand UO_1277 (O_1277,N_19540,N_19731);
xnor UO_1278 (O_1278,N_19549,N_19654);
nor UO_1279 (O_1279,N_19380,N_19289);
and UO_1280 (O_1280,N_19426,N_19126);
nand UO_1281 (O_1281,N_19967,N_19678);
nor UO_1282 (O_1282,N_19148,N_19734);
nand UO_1283 (O_1283,N_19051,N_19879);
and UO_1284 (O_1284,N_19212,N_19138);
and UO_1285 (O_1285,N_19962,N_19843);
nor UO_1286 (O_1286,N_19990,N_19162);
nor UO_1287 (O_1287,N_19423,N_19503);
xnor UO_1288 (O_1288,N_19917,N_19151);
xor UO_1289 (O_1289,N_19705,N_19913);
or UO_1290 (O_1290,N_19869,N_19207);
or UO_1291 (O_1291,N_19360,N_19026);
xor UO_1292 (O_1292,N_19132,N_19956);
xor UO_1293 (O_1293,N_19962,N_19123);
nand UO_1294 (O_1294,N_19290,N_19400);
and UO_1295 (O_1295,N_19837,N_19111);
or UO_1296 (O_1296,N_19236,N_19314);
xnor UO_1297 (O_1297,N_19101,N_19715);
or UO_1298 (O_1298,N_19934,N_19076);
nor UO_1299 (O_1299,N_19760,N_19258);
and UO_1300 (O_1300,N_19344,N_19120);
nor UO_1301 (O_1301,N_19132,N_19906);
nand UO_1302 (O_1302,N_19625,N_19822);
or UO_1303 (O_1303,N_19385,N_19460);
nor UO_1304 (O_1304,N_19537,N_19505);
xnor UO_1305 (O_1305,N_19943,N_19182);
and UO_1306 (O_1306,N_19543,N_19506);
xnor UO_1307 (O_1307,N_19848,N_19065);
or UO_1308 (O_1308,N_19730,N_19228);
xor UO_1309 (O_1309,N_19261,N_19530);
nor UO_1310 (O_1310,N_19163,N_19130);
nor UO_1311 (O_1311,N_19822,N_19634);
xor UO_1312 (O_1312,N_19148,N_19184);
or UO_1313 (O_1313,N_19180,N_19009);
or UO_1314 (O_1314,N_19479,N_19135);
nor UO_1315 (O_1315,N_19521,N_19176);
nand UO_1316 (O_1316,N_19792,N_19231);
and UO_1317 (O_1317,N_19738,N_19356);
xor UO_1318 (O_1318,N_19076,N_19529);
xor UO_1319 (O_1319,N_19855,N_19282);
or UO_1320 (O_1320,N_19278,N_19062);
nand UO_1321 (O_1321,N_19121,N_19778);
and UO_1322 (O_1322,N_19411,N_19789);
or UO_1323 (O_1323,N_19119,N_19432);
or UO_1324 (O_1324,N_19968,N_19326);
or UO_1325 (O_1325,N_19268,N_19331);
or UO_1326 (O_1326,N_19207,N_19039);
or UO_1327 (O_1327,N_19516,N_19903);
xnor UO_1328 (O_1328,N_19137,N_19225);
nand UO_1329 (O_1329,N_19344,N_19762);
nor UO_1330 (O_1330,N_19808,N_19337);
or UO_1331 (O_1331,N_19363,N_19254);
nand UO_1332 (O_1332,N_19630,N_19856);
or UO_1333 (O_1333,N_19882,N_19362);
xnor UO_1334 (O_1334,N_19137,N_19300);
nand UO_1335 (O_1335,N_19513,N_19903);
nor UO_1336 (O_1336,N_19535,N_19271);
xnor UO_1337 (O_1337,N_19898,N_19442);
and UO_1338 (O_1338,N_19322,N_19862);
and UO_1339 (O_1339,N_19953,N_19927);
nand UO_1340 (O_1340,N_19319,N_19675);
and UO_1341 (O_1341,N_19677,N_19618);
and UO_1342 (O_1342,N_19138,N_19520);
or UO_1343 (O_1343,N_19136,N_19294);
or UO_1344 (O_1344,N_19236,N_19809);
and UO_1345 (O_1345,N_19898,N_19652);
nand UO_1346 (O_1346,N_19591,N_19628);
xnor UO_1347 (O_1347,N_19617,N_19412);
and UO_1348 (O_1348,N_19831,N_19723);
nor UO_1349 (O_1349,N_19939,N_19439);
xnor UO_1350 (O_1350,N_19405,N_19561);
xnor UO_1351 (O_1351,N_19203,N_19809);
nor UO_1352 (O_1352,N_19534,N_19072);
nor UO_1353 (O_1353,N_19113,N_19639);
or UO_1354 (O_1354,N_19472,N_19832);
and UO_1355 (O_1355,N_19484,N_19284);
xnor UO_1356 (O_1356,N_19837,N_19826);
or UO_1357 (O_1357,N_19541,N_19718);
nor UO_1358 (O_1358,N_19164,N_19953);
and UO_1359 (O_1359,N_19081,N_19098);
nor UO_1360 (O_1360,N_19479,N_19127);
nand UO_1361 (O_1361,N_19278,N_19436);
and UO_1362 (O_1362,N_19514,N_19553);
or UO_1363 (O_1363,N_19984,N_19496);
nand UO_1364 (O_1364,N_19282,N_19465);
nor UO_1365 (O_1365,N_19697,N_19583);
xnor UO_1366 (O_1366,N_19580,N_19766);
or UO_1367 (O_1367,N_19223,N_19539);
or UO_1368 (O_1368,N_19786,N_19153);
and UO_1369 (O_1369,N_19196,N_19978);
xor UO_1370 (O_1370,N_19034,N_19831);
nand UO_1371 (O_1371,N_19916,N_19497);
xor UO_1372 (O_1372,N_19515,N_19996);
and UO_1373 (O_1373,N_19212,N_19670);
nand UO_1374 (O_1374,N_19183,N_19646);
or UO_1375 (O_1375,N_19129,N_19870);
nor UO_1376 (O_1376,N_19279,N_19329);
nand UO_1377 (O_1377,N_19952,N_19504);
nor UO_1378 (O_1378,N_19079,N_19085);
xor UO_1379 (O_1379,N_19237,N_19427);
and UO_1380 (O_1380,N_19665,N_19409);
or UO_1381 (O_1381,N_19322,N_19252);
or UO_1382 (O_1382,N_19712,N_19947);
nand UO_1383 (O_1383,N_19917,N_19056);
or UO_1384 (O_1384,N_19528,N_19054);
and UO_1385 (O_1385,N_19907,N_19339);
or UO_1386 (O_1386,N_19568,N_19291);
xor UO_1387 (O_1387,N_19953,N_19888);
xor UO_1388 (O_1388,N_19404,N_19581);
xor UO_1389 (O_1389,N_19840,N_19932);
nor UO_1390 (O_1390,N_19539,N_19235);
nand UO_1391 (O_1391,N_19687,N_19607);
nor UO_1392 (O_1392,N_19671,N_19424);
nor UO_1393 (O_1393,N_19711,N_19545);
nor UO_1394 (O_1394,N_19636,N_19671);
or UO_1395 (O_1395,N_19855,N_19887);
xnor UO_1396 (O_1396,N_19570,N_19001);
xor UO_1397 (O_1397,N_19209,N_19192);
or UO_1398 (O_1398,N_19904,N_19913);
and UO_1399 (O_1399,N_19299,N_19686);
nand UO_1400 (O_1400,N_19842,N_19460);
or UO_1401 (O_1401,N_19683,N_19556);
and UO_1402 (O_1402,N_19739,N_19369);
nand UO_1403 (O_1403,N_19048,N_19933);
nand UO_1404 (O_1404,N_19057,N_19529);
and UO_1405 (O_1405,N_19986,N_19119);
and UO_1406 (O_1406,N_19223,N_19972);
xnor UO_1407 (O_1407,N_19197,N_19792);
or UO_1408 (O_1408,N_19126,N_19589);
xnor UO_1409 (O_1409,N_19234,N_19036);
nor UO_1410 (O_1410,N_19719,N_19553);
or UO_1411 (O_1411,N_19352,N_19973);
and UO_1412 (O_1412,N_19733,N_19393);
nor UO_1413 (O_1413,N_19608,N_19523);
xnor UO_1414 (O_1414,N_19849,N_19688);
or UO_1415 (O_1415,N_19898,N_19887);
nor UO_1416 (O_1416,N_19411,N_19481);
nand UO_1417 (O_1417,N_19260,N_19803);
and UO_1418 (O_1418,N_19953,N_19056);
xnor UO_1419 (O_1419,N_19516,N_19910);
nor UO_1420 (O_1420,N_19446,N_19171);
and UO_1421 (O_1421,N_19384,N_19150);
and UO_1422 (O_1422,N_19869,N_19055);
nor UO_1423 (O_1423,N_19889,N_19210);
xnor UO_1424 (O_1424,N_19703,N_19456);
xnor UO_1425 (O_1425,N_19317,N_19729);
nor UO_1426 (O_1426,N_19137,N_19856);
xor UO_1427 (O_1427,N_19516,N_19384);
and UO_1428 (O_1428,N_19687,N_19811);
xnor UO_1429 (O_1429,N_19113,N_19526);
xor UO_1430 (O_1430,N_19315,N_19881);
and UO_1431 (O_1431,N_19338,N_19335);
xnor UO_1432 (O_1432,N_19308,N_19617);
xor UO_1433 (O_1433,N_19564,N_19749);
xnor UO_1434 (O_1434,N_19149,N_19393);
and UO_1435 (O_1435,N_19365,N_19834);
xnor UO_1436 (O_1436,N_19688,N_19228);
and UO_1437 (O_1437,N_19848,N_19695);
xnor UO_1438 (O_1438,N_19300,N_19345);
nand UO_1439 (O_1439,N_19646,N_19639);
nand UO_1440 (O_1440,N_19659,N_19342);
and UO_1441 (O_1441,N_19176,N_19851);
xnor UO_1442 (O_1442,N_19357,N_19640);
or UO_1443 (O_1443,N_19610,N_19836);
nand UO_1444 (O_1444,N_19326,N_19145);
and UO_1445 (O_1445,N_19842,N_19791);
and UO_1446 (O_1446,N_19201,N_19965);
nand UO_1447 (O_1447,N_19525,N_19731);
and UO_1448 (O_1448,N_19904,N_19678);
and UO_1449 (O_1449,N_19218,N_19917);
nor UO_1450 (O_1450,N_19582,N_19797);
nand UO_1451 (O_1451,N_19739,N_19879);
nor UO_1452 (O_1452,N_19614,N_19145);
or UO_1453 (O_1453,N_19345,N_19537);
nand UO_1454 (O_1454,N_19749,N_19191);
nand UO_1455 (O_1455,N_19752,N_19674);
xnor UO_1456 (O_1456,N_19100,N_19692);
nand UO_1457 (O_1457,N_19662,N_19214);
xor UO_1458 (O_1458,N_19402,N_19031);
nor UO_1459 (O_1459,N_19163,N_19357);
and UO_1460 (O_1460,N_19712,N_19604);
nor UO_1461 (O_1461,N_19396,N_19122);
nand UO_1462 (O_1462,N_19097,N_19106);
nand UO_1463 (O_1463,N_19863,N_19899);
and UO_1464 (O_1464,N_19225,N_19834);
and UO_1465 (O_1465,N_19133,N_19726);
xnor UO_1466 (O_1466,N_19671,N_19685);
xnor UO_1467 (O_1467,N_19389,N_19608);
nor UO_1468 (O_1468,N_19938,N_19726);
xor UO_1469 (O_1469,N_19903,N_19443);
nor UO_1470 (O_1470,N_19998,N_19920);
or UO_1471 (O_1471,N_19896,N_19731);
and UO_1472 (O_1472,N_19808,N_19343);
and UO_1473 (O_1473,N_19070,N_19597);
or UO_1474 (O_1474,N_19882,N_19686);
nand UO_1475 (O_1475,N_19066,N_19828);
nand UO_1476 (O_1476,N_19865,N_19576);
xor UO_1477 (O_1477,N_19683,N_19128);
and UO_1478 (O_1478,N_19125,N_19189);
nor UO_1479 (O_1479,N_19896,N_19960);
nor UO_1480 (O_1480,N_19862,N_19608);
xor UO_1481 (O_1481,N_19443,N_19518);
nor UO_1482 (O_1482,N_19610,N_19250);
or UO_1483 (O_1483,N_19318,N_19852);
nor UO_1484 (O_1484,N_19519,N_19946);
nor UO_1485 (O_1485,N_19634,N_19207);
nand UO_1486 (O_1486,N_19526,N_19366);
nor UO_1487 (O_1487,N_19500,N_19797);
xnor UO_1488 (O_1488,N_19178,N_19475);
nand UO_1489 (O_1489,N_19227,N_19871);
nand UO_1490 (O_1490,N_19420,N_19365);
and UO_1491 (O_1491,N_19672,N_19380);
xor UO_1492 (O_1492,N_19747,N_19317);
nor UO_1493 (O_1493,N_19093,N_19997);
nor UO_1494 (O_1494,N_19361,N_19419);
xnor UO_1495 (O_1495,N_19212,N_19990);
xnor UO_1496 (O_1496,N_19257,N_19807);
or UO_1497 (O_1497,N_19054,N_19467);
and UO_1498 (O_1498,N_19019,N_19356);
xnor UO_1499 (O_1499,N_19236,N_19170);
nand UO_1500 (O_1500,N_19620,N_19481);
nand UO_1501 (O_1501,N_19301,N_19150);
nor UO_1502 (O_1502,N_19584,N_19687);
xnor UO_1503 (O_1503,N_19639,N_19688);
and UO_1504 (O_1504,N_19228,N_19287);
nand UO_1505 (O_1505,N_19885,N_19163);
nor UO_1506 (O_1506,N_19318,N_19756);
nand UO_1507 (O_1507,N_19231,N_19577);
nand UO_1508 (O_1508,N_19732,N_19525);
nand UO_1509 (O_1509,N_19922,N_19137);
or UO_1510 (O_1510,N_19924,N_19427);
xor UO_1511 (O_1511,N_19071,N_19713);
and UO_1512 (O_1512,N_19942,N_19968);
or UO_1513 (O_1513,N_19965,N_19254);
nor UO_1514 (O_1514,N_19959,N_19711);
or UO_1515 (O_1515,N_19782,N_19082);
and UO_1516 (O_1516,N_19386,N_19187);
nand UO_1517 (O_1517,N_19716,N_19308);
nor UO_1518 (O_1518,N_19695,N_19717);
nor UO_1519 (O_1519,N_19064,N_19882);
xor UO_1520 (O_1520,N_19132,N_19848);
nor UO_1521 (O_1521,N_19526,N_19497);
nand UO_1522 (O_1522,N_19051,N_19630);
or UO_1523 (O_1523,N_19966,N_19014);
and UO_1524 (O_1524,N_19553,N_19794);
nand UO_1525 (O_1525,N_19638,N_19523);
xnor UO_1526 (O_1526,N_19799,N_19039);
or UO_1527 (O_1527,N_19879,N_19832);
and UO_1528 (O_1528,N_19822,N_19739);
nand UO_1529 (O_1529,N_19064,N_19296);
nor UO_1530 (O_1530,N_19983,N_19602);
or UO_1531 (O_1531,N_19310,N_19943);
or UO_1532 (O_1532,N_19134,N_19194);
nand UO_1533 (O_1533,N_19306,N_19514);
nand UO_1534 (O_1534,N_19376,N_19184);
nor UO_1535 (O_1535,N_19817,N_19015);
nand UO_1536 (O_1536,N_19560,N_19368);
or UO_1537 (O_1537,N_19068,N_19210);
nor UO_1538 (O_1538,N_19062,N_19177);
nand UO_1539 (O_1539,N_19946,N_19082);
and UO_1540 (O_1540,N_19633,N_19813);
nand UO_1541 (O_1541,N_19002,N_19540);
or UO_1542 (O_1542,N_19300,N_19152);
nor UO_1543 (O_1543,N_19680,N_19313);
or UO_1544 (O_1544,N_19626,N_19505);
nor UO_1545 (O_1545,N_19120,N_19944);
nand UO_1546 (O_1546,N_19526,N_19775);
and UO_1547 (O_1547,N_19457,N_19914);
or UO_1548 (O_1548,N_19142,N_19137);
nor UO_1549 (O_1549,N_19060,N_19429);
nand UO_1550 (O_1550,N_19946,N_19124);
or UO_1551 (O_1551,N_19248,N_19201);
nand UO_1552 (O_1552,N_19954,N_19620);
xnor UO_1553 (O_1553,N_19860,N_19056);
nand UO_1554 (O_1554,N_19226,N_19503);
nand UO_1555 (O_1555,N_19093,N_19128);
or UO_1556 (O_1556,N_19330,N_19836);
xor UO_1557 (O_1557,N_19304,N_19478);
nor UO_1558 (O_1558,N_19743,N_19375);
nand UO_1559 (O_1559,N_19537,N_19573);
nand UO_1560 (O_1560,N_19798,N_19845);
nand UO_1561 (O_1561,N_19424,N_19850);
nand UO_1562 (O_1562,N_19111,N_19330);
or UO_1563 (O_1563,N_19786,N_19001);
nor UO_1564 (O_1564,N_19369,N_19439);
xor UO_1565 (O_1565,N_19251,N_19308);
nand UO_1566 (O_1566,N_19899,N_19832);
or UO_1567 (O_1567,N_19841,N_19031);
nand UO_1568 (O_1568,N_19888,N_19938);
and UO_1569 (O_1569,N_19818,N_19341);
nand UO_1570 (O_1570,N_19050,N_19093);
and UO_1571 (O_1571,N_19569,N_19539);
nand UO_1572 (O_1572,N_19768,N_19464);
nor UO_1573 (O_1573,N_19297,N_19011);
and UO_1574 (O_1574,N_19014,N_19376);
and UO_1575 (O_1575,N_19695,N_19759);
nor UO_1576 (O_1576,N_19796,N_19626);
nand UO_1577 (O_1577,N_19394,N_19592);
and UO_1578 (O_1578,N_19038,N_19735);
or UO_1579 (O_1579,N_19501,N_19883);
or UO_1580 (O_1580,N_19268,N_19582);
or UO_1581 (O_1581,N_19018,N_19454);
nand UO_1582 (O_1582,N_19264,N_19574);
nor UO_1583 (O_1583,N_19616,N_19590);
nand UO_1584 (O_1584,N_19403,N_19881);
nand UO_1585 (O_1585,N_19132,N_19596);
or UO_1586 (O_1586,N_19891,N_19315);
and UO_1587 (O_1587,N_19021,N_19963);
xnor UO_1588 (O_1588,N_19249,N_19814);
or UO_1589 (O_1589,N_19849,N_19047);
nand UO_1590 (O_1590,N_19447,N_19045);
and UO_1591 (O_1591,N_19507,N_19013);
xnor UO_1592 (O_1592,N_19904,N_19820);
and UO_1593 (O_1593,N_19730,N_19128);
xor UO_1594 (O_1594,N_19864,N_19065);
nand UO_1595 (O_1595,N_19884,N_19546);
nor UO_1596 (O_1596,N_19155,N_19587);
and UO_1597 (O_1597,N_19727,N_19587);
nand UO_1598 (O_1598,N_19269,N_19973);
and UO_1599 (O_1599,N_19012,N_19006);
nor UO_1600 (O_1600,N_19447,N_19638);
and UO_1601 (O_1601,N_19818,N_19568);
and UO_1602 (O_1602,N_19960,N_19342);
xor UO_1603 (O_1603,N_19857,N_19627);
or UO_1604 (O_1604,N_19151,N_19222);
and UO_1605 (O_1605,N_19077,N_19755);
or UO_1606 (O_1606,N_19835,N_19942);
nor UO_1607 (O_1607,N_19966,N_19176);
nor UO_1608 (O_1608,N_19772,N_19559);
and UO_1609 (O_1609,N_19115,N_19050);
nor UO_1610 (O_1610,N_19843,N_19288);
nand UO_1611 (O_1611,N_19853,N_19832);
and UO_1612 (O_1612,N_19277,N_19730);
and UO_1613 (O_1613,N_19281,N_19166);
nor UO_1614 (O_1614,N_19082,N_19336);
nor UO_1615 (O_1615,N_19637,N_19569);
and UO_1616 (O_1616,N_19549,N_19300);
nand UO_1617 (O_1617,N_19230,N_19228);
xor UO_1618 (O_1618,N_19249,N_19345);
xor UO_1619 (O_1619,N_19691,N_19200);
and UO_1620 (O_1620,N_19447,N_19562);
xnor UO_1621 (O_1621,N_19663,N_19460);
nor UO_1622 (O_1622,N_19385,N_19787);
or UO_1623 (O_1623,N_19364,N_19133);
or UO_1624 (O_1624,N_19964,N_19452);
or UO_1625 (O_1625,N_19846,N_19111);
nand UO_1626 (O_1626,N_19957,N_19640);
xor UO_1627 (O_1627,N_19764,N_19143);
xor UO_1628 (O_1628,N_19686,N_19324);
and UO_1629 (O_1629,N_19975,N_19790);
and UO_1630 (O_1630,N_19524,N_19662);
nand UO_1631 (O_1631,N_19016,N_19839);
and UO_1632 (O_1632,N_19086,N_19615);
xnor UO_1633 (O_1633,N_19662,N_19073);
nand UO_1634 (O_1634,N_19411,N_19868);
nor UO_1635 (O_1635,N_19432,N_19197);
nor UO_1636 (O_1636,N_19643,N_19201);
nor UO_1637 (O_1637,N_19691,N_19689);
nand UO_1638 (O_1638,N_19151,N_19896);
and UO_1639 (O_1639,N_19421,N_19365);
nor UO_1640 (O_1640,N_19185,N_19519);
xnor UO_1641 (O_1641,N_19036,N_19323);
nor UO_1642 (O_1642,N_19996,N_19685);
nand UO_1643 (O_1643,N_19618,N_19416);
nor UO_1644 (O_1644,N_19655,N_19535);
nand UO_1645 (O_1645,N_19207,N_19740);
nand UO_1646 (O_1646,N_19115,N_19093);
nand UO_1647 (O_1647,N_19889,N_19402);
nor UO_1648 (O_1648,N_19466,N_19150);
nand UO_1649 (O_1649,N_19596,N_19703);
or UO_1650 (O_1650,N_19075,N_19520);
xnor UO_1651 (O_1651,N_19653,N_19621);
xnor UO_1652 (O_1652,N_19948,N_19882);
xor UO_1653 (O_1653,N_19628,N_19875);
nor UO_1654 (O_1654,N_19501,N_19531);
xor UO_1655 (O_1655,N_19423,N_19164);
nand UO_1656 (O_1656,N_19435,N_19740);
xor UO_1657 (O_1657,N_19566,N_19660);
xnor UO_1658 (O_1658,N_19399,N_19833);
or UO_1659 (O_1659,N_19560,N_19815);
nor UO_1660 (O_1660,N_19640,N_19847);
nor UO_1661 (O_1661,N_19584,N_19702);
xnor UO_1662 (O_1662,N_19588,N_19999);
nand UO_1663 (O_1663,N_19476,N_19280);
xnor UO_1664 (O_1664,N_19803,N_19014);
and UO_1665 (O_1665,N_19104,N_19358);
nor UO_1666 (O_1666,N_19366,N_19892);
nor UO_1667 (O_1667,N_19966,N_19811);
and UO_1668 (O_1668,N_19363,N_19634);
or UO_1669 (O_1669,N_19209,N_19076);
nor UO_1670 (O_1670,N_19871,N_19329);
xor UO_1671 (O_1671,N_19911,N_19670);
nor UO_1672 (O_1672,N_19633,N_19739);
nor UO_1673 (O_1673,N_19169,N_19319);
and UO_1674 (O_1674,N_19913,N_19304);
nor UO_1675 (O_1675,N_19743,N_19358);
or UO_1676 (O_1676,N_19278,N_19610);
nand UO_1677 (O_1677,N_19364,N_19377);
and UO_1678 (O_1678,N_19402,N_19164);
nand UO_1679 (O_1679,N_19348,N_19266);
and UO_1680 (O_1680,N_19436,N_19564);
and UO_1681 (O_1681,N_19179,N_19093);
and UO_1682 (O_1682,N_19790,N_19129);
nand UO_1683 (O_1683,N_19589,N_19920);
nor UO_1684 (O_1684,N_19758,N_19680);
xor UO_1685 (O_1685,N_19026,N_19925);
xor UO_1686 (O_1686,N_19105,N_19709);
or UO_1687 (O_1687,N_19011,N_19797);
or UO_1688 (O_1688,N_19014,N_19128);
nand UO_1689 (O_1689,N_19626,N_19982);
nor UO_1690 (O_1690,N_19571,N_19097);
nand UO_1691 (O_1691,N_19569,N_19697);
nor UO_1692 (O_1692,N_19678,N_19108);
and UO_1693 (O_1693,N_19246,N_19060);
or UO_1694 (O_1694,N_19389,N_19270);
and UO_1695 (O_1695,N_19639,N_19498);
nand UO_1696 (O_1696,N_19592,N_19241);
and UO_1697 (O_1697,N_19289,N_19342);
xnor UO_1698 (O_1698,N_19747,N_19620);
or UO_1699 (O_1699,N_19394,N_19619);
or UO_1700 (O_1700,N_19970,N_19790);
nor UO_1701 (O_1701,N_19362,N_19678);
nand UO_1702 (O_1702,N_19200,N_19249);
or UO_1703 (O_1703,N_19941,N_19680);
nor UO_1704 (O_1704,N_19594,N_19302);
xor UO_1705 (O_1705,N_19516,N_19686);
nand UO_1706 (O_1706,N_19599,N_19023);
nor UO_1707 (O_1707,N_19694,N_19966);
or UO_1708 (O_1708,N_19019,N_19347);
xnor UO_1709 (O_1709,N_19268,N_19974);
nand UO_1710 (O_1710,N_19007,N_19711);
and UO_1711 (O_1711,N_19293,N_19386);
and UO_1712 (O_1712,N_19798,N_19525);
or UO_1713 (O_1713,N_19739,N_19350);
and UO_1714 (O_1714,N_19748,N_19452);
nor UO_1715 (O_1715,N_19530,N_19254);
nand UO_1716 (O_1716,N_19709,N_19442);
and UO_1717 (O_1717,N_19000,N_19620);
xnor UO_1718 (O_1718,N_19653,N_19724);
nor UO_1719 (O_1719,N_19928,N_19101);
or UO_1720 (O_1720,N_19340,N_19369);
and UO_1721 (O_1721,N_19242,N_19595);
nand UO_1722 (O_1722,N_19823,N_19756);
nand UO_1723 (O_1723,N_19103,N_19041);
or UO_1724 (O_1724,N_19591,N_19235);
or UO_1725 (O_1725,N_19021,N_19600);
nand UO_1726 (O_1726,N_19206,N_19985);
nor UO_1727 (O_1727,N_19453,N_19722);
xnor UO_1728 (O_1728,N_19681,N_19004);
nor UO_1729 (O_1729,N_19762,N_19293);
or UO_1730 (O_1730,N_19569,N_19722);
or UO_1731 (O_1731,N_19260,N_19303);
xor UO_1732 (O_1732,N_19351,N_19216);
and UO_1733 (O_1733,N_19526,N_19834);
nand UO_1734 (O_1734,N_19116,N_19880);
and UO_1735 (O_1735,N_19814,N_19908);
nor UO_1736 (O_1736,N_19852,N_19013);
and UO_1737 (O_1737,N_19043,N_19547);
xnor UO_1738 (O_1738,N_19668,N_19948);
and UO_1739 (O_1739,N_19359,N_19924);
or UO_1740 (O_1740,N_19863,N_19054);
nor UO_1741 (O_1741,N_19046,N_19175);
nand UO_1742 (O_1742,N_19824,N_19753);
or UO_1743 (O_1743,N_19901,N_19051);
xor UO_1744 (O_1744,N_19791,N_19733);
or UO_1745 (O_1745,N_19572,N_19858);
and UO_1746 (O_1746,N_19073,N_19210);
and UO_1747 (O_1747,N_19618,N_19966);
nor UO_1748 (O_1748,N_19963,N_19408);
or UO_1749 (O_1749,N_19980,N_19430);
nor UO_1750 (O_1750,N_19290,N_19655);
or UO_1751 (O_1751,N_19638,N_19474);
and UO_1752 (O_1752,N_19067,N_19994);
and UO_1753 (O_1753,N_19953,N_19949);
nand UO_1754 (O_1754,N_19982,N_19999);
nor UO_1755 (O_1755,N_19531,N_19929);
xor UO_1756 (O_1756,N_19435,N_19700);
xor UO_1757 (O_1757,N_19967,N_19539);
xnor UO_1758 (O_1758,N_19910,N_19861);
nand UO_1759 (O_1759,N_19724,N_19558);
and UO_1760 (O_1760,N_19751,N_19675);
nor UO_1761 (O_1761,N_19577,N_19961);
xor UO_1762 (O_1762,N_19546,N_19651);
and UO_1763 (O_1763,N_19963,N_19707);
nor UO_1764 (O_1764,N_19670,N_19607);
xnor UO_1765 (O_1765,N_19457,N_19088);
or UO_1766 (O_1766,N_19385,N_19487);
and UO_1767 (O_1767,N_19504,N_19923);
nor UO_1768 (O_1768,N_19935,N_19680);
xnor UO_1769 (O_1769,N_19099,N_19063);
nand UO_1770 (O_1770,N_19294,N_19899);
nor UO_1771 (O_1771,N_19973,N_19112);
xor UO_1772 (O_1772,N_19248,N_19746);
xor UO_1773 (O_1773,N_19667,N_19174);
nand UO_1774 (O_1774,N_19753,N_19175);
or UO_1775 (O_1775,N_19672,N_19595);
nand UO_1776 (O_1776,N_19447,N_19320);
nor UO_1777 (O_1777,N_19109,N_19797);
or UO_1778 (O_1778,N_19118,N_19641);
xnor UO_1779 (O_1779,N_19418,N_19642);
or UO_1780 (O_1780,N_19161,N_19893);
and UO_1781 (O_1781,N_19570,N_19713);
or UO_1782 (O_1782,N_19048,N_19094);
or UO_1783 (O_1783,N_19175,N_19719);
xor UO_1784 (O_1784,N_19919,N_19329);
xnor UO_1785 (O_1785,N_19802,N_19848);
nor UO_1786 (O_1786,N_19760,N_19525);
xor UO_1787 (O_1787,N_19913,N_19813);
and UO_1788 (O_1788,N_19383,N_19328);
or UO_1789 (O_1789,N_19133,N_19247);
and UO_1790 (O_1790,N_19548,N_19401);
and UO_1791 (O_1791,N_19330,N_19994);
nand UO_1792 (O_1792,N_19537,N_19199);
and UO_1793 (O_1793,N_19678,N_19109);
nor UO_1794 (O_1794,N_19831,N_19076);
xor UO_1795 (O_1795,N_19831,N_19063);
and UO_1796 (O_1796,N_19779,N_19682);
and UO_1797 (O_1797,N_19217,N_19804);
nor UO_1798 (O_1798,N_19358,N_19317);
or UO_1799 (O_1799,N_19894,N_19900);
nor UO_1800 (O_1800,N_19186,N_19004);
nand UO_1801 (O_1801,N_19806,N_19579);
or UO_1802 (O_1802,N_19325,N_19457);
nor UO_1803 (O_1803,N_19330,N_19433);
nor UO_1804 (O_1804,N_19867,N_19716);
and UO_1805 (O_1805,N_19226,N_19702);
and UO_1806 (O_1806,N_19347,N_19523);
xnor UO_1807 (O_1807,N_19203,N_19812);
or UO_1808 (O_1808,N_19256,N_19542);
nand UO_1809 (O_1809,N_19961,N_19552);
nor UO_1810 (O_1810,N_19516,N_19436);
nand UO_1811 (O_1811,N_19365,N_19564);
and UO_1812 (O_1812,N_19110,N_19447);
or UO_1813 (O_1813,N_19693,N_19385);
or UO_1814 (O_1814,N_19549,N_19204);
nand UO_1815 (O_1815,N_19059,N_19549);
or UO_1816 (O_1816,N_19183,N_19712);
nor UO_1817 (O_1817,N_19246,N_19682);
nor UO_1818 (O_1818,N_19735,N_19800);
or UO_1819 (O_1819,N_19469,N_19459);
nor UO_1820 (O_1820,N_19761,N_19204);
and UO_1821 (O_1821,N_19040,N_19883);
nor UO_1822 (O_1822,N_19901,N_19220);
nand UO_1823 (O_1823,N_19937,N_19157);
or UO_1824 (O_1824,N_19994,N_19946);
or UO_1825 (O_1825,N_19183,N_19564);
nand UO_1826 (O_1826,N_19863,N_19348);
or UO_1827 (O_1827,N_19318,N_19640);
xor UO_1828 (O_1828,N_19115,N_19136);
xnor UO_1829 (O_1829,N_19056,N_19594);
and UO_1830 (O_1830,N_19885,N_19231);
and UO_1831 (O_1831,N_19778,N_19214);
or UO_1832 (O_1832,N_19228,N_19573);
and UO_1833 (O_1833,N_19855,N_19758);
nor UO_1834 (O_1834,N_19532,N_19372);
and UO_1835 (O_1835,N_19100,N_19205);
nor UO_1836 (O_1836,N_19479,N_19476);
or UO_1837 (O_1837,N_19387,N_19938);
nor UO_1838 (O_1838,N_19651,N_19661);
nor UO_1839 (O_1839,N_19159,N_19781);
xor UO_1840 (O_1840,N_19795,N_19474);
nand UO_1841 (O_1841,N_19156,N_19419);
and UO_1842 (O_1842,N_19872,N_19037);
or UO_1843 (O_1843,N_19659,N_19242);
or UO_1844 (O_1844,N_19398,N_19095);
nand UO_1845 (O_1845,N_19018,N_19426);
and UO_1846 (O_1846,N_19772,N_19088);
and UO_1847 (O_1847,N_19260,N_19063);
nand UO_1848 (O_1848,N_19237,N_19684);
nand UO_1849 (O_1849,N_19078,N_19070);
and UO_1850 (O_1850,N_19286,N_19513);
or UO_1851 (O_1851,N_19745,N_19023);
or UO_1852 (O_1852,N_19132,N_19476);
or UO_1853 (O_1853,N_19109,N_19591);
nor UO_1854 (O_1854,N_19738,N_19281);
nand UO_1855 (O_1855,N_19700,N_19297);
or UO_1856 (O_1856,N_19329,N_19162);
nand UO_1857 (O_1857,N_19509,N_19663);
nor UO_1858 (O_1858,N_19634,N_19732);
nor UO_1859 (O_1859,N_19374,N_19829);
xnor UO_1860 (O_1860,N_19419,N_19802);
or UO_1861 (O_1861,N_19492,N_19282);
nor UO_1862 (O_1862,N_19245,N_19884);
xor UO_1863 (O_1863,N_19436,N_19096);
and UO_1864 (O_1864,N_19576,N_19875);
nand UO_1865 (O_1865,N_19223,N_19639);
nor UO_1866 (O_1866,N_19765,N_19145);
nand UO_1867 (O_1867,N_19187,N_19470);
and UO_1868 (O_1868,N_19228,N_19510);
and UO_1869 (O_1869,N_19384,N_19643);
or UO_1870 (O_1870,N_19579,N_19722);
xor UO_1871 (O_1871,N_19816,N_19748);
nand UO_1872 (O_1872,N_19516,N_19087);
and UO_1873 (O_1873,N_19244,N_19188);
xnor UO_1874 (O_1874,N_19562,N_19542);
xnor UO_1875 (O_1875,N_19606,N_19355);
xor UO_1876 (O_1876,N_19264,N_19008);
and UO_1877 (O_1877,N_19683,N_19141);
and UO_1878 (O_1878,N_19279,N_19697);
nand UO_1879 (O_1879,N_19688,N_19609);
xor UO_1880 (O_1880,N_19759,N_19400);
nand UO_1881 (O_1881,N_19024,N_19350);
nand UO_1882 (O_1882,N_19778,N_19912);
nand UO_1883 (O_1883,N_19605,N_19851);
or UO_1884 (O_1884,N_19411,N_19224);
nor UO_1885 (O_1885,N_19586,N_19365);
or UO_1886 (O_1886,N_19834,N_19178);
xor UO_1887 (O_1887,N_19074,N_19182);
and UO_1888 (O_1888,N_19668,N_19579);
and UO_1889 (O_1889,N_19001,N_19032);
nand UO_1890 (O_1890,N_19065,N_19707);
and UO_1891 (O_1891,N_19212,N_19238);
or UO_1892 (O_1892,N_19620,N_19125);
and UO_1893 (O_1893,N_19045,N_19999);
xnor UO_1894 (O_1894,N_19301,N_19950);
nor UO_1895 (O_1895,N_19295,N_19843);
nor UO_1896 (O_1896,N_19055,N_19888);
nand UO_1897 (O_1897,N_19383,N_19708);
and UO_1898 (O_1898,N_19983,N_19288);
or UO_1899 (O_1899,N_19226,N_19449);
nand UO_1900 (O_1900,N_19393,N_19949);
xor UO_1901 (O_1901,N_19917,N_19087);
nand UO_1902 (O_1902,N_19052,N_19300);
and UO_1903 (O_1903,N_19635,N_19093);
xnor UO_1904 (O_1904,N_19333,N_19715);
xnor UO_1905 (O_1905,N_19461,N_19993);
nor UO_1906 (O_1906,N_19604,N_19529);
nor UO_1907 (O_1907,N_19271,N_19809);
and UO_1908 (O_1908,N_19403,N_19240);
xor UO_1909 (O_1909,N_19471,N_19078);
and UO_1910 (O_1910,N_19152,N_19135);
nand UO_1911 (O_1911,N_19239,N_19508);
or UO_1912 (O_1912,N_19531,N_19534);
nand UO_1913 (O_1913,N_19467,N_19666);
xor UO_1914 (O_1914,N_19287,N_19422);
or UO_1915 (O_1915,N_19980,N_19835);
nor UO_1916 (O_1916,N_19875,N_19511);
nand UO_1917 (O_1917,N_19082,N_19715);
or UO_1918 (O_1918,N_19725,N_19635);
xor UO_1919 (O_1919,N_19334,N_19934);
and UO_1920 (O_1920,N_19614,N_19218);
xnor UO_1921 (O_1921,N_19529,N_19405);
and UO_1922 (O_1922,N_19450,N_19272);
xor UO_1923 (O_1923,N_19649,N_19627);
nor UO_1924 (O_1924,N_19615,N_19985);
nand UO_1925 (O_1925,N_19085,N_19402);
xnor UO_1926 (O_1926,N_19867,N_19161);
or UO_1927 (O_1927,N_19679,N_19425);
or UO_1928 (O_1928,N_19419,N_19776);
xor UO_1929 (O_1929,N_19771,N_19168);
nor UO_1930 (O_1930,N_19462,N_19020);
xor UO_1931 (O_1931,N_19264,N_19704);
or UO_1932 (O_1932,N_19517,N_19030);
xor UO_1933 (O_1933,N_19578,N_19036);
or UO_1934 (O_1934,N_19184,N_19880);
nor UO_1935 (O_1935,N_19848,N_19049);
or UO_1936 (O_1936,N_19097,N_19972);
or UO_1937 (O_1937,N_19100,N_19014);
or UO_1938 (O_1938,N_19500,N_19905);
nand UO_1939 (O_1939,N_19324,N_19973);
or UO_1940 (O_1940,N_19929,N_19814);
and UO_1941 (O_1941,N_19621,N_19691);
nand UO_1942 (O_1942,N_19159,N_19261);
or UO_1943 (O_1943,N_19976,N_19821);
and UO_1944 (O_1944,N_19138,N_19178);
xnor UO_1945 (O_1945,N_19273,N_19255);
nand UO_1946 (O_1946,N_19882,N_19757);
xor UO_1947 (O_1947,N_19966,N_19218);
and UO_1948 (O_1948,N_19629,N_19030);
nor UO_1949 (O_1949,N_19432,N_19638);
xor UO_1950 (O_1950,N_19239,N_19118);
nor UO_1951 (O_1951,N_19568,N_19472);
nor UO_1952 (O_1952,N_19474,N_19663);
nand UO_1953 (O_1953,N_19660,N_19738);
or UO_1954 (O_1954,N_19928,N_19896);
nor UO_1955 (O_1955,N_19308,N_19136);
nor UO_1956 (O_1956,N_19558,N_19760);
nor UO_1957 (O_1957,N_19154,N_19376);
nand UO_1958 (O_1958,N_19272,N_19879);
nand UO_1959 (O_1959,N_19465,N_19381);
nand UO_1960 (O_1960,N_19112,N_19956);
and UO_1961 (O_1961,N_19626,N_19145);
and UO_1962 (O_1962,N_19415,N_19892);
nand UO_1963 (O_1963,N_19661,N_19886);
nand UO_1964 (O_1964,N_19511,N_19870);
xor UO_1965 (O_1965,N_19027,N_19848);
xor UO_1966 (O_1966,N_19394,N_19790);
nand UO_1967 (O_1967,N_19316,N_19587);
nand UO_1968 (O_1968,N_19461,N_19910);
nand UO_1969 (O_1969,N_19751,N_19059);
and UO_1970 (O_1970,N_19144,N_19815);
and UO_1971 (O_1971,N_19373,N_19442);
and UO_1972 (O_1972,N_19458,N_19542);
xor UO_1973 (O_1973,N_19735,N_19089);
nand UO_1974 (O_1974,N_19859,N_19479);
or UO_1975 (O_1975,N_19250,N_19643);
and UO_1976 (O_1976,N_19884,N_19886);
nor UO_1977 (O_1977,N_19759,N_19939);
and UO_1978 (O_1978,N_19944,N_19812);
or UO_1979 (O_1979,N_19463,N_19060);
or UO_1980 (O_1980,N_19752,N_19204);
nand UO_1981 (O_1981,N_19733,N_19243);
nor UO_1982 (O_1982,N_19402,N_19876);
and UO_1983 (O_1983,N_19691,N_19033);
or UO_1984 (O_1984,N_19925,N_19099);
nor UO_1985 (O_1985,N_19328,N_19913);
xnor UO_1986 (O_1986,N_19515,N_19462);
nand UO_1987 (O_1987,N_19141,N_19316);
nor UO_1988 (O_1988,N_19466,N_19960);
and UO_1989 (O_1989,N_19655,N_19734);
xor UO_1990 (O_1990,N_19595,N_19966);
nor UO_1991 (O_1991,N_19877,N_19821);
nor UO_1992 (O_1992,N_19073,N_19710);
nand UO_1993 (O_1993,N_19789,N_19055);
and UO_1994 (O_1994,N_19721,N_19279);
and UO_1995 (O_1995,N_19390,N_19356);
nor UO_1996 (O_1996,N_19101,N_19157);
nor UO_1997 (O_1997,N_19893,N_19247);
or UO_1998 (O_1998,N_19153,N_19610);
nand UO_1999 (O_1999,N_19244,N_19439);
xor UO_2000 (O_2000,N_19096,N_19348);
nand UO_2001 (O_2001,N_19340,N_19025);
nand UO_2002 (O_2002,N_19785,N_19560);
nor UO_2003 (O_2003,N_19465,N_19645);
or UO_2004 (O_2004,N_19304,N_19484);
and UO_2005 (O_2005,N_19444,N_19803);
xor UO_2006 (O_2006,N_19022,N_19182);
nor UO_2007 (O_2007,N_19031,N_19256);
nand UO_2008 (O_2008,N_19629,N_19005);
xnor UO_2009 (O_2009,N_19712,N_19602);
xor UO_2010 (O_2010,N_19067,N_19210);
xor UO_2011 (O_2011,N_19867,N_19979);
nand UO_2012 (O_2012,N_19609,N_19776);
nand UO_2013 (O_2013,N_19091,N_19460);
nor UO_2014 (O_2014,N_19341,N_19822);
and UO_2015 (O_2015,N_19327,N_19697);
or UO_2016 (O_2016,N_19263,N_19952);
nor UO_2017 (O_2017,N_19140,N_19739);
and UO_2018 (O_2018,N_19768,N_19580);
and UO_2019 (O_2019,N_19365,N_19521);
nand UO_2020 (O_2020,N_19725,N_19903);
and UO_2021 (O_2021,N_19145,N_19633);
nand UO_2022 (O_2022,N_19208,N_19950);
xor UO_2023 (O_2023,N_19310,N_19997);
and UO_2024 (O_2024,N_19623,N_19935);
nor UO_2025 (O_2025,N_19217,N_19027);
xnor UO_2026 (O_2026,N_19551,N_19435);
xor UO_2027 (O_2027,N_19267,N_19919);
xor UO_2028 (O_2028,N_19022,N_19596);
xnor UO_2029 (O_2029,N_19920,N_19008);
nor UO_2030 (O_2030,N_19797,N_19964);
or UO_2031 (O_2031,N_19117,N_19604);
and UO_2032 (O_2032,N_19946,N_19668);
nand UO_2033 (O_2033,N_19200,N_19658);
and UO_2034 (O_2034,N_19861,N_19639);
or UO_2035 (O_2035,N_19951,N_19870);
nor UO_2036 (O_2036,N_19189,N_19498);
nand UO_2037 (O_2037,N_19060,N_19084);
xor UO_2038 (O_2038,N_19305,N_19370);
nand UO_2039 (O_2039,N_19213,N_19852);
nor UO_2040 (O_2040,N_19380,N_19137);
xnor UO_2041 (O_2041,N_19971,N_19894);
nand UO_2042 (O_2042,N_19230,N_19341);
nor UO_2043 (O_2043,N_19501,N_19543);
nand UO_2044 (O_2044,N_19603,N_19264);
xnor UO_2045 (O_2045,N_19800,N_19240);
xor UO_2046 (O_2046,N_19828,N_19487);
xnor UO_2047 (O_2047,N_19368,N_19638);
xnor UO_2048 (O_2048,N_19019,N_19981);
or UO_2049 (O_2049,N_19426,N_19626);
and UO_2050 (O_2050,N_19691,N_19886);
and UO_2051 (O_2051,N_19214,N_19378);
and UO_2052 (O_2052,N_19024,N_19167);
or UO_2053 (O_2053,N_19606,N_19318);
or UO_2054 (O_2054,N_19916,N_19730);
xor UO_2055 (O_2055,N_19723,N_19693);
xor UO_2056 (O_2056,N_19025,N_19985);
nor UO_2057 (O_2057,N_19688,N_19647);
and UO_2058 (O_2058,N_19026,N_19157);
nand UO_2059 (O_2059,N_19323,N_19110);
nor UO_2060 (O_2060,N_19595,N_19683);
and UO_2061 (O_2061,N_19492,N_19092);
nor UO_2062 (O_2062,N_19537,N_19898);
nand UO_2063 (O_2063,N_19869,N_19844);
xor UO_2064 (O_2064,N_19410,N_19711);
xnor UO_2065 (O_2065,N_19910,N_19162);
xor UO_2066 (O_2066,N_19149,N_19585);
nand UO_2067 (O_2067,N_19399,N_19856);
nor UO_2068 (O_2068,N_19132,N_19644);
or UO_2069 (O_2069,N_19153,N_19195);
or UO_2070 (O_2070,N_19377,N_19402);
nor UO_2071 (O_2071,N_19089,N_19585);
and UO_2072 (O_2072,N_19372,N_19942);
nand UO_2073 (O_2073,N_19933,N_19069);
xor UO_2074 (O_2074,N_19759,N_19651);
and UO_2075 (O_2075,N_19123,N_19183);
nor UO_2076 (O_2076,N_19597,N_19142);
nand UO_2077 (O_2077,N_19981,N_19361);
nor UO_2078 (O_2078,N_19391,N_19107);
or UO_2079 (O_2079,N_19013,N_19220);
xnor UO_2080 (O_2080,N_19297,N_19035);
xnor UO_2081 (O_2081,N_19995,N_19036);
or UO_2082 (O_2082,N_19677,N_19667);
nand UO_2083 (O_2083,N_19261,N_19112);
and UO_2084 (O_2084,N_19685,N_19519);
nor UO_2085 (O_2085,N_19471,N_19809);
and UO_2086 (O_2086,N_19115,N_19529);
xor UO_2087 (O_2087,N_19839,N_19745);
or UO_2088 (O_2088,N_19368,N_19766);
or UO_2089 (O_2089,N_19583,N_19737);
or UO_2090 (O_2090,N_19119,N_19019);
nand UO_2091 (O_2091,N_19888,N_19144);
nor UO_2092 (O_2092,N_19365,N_19182);
or UO_2093 (O_2093,N_19259,N_19498);
nand UO_2094 (O_2094,N_19965,N_19684);
nand UO_2095 (O_2095,N_19583,N_19674);
nand UO_2096 (O_2096,N_19985,N_19971);
nor UO_2097 (O_2097,N_19466,N_19974);
and UO_2098 (O_2098,N_19149,N_19432);
or UO_2099 (O_2099,N_19686,N_19550);
nor UO_2100 (O_2100,N_19535,N_19645);
nand UO_2101 (O_2101,N_19302,N_19446);
xnor UO_2102 (O_2102,N_19353,N_19597);
xnor UO_2103 (O_2103,N_19059,N_19900);
xor UO_2104 (O_2104,N_19914,N_19668);
xnor UO_2105 (O_2105,N_19899,N_19196);
and UO_2106 (O_2106,N_19791,N_19314);
xor UO_2107 (O_2107,N_19443,N_19954);
xnor UO_2108 (O_2108,N_19903,N_19363);
nor UO_2109 (O_2109,N_19536,N_19215);
nor UO_2110 (O_2110,N_19471,N_19323);
nor UO_2111 (O_2111,N_19593,N_19464);
nor UO_2112 (O_2112,N_19272,N_19755);
nor UO_2113 (O_2113,N_19278,N_19433);
and UO_2114 (O_2114,N_19845,N_19825);
xor UO_2115 (O_2115,N_19125,N_19972);
and UO_2116 (O_2116,N_19222,N_19841);
nand UO_2117 (O_2117,N_19618,N_19573);
and UO_2118 (O_2118,N_19335,N_19319);
or UO_2119 (O_2119,N_19549,N_19605);
nand UO_2120 (O_2120,N_19657,N_19343);
xor UO_2121 (O_2121,N_19595,N_19377);
xnor UO_2122 (O_2122,N_19799,N_19441);
nor UO_2123 (O_2123,N_19722,N_19388);
xor UO_2124 (O_2124,N_19809,N_19303);
and UO_2125 (O_2125,N_19076,N_19799);
and UO_2126 (O_2126,N_19808,N_19986);
or UO_2127 (O_2127,N_19356,N_19134);
and UO_2128 (O_2128,N_19651,N_19081);
nor UO_2129 (O_2129,N_19681,N_19081);
and UO_2130 (O_2130,N_19620,N_19494);
and UO_2131 (O_2131,N_19681,N_19228);
and UO_2132 (O_2132,N_19132,N_19668);
nand UO_2133 (O_2133,N_19353,N_19588);
nor UO_2134 (O_2134,N_19002,N_19301);
nor UO_2135 (O_2135,N_19317,N_19091);
xor UO_2136 (O_2136,N_19818,N_19271);
nor UO_2137 (O_2137,N_19501,N_19206);
nor UO_2138 (O_2138,N_19213,N_19311);
or UO_2139 (O_2139,N_19255,N_19116);
or UO_2140 (O_2140,N_19485,N_19280);
nand UO_2141 (O_2141,N_19051,N_19496);
or UO_2142 (O_2142,N_19746,N_19845);
or UO_2143 (O_2143,N_19786,N_19496);
xnor UO_2144 (O_2144,N_19321,N_19696);
and UO_2145 (O_2145,N_19682,N_19375);
and UO_2146 (O_2146,N_19776,N_19509);
xor UO_2147 (O_2147,N_19988,N_19339);
or UO_2148 (O_2148,N_19512,N_19039);
xor UO_2149 (O_2149,N_19798,N_19215);
and UO_2150 (O_2150,N_19883,N_19468);
xnor UO_2151 (O_2151,N_19687,N_19826);
xnor UO_2152 (O_2152,N_19165,N_19338);
and UO_2153 (O_2153,N_19911,N_19223);
and UO_2154 (O_2154,N_19396,N_19629);
or UO_2155 (O_2155,N_19907,N_19558);
nand UO_2156 (O_2156,N_19554,N_19893);
nor UO_2157 (O_2157,N_19178,N_19427);
nor UO_2158 (O_2158,N_19006,N_19802);
or UO_2159 (O_2159,N_19526,N_19841);
nor UO_2160 (O_2160,N_19957,N_19516);
or UO_2161 (O_2161,N_19576,N_19849);
or UO_2162 (O_2162,N_19767,N_19115);
nor UO_2163 (O_2163,N_19743,N_19123);
or UO_2164 (O_2164,N_19573,N_19464);
nor UO_2165 (O_2165,N_19715,N_19220);
or UO_2166 (O_2166,N_19997,N_19278);
nand UO_2167 (O_2167,N_19333,N_19368);
and UO_2168 (O_2168,N_19951,N_19759);
xnor UO_2169 (O_2169,N_19145,N_19196);
nand UO_2170 (O_2170,N_19773,N_19304);
and UO_2171 (O_2171,N_19309,N_19458);
nor UO_2172 (O_2172,N_19014,N_19844);
nand UO_2173 (O_2173,N_19618,N_19952);
nand UO_2174 (O_2174,N_19645,N_19456);
xnor UO_2175 (O_2175,N_19425,N_19409);
xnor UO_2176 (O_2176,N_19553,N_19294);
or UO_2177 (O_2177,N_19735,N_19670);
xnor UO_2178 (O_2178,N_19773,N_19377);
nor UO_2179 (O_2179,N_19750,N_19125);
and UO_2180 (O_2180,N_19762,N_19435);
xnor UO_2181 (O_2181,N_19742,N_19586);
or UO_2182 (O_2182,N_19655,N_19243);
nand UO_2183 (O_2183,N_19959,N_19592);
nand UO_2184 (O_2184,N_19071,N_19198);
nand UO_2185 (O_2185,N_19479,N_19704);
xor UO_2186 (O_2186,N_19975,N_19401);
or UO_2187 (O_2187,N_19837,N_19110);
nor UO_2188 (O_2188,N_19552,N_19251);
xor UO_2189 (O_2189,N_19604,N_19037);
xnor UO_2190 (O_2190,N_19523,N_19029);
or UO_2191 (O_2191,N_19485,N_19790);
nor UO_2192 (O_2192,N_19726,N_19067);
nand UO_2193 (O_2193,N_19151,N_19703);
nor UO_2194 (O_2194,N_19471,N_19838);
nand UO_2195 (O_2195,N_19511,N_19095);
nand UO_2196 (O_2196,N_19580,N_19885);
and UO_2197 (O_2197,N_19040,N_19246);
xor UO_2198 (O_2198,N_19034,N_19811);
and UO_2199 (O_2199,N_19934,N_19451);
xor UO_2200 (O_2200,N_19803,N_19954);
or UO_2201 (O_2201,N_19565,N_19669);
nand UO_2202 (O_2202,N_19367,N_19646);
nand UO_2203 (O_2203,N_19323,N_19621);
nand UO_2204 (O_2204,N_19195,N_19733);
nor UO_2205 (O_2205,N_19456,N_19266);
or UO_2206 (O_2206,N_19622,N_19519);
and UO_2207 (O_2207,N_19438,N_19838);
and UO_2208 (O_2208,N_19063,N_19247);
and UO_2209 (O_2209,N_19398,N_19836);
nor UO_2210 (O_2210,N_19786,N_19667);
and UO_2211 (O_2211,N_19430,N_19446);
and UO_2212 (O_2212,N_19491,N_19735);
xnor UO_2213 (O_2213,N_19159,N_19377);
nor UO_2214 (O_2214,N_19987,N_19358);
or UO_2215 (O_2215,N_19295,N_19301);
xor UO_2216 (O_2216,N_19170,N_19899);
and UO_2217 (O_2217,N_19146,N_19277);
and UO_2218 (O_2218,N_19461,N_19793);
or UO_2219 (O_2219,N_19162,N_19309);
nor UO_2220 (O_2220,N_19452,N_19907);
and UO_2221 (O_2221,N_19858,N_19013);
xnor UO_2222 (O_2222,N_19857,N_19919);
xor UO_2223 (O_2223,N_19274,N_19586);
and UO_2224 (O_2224,N_19158,N_19992);
or UO_2225 (O_2225,N_19785,N_19643);
xor UO_2226 (O_2226,N_19238,N_19413);
xor UO_2227 (O_2227,N_19481,N_19858);
nor UO_2228 (O_2228,N_19793,N_19800);
nor UO_2229 (O_2229,N_19929,N_19453);
xnor UO_2230 (O_2230,N_19843,N_19948);
nand UO_2231 (O_2231,N_19791,N_19983);
nor UO_2232 (O_2232,N_19286,N_19238);
or UO_2233 (O_2233,N_19539,N_19184);
or UO_2234 (O_2234,N_19499,N_19006);
xnor UO_2235 (O_2235,N_19220,N_19198);
or UO_2236 (O_2236,N_19619,N_19921);
nand UO_2237 (O_2237,N_19319,N_19149);
and UO_2238 (O_2238,N_19581,N_19481);
nand UO_2239 (O_2239,N_19252,N_19728);
xnor UO_2240 (O_2240,N_19421,N_19640);
or UO_2241 (O_2241,N_19885,N_19826);
nand UO_2242 (O_2242,N_19167,N_19955);
xor UO_2243 (O_2243,N_19469,N_19941);
nand UO_2244 (O_2244,N_19596,N_19199);
nor UO_2245 (O_2245,N_19247,N_19984);
xnor UO_2246 (O_2246,N_19892,N_19139);
and UO_2247 (O_2247,N_19603,N_19718);
nor UO_2248 (O_2248,N_19380,N_19536);
xor UO_2249 (O_2249,N_19732,N_19376);
and UO_2250 (O_2250,N_19736,N_19478);
nor UO_2251 (O_2251,N_19398,N_19446);
nor UO_2252 (O_2252,N_19575,N_19340);
or UO_2253 (O_2253,N_19265,N_19886);
nor UO_2254 (O_2254,N_19541,N_19252);
nand UO_2255 (O_2255,N_19484,N_19795);
xnor UO_2256 (O_2256,N_19484,N_19769);
and UO_2257 (O_2257,N_19720,N_19095);
or UO_2258 (O_2258,N_19888,N_19110);
nor UO_2259 (O_2259,N_19608,N_19226);
and UO_2260 (O_2260,N_19782,N_19635);
xnor UO_2261 (O_2261,N_19423,N_19921);
nand UO_2262 (O_2262,N_19467,N_19502);
nand UO_2263 (O_2263,N_19041,N_19002);
nor UO_2264 (O_2264,N_19237,N_19978);
and UO_2265 (O_2265,N_19575,N_19692);
xor UO_2266 (O_2266,N_19624,N_19409);
or UO_2267 (O_2267,N_19950,N_19387);
nor UO_2268 (O_2268,N_19144,N_19455);
and UO_2269 (O_2269,N_19882,N_19625);
xnor UO_2270 (O_2270,N_19403,N_19592);
nor UO_2271 (O_2271,N_19539,N_19916);
xor UO_2272 (O_2272,N_19246,N_19260);
and UO_2273 (O_2273,N_19355,N_19169);
nand UO_2274 (O_2274,N_19492,N_19151);
nor UO_2275 (O_2275,N_19283,N_19176);
xor UO_2276 (O_2276,N_19469,N_19488);
xor UO_2277 (O_2277,N_19781,N_19094);
xnor UO_2278 (O_2278,N_19495,N_19057);
nor UO_2279 (O_2279,N_19044,N_19590);
or UO_2280 (O_2280,N_19066,N_19952);
nor UO_2281 (O_2281,N_19008,N_19243);
nand UO_2282 (O_2282,N_19382,N_19541);
nor UO_2283 (O_2283,N_19282,N_19414);
xor UO_2284 (O_2284,N_19331,N_19454);
nand UO_2285 (O_2285,N_19302,N_19941);
nor UO_2286 (O_2286,N_19603,N_19859);
nand UO_2287 (O_2287,N_19051,N_19629);
xnor UO_2288 (O_2288,N_19769,N_19577);
xor UO_2289 (O_2289,N_19282,N_19280);
nand UO_2290 (O_2290,N_19515,N_19517);
nor UO_2291 (O_2291,N_19514,N_19880);
nor UO_2292 (O_2292,N_19478,N_19841);
nand UO_2293 (O_2293,N_19774,N_19299);
or UO_2294 (O_2294,N_19610,N_19662);
and UO_2295 (O_2295,N_19124,N_19176);
xor UO_2296 (O_2296,N_19741,N_19242);
nor UO_2297 (O_2297,N_19720,N_19656);
xor UO_2298 (O_2298,N_19063,N_19508);
nor UO_2299 (O_2299,N_19648,N_19544);
or UO_2300 (O_2300,N_19358,N_19124);
nand UO_2301 (O_2301,N_19953,N_19233);
and UO_2302 (O_2302,N_19715,N_19271);
nand UO_2303 (O_2303,N_19428,N_19838);
nor UO_2304 (O_2304,N_19525,N_19249);
and UO_2305 (O_2305,N_19198,N_19421);
or UO_2306 (O_2306,N_19653,N_19745);
and UO_2307 (O_2307,N_19878,N_19991);
nor UO_2308 (O_2308,N_19991,N_19251);
and UO_2309 (O_2309,N_19729,N_19895);
and UO_2310 (O_2310,N_19672,N_19684);
xnor UO_2311 (O_2311,N_19389,N_19722);
or UO_2312 (O_2312,N_19907,N_19109);
nand UO_2313 (O_2313,N_19034,N_19783);
xor UO_2314 (O_2314,N_19725,N_19710);
and UO_2315 (O_2315,N_19105,N_19728);
nor UO_2316 (O_2316,N_19706,N_19189);
xor UO_2317 (O_2317,N_19464,N_19023);
and UO_2318 (O_2318,N_19152,N_19983);
and UO_2319 (O_2319,N_19539,N_19286);
and UO_2320 (O_2320,N_19884,N_19185);
nand UO_2321 (O_2321,N_19733,N_19435);
nand UO_2322 (O_2322,N_19944,N_19140);
or UO_2323 (O_2323,N_19002,N_19915);
nor UO_2324 (O_2324,N_19735,N_19829);
or UO_2325 (O_2325,N_19205,N_19676);
or UO_2326 (O_2326,N_19638,N_19333);
or UO_2327 (O_2327,N_19848,N_19524);
or UO_2328 (O_2328,N_19159,N_19504);
nand UO_2329 (O_2329,N_19001,N_19681);
xor UO_2330 (O_2330,N_19957,N_19744);
nand UO_2331 (O_2331,N_19286,N_19961);
or UO_2332 (O_2332,N_19372,N_19416);
xor UO_2333 (O_2333,N_19481,N_19582);
xor UO_2334 (O_2334,N_19096,N_19540);
nand UO_2335 (O_2335,N_19872,N_19847);
or UO_2336 (O_2336,N_19560,N_19969);
or UO_2337 (O_2337,N_19909,N_19104);
and UO_2338 (O_2338,N_19936,N_19221);
xor UO_2339 (O_2339,N_19964,N_19388);
and UO_2340 (O_2340,N_19480,N_19355);
nand UO_2341 (O_2341,N_19567,N_19177);
and UO_2342 (O_2342,N_19253,N_19353);
or UO_2343 (O_2343,N_19088,N_19874);
xor UO_2344 (O_2344,N_19354,N_19867);
or UO_2345 (O_2345,N_19919,N_19705);
or UO_2346 (O_2346,N_19159,N_19133);
and UO_2347 (O_2347,N_19368,N_19354);
nor UO_2348 (O_2348,N_19368,N_19960);
or UO_2349 (O_2349,N_19763,N_19682);
or UO_2350 (O_2350,N_19008,N_19815);
nor UO_2351 (O_2351,N_19716,N_19499);
nand UO_2352 (O_2352,N_19121,N_19130);
xor UO_2353 (O_2353,N_19089,N_19536);
nor UO_2354 (O_2354,N_19461,N_19849);
and UO_2355 (O_2355,N_19522,N_19769);
nand UO_2356 (O_2356,N_19889,N_19057);
nor UO_2357 (O_2357,N_19995,N_19129);
nor UO_2358 (O_2358,N_19465,N_19499);
or UO_2359 (O_2359,N_19226,N_19206);
nor UO_2360 (O_2360,N_19981,N_19656);
nand UO_2361 (O_2361,N_19772,N_19018);
or UO_2362 (O_2362,N_19140,N_19362);
xor UO_2363 (O_2363,N_19466,N_19110);
nor UO_2364 (O_2364,N_19732,N_19439);
and UO_2365 (O_2365,N_19992,N_19965);
nand UO_2366 (O_2366,N_19984,N_19003);
or UO_2367 (O_2367,N_19895,N_19801);
or UO_2368 (O_2368,N_19415,N_19080);
and UO_2369 (O_2369,N_19019,N_19609);
nor UO_2370 (O_2370,N_19881,N_19556);
nor UO_2371 (O_2371,N_19483,N_19903);
or UO_2372 (O_2372,N_19487,N_19769);
or UO_2373 (O_2373,N_19533,N_19138);
or UO_2374 (O_2374,N_19057,N_19887);
xor UO_2375 (O_2375,N_19988,N_19061);
nand UO_2376 (O_2376,N_19901,N_19396);
and UO_2377 (O_2377,N_19755,N_19603);
xor UO_2378 (O_2378,N_19136,N_19874);
xor UO_2379 (O_2379,N_19913,N_19517);
or UO_2380 (O_2380,N_19511,N_19527);
xnor UO_2381 (O_2381,N_19373,N_19909);
xnor UO_2382 (O_2382,N_19600,N_19435);
xnor UO_2383 (O_2383,N_19515,N_19951);
and UO_2384 (O_2384,N_19876,N_19061);
or UO_2385 (O_2385,N_19376,N_19492);
nand UO_2386 (O_2386,N_19513,N_19676);
nand UO_2387 (O_2387,N_19851,N_19680);
or UO_2388 (O_2388,N_19287,N_19853);
nand UO_2389 (O_2389,N_19372,N_19978);
xnor UO_2390 (O_2390,N_19716,N_19125);
and UO_2391 (O_2391,N_19416,N_19065);
and UO_2392 (O_2392,N_19488,N_19008);
nand UO_2393 (O_2393,N_19590,N_19130);
nor UO_2394 (O_2394,N_19005,N_19863);
nor UO_2395 (O_2395,N_19972,N_19718);
or UO_2396 (O_2396,N_19716,N_19868);
nand UO_2397 (O_2397,N_19329,N_19096);
nor UO_2398 (O_2398,N_19548,N_19253);
xor UO_2399 (O_2399,N_19414,N_19660);
nand UO_2400 (O_2400,N_19087,N_19190);
nor UO_2401 (O_2401,N_19555,N_19931);
xor UO_2402 (O_2402,N_19414,N_19531);
and UO_2403 (O_2403,N_19243,N_19598);
nor UO_2404 (O_2404,N_19798,N_19683);
or UO_2405 (O_2405,N_19432,N_19862);
nand UO_2406 (O_2406,N_19810,N_19519);
nor UO_2407 (O_2407,N_19453,N_19446);
and UO_2408 (O_2408,N_19807,N_19987);
nor UO_2409 (O_2409,N_19880,N_19663);
nor UO_2410 (O_2410,N_19864,N_19739);
and UO_2411 (O_2411,N_19928,N_19591);
or UO_2412 (O_2412,N_19665,N_19145);
or UO_2413 (O_2413,N_19018,N_19119);
and UO_2414 (O_2414,N_19631,N_19398);
and UO_2415 (O_2415,N_19416,N_19976);
and UO_2416 (O_2416,N_19193,N_19187);
xor UO_2417 (O_2417,N_19723,N_19302);
or UO_2418 (O_2418,N_19184,N_19235);
nand UO_2419 (O_2419,N_19230,N_19350);
nor UO_2420 (O_2420,N_19527,N_19492);
nand UO_2421 (O_2421,N_19910,N_19376);
or UO_2422 (O_2422,N_19615,N_19931);
nor UO_2423 (O_2423,N_19344,N_19330);
and UO_2424 (O_2424,N_19768,N_19127);
and UO_2425 (O_2425,N_19394,N_19223);
and UO_2426 (O_2426,N_19950,N_19861);
or UO_2427 (O_2427,N_19658,N_19066);
and UO_2428 (O_2428,N_19728,N_19300);
and UO_2429 (O_2429,N_19956,N_19847);
and UO_2430 (O_2430,N_19440,N_19668);
and UO_2431 (O_2431,N_19296,N_19862);
nor UO_2432 (O_2432,N_19696,N_19453);
xor UO_2433 (O_2433,N_19490,N_19481);
and UO_2434 (O_2434,N_19631,N_19199);
or UO_2435 (O_2435,N_19702,N_19061);
nand UO_2436 (O_2436,N_19371,N_19637);
and UO_2437 (O_2437,N_19550,N_19878);
nor UO_2438 (O_2438,N_19983,N_19960);
xnor UO_2439 (O_2439,N_19599,N_19915);
xnor UO_2440 (O_2440,N_19683,N_19604);
or UO_2441 (O_2441,N_19812,N_19015);
or UO_2442 (O_2442,N_19675,N_19125);
xor UO_2443 (O_2443,N_19998,N_19919);
and UO_2444 (O_2444,N_19275,N_19695);
xor UO_2445 (O_2445,N_19139,N_19405);
xor UO_2446 (O_2446,N_19832,N_19252);
and UO_2447 (O_2447,N_19006,N_19447);
nor UO_2448 (O_2448,N_19755,N_19578);
or UO_2449 (O_2449,N_19746,N_19397);
and UO_2450 (O_2450,N_19256,N_19250);
and UO_2451 (O_2451,N_19017,N_19617);
or UO_2452 (O_2452,N_19955,N_19785);
and UO_2453 (O_2453,N_19807,N_19395);
nor UO_2454 (O_2454,N_19003,N_19762);
xor UO_2455 (O_2455,N_19692,N_19992);
nor UO_2456 (O_2456,N_19077,N_19575);
or UO_2457 (O_2457,N_19938,N_19835);
xor UO_2458 (O_2458,N_19921,N_19469);
or UO_2459 (O_2459,N_19608,N_19485);
and UO_2460 (O_2460,N_19628,N_19885);
xnor UO_2461 (O_2461,N_19175,N_19351);
nand UO_2462 (O_2462,N_19928,N_19342);
and UO_2463 (O_2463,N_19130,N_19663);
xor UO_2464 (O_2464,N_19504,N_19918);
or UO_2465 (O_2465,N_19395,N_19066);
or UO_2466 (O_2466,N_19554,N_19346);
and UO_2467 (O_2467,N_19993,N_19913);
or UO_2468 (O_2468,N_19404,N_19054);
or UO_2469 (O_2469,N_19722,N_19404);
nand UO_2470 (O_2470,N_19094,N_19925);
nor UO_2471 (O_2471,N_19370,N_19749);
xor UO_2472 (O_2472,N_19703,N_19267);
or UO_2473 (O_2473,N_19350,N_19475);
and UO_2474 (O_2474,N_19329,N_19225);
nand UO_2475 (O_2475,N_19480,N_19104);
nor UO_2476 (O_2476,N_19050,N_19231);
nor UO_2477 (O_2477,N_19780,N_19179);
nand UO_2478 (O_2478,N_19639,N_19649);
nor UO_2479 (O_2479,N_19399,N_19589);
nand UO_2480 (O_2480,N_19986,N_19681);
nor UO_2481 (O_2481,N_19012,N_19698);
nand UO_2482 (O_2482,N_19668,N_19388);
or UO_2483 (O_2483,N_19437,N_19710);
xor UO_2484 (O_2484,N_19686,N_19798);
nand UO_2485 (O_2485,N_19230,N_19110);
nor UO_2486 (O_2486,N_19260,N_19720);
or UO_2487 (O_2487,N_19134,N_19080);
xnor UO_2488 (O_2488,N_19735,N_19135);
xnor UO_2489 (O_2489,N_19169,N_19624);
nor UO_2490 (O_2490,N_19633,N_19891);
xor UO_2491 (O_2491,N_19175,N_19287);
xnor UO_2492 (O_2492,N_19660,N_19612);
and UO_2493 (O_2493,N_19555,N_19475);
and UO_2494 (O_2494,N_19017,N_19493);
nor UO_2495 (O_2495,N_19093,N_19016);
xor UO_2496 (O_2496,N_19086,N_19702);
xor UO_2497 (O_2497,N_19164,N_19989);
and UO_2498 (O_2498,N_19912,N_19477);
nand UO_2499 (O_2499,N_19243,N_19999);
endmodule