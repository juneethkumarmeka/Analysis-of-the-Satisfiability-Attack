module basic_500_3000_500_60_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_235,In_285);
or U1 (N_1,In_193,In_173);
xnor U2 (N_2,In_280,In_465);
and U3 (N_3,In_141,In_375);
nand U4 (N_4,In_300,In_403);
nand U5 (N_5,In_314,In_263);
or U6 (N_6,In_367,In_80);
and U7 (N_7,In_443,In_304);
nor U8 (N_8,In_196,In_366);
or U9 (N_9,In_311,In_395);
or U10 (N_10,In_270,In_117);
nand U11 (N_11,In_298,In_237);
nand U12 (N_12,In_136,In_12);
nand U13 (N_13,In_355,In_50);
and U14 (N_14,In_137,In_215);
nand U15 (N_15,In_216,In_174);
nand U16 (N_16,In_209,In_8);
nor U17 (N_17,In_428,In_365);
or U18 (N_18,In_2,In_369);
and U19 (N_19,In_473,In_218);
nand U20 (N_20,In_13,In_75);
nor U21 (N_21,In_37,In_98);
nand U22 (N_22,In_373,In_497);
or U23 (N_23,In_390,In_214);
nand U24 (N_24,In_84,In_289);
or U25 (N_25,In_102,In_64);
and U26 (N_26,In_199,In_406);
or U27 (N_27,In_422,In_415);
xor U28 (N_28,In_339,In_192);
and U29 (N_29,In_79,In_125);
and U30 (N_30,In_330,In_3);
or U31 (N_31,In_161,In_150);
nor U32 (N_32,In_7,In_187);
or U33 (N_33,In_316,In_165);
or U34 (N_34,In_97,In_88);
nor U35 (N_35,In_38,In_43);
or U36 (N_36,In_156,In_59);
or U37 (N_37,In_31,In_384);
nand U38 (N_38,In_434,In_106);
xnor U39 (N_39,In_85,In_456);
or U40 (N_40,In_252,In_198);
nand U41 (N_41,In_206,In_423);
nand U42 (N_42,In_387,In_421);
nor U43 (N_43,In_128,In_34);
or U44 (N_44,In_66,In_19);
nor U45 (N_45,In_377,In_323);
nand U46 (N_46,In_112,In_155);
nor U47 (N_47,In_472,In_120);
and U48 (N_48,In_325,In_114);
nand U49 (N_49,In_474,In_337);
and U50 (N_50,In_20,In_310);
or U51 (N_51,In_246,In_36);
or U52 (N_52,In_479,In_159);
or U53 (N_53,In_460,In_4);
nor U54 (N_54,In_457,In_210);
and U55 (N_55,In_255,In_205);
or U56 (N_56,In_5,N_15);
or U57 (N_57,In_54,In_27);
nor U58 (N_58,In_153,In_332);
nand U59 (N_59,In_291,In_445);
and U60 (N_60,In_105,In_96);
and U61 (N_61,N_48,In_33);
nand U62 (N_62,In_267,In_327);
or U63 (N_63,In_251,In_394);
nor U64 (N_64,In_25,In_130);
nor U65 (N_65,In_249,In_135);
nand U66 (N_66,In_78,N_30);
nor U67 (N_67,In_157,In_48);
or U68 (N_68,In_259,In_308);
nor U69 (N_69,In_348,In_55);
nor U70 (N_70,In_162,In_121);
or U71 (N_71,In_132,In_74);
and U72 (N_72,In_463,N_10);
nand U73 (N_73,In_49,In_295);
nor U74 (N_74,In_283,N_18);
nor U75 (N_75,In_356,In_454);
nor U76 (N_76,In_405,In_494);
or U77 (N_77,In_306,In_35);
or U78 (N_78,In_233,In_389);
nor U79 (N_79,In_475,In_69);
nand U80 (N_80,In_315,In_363);
nand U81 (N_81,In_212,In_116);
nand U82 (N_82,In_499,N_5);
nor U83 (N_83,In_274,N_1);
nand U84 (N_84,In_317,In_437);
nand U85 (N_85,In_73,In_119);
nor U86 (N_86,In_224,In_410);
nand U87 (N_87,In_213,In_253);
or U88 (N_88,In_359,In_420);
nand U89 (N_89,In_228,In_110);
nor U90 (N_90,In_440,In_483);
or U91 (N_91,N_40,In_368);
nand U92 (N_92,In_493,In_232);
nor U93 (N_93,In_399,In_379);
and U94 (N_94,In_430,In_133);
nand U95 (N_95,In_427,In_63);
nand U96 (N_96,In_186,In_262);
nor U97 (N_97,In_487,In_383);
nand U98 (N_98,In_417,N_0);
nor U99 (N_99,In_294,In_413);
nand U100 (N_100,In_385,In_335);
and U101 (N_101,In_482,N_57);
and U102 (N_102,N_92,In_189);
nand U103 (N_103,In_15,In_240);
nor U104 (N_104,In_83,In_14);
nand U105 (N_105,In_392,In_123);
nand U106 (N_106,In_435,In_416);
nor U107 (N_107,N_59,In_201);
or U108 (N_108,N_36,In_490);
and U109 (N_109,In_451,N_4);
nor U110 (N_110,In_361,In_245);
and U111 (N_111,N_27,N_74);
and U112 (N_112,In_127,In_239);
nand U113 (N_113,In_190,N_81);
nor U114 (N_114,N_21,In_424);
nor U115 (N_115,In_269,In_197);
nor U116 (N_116,In_146,In_352);
nor U117 (N_117,In_380,In_254);
nor U118 (N_118,N_87,In_21);
and U119 (N_119,In_113,In_154);
and U120 (N_120,N_35,In_93);
nand U121 (N_121,N_62,In_202);
and U122 (N_122,In_400,In_293);
and U123 (N_123,N_76,In_476);
nand U124 (N_124,In_183,In_250);
nand U125 (N_125,In_271,N_38);
nor U126 (N_126,In_126,In_203);
and U127 (N_127,In_452,In_24);
nor U128 (N_128,N_22,In_322);
nand U129 (N_129,N_50,In_324);
nor U130 (N_130,N_14,N_96);
nor U131 (N_131,In_182,In_360);
nor U132 (N_132,In_195,In_211);
and U133 (N_133,In_151,In_370);
nor U134 (N_134,In_458,In_53);
nor U135 (N_135,In_168,N_28);
nand U136 (N_136,In_6,In_477);
and U137 (N_137,In_260,In_343);
and U138 (N_138,In_188,N_80);
and U139 (N_139,N_17,In_222);
nand U140 (N_140,In_450,In_70);
and U141 (N_141,In_408,In_71);
and U142 (N_142,In_30,In_495);
nand U143 (N_143,N_43,N_9);
nor U144 (N_144,In_47,N_58);
or U145 (N_145,In_234,In_144);
or U146 (N_146,In_362,N_16);
nor U147 (N_147,In_286,In_398);
nand U148 (N_148,In_175,In_200);
nand U149 (N_149,In_23,In_277);
and U150 (N_150,In_1,N_100);
nand U151 (N_151,In_320,N_108);
and U152 (N_152,In_409,In_22);
nor U153 (N_153,In_459,In_299);
or U154 (N_154,In_393,In_426);
nor U155 (N_155,N_132,N_53);
and U156 (N_156,In_76,N_149);
nor U157 (N_157,In_118,In_122);
and U158 (N_158,In_171,In_347);
nand U159 (N_159,N_140,In_404);
nand U160 (N_160,N_85,In_436);
and U161 (N_161,N_42,In_229);
nor U162 (N_162,In_107,N_11);
nand U163 (N_163,N_12,In_185);
xnor U164 (N_164,N_23,N_65);
or U165 (N_165,In_328,In_492);
nand U166 (N_166,N_95,In_449);
or U167 (N_167,In_484,In_194);
nor U168 (N_168,In_431,In_284);
and U169 (N_169,N_56,In_301);
or U170 (N_170,N_60,In_414);
or U171 (N_171,In_276,In_433);
nand U172 (N_172,In_464,N_116);
nand U173 (N_173,In_344,In_397);
or U174 (N_174,N_120,In_396);
and U175 (N_175,In_108,In_138);
and U176 (N_176,In_318,N_147);
or U177 (N_177,N_98,N_110);
nor U178 (N_178,In_147,In_331);
and U179 (N_179,In_86,N_148);
nor U180 (N_180,N_107,In_100);
or U181 (N_181,In_103,N_138);
nand U182 (N_182,In_358,N_121);
or U183 (N_183,In_39,In_401);
and U184 (N_184,In_104,N_139);
and U185 (N_185,In_230,In_419);
or U186 (N_186,In_45,In_378);
and U187 (N_187,In_382,N_142);
nor U188 (N_188,In_208,In_371);
and U189 (N_189,In_461,In_241);
and U190 (N_190,N_117,In_256);
nand U191 (N_191,In_388,In_17);
or U192 (N_192,In_444,In_455);
xor U193 (N_193,In_264,N_25);
or U194 (N_194,N_88,In_496);
or U195 (N_195,In_16,In_288);
and U196 (N_196,N_86,In_28);
and U197 (N_197,In_225,In_468);
or U198 (N_198,N_61,In_124);
or U199 (N_199,In_160,In_134);
nor U200 (N_200,In_462,N_141);
or U201 (N_201,In_471,In_91);
or U202 (N_202,In_296,N_90);
and U203 (N_203,N_131,N_69);
or U204 (N_204,In_470,In_65);
nand U205 (N_205,N_68,In_488);
or U206 (N_206,In_244,N_186);
nor U207 (N_207,N_73,In_9);
and U208 (N_208,In_257,N_44);
and U209 (N_209,N_172,In_350);
xnor U210 (N_210,In_176,In_439);
or U211 (N_211,N_99,In_302);
and U212 (N_212,N_34,N_105);
and U213 (N_213,In_184,In_207);
nor U214 (N_214,N_176,In_340);
nand U215 (N_215,N_51,In_341);
or U216 (N_216,N_29,In_204);
nand U217 (N_217,N_170,In_447);
and U218 (N_218,N_163,N_133);
nand U219 (N_219,N_125,N_89);
nor U220 (N_220,In_41,In_219);
or U221 (N_221,N_79,In_61);
or U222 (N_222,In_334,In_411);
and U223 (N_223,N_192,In_307);
nor U224 (N_224,In_469,N_181);
and U225 (N_225,N_97,N_93);
nor U226 (N_226,In_51,In_172);
xor U227 (N_227,N_8,N_145);
and U228 (N_228,N_166,In_467);
nand U229 (N_229,In_217,In_478);
nor U230 (N_230,In_489,N_111);
nand U231 (N_231,In_72,In_129);
and U232 (N_232,N_54,N_157);
and U233 (N_233,N_182,In_143);
nand U234 (N_234,In_170,N_197);
nor U235 (N_235,In_305,N_196);
and U236 (N_236,In_167,N_143);
nor U237 (N_237,N_164,In_261);
and U238 (N_238,In_231,N_83);
or U239 (N_239,N_144,In_418);
nor U240 (N_240,In_177,N_137);
nand U241 (N_241,In_158,In_92);
nor U242 (N_242,In_412,In_491);
nand U243 (N_243,In_272,N_115);
and U244 (N_244,N_180,N_199);
nand U245 (N_245,N_102,In_429);
nand U246 (N_246,N_67,In_345);
and U247 (N_247,In_247,In_221);
and U248 (N_248,In_407,N_185);
nand U249 (N_249,In_312,N_31);
and U250 (N_250,In_111,In_220);
or U251 (N_251,In_166,In_275);
or U252 (N_252,In_32,N_104);
or U253 (N_253,In_139,In_226);
nor U254 (N_254,N_198,N_128);
nor U255 (N_255,In_346,In_140);
nor U256 (N_256,In_145,In_376);
or U257 (N_257,In_268,N_150);
nand U258 (N_258,In_321,N_179);
nor U259 (N_259,N_154,N_194);
nor U260 (N_260,In_101,In_90);
or U261 (N_261,In_364,N_201);
and U262 (N_262,N_231,N_243);
nand U263 (N_263,N_106,N_24);
nand U264 (N_264,In_178,In_372);
and U265 (N_265,In_142,N_118);
and U266 (N_266,N_63,N_153);
nor U267 (N_267,In_448,In_18);
and U268 (N_268,In_223,N_227);
or U269 (N_269,In_67,In_57);
and U270 (N_270,In_56,In_248);
and U271 (N_271,In_10,N_13);
and U272 (N_272,N_211,N_204);
or U273 (N_273,N_2,In_386);
and U274 (N_274,N_217,N_177);
and U275 (N_275,In_309,N_225);
nor U276 (N_276,In_115,In_0);
nand U277 (N_277,N_190,In_68);
nand U278 (N_278,N_20,In_297);
and U279 (N_279,N_39,In_354);
nand U280 (N_280,N_112,N_103);
nor U281 (N_281,N_242,N_205);
and U282 (N_282,In_303,N_214);
and U283 (N_283,N_151,In_453);
nor U284 (N_284,In_40,N_241);
nor U285 (N_285,N_174,N_49);
or U286 (N_286,N_200,N_208);
nand U287 (N_287,In_243,In_148);
or U288 (N_288,N_240,In_336);
and U289 (N_289,N_213,N_169);
nand U290 (N_290,In_77,In_273);
nand U291 (N_291,N_126,N_124);
nor U292 (N_292,N_233,N_158);
or U293 (N_293,N_187,N_41);
or U294 (N_294,In_438,N_32);
and U295 (N_295,N_75,In_442);
or U296 (N_296,N_220,In_402);
nand U297 (N_297,N_70,N_171);
nor U298 (N_298,N_77,N_152);
nor U299 (N_299,In_164,In_58);
xnor U300 (N_300,N_3,N_247);
nor U301 (N_301,In_169,In_381);
and U302 (N_302,N_202,N_155);
or U303 (N_303,N_284,In_480);
and U304 (N_304,In_179,N_258);
nand U305 (N_305,N_299,N_266);
nand U306 (N_306,N_239,In_446);
nor U307 (N_307,N_160,In_498);
nor U308 (N_308,N_275,N_191);
nor U309 (N_309,N_215,In_26);
or U310 (N_310,N_184,N_290);
nor U311 (N_311,In_374,N_210);
and U312 (N_312,In_95,In_342);
and U313 (N_313,N_251,N_26);
and U314 (N_314,N_216,In_109);
and U315 (N_315,In_265,In_81);
nand U316 (N_316,N_101,N_272);
and U317 (N_317,N_249,N_55);
and U318 (N_318,N_113,In_152);
nand U319 (N_319,N_203,N_52);
nor U320 (N_320,N_156,N_223);
nor U321 (N_321,N_235,N_298);
or U322 (N_322,N_254,In_391);
or U323 (N_323,N_159,N_123);
and U324 (N_324,In_353,N_168);
and U325 (N_325,In_163,N_6);
and U326 (N_326,N_269,In_46);
and U327 (N_327,N_193,N_206);
and U328 (N_328,In_290,N_134);
and U329 (N_329,N_183,N_189);
or U330 (N_330,N_130,N_218);
or U331 (N_331,In_149,N_221);
or U332 (N_332,N_122,In_441);
xnor U333 (N_333,N_271,N_47);
or U334 (N_334,N_78,N_82);
and U335 (N_335,N_33,N_244);
nand U336 (N_336,In_313,N_222);
nand U337 (N_337,In_349,In_287);
nand U338 (N_338,N_136,N_219);
and U339 (N_339,In_62,N_91);
nor U340 (N_340,In_60,N_281);
nand U341 (N_341,In_42,N_37);
or U342 (N_342,In_82,N_256);
nand U343 (N_343,N_232,N_229);
or U344 (N_344,N_276,N_277);
nor U345 (N_345,N_293,N_267);
or U346 (N_346,In_281,N_165);
nor U347 (N_347,N_175,N_257);
nor U348 (N_348,In_319,In_191);
nand U349 (N_349,In_258,N_294);
or U350 (N_350,N_296,N_255);
nand U351 (N_351,N_94,N_332);
and U352 (N_352,In_94,N_318);
nor U353 (N_353,N_234,In_326);
nor U354 (N_354,N_119,In_333);
and U355 (N_355,N_334,N_270);
and U356 (N_356,N_308,N_135);
or U357 (N_357,N_348,In_180);
nand U358 (N_358,N_146,N_84);
or U359 (N_359,In_279,In_485);
nor U360 (N_360,N_209,N_311);
nor U361 (N_361,N_72,N_273);
and U362 (N_362,N_288,N_129);
nor U363 (N_363,N_291,In_181);
or U364 (N_364,N_336,N_321);
or U365 (N_365,N_283,N_228);
and U366 (N_366,N_167,N_64);
or U367 (N_367,N_319,N_302);
nor U368 (N_368,N_268,N_320);
or U369 (N_369,N_304,N_330);
and U370 (N_370,N_301,In_338);
or U371 (N_371,N_248,In_329);
nand U372 (N_372,N_323,N_7);
or U373 (N_373,N_341,N_340);
nand U374 (N_374,N_345,N_114);
and U375 (N_375,N_173,N_260);
or U376 (N_376,In_351,N_286);
and U377 (N_377,N_324,N_226);
nor U378 (N_378,N_224,N_127);
nand U379 (N_379,In_238,N_188);
or U380 (N_380,N_282,In_486);
nand U381 (N_381,N_45,N_245);
and U382 (N_382,In_44,N_305);
nor U383 (N_383,N_71,N_287);
nand U384 (N_384,N_252,In_52);
or U385 (N_385,N_238,N_212);
or U386 (N_386,N_325,N_262);
nand U387 (N_387,N_313,In_425);
or U388 (N_388,N_316,N_161);
nor U389 (N_389,N_295,In_11);
and U390 (N_390,N_317,N_261);
nor U391 (N_391,N_339,N_322);
nor U392 (N_392,N_109,N_19);
nor U393 (N_393,In_87,N_178);
nand U394 (N_394,N_280,N_309);
or U395 (N_395,N_289,N_285);
or U396 (N_396,N_162,In_481);
xnor U397 (N_397,N_315,N_195);
nand U398 (N_398,N_274,N_259);
nor U399 (N_399,N_230,N_297);
xor U400 (N_400,N_355,N_337);
nand U401 (N_401,N_300,N_331);
nand U402 (N_402,N_312,N_307);
nand U403 (N_403,N_343,N_314);
nand U404 (N_404,N_354,N_381);
or U405 (N_405,N_326,N_375);
nor U406 (N_406,N_346,N_46);
and U407 (N_407,N_398,N_376);
or U408 (N_408,N_394,In_236);
or U409 (N_409,N_265,In_432);
and U410 (N_410,N_385,N_357);
and U411 (N_411,N_368,N_379);
nand U412 (N_412,N_396,N_374);
and U413 (N_413,In_29,N_328);
nand U414 (N_414,N_350,N_253);
and U415 (N_415,N_263,N_360);
nand U416 (N_416,N_393,In_466);
nor U417 (N_417,N_395,N_386);
and U418 (N_418,In_131,In_242);
nor U419 (N_419,In_99,N_236);
and U420 (N_420,N_391,N_384);
and U421 (N_421,In_357,N_382);
and U422 (N_422,N_358,N_66);
or U423 (N_423,N_363,N_278);
and U424 (N_424,N_370,N_369);
and U425 (N_425,N_389,N_303);
or U426 (N_426,N_392,In_89);
and U427 (N_427,N_377,N_383);
xnor U428 (N_428,N_292,In_282);
and U429 (N_429,N_342,N_327);
and U430 (N_430,N_353,N_371);
or U431 (N_431,N_250,N_378);
nand U432 (N_432,N_364,N_347);
nor U433 (N_433,N_356,In_227);
or U434 (N_434,N_397,N_329);
nand U435 (N_435,N_344,N_361);
and U436 (N_436,N_306,N_380);
or U437 (N_437,N_390,In_292);
nand U438 (N_438,N_237,N_246);
and U439 (N_439,N_388,N_373);
or U440 (N_440,N_264,N_335);
or U441 (N_441,N_387,In_278);
or U442 (N_442,N_338,N_349);
and U443 (N_443,N_359,N_333);
or U444 (N_444,N_366,N_351);
nand U445 (N_445,N_362,In_266);
nor U446 (N_446,N_207,N_310);
and U447 (N_447,N_367,N_279);
and U448 (N_448,N_399,N_365);
nand U449 (N_449,N_372,N_352);
or U450 (N_450,N_443,N_425);
nor U451 (N_451,N_404,N_440);
nand U452 (N_452,N_412,N_424);
nor U453 (N_453,N_442,N_417);
nand U454 (N_454,N_436,N_421);
and U455 (N_455,N_439,N_433);
nand U456 (N_456,N_407,N_441);
or U457 (N_457,N_422,N_448);
nor U458 (N_458,N_449,N_408);
and U459 (N_459,N_410,N_405);
nand U460 (N_460,N_438,N_413);
nor U461 (N_461,N_423,N_401);
and U462 (N_462,N_428,N_429);
nand U463 (N_463,N_434,N_409);
nand U464 (N_464,N_427,N_403);
or U465 (N_465,N_414,N_430);
and U466 (N_466,N_416,N_444);
or U467 (N_467,N_402,N_411);
and U468 (N_468,N_426,N_420);
and U469 (N_469,N_431,N_406);
or U470 (N_470,N_418,N_437);
or U471 (N_471,N_419,N_446);
nor U472 (N_472,N_447,N_432);
or U473 (N_473,N_445,N_415);
or U474 (N_474,N_435,N_400);
nand U475 (N_475,N_422,N_420);
nand U476 (N_476,N_409,N_440);
nand U477 (N_477,N_448,N_431);
or U478 (N_478,N_443,N_416);
and U479 (N_479,N_407,N_414);
and U480 (N_480,N_419,N_412);
and U481 (N_481,N_419,N_414);
or U482 (N_482,N_443,N_441);
nor U483 (N_483,N_447,N_413);
or U484 (N_484,N_421,N_407);
nand U485 (N_485,N_435,N_405);
and U486 (N_486,N_441,N_418);
nand U487 (N_487,N_420,N_441);
or U488 (N_488,N_415,N_414);
or U489 (N_489,N_414,N_402);
nand U490 (N_490,N_401,N_407);
nand U491 (N_491,N_403,N_410);
nor U492 (N_492,N_425,N_430);
nand U493 (N_493,N_419,N_429);
nor U494 (N_494,N_432,N_401);
nor U495 (N_495,N_431,N_400);
nor U496 (N_496,N_417,N_444);
nor U497 (N_497,N_405,N_420);
nand U498 (N_498,N_429,N_431);
or U499 (N_499,N_417,N_425);
nand U500 (N_500,N_492,N_464);
and U501 (N_501,N_461,N_498);
and U502 (N_502,N_472,N_479);
or U503 (N_503,N_469,N_477);
nand U504 (N_504,N_494,N_476);
nor U505 (N_505,N_473,N_485);
and U506 (N_506,N_491,N_490);
or U507 (N_507,N_474,N_456);
nor U508 (N_508,N_486,N_482);
nand U509 (N_509,N_470,N_468);
nor U510 (N_510,N_450,N_496);
nand U511 (N_511,N_493,N_481);
or U512 (N_512,N_465,N_457);
nor U513 (N_513,N_454,N_488);
nor U514 (N_514,N_483,N_475);
nand U515 (N_515,N_471,N_480);
and U516 (N_516,N_467,N_478);
and U517 (N_517,N_463,N_466);
nand U518 (N_518,N_460,N_459);
and U519 (N_519,N_462,N_453);
or U520 (N_520,N_499,N_495);
and U521 (N_521,N_497,N_458);
and U522 (N_522,N_451,N_452);
and U523 (N_523,N_484,N_489);
and U524 (N_524,N_487,N_455);
or U525 (N_525,N_451,N_455);
nand U526 (N_526,N_460,N_474);
or U527 (N_527,N_469,N_484);
and U528 (N_528,N_469,N_488);
or U529 (N_529,N_499,N_476);
and U530 (N_530,N_498,N_482);
or U531 (N_531,N_464,N_498);
nand U532 (N_532,N_459,N_462);
and U533 (N_533,N_451,N_498);
or U534 (N_534,N_472,N_461);
nand U535 (N_535,N_468,N_466);
nor U536 (N_536,N_498,N_477);
nand U537 (N_537,N_476,N_477);
or U538 (N_538,N_491,N_462);
or U539 (N_539,N_454,N_489);
nand U540 (N_540,N_493,N_456);
and U541 (N_541,N_465,N_453);
and U542 (N_542,N_498,N_476);
nand U543 (N_543,N_480,N_469);
and U544 (N_544,N_470,N_451);
and U545 (N_545,N_479,N_458);
and U546 (N_546,N_480,N_492);
nor U547 (N_547,N_493,N_497);
or U548 (N_548,N_463,N_485);
nand U549 (N_549,N_495,N_492);
or U550 (N_550,N_513,N_527);
and U551 (N_551,N_541,N_508);
nand U552 (N_552,N_517,N_547);
nand U553 (N_553,N_539,N_536);
or U554 (N_554,N_531,N_544);
nand U555 (N_555,N_514,N_523);
nor U556 (N_556,N_528,N_537);
and U557 (N_557,N_545,N_504);
nor U558 (N_558,N_515,N_533);
and U559 (N_559,N_525,N_524);
nor U560 (N_560,N_538,N_518);
nand U561 (N_561,N_530,N_510);
nor U562 (N_562,N_500,N_507);
nand U563 (N_563,N_520,N_540);
xnor U564 (N_564,N_521,N_502);
or U565 (N_565,N_526,N_503);
nor U566 (N_566,N_506,N_501);
and U567 (N_567,N_534,N_505);
and U568 (N_568,N_532,N_549);
nor U569 (N_569,N_512,N_522);
nor U570 (N_570,N_548,N_542);
nor U571 (N_571,N_546,N_535);
xor U572 (N_572,N_543,N_516);
and U573 (N_573,N_519,N_509);
or U574 (N_574,N_511,N_529);
and U575 (N_575,N_523,N_526);
and U576 (N_576,N_543,N_509);
and U577 (N_577,N_512,N_521);
nand U578 (N_578,N_525,N_547);
nand U579 (N_579,N_510,N_517);
or U580 (N_580,N_525,N_540);
or U581 (N_581,N_542,N_529);
nor U582 (N_582,N_536,N_508);
nor U583 (N_583,N_516,N_508);
or U584 (N_584,N_533,N_504);
and U585 (N_585,N_519,N_503);
or U586 (N_586,N_543,N_514);
nor U587 (N_587,N_513,N_544);
nand U588 (N_588,N_547,N_535);
or U589 (N_589,N_536,N_504);
and U590 (N_590,N_519,N_547);
nand U591 (N_591,N_542,N_507);
nand U592 (N_592,N_544,N_529);
nand U593 (N_593,N_510,N_546);
nand U594 (N_594,N_523,N_529);
or U595 (N_595,N_505,N_509);
nand U596 (N_596,N_504,N_507);
nor U597 (N_597,N_539,N_526);
nor U598 (N_598,N_523,N_500);
and U599 (N_599,N_538,N_504);
nand U600 (N_600,N_590,N_592);
or U601 (N_601,N_563,N_598);
nand U602 (N_602,N_589,N_585);
or U603 (N_603,N_568,N_558);
or U604 (N_604,N_583,N_565);
and U605 (N_605,N_569,N_557);
nor U606 (N_606,N_580,N_582);
or U607 (N_607,N_571,N_560);
nor U608 (N_608,N_562,N_564);
or U609 (N_609,N_593,N_599);
nand U610 (N_610,N_595,N_566);
nand U611 (N_611,N_579,N_573);
and U612 (N_612,N_597,N_554);
nand U613 (N_613,N_581,N_551);
nor U614 (N_614,N_596,N_572);
or U615 (N_615,N_584,N_556);
and U616 (N_616,N_587,N_570);
nor U617 (N_617,N_591,N_574);
nand U618 (N_618,N_586,N_594);
and U619 (N_619,N_550,N_588);
nor U620 (N_620,N_552,N_561);
nand U621 (N_621,N_553,N_555);
and U622 (N_622,N_576,N_575);
nor U623 (N_623,N_567,N_577);
nand U624 (N_624,N_578,N_559);
nand U625 (N_625,N_588,N_574);
and U626 (N_626,N_586,N_589);
or U627 (N_627,N_591,N_577);
or U628 (N_628,N_584,N_592);
nand U629 (N_629,N_560,N_551);
nor U630 (N_630,N_573,N_597);
or U631 (N_631,N_583,N_552);
nor U632 (N_632,N_595,N_570);
nor U633 (N_633,N_551,N_553);
and U634 (N_634,N_559,N_555);
and U635 (N_635,N_590,N_551);
and U636 (N_636,N_599,N_574);
or U637 (N_637,N_559,N_556);
nand U638 (N_638,N_571,N_563);
nand U639 (N_639,N_599,N_589);
and U640 (N_640,N_577,N_585);
or U641 (N_641,N_592,N_556);
and U642 (N_642,N_558,N_597);
nor U643 (N_643,N_577,N_552);
nor U644 (N_644,N_578,N_580);
or U645 (N_645,N_557,N_581);
or U646 (N_646,N_557,N_561);
nor U647 (N_647,N_576,N_551);
nand U648 (N_648,N_575,N_594);
nand U649 (N_649,N_551,N_579);
and U650 (N_650,N_626,N_632);
or U651 (N_651,N_624,N_610);
or U652 (N_652,N_623,N_619);
nand U653 (N_653,N_600,N_641);
or U654 (N_654,N_643,N_627);
and U655 (N_655,N_630,N_649);
nor U656 (N_656,N_604,N_606);
nand U657 (N_657,N_618,N_602);
or U658 (N_658,N_640,N_638);
or U659 (N_659,N_634,N_646);
or U660 (N_660,N_635,N_628);
nor U661 (N_661,N_636,N_612);
nand U662 (N_662,N_629,N_607);
and U663 (N_663,N_609,N_603);
or U664 (N_664,N_642,N_621);
and U665 (N_665,N_625,N_648);
and U666 (N_666,N_622,N_620);
nor U667 (N_667,N_614,N_605);
or U668 (N_668,N_644,N_645);
nor U669 (N_669,N_617,N_639);
nand U670 (N_670,N_616,N_613);
or U671 (N_671,N_637,N_608);
nand U672 (N_672,N_601,N_647);
and U673 (N_673,N_633,N_611);
and U674 (N_674,N_631,N_615);
or U675 (N_675,N_607,N_626);
or U676 (N_676,N_625,N_629);
or U677 (N_677,N_634,N_609);
or U678 (N_678,N_627,N_615);
nand U679 (N_679,N_629,N_600);
nor U680 (N_680,N_603,N_620);
nor U681 (N_681,N_616,N_603);
or U682 (N_682,N_627,N_617);
nor U683 (N_683,N_629,N_619);
and U684 (N_684,N_605,N_616);
and U685 (N_685,N_641,N_622);
nand U686 (N_686,N_638,N_609);
nand U687 (N_687,N_610,N_604);
nor U688 (N_688,N_638,N_634);
nand U689 (N_689,N_612,N_646);
or U690 (N_690,N_608,N_603);
or U691 (N_691,N_639,N_607);
nor U692 (N_692,N_635,N_623);
or U693 (N_693,N_633,N_640);
or U694 (N_694,N_615,N_611);
or U695 (N_695,N_607,N_617);
nand U696 (N_696,N_643,N_610);
nand U697 (N_697,N_617,N_619);
or U698 (N_698,N_622,N_631);
nand U699 (N_699,N_612,N_625);
or U700 (N_700,N_662,N_697);
or U701 (N_701,N_671,N_675);
and U702 (N_702,N_683,N_693);
nor U703 (N_703,N_684,N_650);
or U704 (N_704,N_695,N_664);
or U705 (N_705,N_677,N_690);
nor U706 (N_706,N_694,N_669);
or U707 (N_707,N_656,N_670);
or U708 (N_708,N_667,N_685);
or U709 (N_709,N_660,N_666);
nand U710 (N_710,N_692,N_679);
or U711 (N_711,N_680,N_682);
nand U712 (N_712,N_681,N_699);
or U713 (N_713,N_651,N_673);
nand U714 (N_714,N_691,N_676);
nand U715 (N_715,N_659,N_665);
and U716 (N_716,N_655,N_696);
and U717 (N_717,N_686,N_678);
or U718 (N_718,N_698,N_672);
nand U719 (N_719,N_653,N_689);
nand U720 (N_720,N_674,N_663);
nor U721 (N_721,N_668,N_687);
nand U722 (N_722,N_661,N_688);
nor U723 (N_723,N_654,N_658);
or U724 (N_724,N_657,N_652);
nor U725 (N_725,N_652,N_691);
nand U726 (N_726,N_694,N_698);
and U727 (N_727,N_664,N_655);
nor U728 (N_728,N_660,N_694);
or U729 (N_729,N_687,N_693);
nand U730 (N_730,N_680,N_652);
nand U731 (N_731,N_661,N_669);
nor U732 (N_732,N_667,N_663);
or U733 (N_733,N_678,N_661);
nand U734 (N_734,N_687,N_680);
or U735 (N_735,N_697,N_655);
or U736 (N_736,N_679,N_690);
nand U737 (N_737,N_656,N_658);
nor U738 (N_738,N_666,N_698);
nor U739 (N_739,N_656,N_659);
or U740 (N_740,N_674,N_665);
nand U741 (N_741,N_667,N_657);
or U742 (N_742,N_684,N_656);
nor U743 (N_743,N_679,N_660);
and U744 (N_744,N_653,N_651);
or U745 (N_745,N_672,N_662);
and U746 (N_746,N_665,N_672);
nor U747 (N_747,N_662,N_651);
or U748 (N_748,N_659,N_668);
and U749 (N_749,N_669,N_670);
and U750 (N_750,N_715,N_719);
or U751 (N_751,N_705,N_743);
or U752 (N_752,N_708,N_704);
nand U753 (N_753,N_732,N_726);
and U754 (N_754,N_748,N_728);
nor U755 (N_755,N_747,N_700);
nor U756 (N_756,N_742,N_731);
and U757 (N_757,N_744,N_717);
and U758 (N_758,N_723,N_701);
nand U759 (N_759,N_736,N_734);
nor U760 (N_760,N_725,N_724);
and U761 (N_761,N_720,N_718);
nand U762 (N_762,N_714,N_707);
nor U763 (N_763,N_721,N_702);
nor U764 (N_764,N_740,N_722);
and U765 (N_765,N_727,N_730);
or U766 (N_766,N_709,N_733);
or U767 (N_767,N_735,N_746);
xor U768 (N_768,N_711,N_741);
and U769 (N_769,N_712,N_739);
and U770 (N_770,N_713,N_716);
or U771 (N_771,N_729,N_703);
xnor U772 (N_772,N_710,N_706);
or U773 (N_773,N_737,N_738);
or U774 (N_774,N_745,N_749);
nand U775 (N_775,N_732,N_728);
and U776 (N_776,N_704,N_700);
or U777 (N_777,N_703,N_716);
nor U778 (N_778,N_739,N_735);
nor U779 (N_779,N_737,N_718);
nand U780 (N_780,N_729,N_722);
and U781 (N_781,N_732,N_721);
or U782 (N_782,N_732,N_747);
nor U783 (N_783,N_743,N_701);
or U784 (N_784,N_735,N_713);
or U785 (N_785,N_717,N_722);
nand U786 (N_786,N_724,N_720);
nor U787 (N_787,N_716,N_704);
nor U788 (N_788,N_710,N_726);
or U789 (N_789,N_747,N_726);
or U790 (N_790,N_701,N_748);
nand U791 (N_791,N_700,N_735);
or U792 (N_792,N_748,N_718);
or U793 (N_793,N_707,N_718);
nand U794 (N_794,N_729,N_716);
or U795 (N_795,N_746,N_703);
nand U796 (N_796,N_725,N_715);
nor U797 (N_797,N_730,N_719);
xor U798 (N_798,N_744,N_707);
nor U799 (N_799,N_720,N_748);
or U800 (N_800,N_798,N_756);
nand U801 (N_801,N_754,N_774);
or U802 (N_802,N_790,N_773);
and U803 (N_803,N_799,N_751);
nor U804 (N_804,N_796,N_784);
nand U805 (N_805,N_775,N_763);
and U806 (N_806,N_779,N_788);
nand U807 (N_807,N_759,N_757);
nor U808 (N_808,N_753,N_791);
nand U809 (N_809,N_766,N_772);
and U810 (N_810,N_797,N_762);
nand U811 (N_811,N_769,N_783);
nor U812 (N_812,N_777,N_782);
or U813 (N_813,N_760,N_764);
and U814 (N_814,N_770,N_761);
and U815 (N_815,N_767,N_758);
nand U816 (N_816,N_750,N_752);
and U817 (N_817,N_778,N_776);
and U818 (N_818,N_793,N_795);
and U819 (N_819,N_781,N_786);
nor U820 (N_820,N_780,N_765);
nor U821 (N_821,N_792,N_768);
nand U822 (N_822,N_785,N_755);
and U823 (N_823,N_794,N_789);
nor U824 (N_824,N_771,N_787);
or U825 (N_825,N_775,N_759);
nor U826 (N_826,N_799,N_769);
nor U827 (N_827,N_786,N_793);
or U828 (N_828,N_755,N_777);
or U829 (N_829,N_791,N_798);
and U830 (N_830,N_778,N_762);
nand U831 (N_831,N_760,N_770);
or U832 (N_832,N_759,N_755);
and U833 (N_833,N_756,N_772);
nand U834 (N_834,N_776,N_785);
nor U835 (N_835,N_767,N_786);
and U836 (N_836,N_770,N_753);
nor U837 (N_837,N_760,N_781);
nand U838 (N_838,N_791,N_788);
or U839 (N_839,N_757,N_762);
nor U840 (N_840,N_769,N_784);
nor U841 (N_841,N_758,N_786);
or U842 (N_842,N_751,N_794);
or U843 (N_843,N_789,N_797);
or U844 (N_844,N_758,N_761);
nor U845 (N_845,N_770,N_793);
and U846 (N_846,N_762,N_789);
nand U847 (N_847,N_767,N_793);
and U848 (N_848,N_779,N_756);
and U849 (N_849,N_796,N_774);
or U850 (N_850,N_807,N_806);
and U851 (N_851,N_805,N_803);
and U852 (N_852,N_835,N_824);
and U853 (N_853,N_844,N_831);
or U854 (N_854,N_812,N_817);
and U855 (N_855,N_818,N_839);
nor U856 (N_856,N_816,N_825);
and U857 (N_857,N_810,N_800);
and U858 (N_858,N_801,N_841);
and U859 (N_859,N_809,N_813);
nand U860 (N_860,N_820,N_832);
and U861 (N_861,N_834,N_804);
nor U862 (N_862,N_829,N_827);
and U863 (N_863,N_837,N_849);
nor U864 (N_864,N_814,N_833);
and U865 (N_865,N_815,N_846);
nor U866 (N_866,N_808,N_840);
and U867 (N_867,N_819,N_838);
nand U868 (N_868,N_811,N_836);
nor U869 (N_869,N_842,N_830);
nand U870 (N_870,N_843,N_821);
nor U871 (N_871,N_822,N_845);
nand U872 (N_872,N_828,N_848);
nand U873 (N_873,N_826,N_823);
nand U874 (N_874,N_847,N_802);
or U875 (N_875,N_820,N_818);
nor U876 (N_876,N_805,N_834);
nand U877 (N_877,N_835,N_833);
nand U878 (N_878,N_800,N_841);
and U879 (N_879,N_812,N_844);
nor U880 (N_880,N_812,N_806);
or U881 (N_881,N_803,N_832);
nor U882 (N_882,N_809,N_817);
nor U883 (N_883,N_840,N_842);
nor U884 (N_884,N_840,N_807);
nand U885 (N_885,N_822,N_829);
nor U886 (N_886,N_833,N_827);
or U887 (N_887,N_828,N_815);
and U888 (N_888,N_805,N_814);
or U889 (N_889,N_801,N_846);
nand U890 (N_890,N_821,N_844);
and U891 (N_891,N_802,N_825);
nand U892 (N_892,N_815,N_849);
and U893 (N_893,N_818,N_801);
and U894 (N_894,N_802,N_816);
nor U895 (N_895,N_803,N_828);
and U896 (N_896,N_806,N_814);
and U897 (N_897,N_849,N_825);
and U898 (N_898,N_810,N_847);
and U899 (N_899,N_811,N_810);
and U900 (N_900,N_854,N_891);
or U901 (N_901,N_857,N_862);
xnor U902 (N_902,N_851,N_896);
nor U903 (N_903,N_886,N_898);
or U904 (N_904,N_885,N_882);
nor U905 (N_905,N_850,N_888);
and U906 (N_906,N_893,N_859);
and U907 (N_907,N_863,N_892);
or U908 (N_908,N_884,N_856);
or U909 (N_909,N_880,N_897);
or U910 (N_910,N_861,N_858);
and U911 (N_911,N_887,N_879);
and U912 (N_912,N_878,N_871);
nor U913 (N_913,N_873,N_899);
and U914 (N_914,N_868,N_864);
or U915 (N_915,N_874,N_875);
or U916 (N_916,N_852,N_872);
or U917 (N_917,N_894,N_867);
or U918 (N_918,N_870,N_877);
and U919 (N_919,N_860,N_890);
and U920 (N_920,N_876,N_853);
nand U921 (N_921,N_881,N_889);
nand U922 (N_922,N_865,N_855);
and U923 (N_923,N_883,N_866);
or U924 (N_924,N_869,N_895);
nand U925 (N_925,N_875,N_856);
nand U926 (N_926,N_896,N_861);
nor U927 (N_927,N_895,N_889);
and U928 (N_928,N_879,N_880);
or U929 (N_929,N_871,N_851);
nand U930 (N_930,N_893,N_888);
nand U931 (N_931,N_889,N_890);
or U932 (N_932,N_875,N_868);
nand U933 (N_933,N_879,N_876);
and U934 (N_934,N_895,N_882);
and U935 (N_935,N_850,N_862);
nor U936 (N_936,N_894,N_893);
and U937 (N_937,N_879,N_861);
or U938 (N_938,N_888,N_856);
or U939 (N_939,N_858,N_863);
nor U940 (N_940,N_884,N_878);
and U941 (N_941,N_852,N_889);
nand U942 (N_942,N_872,N_886);
nor U943 (N_943,N_866,N_893);
nor U944 (N_944,N_864,N_897);
xor U945 (N_945,N_898,N_895);
and U946 (N_946,N_899,N_877);
and U947 (N_947,N_883,N_857);
nor U948 (N_948,N_885,N_884);
nor U949 (N_949,N_872,N_875);
and U950 (N_950,N_909,N_916);
and U951 (N_951,N_901,N_920);
nand U952 (N_952,N_915,N_935);
nor U953 (N_953,N_911,N_926);
nand U954 (N_954,N_934,N_902);
and U955 (N_955,N_943,N_927);
or U956 (N_956,N_900,N_925);
and U957 (N_957,N_914,N_905);
or U958 (N_958,N_907,N_918);
or U959 (N_959,N_903,N_908);
nand U960 (N_960,N_942,N_919);
nand U961 (N_961,N_941,N_922);
nand U962 (N_962,N_937,N_944);
and U963 (N_963,N_923,N_945);
or U964 (N_964,N_906,N_912);
or U965 (N_965,N_930,N_921);
and U966 (N_966,N_946,N_924);
nand U967 (N_967,N_917,N_939);
nor U968 (N_968,N_932,N_929);
and U969 (N_969,N_938,N_933);
and U970 (N_970,N_913,N_948);
or U971 (N_971,N_940,N_910);
and U972 (N_972,N_904,N_947);
and U973 (N_973,N_949,N_931);
or U974 (N_974,N_928,N_936);
nor U975 (N_975,N_948,N_918);
or U976 (N_976,N_945,N_906);
nor U977 (N_977,N_905,N_922);
nor U978 (N_978,N_945,N_922);
or U979 (N_979,N_927,N_900);
and U980 (N_980,N_948,N_947);
nor U981 (N_981,N_941,N_900);
nor U982 (N_982,N_904,N_913);
nor U983 (N_983,N_926,N_923);
and U984 (N_984,N_945,N_936);
nand U985 (N_985,N_934,N_929);
and U986 (N_986,N_928,N_916);
nand U987 (N_987,N_933,N_914);
nand U988 (N_988,N_914,N_904);
and U989 (N_989,N_920,N_925);
and U990 (N_990,N_921,N_925);
or U991 (N_991,N_903,N_912);
or U992 (N_992,N_921,N_940);
nor U993 (N_993,N_923,N_900);
or U994 (N_994,N_922,N_909);
or U995 (N_995,N_908,N_946);
nand U996 (N_996,N_914,N_907);
or U997 (N_997,N_940,N_949);
and U998 (N_998,N_901,N_908);
or U999 (N_999,N_927,N_914);
nor U1000 (N_1000,N_995,N_954);
or U1001 (N_1001,N_996,N_980);
nand U1002 (N_1002,N_976,N_971);
nor U1003 (N_1003,N_950,N_990);
nand U1004 (N_1004,N_960,N_970);
nand U1005 (N_1005,N_987,N_968);
nor U1006 (N_1006,N_963,N_994);
nor U1007 (N_1007,N_955,N_964);
nor U1008 (N_1008,N_974,N_959);
and U1009 (N_1009,N_975,N_969);
nand U1010 (N_1010,N_951,N_956);
nor U1011 (N_1011,N_984,N_966);
or U1012 (N_1012,N_973,N_988);
nand U1013 (N_1013,N_991,N_962);
and U1014 (N_1014,N_972,N_979);
nand U1015 (N_1015,N_997,N_967);
nor U1016 (N_1016,N_953,N_989);
nor U1017 (N_1017,N_965,N_981);
or U1018 (N_1018,N_999,N_958);
nor U1019 (N_1019,N_986,N_998);
nor U1020 (N_1020,N_992,N_982);
nor U1021 (N_1021,N_983,N_961);
or U1022 (N_1022,N_977,N_952);
nand U1023 (N_1023,N_993,N_957);
nor U1024 (N_1024,N_985,N_978);
or U1025 (N_1025,N_974,N_982);
nor U1026 (N_1026,N_981,N_967);
nor U1027 (N_1027,N_980,N_961);
nand U1028 (N_1028,N_983,N_976);
and U1029 (N_1029,N_999,N_989);
and U1030 (N_1030,N_962,N_978);
and U1031 (N_1031,N_952,N_955);
nor U1032 (N_1032,N_978,N_997);
nand U1033 (N_1033,N_971,N_969);
and U1034 (N_1034,N_997,N_950);
nand U1035 (N_1035,N_976,N_956);
or U1036 (N_1036,N_963,N_959);
and U1037 (N_1037,N_979,N_995);
and U1038 (N_1038,N_962,N_959);
nand U1039 (N_1039,N_979,N_965);
or U1040 (N_1040,N_998,N_967);
nor U1041 (N_1041,N_973,N_990);
nand U1042 (N_1042,N_992,N_966);
nor U1043 (N_1043,N_963,N_989);
nand U1044 (N_1044,N_966,N_955);
nand U1045 (N_1045,N_954,N_955);
nand U1046 (N_1046,N_966,N_976);
or U1047 (N_1047,N_976,N_980);
or U1048 (N_1048,N_953,N_950);
nor U1049 (N_1049,N_989,N_977);
or U1050 (N_1050,N_1013,N_1036);
or U1051 (N_1051,N_1038,N_1039);
nor U1052 (N_1052,N_1028,N_1035);
nor U1053 (N_1053,N_1045,N_1009);
nand U1054 (N_1054,N_1021,N_1034);
nand U1055 (N_1055,N_1043,N_1000);
or U1056 (N_1056,N_1026,N_1031);
and U1057 (N_1057,N_1006,N_1010);
nor U1058 (N_1058,N_1001,N_1046);
or U1059 (N_1059,N_1004,N_1012);
nand U1060 (N_1060,N_1044,N_1023);
nand U1061 (N_1061,N_1015,N_1033);
nand U1062 (N_1062,N_1011,N_1027);
or U1063 (N_1063,N_1020,N_1014);
nand U1064 (N_1064,N_1017,N_1007);
nand U1065 (N_1065,N_1019,N_1016);
and U1066 (N_1066,N_1032,N_1041);
nor U1067 (N_1067,N_1002,N_1037);
xor U1068 (N_1068,N_1049,N_1025);
nand U1069 (N_1069,N_1005,N_1018);
or U1070 (N_1070,N_1047,N_1008);
nand U1071 (N_1071,N_1029,N_1040);
nand U1072 (N_1072,N_1003,N_1030);
or U1073 (N_1073,N_1042,N_1022);
and U1074 (N_1074,N_1024,N_1048);
or U1075 (N_1075,N_1028,N_1033);
or U1076 (N_1076,N_1030,N_1031);
and U1077 (N_1077,N_1033,N_1021);
nand U1078 (N_1078,N_1038,N_1005);
nor U1079 (N_1079,N_1031,N_1015);
nand U1080 (N_1080,N_1017,N_1016);
nand U1081 (N_1081,N_1026,N_1010);
nor U1082 (N_1082,N_1041,N_1049);
nand U1083 (N_1083,N_1012,N_1044);
nor U1084 (N_1084,N_1028,N_1037);
nor U1085 (N_1085,N_1018,N_1035);
or U1086 (N_1086,N_1006,N_1029);
nor U1087 (N_1087,N_1042,N_1033);
or U1088 (N_1088,N_1007,N_1044);
nor U1089 (N_1089,N_1002,N_1029);
nor U1090 (N_1090,N_1012,N_1036);
and U1091 (N_1091,N_1044,N_1009);
and U1092 (N_1092,N_1002,N_1024);
and U1093 (N_1093,N_1045,N_1013);
nand U1094 (N_1094,N_1016,N_1015);
or U1095 (N_1095,N_1039,N_1011);
or U1096 (N_1096,N_1043,N_1016);
nor U1097 (N_1097,N_1036,N_1044);
nor U1098 (N_1098,N_1043,N_1041);
nor U1099 (N_1099,N_1049,N_1031);
or U1100 (N_1100,N_1085,N_1079);
and U1101 (N_1101,N_1073,N_1090);
nand U1102 (N_1102,N_1087,N_1069);
xor U1103 (N_1103,N_1076,N_1063);
nand U1104 (N_1104,N_1050,N_1061);
and U1105 (N_1105,N_1093,N_1088);
nor U1106 (N_1106,N_1099,N_1089);
and U1107 (N_1107,N_1097,N_1059);
and U1108 (N_1108,N_1064,N_1078);
nand U1109 (N_1109,N_1056,N_1057);
nor U1110 (N_1110,N_1054,N_1081);
nand U1111 (N_1111,N_1068,N_1082);
or U1112 (N_1112,N_1075,N_1074);
nor U1113 (N_1113,N_1072,N_1053);
or U1114 (N_1114,N_1066,N_1080);
nor U1115 (N_1115,N_1077,N_1084);
or U1116 (N_1116,N_1071,N_1060);
nand U1117 (N_1117,N_1051,N_1091);
or U1118 (N_1118,N_1067,N_1058);
and U1119 (N_1119,N_1070,N_1098);
nor U1120 (N_1120,N_1062,N_1086);
nor U1121 (N_1121,N_1095,N_1083);
nand U1122 (N_1122,N_1092,N_1052);
nand U1123 (N_1123,N_1055,N_1065);
and U1124 (N_1124,N_1094,N_1096);
or U1125 (N_1125,N_1077,N_1080);
nand U1126 (N_1126,N_1081,N_1071);
and U1127 (N_1127,N_1092,N_1088);
and U1128 (N_1128,N_1075,N_1087);
nor U1129 (N_1129,N_1059,N_1088);
nor U1130 (N_1130,N_1072,N_1063);
or U1131 (N_1131,N_1094,N_1077);
or U1132 (N_1132,N_1054,N_1091);
and U1133 (N_1133,N_1062,N_1055);
nor U1134 (N_1134,N_1074,N_1087);
and U1135 (N_1135,N_1095,N_1062);
and U1136 (N_1136,N_1077,N_1064);
or U1137 (N_1137,N_1055,N_1053);
nand U1138 (N_1138,N_1098,N_1061);
or U1139 (N_1139,N_1069,N_1054);
and U1140 (N_1140,N_1096,N_1060);
nor U1141 (N_1141,N_1083,N_1075);
or U1142 (N_1142,N_1099,N_1080);
or U1143 (N_1143,N_1094,N_1067);
or U1144 (N_1144,N_1059,N_1077);
and U1145 (N_1145,N_1058,N_1086);
nor U1146 (N_1146,N_1054,N_1072);
nor U1147 (N_1147,N_1075,N_1095);
or U1148 (N_1148,N_1073,N_1084);
and U1149 (N_1149,N_1067,N_1096);
nor U1150 (N_1150,N_1123,N_1103);
nand U1151 (N_1151,N_1130,N_1133);
and U1152 (N_1152,N_1134,N_1127);
nor U1153 (N_1153,N_1139,N_1114);
and U1154 (N_1154,N_1104,N_1138);
nand U1155 (N_1155,N_1118,N_1107);
or U1156 (N_1156,N_1129,N_1105);
nor U1157 (N_1157,N_1111,N_1115);
nand U1158 (N_1158,N_1116,N_1121);
or U1159 (N_1159,N_1148,N_1110);
or U1160 (N_1160,N_1146,N_1113);
nor U1161 (N_1161,N_1137,N_1119);
and U1162 (N_1162,N_1135,N_1101);
and U1163 (N_1163,N_1108,N_1100);
nand U1164 (N_1164,N_1131,N_1147);
or U1165 (N_1165,N_1141,N_1125);
nand U1166 (N_1166,N_1109,N_1145);
or U1167 (N_1167,N_1120,N_1143);
nor U1168 (N_1168,N_1132,N_1126);
or U1169 (N_1169,N_1106,N_1136);
nand U1170 (N_1170,N_1149,N_1112);
or U1171 (N_1171,N_1122,N_1124);
nand U1172 (N_1172,N_1140,N_1142);
nor U1173 (N_1173,N_1128,N_1144);
nor U1174 (N_1174,N_1102,N_1117);
nor U1175 (N_1175,N_1149,N_1102);
nand U1176 (N_1176,N_1112,N_1145);
or U1177 (N_1177,N_1146,N_1131);
nor U1178 (N_1178,N_1103,N_1102);
and U1179 (N_1179,N_1130,N_1134);
nand U1180 (N_1180,N_1124,N_1140);
and U1181 (N_1181,N_1132,N_1106);
or U1182 (N_1182,N_1102,N_1115);
and U1183 (N_1183,N_1139,N_1106);
or U1184 (N_1184,N_1103,N_1132);
nor U1185 (N_1185,N_1115,N_1124);
and U1186 (N_1186,N_1149,N_1134);
nor U1187 (N_1187,N_1143,N_1116);
and U1188 (N_1188,N_1112,N_1128);
nor U1189 (N_1189,N_1131,N_1128);
or U1190 (N_1190,N_1108,N_1147);
nand U1191 (N_1191,N_1108,N_1146);
nor U1192 (N_1192,N_1130,N_1122);
nand U1193 (N_1193,N_1114,N_1122);
nand U1194 (N_1194,N_1137,N_1124);
nand U1195 (N_1195,N_1101,N_1104);
nor U1196 (N_1196,N_1115,N_1141);
nand U1197 (N_1197,N_1121,N_1137);
nand U1198 (N_1198,N_1144,N_1138);
nor U1199 (N_1199,N_1146,N_1102);
nor U1200 (N_1200,N_1180,N_1172);
nor U1201 (N_1201,N_1197,N_1165);
and U1202 (N_1202,N_1156,N_1161);
nor U1203 (N_1203,N_1153,N_1193);
nand U1204 (N_1204,N_1168,N_1150);
nor U1205 (N_1205,N_1155,N_1175);
xnor U1206 (N_1206,N_1179,N_1159);
and U1207 (N_1207,N_1171,N_1158);
and U1208 (N_1208,N_1160,N_1181);
nor U1209 (N_1209,N_1162,N_1188);
nor U1210 (N_1210,N_1189,N_1170);
xnor U1211 (N_1211,N_1191,N_1176);
nand U1212 (N_1212,N_1183,N_1190);
nor U1213 (N_1213,N_1195,N_1182);
and U1214 (N_1214,N_1174,N_1199);
and U1215 (N_1215,N_1157,N_1187);
nand U1216 (N_1216,N_1152,N_1167);
xnor U1217 (N_1217,N_1186,N_1184);
and U1218 (N_1218,N_1192,N_1177);
nand U1219 (N_1219,N_1196,N_1169);
nor U1220 (N_1220,N_1166,N_1163);
or U1221 (N_1221,N_1173,N_1194);
or U1222 (N_1222,N_1154,N_1198);
nand U1223 (N_1223,N_1151,N_1164);
and U1224 (N_1224,N_1178,N_1185);
or U1225 (N_1225,N_1195,N_1167);
nand U1226 (N_1226,N_1189,N_1179);
nor U1227 (N_1227,N_1164,N_1170);
or U1228 (N_1228,N_1191,N_1153);
nor U1229 (N_1229,N_1195,N_1172);
or U1230 (N_1230,N_1178,N_1176);
nor U1231 (N_1231,N_1171,N_1176);
or U1232 (N_1232,N_1198,N_1177);
nand U1233 (N_1233,N_1187,N_1151);
nand U1234 (N_1234,N_1184,N_1187);
nand U1235 (N_1235,N_1156,N_1150);
and U1236 (N_1236,N_1196,N_1172);
nand U1237 (N_1237,N_1194,N_1191);
and U1238 (N_1238,N_1161,N_1196);
or U1239 (N_1239,N_1156,N_1171);
and U1240 (N_1240,N_1167,N_1176);
and U1241 (N_1241,N_1198,N_1161);
and U1242 (N_1242,N_1186,N_1155);
nand U1243 (N_1243,N_1165,N_1163);
or U1244 (N_1244,N_1165,N_1194);
and U1245 (N_1245,N_1150,N_1167);
nor U1246 (N_1246,N_1188,N_1150);
nor U1247 (N_1247,N_1188,N_1171);
and U1248 (N_1248,N_1177,N_1159);
xnor U1249 (N_1249,N_1188,N_1168);
or U1250 (N_1250,N_1248,N_1242);
nand U1251 (N_1251,N_1226,N_1236);
or U1252 (N_1252,N_1206,N_1214);
nor U1253 (N_1253,N_1241,N_1239);
or U1254 (N_1254,N_1213,N_1220);
nand U1255 (N_1255,N_1212,N_1208);
or U1256 (N_1256,N_1218,N_1221);
or U1257 (N_1257,N_1205,N_1233);
nand U1258 (N_1258,N_1202,N_1222);
or U1259 (N_1259,N_1216,N_1201);
or U1260 (N_1260,N_1234,N_1244);
nand U1261 (N_1261,N_1215,N_1231);
or U1262 (N_1262,N_1217,N_1227);
or U1263 (N_1263,N_1228,N_1243);
or U1264 (N_1264,N_1230,N_1210);
nor U1265 (N_1265,N_1249,N_1240);
or U1266 (N_1266,N_1209,N_1235);
and U1267 (N_1267,N_1245,N_1203);
nor U1268 (N_1268,N_1229,N_1211);
nand U1269 (N_1269,N_1207,N_1224);
nor U1270 (N_1270,N_1232,N_1247);
nand U1271 (N_1271,N_1223,N_1204);
nor U1272 (N_1272,N_1246,N_1238);
and U1273 (N_1273,N_1225,N_1219);
or U1274 (N_1274,N_1237,N_1200);
or U1275 (N_1275,N_1228,N_1220);
nand U1276 (N_1276,N_1213,N_1210);
and U1277 (N_1277,N_1232,N_1211);
nor U1278 (N_1278,N_1216,N_1247);
and U1279 (N_1279,N_1242,N_1209);
and U1280 (N_1280,N_1202,N_1235);
nor U1281 (N_1281,N_1230,N_1213);
nor U1282 (N_1282,N_1201,N_1243);
nand U1283 (N_1283,N_1237,N_1216);
or U1284 (N_1284,N_1242,N_1218);
nand U1285 (N_1285,N_1207,N_1249);
nor U1286 (N_1286,N_1207,N_1237);
nor U1287 (N_1287,N_1223,N_1236);
and U1288 (N_1288,N_1246,N_1222);
nand U1289 (N_1289,N_1241,N_1249);
nand U1290 (N_1290,N_1231,N_1226);
and U1291 (N_1291,N_1205,N_1240);
and U1292 (N_1292,N_1204,N_1241);
and U1293 (N_1293,N_1230,N_1207);
or U1294 (N_1294,N_1211,N_1228);
and U1295 (N_1295,N_1206,N_1203);
nand U1296 (N_1296,N_1218,N_1207);
nand U1297 (N_1297,N_1212,N_1215);
nand U1298 (N_1298,N_1200,N_1244);
or U1299 (N_1299,N_1201,N_1232);
and U1300 (N_1300,N_1258,N_1284);
nor U1301 (N_1301,N_1272,N_1288);
xor U1302 (N_1302,N_1292,N_1295);
nand U1303 (N_1303,N_1260,N_1294);
nand U1304 (N_1304,N_1255,N_1265);
nand U1305 (N_1305,N_1285,N_1250);
and U1306 (N_1306,N_1263,N_1261);
nor U1307 (N_1307,N_1290,N_1270);
nand U1308 (N_1308,N_1256,N_1286);
nor U1309 (N_1309,N_1271,N_1276);
and U1310 (N_1310,N_1253,N_1297);
xor U1311 (N_1311,N_1283,N_1298);
and U1312 (N_1312,N_1264,N_1282);
or U1313 (N_1313,N_1277,N_1279);
and U1314 (N_1314,N_1281,N_1269);
nor U1315 (N_1315,N_1287,N_1257);
or U1316 (N_1316,N_1268,N_1278);
nand U1317 (N_1317,N_1293,N_1251);
and U1318 (N_1318,N_1291,N_1267);
and U1319 (N_1319,N_1299,N_1296);
or U1320 (N_1320,N_1274,N_1280);
or U1321 (N_1321,N_1262,N_1289);
nand U1322 (N_1322,N_1259,N_1275);
and U1323 (N_1323,N_1273,N_1254);
and U1324 (N_1324,N_1266,N_1252);
nand U1325 (N_1325,N_1278,N_1265);
and U1326 (N_1326,N_1291,N_1283);
nand U1327 (N_1327,N_1283,N_1261);
nand U1328 (N_1328,N_1271,N_1275);
nor U1329 (N_1329,N_1252,N_1291);
and U1330 (N_1330,N_1289,N_1263);
or U1331 (N_1331,N_1286,N_1255);
or U1332 (N_1332,N_1265,N_1277);
or U1333 (N_1333,N_1260,N_1258);
nor U1334 (N_1334,N_1272,N_1287);
nor U1335 (N_1335,N_1279,N_1255);
nand U1336 (N_1336,N_1284,N_1281);
and U1337 (N_1337,N_1274,N_1285);
and U1338 (N_1338,N_1274,N_1296);
or U1339 (N_1339,N_1266,N_1268);
and U1340 (N_1340,N_1280,N_1268);
nor U1341 (N_1341,N_1277,N_1258);
nand U1342 (N_1342,N_1284,N_1294);
and U1343 (N_1343,N_1251,N_1288);
or U1344 (N_1344,N_1293,N_1261);
or U1345 (N_1345,N_1299,N_1285);
nor U1346 (N_1346,N_1251,N_1265);
nor U1347 (N_1347,N_1250,N_1275);
or U1348 (N_1348,N_1257,N_1278);
nand U1349 (N_1349,N_1254,N_1286);
or U1350 (N_1350,N_1332,N_1340);
nand U1351 (N_1351,N_1345,N_1306);
and U1352 (N_1352,N_1325,N_1304);
nand U1353 (N_1353,N_1323,N_1337);
nor U1354 (N_1354,N_1320,N_1348);
nor U1355 (N_1355,N_1305,N_1335);
nor U1356 (N_1356,N_1342,N_1317);
or U1357 (N_1357,N_1327,N_1338);
xor U1358 (N_1358,N_1310,N_1349);
or U1359 (N_1359,N_1334,N_1344);
xnor U1360 (N_1360,N_1301,N_1308);
nand U1361 (N_1361,N_1329,N_1322);
nor U1362 (N_1362,N_1302,N_1314);
nand U1363 (N_1363,N_1319,N_1312);
and U1364 (N_1364,N_1316,N_1347);
and U1365 (N_1365,N_1341,N_1307);
nor U1366 (N_1366,N_1321,N_1333);
or U1367 (N_1367,N_1309,N_1346);
and U1368 (N_1368,N_1328,N_1326);
nor U1369 (N_1369,N_1336,N_1331);
and U1370 (N_1370,N_1311,N_1343);
and U1371 (N_1371,N_1339,N_1300);
and U1372 (N_1372,N_1313,N_1318);
and U1373 (N_1373,N_1315,N_1324);
nor U1374 (N_1374,N_1330,N_1303);
nand U1375 (N_1375,N_1307,N_1313);
nand U1376 (N_1376,N_1304,N_1307);
or U1377 (N_1377,N_1303,N_1318);
and U1378 (N_1378,N_1328,N_1322);
or U1379 (N_1379,N_1307,N_1340);
and U1380 (N_1380,N_1342,N_1316);
nand U1381 (N_1381,N_1306,N_1342);
and U1382 (N_1382,N_1322,N_1305);
and U1383 (N_1383,N_1338,N_1331);
or U1384 (N_1384,N_1341,N_1318);
or U1385 (N_1385,N_1329,N_1316);
nand U1386 (N_1386,N_1315,N_1317);
nor U1387 (N_1387,N_1341,N_1301);
or U1388 (N_1388,N_1334,N_1316);
or U1389 (N_1389,N_1345,N_1309);
and U1390 (N_1390,N_1304,N_1328);
nor U1391 (N_1391,N_1327,N_1330);
nor U1392 (N_1392,N_1348,N_1335);
and U1393 (N_1393,N_1348,N_1336);
nor U1394 (N_1394,N_1303,N_1339);
nand U1395 (N_1395,N_1303,N_1324);
nor U1396 (N_1396,N_1323,N_1339);
nand U1397 (N_1397,N_1328,N_1303);
xor U1398 (N_1398,N_1337,N_1339);
nand U1399 (N_1399,N_1335,N_1323);
nand U1400 (N_1400,N_1362,N_1376);
nor U1401 (N_1401,N_1350,N_1375);
nand U1402 (N_1402,N_1386,N_1378);
nand U1403 (N_1403,N_1351,N_1389);
nand U1404 (N_1404,N_1356,N_1373);
or U1405 (N_1405,N_1398,N_1397);
nand U1406 (N_1406,N_1391,N_1353);
or U1407 (N_1407,N_1359,N_1394);
or U1408 (N_1408,N_1358,N_1383);
nand U1409 (N_1409,N_1399,N_1361);
nand U1410 (N_1410,N_1372,N_1379);
or U1411 (N_1411,N_1352,N_1382);
or U1412 (N_1412,N_1384,N_1392);
nand U1413 (N_1413,N_1370,N_1390);
or U1414 (N_1414,N_1355,N_1363);
nor U1415 (N_1415,N_1368,N_1360);
or U1416 (N_1416,N_1369,N_1374);
nand U1417 (N_1417,N_1381,N_1377);
nor U1418 (N_1418,N_1371,N_1395);
or U1419 (N_1419,N_1380,N_1364);
and U1420 (N_1420,N_1385,N_1366);
or U1421 (N_1421,N_1367,N_1365);
nand U1422 (N_1422,N_1387,N_1393);
or U1423 (N_1423,N_1396,N_1357);
and U1424 (N_1424,N_1388,N_1354);
nand U1425 (N_1425,N_1376,N_1393);
or U1426 (N_1426,N_1364,N_1369);
nand U1427 (N_1427,N_1397,N_1389);
xnor U1428 (N_1428,N_1369,N_1365);
or U1429 (N_1429,N_1364,N_1366);
or U1430 (N_1430,N_1355,N_1370);
or U1431 (N_1431,N_1358,N_1376);
nor U1432 (N_1432,N_1358,N_1359);
nand U1433 (N_1433,N_1373,N_1394);
or U1434 (N_1434,N_1382,N_1378);
or U1435 (N_1435,N_1370,N_1358);
nand U1436 (N_1436,N_1361,N_1352);
nor U1437 (N_1437,N_1360,N_1379);
nor U1438 (N_1438,N_1350,N_1384);
or U1439 (N_1439,N_1394,N_1367);
and U1440 (N_1440,N_1377,N_1363);
and U1441 (N_1441,N_1396,N_1395);
and U1442 (N_1442,N_1384,N_1353);
or U1443 (N_1443,N_1363,N_1379);
nor U1444 (N_1444,N_1353,N_1398);
nand U1445 (N_1445,N_1364,N_1360);
nor U1446 (N_1446,N_1388,N_1380);
and U1447 (N_1447,N_1383,N_1399);
nor U1448 (N_1448,N_1377,N_1390);
nand U1449 (N_1449,N_1387,N_1375);
xnor U1450 (N_1450,N_1439,N_1401);
nand U1451 (N_1451,N_1410,N_1403);
and U1452 (N_1452,N_1411,N_1427);
nand U1453 (N_1453,N_1443,N_1445);
nor U1454 (N_1454,N_1423,N_1415);
nand U1455 (N_1455,N_1425,N_1446);
or U1456 (N_1456,N_1407,N_1421);
nor U1457 (N_1457,N_1419,N_1412);
and U1458 (N_1458,N_1431,N_1442);
or U1459 (N_1459,N_1440,N_1405);
or U1460 (N_1460,N_1432,N_1417);
nor U1461 (N_1461,N_1429,N_1402);
nand U1462 (N_1462,N_1418,N_1434);
nand U1463 (N_1463,N_1404,N_1400);
nor U1464 (N_1464,N_1424,N_1420);
and U1465 (N_1465,N_1428,N_1409);
or U1466 (N_1466,N_1437,N_1441);
nand U1467 (N_1467,N_1448,N_1438);
or U1468 (N_1468,N_1426,N_1414);
or U1469 (N_1469,N_1435,N_1444);
or U1470 (N_1470,N_1413,N_1422);
or U1471 (N_1471,N_1447,N_1408);
nor U1472 (N_1472,N_1406,N_1436);
nor U1473 (N_1473,N_1430,N_1433);
nand U1474 (N_1474,N_1416,N_1449);
and U1475 (N_1475,N_1433,N_1401);
or U1476 (N_1476,N_1444,N_1415);
and U1477 (N_1477,N_1419,N_1447);
nor U1478 (N_1478,N_1432,N_1431);
and U1479 (N_1479,N_1406,N_1434);
or U1480 (N_1480,N_1406,N_1430);
or U1481 (N_1481,N_1410,N_1412);
and U1482 (N_1482,N_1448,N_1433);
or U1483 (N_1483,N_1421,N_1438);
nand U1484 (N_1484,N_1424,N_1435);
and U1485 (N_1485,N_1442,N_1444);
nand U1486 (N_1486,N_1440,N_1402);
nor U1487 (N_1487,N_1437,N_1426);
nand U1488 (N_1488,N_1414,N_1405);
or U1489 (N_1489,N_1401,N_1403);
and U1490 (N_1490,N_1406,N_1438);
nor U1491 (N_1491,N_1428,N_1419);
nand U1492 (N_1492,N_1441,N_1404);
nand U1493 (N_1493,N_1449,N_1419);
or U1494 (N_1494,N_1430,N_1419);
nor U1495 (N_1495,N_1432,N_1402);
nor U1496 (N_1496,N_1429,N_1433);
or U1497 (N_1497,N_1411,N_1432);
nand U1498 (N_1498,N_1431,N_1438);
and U1499 (N_1499,N_1430,N_1412);
and U1500 (N_1500,N_1494,N_1466);
or U1501 (N_1501,N_1459,N_1474);
and U1502 (N_1502,N_1455,N_1477);
nor U1503 (N_1503,N_1489,N_1483);
and U1504 (N_1504,N_1493,N_1463);
or U1505 (N_1505,N_1464,N_1487);
nor U1506 (N_1506,N_1465,N_1453);
nor U1507 (N_1507,N_1462,N_1499);
or U1508 (N_1508,N_1469,N_1458);
nand U1509 (N_1509,N_1498,N_1486);
nand U1510 (N_1510,N_1456,N_1476);
and U1511 (N_1511,N_1467,N_1480);
nor U1512 (N_1512,N_1479,N_1490);
and U1513 (N_1513,N_1478,N_1482);
and U1514 (N_1514,N_1460,N_1473);
nand U1515 (N_1515,N_1472,N_1475);
nor U1516 (N_1516,N_1497,N_1450);
and U1517 (N_1517,N_1471,N_1468);
nor U1518 (N_1518,N_1451,N_1461);
and U1519 (N_1519,N_1484,N_1481);
nand U1520 (N_1520,N_1496,N_1488);
nand U1521 (N_1521,N_1491,N_1454);
nand U1522 (N_1522,N_1495,N_1457);
nand U1523 (N_1523,N_1492,N_1485);
nor U1524 (N_1524,N_1452,N_1470);
or U1525 (N_1525,N_1463,N_1471);
or U1526 (N_1526,N_1496,N_1481);
and U1527 (N_1527,N_1451,N_1459);
nor U1528 (N_1528,N_1466,N_1486);
nor U1529 (N_1529,N_1450,N_1453);
nor U1530 (N_1530,N_1454,N_1481);
nor U1531 (N_1531,N_1477,N_1454);
nor U1532 (N_1532,N_1467,N_1469);
nand U1533 (N_1533,N_1486,N_1453);
nor U1534 (N_1534,N_1474,N_1470);
and U1535 (N_1535,N_1469,N_1471);
nand U1536 (N_1536,N_1487,N_1456);
nor U1537 (N_1537,N_1492,N_1469);
and U1538 (N_1538,N_1494,N_1468);
nor U1539 (N_1539,N_1476,N_1499);
or U1540 (N_1540,N_1490,N_1481);
nor U1541 (N_1541,N_1468,N_1491);
nor U1542 (N_1542,N_1483,N_1454);
or U1543 (N_1543,N_1494,N_1489);
or U1544 (N_1544,N_1481,N_1474);
or U1545 (N_1545,N_1489,N_1473);
or U1546 (N_1546,N_1477,N_1472);
nor U1547 (N_1547,N_1495,N_1478);
xor U1548 (N_1548,N_1478,N_1450);
or U1549 (N_1549,N_1496,N_1499);
nand U1550 (N_1550,N_1515,N_1536);
nand U1551 (N_1551,N_1514,N_1531);
or U1552 (N_1552,N_1507,N_1539);
nand U1553 (N_1553,N_1524,N_1504);
or U1554 (N_1554,N_1525,N_1521);
and U1555 (N_1555,N_1519,N_1543);
nor U1556 (N_1556,N_1510,N_1532);
and U1557 (N_1557,N_1542,N_1506);
nor U1558 (N_1558,N_1503,N_1546);
or U1559 (N_1559,N_1520,N_1501);
or U1560 (N_1560,N_1540,N_1513);
and U1561 (N_1561,N_1508,N_1527);
and U1562 (N_1562,N_1511,N_1541);
nor U1563 (N_1563,N_1535,N_1516);
or U1564 (N_1564,N_1534,N_1522);
or U1565 (N_1565,N_1545,N_1505);
nand U1566 (N_1566,N_1526,N_1517);
and U1567 (N_1567,N_1537,N_1548);
or U1568 (N_1568,N_1538,N_1533);
nand U1569 (N_1569,N_1547,N_1502);
nand U1570 (N_1570,N_1500,N_1523);
and U1571 (N_1571,N_1549,N_1509);
nor U1572 (N_1572,N_1512,N_1529);
nor U1573 (N_1573,N_1518,N_1530);
nor U1574 (N_1574,N_1544,N_1528);
and U1575 (N_1575,N_1504,N_1543);
and U1576 (N_1576,N_1522,N_1523);
and U1577 (N_1577,N_1518,N_1545);
nor U1578 (N_1578,N_1500,N_1527);
or U1579 (N_1579,N_1514,N_1526);
or U1580 (N_1580,N_1529,N_1525);
nor U1581 (N_1581,N_1528,N_1532);
and U1582 (N_1582,N_1513,N_1524);
nand U1583 (N_1583,N_1513,N_1512);
nor U1584 (N_1584,N_1533,N_1509);
and U1585 (N_1585,N_1502,N_1529);
nand U1586 (N_1586,N_1526,N_1522);
nand U1587 (N_1587,N_1538,N_1536);
and U1588 (N_1588,N_1501,N_1546);
nand U1589 (N_1589,N_1530,N_1539);
or U1590 (N_1590,N_1519,N_1506);
nor U1591 (N_1591,N_1530,N_1525);
and U1592 (N_1592,N_1517,N_1523);
nand U1593 (N_1593,N_1507,N_1532);
nand U1594 (N_1594,N_1522,N_1515);
nor U1595 (N_1595,N_1502,N_1518);
nand U1596 (N_1596,N_1509,N_1526);
nand U1597 (N_1597,N_1514,N_1506);
nand U1598 (N_1598,N_1503,N_1523);
and U1599 (N_1599,N_1510,N_1536);
and U1600 (N_1600,N_1570,N_1565);
nor U1601 (N_1601,N_1592,N_1584);
and U1602 (N_1602,N_1596,N_1585);
nand U1603 (N_1603,N_1593,N_1589);
and U1604 (N_1604,N_1590,N_1598);
xnor U1605 (N_1605,N_1551,N_1552);
or U1606 (N_1606,N_1556,N_1564);
and U1607 (N_1607,N_1597,N_1574);
nor U1608 (N_1608,N_1571,N_1569);
nand U1609 (N_1609,N_1583,N_1587);
nand U1610 (N_1610,N_1554,N_1560);
or U1611 (N_1611,N_1563,N_1591);
nand U1612 (N_1612,N_1557,N_1553);
nand U1613 (N_1613,N_1575,N_1572);
and U1614 (N_1614,N_1588,N_1580);
and U1615 (N_1615,N_1579,N_1599);
or U1616 (N_1616,N_1582,N_1566);
nand U1617 (N_1617,N_1568,N_1594);
or U1618 (N_1618,N_1562,N_1559);
or U1619 (N_1619,N_1576,N_1581);
and U1620 (N_1620,N_1586,N_1558);
nor U1621 (N_1621,N_1573,N_1561);
nand U1622 (N_1622,N_1578,N_1577);
or U1623 (N_1623,N_1595,N_1555);
or U1624 (N_1624,N_1567,N_1550);
and U1625 (N_1625,N_1595,N_1588);
nand U1626 (N_1626,N_1592,N_1560);
nor U1627 (N_1627,N_1575,N_1585);
nand U1628 (N_1628,N_1582,N_1556);
and U1629 (N_1629,N_1581,N_1597);
or U1630 (N_1630,N_1572,N_1592);
and U1631 (N_1631,N_1586,N_1583);
nor U1632 (N_1632,N_1572,N_1561);
nor U1633 (N_1633,N_1574,N_1562);
nor U1634 (N_1634,N_1573,N_1584);
nor U1635 (N_1635,N_1593,N_1559);
nor U1636 (N_1636,N_1580,N_1560);
nand U1637 (N_1637,N_1579,N_1596);
and U1638 (N_1638,N_1553,N_1585);
nor U1639 (N_1639,N_1595,N_1550);
nor U1640 (N_1640,N_1596,N_1595);
nor U1641 (N_1641,N_1596,N_1591);
nand U1642 (N_1642,N_1591,N_1597);
or U1643 (N_1643,N_1593,N_1556);
nor U1644 (N_1644,N_1553,N_1592);
and U1645 (N_1645,N_1586,N_1553);
nand U1646 (N_1646,N_1582,N_1565);
and U1647 (N_1647,N_1594,N_1575);
nand U1648 (N_1648,N_1562,N_1592);
nor U1649 (N_1649,N_1565,N_1588);
or U1650 (N_1650,N_1642,N_1647);
nor U1651 (N_1651,N_1620,N_1605);
nand U1652 (N_1652,N_1629,N_1638);
nor U1653 (N_1653,N_1631,N_1607);
and U1654 (N_1654,N_1633,N_1627);
and U1655 (N_1655,N_1635,N_1639);
nor U1656 (N_1656,N_1628,N_1649);
nor U1657 (N_1657,N_1621,N_1637);
nand U1658 (N_1658,N_1624,N_1604);
and U1659 (N_1659,N_1646,N_1600);
and U1660 (N_1660,N_1645,N_1610);
nand U1661 (N_1661,N_1613,N_1616);
nor U1662 (N_1662,N_1612,N_1643);
nand U1663 (N_1663,N_1618,N_1640);
nand U1664 (N_1664,N_1625,N_1644);
or U1665 (N_1665,N_1619,N_1615);
nand U1666 (N_1666,N_1608,N_1632);
xor U1667 (N_1667,N_1609,N_1622);
and U1668 (N_1668,N_1641,N_1626);
nand U1669 (N_1669,N_1630,N_1648);
or U1670 (N_1670,N_1602,N_1606);
nand U1671 (N_1671,N_1617,N_1603);
and U1672 (N_1672,N_1634,N_1614);
and U1673 (N_1673,N_1601,N_1623);
nand U1674 (N_1674,N_1611,N_1636);
and U1675 (N_1675,N_1646,N_1610);
and U1676 (N_1676,N_1632,N_1614);
or U1677 (N_1677,N_1600,N_1639);
or U1678 (N_1678,N_1647,N_1637);
or U1679 (N_1679,N_1610,N_1607);
nand U1680 (N_1680,N_1607,N_1616);
nor U1681 (N_1681,N_1607,N_1629);
nor U1682 (N_1682,N_1628,N_1625);
nor U1683 (N_1683,N_1644,N_1624);
nor U1684 (N_1684,N_1619,N_1649);
nand U1685 (N_1685,N_1619,N_1617);
and U1686 (N_1686,N_1610,N_1611);
and U1687 (N_1687,N_1649,N_1622);
or U1688 (N_1688,N_1607,N_1602);
and U1689 (N_1689,N_1632,N_1603);
nand U1690 (N_1690,N_1625,N_1623);
nor U1691 (N_1691,N_1644,N_1640);
or U1692 (N_1692,N_1638,N_1632);
or U1693 (N_1693,N_1641,N_1627);
nor U1694 (N_1694,N_1607,N_1649);
nor U1695 (N_1695,N_1609,N_1636);
or U1696 (N_1696,N_1644,N_1627);
or U1697 (N_1697,N_1635,N_1633);
nor U1698 (N_1698,N_1613,N_1628);
or U1699 (N_1699,N_1634,N_1627);
xnor U1700 (N_1700,N_1693,N_1676);
and U1701 (N_1701,N_1667,N_1684);
or U1702 (N_1702,N_1655,N_1677);
or U1703 (N_1703,N_1654,N_1696);
and U1704 (N_1704,N_1666,N_1690);
nor U1705 (N_1705,N_1675,N_1672);
nor U1706 (N_1706,N_1664,N_1686);
nor U1707 (N_1707,N_1662,N_1680);
nor U1708 (N_1708,N_1685,N_1658);
xor U1709 (N_1709,N_1678,N_1697);
nor U1710 (N_1710,N_1687,N_1665);
or U1711 (N_1711,N_1695,N_1674);
nor U1712 (N_1712,N_1688,N_1689);
and U1713 (N_1713,N_1650,N_1694);
or U1714 (N_1714,N_1653,N_1652);
and U1715 (N_1715,N_1656,N_1660);
nor U1716 (N_1716,N_1663,N_1698);
nand U1717 (N_1717,N_1657,N_1661);
nor U1718 (N_1718,N_1668,N_1681);
or U1719 (N_1719,N_1671,N_1670);
nand U1720 (N_1720,N_1679,N_1651);
or U1721 (N_1721,N_1683,N_1682);
or U1722 (N_1722,N_1669,N_1673);
nand U1723 (N_1723,N_1691,N_1659);
or U1724 (N_1724,N_1699,N_1692);
and U1725 (N_1725,N_1663,N_1673);
and U1726 (N_1726,N_1692,N_1689);
xor U1727 (N_1727,N_1666,N_1678);
nor U1728 (N_1728,N_1694,N_1670);
and U1729 (N_1729,N_1688,N_1670);
xor U1730 (N_1730,N_1682,N_1674);
nand U1731 (N_1731,N_1658,N_1697);
nor U1732 (N_1732,N_1658,N_1670);
or U1733 (N_1733,N_1683,N_1692);
nor U1734 (N_1734,N_1688,N_1690);
and U1735 (N_1735,N_1691,N_1650);
and U1736 (N_1736,N_1656,N_1693);
nand U1737 (N_1737,N_1680,N_1664);
nor U1738 (N_1738,N_1696,N_1675);
or U1739 (N_1739,N_1697,N_1669);
or U1740 (N_1740,N_1697,N_1691);
and U1741 (N_1741,N_1695,N_1676);
nor U1742 (N_1742,N_1683,N_1694);
nand U1743 (N_1743,N_1657,N_1674);
and U1744 (N_1744,N_1653,N_1672);
nand U1745 (N_1745,N_1654,N_1688);
and U1746 (N_1746,N_1677,N_1692);
xnor U1747 (N_1747,N_1686,N_1661);
and U1748 (N_1748,N_1659,N_1653);
nor U1749 (N_1749,N_1687,N_1660);
nand U1750 (N_1750,N_1703,N_1727);
nor U1751 (N_1751,N_1717,N_1706);
nor U1752 (N_1752,N_1713,N_1705);
and U1753 (N_1753,N_1726,N_1743);
and U1754 (N_1754,N_1730,N_1710);
nor U1755 (N_1755,N_1734,N_1736);
and U1756 (N_1756,N_1746,N_1716);
nor U1757 (N_1757,N_1745,N_1724);
and U1758 (N_1758,N_1725,N_1731);
nand U1759 (N_1759,N_1735,N_1739);
nand U1760 (N_1760,N_1715,N_1729);
or U1761 (N_1761,N_1748,N_1742);
nor U1762 (N_1762,N_1749,N_1722);
or U1763 (N_1763,N_1711,N_1747);
and U1764 (N_1764,N_1700,N_1737);
nor U1765 (N_1765,N_1701,N_1709);
nor U1766 (N_1766,N_1740,N_1733);
nor U1767 (N_1767,N_1728,N_1720);
nand U1768 (N_1768,N_1712,N_1738);
or U1769 (N_1769,N_1744,N_1721);
and U1770 (N_1770,N_1719,N_1741);
nor U1771 (N_1771,N_1704,N_1702);
xnor U1772 (N_1772,N_1708,N_1732);
nor U1773 (N_1773,N_1714,N_1718);
or U1774 (N_1774,N_1723,N_1707);
or U1775 (N_1775,N_1730,N_1702);
and U1776 (N_1776,N_1740,N_1700);
and U1777 (N_1777,N_1705,N_1703);
or U1778 (N_1778,N_1705,N_1748);
nor U1779 (N_1779,N_1708,N_1717);
nand U1780 (N_1780,N_1720,N_1741);
or U1781 (N_1781,N_1717,N_1715);
and U1782 (N_1782,N_1715,N_1749);
nand U1783 (N_1783,N_1739,N_1716);
nor U1784 (N_1784,N_1739,N_1748);
nand U1785 (N_1785,N_1701,N_1712);
and U1786 (N_1786,N_1700,N_1702);
nand U1787 (N_1787,N_1740,N_1715);
and U1788 (N_1788,N_1728,N_1730);
or U1789 (N_1789,N_1717,N_1719);
or U1790 (N_1790,N_1741,N_1713);
or U1791 (N_1791,N_1738,N_1707);
nor U1792 (N_1792,N_1744,N_1707);
and U1793 (N_1793,N_1726,N_1723);
nor U1794 (N_1794,N_1729,N_1709);
nand U1795 (N_1795,N_1729,N_1714);
or U1796 (N_1796,N_1745,N_1712);
nor U1797 (N_1797,N_1722,N_1743);
nor U1798 (N_1798,N_1705,N_1739);
nor U1799 (N_1799,N_1749,N_1713);
and U1800 (N_1800,N_1774,N_1782);
and U1801 (N_1801,N_1751,N_1786);
nor U1802 (N_1802,N_1783,N_1770);
nand U1803 (N_1803,N_1775,N_1757);
and U1804 (N_1804,N_1787,N_1789);
nor U1805 (N_1805,N_1756,N_1750);
nor U1806 (N_1806,N_1766,N_1761);
or U1807 (N_1807,N_1753,N_1798);
and U1808 (N_1808,N_1779,N_1758);
nor U1809 (N_1809,N_1765,N_1796);
or U1810 (N_1810,N_1772,N_1778);
and U1811 (N_1811,N_1791,N_1773);
nor U1812 (N_1812,N_1768,N_1780);
nand U1813 (N_1813,N_1777,N_1794);
nand U1814 (N_1814,N_1759,N_1767);
nand U1815 (N_1815,N_1771,N_1763);
or U1816 (N_1816,N_1788,N_1792);
nor U1817 (N_1817,N_1781,N_1754);
and U1818 (N_1818,N_1776,N_1793);
nor U1819 (N_1819,N_1769,N_1760);
or U1820 (N_1820,N_1755,N_1795);
or U1821 (N_1821,N_1752,N_1785);
or U1822 (N_1822,N_1790,N_1797);
and U1823 (N_1823,N_1762,N_1764);
and U1824 (N_1824,N_1799,N_1784);
and U1825 (N_1825,N_1774,N_1783);
xor U1826 (N_1826,N_1772,N_1770);
or U1827 (N_1827,N_1792,N_1797);
and U1828 (N_1828,N_1786,N_1778);
and U1829 (N_1829,N_1763,N_1776);
and U1830 (N_1830,N_1759,N_1761);
nor U1831 (N_1831,N_1796,N_1763);
or U1832 (N_1832,N_1756,N_1779);
nor U1833 (N_1833,N_1797,N_1782);
nand U1834 (N_1834,N_1756,N_1753);
or U1835 (N_1835,N_1768,N_1791);
or U1836 (N_1836,N_1769,N_1790);
nand U1837 (N_1837,N_1750,N_1791);
nand U1838 (N_1838,N_1762,N_1794);
xnor U1839 (N_1839,N_1758,N_1775);
nor U1840 (N_1840,N_1757,N_1767);
or U1841 (N_1841,N_1757,N_1769);
and U1842 (N_1842,N_1795,N_1798);
and U1843 (N_1843,N_1763,N_1784);
and U1844 (N_1844,N_1776,N_1798);
or U1845 (N_1845,N_1788,N_1752);
nand U1846 (N_1846,N_1753,N_1784);
nand U1847 (N_1847,N_1765,N_1795);
or U1848 (N_1848,N_1791,N_1796);
and U1849 (N_1849,N_1776,N_1784);
nor U1850 (N_1850,N_1837,N_1803);
and U1851 (N_1851,N_1815,N_1808);
nand U1852 (N_1852,N_1840,N_1804);
and U1853 (N_1853,N_1836,N_1819);
or U1854 (N_1854,N_1832,N_1818);
and U1855 (N_1855,N_1807,N_1847);
and U1856 (N_1856,N_1805,N_1846);
nor U1857 (N_1857,N_1849,N_1831);
or U1858 (N_1858,N_1834,N_1813);
nor U1859 (N_1859,N_1821,N_1806);
nand U1860 (N_1860,N_1800,N_1833);
and U1861 (N_1861,N_1845,N_1839);
nand U1862 (N_1862,N_1844,N_1828);
nor U1863 (N_1863,N_1835,N_1841);
nand U1864 (N_1864,N_1811,N_1824);
nand U1865 (N_1865,N_1822,N_1830);
nand U1866 (N_1866,N_1829,N_1827);
nand U1867 (N_1867,N_1812,N_1801);
nand U1868 (N_1868,N_1817,N_1838);
nor U1869 (N_1869,N_1848,N_1825);
nand U1870 (N_1870,N_1823,N_1814);
and U1871 (N_1871,N_1826,N_1809);
or U1872 (N_1872,N_1843,N_1810);
nor U1873 (N_1873,N_1802,N_1820);
or U1874 (N_1874,N_1842,N_1816);
or U1875 (N_1875,N_1835,N_1816);
nand U1876 (N_1876,N_1810,N_1818);
or U1877 (N_1877,N_1819,N_1831);
nor U1878 (N_1878,N_1805,N_1837);
or U1879 (N_1879,N_1842,N_1812);
and U1880 (N_1880,N_1839,N_1837);
nand U1881 (N_1881,N_1829,N_1805);
or U1882 (N_1882,N_1816,N_1825);
and U1883 (N_1883,N_1810,N_1822);
nor U1884 (N_1884,N_1811,N_1828);
nand U1885 (N_1885,N_1805,N_1810);
or U1886 (N_1886,N_1845,N_1811);
nor U1887 (N_1887,N_1839,N_1806);
or U1888 (N_1888,N_1814,N_1801);
nor U1889 (N_1889,N_1837,N_1815);
nand U1890 (N_1890,N_1823,N_1829);
or U1891 (N_1891,N_1835,N_1809);
or U1892 (N_1892,N_1815,N_1846);
nor U1893 (N_1893,N_1811,N_1820);
nor U1894 (N_1894,N_1848,N_1821);
nor U1895 (N_1895,N_1825,N_1815);
and U1896 (N_1896,N_1823,N_1842);
nor U1897 (N_1897,N_1836,N_1808);
nand U1898 (N_1898,N_1838,N_1849);
nand U1899 (N_1899,N_1803,N_1810);
or U1900 (N_1900,N_1894,N_1878);
nand U1901 (N_1901,N_1890,N_1897);
nor U1902 (N_1902,N_1899,N_1852);
xnor U1903 (N_1903,N_1850,N_1857);
or U1904 (N_1904,N_1874,N_1865);
and U1905 (N_1905,N_1873,N_1856);
nor U1906 (N_1906,N_1863,N_1858);
and U1907 (N_1907,N_1884,N_1853);
or U1908 (N_1908,N_1886,N_1892);
or U1909 (N_1909,N_1891,N_1870);
nand U1910 (N_1910,N_1872,N_1866);
nor U1911 (N_1911,N_1861,N_1859);
nand U1912 (N_1912,N_1895,N_1880);
nand U1913 (N_1913,N_1887,N_1862);
nand U1914 (N_1914,N_1869,N_1885);
nand U1915 (N_1915,N_1868,N_1876);
nand U1916 (N_1916,N_1893,N_1855);
or U1917 (N_1917,N_1871,N_1879);
or U1918 (N_1918,N_1877,N_1851);
nand U1919 (N_1919,N_1888,N_1864);
or U1920 (N_1920,N_1881,N_1882);
and U1921 (N_1921,N_1883,N_1854);
nor U1922 (N_1922,N_1896,N_1875);
or U1923 (N_1923,N_1867,N_1860);
and U1924 (N_1924,N_1898,N_1889);
nor U1925 (N_1925,N_1856,N_1881);
or U1926 (N_1926,N_1883,N_1856);
or U1927 (N_1927,N_1886,N_1897);
and U1928 (N_1928,N_1898,N_1866);
nor U1929 (N_1929,N_1889,N_1856);
and U1930 (N_1930,N_1854,N_1857);
nand U1931 (N_1931,N_1881,N_1864);
or U1932 (N_1932,N_1876,N_1869);
nand U1933 (N_1933,N_1896,N_1886);
nor U1934 (N_1934,N_1884,N_1852);
or U1935 (N_1935,N_1864,N_1870);
nand U1936 (N_1936,N_1884,N_1854);
nor U1937 (N_1937,N_1894,N_1855);
nor U1938 (N_1938,N_1879,N_1868);
nor U1939 (N_1939,N_1898,N_1854);
nand U1940 (N_1940,N_1878,N_1884);
and U1941 (N_1941,N_1850,N_1852);
nor U1942 (N_1942,N_1852,N_1870);
nor U1943 (N_1943,N_1875,N_1893);
nor U1944 (N_1944,N_1853,N_1893);
and U1945 (N_1945,N_1890,N_1853);
nand U1946 (N_1946,N_1859,N_1880);
and U1947 (N_1947,N_1851,N_1889);
or U1948 (N_1948,N_1882,N_1870);
nor U1949 (N_1949,N_1853,N_1877);
xor U1950 (N_1950,N_1916,N_1931);
nand U1951 (N_1951,N_1926,N_1914);
and U1952 (N_1952,N_1929,N_1937);
and U1953 (N_1953,N_1910,N_1928);
nand U1954 (N_1954,N_1923,N_1920);
or U1955 (N_1955,N_1949,N_1903);
and U1956 (N_1956,N_1927,N_1941);
or U1957 (N_1957,N_1924,N_1934);
nand U1958 (N_1958,N_1945,N_1913);
nand U1959 (N_1959,N_1947,N_1900);
nor U1960 (N_1960,N_1948,N_1922);
nand U1961 (N_1961,N_1912,N_1909);
or U1962 (N_1962,N_1911,N_1943);
or U1963 (N_1963,N_1942,N_1939);
nor U1964 (N_1964,N_1908,N_1946);
or U1965 (N_1965,N_1906,N_1904);
nor U1966 (N_1966,N_1940,N_1915);
and U1967 (N_1967,N_1907,N_1919);
or U1968 (N_1968,N_1918,N_1917);
nand U1969 (N_1969,N_1902,N_1932);
nor U1970 (N_1970,N_1930,N_1901);
and U1971 (N_1971,N_1933,N_1925);
and U1972 (N_1972,N_1936,N_1935);
nor U1973 (N_1973,N_1944,N_1905);
or U1974 (N_1974,N_1938,N_1921);
nand U1975 (N_1975,N_1944,N_1929);
nor U1976 (N_1976,N_1941,N_1935);
nor U1977 (N_1977,N_1932,N_1924);
nand U1978 (N_1978,N_1942,N_1902);
nor U1979 (N_1979,N_1929,N_1909);
and U1980 (N_1980,N_1904,N_1940);
or U1981 (N_1981,N_1933,N_1901);
and U1982 (N_1982,N_1916,N_1911);
nor U1983 (N_1983,N_1941,N_1909);
or U1984 (N_1984,N_1907,N_1925);
nor U1985 (N_1985,N_1904,N_1930);
or U1986 (N_1986,N_1910,N_1946);
nand U1987 (N_1987,N_1927,N_1901);
and U1988 (N_1988,N_1945,N_1925);
or U1989 (N_1989,N_1902,N_1916);
nand U1990 (N_1990,N_1945,N_1938);
nor U1991 (N_1991,N_1926,N_1945);
and U1992 (N_1992,N_1944,N_1906);
nor U1993 (N_1993,N_1918,N_1940);
or U1994 (N_1994,N_1946,N_1940);
and U1995 (N_1995,N_1948,N_1925);
nor U1996 (N_1996,N_1923,N_1944);
or U1997 (N_1997,N_1904,N_1914);
nand U1998 (N_1998,N_1935,N_1932);
and U1999 (N_1999,N_1905,N_1938);
and U2000 (N_2000,N_1973,N_1965);
and U2001 (N_2001,N_1979,N_1989);
nand U2002 (N_2002,N_1974,N_1959);
nor U2003 (N_2003,N_1958,N_1992);
and U2004 (N_2004,N_1957,N_1999);
or U2005 (N_2005,N_1985,N_1978);
nand U2006 (N_2006,N_1955,N_1987);
nand U2007 (N_2007,N_1995,N_1986);
or U2008 (N_2008,N_1983,N_1954);
nand U2009 (N_2009,N_1975,N_1969);
and U2010 (N_2010,N_1956,N_1951);
nor U2011 (N_2011,N_1982,N_1964);
and U2012 (N_2012,N_1966,N_1984);
and U2013 (N_2013,N_1990,N_1950);
nor U2014 (N_2014,N_1993,N_1996);
nand U2015 (N_2015,N_1970,N_1953);
or U2016 (N_2016,N_1976,N_1972);
and U2017 (N_2017,N_1988,N_1971);
nand U2018 (N_2018,N_1994,N_1991);
and U2019 (N_2019,N_1960,N_1980);
and U2020 (N_2020,N_1998,N_1967);
nor U2021 (N_2021,N_1961,N_1997);
nor U2022 (N_2022,N_1977,N_1952);
or U2023 (N_2023,N_1963,N_1968);
and U2024 (N_2024,N_1981,N_1962);
or U2025 (N_2025,N_1974,N_1975);
or U2026 (N_2026,N_1963,N_1961);
and U2027 (N_2027,N_1950,N_1998);
or U2028 (N_2028,N_1987,N_1973);
nand U2029 (N_2029,N_1974,N_1986);
nor U2030 (N_2030,N_1952,N_1964);
and U2031 (N_2031,N_1998,N_1951);
nand U2032 (N_2032,N_1957,N_1964);
or U2033 (N_2033,N_1981,N_1980);
and U2034 (N_2034,N_1959,N_1960);
nand U2035 (N_2035,N_1999,N_1951);
and U2036 (N_2036,N_1990,N_1960);
nand U2037 (N_2037,N_1988,N_1954);
and U2038 (N_2038,N_1996,N_1987);
nand U2039 (N_2039,N_1965,N_1975);
nor U2040 (N_2040,N_1989,N_1953);
and U2041 (N_2041,N_1981,N_1985);
and U2042 (N_2042,N_1983,N_1985);
and U2043 (N_2043,N_1998,N_1996);
and U2044 (N_2044,N_1952,N_1960);
nor U2045 (N_2045,N_1989,N_1978);
nand U2046 (N_2046,N_1965,N_1972);
or U2047 (N_2047,N_1968,N_1978);
or U2048 (N_2048,N_1997,N_1994);
nand U2049 (N_2049,N_1982,N_1970);
or U2050 (N_2050,N_2021,N_2030);
nor U2051 (N_2051,N_2027,N_2015);
and U2052 (N_2052,N_2019,N_2009);
or U2053 (N_2053,N_2006,N_2026);
nand U2054 (N_2054,N_2020,N_2002);
nand U2055 (N_2055,N_2043,N_2038);
and U2056 (N_2056,N_2013,N_2047);
nand U2057 (N_2057,N_2035,N_2025);
nand U2058 (N_2058,N_2016,N_2040);
or U2059 (N_2059,N_2007,N_2008);
nand U2060 (N_2060,N_2028,N_2014);
and U2061 (N_2061,N_2024,N_2037);
and U2062 (N_2062,N_2033,N_2023);
nor U2063 (N_2063,N_2005,N_2018);
nand U2064 (N_2064,N_2010,N_2003);
nand U2065 (N_2065,N_2048,N_2017);
nand U2066 (N_2066,N_2012,N_2001);
nand U2067 (N_2067,N_2045,N_2044);
or U2068 (N_2068,N_2042,N_2049);
nand U2069 (N_2069,N_2034,N_2004);
nor U2070 (N_2070,N_2046,N_2032);
nor U2071 (N_2071,N_2039,N_2031);
nand U2072 (N_2072,N_2036,N_2029);
or U2073 (N_2073,N_2000,N_2011);
nor U2074 (N_2074,N_2022,N_2041);
nand U2075 (N_2075,N_2022,N_2019);
nor U2076 (N_2076,N_2003,N_2028);
and U2077 (N_2077,N_2011,N_2014);
nand U2078 (N_2078,N_2032,N_2012);
or U2079 (N_2079,N_2020,N_2007);
or U2080 (N_2080,N_2026,N_2019);
and U2081 (N_2081,N_2016,N_2037);
nand U2082 (N_2082,N_2045,N_2015);
nor U2083 (N_2083,N_2001,N_2023);
nor U2084 (N_2084,N_2002,N_2046);
nor U2085 (N_2085,N_2045,N_2023);
and U2086 (N_2086,N_2007,N_2012);
and U2087 (N_2087,N_2032,N_2035);
or U2088 (N_2088,N_2013,N_2000);
nand U2089 (N_2089,N_2047,N_2021);
or U2090 (N_2090,N_2043,N_2026);
nand U2091 (N_2091,N_2037,N_2033);
and U2092 (N_2092,N_2028,N_2022);
nand U2093 (N_2093,N_2015,N_2034);
nand U2094 (N_2094,N_2029,N_2002);
or U2095 (N_2095,N_2035,N_2049);
or U2096 (N_2096,N_2034,N_2039);
xor U2097 (N_2097,N_2045,N_2040);
or U2098 (N_2098,N_2015,N_2043);
and U2099 (N_2099,N_2031,N_2026);
nor U2100 (N_2100,N_2079,N_2084);
nor U2101 (N_2101,N_2059,N_2097);
and U2102 (N_2102,N_2094,N_2090);
and U2103 (N_2103,N_2052,N_2068);
nand U2104 (N_2104,N_2099,N_2095);
and U2105 (N_2105,N_2083,N_2064);
nand U2106 (N_2106,N_2063,N_2065);
or U2107 (N_2107,N_2054,N_2091);
nand U2108 (N_2108,N_2060,N_2069);
or U2109 (N_2109,N_2075,N_2087);
nand U2110 (N_2110,N_2092,N_2061);
nand U2111 (N_2111,N_2074,N_2081);
and U2112 (N_2112,N_2057,N_2076);
nor U2113 (N_2113,N_2096,N_2085);
nand U2114 (N_2114,N_2071,N_2073);
or U2115 (N_2115,N_2070,N_2072);
or U2116 (N_2116,N_2056,N_2098);
or U2117 (N_2117,N_2078,N_2051);
and U2118 (N_2118,N_2093,N_2050);
or U2119 (N_2119,N_2066,N_2082);
nor U2120 (N_2120,N_2053,N_2088);
or U2121 (N_2121,N_2086,N_2067);
nand U2122 (N_2122,N_2062,N_2080);
and U2123 (N_2123,N_2058,N_2089);
nand U2124 (N_2124,N_2077,N_2055);
nand U2125 (N_2125,N_2068,N_2085);
or U2126 (N_2126,N_2072,N_2096);
and U2127 (N_2127,N_2071,N_2064);
nor U2128 (N_2128,N_2088,N_2066);
or U2129 (N_2129,N_2083,N_2057);
nor U2130 (N_2130,N_2074,N_2096);
nand U2131 (N_2131,N_2098,N_2059);
nand U2132 (N_2132,N_2098,N_2087);
or U2133 (N_2133,N_2053,N_2076);
nand U2134 (N_2134,N_2059,N_2099);
or U2135 (N_2135,N_2058,N_2069);
xor U2136 (N_2136,N_2054,N_2095);
nand U2137 (N_2137,N_2058,N_2061);
and U2138 (N_2138,N_2051,N_2070);
nand U2139 (N_2139,N_2080,N_2097);
and U2140 (N_2140,N_2084,N_2072);
nor U2141 (N_2141,N_2073,N_2070);
and U2142 (N_2142,N_2076,N_2074);
nor U2143 (N_2143,N_2061,N_2068);
or U2144 (N_2144,N_2053,N_2098);
or U2145 (N_2145,N_2096,N_2056);
nor U2146 (N_2146,N_2062,N_2087);
nand U2147 (N_2147,N_2081,N_2084);
nand U2148 (N_2148,N_2057,N_2088);
and U2149 (N_2149,N_2050,N_2069);
nand U2150 (N_2150,N_2141,N_2148);
and U2151 (N_2151,N_2138,N_2111);
nor U2152 (N_2152,N_2122,N_2139);
nor U2153 (N_2153,N_2103,N_2114);
or U2154 (N_2154,N_2124,N_2126);
or U2155 (N_2155,N_2134,N_2147);
nor U2156 (N_2156,N_2131,N_2132);
or U2157 (N_2157,N_2146,N_2125);
nand U2158 (N_2158,N_2106,N_2127);
and U2159 (N_2159,N_2115,N_2133);
nor U2160 (N_2160,N_2107,N_2144);
and U2161 (N_2161,N_2102,N_2130);
nand U2162 (N_2162,N_2117,N_2136);
nand U2163 (N_2163,N_2105,N_2104);
or U2164 (N_2164,N_2120,N_2112);
or U2165 (N_2165,N_2118,N_2129);
or U2166 (N_2166,N_2145,N_2123);
nand U2167 (N_2167,N_2108,N_2143);
and U2168 (N_2168,N_2116,N_2137);
nand U2169 (N_2169,N_2142,N_2135);
and U2170 (N_2170,N_2101,N_2119);
nand U2171 (N_2171,N_2140,N_2109);
or U2172 (N_2172,N_2121,N_2149);
nor U2173 (N_2173,N_2128,N_2100);
nand U2174 (N_2174,N_2110,N_2113);
or U2175 (N_2175,N_2112,N_2141);
nand U2176 (N_2176,N_2140,N_2111);
or U2177 (N_2177,N_2127,N_2110);
or U2178 (N_2178,N_2135,N_2139);
and U2179 (N_2179,N_2119,N_2141);
nand U2180 (N_2180,N_2111,N_2145);
nand U2181 (N_2181,N_2149,N_2140);
and U2182 (N_2182,N_2143,N_2138);
nor U2183 (N_2183,N_2104,N_2113);
nor U2184 (N_2184,N_2106,N_2117);
nor U2185 (N_2185,N_2117,N_2125);
and U2186 (N_2186,N_2105,N_2134);
or U2187 (N_2187,N_2111,N_2139);
nor U2188 (N_2188,N_2148,N_2101);
nor U2189 (N_2189,N_2113,N_2121);
and U2190 (N_2190,N_2112,N_2124);
or U2191 (N_2191,N_2100,N_2144);
xnor U2192 (N_2192,N_2141,N_2126);
and U2193 (N_2193,N_2124,N_2108);
nand U2194 (N_2194,N_2122,N_2109);
and U2195 (N_2195,N_2101,N_2126);
or U2196 (N_2196,N_2147,N_2125);
or U2197 (N_2197,N_2139,N_2116);
or U2198 (N_2198,N_2106,N_2142);
nor U2199 (N_2199,N_2113,N_2139);
nor U2200 (N_2200,N_2160,N_2181);
or U2201 (N_2201,N_2165,N_2176);
nand U2202 (N_2202,N_2152,N_2161);
and U2203 (N_2203,N_2196,N_2177);
or U2204 (N_2204,N_2180,N_2187);
or U2205 (N_2205,N_2193,N_2171);
and U2206 (N_2206,N_2199,N_2184);
or U2207 (N_2207,N_2179,N_2197);
nand U2208 (N_2208,N_2163,N_2158);
nor U2209 (N_2209,N_2154,N_2175);
nor U2210 (N_2210,N_2155,N_2166);
nor U2211 (N_2211,N_2153,N_2188);
and U2212 (N_2212,N_2182,N_2183);
and U2213 (N_2213,N_2191,N_2151);
and U2214 (N_2214,N_2173,N_2157);
and U2215 (N_2215,N_2150,N_2162);
nand U2216 (N_2216,N_2192,N_2186);
or U2217 (N_2217,N_2156,N_2198);
or U2218 (N_2218,N_2168,N_2185);
nor U2219 (N_2219,N_2172,N_2189);
and U2220 (N_2220,N_2174,N_2178);
and U2221 (N_2221,N_2164,N_2159);
nand U2222 (N_2222,N_2194,N_2167);
nor U2223 (N_2223,N_2169,N_2170);
nand U2224 (N_2224,N_2195,N_2190);
or U2225 (N_2225,N_2199,N_2189);
nand U2226 (N_2226,N_2186,N_2179);
and U2227 (N_2227,N_2194,N_2175);
and U2228 (N_2228,N_2194,N_2151);
nor U2229 (N_2229,N_2155,N_2187);
or U2230 (N_2230,N_2165,N_2173);
nor U2231 (N_2231,N_2166,N_2170);
and U2232 (N_2232,N_2193,N_2195);
and U2233 (N_2233,N_2151,N_2152);
or U2234 (N_2234,N_2182,N_2179);
or U2235 (N_2235,N_2164,N_2156);
nand U2236 (N_2236,N_2156,N_2167);
nor U2237 (N_2237,N_2164,N_2181);
nor U2238 (N_2238,N_2195,N_2192);
nand U2239 (N_2239,N_2167,N_2174);
and U2240 (N_2240,N_2183,N_2190);
nor U2241 (N_2241,N_2163,N_2151);
and U2242 (N_2242,N_2195,N_2182);
or U2243 (N_2243,N_2192,N_2165);
and U2244 (N_2244,N_2188,N_2181);
and U2245 (N_2245,N_2193,N_2190);
nor U2246 (N_2246,N_2184,N_2188);
nor U2247 (N_2247,N_2186,N_2188);
nand U2248 (N_2248,N_2193,N_2165);
nor U2249 (N_2249,N_2168,N_2179);
and U2250 (N_2250,N_2238,N_2212);
nand U2251 (N_2251,N_2224,N_2213);
and U2252 (N_2252,N_2208,N_2237);
nor U2253 (N_2253,N_2246,N_2203);
nand U2254 (N_2254,N_2200,N_2220);
nand U2255 (N_2255,N_2229,N_2245);
nand U2256 (N_2256,N_2234,N_2227);
nand U2257 (N_2257,N_2247,N_2210);
nand U2258 (N_2258,N_2241,N_2211);
nand U2259 (N_2259,N_2235,N_2230);
or U2260 (N_2260,N_2207,N_2202);
or U2261 (N_2261,N_2223,N_2236);
or U2262 (N_2262,N_2204,N_2201);
nand U2263 (N_2263,N_2226,N_2218);
nor U2264 (N_2264,N_2242,N_2222);
nor U2265 (N_2265,N_2206,N_2233);
and U2266 (N_2266,N_2232,N_2205);
nor U2267 (N_2267,N_2248,N_2221);
nor U2268 (N_2268,N_2243,N_2239);
and U2269 (N_2269,N_2219,N_2216);
nand U2270 (N_2270,N_2214,N_2209);
nor U2271 (N_2271,N_2249,N_2225);
or U2272 (N_2272,N_2240,N_2215);
or U2273 (N_2273,N_2217,N_2228);
nor U2274 (N_2274,N_2244,N_2231);
and U2275 (N_2275,N_2227,N_2230);
nand U2276 (N_2276,N_2226,N_2242);
and U2277 (N_2277,N_2206,N_2239);
nor U2278 (N_2278,N_2214,N_2213);
xnor U2279 (N_2279,N_2204,N_2243);
or U2280 (N_2280,N_2202,N_2239);
and U2281 (N_2281,N_2218,N_2224);
nand U2282 (N_2282,N_2244,N_2247);
nor U2283 (N_2283,N_2238,N_2240);
and U2284 (N_2284,N_2235,N_2242);
and U2285 (N_2285,N_2219,N_2230);
nor U2286 (N_2286,N_2242,N_2245);
nand U2287 (N_2287,N_2234,N_2243);
and U2288 (N_2288,N_2245,N_2232);
nand U2289 (N_2289,N_2233,N_2241);
nand U2290 (N_2290,N_2228,N_2210);
nand U2291 (N_2291,N_2232,N_2218);
or U2292 (N_2292,N_2244,N_2242);
nand U2293 (N_2293,N_2235,N_2203);
nand U2294 (N_2294,N_2211,N_2240);
nor U2295 (N_2295,N_2204,N_2239);
nor U2296 (N_2296,N_2211,N_2246);
nand U2297 (N_2297,N_2229,N_2239);
or U2298 (N_2298,N_2200,N_2238);
and U2299 (N_2299,N_2240,N_2221);
nand U2300 (N_2300,N_2275,N_2294);
nand U2301 (N_2301,N_2289,N_2261);
and U2302 (N_2302,N_2251,N_2254);
or U2303 (N_2303,N_2272,N_2288);
or U2304 (N_2304,N_2271,N_2298);
nor U2305 (N_2305,N_2290,N_2255);
or U2306 (N_2306,N_2286,N_2287);
nand U2307 (N_2307,N_2264,N_2268);
nor U2308 (N_2308,N_2276,N_2267);
and U2309 (N_2309,N_2259,N_2280);
nand U2310 (N_2310,N_2282,N_2296);
xnor U2311 (N_2311,N_2292,N_2266);
and U2312 (N_2312,N_2284,N_2278);
or U2313 (N_2313,N_2256,N_2277);
nor U2314 (N_2314,N_2250,N_2291);
nor U2315 (N_2315,N_2262,N_2257);
nand U2316 (N_2316,N_2252,N_2263);
and U2317 (N_2317,N_2297,N_2258);
and U2318 (N_2318,N_2285,N_2269);
and U2319 (N_2319,N_2265,N_2273);
nand U2320 (N_2320,N_2274,N_2295);
and U2321 (N_2321,N_2270,N_2283);
and U2322 (N_2322,N_2260,N_2293);
or U2323 (N_2323,N_2281,N_2299);
or U2324 (N_2324,N_2279,N_2253);
nor U2325 (N_2325,N_2259,N_2258);
or U2326 (N_2326,N_2288,N_2256);
or U2327 (N_2327,N_2270,N_2261);
and U2328 (N_2328,N_2267,N_2286);
or U2329 (N_2329,N_2275,N_2259);
or U2330 (N_2330,N_2277,N_2292);
nand U2331 (N_2331,N_2281,N_2259);
xor U2332 (N_2332,N_2297,N_2277);
and U2333 (N_2333,N_2265,N_2291);
and U2334 (N_2334,N_2293,N_2297);
or U2335 (N_2335,N_2274,N_2283);
nor U2336 (N_2336,N_2276,N_2287);
nand U2337 (N_2337,N_2269,N_2280);
nor U2338 (N_2338,N_2288,N_2273);
nor U2339 (N_2339,N_2284,N_2250);
or U2340 (N_2340,N_2273,N_2285);
nor U2341 (N_2341,N_2295,N_2263);
or U2342 (N_2342,N_2257,N_2281);
and U2343 (N_2343,N_2271,N_2253);
or U2344 (N_2344,N_2284,N_2254);
or U2345 (N_2345,N_2291,N_2277);
and U2346 (N_2346,N_2253,N_2291);
or U2347 (N_2347,N_2298,N_2283);
nand U2348 (N_2348,N_2252,N_2253);
and U2349 (N_2349,N_2250,N_2283);
and U2350 (N_2350,N_2313,N_2315);
or U2351 (N_2351,N_2303,N_2322);
xor U2352 (N_2352,N_2346,N_2312);
or U2353 (N_2353,N_2307,N_2302);
and U2354 (N_2354,N_2304,N_2338);
nand U2355 (N_2355,N_2335,N_2331);
nand U2356 (N_2356,N_2301,N_2316);
or U2357 (N_2357,N_2344,N_2311);
and U2358 (N_2358,N_2349,N_2323);
and U2359 (N_2359,N_2300,N_2345);
or U2360 (N_2360,N_2347,N_2339);
nor U2361 (N_2361,N_2333,N_2348);
or U2362 (N_2362,N_2327,N_2318);
or U2363 (N_2363,N_2343,N_2334);
and U2364 (N_2364,N_2324,N_2336);
or U2365 (N_2365,N_2337,N_2309);
nor U2366 (N_2366,N_2306,N_2332);
or U2367 (N_2367,N_2340,N_2308);
nand U2368 (N_2368,N_2314,N_2329);
and U2369 (N_2369,N_2310,N_2305);
nor U2370 (N_2370,N_2330,N_2320);
and U2371 (N_2371,N_2319,N_2321);
or U2372 (N_2372,N_2317,N_2341);
nor U2373 (N_2373,N_2325,N_2326);
nand U2374 (N_2374,N_2328,N_2342);
and U2375 (N_2375,N_2332,N_2317);
nand U2376 (N_2376,N_2335,N_2312);
or U2377 (N_2377,N_2306,N_2320);
and U2378 (N_2378,N_2348,N_2346);
nor U2379 (N_2379,N_2332,N_2345);
nand U2380 (N_2380,N_2339,N_2321);
nand U2381 (N_2381,N_2349,N_2343);
or U2382 (N_2382,N_2316,N_2305);
nand U2383 (N_2383,N_2324,N_2303);
or U2384 (N_2384,N_2303,N_2304);
nand U2385 (N_2385,N_2334,N_2346);
nor U2386 (N_2386,N_2335,N_2334);
nor U2387 (N_2387,N_2300,N_2304);
or U2388 (N_2388,N_2300,N_2323);
nand U2389 (N_2389,N_2333,N_2349);
nand U2390 (N_2390,N_2327,N_2341);
or U2391 (N_2391,N_2341,N_2335);
or U2392 (N_2392,N_2308,N_2312);
or U2393 (N_2393,N_2344,N_2340);
nor U2394 (N_2394,N_2328,N_2311);
nand U2395 (N_2395,N_2311,N_2329);
or U2396 (N_2396,N_2343,N_2332);
nand U2397 (N_2397,N_2334,N_2306);
nand U2398 (N_2398,N_2322,N_2314);
nand U2399 (N_2399,N_2311,N_2304);
nand U2400 (N_2400,N_2365,N_2395);
or U2401 (N_2401,N_2392,N_2379);
and U2402 (N_2402,N_2376,N_2374);
or U2403 (N_2403,N_2355,N_2352);
nand U2404 (N_2404,N_2354,N_2386);
nand U2405 (N_2405,N_2362,N_2351);
or U2406 (N_2406,N_2389,N_2381);
or U2407 (N_2407,N_2364,N_2357);
nand U2408 (N_2408,N_2353,N_2373);
or U2409 (N_2409,N_2394,N_2382);
or U2410 (N_2410,N_2380,N_2359);
nor U2411 (N_2411,N_2385,N_2360);
and U2412 (N_2412,N_2377,N_2363);
or U2413 (N_2413,N_2370,N_2388);
or U2414 (N_2414,N_2367,N_2361);
or U2415 (N_2415,N_2391,N_2384);
or U2416 (N_2416,N_2368,N_2366);
and U2417 (N_2417,N_2383,N_2397);
or U2418 (N_2418,N_2393,N_2378);
nor U2419 (N_2419,N_2387,N_2369);
nand U2420 (N_2420,N_2371,N_2375);
and U2421 (N_2421,N_2356,N_2358);
nand U2422 (N_2422,N_2372,N_2390);
and U2423 (N_2423,N_2399,N_2398);
or U2424 (N_2424,N_2350,N_2396);
or U2425 (N_2425,N_2397,N_2369);
nand U2426 (N_2426,N_2373,N_2384);
nand U2427 (N_2427,N_2375,N_2390);
and U2428 (N_2428,N_2360,N_2374);
nor U2429 (N_2429,N_2385,N_2378);
or U2430 (N_2430,N_2387,N_2388);
or U2431 (N_2431,N_2353,N_2388);
nand U2432 (N_2432,N_2363,N_2370);
nand U2433 (N_2433,N_2358,N_2381);
nor U2434 (N_2434,N_2360,N_2358);
nand U2435 (N_2435,N_2379,N_2370);
nor U2436 (N_2436,N_2384,N_2399);
nand U2437 (N_2437,N_2380,N_2365);
or U2438 (N_2438,N_2367,N_2356);
nor U2439 (N_2439,N_2350,N_2374);
nand U2440 (N_2440,N_2356,N_2382);
nor U2441 (N_2441,N_2363,N_2365);
and U2442 (N_2442,N_2386,N_2376);
and U2443 (N_2443,N_2371,N_2384);
nand U2444 (N_2444,N_2361,N_2360);
nor U2445 (N_2445,N_2389,N_2353);
nand U2446 (N_2446,N_2388,N_2391);
and U2447 (N_2447,N_2385,N_2394);
nor U2448 (N_2448,N_2392,N_2360);
nand U2449 (N_2449,N_2361,N_2354);
nor U2450 (N_2450,N_2430,N_2422);
nor U2451 (N_2451,N_2441,N_2404);
and U2452 (N_2452,N_2411,N_2412);
or U2453 (N_2453,N_2424,N_2406);
nand U2454 (N_2454,N_2447,N_2428);
and U2455 (N_2455,N_2416,N_2449);
nand U2456 (N_2456,N_2420,N_2407);
nand U2457 (N_2457,N_2409,N_2437);
nor U2458 (N_2458,N_2442,N_2425);
or U2459 (N_2459,N_2429,N_2415);
nor U2460 (N_2460,N_2410,N_2438);
nor U2461 (N_2461,N_2408,N_2444);
and U2462 (N_2462,N_2434,N_2427);
or U2463 (N_2463,N_2433,N_2419);
or U2464 (N_2464,N_2448,N_2421);
xnor U2465 (N_2465,N_2423,N_2440);
xnor U2466 (N_2466,N_2445,N_2436);
or U2467 (N_2467,N_2426,N_2446);
or U2468 (N_2468,N_2417,N_2400);
nand U2469 (N_2469,N_2435,N_2403);
nor U2470 (N_2470,N_2401,N_2431);
or U2471 (N_2471,N_2418,N_2439);
nor U2472 (N_2472,N_2402,N_2432);
nand U2473 (N_2473,N_2405,N_2443);
and U2474 (N_2474,N_2414,N_2413);
nand U2475 (N_2475,N_2413,N_2417);
nor U2476 (N_2476,N_2428,N_2449);
nand U2477 (N_2477,N_2443,N_2444);
nor U2478 (N_2478,N_2449,N_2403);
and U2479 (N_2479,N_2409,N_2426);
or U2480 (N_2480,N_2418,N_2447);
nor U2481 (N_2481,N_2426,N_2404);
nor U2482 (N_2482,N_2417,N_2446);
nor U2483 (N_2483,N_2410,N_2414);
and U2484 (N_2484,N_2433,N_2447);
nor U2485 (N_2485,N_2434,N_2400);
or U2486 (N_2486,N_2434,N_2430);
or U2487 (N_2487,N_2433,N_2416);
nor U2488 (N_2488,N_2436,N_2444);
nor U2489 (N_2489,N_2408,N_2425);
and U2490 (N_2490,N_2435,N_2444);
and U2491 (N_2491,N_2437,N_2444);
or U2492 (N_2492,N_2404,N_2406);
or U2493 (N_2493,N_2403,N_2429);
nor U2494 (N_2494,N_2416,N_2425);
nand U2495 (N_2495,N_2431,N_2403);
nand U2496 (N_2496,N_2417,N_2442);
nand U2497 (N_2497,N_2438,N_2411);
nand U2498 (N_2498,N_2435,N_2418);
or U2499 (N_2499,N_2400,N_2423);
nand U2500 (N_2500,N_2458,N_2495);
or U2501 (N_2501,N_2472,N_2455);
or U2502 (N_2502,N_2477,N_2467);
and U2503 (N_2503,N_2479,N_2493);
or U2504 (N_2504,N_2463,N_2487);
nand U2505 (N_2505,N_2466,N_2454);
and U2506 (N_2506,N_2489,N_2451);
and U2507 (N_2507,N_2482,N_2498);
nor U2508 (N_2508,N_2453,N_2462);
or U2509 (N_2509,N_2484,N_2471);
nor U2510 (N_2510,N_2457,N_2474);
and U2511 (N_2511,N_2452,N_2492);
and U2512 (N_2512,N_2465,N_2478);
nand U2513 (N_2513,N_2464,N_2483);
and U2514 (N_2514,N_2470,N_2497);
nand U2515 (N_2515,N_2496,N_2468);
nand U2516 (N_2516,N_2475,N_2490);
nor U2517 (N_2517,N_2494,N_2456);
or U2518 (N_2518,N_2461,N_2460);
nand U2519 (N_2519,N_2485,N_2491);
nor U2520 (N_2520,N_2476,N_2481);
and U2521 (N_2521,N_2450,N_2499);
or U2522 (N_2522,N_2459,N_2486);
and U2523 (N_2523,N_2473,N_2480);
and U2524 (N_2524,N_2488,N_2469);
nand U2525 (N_2525,N_2479,N_2481);
and U2526 (N_2526,N_2494,N_2498);
xor U2527 (N_2527,N_2498,N_2458);
and U2528 (N_2528,N_2450,N_2460);
or U2529 (N_2529,N_2454,N_2479);
or U2530 (N_2530,N_2493,N_2465);
or U2531 (N_2531,N_2470,N_2474);
nand U2532 (N_2532,N_2455,N_2471);
nor U2533 (N_2533,N_2469,N_2492);
nand U2534 (N_2534,N_2464,N_2495);
nand U2535 (N_2535,N_2469,N_2455);
nand U2536 (N_2536,N_2463,N_2451);
or U2537 (N_2537,N_2487,N_2491);
or U2538 (N_2538,N_2478,N_2456);
and U2539 (N_2539,N_2476,N_2477);
and U2540 (N_2540,N_2457,N_2483);
or U2541 (N_2541,N_2454,N_2491);
or U2542 (N_2542,N_2490,N_2459);
nand U2543 (N_2543,N_2456,N_2486);
or U2544 (N_2544,N_2462,N_2472);
nand U2545 (N_2545,N_2481,N_2495);
nor U2546 (N_2546,N_2472,N_2498);
or U2547 (N_2547,N_2493,N_2495);
nor U2548 (N_2548,N_2499,N_2460);
or U2549 (N_2549,N_2451,N_2457);
or U2550 (N_2550,N_2527,N_2521);
and U2551 (N_2551,N_2511,N_2505);
nor U2552 (N_2552,N_2519,N_2502);
and U2553 (N_2553,N_2534,N_2501);
and U2554 (N_2554,N_2536,N_2529);
or U2555 (N_2555,N_2532,N_2528);
nand U2556 (N_2556,N_2520,N_2541);
and U2557 (N_2557,N_2509,N_2537);
or U2558 (N_2558,N_2514,N_2517);
or U2559 (N_2559,N_2546,N_2510);
or U2560 (N_2560,N_2543,N_2533);
and U2561 (N_2561,N_2538,N_2516);
nor U2562 (N_2562,N_2530,N_2500);
nand U2563 (N_2563,N_2504,N_2513);
nor U2564 (N_2564,N_2548,N_2531);
or U2565 (N_2565,N_2525,N_2507);
nand U2566 (N_2566,N_2544,N_2547);
or U2567 (N_2567,N_2522,N_2512);
nand U2568 (N_2568,N_2503,N_2526);
xor U2569 (N_2569,N_2508,N_2506);
and U2570 (N_2570,N_2542,N_2545);
or U2571 (N_2571,N_2524,N_2523);
nand U2572 (N_2572,N_2549,N_2518);
or U2573 (N_2573,N_2540,N_2535);
nor U2574 (N_2574,N_2539,N_2515);
nand U2575 (N_2575,N_2518,N_2516);
or U2576 (N_2576,N_2528,N_2522);
or U2577 (N_2577,N_2521,N_2511);
nor U2578 (N_2578,N_2532,N_2507);
nor U2579 (N_2579,N_2502,N_2530);
nor U2580 (N_2580,N_2543,N_2529);
and U2581 (N_2581,N_2536,N_2502);
and U2582 (N_2582,N_2506,N_2529);
or U2583 (N_2583,N_2532,N_2522);
nand U2584 (N_2584,N_2504,N_2537);
and U2585 (N_2585,N_2505,N_2528);
nor U2586 (N_2586,N_2532,N_2537);
and U2587 (N_2587,N_2526,N_2521);
nand U2588 (N_2588,N_2508,N_2531);
nand U2589 (N_2589,N_2519,N_2503);
and U2590 (N_2590,N_2523,N_2522);
nand U2591 (N_2591,N_2537,N_2533);
and U2592 (N_2592,N_2542,N_2502);
xor U2593 (N_2593,N_2513,N_2527);
and U2594 (N_2594,N_2544,N_2541);
nor U2595 (N_2595,N_2528,N_2545);
or U2596 (N_2596,N_2517,N_2544);
or U2597 (N_2597,N_2524,N_2502);
or U2598 (N_2598,N_2534,N_2521);
and U2599 (N_2599,N_2509,N_2514);
nand U2600 (N_2600,N_2591,N_2554);
and U2601 (N_2601,N_2564,N_2566);
and U2602 (N_2602,N_2593,N_2573);
or U2603 (N_2603,N_2589,N_2571);
nor U2604 (N_2604,N_2568,N_2596);
nor U2605 (N_2605,N_2561,N_2550);
or U2606 (N_2606,N_2576,N_2588);
and U2607 (N_2607,N_2563,N_2580);
nand U2608 (N_2608,N_2553,N_2572);
and U2609 (N_2609,N_2569,N_2599);
nor U2610 (N_2610,N_2595,N_2598);
nand U2611 (N_2611,N_2575,N_2555);
nor U2612 (N_2612,N_2581,N_2585);
or U2613 (N_2613,N_2590,N_2584);
nor U2614 (N_2614,N_2577,N_2583);
nor U2615 (N_2615,N_2558,N_2570);
nor U2616 (N_2616,N_2559,N_2594);
nor U2617 (N_2617,N_2592,N_2579);
nand U2618 (N_2618,N_2578,N_2574);
nand U2619 (N_2619,N_2557,N_2565);
and U2620 (N_2620,N_2586,N_2556);
or U2621 (N_2621,N_2582,N_2551);
nand U2622 (N_2622,N_2597,N_2587);
or U2623 (N_2623,N_2567,N_2560);
nand U2624 (N_2624,N_2562,N_2552);
nand U2625 (N_2625,N_2556,N_2587);
nor U2626 (N_2626,N_2585,N_2572);
nand U2627 (N_2627,N_2575,N_2559);
or U2628 (N_2628,N_2564,N_2572);
nand U2629 (N_2629,N_2550,N_2552);
and U2630 (N_2630,N_2577,N_2575);
or U2631 (N_2631,N_2579,N_2566);
or U2632 (N_2632,N_2554,N_2595);
nand U2633 (N_2633,N_2560,N_2555);
or U2634 (N_2634,N_2577,N_2562);
nand U2635 (N_2635,N_2555,N_2577);
or U2636 (N_2636,N_2561,N_2577);
and U2637 (N_2637,N_2590,N_2566);
nor U2638 (N_2638,N_2575,N_2580);
or U2639 (N_2639,N_2580,N_2573);
nand U2640 (N_2640,N_2573,N_2557);
or U2641 (N_2641,N_2590,N_2575);
nor U2642 (N_2642,N_2550,N_2588);
xor U2643 (N_2643,N_2553,N_2590);
or U2644 (N_2644,N_2594,N_2593);
and U2645 (N_2645,N_2583,N_2582);
and U2646 (N_2646,N_2578,N_2590);
nor U2647 (N_2647,N_2561,N_2562);
or U2648 (N_2648,N_2577,N_2572);
nand U2649 (N_2649,N_2555,N_2595);
nor U2650 (N_2650,N_2611,N_2640);
and U2651 (N_2651,N_2632,N_2623);
or U2652 (N_2652,N_2613,N_2605);
or U2653 (N_2653,N_2644,N_2647);
nand U2654 (N_2654,N_2646,N_2628);
or U2655 (N_2655,N_2630,N_2600);
nor U2656 (N_2656,N_2635,N_2636);
nor U2657 (N_2657,N_2638,N_2604);
nor U2658 (N_2658,N_2607,N_2634);
and U2659 (N_2659,N_2641,N_2602);
and U2660 (N_2660,N_2624,N_2615);
and U2661 (N_2661,N_2631,N_2642);
nand U2662 (N_2662,N_2614,N_2627);
nand U2663 (N_2663,N_2648,N_2608);
nand U2664 (N_2664,N_2620,N_2609);
and U2665 (N_2665,N_2601,N_2633);
nand U2666 (N_2666,N_2625,N_2621);
xnor U2667 (N_2667,N_2649,N_2622);
or U2668 (N_2668,N_2626,N_2603);
and U2669 (N_2669,N_2629,N_2606);
and U2670 (N_2670,N_2618,N_2643);
nand U2671 (N_2671,N_2616,N_2610);
or U2672 (N_2672,N_2639,N_2637);
or U2673 (N_2673,N_2619,N_2645);
and U2674 (N_2674,N_2612,N_2617);
nor U2675 (N_2675,N_2639,N_2612);
and U2676 (N_2676,N_2643,N_2609);
and U2677 (N_2677,N_2634,N_2642);
nand U2678 (N_2678,N_2640,N_2619);
or U2679 (N_2679,N_2618,N_2649);
nor U2680 (N_2680,N_2633,N_2604);
nand U2681 (N_2681,N_2600,N_2608);
or U2682 (N_2682,N_2634,N_2620);
nand U2683 (N_2683,N_2633,N_2637);
or U2684 (N_2684,N_2602,N_2617);
nor U2685 (N_2685,N_2625,N_2646);
nor U2686 (N_2686,N_2614,N_2638);
nor U2687 (N_2687,N_2615,N_2643);
xnor U2688 (N_2688,N_2610,N_2617);
or U2689 (N_2689,N_2620,N_2645);
or U2690 (N_2690,N_2623,N_2618);
nor U2691 (N_2691,N_2604,N_2625);
and U2692 (N_2692,N_2616,N_2628);
nor U2693 (N_2693,N_2604,N_2648);
and U2694 (N_2694,N_2634,N_2639);
xor U2695 (N_2695,N_2611,N_2625);
and U2696 (N_2696,N_2645,N_2627);
or U2697 (N_2697,N_2612,N_2622);
xor U2698 (N_2698,N_2627,N_2618);
nor U2699 (N_2699,N_2637,N_2649);
nor U2700 (N_2700,N_2664,N_2684);
nor U2701 (N_2701,N_2693,N_2656);
or U2702 (N_2702,N_2686,N_2651);
nand U2703 (N_2703,N_2653,N_2668);
nor U2704 (N_2704,N_2687,N_2663);
or U2705 (N_2705,N_2690,N_2671);
nor U2706 (N_2706,N_2679,N_2660);
and U2707 (N_2707,N_2675,N_2692);
xnor U2708 (N_2708,N_2677,N_2657);
or U2709 (N_2709,N_2691,N_2670);
nand U2710 (N_2710,N_2652,N_2669);
or U2711 (N_2711,N_2694,N_2685);
nand U2712 (N_2712,N_2665,N_2658);
or U2713 (N_2713,N_2695,N_2696);
and U2714 (N_2714,N_2662,N_2681);
nand U2715 (N_2715,N_2689,N_2650);
and U2716 (N_2716,N_2688,N_2697);
nor U2717 (N_2717,N_2683,N_2674);
and U2718 (N_2718,N_2698,N_2661);
or U2719 (N_2719,N_2673,N_2699);
and U2720 (N_2720,N_2666,N_2655);
nand U2721 (N_2721,N_2680,N_2682);
nand U2722 (N_2722,N_2672,N_2676);
nand U2723 (N_2723,N_2667,N_2659);
nor U2724 (N_2724,N_2678,N_2654);
and U2725 (N_2725,N_2659,N_2680);
nor U2726 (N_2726,N_2666,N_2695);
or U2727 (N_2727,N_2660,N_2668);
nand U2728 (N_2728,N_2671,N_2672);
or U2729 (N_2729,N_2668,N_2680);
nand U2730 (N_2730,N_2676,N_2681);
nor U2731 (N_2731,N_2666,N_2674);
or U2732 (N_2732,N_2670,N_2679);
and U2733 (N_2733,N_2699,N_2676);
and U2734 (N_2734,N_2663,N_2662);
nand U2735 (N_2735,N_2691,N_2693);
nand U2736 (N_2736,N_2661,N_2686);
nand U2737 (N_2737,N_2663,N_2691);
or U2738 (N_2738,N_2690,N_2686);
nor U2739 (N_2739,N_2683,N_2693);
and U2740 (N_2740,N_2682,N_2676);
and U2741 (N_2741,N_2697,N_2692);
xnor U2742 (N_2742,N_2661,N_2679);
nor U2743 (N_2743,N_2666,N_2659);
and U2744 (N_2744,N_2690,N_2681);
or U2745 (N_2745,N_2684,N_2654);
or U2746 (N_2746,N_2692,N_2695);
nor U2747 (N_2747,N_2658,N_2667);
xor U2748 (N_2748,N_2688,N_2696);
nand U2749 (N_2749,N_2650,N_2677);
and U2750 (N_2750,N_2714,N_2721);
nand U2751 (N_2751,N_2703,N_2732);
nor U2752 (N_2752,N_2710,N_2735);
nor U2753 (N_2753,N_2746,N_2728);
nand U2754 (N_2754,N_2743,N_2711);
nor U2755 (N_2755,N_2704,N_2731);
nor U2756 (N_2756,N_2707,N_2744);
nor U2757 (N_2757,N_2737,N_2713);
or U2758 (N_2758,N_2701,N_2712);
nand U2759 (N_2759,N_2733,N_2700);
nand U2760 (N_2760,N_2738,N_2740);
or U2761 (N_2761,N_2725,N_2723);
and U2762 (N_2762,N_2742,N_2708);
nor U2763 (N_2763,N_2729,N_2739);
nor U2764 (N_2764,N_2734,N_2736);
and U2765 (N_2765,N_2716,N_2727);
or U2766 (N_2766,N_2719,N_2741);
and U2767 (N_2767,N_2747,N_2745);
nand U2768 (N_2768,N_2722,N_2702);
or U2769 (N_2769,N_2705,N_2720);
and U2770 (N_2770,N_2718,N_2730);
and U2771 (N_2771,N_2717,N_2715);
and U2772 (N_2772,N_2748,N_2726);
nor U2773 (N_2773,N_2709,N_2724);
nor U2774 (N_2774,N_2749,N_2706);
and U2775 (N_2775,N_2717,N_2700);
nand U2776 (N_2776,N_2739,N_2731);
nor U2777 (N_2777,N_2742,N_2726);
nor U2778 (N_2778,N_2701,N_2717);
or U2779 (N_2779,N_2732,N_2707);
nor U2780 (N_2780,N_2720,N_2738);
nand U2781 (N_2781,N_2708,N_2707);
nor U2782 (N_2782,N_2709,N_2708);
and U2783 (N_2783,N_2747,N_2739);
nor U2784 (N_2784,N_2736,N_2714);
nor U2785 (N_2785,N_2715,N_2705);
or U2786 (N_2786,N_2723,N_2730);
nor U2787 (N_2787,N_2718,N_2748);
nand U2788 (N_2788,N_2742,N_2705);
nor U2789 (N_2789,N_2748,N_2700);
nand U2790 (N_2790,N_2701,N_2747);
and U2791 (N_2791,N_2734,N_2723);
nand U2792 (N_2792,N_2723,N_2700);
nor U2793 (N_2793,N_2707,N_2719);
nand U2794 (N_2794,N_2704,N_2723);
or U2795 (N_2795,N_2746,N_2709);
nor U2796 (N_2796,N_2717,N_2739);
nand U2797 (N_2797,N_2748,N_2725);
or U2798 (N_2798,N_2719,N_2742);
and U2799 (N_2799,N_2713,N_2738);
and U2800 (N_2800,N_2781,N_2779);
nand U2801 (N_2801,N_2776,N_2790);
or U2802 (N_2802,N_2775,N_2773);
xor U2803 (N_2803,N_2766,N_2756);
or U2804 (N_2804,N_2789,N_2795);
nor U2805 (N_2805,N_2770,N_2778);
and U2806 (N_2806,N_2758,N_2771);
and U2807 (N_2807,N_2754,N_2796);
xor U2808 (N_2808,N_2791,N_2782);
or U2809 (N_2809,N_2799,N_2780);
nand U2810 (N_2810,N_2797,N_2769);
or U2811 (N_2811,N_2753,N_2772);
nor U2812 (N_2812,N_2786,N_2751);
or U2813 (N_2813,N_2783,N_2785);
and U2814 (N_2814,N_2764,N_2784);
and U2815 (N_2815,N_2752,N_2762);
nor U2816 (N_2816,N_2787,N_2792);
nand U2817 (N_2817,N_2761,N_2777);
and U2818 (N_2818,N_2765,N_2759);
xnor U2819 (N_2819,N_2788,N_2750);
or U2820 (N_2820,N_2774,N_2768);
and U2821 (N_2821,N_2757,N_2760);
nand U2822 (N_2822,N_2798,N_2755);
nand U2823 (N_2823,N_2793,N_2794);
nor U2824 (N_2824,N_2763,N_2767);
nor U2825 (N_2825,N_2752,N_2773);
nand U2826 (N_2826,N_2768,N_2798);
nor U2827 (N_2827,N_2760,N_2792);
and U2828 (N_2828,N_2757,N_2777);
or U2829 (N_2829,N_2762,N_2753);
and U2830 (N_2830,N_2771,N_2752);
nor U2831 (N_2831,N_2789,N_2752);
nand U2832 (N_2832,N_2764,N_2780);
nor U2833 (N_2833,N_2796,N_2760);
nor U2834 (N_2834,N_2789,N_2787);
nand U2835 (N_2835,N_2762,N_2794);
or U2836 (N_2836,N_2778,N_2786);
nor U2837 (N_2837,N_2791,N_2799);
or U2838 (N_2838,N_2784,N_2779);
and U2839 (N_2839,N_2763,N_2792);
nand U2840 (N_2840,N_2766,N_2798);
or U2841 (N_2841,N_2760,N_2791);
nor U2842 (N_2842,N_2761,N_2795);
and U2843 (N_2843,N_2776,N_2762);
and U2844 (N_2844,N_2783,N_2778);
nand U2845 (N_2845,N_2767,N_2792);
nor U2846 (N_2846,N_2750,N_2759);
nand U2847 (N_2847,N_2797,N_2784);
nand U2848 (N_2848,N_2783,N_2786);
or U2849 (N_2849,N_2772,N_2781);
and U2850 (N_2850,N_2835,N_2818);
or U2851 (N_2851,N_2802,N_2803);
nor U2852 (N_2852,N_2821,N_2810);
or U2853 (N_2853,N_2807,N_2813);
nand U2854 (N_2854,N_2828,N_2805);
nand U2855 (N_2855,N_2811,N_2846);
and U2856 (N_2856,N_2801,N_2838);
or U2857 (N_2857,N_2827,N_2814);
nand U2858 (N_2858,N_2831,N_2808);
or U2859 (N_2859,N_2840,N_2816);
and U2860 (N_2860,N_2812,N_2815);
nor U2861 (N_2861,N_2804,N_2829);
or U2862 (N_2862,N_2825,N_2832);
nor U2863 (N_2863,N_2822,N_2823);
nand U2864 (N_2864,N_2849,N_2834);
or U2865 (N_2865,N_2833,N_2809);
nand U2866 (N_2866,N_2836,N_2820);
or U2867 (N_2867,N_2817,N_2826);
nor U2868 (N_2868,N_2848,N_2843);
or U2869 (N_2869,N_2845,N_2842);
or U2870 (N_2870,N_2847,N_2830);
nor U2871 (N_2871,N_2824,N_2819);
nand U2872 (N_2872,N_2844,N_2837);
nor U2873 (N_2873,N_2841,N_2806);
nand U2874 (N_2874,N_2839,N_2800);
and U2875 (N_2875,N_2823,N_2821);
nand U2876 (N_2876,N_2838,N_2833);
or U2877 (N_2877,N_2816,N_2848);
nand U2878 (N_2878,N_2815,N_2831);
and U2879 (N_2879,N_2842,N_2800);
nor U2880 (N_2880,N_2813,N_2820);
nor U2881 (N_2881,N_2815,N_2825);
or U2882 (N_2882,N_2813,N_2834);
nand U2883 (N_2883,N_2804,N_2820);
nand U2884 (N_2884,N_2828,N_2835);
or U2885 (N_2885,N_2846,N_2842);
nor U2886 (N_2886,N_2817,N_2822);
and U2887 (N_2887,N_2841,N_2814);
nor U2888 (N_2888,N_2804,N_2837);
nand U2889 (N_2889,N_2848,N_2840);
nand U2890 (N_2890,N_2811,N_2835);
or U2891 (N_2891,N_2810,N_2826);
and U2892 (N_2892,N_2847,N_2837);
nor U2893 (N_2893,N_2813,N_2826);
and U2894 (N_2894,N_2817,N_2819);
nand U2895 (N_2895,N_2809,N_2844);
or U2896 (N_2896,N_2817,N_2843);
nor U2897 (N_2897,N_2827,N_2838);
and U2898 (N_2898,N_2802,N_2812);
and U2899 (N_2899,N_2838,N_2817);
nand U2900 (N_2900,N_2853,N_2893);
nand U2901 (N_2901,N_2864,N_2857);
nand U2902 (N_2902,N_2852,N_2858);
or U2903 (N_2903,N_2891,N_2861);
or U2904 (N_2904,N_2882,N_2877);
or U2905 (N_2905,N_2883,N_2867);
or U2906 (N_2906,N_2863,N_2874);
nand U2907 (N_2907,N_2855,N_2854);
nand U2908 (N_2908,N_2879,N_2887);
nand U2909 (N_2909,N_2881,N_2856);
nor U2910 (N_2910,N_2860,N_2869);
or U2911 (N_2911,N_2851,N_2884);
nand U2912 (N_2912,N_2871,N_2896);
nand U2913 (N_2913,N_2894,N_2870);
or U2914 (N_2914,N_2866,N_2892);
nand U2915 (N_2915,N_2895,N_2885);
or U2916 (N_2916,N_2865,N_2888);
nand U2917 (N_2917,N_2880,N_2862);
nor U2918 (N_2918,N_2875,N_2872);
or U2919 (N_2919,N_2859,N_2876);
or U2920 (N_2920,N_2897,N_2898);
and U2921 (N_2921,N_2889,N_2873);
or U2922 (N_2922,N_2878,N_2890);
nand U2923 (N_2923,N_2899,N_2868);
or U2924 (N_2924,N_2886,N_2850);
or U2925 (N_2925,N_2871,N_2879);
nand U2926 (N_2926,N_2853,N_2864);
and U2927 (N_2927,N_2860,N_2872);
nand U2928 (N_2928,N_2878,N_2879);
nand U2929 (N_2929,N_2896,N_2894);
or U2930 (N_2930,N_2852,N_2881);
nand U2931 (N_2931,N_2897,N_2873);
nor U2932 (N_2932,N_2874,N_2857);
nand U2933 (N_2933,N_2891,N_2892);
or U2934 (N_2934,N_2885,N_2850);
and U2935 (N_2935,N_2897,N_2855);
nor U2936 (N_2936,N_2853,N_2872);
nand U2937 (N_2937,N_2880,N_2860);
or U2938 (N_2938,N_2874,N_2888);
nand U2939 (N_2939,N_2869,N_2885);
nor U2940 (N_2940,N_2888,N_2884);
or U2941 (N_2941,N_2864,N_2855);
nand U2942 (N_2942,N_2876,N_2863);
nor U2943 (N_2943,N_2854,N_2888);
and U2944 (N_2944,N_2862,N_2871);
and U2945 (N_2945,N_2873,N_2884);
or U2946 (N_2946,N_2865,N_2863);
and U2947 (N_2947,N_2887,N_2866);
or U2948 (N_2948,N_2880,N_2886);
or U2949 (N_2949,N_2898,N_2892);
and U2950 (N_2950,N_2939,N_2911);
nor U2951 (N_2951,N_2942,N_2902);
and U2952 (N_2952,N_2930,N_2910);
and U2953 (N_2953,N_2937,N_2945);
nor U2954 (N_2954,N_2940,N_2923);
and U2955 (N_2955,N_2903,N_2912);
or U2956 (N_2956,N_2949,N_2909);
nand U2957 (N_2957,N_2900,N_2914);
and U2958 (N_2958,N_2928,N_2905);
nor U2959 (N_2959,N_2929,N_2904);
or U2960 (N_2960,N_2944,N_2917);
or U2961 (N_2961,N_2906,N_2922);
or U2962 (N_2962,N_2931,N_2915);
or U2963 (N_2963,N_2936,N_2925);
or U2964 (N_2964,N_2901,N_2947);
nand U2965 (N_2965,N_2934,N_2946);
and U2966 (N_2966,N_2916,N_2935);
nor U2967 (N_2967,N_2919,N_2932);
and U2968 (N_2968,N_2908,N_2948);
nand U2969 (N_2969,N_2927,N_2941);
and U2970 (N_2970,N_2907,N_2918);
or U2971 (N_2971,N_2924,N_2943);
nor U2972 (N_2972,N_2938,N_2920);
and U2973 (N_2973,N_2913,N_2921);
nand U2974 (N_2974,N_2926,N_2933);
nor U2975 (N_2975,N_2909,N_2936);
nand U2976 (N_2976,N_2944,N_2942);
or U2977 (N_2977,N_2948,N_2940);
or U2978 (N_2978,N_2936,N_2910);
and U2979 (N_2979,N_2916,N_2944);
and U2980 (N_2980,N_2902,N_2934);
nand U2981 (N_2981,N_2912,N_2933);
nor U2982 (N_2982,N_2904,N_2900);
or U2983 (N_2983,N_2908,N_2900);
or U2984 (N_2984,N_2949,N_2928);
or U2985 (N_2985,N_2946,N_2922);
or U2986 (N_2986,N_2926,N_2920);
and U2987 (N_2987,N_2942,N_2936);
and U2988 (N_2988,N_2929,N_2924);
nand U2989 (N_2989,N_2946,N_2940);
nand U2990 (N_2990,N_2910,N_2937);
nand U2991 (N_2991,N_2947,N_2917);
or U2992 (N_2992,N_2911,N_2925);
nand U2993 (N_2993,N_2941,N_2948);
nor U2994 (N_2994,N_2907,N_2917);
nand U2995 (N_2995,N_2932,N_2936);
nor U2996 (N_2996,N_2930,N_2900);
nor U2997 (N_2997,N_2920,N_2929);
and U2998 (N_2998,N_2924,N_2911);
or U2999 (N_2999,N_2936,N_2902);
and UO_0 (O_0,N_2983,N_2958);
nor UO_1 (O_1,N_2961,N_2970);
nor UO_2 (O_2,N_2965,N_2978);
or UO_3 (O_3,N_2950,N_2967);
or UO_4 (O_4,N_2952,N_2962);
nor UO_5 (O_5,N_2968,N_2982);
or UO_6 (O_6,N_2997,N_2992);
and UO_7 (O_7,N_2975,N_2986);
nor UO_8 (O_8,N_2953,N_2984);
nor UO_9 (O_9,N_2951,N_2990);
nor UO_10 (O_10,N_2976,N_2998);
nor UO_11 (O_11,N_2980,N_2994);
or UO_12 (O_12,N_2972,N_2966);
nand UO_13 (O_13,N_2988,N_2993);
and UO_14 (O_14,N_2973,N_2956);
and UO_15 (O_15,N_2969,N_2985);
nand UO_16 (O_16,N_2957,N_2989);
nor UO_17 (O_17,N_2995,N_2954);
nor UO_18 (O_18,N_2977,N_2981);
xor UO_19 (O_19,N_2955,N_2964);
or UO_20 (O_20,N_2960,N_2987);
and UO_21 (O_21,N_2999,N_2959);
nor UO_22 (O_22,N_2996,N_2974);
and UO_23 (O_23,N_2971,N_2991);
nor UO_24 (O_24,N_2963,N_2979);
nand UO_25 (O_25,N_2995,N_2986);
nor UO_26 (O_26,N_2963,N_2990);
or UO_27 (O_27,N_2987,N_2959);
or UO_28 (O_28,N_2982,N_2991);
and UO_29 (O_29,N_2990,N_2986);
nor UO_30 (O_30,N_2974,N_2984);
nand UO_31 (O_31,N_2995,N_2964);
nor UO_32 (O_32,N_2954,N_2982);
nor UO_33 (O_33,N_2998,N_2977);
nor UO_34 (O_34,N_2975,N_2989);
nand UO_35 (O_35,N_2974,N_2950);
and UO_36 (O_36,N_2957,N_2999);
and UO_37 (O_37,N_2996,N_2955);
or UO_38 (O_38,N_2958,N_2984);
and UO_39 (O_39,N_2958,N_2998);
or UO_40 (O_40,N_2967,N_2964);
and UO_41 (O_41,N_2966,N_2953);
and UO_42 (O_42,N_2954,N_2959);
nand UO_43 (O_43,N_2979,N_2985);
or UO_44 (O_44,N_2978,N_2959);
and UO_45 (O_45,N_2952,N_2954);
nor UO_46 (O_46,N_2981,N_2968);
nor UO_47 (O_47,N_2999,N_2997);
or UO_48 (O_48,N_2997,N_2970);
or UO_49 (O_49,N_2994,N_2961);
nand UO_50 (O_50,N_2995,N_2952);
nand UO_51 (O_51,N_2956,N_2960);
and UO_52 (O_52,N_2982,N_2996);
nor UO_53 (O_53,N_2957,N_2953);
nor UO_54 (O_54,N_2970,N_2985);
and UO_55 (O_55,N_2952,N_2961);
nor UO_56 (O_56,N_2962,N_2965);
or UO_57 (O_57,N_2967,N_2977);
nand UO_58 (O_58,N_2951,N_2997);
nand UO_59 (O_59,N_2951,N_2987);
or UO_60 (O_60,N_2984,N_2959);
nand UO_61 (O_61,N_2951,N_2976);
nand UO_62 (O_62,N_2984,N_2955);
nand UO_63 (O_63,N_2997,N_2995);
nand UO_64 (O_64,N_2952,N_2987);
and UO_65 (O_65,N_2984,N_2970);
nor UO_66 (O_66,N_2954,N_2973);
and UO_67 (O_67,N_2999,N_2960);
or UO_68 (O_68,N_2952,N_2970);
or UO_69 (O_69,N_2993,N_2983);
and UO_70 (O_70,N_2985,N_2989);
nand UO_71 (O_71,N_2997,N_2965);
and UO_72 (O_72,N_2983,N_2996);
or UO_73 (O_73,N_2952,N_2977);
and UO_74 (O_74,N_2983,N_2982);
nand UO_75 (O_75,N_2997,N_2955);
or UO_76 (O_76,N_2975,N_2971);
nor UO_77 (O_77,N_2988,N_2986);
or UO_78 (O_78,N_2989,N_2950);
nor UO_79 (O_79,N_2952,N_2963);
nand UO_80 (O_80,N_2973,N_2999);
nor UO_81 (O_81,N_2966,N_2973);
nand UO_82 (O_82,N_2968,N_2955);
xnor UO_83 (O_83,N_2951,N_2960);
or UO_84 (O_84,N_2996,N_2989);
and UO_85 (O_85,N_2960,N_2950);
or UO_86 (O_86,N_2979,N_2960);
nand UO_87 (O_87,N_2999,N_2969);
nand UO_88 (O_88,N_2981,N_2979);
and UO_89 (O_89,N_2974,N_2958);
and UO_90 (O_90,N_2997,N_2974);
and UO_91 (O_91,N_2999,N_2967);
or UO_92 (O_92,N_2972,N_2996);
nand UO_93 (O_93,N_2971,N_2970);
and UO_94 (O_94,N_2982,N_2969);
or UO_95 (O_95,N_2963,N_2955);
nor UO_96 (O_96,N_2967,N_2963);
nand UO_97 (O_97,N_2993,N_2985);
nand UO_98 (O_98,N_2990,N_2984);
or UO_99 (O_99,N_2951,N_2958);
nand UO_100 (O_100,N_2970,N_2956);
nand UO_101 (O_101,N_2982,N_2974);
nor UO_102 (O_102,N_2970,N_2998);
and UO_103 (O_103,N_2995,N_2979);
and UO_104 (O_104,N_2983,N_2956);
or UO_105 (O_105,N_2995,N_2970);
nor UO_106 (O_106,N_2996,N_2984);
and UO_107 (O_107,N_2973,N_2988);
nand UO_108 (O_108,N_2982,N_2987);
and UO_109 (O_109,N_2987,N_2977);
or UO_110 (O_110,N_2990,N_2994);
nor UO_111 (O_111,N_2966,N_2983);
nor UO_112 (O_112,N_2978,N_2974);
or UO_113 (O_113,N_2969,N_2950);
nand UO_114 (O_114,N_2974,N_2965);
and UO_115 (O_115,N_2975,N_2988);
nor UO_116 (O_116,N_2955,N_2985);
and UO_117 (O_117,N_2984,N_2979);
nor UO_118 (O_118,N_2995,N_2961);
nand UO_119 (O_119,N_2983,N_2979);
nor UO_120 (O_120,N_2969,N_2980);
nand UO_121 (O_121,N_2974,N_2971);
and UO_122 (O_122,N_2978,N_2996);
and UO_123 (O_123,N_2958,N_2982);
and UO_124 (O_124,N_2977,N_2997);
nor UO_125 (O_125,N_2983,N_2969);
or UO_126 (O_126,N_2998,N_2980);
or UO_127 (O_127,N_2997,N_2960);
and UO_128 (O_128,N_2963,N_2957);
and UO_129 (O_129,N_2966,N_2959);
nand UO_130 (O_130,N_2968,N_2984);
or UO_131 (O_131,N_2982,N_2963);
nor UO_132 (O_132,N_2990,N_2957);
nand UO_133 (O_133,N_2971,N_2973);
nor UO_134 (O_134,N_2953,N_2994);
nor UO_135 (O_135,N_2998,N_2995);
nor UO_136 (O_136,N_2971,N_2950);
or UO_137 (O_137,N_2973,N_2968);
nor UO_138 (O_138,N_2974,N_2968);
nand UO_139 (O_139,N_2956,N_2985);
nor UO_140 (O_140,N_2979,N_2973);
and UO_141 (O_141,N_2964,N_2986);
or UO_142 (O_142,N_2989,N_2987);
nor UO_143 (O_143,N_2955,N_2981);
nor UO_144 (O_144,N_2987,N_2998);
or UO_145 (O_145,N_2982,N_2986);
nor UO_146 (O_146,N_2958,N_2950);
and UO_147 (O_147,N_2966,N_2985);
nor UO_148 (O_148,N_2987,N_2990);
or UO_149 (O_149,N_2998,N_2964);
nor UO_150 (O_150,N_2992,N_2977);
and UO_151 (O_151,N_2969,N_2951);
nand UO_152 (O_152,N_2993,N_2976);
and UO_153 (O_153,N_2976,N_2969);
nor UO_154 (O_154,N_2961,N_2964);
and UO_155 (O_155,N_2986,N_2962);
nand UO_156 (O_156,N_2953,N_2955);
nor UO_157 (O_157,N_2995,N_2975);
and UO_158 (O_158,N_2987,N_2991);
nor UO_159 (O_159,N_2975,N_2973);
nor UO_160 (O_160,N_2985,N_2962);
and UO_161 (O_161,N_2992,N_2988);
nand UO_162 (O_162,N_2971,N_2983);
nand UO_163 (O_163,N_2990,N_2989);
and UO_164 (O_164,N_2996,N_2994);
nand UO_165 (O_165,N_2983,N_2997);
nand UO_166 (O_166,N_2960,N_2992);
nand UO_167 (O_167,N_2960,N_2976);
nand UO_168 (O_168,N_2951,N_2954);
nand UO_169 (O_169,N_2953,N_2997);
and UO_170 (O_170,N_2975,N_2955);
and UO_171 (O_171,N_2974,N_2983);
nor UO_172 (O_172,N_2963,N_2985);
and UO_173 (O_173,N_2969,N_2997);
or UO_174 (O_174,N_2966,N_2984);
or UO_175 (O_175,N_2978,N_2968);
or UO_176 (O_176,N_2982,N_2972);
and UO_177 (O_177,N_2950,N_2954);
nand UO_178 (O_178,N_2984,N_2973);
and UO_179 (O_179,N_2964,N_2973);
nand UO_180 (O_180,N_2958,N_2969);
nand UO_181 (O_181,N_2974,N_2957);
or UO_182 (O_182,N_2986,N_2985);
nand UO_183 (O_183,N_2995,N_2950);
nor UO_184 (O_184,N_2994,N_2995);
nand UO_185 (O_185,N_2998,N_2954);
and UO_186 (O_186,N_2974,N_2991);
nor UO_187 (O_187,N_2973,N_2986);
and UO_188 (O_188,N_2963,N_2994);
nor UO_189 (O_189,N_2950,N_2990);
and UO_190 (O_190,N_2964,N_2958);
nor UO_191 (O_191,N_2994,N_2972);
nand UO_192 (O_192,N_2978,N_2993);
and UO_193 (O_193,N_2961,N_2956);
or UO_194 (O_194,N_2990,N_2952);
or UO_195 (O_195,N_2966,N_2975);
nor UO_196 (O_196,N_2956,N_2975);
nand UO_197 (O_197,N_2957,N_2988);
and UO_198 (O_198,N_2985,N_2998);
nor UO_199 (O_199,N_2957,N_2950);
or UO_200 (O_200,N_2990,N_2970);
and UO_201 (O_201,N_2970,N_2965);
or UO_202 (O_202,N_2974,N_2955);
nor UO_203 (O_203,N_2992,N_2986);
nand UO_204 (O_204,N_2977,N_2982);
and UO_205 (O_205,N_2964,N_2988);
and UO_206 (O_206,N_2959,N_2970);
nor UO_207 (O_207,N_2951,N_2955);
nor UO_208 (O_208,N_2986,N_2977);
and UO_209 (O_209,N_2986,N_2989);
nand UO_210 (O_210,N_2960,N_2995);
nand UO_211 (O_211,N_2953,N_2990);
nor UO_212 (O_212,N_2963,N_2961);
nor UO_213 (O_213,N_2980,N_2991);
nor UO_214 (O_214,N_2951,N_2974);
or UO_215 (O_215,N_2974,N_2963);
nor UO_216 (O_216,N_2998,N_2978);
and UO_217 (O_217,N_2986,N_2970);
and UO_218 (O_218,N_2983,N_2989);
or UO_219 (O_219,N_2991,N_2996);
nand UO_220 (O_220,N_2989,N_2959);
or UO_221 (O_221,N_2953,N_2993);
and UO_222 (O_222,N_2994,N_2965);
nand UO_223 (O_223,N_2962,N_2950);
nor UO_224 (O_224,N_2956,N_2998);
or UO_225 (O_225,N_2979,N_2987);
or UO_226 (O_226,N_2978,N_2983);
nand UO_227 (O_227,N_2990,N_2979);
nor UO_228 (O_228,N_2992,N_2972);
and UO_229 (O_229,N_2956,N_2954);
nor UO_230 (O_230,N_2960,N_2974);
nand UO_231 (O_231,N_2968,N_2950);
nor UO_232 (O_232,N_2971,N_2988);
nor UO_233 (O_233,N_2957,N_2959);
nor UO_234 (O_234,N_2957,N_2970);
nor UO_235 (O_235,N_2957,N_2961);
and UO_236 (O_236,N_2996,N_2950);
xnor UO_237 (O_237,N_2985,N_2957);
and UO_238 (O_238,N_2999,N_2995);
and UO_239 (O_239,N_2960,N_2978);
and UO_240 (O_240,N_2993,N_2977);
and UO_241 (O_241,N_2996,N_2995);
and UO_242 (O_242,N_2972,N_2989);
nand UO_243 (O_243,N_2987,N_2964);
and UO_244 (O_244,N_2990,N_2971);
nand UO_245 (O_245,N_2984,N_2988);
or UO_246 (O_246,N_2984,N_2999);
nor UO_247 (O_247,N_2975,N_2992);
or UO_248 (O_248,N_2997,N_2988);
or UO_249 (O_249,N_2967,N_2984);
nor UO_250 (O_250,N_2962,N_2988);
nor UO_251 (O_251,N_2991,N_2983);
and UO_252 (O_252,N_2954,N_2986);
or UO_253 (O_253,N_2990,N_2969);
nor UO_254 (O_254,N_2985,N_2999);
or UO_255 (O_255,N_2971,N_2968);
and UO_256 (O_256,N_2956,N_2991);
and UO_257 (O_257,N_2979,N_2999);
nand UO_258 (O_258,N_2971,N_2956);
nor UO_259 (O_259,N_2992,N_2973);
nand UO_260 (O_260,N_2971,N_2951);
nand UO_261 (O_261,N_2960,N_2990);
and UO_262 (O_262,N_2965,N_2971);
or UO_263 (O_263,N_2976,N_2959);
and UO_264 (O_264,N_2992,N_2951);
and UO_265 (O_265,N_2989,N_2963);
or UO_266 (O_266,N_2987,N_2986);
or UO_267 (O_267,N_2986,N_2978);
nand UO_268 (O_268,N_2975,N_2964);
and UO_269 (O_269,N_2966,N_2991);
or UO_270 (O_270,N_2964,N_2972);
nor UO_271 (O_271,N_2958,N_2977);
nor UO_272 (O_272,N_2951,N_2979);
and UO_273 (O_273,N_2968,N_2962);
nor UO_274 (O_274,N_2953,N_2963);
or UO_275 (O_275,N_2965,N_2980);
nand UO_276 (O_276,N_2994,N_2978);
nand UO_277 (O_277,N_2956,N_2980);
or UO_278 (O_278,N_2993,N_2966);
nand UO_279 (O_279,N_2950,N_2997);
or UO_280 (O_280,N_2970,N_2964);
or UO_281 (O_281,N_2957,N_2973);
or UO_282 (O_282,N_2955,N_2995);
nand UO_283 (O_283,N_2980,N_2972);
nand UO_284 (O_284,N_2991,N_2990);
and UO_285 (O_285,N_2974,N_2990);
nand UO_286 (O_286,N_2971,N_2963);
and UO_287 (O_287,N_2999,N_2966);
nor UO_288 (O_288,N_2975,N_2981);
nand UO_289 (O_289,N_2959,N_2979);
and UO_290 (O_290,N_2989,N_2988);
or UO_291 (O_291,N_2952,N_2986);
nor UO_292 (O_292,N_2975,N_2976);
nor UO_293 (O_293,N_2968,N_2986);
nand UO_294 (O_294,N_2953,N_2987);
and UO_295 (O_295,N_2995,N_2988);
nor UO_296 (O_296,N_2961,N_2968);
and UO_297 (O_297,N_2978,N_2981);
nor UO_298 (O_298,N_2977,N_2959);
nor UO_299 (O_299,N_2955,N_2989);
nand UO_300 (O_300,N_2959,N_2965);
nand UO_301 (O_301,N_2971,N_2984);
nor UO_302 (O_302,N_2995,N_2980);
nor UO_303 (O_303,N_2975,N_2978);
and UO_304 (O_304,N_2970,N_2992);
nor UO_305 (O_305,N_2951,N_2968);
or UO_306 (O_306,N_2999,N_2983);
and UO_307 (O_307,N_2978,N_2979);
or UO_308 (O_308,N_2967,N_2968);
or UO_309 (O_309,N_2951,N_2956);
and UO_310 (O_310,N_2985,N_2994);
nor UO_311 (O_311,N_2968,N_2985);
nor UO_312 (O_312,N_2971,N_2981);
nand UO_313 (O_313,N_2968,N_2954);
nand UO_314 (O_314,N_2960,N_2985);
or UO_315 (O_315,N_2967,N_2990);
nand UO_316 (O_316,N_2982,N_2959);
xnor UO_317 (O_317,N_2959,N_2994);
nor UO_318 (O_318,N_2998,N_2969);
nand UO_319 (O_319,N_2999,N_2994);
or UO_320 (O_320,N_2975,N_2969);
and UO_321 (O_321,N_2958,N_2994);
nor UO_322 (O_322,N_2976,N_2950);
and UO_323 (O_323,N_2973,N_2982);
nand UO_324 (O_324,N_2984,N_2993);
nor UO_325 (O_325,N_2975,N_2961);
or UO_326 (O_326,N_2997,N_2979);
nor UO_327 (O_327,N_2952,N_2974);
and UO_328 (O_328,N_2952,N_2971);
nand UO_329 (O_329,N_2962,N_2979);
or UO_330 (O_330,N_2999,N_2962);
or UO_331 (O_331,N_2988,N_2994);
nand UO_332 (O_332,N_2981,N_2976);
and UO_333 (O_333,N_2960,N_2982);
nand UO_334 (O_334,N_2980,N_2996);
nand UO_335 (O_335,N_2996,N_2990);
nor UO_336 (O_336,N_2965,N_2993);
and UO_337 (O_337,N_2977,N_2960);
nand UO_338 (O_338,N_2992,N_2964);
nand UO_339 (O_339,N_2985,N_2980);
nor UO_340 (O_340,N_2976,N_2989);
nor UO_341 (O_341,N_2996,N_2986);
or UO_342 (O_342,N_2962,N_2984);
and UO_343 (O_343,N_2977,N_2974);
nor UO_344 (O_344,N_2975,N_2950);
nand UO_345 (O_345,N_2989,N_2969);
nand UO_346 (O_346,N_2995,N_2971);
or UO_347 (O_347,N_2953,N_2954);
nor UO_348 (O_348,N_2976,N_2982);
or UO_349 (O_349,N_2957,N_2969);
nor UO_350 (O_350,N_2968,N_2996);
nor UO_351 (O_351,N_2976,N_2955);
or UO_352 (O_352,N_2963,N_2958);
nor UO_353 (O_353,N_2979,N_2986);
nand UO_354 (O_354,N_2959,N_2996);
or UO_355 (O_355,N_2971,N_2964);
and UO_356 (O_356,N_2984,N_2983);
or UO_357 (O_357,N_2973,N_2987);
or UO_358 (O_358,N_2962,N_2972);
nand UO_359 (O_359,N_2959,N_2950);
nand UO_360 (O_360,N_2955,N_2957);
or UO_361 (O_361,N_2972,N_2955);
and UO_362 (O_362,N_2997,N_2972);
and UO_363 (O_363,N_2967,N_2956);
nand UO_364 (O_364,N_2995,N_2978);
nor UO_365 (O_365,N_2986,N_2998);
nor UO_366 (O_366,N_2958,N_2988);
nor UO_367 (O_367,N_2962,N_2959);
nand UO_368 (O_368,N_2967,N_2992);
or UO_369 (O_369,N_2995,N_2966);
nand UO_370 (O_370,N_2980,N_2981);
or UO_371 (O_371,N_2995,N_2985);
nor UO_372 (O_372,N_2970,N_2987);
nor UO_373 (O_373,N_2951,N_2959);
or UO_374 (O_374,N_2953,N_2988);
or UO_375 (O_375,N_2984,N_2980);
nand UO_376 (O_376,N_2967,N_2974);
or UO_377 (O_377,N_2955,N_2986);
nor UO_378 (O_378,N_2988,N_2966);
nor UO_379 (O_379,N_2963,N_2987);
and UO_380 (O_380,N_2980,N_2977);
nand UO_381 (O_381,N_2992,N_2995);
and UO_382 (O_382,N_2952,N_2960);
nor UO_383 (O_383,N_2962,N_2961);
nand UO_384 (O_384,N_2977,N_2996);
or UO_385 (O_385,N_2984,N_2972);
xnor UO_386 (O_386,N_2965,N_2975);
and UO_387 (O_387,N_2992,N_2983);
and UO_388 (O_388,N_2998,N_2983);
xnor UO_389 (O_389,N_2955,N_2992);
and UO_390 (O_390,N_2960,N_2975);
nor UO_391 (O_391,N_2979,N_2996);
and UO_392 (O_392,N_2951,N_2999);
nor UO_393 (O_393,N_2965,N_2956);
and UO_394 (O_394,N_2961,N_2969);
nand UO_395 (O_395,N_2981,N_2965);
nor UO_396 (O_396,N_2968,N_2989);
xor UO_397 (O_397,N_2975,N_2967);
or UO_398 (O_398,N_2968,N_2977);
and UO_399 (O_399,N_2968,N_2979);
nor UO_400 (O_400,N_2957,N_2980);
nor UO_401 (O_401,N_2992,N_2996);
and UO_402 (O_402,N_2970,N_2976);
nand UO_403 (O_403,N_2960,N_2959);
or UO_404 (O_404,N_2975,N_2968);
nor UO_405 (O_405,N_2961,N_2992);
or UO_406 (O_406,N_2968,N_2991);
or UO_407 (O_407,N_2983,N_2965);
or UO_408 (O_408,N_2978,N_2971);
nand UO_409 (O_409,N_2984,N_2977);
and UO_410 (O_410,N_2981,N_2950);
nor UO_411 (O_411,N_2974,N_2987);
and UO_412 (O_412,N_2957,N_2986);
or UO_413 (O_413,N_2954,N_2977);
nor UO_414 (O_414,N_2965,N_2979);
and UO_415 (O_415,N_2959,N_2963);
nand UO_416 (O_416,N_2966,N_2992);
nand UO_417 (O_417,N_2957,N_2994);
nor UO_418 (O_418,N_2968,N_2956);
nor UO_419 (O_419,N_2951,N_2967);
nand UO_420 (O_420,N_2964,N_2984);
or UO_421 (O_421,N_2969,N_2970);
nand UO_422 (O_422,N_2991,N_2994);
and UO_423 (O_423,N_2969,N_2974);
and UO_424 (O_424,N_2982,N_2979);
or UO_425 (O_425,N_2966,N_2970);
nand UO_426 (O_426,N_2992,N_2965);
or UO_427 (O_427,N_2991,N_2998);
nor UO_428 (O_428,N_2999,N_2987);
nor UO_429 (O_429,N_2954,N_2999);
nor UO_430 (O_430,N_2985,N_2954);
xor UO_431 (O_431,N_2972,N_2968);
or UO_432 (O_432,N_2965,N_2961);
nand UO_433 (O_433,N_2954,N_2958);
or UO_434 (O_434,N_2961,N_2966);
and UO_435 (O_435,N_2976,N_2984);
nor UO_436 (O_436,N_2962,N_2987);
and UO_437 (O_437,N_2951,N_2988);
or UO_438 (O_438,N_2956,N_2986);
and UO_439 (O_439,N_2993,N_2995);
or UO_440 (O_440,N_2963,N_2995);
nand UO_441 (O_441,N_2971,N_2986);
nor UO_442 (O_442,N_2982,N_2975);
xor UO_443 (O_443,N_2987,N_2983);
and UO_444 (O_444,N_2950,N_2979);
nand UO_445 (O_445,N_2975,N_2951);
or UO_446 (O_446,N_2980,N_2993);
nor UO_447 (O_447,N_2987,N_2971);
nor UO_448 (O_448,N_2954,N_2979);
or UO_449 (O_449,N_2962,N_2957);
nand UO_450 (O_450,N_2978,N_2989);
and UO_451 (O_451,N_2999,N_2972);
or UO_452 (O_452,N_2973,N_2996);
and UO_453 (O_453,N_2962,N_2960);
or UO_454 (O_454,N_2979,N_2988);
and UO_455 (O_455,N_2951,N_2978);
nor UO_456 (O_456,N_2991,N_2973);
nor UO_457 (O_457,N_2988,N_2969);
nor UO_458 (O_458,N_2964,N_2993);
nor UO_459 (O_459,N_2983,N_2955);
nor UO_460 (O_460,N_2990,N_2975);
nand UO_461 (O_461,N_2991,N_2954);
or UO_462 (O_462,N_2970,N_2981);
and UO_463 (O_463,N_2969,N_2978);
and UO_464 (O_464,N_2963,N_2976);
nand UO_465 (O_465,N_2955,N_2960);
nand UO_466 (O_466,N_2993,N_2961);
nand UO_467 (O_467,N_2950,N_2966);
nand UO_468 (O_468,N_2981,N_2963);
nor UO_469 (O_469,N_2962,N_2958);
and UO_470 (O_470,N_2996,N_2951);
nor UO_471 (O_471,N_2993,N_2989);
or UO_472 (O_472,N_2962,N_2955);
or UO_473 (O_473,N_2958,N_2980);
nand UO_474 (O_474,N_2991,N_2997);
or UO_475 (O_475,N_2977,N_2999);
nand UO_476 (O_476,N_2957,N_2951);
or UO_477 (O_477,N_2968,N_2953);
nand UO_478 (O_478,N_2973,N_2950);
nor UO_479 (O_479,N_2990,N_2985);
or UO_480 (O_480,N_2955,N_2969);
nand UO_481 (O_481,N_2987,N_2993);
and UO_482 (O_482,N_2952,N_2993);
nand UO_483 (O_483,N_2984,N_2957);
nor UO_484 (O_484,N_2983,N_2981);
or UO_485 (O_485,N_2977,N_2961);
or UO_486 (O_486,N_2960,N_2972);
nor UO_487 (O_487,N_2990,N_2962);
nor UO_488 (O_488,N_2976,N_2962);
nand UO_489 (O_489,N_2990,N_2955);
and UO_490 (O_490,N_2976,N_2956);
nor UO_491 (O_491,N_2972,N_2953);
nor UO_492 (O_492,N_2968,N_2987);
nor UO_493 (O_493,N_2974,N_2976);
nor UO_494 (O_494,N_2993,N_2994);
nand UO_495 (O_495,N_2985,N_2988);
or UO_496 (O_496,N_2968,N_2964);
nand UO_497 (O_497,N_2985,N_2992);
or UO_498 (O_498,N_2958,N_2968);
and UO_499 (O_499,N_2988,N_2952);
endmodule