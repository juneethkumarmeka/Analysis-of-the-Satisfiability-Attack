module basic_500_3000_500_50_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_23,In_89);
or U1 (N_1,In_352,In_270);
nor U2 (N_2,In_484,In_176);
nor U3 (N_3,In_34,In_340);
and U4 (N_4,In_373,In_372);
and U5 (N_5,In_240,In_108);
and U6 (N_6,In_364,In_298);
nand U7 (N_7,In_274,In_279);
and U8 (N_8,In_113,In_162);
nand U9 (N_9,In_343,In_407);
nand U10 (N_10,In_62,In_481);
or U11 (N_11,In_130,In_151);
and U12 (N_12,In_102,In_485);
nor U13 (N_13,In_308,In_375);
or U14 (N_14,In_290,In_150);
or U15 (N_15,In_207,In_88);
and U16 (N_16,In_280,In_226);
and U17 (N_17,In_365,In_330);
nor U18 (N_18,In_224,In_15);
nor U19 (N_19,In_75,In_216);
and U20 (N_20,In_268,In_237);
or U21 (N_21,In_106,In_384);
or U22 (N_22,In_492,In_38);
or U23 (N_23,In_49,In_295);
nand U24 (N_24,In_168,In_21);
nand U25 (N_25,In_129,In_263);
nor U26 (N_26,In_190,In_385);
nor U27 (N_27,In_149,In_46);
and U28 (N_28,In_284,In_164);
nand U29 (N_29,In_60,In_70);
nor U30 (N_30,In_173,In_366);
or U31 (N_31,In_73,In_29);
nand U32 (N_32,In_165,In_497);
and U33 (N_33,In_255,In_14);
and U34 (N_34,In_401,In_71);
nand U35 (N_35,In_12,In_256);
or U36 (N_36,In_454,In_283);
and U37 (N_37,In_86,In_369);
or U38 (N_38,In_241,In_194);
nand U39 (N_39,In_299,In_235);
and U40 (N_40,In_178,In_473);
and U41 (N_41,In_97,In_7);
nor U42 (N_42,In_467,In_486);
nand U43 (N_43,In_309,In_30);
nor U44 (N_44,In_57,In_192);
and U45 (N_45,In_383,In_8);
nand U46 (N_46,In_121,In_348);
nor U47 (N_47,In_307,In_482);
nor U48 (N_48,In_193,In_6);
or U49 (N_49,In_41,In_291);
or U50 (N_50,In_425,In_206);
and U51 (N_51,In_344,In_58);
or U52 (N_52,In_297,In_402);
nor U53 (N_53,In_212,In_392);
or U54 (N_54,In_345,In_25);
nand U55 (N_55,In_128,In_154);
and U56 (N_56,In_431,In_438);
or U57 (N_57,In_358,In_213);
and U58 (N_58,In_488,In_3);
nand U59 (N_59,In_219,In_91);
nor U60 (N_60,In_257,N_57);
nand U61 (N_61,In_109,In_361);
and U62 (N_62,In_227,In_363);
nand U63 (N_63,In_144,N_51);
nand U64 (N_64,In_292,N_6);
or U65 (N_65,In_273,In_107);
nor U66 (N_66,In_76,In_323);
or U67 (N_67,In_447,N_10);
nand U68 (N_68,In_248,In_136);
or U69 (N_69,In_67,In_215);
or U70 (N_70,N_32,N_23);
nand U71 (N_71,In_317,In_288);
nand U72 (N_72,In_305,In_245);
or U73 (N_73,In_155,In_196);
and U74 (N_74,In_301,In_259);
and U75 (N_75,In_205,In_440);
nor U76 (N_76,In_261,In_442);
or U77 (N_77,In_478,In_35);
nor U78 (N_78,In_477,In_499);
nand U79 (N_79,N_19,In_443);
nor U80 (N_80,In_156,In_479);
or U81 (N_81,In_388,In_430);
nand U82 (N_82,In_476,In_448);
or U83 (N_83,In_233,In_318);
or U84 (N_84,In_355,In_230);
or U85 (N_85,In_396,In_329);
or U86 (N_86,In_40,In_174);
nor U87 (N_87,In_445,In_169);
and U88 (N_88,In_367,N_9);
or U89 (N_89,In_72,In_428);
nor U90 (N_90,In_455,In_390);
nand U91 (N_91,N_20,In_487);
nor U92 (N_92,In_313,In_422);
nand U93 (N_93,In_350,In_44);
or U94 (N_94,In_400,In_379);
or U95 (N_95,In_416,In_163);
nor U96 (N_96,In_118,N_15);
and U97 (N_97,In_414,In_316);
nand U98 (N_98,N_34,N_17);
nand U99 (N_99,In_179,In_380);
or U100 (N_100,N_22,In_20);
nand U101 (N_101,In_258,In_63);
or U102 (N_102,In_244,In_483);
nor U103 (N_103,In_47,In_335);
nand U104 (N_104,N_21,N_43);
nor U105 (N_105,In_36,N_45);
or U106 (N_106,In_278,In_22);
or U107 (N_107,In_115,In_286);
and U108 (N_108,N_18,In_126);
nor U109 (N_109,N_48,In_466);
or U110 (N_110,N_27,In_338);
nor U111 (N_111,In_320,In_419);
nand U112 (N_112,In_493,In_457);
nor U113 (N_113,In_300,In_210);
and U114 (N_114,In_269,In_27);
nor U115 (N_115,In_267,In_306);
nor U116 (N_116,In_112,In_246);
nor U117 (N_117,In_104,In_145);
nand U118 (N_118,In_98,In_54);
and U119 (N_119,In_354,In_140);
or U120 (N_120,N_3,In_322);
and U121 (N_121,N_64,In_398);
nor U122 (N_122,N_107,In_209);
and U123 (N_123,In_158,In_99);
nand U124 (N_124,N_49,In_195);
nor U125 (N_125,In_347,N_56);
and U126 (N_126,In_303,In_90);
and U127 (N_127,N_67,In_408);
and U128 (N_128,N_14,In_336);
nor U129 (N_129,In_79,N_80);
nand U130 (N_130,In_198,N_119);
or U131 (N_131,In_395,In_332);
and U132 (N_132,N_93,In_101);
nand U133 (N_133,In_418,In_185);
nor U134 (N_134,In_143,In_362);
and U135 (N_135,In_378,N_59);
nor U136 (N_136,In_417,In_432);
nor U137 (N_137,N_70,N_105);
and U138 (N_138,N_87,In_472);
and U139 (N_139,In_464,In_328);
or U140 (N_140,In_65,N_76);
nand U141 (N_141,In_394,In_223);
or U142 (N_142,In_489,In_87);
nand U143 (N_143,In_100,N_36);
nor U144 (N_144,In_161,In_311);
or U145 (N_145,N_42,In_69);
nor U146 (N_146,In_287,In_85);
nand U147 (N_147,In_264,In_220);
and U148 (N_148,N_61,In_214);
nand U149 (N_149,In_229,In_420);
and U150 (N_150,In_312,In_39);
or U151 (N_151,In_19,In_197);
nor U152 (N_152,N_94,In_433);
nand U153 (N_153,N_95,In_359);
and U154 (N_154,In_360,In_412);
nor U155 (N_155,N_99,In_200);
and U156 (N_156,N_39,In_225);
and U157 (N_157,In_387,In_95);
nor U158 (N_158,In_314,In_139);
or U159 (N_159,N_118,N_65);
and U160 (N_160,N_109,In_349);
or U161 (N_161,N_2,In_441);
nor U162 (N_162,In_242,In_238);
xor U163 (N_163,In_453,In_333);
and U164 (N_164,In_451,In_111);
nand U165 (N_165,N_72,In_61);
nor U166 (N_166,N_101,N_113);
and U167 (N_167,In_249,N_54);
or U168 (N_168,In_495,N_106);
or U169 (N_169,N_58,N_1);
and U170 (N_170,In_117,In_208);
and U171 (N_171,In_435,In_370);
or U172 (N_172,In_382,In_204);
and U173 (N_173,In_404,In_181);
and U174 (N_174,In_399,In_296);
and U175 (N_175,In_351,N_41);
nor U176 (N_176,In_427,In_342);
nand U177 (N_177,N_46,In_135);
nor U178 (N_178,In_217,N_82);
nand U179 (N_179,In_371,In_64);
nor U180 (N_180,N_133,N_7);
or U181 (N_181,N_83,N_37);
and U182 (N_182,N_69,N_172);
or U183 (N_183,N_171,N_81);
nand U184 (N_184,In_74,In_429);
nand U185 (N_185,N_104,N_111);
nand U186 (N_186,N_60,In_153);
or U187 (N_187,In_397,N_130);
or U188 (N_188,N_73,In_105);
nor U189 (N_189,In_232,N_124);
nand U190 (N_190,N_47,In_250);
nand U191 (N_191,In_449,In_157);
nor U192 (N_192,In_187,N_12);
or U193 (N_193,In_77,In_134);
nand U194 (N_194,In_452,In_1);
nand U195 (N_195,In_203,N_167);
and U196 (N_196,N_121,In_170);
and U197 (N_197,In_302,N_166);
or U198 (N_198,N_163,N_127);
nand U199 (N_199,N_175,N_128);
and U200 (N_200,N_148,In_17);
or U201 (N_201,In_281,N_98);
or U202 (N_202,In_131,In_147);
or U203 (N_203,N_144,N_178);
nor U204 (N_204,In_247,N_66);
nand U205 (N_205,N_102,In_463);
or U206 (N_206,In_450,N_160);
nor U207 (N_207,N_164,In_459);
nor U208 (N_208,In_183,N_40);
or U209 (N_209,N_84,N_92);
nand U210 (N_210,N_16,In_446);
nor U211 (N_211,N_86,In_337);
nand U212 (N_212,In_491,N_52);
nand U213 (N_213,N_74,In_33);
and U214 (N_214,In_490,N_31);
nand U215 (N_215,In_51,N_151);
nand U216 (N_216,N_162,In_146);
nand U217 (N_217,In_469,In_480);
or U218 (N_218,In_357,In_346);
nand U219 (N_219,In_377,N_136);
nor U220 (N_220,In_439,In_48);
nand U221 (N_221,In_253,In_78);
nor U222 (N_222,In_11,N_140);
nor U223 (N_223,In_326,In_436);
or U224 (N_224,In_16,In_218);
nand U225 (N_225,In_138,N_115);
or U226 (N_226,In_325,N_131);
and U227 (N_227,In_334,In_132);
or U228 (N_228,In_94,In_353);
and U229 (N_229,In_13,In_166);
nand U230 (N_230,In_389,In_368);
nand U231 (N_231,In_356,In_172);
nand U232 (N_232,N_176,In_103);
nand U233 (N_233,In_411,In_114);
nand U234 (N_234,In_222,In_9);
and U235 (N_235,In_122,N_30);
and U236 (N_236,N_145,In_260);
nor U237 (N_237,In_434,N_71);
nor U238 (N_238,N_141,N_125);
and U239 (N_239,N_152,In_470);
or U240 (N_240,N_238,N_150);
or U241 (N_241,N_165,N_139);
nand U242 (N_242,In_293,N_221);
and U243 (N_243,N_183,N_185);
and U244 (N_244,In_127,N_181);
and U245 (N_245,In_423,N_38);
or U246 (N_246,N_224,N_169);
nand U247 (N_247,N_218,N_63);
nand U248 (N_248,N_220,In_386);
or U249 (N_249,N_33,In_80);
and U250 (N_250,N_198,N_225);
and U251 (N_251,N_62,N_147);
or U252 (N_252,N_138,In_496);
nor U253 (N_253,N_123,N_210);
or U254 (N_254,N_53,N_195);
or U255 (N_255,N_126,In_409);
nor U256 (N_256,In_254,In_188);
and U257 (N_257,In_374,N_88);
nor U258 (N_258,N_186,In_18);
and U259 (N_259,In_424,In_304);
or U260 (N_260,N_193,In_211);
or U261 (N_261,In_494,In_124);
nor U262 (N_262,In_82,N_222);
or U263 (N_263,N_154,In_31);
and U264 (N_264,N_213,In_68);
nor U265 (N_265,In_271,In_160);
and U266 (N_266,In_2,N_188);
nand U267 (N_267,N_4,N_29);
nor U268 (N_268,In_52,In_81);
nand U269 (N_269,In_26,N_78);
nand U270 (N_270,In_285,N_13);
or U271 (N_271,In_191,In_236);
nor U272 (N_272,In_180,N_0);
and U273 (N_273,In_120,In_125);
nor U274 (N_274,N_142,N_208);
nand U275 (N_275,In_465,In_275);
nand U276 (N_276,N_44,N_199);
or U277 (N_277,N_201,N_96);
nor U278 (N_278,N_206,In_426);
or U279 (N_279,In_458,In_171);
nor U280 (N_280,N_143,N_235);
nor U281 (N_281,In_252,N_5);
or U282 (N_282,N_233,N_112);
nor U283 (N_283,N_227,In_5);
and U284 (N_284,In_498,In_410);
nor U285 (N_285,In_437,In_381);
xnor U286 (N_286,In_32,In_315);
and U287 (N_287,In_475,N_189);
nand U288 (N_288,In_277,In_276);
and U289 (N_289,In_110,N_28);
nand U290 (N_290,N_192,In_50);
nor U291 (N_291,N_226,In_221);
or U292 (N_292,N_180,In_310);
nand U293 (N_293,N_24,N_137);
or U294 (N_294,N_223,N_232);
nor U295 (N_295,In_201,In_339);
or U296 (N_296,In_460,In_444);
and U297 (N_297,In_0,In_55);
nand U298 (N_298,N_209,N_122);
nor U299 (N_299,N_239,In_133);
or U300 (N_300,In_243,N_204);
nand U301 (N_301,N_157,N_217);
nor U302 (N_302,N_77,N_229);
nor U303 (N_303,N_91,In_289);
nor U304 (N_304,N_191,N_270);
nand U305 (N_305,N_292,In_141);
nor U306 (N_306,In_93,In_24);
nor U307 (N_307,N_117,In_231);
and U308 (N_308,N_294,In_319);
nand U309 (N_309,N_241,In_116);
or U310 (N_310,N_255,In_142);
nor U311 (N_311,In_123,In_456);
nor U312 (N_312,N_264,In_462);
and U313 (N_313,N_212,N_153);
nand U314 (N_314,N_25,N_214);
or U315 (N_315,N_149,N_35);
nand U316 (N_316,N_168,N_120);
or U317 (N_317,N_159,N_251);
xnor U318 (N_318,N_100,In_324);
or U319 (N_319,In_228,N_293);
and U320 (N_320,N_252,In_331);
nand U321 (N_321,N_196,N_85);
and U322 (N_322,In_159,N_190);
or U323 (N_323,In_471,N_161);
nand U324 (N_324,In_415,N_55);
and U325 (N_325,In_148,N_135);
or U326 (N_326,N_116,N_194);
or U327 (N_327,In_202,In_393);
nand U328 (N_328,N_103,In_272);
nor U329 (N_329,In_239,In_376);
or U330 (N_330,N_242,N_281);
and U331 (N_331,N_97,N_240);
nor U332 (N_332,In_294,N_187);
nor U333 (N_333,N_272,N_257);
nand U334 (N_334,N_266,N_243);
nor U335 (N_335,N_202,N_231);
or U336 (N_336,N_253,N_275);
and U337 (N_337,N_200,In_474);
nor U338 (N_338,In_403,In_266);
nor U339 (N_339,N_170,N_268);
nand U340 (N_340,In_421,In_461);
nand U341 (N_341,N_263,In_10);
or U342 (N_342,In_53,In_83);
and U343 (N_343,N_265,N_205);
and U344 (N_344,In_189,In_42);
nand U345 (N_345,In_119,N_211);
nand U346 (N_346,N_289,N_158);
nor U347 (N_347,N_173,N_273);
nor U348 (N_348,N_236,N_108);
or U349 (N_349,In_341,N_132);
or U350 (N_350,N_75,N_267);
and U351 (N_351,N_234,N_244);
nand U352 (N_352,N_50,In_37);
nor U353 (N_353,N_249,In_4);
xnor U354 (N_354,N_79,In_321);
or U355 (N_355,In_234,N_8);
nor U356 (N_356,N_295,N_284);
nand U357 (N_357,In_327,In_43);
nand U358 (N_358,In_391,In_262);
nor U359 (N_359,In_28,N_11);
nand U360 (N_360,In_45,In_265);
or U361 (N_361,In_413,N_297);
and U362 (N_362,N_278,N_207);
or U363 (N_363,In_405,In_184);
nor U364 (N_364,N_356,In_84);
nor U365 (N_365,N_110,N_254);
nand U366 (N_366,N_352,N_260);
and U367 (N_367,N_337,N_330);
or U368 (N_368,N_89,N_179);
nand U369 (N_369,N_325,N_338);
or U370 (N_370,N_182,N_301);
nor U371 (N_371,N_298,N_343);
or U372 (N_372,N_219,N_304);
or U373 (N_373,N_246,N_339);
nand U374 (N_374,N_315,N_318);
or U375 (N_375,N_287,N_331);
nand U376 (N_376,N_358,In_152);
or U377 (N_377,N_250,N_353);
and U378 (N_378,N_259,N_286);
nor U379 (N_379,N_346,N_335);
or U380 (N_380,N_319,N_134);
or U381 (N_381,In_92,N_334);
and U382 (N_382,N_271,In_468);
and U383 (N_383,N_332,N_261);
and U384 (N_384,N_317,N_296);
and U385 (N_385,N_312,N_344);
nand U386 (N_386,N_329,N_129);
or U387 (N_387,N_307,N_341);
or U388 (N_388,In_66,In_59);
nand U389 (N_389,N_228,N_350);
nor U390 (N_390,In_56,N_326);
nand U391 (N_391,N_354,N_245);
nor U392 (N_392,N_327,N_345);
or U393 (N_393,N_26,N_237);
and U394 (N_394,N_174,N_156);
and U395 (N_395,N_283,N_290);
and U396 (N_396,N_316,N_333);
xnor U397 (N_397,N_114,N_305);
nand U398 (N_398,In_175,N_262);
nor U399 (N_399,N_277,N_303);
or U400 (N_400,N_340,In_199);
or U401 (N_401,N_216,In_96);
nand U402 (N_402,N_215,N_314);
or U403 (N_403,N_258,N_248);
nor U404 (N_404,N_280,N_269);
or U405 (N_405,N_320,In_167);
nor U406 (N_406,N_336,N_282);
nor U407 (N_407,N_276,N_90);
and U408 (N_408,In_251,N_355);
nor U409 (N_409,In_137,N_177);
and U410 (N_410,N_328,N_300);
or U411 (N_411,N_203,In_177);
nand U412 (N_412,In_186,N_324);
or U413 (N_413,N_347,N_351);
and U414 (N_414,N_321,N_230);
and U415 (N_415,N_349,N_279);
nor U416 (N_416,In_406,N_322);
nor U417 (N_417,N_308,In_282);
and U418 (N_418,In_182,N_309);
nand U419 (N_419,N_291,N_146);
nand U420 (N_420,N_395,N_361);
or U421 (N_421,N_247,N_378);
nand U422 (N_422,N_392,N_381);
or U423 (N_423,N_419,N_363);
nand U424 (N_424,N_348,N_416);
nand U425 (N_425,N_417,N_374);
and U426 (N_426,N_385,N_302);
or U427 (N_427,N_373,N_376);
or U428 (N_428,N_394,N_367);
nor U429 (N_429,N_403,N_405);
or U430 (N_430,N_408,N_411);
nor U431 (N_431,N_274,N_323);
nor U432 (N_432,N_389,N_371);
xor U433 (N_433,N_256,N_397);
and U434 (N_434,N_418,N_401);
or U435 (N_435,N_413,N_409);
nor U436 (N_436,N_366,N_313);
xnor U437 (N_437,N_368,N_406);
nand U438 (N_438,N_375,N_391);
and U439 (N_439,N_410,N_342);
and U440 (N_440,N_384,N_357);
nor U441 (N_441,N_379,N_380);
and U442 (N_442,N_415,N_365);
and U443 (N_443,N_68,N_359);
nand U444 (N_444,N_390,N_400);
nand U445 (N_445,N_396,N_382);
and U446 (N_446,N_388,N_299);
nand U447 (N_447,N_414,N_362);
and U448 (N_448,N_398,N_155);
or U449 (N_449,N_387,N_393);
nand U450 (N_450,N_369,N_370);
and U451 (N_451,N_306,N_399);
nand U452 (N_452,N_402,N_383);
nand U453 (N_453,N_386,N_372);
and U454 (N_454,N_360,N_407);
and U455 (N_455,N_412,N_364);
nand U456 (N_456,N_288,N_285);
nand U457 (N_457,N_404,N_310);
and U458 (N_458,N_377,N_311);
nor U459 (N_459,N_197,N_184);
nand U460 (N_460,N_418,N_311);
nand U461 (N_461,N_412,N_368);
nand U462 (N_462,N_376,N_348);
or U463 (N_463,N_377,N_360);
nor U464 (N_464,N_371,N_396);
nand U465 (N_465,N_403,N_302);
nand U466 (N_466,N_386,N_416);
or U467 (N_467,N_342,N_383);
nand U468 (N_468,N_394,N_380);
or U469 (N_469,N_299,N_391);
and U470 (N_470,N_405,N_376);
or U471 (N_471,N_392,N_68);
and U472 (N_472,N_376,N_310);
and U473 (N_473,N_384,N_413);
and U474 (N_474,N_419,N_360);
or U475 (N_475,N_394,N_408);
nor U476 (N_476,N_364,N_313);
nand U477 (N_477,N_323,N_371);
xor U478 (N_478,N_387,N_408);
xor U479 (N_479,N_288,N_370);
and U480 (N_480,N_443,N_460);
nand U481 (N_481,N_433,N_461);
nand U482 (N_482,N_477,N_442);
and U483 (N_483,N_421,N_470);
or U484 (N_484,N_438,N_434);
or U485 (N_485,N_431,N_445);
or U486 (N_486,N_444,N_472);
or U487 (N_487,N_458,N_475);
nor U488 (N_488,N_429,N_450);
nor U489 (N_489,N_466,N_435);
or U490 (N_490,N_422,N_441);
and U491 (N_491,N_423,N_427);
xor U492 (N_492,N_463,N_439);
nor U493 (N_493,N_424,N_430);
nand U494 (N_494,N_454,N_457);
and U495 (N_495,N_428,N_459);
and U496 (N_496,N_432,N_467);
nand U497 (N_497,N_420,N_436);
nor U498 (N_498,N_468,N_437);
or U499 (N_499,N_476,N_469);
nand U500 (N_500,N_455,N_474);
nor U501 (N_501,N_452,N_440);
and U502 (N_502,N_462,N_446);
nor U503 (N_503,N_464,N_449);
nor U504 (N_504,N_456,N_479);
and U505 (N_505,N_478,N_451);
or U506 (N_506,N_425,N_453);
nand U507 (N_507,N_471,N_448);
and U508 (N_508,N_473,N_465);
nand U509 (N_509,N_426,N_447);
and U510 (N_510,N_431,N_472);
or U511 (N_511,N_441,N_464);
or U512 (N_512,N_423,N_477);
nand U513 (N_513,N_449,N_451);
nand U514 (N_514,N_434,N_468);
nand U515 (N_515,N_477,N_447);
nor U516 (N_516,N_424,N_479);
nand U517 (N_517,N_430,N_426);
and U518 (N_518,N_420,N_433);
nand U519 (N_519,N_450,N_431);
nand U520 (N_520,N_422,N_457);
nand U521 (N_521,N_469,N_474);
nor U522 (N_522,N_448,N_444);
nor U523 (N_523,N_436,N_475);
or U524 (N_524,N_469,N_453);
nand U525 (N_525,N_432,N_478);
nor U526 (N_526,N_476,N_426);
or U527 (N_527,N_446,N_450);
nand U528 (N_528,N_435,N_432);
nor U529 (N_529,N_466,N_424);
nand U530 (N_530,N_434,N_467);
or U531 (N_531,N_421,N_448);
and U532 (N_532,N_441,N_426);
or U533 (N_533,N_443,N_453);
and U534 (N_534,N_444,N_453);
nand U535 (N_535,N_474,N_465);
and U536 (N_536,N_454,N_432);
and U537 (N_537,N_421,N_441);
nor U538 (N_538,N_451,N_425);
nor U539 (N_539,N_439,N_450);
nand U540 (N_540,N_510,N_491);
nand U541 (N_541,N_493,N_529);
nor U542 (N_542,N_521,N_503);
or U543 (N_543,N_492,N_527);
or U544 (N_544,N_496,N_505);
or U545 (N_545,N_502,N_499);
nor U546 (N_546,N_504,N_517);
nor U547 (N_547,N_531,N_532);
and U548 (N_548,N_538,N_513);
nand U549 (N_549,N_518,N_520);
or U550 (N_550,N_501,N_526);
or U551 (N_551,N_486,N_489);
and U552 (N_552,N_481,N_482);
and U553 (N_553,N_483,N_516);
nor U554 (N_554,N_507,N_537);
nand U555 (N_555,N_497,N_511);
or U556 (N_556,N_515,N_512);
nand U557 (N_557,N_500,N_530);
and U558 (N_558,N_533,N_519);
nor U559 (N_559,N_514,N_535);
or U560 (N_560,N_523,N_498);
nand U561 (N_561,N_524,N_539);
nand U562 (N_562,N_508,N_485);
and U563 (N_563,N_522,N_487);
nand U564 (N_564,N_490,N_495);
nand U565 (N_565,N_484,N_528);
and U566 (N_566,N_480,N_488);
nor U567 (N_567,N_525,N_509);
nand U568 (N_568,N_494,N_506);
nand U569 (N_569,N_536,N_534);
nor U570 (N_570,N_487,N_516);
nor U571 (N_571,N_495,N_523);
nor U572 (N_572,N_484,N_525);
nand U573 (N_573,N_502,N_486);
and U574 (N_574,N_480,N_514);
or U575 (N_575,N_507,N_506);
nor U576 (N_576,N_536,N_492);
nor U577 (N_577,N_525,N_480);
nand U578 (N_578,N_494,N_535);
and U579 (N_579,N_507,N_487);
and U580 (N_580,N_530,N_508);
or U581 (N_581,N_539,N_538);
or U582 (N_582,N_500,N_502);
nor U583 (N_583,N_492,N_482);
nor U584 (N_584,N_504,N_491);
nand U585 (N_585,N_502,N_509);
and U586 (N_586,N_506,N_486);
nand U587 (N_587,N_522,N_481);
and U588 (N_588,N_485,N_491);
nand U589 (N_589,N_526,N_537);
or U590 (N_590,N_492,N_487);
nor U591 (N_591,N_535,N_512);
nand U592 (N_592,N_526,N_509);
xor U593 (N_593,N_516,N_492);
nand U594 (N_594,N_508,N_510);
nor U595 (N_595,N_489,N_488);
or U596 (N_596,N_486,N_513);
and U597 (N_597,N_497,N_499);
nand U598 (N_598,N_495,N_502);
nand U599 (N_599,N_504,N_527);
or U600 (N_600,N_552,N_578);
nor U601 (N_601,N_561,N_574);
nand U602 (N_602,N_582,N_579);
and U603 (N_603,N_587,N_599);
nand U604 (N_604,N_545,N_557);
nor U605 (N_605,N_543,N_580);
nand U606 (N_606,N_584,N_559);
and U607 (N_607,N_546,N_565);
or U608 (N_608,N_590,N_575);
nand U609 (N_609,N_598,N_594);
or U610 (N_610,N_577,N_572);
nor U611 (N_611,N_585,N_547);
nand U612 (N_612,N_550,N_562);
and U613 (N_613,N_560,N_570);
and U614 (N_614,N_576,N_583);
nand U615 (N_615,N_568,N_573);
nand U616 (N_616,N_566,N_592);
nand U617 (N_617,N_548,N_549);
or U618 (N_618,N_541,N_544);
or U619 (N_619,N_591,N_555);
nand U620 (N_620,N_556,N_554);
or U621 (N_621,N_596,N_558);
or U622 (N_622,N_586,N_542);
nand U623 (N_623,N_564,N_563);
or U624 (N_624,N_551,N_569);
or U625 (N_625,N_553,N_595);
nor U626 (N_626,N_593,N_567);
xor U627 (N_627,N_581,N_589);
or U628 (N_628,N_540,N_588);
and U629 (N_629,N_571,N_597);
nor U630 (N_630,N_573,N_551);
nand U631 (N_631,N_545,N_555);
nand U632 (N_632,N_541,N_551);
and U633 (N_633,N_591,N_599);
or U634 (N_634,N_548,N_588);
and U635 (N_635,N_598,N_558);
nor U636 (N_636,N_568,N_591);
nor U637 (N_637,N_596,N_547);
nor U638 (N_638,N_559,N_548);
nor U639 (N_639,N_560,N_544);
nor U640 (N_640,N_555,N_575);
or U641 (N_641,N_563,N_572);
nor U642 (N_642,N_555,N_571);
nor U643 (N_643,N_578,N_596);
nand U644 (N_644,N_560,N_598);
nand U645 (N_645,N_540,N_549);
nor U646 (N_646,N_565,N_559);
nand U647 (N_647,N_542,N_553);
nand U648 (N_648,N_555,N_552);
nor U649 (N_649,N_585,N_557);
nand U650 (N_650,N_551,N_597);
nand U651 (N_651,N_575,N_540);
and U652 (N_652,N_578,N_579);
or U653 (N_653,N_555,N_567);
nand U654 (N_654,N_594,N_560);
nand U655 (N_655,N_594,N_554);
nand U656 (N_656,N_591,N_540);
nor U657 (N_657,N_592,N_578);
nand U658 (N_658,N_560,N_563);
nor U659 (N_659,N_576,N_542);
and U660 (N_660,N_641,N_644);
nor U661 (N_661,N_647,N_637);
or U662 (N_662,N_654,N_652);
nor U663 (N_663,N_614,N_643);
nor U664 (N_664,N_646,N_656);
nand U665 (N_665,N_618,N_611);
and U666 (N_666,N_617,N_602);
and U667 (N_667,N_604,N_621);
nor U668 (N_668,N_651,N_648);
nand U669 (N_669,N_619,N_607);
nand U670 (N_670,N_638,N_632);
and U671 (N_671,N_650,N_645);
nor U672 (N_672,N_636,N_624);
or U673 (N_673,N_626,N_612);
nor U674 (N_674,N_629,N_601);
nand U675 (N_675,N_630,N_610);
and U676 (N_676,N_631,N_605);
or U677 (N_677,N_657,N_603);
xnor U678 (N_678,N_655,N_625);
and U679 (N_679,N_633,N_649);
nor U680 (N_680,N_608,N_616);
nor U681 (N_681,N_609,N_606);
nand U682 (N_682,N_627,N_659);
nor U683 (N_683,N_639,N_634);
or U684 (N_684,N_628,N_642);
and U685 (N_685,N_615,N_613);
and U686 (N_686,N_622,N_640);
and U687 (N_687,N_658,N_653);
and U688 (N_688,N_623,N_600);
nand U689 (N_689,N_635,N_620);
nand U690 (N_690,N_619,N_612);
and U691 (N_691,N_640,N_600);
and U692 (N_692,N_656,N_618);
or U693 (N_693,N_649,N_627);
and U694 (N_694,N_642,N_625);
and U695 (N_695,N_638,N_639);
or U696 (N_696,N_601,N_607);
nand U697 (N_697,N_603,N_600);
and U698 (N_698,N_620,N_641);
or U699 (N_699,N_654,N_649);
and U700 (N_700,N_651,N_629);
nand U701 (N_701,N_609,N_646);
or U702 (N_702,N_602,N_648);
nor U703 (N_703,N_635,N_622);
and U704 (N_704,N_602,N_608);
nor U705 (N_705,N_631,N_627);
nand U706 (N_706,N_612,N_610);
and U707 (N_707,N_647,N_609);
nor U708 (N_708,N_615,N_610);
or U709 (N_709,N_642,N_633);
or U710 (N_710,N_610,N_619);
or U711 (N_711,N_606,N_614);
nand U712 (N_712,N_644,N_610);
or U713 (N_713,N_616,N_610);
nand U714 (N_714,N_634,N_644);
nor U715 (N_715,N_636,N_625);
and U716 (N_716,N_603,N_630);
or U717 (N_717,N_639,N_621);
nand U718 (N_718,N_631,N_652);
nor U719 (N_719,N_638,N_658);
or U720 (N_720,N_667,N_702);
nor U721 (N_721,N_700,N_674);
nor U722 (N_722,N_680,N_698);
and U723 (N_723,N_707,N_701);
or U724 (N_724,N_675,N_694);
nand U725 (N_725,N_664,N_669);
nand U726 (N_726,N_677,N_705);
nand U727 (N_727,N_709,N_693);
or U728 (N_728,N_717,N_699);
nand U729 (N_729,N_665,N_704);
nand U730 (N_730,N_714,N_718);
and U731 (N_731,N_706,N_692);
nand U732 (N_732,N_689,N_712);
nor U733 (N_733,N_703,N_661);
nor U734 (N_734,N_690,N_682);
or U735 (N_735,N_684,N_670);
or U736 (N_736,N_713,N_688);
and U737 (N_737,N_719,N_673);
nor U738 (N_738,N_687,N_696);
nor U739 (N_739,N_683,N_691);
and U740 (N_740,N_668,N_708);
nand U741 (N_741,N_695,N_685);
and U742 (N_742,N_710,N_681);
and U743 (N_743,N_711,N_672);
and U744 (N_744,N_660,N_679);
nor U745 (N_745,N_678,N_666);
nor U746 (N_746,N_663,N_686);
nor U747 (N_747,N_676,N_697);
and U748 (N_748,N_716,N_662);
nor U749 (N_749,N_671,N_715);
nand U750 (N_750,N_710,N_695);
or U751 (N_751,N_682,N_684);
nand U752 (N_752,N_701,N_717);
nor U753 (N_753,N_719,N_662);
or U754 (N_754,N_678,N_697);
nand U755 (N_755,N_708,N_716);
nand U756 (N_756,N_695,N_660);
and U757 (N_757,N_684,N_715);
and U758 (N_758,N_672,N_686);
or U759 (N_759,N_678,N_690);
and U760 (N_760,N_693,N_697);
nor U761 (N_761,N_691,N_665);
nand U762 (N_762,N_698,N_706);
or U763 (N_763,N_718,N_688);
and U764 (N_764,N_662,N_709);
or U765 (N_765,N_712,N_680);
or U766 (N_766,N_665,N_687);
or U767 (N_767,N_678,N_714);
and U768 (N_768,N_679,N_718);
and U769 (N_769,N_713,N_665);
nand U770 (N_770,N_715,N_709);
nor U771 (N_771,N_676,N_709);
nand U772 (N_772,N_674,N_693);
and U773 (N_773,N_687,N_714);
nand U774 (N_774,N_709,N_698);
nor U775 (N_775,N_673,N_712);
and U776 (N_776,N_719,N_705);
and U777 (N_777,N_689,N_663);
nand U778 (N_778,N_673,N_682);
nor U779 (N_779,N_713,N_698);
nor U780 (N_780,N_775,N_778);
and U781 (N_781,N_735,N_771);
nand U782 (N_782,N_755,N_752);
or U783 (N_783,N_759,N_731);
and U784 (N_784,N_776,N_764);
or U785 (N_785,N_734,N_725);
nand U786 (N_786,N_777,N_772);
or U787 (N_787,N_732,N_741);
or U788 (N_788,N_761,N_763);
nor U789 (N_789,N_742,N_758);
and U790 (N_790,N_743,N_748);
nor U791 (N_791,N_723,N_756);
nor U792 (N_792,N_720,N_738);
nor U793 (N_793,N_728,N_751);
and U794 (N_794,N_750,N_767);
or U795 (N_795,N_745,N_724);
nor U796 (N_796,N_774,N_722);
and U797 (N_797,N_729,N_766);
and U798 (N_798,N_733,N_773);
nand U799 (N_799,N_760,N_765);
and U800 (N_800,N_740,N_737);
and U801 (N_801,N_736,N_726);
nand U802 (N_802,N_749,N_730);
nand U803 (N_803,N_768,N_744);
nand U804 (N_804,N_746,N_753);
and U805 (N_805,N_770,N_754);
nor U806 (N_806,N_762,N_779);
and U807 (N_807,N_721,N_747);
or U808 (N_808,N_769,N_757);
or U809 (N_809,N_727,N_739);
nand U810 (N_810,N_730,N_740);
nor U811 (N_811,N_764,N_778);
and U812 (N_812,N_721,N_772);
nand U813 (N_813,N_770,N_772);
nor U814 (N_814,N_725,N_739);
nor U815 (N_815,N_758,N_768);
nand U816 (N_816,N_732,N_745);
and U817 (N_817,N_748,N_732);
and U818 (N_818,N_758,N_770);
nor U819 (N_819,N_724,N_732);
or U820 (N_820,N_752,N_774);
nor U821 (N_821,N_724,N_737);
or U822 (N_822,N_768,N_749);
or U823 (N_823,N_763,N_732);
nand U824 (N_824,N_732,N_744);
nand U825 (N_825,N_749,N_763);
nand U826 (N_826,N_727,N_776);
or U827 (N_827,N_774,N_735);
nand U828 (N_828,N_760,N_756);
and U829 (N_829,N_769,N_770);
nand U830 (N_830,N_733,N_750);
or U831 (N_831,N_737,N_779);
nand U832 (N_832,N_761,N_733);
nand U833 (N_833,N_736,N_779);
nor U834 (N_834,N_775,N_751);
or U835 (N_835,N_767,N_738);
nor U836 (N_836,N_763,N_769);
or U837 (N_837,N_766,N_731);
and U838 (N_838,N_742,N_748);
and U839 (N_839,N_721,N_748);
nand U840 (N_840,N_816,N_803);
nor U841 (N_841,N_823,N_818);
nand U842 (N_842,N_808,N_833);
and U843 (N_843,N_809,N_835);
nand U844 (N_844,N_800,N_798);
nor U845 (N_845,N_789,N_782);
nor U846 (N_846,N_792,N_806);
and U847 (N_847,N_826,N_804);
nand U848 (N_848,N_797,N_828);
nand U849 (N_849,N_802,N_785);
nor U850 (N_850,N_813,N_831);
nand U851 (N_851,N_834,N_791);
or U852 (N_852,N_783,N_786);
or U853 (N_853,N_815,N_824);
nand U854 (N_854,N_781,N_829);
nand U855 (N_855,N_812,N_790);
nand U856 (N_856,N_788,N_832);
or U857 (N_857,N_787,N_794);
and U858 (N_858,N_795,N_793);
nand U859 (N_859,N_839,N_822);
nor U860 (N_860,N_821,N_827);
nand U861 (N_861,N_801,N_780);
nand U862 (N_862,N_814,N_820);
nor U863 (N_863,N_837,N_807);
or U864 (N_864,N_796,N_838);
nor U865 (N_865,N_817,N_799);
nor U866 (N_866,N_830,N_805);
xnor U867 (N_867,N_825,N_819);
nand U868 (N_868,N_784,N_811);
nand U869 (N_869,N_836,N_810);
and U870 (N_870,N_780,N_835);
xnor U871 (N_871,N_802,N_787);
or U872 (N_872,N_793,N_831);
nand U873 (N_873,N_815,N_801);
or U874 (N_874,N_820,N_808);
nand U875 (N_875,N_782,N_791);
nor U876 (N_876,N_825,N_838);
nand U877 (N_877,N_792,N_802);
nor U878 (N_878,N_794,N_839);
nor U879 (N_879,N_838,N_809);
and U880 (N_880,N_809,N_819);
and U881 (N_881,N_809,N_805);
or U882 (N_882,N_830,N_838);
or U883 (N_883,N_799,N_786);
nor U884 (N_884,N_806,N_788);
nor U885 (N_885,N_786,N_789);
or U886 (N_886,N_813,N_796);
or U887 (N_887,N_819,N_827);
and U888 (N_888,N_832,N_793);
and U889 (N_889,N_839,N_820);
or U890 (N_890,N_784,N_830);
nor U891 (N_891,N_781,N_797);
nor U892 (N_892,N_810,N_784);
nand U893 (N_893,N_799,N_807);
nor U894 (N_894,N_781,N_801);
nor U895 (N_895,N_801,N_825);
or U896 (N_896,N_818,N_830);
nand U897 (N_897,N_822,N_823);
or U898 (N_898,N_810,N_782);
or U899 (N_899,N_792,N_787);
or U900 (N_900,N_846,N_893);
and U901 (N_901,N_859,N_897);
nor U902 (N_902,N_862,N_843);
nor U903 (N_903,N_891,N_892);
or U904 (N_904,N_879,N_850);
nor U905 (N_905,N_852,N_863);
and U906 (N_906,N_844,N_881);
nand U907 (N_907,N_883,N_871);
nor U908 (N_908,N_853,N_894);
nor U909 (N_909,N_842,N_847);
or U910 (N_910,N_870,N_882);
and U911 (N_911,N_861,N_899);
nor U912 (N_912,N_840,N_865);
or U913 (N_913,N_886,N_854);
and U914 (N_914,N_898,N_855);
and U915 (N_915,N_841,N_849);
or U916 (N_916,N_880,N_872);
or U917 (N_917,N_876,N_889);
and U918 (N_918,N_857,N_885);
or U919 (N_919,N_848,N_874);
and U920 (N_920,N_888,N_851);
or U921 (N_921,N_890,N_896);
nand U922 (N_922,N_869,N_877);
nor U923 (N_923,N_887,N_868);
nand U924 (N_924,N_875,N_895);
nand U925 (N_925,N_845,N_867);
nor U926 (N_926,N_866,N_858);
nand U927 (N_927,N_878,N_856);
nor U928 (N_928,N_864,N_860);
nand U929 (N_929,N_884,N_873);
nor U930 (N_930,N_873,N_891);
or U931 (N_931,N_883,N_895);
and U932 (N_932,N_894,N_860);
and U933 (N_933,N_894,N_899);
or U934 (N_934,N_887,N_848);
nand U935 (N_935,N_851,N_857);
and U936 (N_936,N_859,N_889);
nand U937 (N_937,N_865,N_887);
nor U938 (N_938,N_896,N_891);
or U939 (N_939,N_841,N_851);
or U940 (N_940,N_894,N_861);
xor U941 (N_941,N_864,N_899);
nor U942 (N_942,N_870,N_875);
nor U943 (N_943,N_894,N_845);
and U944 (N_944,N_860,N_892);
nor U945 (N_945,N_861,N_892);
and U946 (N_946,N_887,N_866);
and U947 (N_947,N_858,N_857);
or U948 (N_948,N_850,N_854);
nor U949 (N_949,N_869,N_845);
nand U950 (N_950,N_864,N_858);
or U951 (N_951,N_870,N_895);
and U952 (N_952,N_854,N_851);
or U953 (N_953,N_878,N_888);
nor U954 (N_954,N_845,N_873);
nor U955 (N_955,N_842,N_875);
or U956 (N_956,N_875,N_846);
nor U957 (N_957,N_849,N_876);
nor U958 (N_958,N_893,N_874);
and U959 (N_959,N_866,N_876);
nand U960 (N_960,N_943,N_907);
nor U961 (N_961,N_904,N_917);
and U962 (N_962,N_909,N_941);
nor U963 (N_963,N_958,N_913);
and U964 (N_964,N_927,N_944);
nand U965 (N_965,N_923,N_929);
and U966 (N_966,N_918,N_933);
and U967 (N_967,N_906,N_934);
nor U968 (N_968,N_951,N_928);
or U969 (N_969,N_945,N_919);
and U970 (N_970,N_949,N_946);
nand U971 (N_971,N_957,N_922);
nand U972 (N_972,N_955,N_926);
nand U973 (N_973,N_925,N_905);
and U974 (N_974,N_954,N_920);
or U975 (N_975,N_910,N_947);
nand U976 (N_976,N_939,N_953);
and U977 (N_977,N_938,N_937);
nand U978 (N_978,N_931,N_935);
or U979 (N_979,N_948,N_959);
nor U980 (N_980,N_956,N_908);
or U981 (N_981,N_942,N_936);
nor U982 (N_982,N_932,N_914);
nor U983 (N_983,N_901,N_952);
and U984 (N_984,N_912,N_924);
or U985 (N_985,N_915,N_940);
nand U986 (N_986,N_903,N_916);
nand U987 (N_987,N_930,N_902);
or U988 (N_988,N_921,N_911);
nand U989 (N_989,N_900,N_950);
or U990 (N_990,N_924,N_942);
or U991 (N_991,N_931,N_929);
or U992 (N_992,N_901,N_923);
and U993 (N_993,N_912,N_906);
and U994 (N_994,N_918,N_942);
nand U995 (N_995,N_906,N_929);
nand U996 (N_996,N_934,N_916);
nand U997 (N_997,N_939,N_931);
xnor U998 (N_998,N_922,N_919);
or U999 (N_999,N_954,N_943);
and U1000 (N_1000,N_946,N_915);
and U1001 (N_1001,N_922,N_910);
nand U1002 (N_1002,N_930,N_911);
or U1003 (N_1003,N_937,N_936);
and U1004 (N_1004,N_907,N_916);
and U1005 (N_1005,N_905,N_959);
nand U1006 (N_1006,N_930,N_921);
or U1007 (N_1007,N_940,N_903);
or U1008 (N_1008,N_924,N_928);
nand U1009 (N_1009,N_906,N_940);
or U1010 (N_1010,N_958,N_906);
and U1011 (N_1011,N_948,N_904);
nand U1012 (N_1012,N_931,N_938);
nand U1013 (N_1013,N_929,N_949);
or U1014 (N_1014,N_955,N_922);
nand U1015 (N_1015,N_931,N_955);
and U1016 (N_1016,N_936,N_907);
and U1017 (N_1017,N_939,N_946);
and U1018 (N_1018,N_915,N_929);
nand U1019 (N_1019,N_947,N_942);
nand U1020 (N_1020,N_971,N_975);
and U1021 (N_1021,N_1018,N_1010);
or U1022 (N_1022,N_977,N_986);
or U1023 (N_1023,N_978,N_960);
nor U1024 (N_1024,N_999,N_991);
or U1025 (N_1025,N_964,N_990);
nand U1026 (N_1026,N_994,N_961);
and U1027 (N_1027,N_976,N_965);
nand U1028 (N_1028,N_968,N_983);
or U1029 (N_1029,N_1001,N_988);
nor U1030 (N_1030,N_985,N_1003);
nor U1031 (N_1031,N_1004,N_989);
nand U1032 (N_1032,N_1005,N_1000);
nand U1033 (N_1033,N_984,N_993);
nor U1034 (N_1034,N_970,N_1013);
and U1035 (N_1035,N_1002,N_1008);
nand U1036 (N_1036,N_1017,N_996);
nand U1037 (N_1037,N_966,N_982);
or U1038 (N_1038,N_1007,N_1012);
or U1039 (N_1039,N_992,N_1016);
and U1040 (N_1040,N_1015,N_995);
and U1041 (N_1041,N_969,N_980);
nand U1042 (N_1042,N_974,N_1011);
and U1043 (N_1043,N_973,N_997);
xor U1044 (N_1044,N_998,N_1019);
nor U1045 (N_1045,N_979,N_987);
nand U1046 (N_1046,N_1006,N_972);
and U1047 (N_1047,N_962,N_963);
nand U1048 (N_1048,N_981,N_1009);
nor U1049 (N_1049,N_967,N_1014);
nor U1050 (N_1050,N_1010,N_981);
nand U1051 (N_1051,N_1007,N_964);
nand U1052 (N_1052,N_971,N_980);
or U1053 (N_1053,N_976,N_1009);
nor U1054 (N_1054,N_981,N_1001);
nor U1055 (N_1055,N_972,N_1002);
nand U1056 (N_1056,N_976,N_1013);
or U1057 (N_1057,N_1000,N_993);
and U1058 (N_1058,N_973,N_1005);
or U1059 (N_1059,N_965,N_1016);
nor U1060 (N_1060,N_1008,N_981);
nand U1061 (N_1061,N_973,N_965);
and U1062 (N_1062,N_972,N_1003);
nand U1063 (N_1063,N_970,N_983);
and U1064 (N_1064,N_969,N_1012);
nor U1065 (N_1065,N_1002,N_1004);
and U1066 (N_1066,N_992,N_971);
and U1067 (N_1067,N_974,N_993);
and U1068 (N_1068,N_1007,N_997);
nor U1069 (N_1069,N_1019,N_1003);
nand U1070 (N_1070,N_981,N_985);
nor U1071 (N_1071,N_974,N_1005);
and U1072 (N_1072,N_982,N_961);
nand U1073 (N_1073,N_972,N_960);
nor U1074 (N_1074,N_1007,N_991);
nor U1075 (N_1075,N_969,N_1002);
nor U1076 (N_1076,N_995,N_983);
and U1077 (N_1077,N_1007,N_966);
nand U1078 (N_1078,N_978,N_976);
nand U1079 (N_1079,N_976,N_996);
and U1080 (N_1080,N_1079,N_1064);
and U1081 (N_1081,N_1061,N_1026);
or U1082 (N_1082,N_1076,N_1031);
and U1083 (N_1083,N_1058,N_1027);
or U1084 (N_1084,N_1035,N_1078);
nand U1085 (N_1085,N_1074,N_1037);
or U1086 (N_1086,N_1044,N_1071);
and U1087 (N_1087,N_1056,N_1065);
nand U1088 (N_1088,N_1059,N_1039);
nor U1089 (N_1089,N_1030,N_1041);
or U1090 (N_1090,N_1062,N_1077);
nor U1091 (N_1091,N_1068,N_1022);
and U1092 (N_1092,N_1070,N_1038);
nor U1093 (N_1093,N_1052,N_1053);
or U1094 (N_1094,N_1023,N_1032);
nor U1095 (N_1095,N_1048,N_1050);
and U1096 (N_1096,N_1057,N_1029);
nand U1097 (N_1097,N_1055,N_1025);
or U1098 (N_1098,N_1063,N_1028);
nand U1099 (N_1099,N_1046,N_1042);
nand U1100 (N_1100,N_1047,N_1075);
nor U1101 (N_1101,N_1043,N_1034);
and U1102 (N_1102,N_1060,N_1036);
nor U1103 (N_1103,N_1021,N_1051);
nand U1104 (N_1104,N_1069,N_1067);
and U1105 (N_1105,N_1033,N_1024);
nor U1106 (N_1106,N_1040,N_1045);
and U1107 (N_1107,N_1072,N_1020);
nor U1108 (N_1108,N_1054,N_1049);
nand U1109 (N_1109,N_1073,N_1066);
and U1110 (N_1110,N_1036,N_1032);
nand U1111 (N_1111,N_1048,N_1028);
and U1112 (N_1112,N_1043,N_1049);
nand U1113 (N_1113,N_1077,N_1050);
or U1114 (N_1114,N_1021,N_1038);
or U1115 (N_1115,N_1029,N_1058);
nor U1116 (N_1116,N_1027,N_1020);
nor U1117 (N_1117,N_1071,N_1078);
nor U1118 (N_1118,N_1064,N_1055);
nand U1119 (N_1119,N_1037,N_1038);
or U1120 (N_1120,N_1033,N_1026);
nor U1121 (N_1121,N_1065,N_1075);
or U1122 (N_1122,N_1075,N_1022);
nand U1123 (N_1123,N_1031,N_1030);
and U1124 (N_1124,N_1076,N_1058);
nor U1125 (N_1125,N_1054,N_1067);
and U1126 (N_1126,N_1040,N_1069);
nor U1127 (N_1127,N_1070,N_1025);
nand U1128 (N_1128,N_1065,N_1028);
nand U1129 (N_1129,N_1053,N_1059);
nor U1130 (N_1130,N_1032,N_1046);
or U1131 (N_1131,N_1037,N_1028);
and U1132 (N_1132,N_1038,N_1055);
and U1133 (N_1133,N_1041,N_1022);
and U1134 (N_1134,N_1063,N_1041);
and U1135 (N_1135,N_1062,N_1044);
nor U1136 (N_1136,N_1054,N_1041);
and U1137 (N_1137,N_1040,N_1056);
or U1138 (N_1138,N_1043,N_1046);
or U1139 (N_1139,N_1021,N_1022);
or U1140 (N_1140,N_1122,N_1093);
or U1141 (N_1141,N_1133,N_1085);
nor U1142 (N_1142,N_1109,N_1134);
nand U1143 (N_1143,N_1114,N_1111);
and U1144 (N_1144,N_1103,N_1098);
and U1145 (N_1145,N_1135,N_1138);
nand U1146 (N_1146,N_1090,N_1128);
and U1147 (N_1147,N_1082,N_1091);
and U1148 (N_1148,N_1139,N_1112);
and U1149 (N_1149,N_1087,N_1081);
or U1150 (N_1150,N_1097,N_1126);
and U1151 (N_1151,N_1086,N_1106);
and U1152 (N_1152,N_1132,N_1083);
nor U1153 (N_1153,N_1096,N_1123);
or U1154 (N_1154,N_1089,N_1115);
nor U1155 (N_1155,N_1131,N_1100);
nor U1156 (N_1156,N_1119,N_1130);
nor U1157 (N_1157,N_1116,N_1127);
nand U1158 (N_1158,N_1124,N_1102);
and U1159 (N_1159,N_1108,N_1092);
nand U1160 (N_1160,N_1136,N_1117);
or U1161 (N_1161,N_1101,N_1088);
and U1162 (N_1162,N_1120,N_1110);
nor U1163 (N_1163,N_1125,N_1129);
nand U1164 (N_1164,N_1095,N_1105);
and U1165 (N_1165,N_1113,N_1099);
and U1166 (N_1166,N_1084,N_1121);
and U1167 (N_1167,N_1094,N_1137);
nand U1168 (N_1168,N_1118,N_1080);
and U1169 (N_1169,N_1107,N_1104);
nand U1170 (N_1170,N_1109,N_1136);
nand U1171 (N_1171,N_1086,N_1118);
and U1172 (N_1172,N_1104,N_1128);
or U1173 (N_1173,N_1082,N_1109);
and U1174 (N_1174,N_1105,N_1081);
and U1175 (N_1175,N_1122,N_1087);
nor U1176 (N_1176,N_1133,N_1102);
nor U1177 (N_1177,N_1103,N_1105);
or U1178 (N_1178,N_1088,N_1128);
nand U1179 (N_1179,N_1109,N_1107);
nand U1180 (N_1180,N_1111,N_1091);
nand U1181 (N_1181,N_1098,N_1112);
or U1182 (N_1182,N_1104,N_1109);
and U1183 (N_1183,N_1122,N_1114);
or U1184 (N_1184,N_1138,N_1106);
or U1185 (N_1185,N_1080,N_1124);
or U1186 (N_1186,N_1130,N_1124);
or U1187 (N_1187,N_1081,N_1119);
nand U1188 (N_1188,N_1094,N_1126);
nand U1189 (N_1189,N_1127,N_1114);
nand U1190 (N_1190,N_1094,N_1119);
nand U1191 (N_1191,N_1108,N_1090);
nor U1192 (N_1192,N_1124,N_1115);
nor U1193 (N_1193,N_1133,N_1122);
and U1194 (N_1194,N_1128,N_1126);
or U1195 (N_1195,N_1120,N_1112);
nand U1196 (N_1196,N_1127,N_1094);
nand U1197 (N_1197,N_1114,N_1121);
nand U1198 (N_1198,N_1130,N_1109);
nor U1199 (N_1199,N_1129,N_1123);
nand U1200 (N_1200,N_1168,N_1152);
and U1201 (N_1201,N_1194,N_1174);
and U1202 (N_1202,N_1179,N_1164);
or U1203 (N_1203,N_1151,N_1147);
or U1204 (N_1204,N_1160,N_1163);
or U1205 (N_1205,N_1180,N_1143);
nand U1206 (N_1206,N_1150,N_1178);
and U1207 (N_1207,N_1181,N_1198);
or U1208 (N_1208,N_1159,N_1193);
nor U1209 (N_1209,N_1196,N_1182);
and U1210 (N_1210,N_1191,N_1162);
xor U1211 (N_1211,N_1187,N_1173);
or U1212 (N_1212,N_1177,N_1171);
or U1213 (N_1213,N_1145,N_1195);
or U1214 (N_1214,N_1175,N_1183);
nor U1215 (N_1215,N_1157,N_1144);
nand U1216 (N_1216,N_1185,N_1161);
or U1217 (N_1217,N_1142,N_1140);
or U1218 (N_1218,N_1149,N_1148);
and U1219 (N_1219,N_1186,N_1172);
nand U1220 (N_1220,N_1158,N_1188);
and U1221 (N_1221,N_1184,N_1154);
nor U1222 (N_1222,N_1199,N_1197);
and U1223 (N_1223,N_1167,N_1166);
nor U1224 (N_1224,N_1155,N_1141);
or U1225 (N_1225,N_1146,N_1189);
or U1226 (N_1226,N_1190,N_1156);
nor U1227 (N_1227,N_1192,N_1170);
and U1228 (N_1228,N_1165,N_1176);
or U1229 (N_1229,N_1153,N_1169);
or U1230 (N_1230,N_1183,N_1184);
xor U1231 (N_1231,N_1156,N_1151);
nand U1232 (N_1232,N_1199,N_1172);
and U1233 (N_1233,N_1193,N_1192);
and U1234 (N_1234,N_1174,N_1166);
or U1235 (N_1235,N_1158,N_1176);
and U1236 (N_1236,N_1163,N_1157);
and U1237 (N_1237,N_1171,N_1149);
nand U1238 (N_1238,N_1154,N_1198);
and U1239 (N_1239,N_1189,N_1151);
nand U1240 (N_1240,N_1186,N_1198);
nor U1241 (N_1241,N_1147,N_1177);
nand U1242 (N_1242,N_1176,N_1196);
nand U1243 (N_1243,N_1152,N_1157);
nand U1244 (N_1244,N_1177,N_1140);
or U1245 (N_1245,N_1182,N_1167);
nor U1246 (N_1246,N_1149,N_1179);
nor U1247 (N_1247,N_1180,N_1163);
xor U1248 (N_1248,N_1146,N_1192);
nor U1249 (N_1249,N_1141,N_1147);
nor U1250 (N_1250,N_1187,N_1163);
nor U1251 (N_1251,N_1199,N_1188);
and U1252 (N_1252,N_1198,N_1177);
and U1253 (N_1253,N_1193,N_1194);
nor U1254 (N_1254,N_1165,N_1161);
nand U1255 (N_1255,N_1164,N_1189);
nand U1256 (N_1256,N_1153,N_1148);
nor U1257 (N_1257,N_1187,N_1149);
nor U1258 (N_1258,N_1168,N_1174);
nor U1259 (N_1259,N_1158,N_1185);
and U1260 (N_1260,N_1230,N_1222);
nand U1261 (N_1261,N_1232,N_1210);
nor U1262 (N_1262,N_1229,N_1221);
nand U1263 (N_1263,N_1252,N_1231);
or U1264 (N_1264,N_1242,N_1203);
or U1265 (N_1265,N_1225,N_1256);
nor U1266 (N_1266,N_1238,N_1208);
nor U1267 (N_1267,N_1228,N_1202);
nor U1268 (N_1268,N_1255,N_1246);
and U1269 (N_1269,N_1245,N_1209);
and U1270 (N_1270,N_1223,N_1211);
nor U1271 (N_1271,N_1207,N_1244);
and U1272 (N_1272,N_1254,N_1248);
and U1273 (N_1273,N_1234,N_1206);
nor U1274 (N_1274,N_1220,N_1215);
nand U1275 (N_1275,N_1235,N_1205);
nor U1276 (N_1276,N_1251,N_1247);
or U1277 (N_1277,N_1236,N_1216);
nor U1278 (N_1278,N_1241,N_1219);
or U1279 (N_1279,N_1212,N_1259);
nor U1280 (N_1280,N_1224,N_1201);
and U1281 (N_1281,N_1249,N_1214);
nor U1282 (N_1282,N_1227,N_1200);
or U1283 (N_1283,N_1237,N_1217);
nor U1284 (N_1284,N_1204,N_1257);
or U1285 (N_1285,N_1213,N_1243);
or U1286 (N_1286,N_1250,N_1233);
and U1287 (N_1287,N_1226,N_1258);
nor U1288 (N_1288,N_1239,N_1253);
nor U1289 (N_1289,N_1240,N_1218);
and U1290 (N_1290,N_1226,N_1200);
nor U1291 (N_1291,N_1219,N_1211);
nand U1292 (N_1292,N_1234,N_1253);
nand U1293 (N_1293,N_1218,N_1220);
or U1294 (N_1294,N_1240,N_1213);
or U1295 (N_1295,N_1235,N_1221);
or U1296 (N_1296,N_1219,N_1212);
nor U1297 (N_1297,N_1202,N_1227);
and U1298 (N_1298,N_1246,N_1211);
and U1299 (N_1299,N_1247,N_1213);
nand U1300 (N_1300,N_1252,N_1227);
and U1301 (N_1301,N_1244,N_1234);
and U1302 (N_1302,N_1249,N_1207);
nand U1303 (N_1303,N_1203,N_1246);
or U1304 (N_1304,N_1243,N_1235);
nand U1305 (N_1305,N_1235,N_1245);
or U1306 (N_1306,N_1202,N_1240);
nand U1307 (N_1307,N_1247,N_1223);
and U1308 (N_1308,N_1239,N_1256);
xnor U1309 (N_1309,N_1208,N_1212);
nand U1310 (N_1310,N_1220,N_1247);
nand U1311 (N_1311,N_1202,N_1257);
nand U1312 (N_1312,N_1213,N_1253);
and U1313 (N_1313,N_1258,N_1209);
and U1314 (N_1314,N_1207,N_1205);
nand U1315 (N_1315,N_1201,N_1216);
nand U1316 (N_1316,N_1250,N_1222);
and U1317 (N_1317,N_1204,N_1258);
and U1318 (N_1318,N_1240,N_1232);
and U1319 (N_1319,N_1241,N_1240);
nand U1320 (N_1320,N_1267,N_1316);
nor U1321 (N_1321,N_1260,N_1295);
or U1322 (N_1322,N_1299,N_1284);
nor U1323 (N_1323,N_1262,N_1281);
nor U1324 (N_1324,N_1308,N_1268);
nor U1325 (N_1325,N_1301,N_1274);
and U1326 (N_1326,N_1303,N_1311);
or U1327 (N_1327,N_1314,N_1273);
or U1328 (N_1328,N_1271,N_1315);
and U1329 (N_1329,N_1285,N_1309);
nor U1330 (N_1330,N_1287,N_1288);
or U1331 (N_1331,N_1300,N_1317);
nor U1332 (N_1332,N_1283,N_1275);
nand U1333 (N_1333,N_1294,N_1269);
and U1334 (N_1334,N_1261,N_1263);
nor U1335 (N_1335,N_1270,N_1305);
and U1336 (N_1336,N_1318,N_1307);
nor U1337 (N_1337,N_1292,N_1319);
or U1338 (N_1338,N_1291,N_1297);
or U1339 (N_1339,N_1279,N_1277);
and U1340 (N_1340,N_1290,N_1266);
nand U1341 (N_1341,N_1312,N_1265);
or U1342 (N_1342,N_1286,N_1276);
and U1343 (N_1343,N_1278,N_1280);
nand U1344 (N_1344,N_1296,N_1304);
nor U1345 (N_1345,N_1282,N_1272);
nand U1346 (N_1346,N_1289,N_1310);
or U1347 (N_1347,N_1264,N_1302);
nor U1348 (N_1348,N_1293,N_1306);
nor U1349 (N_1349,N_1313,N_1298);
and U1350 (N_1350,N_1285,N_1296);
and U1351 (N_1351,N_1287,N_1289);
nand U1352 (N_1352,N_1313,N_1300);
and U1353 (N_1353,N_1267,N_1290);
and U1354 (N_1354,N_1307,N_1293);
and U1355 (N_1355,N_1284,N_1291);
and U1356 (N_1356,N_1263,N_1291);
or U1357 (N_1357,N_1272,N_1315);
or U1358 (N_1358,N_1269,N_1309);
and U1359 (N_1359,N_1276,N_1275);
nand U1360 (N_1360,N_1311,N_1286);
nor U1361 (N_1361,N_1316,N_1283);
nand U1362 (N_1362,N_1302,N_1305);
and U1363 (N_1363,N_1265,N_1296);
nand U1364 (N_1364,N_1295,N_1314);
nor U1365 (N_1365,N_1272,N_1266);
and U1366 (N_1366,N_1293,N_1283);
or U1367 (N_1367,N_1293,N_1269);
or U1368 (N_1368,N_1304,N_1315);
and U1369 (N_1369,N_1260,N_1301);
nand U1370 (N_1370,N_1280,N_1300);
nor U1371 (N_1371,N_1263,N_1306);
nand U1372 (N_1372,N_1303,N_1305);
nand U1373 (N_1373,N_1311,N_1315);
or U1374 (N_1374,N_1299,N_1273);
and U1375 (N_1375,N_1301,N_1292);
nand U1376 (N_1376,N_1275,N_1297);
or U1377 (N_1377,N_1304,N_1295);
and U1378 (N_1378,N_1317,N_1312);
nor U1379 (N_1379,N_1266,N_1309);
nand U1380 (N_1380,N_1338,N_1326);
or U1381 (N_1381,N_1357,N_1350);
nor U1382 (N_1382,N_1362,N_1361);
nor U1383 (N_1383,N_1367,N_1327);
and U1384 (N_1384,N_1343,N_1377);
or U1385 (N_1385,N_1322,N_1331);
and U1386 (N_1386,N_1368,N_1345);
nand U1387 (N_1387,N_1333,N_1323);
nand U1388 (N_1388,N_1370,N_1352);
or U1389 (N_1389,N_1337,N_1363);
nor U1390 (N_1390,N_1373,N_1360);
or U1391 (N_1391,N_1359,N_1348);
nand U1392 (N_1392,N_1369,N_1379);
and U1393 (N_1393,N_1324,N_1372);
and U1394 (N_1394,N_1332,N_1328);
and U1395 (N_1395,N_1335,N_1341);
nor U1396 (N_1396,N_1325,N_1346);
and U1397 (N_1397,N_1351,N_1320);
nand U1398 (N_1398,N_1354,N_1340);
and U1399 (N_1399,N_1353,N_1365);
and U1400 (N_1400,N_1330,N_1356);
nor U1401 (N_1401,N_1349,N_1347);
nor U1402 (N_1402,N_1376,N_1374);
or U1403 (N_1403,N_1336,N_1355);
and U1404 (N_1404,N_1358,N_1364);
nand U1405 (N_1405,N_1342,N_1375);
xor U1406 (N_1406,N_1344,N_1321);
nand U1407 (N_1407,N_1366,N_1371);
nor U1408 (N_1408,N_1378,N_1339);
nor U1409 (N_1409,N_1329,N_1334);
and U1410 (N_1410,N_1324,N_1330);
and U1411 (N_1411,N_1351,N_1326);
nand U1412 (N_1412,N_1332,N_1336);
or U1413 (N_1413,N_1343,N_1361);
nor U1414 (N_1414,N_1356,N_1365);
nor U1415 (N_1415,N_1324,N_1334);
nor U1416 (N_1416,N_1371,N_1335);
nand U1417 (N_1417,N_1360,N_1320);
nand U1418 (N_1418,N_1342,N_1322);
or U1419 (N_1419,N_1348,N_1323);
and U1420 (N_1420,N_1327,N_1357);
nand U1421 (N_1421,N_1340,N_1322);
or U1422 (N_1422,N_1351,N_1368);
and U1423 (N_1423,N_1376,N_1322);
or U1424 (N_1424,N_1347,N_1351);
xnor U1425 (N_1425,N_1341,N_1324);
or U1426 (N_1426,N_1336,N_1373);
and U1427 (N_1427,N_1349,N_1367);
or U1428 (N_1428,N_1376,N_1344);
and U1429 (N_1429,N_1361,N_1360);
nand U1430 (N_1430,N_1354,N_1375);
nor U1431 (N_1431,N_1358,N_1344);
or U1432 (N_1432,N_1344,N_1348);
nand U1433 (N_1433,N_1345,N_1350);
nor U1434 (N_1434,N_1335,N_1345);
nor U1435 (N_1435,N_1367,N_1378);
nand U1436 (N_1436,N_1345,N_1369);
nor U1437 (N_1437,N_1346,N_1365);
or U1438 (N_1438,N_1320,N_1326);
nand U1439 (N_1439,N_1379,N_1331);
nand U1440 (N_1440,N_1427,N_1410);
nand U1441 (N_1441,N_1424,N_1397);
and U1442 (N_1442,N_1401,N_1385);
nor U1443 (N_1443,N_1409,N_1439);
nor U1444 (N_1444,N_1416,N_1393);
nor U1445 (N_1445,N_1384,N_1413);
and U1446 (N_1446,N_1436,N_1399);
or U1447 (N_1447,N_1387,N_1415);
and U1448 (N_1448,N_1419,N_1433);
nor U1449 (N_1449,N_1435,N_1438);
nor U1450 (N_1450,N_1389,N_1432);
nand U1451 (N_1451,N_1404,N_1411);
and U1452 (N_1452,N_1390,N_1400);
nand U1453 (N_1453,N_1429,N_1434);
or U1454 (N_1454,N_1380,N_1414);
and U1455 (N_1455,N_1386,N_1388);
or U1456 (N_1456,N_1423,N_1422);
or U1457 (N_1457,N_1437,N_1407);
nand U1458 (N_1458,N_1405,N_1381);
nor U1459 (N_1459,N_1382,N_1391);
or U1460 (N_1460,N_1425,N_1421);
or U1461 (N_1461,N_1395,N_1426);
nor U1462 (N_1462,N_1417,N_1412);
and U1463 (N_1463,N_1396,N_1402);
and U1464 (N_1464,N_1398,N_1431);
or U1465 (N_1465,N_1408,N_1394);
nand U1466 (N_1466,N_1392,N_1430);
or U1467 (N_1467,N_1418,N_1403);
and U1468 (N_1468,N_1406,N_1420);
nand U1469 (N_1469,N_1428,N_1383);
or U1470 (N_1470,N_1431,N_1381);
and U1471 (N_1471,N_1424,N_1384);
nor U1472 (N_1472,N_1383,N_1414);
and U1473 (N_1473,N_1402,N_1414);
nor U1474 (N_1474,N_1415,N_1395);
nor U1475 (N_1475,N_1431,N_1387);
nand U1476 (N_1476,N_1415,N_1404);
or U1477 (N_1477,N_1409,N_1385);
and U1478 (N_1478,N_1437,N_1405);
and U1479 (N_1479,N_1437,N_1422);
and U1480 (N_1480,N_1380,N_1404);
and U1481 (N_1481,N_1401,N_1411);
or U1482 (N_1482,N_1426,N_1430);
or U1483 (N_1483,N_1415,N_1410);
nor U1484 (N_1484,N_1395,N_1422);
and U1485 (N_1485,N_1435,N_1414);
or U1486 (N_1486,N_1385,N_1426);
and U1487 (N_1487,N_1426,N_1437);
and U1488 (N_1488,N_1405,N_1397);
or U1489 (N_1489,N_1420,N_1391);
or U1490 (N_1490,N_1415,N_1437);
or U1491 (N_1491,N_1416,N_1424);
or U1492 (N_1492,N_1414,N_1425);
nor U1493 (N_1493,N_1420,N_1427);
xor U1494 (N_1494,N_1438,N_1383);
or U1495 (N_1495,N_1420,N_1395);
nand U1496 (N_1496,N_1412,N_1433);
and U1497 (N_1497,N_1399,N_1398);
nand U1498 (N_1498,N_1388,N_1400);
nand U1499 (N_1499,N_1406,N_1419);
nor U1500 (N_1500,N_1446,N_1480);
xnor U1501 (N_1501,N_1445,N_1465);
xnor U1502 (N_1502,N_1483,N_1440);
or U1503 (N_1503,N_1452,N_1479);
nand U1504 (N_1504,N_1495,N_1494);
nor U1505 (N_1505,N_1449,N_1472);
or U1506 (N_1506,N_1475,N_1498);
and U1507 (N_1507,N_1459,N_1453);
or U1508 (N_1508,N_1471,N_1469);
nor U1509 (N_1509,N_1473,N_1461);
or U1510 (N_1510,N_1474,N_1456);
nand U1511 (N_1511,N_1477,N_1493);
nor U1512 (N_1512,N_1450,N_1488);
nor U1513 (N_1513,N_1476,N_1484);
nor U1514 (N_1514,N_1467,N_1485);
nor U1515 (N_1515,N_1444,N_1447);
nor U1516 (N_1516,N_1490,N_1482);
nor U1517 (N_1517,N_1455,N_1499);
nor U1518 (N_1518,N_1466,N_1468);
nand U1519 (N_1519,N_1491,N_1486);
nand U1520 (N_1520,N_1454,N_1489);
xnor U1521 (N_1521,N_1441,N_1492);
nor U1522 (N_1522,N_1464,N_1442);
and U1523 (N_1523,N_1470,N_1496);
nand U1524 (N_1524,N_1497,N_1443);
and U1525 (N_1525,N_1448,N_1463);
and U1526 (N_1526,N_1481,N_1457);
and U1527 (N_1527,N_1460,N_1451);
or U1528 (N_1528,N_1487,N_1462);
or U1529 (N_1529,N_1458,N_1478);
nand U1530 (N_1530,N_1450,N_1442);
nor U1531 (N_1531,N_1468,N_1485);
and U1532 (N_1532,N_1463,N_1454);
nand U1533 (N_1533,N_1449,N_1446);
or U1534 (N_1534,N_1455,N_1444);
nor U1535 (N_1535,N_1458,N_1491);
or U1536 (N_1536,N_1474,N_1482);
nor U1537 (N_1537,N_1498,N_1491);
nor U1538 (N_1538,N_1496,N_1478);
or U1539 (N_1539,N_1485,N_1480);
nand U1540 (N_1540,N_1459,N_1475);
nand U1541 (N_1541,N_1465,N_1459);
and U1542 (N_1542,N_1480,N_1450);
and U1543 (N_1543,N_1473,N_1478);
nand U1544 (N_1544,N_1453,N_1475);
nor U1545 (N_1545,N_1470,N_1479);
and U1546 (N_1546,N_1477,N_1475);
nor U1547 (N_1547,N_1474,N_1498);
nor U1548 (N_1548,N_1460,N_1463);
and U1549 (N_1549,N_1474,N_1497);
and U1550 (N_1550,N_1441,N_1489);
nand U1551 (N_1551,N_1484,N_1479);
nor U1552 (N_1552,N_1457,N_1453);
or U1553 (N_1553,N_1460,N_1454);
nor U1554 (N_1554,N_1473,N_1453);
and U1555 (N_1555,N_1449,N_1445);
nand U1556 (N_1556,N_1489,N_1456);
nand U1557 (N_1557,N_1487,N_1457);
or U1558 (N_1558,N_1492,N_1461);
nor U1559 (N_1559,N_1487,N_1467);
and U1560 (N_1560,N_1510,N_1548);
nand U1561 (N_1561,N_1554,N_1556);
and U1562 (N_1562,N_1506,N_1502);
nand U1563 (N_1563,N_1518,N_1528);
or U1564 (N_1564,N_1511,N_1516);
and U1565 (N_1565,N_1536,N_1533);
nor U1566 (N_1566,N_1524,N_1553);
or U1567 (N_1567,N_1501,N_1547);
and U1568 (N_1568,N_1549,N_1525);
and U1569 (N_1569,N_1522,N_1517);
or U1570 (N_1570,N_1526,N_1531);
nand U1571 (N_1571,N_1544,N_1551);
nand U1572 (N_1572,N_1535,N_1541);
nor U1573 (N_1573,N_1540,N_1557);
nand U1574 (N_1574,N_1539,N_1552);
nor U1575 (N_1575,N_1508,N_1529);
nor U1576 (N_1576,N_1512,N_1519);
nor U1577 (N_1577,N_1545,N_1555);
and U1578 (N_1578,N_1558,N_1542);
or U1579 (N_1579,N_1513,N_1514);
and U1580 (N_1580,N_1537,N_1503);
and U1581 (N_1581,N_1505,N_1507);
nor U1582 (N_1582,N_1500,N_1543);
nand U1583 (N_1583,N_1538,N_1520);
nor U1584 (N_1584,N_1530,N_1521);
and U1585 (N_1585,N_1550,N_1527);
or U1586 (N_1586,N_1509,N_1534);
nand U1587 (N_1587,N_1532,N_1523);
nor U1588 (N_1588,N_1546,N_1559);
nor U1589 (N_1589,N_1504,N_1515);
nand U1590 (N_1590,N_1554,N_1551);
nor U1591 (N_1591,N_1540,N_1533);
or U1592 (N_1592,N_1556,N_1525);
nand U1593 (N_1593,N_1521,N_1524);
and U1594 (N_1594,N_1518,N_1542);
nand U1595 (N_1595,N_1559,N_1504);
nand U1596 (N_1596,N_1549,N_1559);
nor U1597 (N_1597,N_1518,N_1529);
nand U1598 (N_1598,N_1547,N_1523);
nor U1599 (N_1599,N_1504,N_1516);
or U1600 (N_1600,N_1500,N_1531);
and U1601 (N_1601,N_1504,N_1529);
or U1602 (N_1602,N_1516,N_1558);
and U1603 (N_1603,N_1526,N_1537);
nor U1604 (N_1604,N_1512,N_1505);
and U1605 (N_1605,N_1520,N_1554);
nor U1606 (N_1606,N_1515,N_1501);
nor U1607 (N_1607,N_1514,N_1554);
nor U1608 (N_1608,N_1503,N_1541);
nand U1609 (N_1609,N_1521,N_1504);
or U1610 (N_1610,N_1535,N_1509);
and U1611 (N_1611,N_1501,N_1518);
and U1612 (N_1612,N_1543,N_1503);
nand U1613 (N_1613,N_1500,N_1505);
or U1614 (N_1614,N_1541,N_1554);
nand U1615 (N_1615,N_1519,N_1522);
nand U1616 (N_1616,N_1520,N_1529);
nand U1617 (N_1617,N_1553,N_1506);
nand U1618 (N_1618,N_1556,N_1504);
and U1619 (N_1619,N_1531,N_1553);
or U1620 (N_1620,N_1603,N_1566);
nor U1621 (N_1621,N_1601,N_1611);
or U1622 (N_1622,N_1616,N_1573);
nor U1623 (N_1623,N_1599,N_1590);
or U1624 (N_1624,N_1585,N_1568);
or U1625 (N_1625,N_1600,N_1577);
or U1626 (N_1626,N_1607,N_1589);
nor U1627 (N_1627,N_1579,N_1564);
nor U1628 (N_1628,N_1612,N_1560);
and U1629 (N_1629,N_1615,N_1609);
nand U1630 (N_1630,N_1576,N_1593);
or U1631 (N_1631,N_1596,N_1597);
and U1632 (N_1632,N_1581,N_1582);
nand U1633 (N_1633,N_1604,N_1569);
nor U1634 (N_1634,N_1578,N_1591);
nand U1635 (N_1635,N_1610,N_1617);
nand U1636 (N_1636,N_1588,N_1563);
nor U1637 (N_1637,N_1614,N_1574);
nor U1638 (N_1638,N_1592,N_1567);
nor U1639 (N_1639,N_1618,N_1598);
nor U1640 (N_1640,N_1594,N_1605);
nor U1641 (N_1641,N_1584,N_1570);
nand U1642 (N_1642,N_1608,N_1561);
nor U1643 (N_1643,N_1572,N_1580);
nor U1644 (N_1644,N_1587,N_1571);
or U1645 (N_1645,N_1583,N_1562);
or U1646 (N_1646,N_1613,N_1575);
or U1647 (N_1647,N_1565,N_1606);
or U1648 (N_1648,N_1602,N_1619);
nor U1649 (N_1649,N_1586,N_1595);
nand U1650 (N_1650,N_1595,N_1561);
and U1651 (N_1651,N_1587,N_1613);
and U1652 (N_1652,N_1591,N_1617);
nor U1653 (N_1653,N_1599,N_1619);
and U1654 (N_1654,N_1619,N_1579);
nor U1655 (N_1655,N_1614,N_1586);
and U1656 (N_1656,N_1592,N_1591);
nor U1657 (N_1657,N_1574,N_1591);
or U1658 (N_1658,N_1599,N_1611);
and U1659 (N_1659,N_1588,N_1580);
or U1660 (N_1660,N_1612,N_1573);
and U1661 (N_1661,N_1580,N_1589);
nand U1662 (N_1662,N_1576,N_1586);
nand U1663 (N_1663,N_1574,N_1599);
nor U1664 (N_1664,N_1596,N_1589);
nand U1665 (N_1665,N_1594,N_1586);
nor U1666 (N_1666,N_1595,N_1589);
nand U1667 (N_1667,N_1608,N_1594);
nand U1668 (N_1668,N_1576,N_1613);
or U1669 (N_1669,N_1571,N_1616);
or U1670 (N_1670,N_1592,N_1613);
and U1671 (N_1671,N_1560,N_1611);
and U1672 (N_1672,N_1566,N_1611);
nand U1673 (N_1673,N_1575,N_1583);
xor U1674 (N_1674,N_1614,N_1565);
and U1675 (N_1675,N_1611,N_1600);
nor U1676 (N_1676,N_1564,N_1585);
or U1677 (N_1677,N_1609,N_1605);
nor U1678 (N_1678,N_1590,N_1613);
nor U1679 (N_1679,N_1597,N_1611);
and U1680 (N_1680,N_1629,N_1637);
or U1681 (N_1681,N_1674,N_1641);
nor U1682 (N_1682,N_1638,N_1649);
or U1683 (N_1683,N_1634,N_1678);
nand U1684 (N_1684,N_1670,N_1679);
nor U1685 (N_1685,N_1625,N_1665);
and U1686 (N_1686,N_1676,N_1653);
nor U1687 (N_1687,N_1640,N_1660);
nor U1688 (N_1688,N_1623,N_1650);
nor U1689 (N_1689,N_1672,N_1632);
or U1690 (N_1690,N_1668,N_1661);
and U1691 (N_1691,N_1666,N_1633);
nand U1692 (N_1692,N_1642,N_1651);
nand U1693 (N_1693,N_1658,N_1624);
and U1694 (N_1694,N_1621,N_1626);
nand U1695 (N_1695,N_1652,N_1627);
and U1696 (N_1696,N_1635,N_1645);
nor U1697 (N_1697,N_1648,N_1669);
nor U1698 (N_1698,N_1664,N_1644);
nand U1699 (N_1699,N_1662,N_1631);
or U1700 (N_1700,N_1663,N_1655);
nand U1701 (N_1701,N_1677,N_1671);
nor U1702 (N_1702,N_1620,N_1630);
or U1703 (N_1703,N_1667,N_1628);
nand U1704 (N_1704,N_1639,N_1636);
nand U1705 (N_1705,N_1656,N_1659);
nand U1706 (N_1706,N_1646,N_1654);
and U1707 (N_1707,N_1657,N_1673);
nor U1708 (N_1708,N_1643,N_1675);
or U1709 (N_1709,N_1622,N_1647);
nor U1710 (N_1710,N_1646,N_1652);
or U1711 (N_1711,N_1662,N_1651);
and U1712 (N_1712,N_1658,N_1629);
nand U1713 (N_1713,N_1653,N_1670);
and U1714 (N_1714,N_1649,N_1637);
nand U1715 (N_1715,N_1649,N_1623);
or U1716 (N_1716,N_1657,N_1653);
and U1717 (N_1717,N_1622,N_1620);
nor U1718 (N_1718,N_1643,N_1662);
nand U1719 (N_1719,N_1665,N_1632);
or U1720 (N_1720,N_1661,N_1625);
nor U1721 (N_1721,N_1679,N_1663);
nand U1722 (N_1722,N_1659,N_1635);
and U1723 (N_1723,N_1622,N_1653);
or U1724 (N_1724,N_1656,N_1674);
nor U1725 (N_1725,N_1657,N_1640);
or U1726 (N_1726,N_1637,N_1627);
and U1727 (N_1727,N_1636,N_1646);
xnor U1728 (N_1728,N_1637,N_1654);
and U1729 (N_1729,N_1638,N_1650);
nor U1730 (N_1730,N_1644,N_1646);
or U1731 (N_1731,N_1660,N_1639);
and U1732 (N_1732,N_1664,N_1621);
nand U1733 (N_1733,N_1623,N_1658);
and U1734 (N_1734,N_1627,N_1678);
nand U1735 (N_1735,N_1673,N_1625);
or U1736 (N_1736,N_1665,N_1644);
or U1737 (N_1737,N_1644,N_1660);
nand U1738 (N_1738,N_1630,N_1640);
nor U1739 (N_1739,N_1630,N_1653);
nor U1740 (N_1740,N_1681,N_1715);
and U1741 (N_1741,N_1682,N_1728);
or U1742 (N_1742,N_1698,N_1687);
nand U1743 (N_1743,N_1720,N_1690);
nor U1744 (N_1744,N_1738,N_1732);
or U1745 (N_1745,N_1694,N_1688);
or U1746 (N_1746,N_1706,N_1729);
nor U1747 (N_1747,N_1691,N_1703);
and U1748 (N_1748,N_1700,N_1734);
nor U1749 (N_1749,N_1718,N_1726);
nand U1750 (N_1750,N_1714,N_1719);
nor U1751 (N_1751,N_1705,N_1696);
nor U1752 (N_1752,N_1685,N_1733);
nand U1753 (N_1753,N_1724,N_1725);
nand U1754 (N_1754,N_1739,N_1727);
or U1755 (N_1755,N_1683,N_1717);
nand U1756 (N_1756,N_1710,N_1692);
nor U1757 (N_1757,N_1735,N_1702);
xor U1758 (N_1758,N_1680,N_1711);
nor U1759 (N_1759,N_1716,N_1736);
nand U1760 (N_1760,N_1695,N_1713);
nand U1761 (N_1761,N_1730,N_1722);
and U1762 (N_1762,N_1731,N_1708);
nand U1763 (N_1763,N_1721,N_1704);
nor U1764 (N_1764,N_1697,N_1699);
nor U1765 (N_1765,N_1689,N_1712);
and U1766 (N_1766,N_1723,N_1684);
nand U1767 (N_1767,N_1737,N_1693);
or U1768 (N_1768,N_1709,N_1707);
nand U1769 (N_1769,N_1686,N_1701);
or U1770 (N_1770,N_1710,N_1698);
nand U1771 (N_1771,N_1715,N_1735);
nand U1772 (N_1772,N_1684,N_1704);
nor U1773 (N_1773,N_1717,N_1728);
or U1774 (N_1774,N_1733,N_1706);
and U1775 (N_1775,N_1724,N_1709);
nor U1776 (N_1776,N_1725,N_1723);
nand U1777 (N_1777,N_1727,N_1685);
and U1778 (N_1778,N_1680,N_1723);
and U1779 (N_1779,N_1731,N_1739);
xnor U1780 (N_1780,N_1696,N_1681);
nor U1781 (N_1781,N_1692,N_1727);
nand U1782 (N_1782,N_1718,N_1683);
nand U1783 (N_1783,N_1739,N_1713);
or U1784 (N_1784,N_1725,N_1718);
nor U1785 (N_1785,N_1701,N_1683);
or U1786 (N_1786,N_1733,N_1693);
nand U1787 (N_1787,N_1694,N_1714);
nand U1788 (N_1788,N_1733,N_1719);
or U1789 (N_1789,N_1722,N_1693);
nor U1790 (N_1790,N_1685,N_1713);
or U1791 (N_1791,N_1700,N_1716);
or U1792 (N_1792,N_1705,N_1698);
nand U1793 (N_1793,N_1722,N_1728);
nor U1794 (N_1794,N_1708,N_1697);
nor U1795 (N_1795,N_1713,N_1735);
nand U1796 (N_1796,N_1702,N_1721);
nor U1797 (N_1797,N_1707,N_1691);
nand U1798 (N_1798,N_1729,N_1724);
nand U1799 (N_1799,N_1682,N_1708);
nor U1800 (N_1800,N_1748,N_1766);
nor U1801 (N_1801,N_1741,N_1798);
nor U1802 (N_1802,N_1753,N_1762);
nand U1803 (N_1803,N_1797,N_1789);
nor U1804 (N_1804,N_1774,N_1767);
and U1805 (N_1805,N_1799,N_1745);
nand U1806 (N_1806,N_1764,N_1749);
and U1807 (N_1807,N_1781,N_1785);
or U1808 (N_1808,N_1787,N_1765);
or U1809 (N_1809,N_1754,N_1791);
nand U1810 (N_1810,N_1757,N_1776);
nor U1811 (N_1811,N_1777,N_1790);
and U1812 (N_1812,N_1763,N_1769);
nor U1813 (N_1813,N_1775,N_1788);
or U1814 (N_1814,N_1759,N_1743);
nand U1815 (N_1815,N_1751,N_1758);
nand U1816 (N_1816,N_1750,N_1770);
nand U1817 (N_1817,N_1752,N_1795);
or U1818 (N_1818,N_1744,N_1792);
nor U1819 (N_1819,N_1756,N_1780);
nand U1820 (N_1820,N_1783,N_1772);
or U1821 (N_1821,N_1796,N_1782);
nand U1822 (N_1822,N_1740,N_1786);
nand U1823 (N_1823,N_1784,N_1779);
nand U1824 (N_1824,N_1773,N_1746);
and U1825 (N_1825,N_1793,N_1747);
or U1826 (N_1826,N_1742,N_1760);
and U1827 (N_1827,N_1768,N_1794);
or U1828 (N_1828,N_1755,N_1778);
or U1829 (N_1829,N_1761,N_1771);
nand U1830 (N_1830,N_1787,N_1792);
nand U1831 (N_1831,N_1784,N_1756);
nor U1832 (N_1832,N_1794,N_1789);
nand U1833 (N_1833,N_1749,N_1760);
or U1834 (N_1834,N_1794,N_1776);
or U1835 (N_1835,N_1754,N_1792);
nand U1836 (N_1836,N_1799,N_1779);
or U1837 (N_1837,N_1759,N_1790);
nand U1838 (N_1838,N_1788,N_1799);
and U1839 (N_1839,N_1746,N_1750);
or U1840 (N_1840,N_1799,N_1778);
and U1841 (N_1841,N_1769,N_1770);
nor U1842 (N_1842,N_1771,N_1791);
or U1843 (N_1843,N_1799,N_1768);
or U1844 (N_1844,N_1748,N_1776);
and U1845 (N_1845,N_1774,N_1795);
nand U1846 (N_1846,N_1786,N_1741);
or U1847 (N_1847,N_1780,N_1761);
xnor U1848 (N_1848,N_1785,N_1788);
nor U1849 (N_1849,N_1768,N_1742);
nand U1850 (N_1850,N_1759,N_1794);
and U1851 (N_1851,N_1775,N_1751);
and U1852 (N_1852,N_1751,N_1746);
nor U1853 (N_1853,N_1795,N_1751);
nand U1854 (N_1854,N_1751,N_1744);
and U1855 (N_1855,N_1764,N_1795);
nor U1856 (N_1856,N_1776,N_1796);
nor U1857 (N_1857,N_1785,N_1777);
and U1858 (N_1858,N_1775,N_1755);
and U1859 (N_1859,N_1781,N_1790);
and U1860 (N_1860,N_1806,N_1848);
or U1861 (N_1861,N_1824,N_1819);
and U1862 (N_1862,N_1803,N_1809);
nor U1863 (N_1863,N_1802,N_1800);
nand U1864 (N_1864,N_1854,N_1823);
and U1865 (N_1865,N_1804,N_1801);
or U1866 (N_1866,N_1846,N_1816);
nand U1867 (N_1867,N_1839,N_1855);
nor U1868 (N_1868,N_1858,N_1838);
nor U1869 (N_1869,N_1812,N_1832);
nand U1870 (N_1870,N_1821,N_1851);
nand U1871 (N_1871,N_1840,N_1825);
and U1872 (N_1872,N_1818,N_1817);
nor U1873 (N_1873,N_1847,N_1859);
nand U1874 (N_1874,N_1811,N_1852);
nor U1875 (N_1875,N_1835,N_1836);
nand U1876 (N_1876,N_1829,N_1810);
nor U1877 (N_1877,N_1826,N_1837);
and U1878 (N_1878,N_1833,N_1827);
and U1879 (N_1879,N_1845,N_1834);
and U1880 (N_1880,N_1853,N_1857);
nor U1881 (N_1881,N_1822,N_1830);
nand U1882 (N_1882,N_1842,N_1841);
or U1883 (N_1883,N_1807,N_1820);
and U1884 (N_1884,N_1856,N_1831);
nand U1885 (N_1885,N_1815,N_1844);
nand U1886 (N_1886,N_1808,N_1828);
or U1887 (N_1887,N_1805,N_1843);
nand U1888 (N_1888,N_1850,N_1849);
nand U1889 (N_1889,N_1814,N_1813);
and U1890 (N_1890,N_1808,N_1852);
nand U1891 (N_1891,N_1848,N_1807);
nor U1892 (N_1892,N_1842,N_1813);
nand U1893 (N_1893,N_1855,N_1829);
nor U1894 (N_1894,N_1857,N_1814);
and U1895 (N_1895,N_1859,N_1827);
nand U1896 (N_1896,N_1839,N_1846);
nor U1897 (N_1897,N_1824,N_1814);
nand U1898 (N_1898,N_1848,N_1840);
xor U1899 (N_1899,N_1837,N_1803);
nand U1900 (N_1900,N_1854,N_1807);
or U1901 (N_1901,N_1846,N_1854);
nand U1902 (N_1902,N_1829,N_1807);
or U1903 (N_1903,N_1815,N_1818);
and U1904 (N_1904,N_1803,N_1821);
nor U1905 (N_1905,N_1848,N_1842);
nand U1906 (N_1906,N_1850,N_1830);
and U1907 (N_1907,N_1811,N_1830);
nor U1908 (N_1908,N_1841,N_1830);
nor U1909 (N_1909,N_1815,N_1822);
nand U1910 (N_1910,N_1821,N_1852);
nor U1911 (N_1911,N_1824,N_1800);
and U1912 (N_1912,N_1831,N_1857);
or U1913 (N_1913,N_1819,N_1853);
or U1914 (N_1914,N_1859,N_1810);
nor U1915 (N_1915,N_1809,N_1851);
nand U1916 (N_1916,N_1813,N_1819);
and U1917 (N_1917,N_1855,N_1804);
or U1918 (N_1918,N_1810,N_1827);
and U1919 (N_1919,N_1842,N_1820);
nor U1920 (N_1920,N_1882,N_1916);
or U1921 (N_1921,N_1904,N_1907);
nand U1922 (N_1922,N_1867,N_1905);
or U1923 (N_1923,N_1886,N_1860);
nor U1924 (N_1924,N_1862,N_1887);
or U1925 (N_1925,N_1875,N_1899);
or U1926 (N_1926,N_1903,N_1911);
nand U1927 (N_1927,N_1913,N_1897);
or U1928 (N_1928,N_1892,N_1863);
or U1929 (N_1929,N_1879,N_1876);
nor U1930 (N_1930,N_1902,N_1865);
nor U1931 (N_1931,N_1910,N_1914);
nand U1932 (N_1932,N_1893,N_1866);
nor U1933 (N_1933,N_1878,N_1900);
and U1934 (N_1934,N_1891,N_1873);
nand U1935 (N_1935,N_1894,N_1880);
and U1936 (N_1936,N_1871,N_1885);
or U1937 (N_1937,N_1881,N_1872);
or U1938 (N_1938,N_1919,N_1918);
nand U1939 (N_1939,N_1917,N_1895);
nand U1940 (N_1940,N_1890,N_1889);
nor U1941 (N_1941,N_1908,N_1915);
or U1942 (N_1942,N_1901,N_1870);
nand U1943 (N_1943,N_1896,N_1874);
and U1944 (N_1944,N_1864,N_1869);
nor U1945 (N_1945,N_1861,N_1883);
or U1946 (N_1946,N_1877,N_1884);
nand U1947 (N_1947,N_1912,N_1898);
or U1948 (N_1948,N_1888,N_1906);
nand U1949 (N_1949,N_1868,N_1909);
nor U1950 (N_1950,N_1877,N_1882);
nor U1951 (N_1951,N_1904,N_1917);
nand U1952 (N_1952,N_1873,N_1872);
and U1953 (N_1953,N_1880,N_1908);
nor U1954 (N_1954,N_1899,N_1882);
nor U1955 (N_1955,N_1864,N_1898);
and U1956 (N_1956,N_1866,N_1884);
and U1957 (N_1957,N_1901,N_1914);
nand U1958 (N_1958,N_1862,N_1918);
nand U1959 (N_1959,N_1880,N_1860);
and U1960 (N_1960,N_1889,N_1918);
or U1961 (N_1961,N_1863,N_1900);
nand U1962 (N_1962,N_1865,N_1889);
or U1963 (N_1963,N_1889,N_1913);
or U1964 (N_1964,N_1906,N_1909);
or U1965 (N_1965,N_1874,N_1881);
nand U1966 (N_1966,N_1874,N_1899);
and U1967 (N_1967,N_1869,N_1897);
or U1968 (N_1968,N_1877,N_1881);
nand U1969 (N_1969,N_1873,N_1913);
and U1970 (N_1970,N_1874,N_1871);
or U1971 (N_1971,N_1887,N_1900);
nand U1972 (N_1972,N_1919,N_1885);
and U1973 (N_1973,N_1861,N_1913);
and U1974 (N_1974,N_1895,N_1915);
nor U1975 (N_1975,N_1895,N_1918);
or U1976 (N_1976,N_1913,N_1866);
and U1977 (N_1977,N_1902,N_1864);
nor U1978 (N_1978,N_1898,N_1875);
nor U1979 (N_1979,N_1861,N_1901);
and U1980 (N_1980,N_1929,N_1973);
and U1981 (N_1981,N_1969,N_1974);
nor U1982 (N_1982,N_1933,N_1928);
and U1983 (N_1983,N_1937,N_1970);
nor U1984 (N_1984,N_1930,N_1953);
nand U1985 (N_1985,N_1952,N_1941);
nor U1986 (N_1986,N_1979,N_1958);
nand U1987 (N_1987,N_1959,N_1966);
and U1988 (N_1988,N_1936,N_1932);
nand U1989 (N_1989,N_1951,N_1939);
or U1990 (N_1990,N_1947,N_1920);
or U1991 (N_1991,N_1922,N_1945);
nand U1992 (N_1992,N_1960,N_1965);
and U1993 (N_1993,N_1967,N_1971);
nand U1994 (N_1994,N_1935,N_1968);
nor U1995 (N_1995,N_1961,N_1946);
nand U1996 (N_1996,N_1963,N_1955);
nand U1997 (N_1997,N_1944,N_1954);
or U1998 (N_1998,N_1925,N_1976);
and U1999 (N_1999,N_1949,N_1938);
nor U2000 (N_2000,N_1923,N_1978);
and U2001 (N_2001,N_1972,N_1956);
nor U2002 (N_2002,N_1940,N_1942);
and U2003 (N_2003,N_1975,N_1934);
or U2004 (N_2004,N_1943,N_1921);
nand U2005 (N_2005,N_1948,N_1950);
and U2006 (N_2006,N_1927,N_1962);
nand U2007 (N_2007,N_1924,N_1977);
or U2008 (N_2008,N_1957,N_1964);
nand U2009 (N_2009,N_1931,N_1926);
nand U2010 (N_2010,N_1925,N_1975);
nor U2011 (N_2011,N_1966,N_1954);
nand U2012 (N_2012,N_1968,N_1972);
or U2013 (N_2013,N_1973,N_1922);
or U2014 (N_2014,N_1978,N_1977);
and U2015 (N_2015,N_1947,N_1972);
nor U2016 (N_2016,N_1973,N_1941);
nand U2017 (N_2017,N_1969,N_1963);
or U2018 (N_2018,N_1926,N_1941);
or U2019 (N_2019,N_1973,N_1920);
or U2020 (N_2020,N_1961,N_1979);
or U2021 (N_2021,N_1965,N_1937);
and U2022 (N_2022,N_1933,N_1967);
nor U2023 (N_2023,N_1963,N_1958);
nand U2024 (N_2024,N_1920,N_1930);
and U2025 (N_2025,N_1948,N_1944);
nand U2026 (N_2026,N_1978,N_1964);
nand U2027 (N_2027,N_1934,N_1952);
or U2028 (N_2028,N_1955,N_1934);
and U2029 (N_2029,N_1930,N_1967);
and U2030 (N_2030,N_1951,N_1959);
nand U2031 (N_2031,N_1959,N_1927);
and U2032 (N_2032,N_1935,N_1970);
nand U2033 (N_2033,N_1926,N_1971);
or U2034 (N_2034,N_1955,N_1972);
or U2035 (N_2035,N_1925,N_1954);
or U2036 (N_2036,N_1965,N_1924);
or U2037 (N_2037,N_1956,N_1959);
or U2038 (N_2038,N_1939,N_1967);
or U2039 (N_2039,N_1955,N_1921);
nand U2040 (N_2040,N_2001,N_1981);
nand U2041 (N_2041,N_1993,N_2011);
or U2042 (N_2042,N_2017,N_1991);
nor U2043 (N_2043,N_2000,N_2009);
or U2044 (N_2044,N_2012,N_1987);
or U2045 (N_2045,N_2028,N_2031);
nor U2046 (N_2046,N_2002,N_2010);
and U2047 (N_2047,N_2007,N_1985);
or U2048 (N_2048,N_2021,N_2008);
nand U2049 (N_2049,N_2016,N_1984);
and U2050 (N_2050,N_2020,N_2023);
nor U2051 (N_2051,N_2014,N_1986);
or U2052 (N_2052,N_2030,N_2024);
nor U2053 (N_2053,N_2004,N_2005);
and U2054 (N_2054,N_2015,N_1999);
or U2055 (N_2055,N_2036,N_2029);
and U2056 (N_2056,N_1997,N_1982);
or U2057 (N_2057,N_2032,N_2013);
nor U2058 (N_2058,N_2026,N_1988);
or U2059 (N_2059,N_2033,N_2022);
or U2060 (N_2060,N_1983,N_2037);
xor U2061 (N_2061,N_2019,N_1994);
and U2062 (N_2062,N_1992,N_2038);
and U2063 (N_2063,N_1980,N_2027);
nor U2064 (N_2064,N_1989,N_2025);
and U2065 (N_2065,N_2039,N_1990);
or U2066 (N_2066,N_2018,N_2034);
nor U2067 (N_2067,N_2003,N_1995);
xnor U2068 (N_2068,N_1998,N_2006);
or U2069 (N_2069,N_1996,N_2035);
or U2070 (N_2070,N_2028,N_1980);
and U2071 (N_2071,N_2020,N_2027);
and U2072 (N_2072,N_2005,N_2018);
nor U2073 (N_2073,N_1989,N_1990);
or U2074 (N_2074,N_2023,N_1987);
nor U2075 (N_2075,N_2029,N_2017);
nor U2076 (N_2076,N_2016,N_1982);
nor U2077 (N_2077,N_1996,N_1980);
nand U2078 (N_2078,N_2000,N_1999);
nor U2079 (N_2079,N_2034,N_1993);
nand U2080 (N_2080,N_2030,N_1991);
and U2081 (N_2081,N_1990,N_2021);
and U2082 (N_2082,N_1985,N_2024);
or U2083 (N_2083,N_1994,N_1983);
and U2084 (N_2084,N_2019,N_2037);
nor U2085 (N_2085,N_2033,N_2008);
or U2086 (N_2086,N_1992,N_2008);
nor U2087 (N_2087,N_1992,N_1988);
nor U2088 (N_2088,N_2026,N_2038);
nor U2089 (N_2089,N_2009,N_2039);
or U2090 (N_2090,N_1998,N_2037);
nor U2091 (N_2091,N_2015,N_2000);
nand U2092 (N_2092,N_1994,N_2015);
and U2093 (N_2093,N_2030,N_2039);
and U2094 (N_2094,N_2000,N_2007);
nor U2095 (N_2095,N_2031,N_2034);
or U2096 (N_2096,N_2009,N_1987);
and U2097 (N_2097,N_2037,N_2015);
nand U2098 (N_2098,N_2018,N_1995);
or U2099 (N_2099,N_1981,N_2038);
nor U2100 (N_2100,N_2046,N_2080);
and U2101 (N_2101,N_2089,N_2059);
or U2102 (N_2102,N_2056,N_2099);
nand U2103 (N_2103,N_2097,N_2062);
nor U2104 (N_2104,N_2068,N_2079);
or U2105 (N_2105,N_2052,N_2081);
nor U2106 (N_2106,N_2091,N_2086);
nand U2107 (N_2107,N_2042,N_2065);
or U2108 (N_2108,N_2058,N_2057);
or U2109 (N_2109,N_2077,N_2092);
and U2110 (N_2110,N_2093,N_2095);
or U2111 (N_2111,N_2041,N_2072);
nand U2112 (N_2112,N_2098,N_2073);
nand U2113 (N_2113,N_2074,N_2070);
nor U2114 (N_2114,N_2050,N_2096);
and U2115 (N_2115,N_2051,N_2083);
nand U2116 (N_2116,N_2084,N_2055);
nand U2117 (N_2117,N_2063,N_2049);
nor U2118 (N_2118,N_2078,N_2067);
nor U2119 (N_2119,N_2090,N_2082);
and U2120 (N_2120,N_2064,N_2040);
and U2121 (N_2121,N_2043,N_2044);
or U2122 (N_2122,N_2087,N_2061);
nand U2123 (N_2123,N_2069,N_2045);
or U2124 (N_2124,N_2053,N_2076);
or U2125 (N_2125,N_2088,N_2085);
nand U2126 (N_2126,N_2048,N_2094);
nand U2127 (N_2127,N_2054,N_2066);
or U2128 (N_2128,N_2075,N_2071);
nand U2129 (N_2129,N_2047,N_2060);
and U2130 (N_2130,N_2050,N_2098);
nand U2131 (N_2131,N_2046,N_2041);
nand U2132 (N_2132,N_2083,N_2098);
and U2133 (N_2133,N_2089,N_2077);
nand U2134 (N_2134,N_2052,N_2073);
nor U2135 (N_2135,N_2063,N_2064);
nor U2136 (N_2136,N_2089,N_2048);
and U2137 (N_2137,N_2072,N_2085);
nor U2138 (N_2138,N_2053,N_2066);
nor U2139 (N_2139,N_2073,N_2050);
nor U2140 (N_2140,N_2047,N_2046);
or U2141 (N_2141,N_2091,N_2085);
or U2142 (N_2142,N_2067,N_2073);
nand U2143 (N_2143,N_2078,N_2045);
and U2144 (N_2144,N_2040,N_2048);
or U2145 (N_2145,N_2097,N_2095);
nor U2146 (N_2146,N_2079,N_2070);
or U2147 (N_2147,N_2097,N_2085);
nand U2148 (N_2148,N_2075,N_2057);
nor U2149 (N_2149,N_2044,N_2048);
nor U2150 (N_2150,N_2062,N_2074);
nor U2151 (N_2151,N_2050,N_2042);
and U2152 (N_2152,N_2086,N_2057);
nand U2153 (N_2153,N_2065,N_2069);
or U2154 (N_2154,N_2047,N_2045);
nor U2155 (N_2155,N_2084,N_2064);
nor U2156 (N_2156,N_2080,N_2089);
or U2157 (N_2157,N_2085,N_2076);
or U2158 (N_2158,N_2086,N_2062);
or U2159 (N_2159,N_2055,N_2067);
nand U2160 (N_2160,N_2110,N_2127);
xor U2161 (N_2161,N_2117,N_2108);
or U2162 (N_2162,N_2120,N_2139);
nor U2163 (N_2163,N_2157,N_2155);
nor U2164 (N_2164,N_2133,N_2104);
and U2165 (N_2165,N_2105,N_2101);
nand U2166 (N_2166,N_2123,N_2134);
nand U2167 (N_2167,N_2150,N_2149);
nor U2168 (N_2168,N_2152,N_2100);
and U2169 (N_2169,N_2112,N_2115);
and U2170 (N_2170,N_2103,N_2121);
and U2171 (N_2171,N_2107,N_2116);
nand U2172 (N_2172,N_2102,N_2137);
and U2173 (N_2173,N_2132,N_2113);
nor U2174 (N_2174,N_2144,N_2111);
or U2175 (N_2175,N_2146,N_2122);
and U2176 (N_2176,N_2143,N_2129);
and U2177 (N_2177,N_2124,N_2126);
or U2178 (N_2178,N_2140,N_2119);
nor U2179 (N_2179,N_2142,N_2153);
nand U2180 (N_2180,N_2125,N_2138);
and U2181 (N_2181,N_2147,N_2151);
and U2182 (N_2182,N_2135,N_2109);
nand U2183 (N_2183,N_2154,N_2148);
nand U2184 (N_2184,N_2128,N_2159);
nor U2185 (N_2185,N_2156,N_2106);
nand U2186 (N_2186,N_2131,N_2145);
and U2187 (N_2187,N_2130,N_2141);
and U2188 (N_2188,N_2114,N_2136);
and U2189 (N_2189,N_2158,N_2118);
nor U2190 (N_2190,N_2107,N_2108);
xnor U2191 (N_2191,N_2105,N_2117);
or U2192 (N_2192,N_2102,N_2159);
nand U2193 (N_2193,N_2159,N_2103);
nor U2194 (N_2194,N_2100,N_2121);
or U2195 (N_2195,N_2115,N_2120);
or U2196 (N_2196,N_2128,N_2153);
nor U2197 (N_2197,N_2115,N_2125);
nand U2198 (N_2198,N_2112,N_2136);
and U2199 (N_2199,N_2106,N_2159);
nand U2200 (N_2200,N_2131,N_2154);
or U2201 (N_2201,N_2126,N_2105);
or U2202 (N_2202,N_2148,N_2157);
or U2203 (N_2203,N_2104,N_2132);
and U2204 (N_2204,N_2138,N_2159);
or U2205 (N_2205,N_2151,N_2101);
nand U2206 (N_2206,N_2156,N_2155);
and U2207 (N_2207,N_2153,N_2124);
nand U2208 (N_2208,N_2147,N_2114);
nor U2209 (N_2209,N_2156,N_2122);
nor U2210 (N_2210,N_2114,N_2146);
nand U2211 (N_2211,N_2138,N_2100);
nor U2212 (N_2212,N_2141,N_2119);
or U2213 (N_2213,N_2120,N_2157);
nand U2214 (N_2214,N_2100,N_2154);
and U2215 (N_2215,N_2150,N_2153);
and U2216 (N_2216,N_2152,N_2125);
or U2217 (N_2217,N_2127,N_2145);
nand U2218 (N_2218,N_2123,N_2143);
and U2219 (N_2219,N_2152,N_2151);
nand U2220 (N_2220,N_2206,N_2161);
or U2221 (N_2221,N_2180,N_2207);
nor U2222 (N_2222,N_2182,N_2205);
nor U2223 (N_2223,N_2211,N_2204);
nor U2224 (N_2224,N_2173,N_2212);
nand U2225 (N_2225,N_2195,N_2210);
and U2226 (N_2226,N_2209,N_2171);
or U2227 (N_2227,N_2213,N_2181);
or U2228 (N_2228,N_2197,N_2187);
nand U2229 (N_2229,N_2189,N_2168);
nor U2230 (N_2230,N_2178,N_2218);
nor U2231 (N_2231,N_2214,N_2183);
and U2232 (N_2232,N_2217,N_2201);
and U2233 (N_2233,N_2194,N_2166);
or U2234 (N_2234,N_2198,N_2164);
nand U2235 (N_2235,N_2193,N_2199);
or U2236 (N_2236,N_2163,N_2190);
and U2237 (N_2237,N_2203,N_2185);
nor U2238 (N_2238,N_2174,N_2184);
nor U2239 (N_2239,N_2196,N_2170);
or U2240 (N_2240,N_2167,N_2215);
nand U2241 (N_2241,N_2192,N_2177);
nor U2242 (N_2242,N_2200,N_2202);
nor U2243 (N_2243,N_2162,N_2160);
or U2244 (N_2244,N_2216,N_2176);
nand U2245 (N_2245,N_2179,N_2175);
and U2246 (N_2246,N_2172,N_2188);
and U2247 (N_2247,N_2169,N_2219);
or U2248 (N_2248,N_2165,N_2186);
nand U2249 (N_2249,N_2208,N_2191);
and U2250 (N_2250,N_2176,N_2173);
nand U2251 (N_2251,N_2163,N_2169);
nor U2252 (N_2252,N_2162,N_2165);
nand U2253 (N_2253,N_2195,N_2214);
nand U2254 (N_2254,N_2206,N_2212);
xnor U2255 (N_2255,N_2208,N_2178);
and U2256 (N_2256,N_2170,N_2197);
nor U2257 (N_2257,N_2207,N_2208);
nand U2258 (N_2258,N_2184,N_2188);
nand U2259 (N_2259,N_2219,N_2212);
and U2260 (N_2260,N_2190,N_2213);
nand U2261 (N_2261,N_2167,N_2213);
and U2262 (N_2262,N_2161,N_2219);
nand U2263 (N_2263,N_2175,N_2188);
and U2264 (N_2264,N_2163,N_2201);
and U2265 (N_2265,N_2183,N_2213);
or U2266 (N_2266,N_2163,N_2214);
nor U2267 (N_2267,N_2203,N_2169);
nor U2268 (N_2268,N_2189,N_2181);
or U2269 (N_2269,N_2161,N_2170);
or U2270 (N_2270,N_2202,N_2179);
nor U2271 (N_2271,N_2160,N_2216);
and U2272 (N_2272,N_2187,N_2162);
nor U2273 (N_2273,N_2219,N_2182);
or U2274 (N_2274,N_2219,N_2168);
nand U2275 (N_2275,N_2164,N_2197);
nand U2276 (N_2276,N_2181,N_2202);
and U2277 (N_2277,N_2207,N_2161);
or U2278 (N_2278,N_2218,N_2212);
or U2279 (N_2279,N_2203,N_2179);
nor U2280 (N_2280,N_2249,N_2240);
and U2281 (N_2281,N_2271,N_2235);
nor U2282 (N_2282,N_2279,N_2232);
or U2283 (N_2283,N_2253,N_2231);
or U2284 (N_2284,N_2242,N_2248);
nor U2285 (N_2285,N_2268,N_2220);
nand U2286 (N_2286,N_2239,N_2270);
nor U2287 (N_2287,N_2233,N_2227);
and U2288 (N_2288,N_2254,N_2269);
nor U2289 (N_2289,N_2229,N_2236);
and U2290 (N_2290,N_2277,N_2225);
and U2291 (N_2291,N_2222,N_2278);
nand U2292 (N_2292,N_2266,N_2265);
and U2293 (N_2293,N_2272,N_2246);
and U2294 (N_2294,N_2274,N_2276);
and U2295 (N_2295,N_2261,N_2238);
nor U2296 (N_2296,N_2252,N_2247);
and U2297 (N_2297,N_2250,N_2257);
or U2298 (N_2298,N_2244,N_2243);
and U2299 (N_2299,N_2267,N_2264);
or U2300 (N_2300,N_2260,N_2273);
or U2301 (N_2301,N_2245,N_2237);
nor U2302 (N_2302,N_2259,N_2241);
and U2303 (N_2303,N_2234,N_2224);
or U2304 (N_2304,N_2230,N_2262);
or U2305 (N_2305,N_2228,N_2221);
nand U2306 (N_2306,N_2226,N_2263);
nor U2307 (N_2307,N_2256,N_2251);
and U2308 (N_2308,N_2275,N_2255);
nand U2309 (N_2309,N_2258,N_2223);
nor U2310 (N_2310,N_2244,N_2247);
nor U2311 (N_2311,N_2259,N_2257);
nor U2312 (N_2312,N_2233,N_2258);
nor U2313 (N_2313,N_2262,N_2250);
nor U2314 (N_2314,N_2273,N_2230);
and U2315 (N_2315,N_2239,N_2279);
and U2316 (N_2316,N_2278,N_2226);
nand U2317 (N_2317,N_2245,N_2233);
and U2318 (N_2318,N_2236,N_2261);
and U2319 (N_2319,N_2233,N_2274);
and U2320 (N_2320,N_2258,N_2236);
or U2321 (N_2321,N_2265,N_2222);
nand U2322 (N_2322,N_2274,N_2245);
nor U2323 (N_2323,N_2249,N_2257);
and U2324 (N_2324,N_2271,N_2267);
or U2325 (N_2325,N_2230,N_2227);
nor U2326 (N_2326,N_2276,N_2256);
or U2327 (N_2327,N_2246,N_2242);
and U2328 (N_2328,N_2225,N_2251);
or U2329 (N_2329,N_2277,N_2245);
nand U2330 (N_2330,N_2279,N_2252);
or U2331 (N_2331,N_2227,N_2224);
or U2332 (N_2332,N_2227,N_2279);
nand U2333 (N_2333,N_2265,N_2278);
nor U2334 (N_2334,N_2243,N_2240);
nand U2335 (N_2335,N_2241,N_2227);
and U2336 (N_2336,N_2253,N_2273);
nor U2337 (N_2337,N_2275,N_2224);
and U2338 (N_2338,N_2252,N_2255);
nor U2339 (N_2339,N_2272,N_2235);
nor U2340 (N_2340,N_2282,N_2297);
and U2341 (N_2341,N_2335,N_2288);
and U2342 (N_2342,N_2334,N_2330);
nor U2343 (N_2343,N_2290,N_2294);
nor U2344 (N_2344,N_2283,N_2293);
and U2345 (N_2345,N_2303,N_2326);
or U2346 (N_2346,N_2329,N_2316);
or U2347 (N_2347,N_2289,N_2323);
or U2348 (N_2348,N_2310,N_2305);
nand U2349 (N_2349,N_2299,N_2317);
nand U2350 (N_2350,N_2281,N_2328);
nor U2351 (N_2351,N_2318,N_2322);
or U2352 (N_2352,N_2309,N_2280);
or U2353 (N_2353,N_2319,N_2298);
nand U2354 (N_2354,N_2333,N_2292);
and U2355 (N_2355,N_2307,N_2291);
and U2356 (N_2356,N_2332,N_2325);
nand U2357 (N_2357,N_2337,N_2300);
or U2358 (N_2358,N_2302,N_2285);
nand U2359 (N_2359,N_2313,N_2311);
nand U2360 (N_2360,N_2321,N_2295);
nand U2361 (N_2361,N_2287,N_2312);
or U2362 (N_2362,N_2284,N_2304);
or U2363 (N_2363,N_2331,N_2314);
or U2364 (N_2364,N_2327,N_2296);
nor U2365 (N_2365,N_2315,N_2306);
nand U2366 (N_2366,N_2320,N_2286);
nor U2367 (N_2367,N_2308,N_2301);
or U2368 (N_2368,N_2324,N_2336);
nor U2369 (N_2369,N_2338,N_2339);
nor U2370 (N_2370,N_2339,N_2318);
nor U2371 (N_2371,N_2334,N_2293);
or U2372 (N_2372,N_2302,N_2309);
or U2373 (N_2373,N_2302,N_2326);
nor U2374 (N_2374,N_2295,N_2338);
nor U2375 (N_2375,N_2290,N_2289);
nor U2376 (N_2376,N_2333,N_2329);
or U2377 (N_2377,N_2316,N_2312);
nand U2378 (N_2378,N_2282,N_2294);
or U2379 (N_2379,N_2333,N_2315);
and U2380 (N_2380,N_2316,N_2305);
nand U2381 (N_2381,N_2337,N_2328);
nand U2382 (N_2382,N_2286,N_2291);
or U2383 (N_2383,N_2339,N_2330);
nor U2384 (N_2384,N_2290,N_2328);
and U2385 (N_2385,N_2330,N_2338);
or U2386 (N_2386,N_2300,N_2317);
or U2387 (N_2387,N_2283,N_2314);
and U2388 (N_2388,N_2312,N_2310);
and U2389 (N_2389,N_2286,N_2308);
nor U2390 (N_2390,N_2328,N_2307);
and U2391 (N_2391,N_2317,N_2336);
nand U2392 (N_2392,N_2318,N_2314);
nand U2393 (N_2393,N_2320,N_2329);
nand U2394 (N_2394,N_2309,N_2336);
and U2395 (N_2395,N_2296,N_2293);
and U2396 (N_2396,N_2291,N_2318);
or U2397 (N_2397,N_2314,N_2324);
nor U2398 (N_2398,N_2303,N_2288);
nor U2399 (N_2399,N_2304,N_2295);
and U2400 (N_2400,N_2387,N_2371);
or U2401 (N_2401,N_2363,N_2396);
or U2402 (N_2402,N_2362,N_2345);
or U2403 (N_2403,N_2388,N_2340);
nor U2404 (N_2404,N_2378,N_2357);
nand U2405 (N_2405,N_2398,N_2384);
and U2406 (N_2406,N_2372,N_2350);
or U2407 (N_2407,N_2375,N_2394);
and U2408 (N_2408,N_2379,N_2392);
xor U2409 (N_2409,N_2352,N_2374);
nand U2410 (N_2410,N_2399,N_2397);
and U2411 (N_2411,N_2391,N_2351);
nor U2412 (N_2412,N_2377,N_2359);
nand U2413 (N_2413,N_2358,N_2369);
or U2414 (N_2414,N_2356,N_2361);
or U2415 (N_2415,N_2390,N_2367);
nand U2416 (N_2416,N_2346,N_2385);
or U2417 (N_2417,N_2341,N_2348);
or U2418 (N_2418,N_2347,N_2365);
nor U2419 (N_2419,N_2344,N_2349);
or U2420 (N_2420,N_2380,N_2366);
nor U2421 (N_2421,N_2386,N_2376);
or U2422 (N_2422,N_2382,N_2353);
nand U2423 (N_2423,N_2383,N_2355);
and U2424 (N_2424,N_2373,N_2360);
nand U2425 (N_2425,N_2395,N_2342);
and U2426 (N_2426,N_2364,N_2389);
nor U2427 (N_2427,N_2370,N_2381);
and U2428 (N_2428,N_2393,N_2368);
and U2429 (N_2429,N_2343,N_2354);
and U2430 (N_2430,N_2398,N_2389);
nor U2431 (N_2431,N_2343,N_2386);
nand U2432 (N_2432,N_2388,N_2348);
nor U2433 (N_2433,N_2389,N_2375);
and U2434 (N_2434,N_2397,N_2341);
or U2435 (N_2435,N_2379,N_2356);
nand U2436 (N_2436,N_2363,N_2340);
and U2437 (N_2437,N_2394,N_2355);
nor U2438 (N_2438,N_2368,N_2378);
and U2439 (N_2439,N_2374,N_2346);
and U2440 (N_2440,N_2347,N_2362);
nor U2441 (N_2441,N_2359,N_2357);
nor U2442 (N_2442,N_2399,N_2349);
or U2443 (N_2443,N_2356,N_2372);
or U2444 (N_2444,N_2389,N_2382);
or U2445 (N_2445,N_2366,N_2355);
or U2446 (N_2446,N_2365,N_2370);
nor U2447 (N_2447,N_2365,N_2393);
or U2448 (N_2448,N_2349,N_2345);
or U2449 (N_2449,N_2369,N_2370);
nor U2450 (N_2450,N_2386,N_2395);
nor U2451 (N_2451,N_2364,N_2377);
or U2452 (N_2452,N_2377,N_2383);
nor U2453 (N_2453,N_2397,N_2392);
nor U2454 (N_2454,N_2370,N_2349);
nor U2455 (N_2455,N_2366,N_2373);
and U2456 (N_2456,N_2366,N_2348);
nor U2457 (N_2457,N_2390,N_2348);
and U2458 (N_2458,N_2387,N_2378);
or U2459 (N_2459,N_2386,N_2358);
and U2460 (N_2460,N_2431,N_2404);
nand U2461 (N_2461,N_2440,N_2452);
nor U2462 (N_2462,N_2453,N_2424);
and U2463 (N_2463,N_2443,N_2425);
and U2464 (N_2464,N_2410,N_2450);
and U2465 (N_2465,N_2421,N_2438);
and U2466 (N_2466,N_2407,N_2418);
and U2467 (N_2467,N_2417,N_2448);
or U2468 (N_2468,N_2400,N_2433);
nand U2469 (N_2469,N_2434,N_2456);
and U2470 (N_2470,N_2432,N_2451);
nor U2471 (N_2471,N_2439,N_2457);
nand U2472 (N_2472,N_2416,N_2428);
nor U2473 (N_2473,N_2401,N_2441);
and U2474 (N_2474,N_2411,N_2436);
or U2475 (N_2475,N_2430,N_2402);
or U2476 (N_2476,N_2445,N_2423);
or U2477 (N_2477,N_2427,N_2454);
nor U2478 (N_2478,N_2426,N_2435);
nand U2479 (N_2479,N_2420,N_2442);
or U2480 (N_2480,N_2458,N_2422);
and U2481 (N_2481,N_2405,N_2403);
nor U2482 (N_2482,N_2437,N_2444);
and U2483 (N_2483,N_2447,N_2414);
or U2484 (N_2484,N_2446,N_2455);
or U2485 (N_2485,N_2409,N_2429);
nand U2486 (N_2486,N_2415,N_2408);
or U2487 (N_2487,N_2413,N_2419);
nor U2488 (N_2488,N_2406,N_2412);
and U2489 (N_2489,N_2459,N_2449);
nor U2490 (N_2490,N_2426,N_2403);
or U2491 (N_2491,N_2455,N_2454);
and U2492 (N_2492,N_2446,N_2450);
nor U2493 (N_2493,N_2418,N_2457);
nor U2494 (N_2494,N_2419,N_2440);
and U2495 (N_2495,N_2409,N_2442);
or U2496 (N_2496,N_2400,N_2429);
nand U2497 (N_2497,N_2450,N_2458);
nor U2498 (N_2498,N_2402,N_2405);
and U2499 (N_2499,N_2421,N_2424);
nor U2500 (N_2500,N_2415,N_2450);
nand U2501 (N_2501,N_2444,N_2428);
or U2502 (N_2502,N_2432,N_2459);
nand U2503 (N_2503,N_2454,N_2420);
or U2504 (N_2504,N_2412,N_2454);
or U2505 (N_2505,N_2426,N_2411);
or U2506 (N_2506,N_2432,N_2408);
and U2507 (N_2507,N_2408,N_2414);
or U2508 (N_2508,N_2430,N_2425);
nor U2509 (N_2509,N_2412,N_2427);
nand U2510 (N_2510,N_2455,N_2448);
nor U2511 (N_2511,N_2447,N_2406);
nand U2512 (N_2512,N_2428,N_2453);
or U2513 (N_2513,N_2437,N_2403);
nor U2514 (N_2514,N_2429,N_2445);
or U2515 (N_2515,N_2444,N_2425);
nor U2516 (N_2516,N_2428,N_2458);
and U2517 (N_2517,N_2409,N_2410);
or U2518 (N_2518,N_2415,N_2428);
nor U2519 (N_2519,N_2450,N_2443);
or U2520 (N_2520,N_2476,N_2474);
and U2521 (N_2521,N_2504,N_2497);
nand U2522 (N_2522,N_2493,N_2463);
or U2523 (N_2523,N_2473,N_2488);
and U2524 (N_2524,N_2515,N_2508);
or U2525 (N_2525,N_2491,N_2477);
nand U2526 (N_2526,N_2518,N_2498);
and U2527 (N_2527,N_2490,N_2467);
and U2528 (N_2528,N_2468,N_2489);
nand U2529 (N_2529,N_2469,N_2479);
and U2530 (N_2530,N_2502,N_2487);
nand U2531 (N_2531,N_2475,N_2505);
or U2532 (N_2532,N_2514,N_2460);
nand U2533 (N_2533,N_2470,N_2486);
nand U2534 (N_2534,N_2500,N_2510);
nor U2535 (N_2535,N_2519,N_2503);
and U2536 (N_2536,N_2501,N_2485);
nand U2537 (N_2537,N_2516,N_2480);
nand U2538 (N_2538,N_2512,N_2509);
nor U2539 (N_2539,N_2511,N_2461);
or U2540 (N_2540,N_2462,N_2517);
nand U2541 (N_2541,N_2472,N_2471);
nand U2542 (N_2542,N_2466,N_2483);
nand U2543 (N_2543,N_2513,N_2464);
or U2544 (N_2544,N_2482,N_2481);
and U2545 (N_2545,N_2492,N_2465);
or U2546 (N_2546,N_2494,N_2478);
nand U2547 (N_2547,N_2495,N_2499);
and U2548 (N_2548,N_2496,N_2507);
and U2549 (N_2549,N_2506,N_2484);
nand U2550 (N_2550,N_2498,N_2475);
or U2551 (N_2551,N_2487,N_2512);
and U2552 (N_2552,N_2466,N_2518);
nand U2553 (N_2553,N_2516,N_2484);
nand U2554 (N_2554,N_2478,N_2493);
nand U2555 (N_2555,N_2517,N_2516);
and U2556 (N_2556,N_2473,N_2474);
and U2557 (N_2557,N_2470,N_2495);
and U2558 (N_2558,N_2510,N_2498);
or U2559 (N_2559,N_2500,N_2502);
xor U2560 (N_2560,N_2478,N_2512);
nor U2561 (N_2561,N_2505,N_2462);
nand U2562 (N_2562,N_2489,N_2479);
and U2563 (N_2563,N_2489,N_2470);
nand U2564 (N_2564,N_2464,N_2460);
nand U2565 (N_2565,N_2496,N_2495);
or U2566 (N_2566,N_2467,N_2502);
and U2567 (N_2567,N_2510,N_2512);
and U2568 (N_2568,N_2505,N_2513);
nand U2569 (N_2569,N_2482,N_2475);
nand U2570 (N_2570,N_2502,N_2460);
or U2571 (N_2571,N_2508,N_2461);
nor U2572 (N_2572,N_2484,N_2488);
or U2573 (N_2573,N_2508,N_2472);
or U2574 (N_2574,N_2496,N_2506);
or U2575 (N_2575,N_2490,N_2482);
nor U2576 (N_2576,N_2500,N_2512);
or U2577 (N_2577,N_2465,N_2463);
or U2578 (N_2578,N_2517,N_2472);
nand U2579 (N_2579,N_2493,N_2483);
nor U2580 (N_2580,N_2562,N_2541);
nor U2581 (N_2581,N_2531,N_2524);
nor U2582 (N_2582,N_2573,N_2546);
and U2583 (N_2583,N_2565,N_2578);
and U2584 (N_2584,N_2576,N_2539);
nor U2585 (N_2585,N_2575,N_2533);
nor U2586 (N_2586,N_2556,N_2547);
and U2587 (N_2587,N_2521,N_2523);
or U2588 (N_2588,N_2554,N_2540);
or U2589 (N_2589,N_2526,N_2529);
nor U2590 (N_2590,N_2548,N_2545);
and U2591 (N_2591,N_2553,N_2564);
and U2592 (N_2592,N_2566,N_2555);
or U2593 (N_2593,N_2550,N_2574);
or U2594 (N_2594,N_2528,N_2544);
nand U2595 (N_2595,N_2560,N_2579);
or U2596 (N_2596,N_2535,N_2568);
nor U2597 (N_2597,N_2549,N_2525);
and U2598 (N_2598,N_2561,N_2532);
or U2599 (N_2599,N_2520,N_2537);
nand U2600 (N_2600,N_2551,N_2572);
nand U2601 (N_2601,N_2569,N_2557);
or U2602 (N_2602,N_2534,N_2522);
and U2603 (N_2603,N_2527,N_2570);
or U2604 (N_2604,N_2542,N_2543);
and U2605 (N_2605,N_2571,N_2538);
or U2606 (N_2606,N_2559,N_2530);
nor U2607 (N_2607,N_2558,N_2567);
or U2608 (N_2608,N_2536,N_2563);
or U2609 (N_2609,N_2552,N_2577);
nor U2610 (N_2610,N_2574,N_2526);
and U2611 (N_2611,N_2560,N_2543);
nor U2612 (N_2612,N_2558,N_2534);
nor U2613 (N_2613,N_2530,N_2563);
nor U2614 (N_2614,N_2543,N_2525);
nor U2615 (N_2615,N_2562,N_2549);
nand U2616 (N_2616,N_2553,N_2556);
xor U2617 (N_2617,N_2575,N_2574);
or U2618 (N_2618,N_2522,N_2567);
and U2619 (N_2619,N_2571,N_2572);
xnor U2620 (N_2620,N_2529,N_2574);
nor U2621 (N_2621,N_2536,N_2557);
nor U2622 (N_2622,N_2565,N_2579);
and U2623 (N_2623,N_2568,N_2576);
nand U2624 (N_2624,N_2564,N_2574);
nor U2625 (N_2625,N_2554,N_2534);
nor U2626 (N_2626,N_2521,N_2562);
and U2627 (N_2627,N_2539,N_2532);
nor U2628 (N_2628,N_2573,N_2529);
and U2629 (N_2629,N_2563,N_2553);
or U2630 (N_2630,N_2568,N_2579);
and U2631 (N_2631,N_2521,N_2524);
and U2632 (N_2632,N_2540,N_2526);
and U2633 (N_2633,N_2524,N_2564);
or U2634 (N_2634,N_2531,N_2565);
nor U2635 (N_2635,N_2550,N_2529);
or U2636 (N_2636,N_2527,N_2561);
or U2637 (N_2637,N_2529,N_2542);
and U2638 (N_2638,N_2578,N_2562);
and U2639 (N_2639,N_2533,N_2562);
or U2640 (N_2640,N_2622,N_2591);
nand U2641 (N_2641,N_2618,N_2623);
or U2642 (N_2642,N_2590,N_2611);
nand U2643 (N_2643,N_2620,N_2634);
nor U2644 (N_2644,N_2639,N_2580);
and U2645 (N_2645,N_2596,N_2624);
nand U2646 (N_2646,N_2599,N_2604);
or U2647 (N_2647,N_2621,N_2638);
nand U2648 (N_2648,N_2595,N_2597);
nand U2649 (N_2649,N_2633,N_2628);
or U2650 (N_2650,N_2593,N_2610);
or U2651 (N_2651,N_2601,N_2632);
and U2652 (N_2652,N_2594,N_2619);
and U2653 (N_2653,N_2617,N_2616);
nor U2654 (N_2654,N_2605,N_2609);
nor U2655 (N_2655,N_2581,N_2603);
or U2656 (N_2656,N_2600,N_2584);
nor U2657 (N_2657,N_2582,N_2607);
nor U2658 (N_2658,N_2636,N_2613);
nor U2659 (N_2659,N_2608,N_2614);
nor U2660 (N_2660,N_2606,N_2631);
nand U2661 (N_2661,N_2586,N_2588);
nor U2662 (N_2662,N_2625,N_2637);
nor U2663 (N_2663,N_2629,N_2602);
nor U2664 (N_2664,N_2585,N_2583);
and U2665 (N_2665,N_2612,N_2635);
or U2666 (N_2666,N_2587,N_2630);
nand U2667 (N_2667,N_2627,N_2615);
nand U2668 (N_2668,N_2589,N_2598);
nor U2669 (N_2669,N_2626,N_2592);
or U2670 (N_2670,N_2592,N_2622);
nor U2671 (N_2671,N_2604,N_2637);
nor U2672 (N_2672,N_2628,N_2623);
nor U2673 (N_2673,N_2626,N_2580);
or U2674 (N_2674,N_2590,N_2615);
or U2675 (N_2675,N_2627,N_2618);
nor U2676 (N_2676,N_2614,N_2584);
nor U2677 (N_2677,N_2637,N_2611);
or U2678 (N_2678,N_2580,N_2637);
or U2679 (N_2679,N_2586,N_2589);
nor U2680 (N_2680,N_2594,N_2626);
nor U2681 (N_2681,N_2633,N_2596);
or U2682 (N_2682,N_2620,N_2616);
nor U2683 (N_2683,N_2613,N_2594);
nor U2684 (N_2684,N_2636,N_2584);
nand U2685 (N_2685,N_2613,N_2626);
nand U2686 (N_2686,N_2633,N_2615);
and U2687 (N_2687,N_2584,N_2638);
or U2688 (N_2688,N_2623,N_2616);
and U2689 (N_2689,N_2620,N_2608);
and U2690 (N_2690,N_2638,N_2596);
or U2691 (N_2691,N_2603,N_2582);
and U2692 (N_2692,N_2625,N_2622);
xnor U2693 (N_2693,N_2628,N_2580);
nand U2694 (N_2694,N_2612,N_2606);
or U2695 (N_2695,N_2630,N_2612);
nor U2696 (N_2696,N_2635,N_2610);
nand U2697 (N_2697,N_2615,N_2628);
and U2698 (N_2698,N_2608,N_2631);
nor U2699 (N_2699,N_2587,N_2586);
nor U2700 (N_2700,N_2655,N_2653);
nand U2701 (N_2701,N_2665,N_2661);
nor U2702 (N_2702,N_2687,N_2693);
nand U2703 (N_2703,N_2647,N_2679);
nand U2704 (N_2704,N_2697,N_2684);
or U2705 (N_2705,N_2671,N_2660);
nor U2706 (N_2706,N_2692,N_2678);
nand U2707 (N_2707,N_2644,N_2664);
nor U2708 (N_2708,N_2645,N_2680);
or U2709 (N_2709,N_2667,N_2681);
and U2710 (N_2710,N_2685,N_2650);
nand U2711 (N_2711,N_2683,N_2662);
nor U2712 (N_2712,N_2657,N_2651);
nand U2713 (N_2713,N_2654,N_2646);
or U2714 (N_2714,N_2691,N_2641);
nor U2715 (N_2715,N_2696,N_2670);
or U2716 (N_2716,N_2642,N_2695);
nor U2717 (N_2717,N_2677,N_2676);
nand U2718 (N_2718,N_2698,N_2675);
nor U2719 (N_2719,N_2674,N_2659);
nand U2720 (N_2720,N_2689,N_2666);
nor U2721 (N_2721,N_2672,N_2656);
or U2722 (N_2722,N_2682,N_2643);
nor U2723 (N_2723,N_2658,N_2699);
or U2724 (N_2724,N_2669,N_2649);
or U2725 (N_2725,N_2648,N_2652);
nor U2726 (N_2726,N_2694,N_2640);
nand U2727 (N_2727,N_2663,N_2668);
or U2728 (N_2728,N_2673,N_2690);
and U2729 (N_2729,N_2688,N_2686);
nand U2730 (N_2730,N_2657,N_2687);
nor U2731 (N_2731,N_2674,N_2684);
nand U2732 (N_2732,N_2671,N_2642);
nand U2733 (N_2733,N_2652,N_2641);
nand U2734 (N_2734,N_2681,N_2672);
or U2735 (N_2735,N_2664,N_2672);
and U2736 (N_2736,N_2664,N_2660);
or U2737 (N_2737,N_2671,N_2641);
nand U2738 (N_2738,N_2696,N_2649);
or U2739 (N_2739,N_2669,N_2660);
nor U2740 (N_2740,N_2666,N_2691);
or U2741 (N_2741,N_2682,N_2641);
nand U2742 (N_2742,N_2660,N_2653);
nor U2743 (N_2743,N_2653,N_2688);
and U2744 (N_2744,N_2671,N_2698);
nor U2745 (N_2745,N_2668,N_2658);
nor U2746 (N_2746,N_2647,N_2652);
nand U2747 (N_2747,N_2689,N_2665);
nand U2748 (N_2748,N_2645,N_2650);
nand U2749 (N_2749,N_2644,N_2686);
and U2750 (N_2750,N_2667,N_2650);
or U2751 (N_2751,N_2681,N_2658);
or U2752 (N_2752,N_2641,N_2676);
nor U2753 (N_2753,N_2689,N_2691);
nor U2754 (N_2754,N_2685,N_2690);
and U2755 (N_2755,N_2679,N_2650);
nor U2756 (N_2756,N_2674,N_2645);
and U2757 (N_2757,N_2695,N_2685);
or U2758 (N_2758,N_2694,N_2647);
nand U2759 (N_2759,N_2699,N_2697);
and U2760 (N_2760,N_2724,N_2711);
nor U2761 (N_2761,N_2706,N_2751);
and U2762 (N_2762,N_2739,N_2733);
nor U2763 (N_2763,N_2709,N_2721);
nand U2764 (N_2764,N_2757,N_2703);
or U2765 (N_2765,N_2720,N_2737);
nor U2766 (N_2766,N_2743,N_2748);
nand U2767 (N_2767,N_2745,N_2734);
or U2768 (N_2768,N_2742,N_2723);
nand U2769 (N_2769,N_2747,N_2740);
and U2770 (N_2770,N_2738,N_2730);
and U2771 (N_2771,N_2722,N_2718);
nand U2772 (N_2772,N_2735,N_2758);
or U2773 (N_2773,N_2713,N_2754);
nand U2774 (N_2774,N_2707,N_2705);
and U2775 (N_2775,N_2719,N_2725);
and U2776 (N_2776,N_2746,N_2752);
nor U2777 (N_2777,N_2716,N_2729);
or U2778 (N_2778,N_2755,N_2727);
or U2779 (N_2779,N_2753,N_2714);
xnor U2780 (N_2780,N_2732,N_2708);
nor U2781 (N_2781,N_2726,N_2744);
nor U2782 (N_2782,N_2717,N_2728);
or U2783 (N_2783,N_2702,N_2701);
or U2784 (N_2784,N_2700,N_2715);
and U2785 (N_2785,N_2741,N_2736);
nor U2786 (N_2786,N_2750,N_2731);
nor U2787 (N_2787,N_2712,N_2759);
and U2788 (N_2788,N_2704,N_2749);
or U2789 (N_2789,N_2710,N_2756);
or U2790 (N_2790,N_2723,N_2744);
and U2791 (N_2791,N_2710,N_2722);
nand U2792 (N_2792,N_2756,N_2755);
nand U2793 (N_2793,N_2759,N_2745);
or U2794 (N_2794,N_2754,N_2733);
and U2795 (N_2795,N_2728,N_2741);
nor U2796 (N_2796,N_2717,N_2709);
and U2797 (N_2797,N_2739,N_2702);
nor U2798 (N_2798,N_2701,N_2749);
nand U2799 (N_2799,N_2707,N_2708);
nor U2800 (N_2800,N_2712,N_2739);
and U2801 (N_2801,N_2730,N_2715);
nor U2802 (N_2802,N_2744,N_2714);
and U2803 (N_2803,N_2728,N_2731);
or U2804 (N_2804,N_2736,N_2745);
or U2805 (N_2805,N_2749,N_2719);
and U2806 (N_2806,N_2758,N_2733);
nor U2807 (N_2807,N_2734,N_2716);
nand U2808 (N_2808,N_2745,N_2751);
or U2809 (N_2809,N_2753,N_2719);
nand U2810 (N_2810,N_2725,N_2716);
nand U2811 (N_2811,N_2739,N_2722);
and U2812 (N_2812,N_2754,N_2719);
nor U2813 (N_2813,N_2708,N_2709);
or U2814 (N_2814,N_2739,N_2730);
or U2815 (N_2815,N_2720,N_2716);
and U2816 (N_2816,N_2750,N_2733);
and U2817 (N_2817,N_2714,N_2720);
or U2818 (N_2818,N_2758,N_2715);
or U2819 (N_2819,N_2746,N_2714);
nand U2820 (N_2820,N_2768,N_2779);
and U2821 (N_2821,N_2787,N_2780);
nor U2822 (N_2822,N_2814,N_2816);
nand U2823 (N_2823,N_2806,N_2774);
and U2824 (N_2824,N_2810,N_2804);
or U2825 (N_2825,N_2772,N_2778);
nor U2826 (N_2826,N_2762,N_2790);
and U2827 (N_2827,N_2770,N_2782);
and U2828 (N_2828,N_2792,N_2785);
and U2829 (N_2829,N_2781,N_2776);
nand U2830 (N_2830,N_2801,N_2773);
and U2831 (N_2831,N_2805,N_2818);
and U2832 (N_2832,N_2794,N_2811);
nor U2833 (N_2833,N_2784,N_2775);
nor U2834 (N_2834,N_2797,N_2767);
xnor U2835 (N_2835,N_2789,N_2764);
nand U2836 (N_2836,N_2793,N_2766);
nand U2837 (N_2837,N_2783,N_2788);
xor U2838 (N_2838,N_2761,N_2760);
nor U2839 (N_2839,N_2813,N_2777);
nand U2840 (N_2840,N_2796,N_2807);
or U2841 (N_2841,N_2798,N_2799);
nor U2842 (N_2842,N_2795,N_2769);
nand U2843 (N_2843,N_2771,N_2809);
and U2844 (N_2844,N_2819,N_2803);
nand U2845 (N_2845,N_2791,N_2817);
nand U2846 (N_2846,N_2800,N_2786);
nand U2847 (N_2847,N_2802,N_2808);
nand U2848 (N_2848,N_2812,N_2765);
and U2849 (N_2849,N_2763,N_2815);
or U2850 (N_2850,N_2813,N_2810);
nor U2851 (N_2851,N_2774,N_2799);
or U2852 (N_2852,N_2803,N_2791);
or U2853 (N_2853,N_2771,N_2766);
or U2854 (N_2854,N_2790,N_2788);
nand U2855 (N_2855,N_2779,N_2801);
or U2856 (N_2856,N_2791,N_2766);
nor U2857 (N_2857,N_2772,N_2807);
and U2858 (N_2858,N_2813,N_2761);
nor U2859 (N_2859,N_2789,N_2781);
or U2860 (N_2860,N_2799,N_2777);
or U2861 (N_2861,N_2787,N_2778);
nor U2862 (N_2862,N_2819,N_2801);
nand U2863 (N_2863,N_2766,N_2806);
and U2864 (N_2864,N_2770,N_2761);
or U2865 (N_2865,N_2780,N_2801);
nor U2866 (N_2866,N_2801,N_2777);
nor U2867 (N_2867,N_2764,N_2781);
or U2868 (N_2868,N_2768,N_2783);
or U2869 (N_2869,N_2803,N_2797);
nand U2870 (N_2870,N_2799,N_2787);
nor U2871 (N_2871,N_2791,N_2800);
nor U2872 (N_2872,N_2817,N_2811);
xnor U2873 (N_2873,N_2775,N_2760);
nand U2874 (N_2874,N_2769,N_2774);
nand U2875 (N_2875,N_2814,N_2795);
and U2876 (N_2876,N_2762,N_2805);
and U2877 (N_2877,N_2794,N_2760);
nand U2878 (N_2878,N_2810,N_2782);
or U2879 (N_2879,N_2760,N_2819);
nand U2880 (N_2880,N_2842,N_2822);
nand U2881 (N_2881,N_2826,N_2873);
or U2882 (N_2882,N_2868,N_2829);
or U2883 (N_2883,N_2851,N_2847);
nand U2884 (N_2884,N_2841,N_2866);
nor U2885 (N_2885,N_2855,N_2840);
and U2886 (N_2886,N_2850,N_2875);
or U2887 (N_2887,N_2835,N_2863);
nand U2888 (N_2888,N_2838,N_2845);
or U2889 (N_2889,N_2879,N_2867);
or U2890 (N_2890,N_2830,N_2849);
or U2891 (N_2891,N_2827,N_2869);
nand U2892 (N_2892,N_2846,N_2859);
or U2893 (N_2893,N_2854,N_2872);
or U2894 (N_2894,N_2862,N_2848);
nand U2895 (N_2895,N_2831,N_2833);
or U2896 (N_2896,N_2857,N_2824);
xor U2897 (N_2897,N_2820,N_2844);
and U2898 (N_2898,N_2837,N_2839);
nor U2899 (N_2899,N_2874,N_2832);
nor U2900 (N_2900,N_2825,N_2821);
and U2901 (N_2901,N_2834,N_2856);
or U2902 (N_2902,N_2860,N_2828);
nor U2903 (N_2903,N_2877,N_2864);
nor U2904 (N_2904,N_2861,N_2853);
nor U2905 (N_2905,N_2858,N_2852);
nand U2906 (N_2906,N_2865,N_2843);
nand U2907 (N_2907,N_2823,N_2876);
nor U2908 (N_2908,N_2871,N_2870);
or U2909 (N_2909,N_2878,N_2836);
or U2910 (N_2910,N_2858,N_2832);
nand U2911 (N_2911,N_2870,N_2860);
nand U2912 (N_2912,N_2872,N_2831);
or U2913 (N_2913,N_2877,N_2857);
or U2914 (N_2914,N_2875,N_2840);
nor U2915 (N_2915,N_2826,N_2833);
nor U2916 (N_2916,N_2862,N_2869);
nor U2917 (N_2917,N_2833,N_2846);
and U2918 (N_2918,N_2858,N_2874);
or U2919 (N_2919,N_2830,N_2851);
nand U2920 (N_2920,N_2850,N_2844);
or U2921 (N_2921,N_2863,N_2866);
and U2922 (N_2922,N_2834,N_2877);
or U2923 (N_2923,N_2836,N_2830);
or U2924 (N_2924,N_2821,N_2837);
or U2925 (N_2925,N_2831,N_2850);
or U2926 (N_2926,N_2822,N_2865);
nand U2927 (N_2927,N_2862,N_2849);
and U2928 (N_2928,N_2871,N_2863);
and U2929 (N_2929,N_2873,N_2877);
and U2930 (N_2930,N_2822,N_2872);
and U2931 (N_2931,N_2862,N_2874);
and U2932 (N_2932,N_2873,N_2874);
and U2933 (N_2933,N_2828,N_2870);
nand U2934 (N_2934,N_2869,N_2867);
nand U2935 (N_2935,N_2867,N_2831);
nand U2936 (N_2936,N_2864,N_2837);
nor U2937 (N_2937,N_2840,N_2876);
nand U2938 (N_2938,N_2840,N_2859);
nor U2939 (N_2939,N_2846,N_2822);
nand U2940 (N_2940,N_2901,N_2924);
nor U2941 (N_2941,N_2923,N_2910);
or U2942 (N_2942,N_2906,N_2926);
and U2943 (N_2943,N_2919,N_2920);
or U2944 (N_2944,N_2897,N_2937);
or U2945 (N_2945,N_2914,N_2928);
or U2946 (N_2946,N_2895,N_2882);
nand U2947 (N_2947,N_2903,N_2905);
nand U2948 (N_2948,N_2908,N_2915);
nor U2949 (N_2949,N_2916,N_2934);
and U2950 (N_2950,N_2912,N_2939);
nor U2951 (N_2951,N_2917,N_2913);
nor U2952 (N_2952,N_2891,N_2911);
or U2953 (N_2953,N_2931,N_2929);
nand U2954 (N_2954,N_2922,N_2907);
nand U2955 (N_2955,N_2899,N_2927);
nand U2956 (N_2956,N_2887,N_2884);
or U2957 (N_2957,N_2909,N_2936);
and U2958 (N_2958,N_2900,N_2935);
nand U2959 (N_2959,N_2896,N_2894);
and U2960 (N_2960,N_2890,N_2930);
and U2961 (N_2961,N_2925,N_2933);
and U2962 (N_2962,N_2886,N_2893);
nand U2963 (N_2963,N_2938,N_2932);
or U2964 (N_2964,N_2888,N_2885);
nor U2965 (N_2965,N_2902,N_2889);
nor U2966 (N_2966,N_2881,N_2883);
nor U2967 (N_2967,N_2921,N_2880);
or U2968 (N_2968,N_2898,N_2892);
nand U2969 (N_2969,N_2904,N_2918);
and U2970 (N_2970,N_2901,N_2906);
nor U2971 (N_2971,N_2918,N_2936);
nor U2972 (N_2972,N_2936,N_2923);
nand U2973 (N_2973,N_2884,N_2906);
nor U2974 (N_2974,N_2928,N_2898);
or U2975 (N_2975,N_2904,N_2910);
xor U2976 (N_2976,N_2880,N_2926);
or U2977 (N_2977,N_2918,N_2937);
nand U2978 (N_2978,N_2930,N_2901);
nand U2979 (N_2979,N_2917,N_2889);
and U2980 (N_2980,N_2897,N_2923);
or U2981 (N_2981,N_2928,N_2909);
nand U2982 (N_2982,N_2910,N_2888);
nor U2983 (N_2983,N_2885,N_2915);
and U2984 (N_2984,N_2926,N_2931);
nor U2985 (N_2985,N_2934,N_2892);
or U2986 (N_2986,N_2896,N_2923);
nor U2987 (N_2987,N_2915,N_2883);
nor U2988 (N_2988,N_2896,N_2911);
and U2989 (N_2989,N_2924,N_2890);
nor U2990 (N_2990,N_2888,N_2925);
or U2991 (N_2991,N_2937,N_2926);
or U2992 (N_2992,N_2892,N_2935);
nand U2993 (N_2993,N_2882,N_2908);
or U2994 (N_2994,N_2903,N_2927);
and U2995 (N_2995,N_2898,N_2933);
nor U2996 (N_2996,N_2931,N_2934);
and U2997 (N_2997,N_2937,N_2932);
and U2998 (N_2998,N_2888,N_2919);
nand U2999 (N_2999,N_2919,N_2890);
and UO_0 (O_0,N_2976,N_2997);
nor UO_1 (O_1,N_2949,N_2973);
nor UO_2 (O_2,N_2967,N_2946);
nand UO_3 (O_3,N_2952,N_2972);
nand UO_4 (O_4,N_2991,N_2969);
or UO_5 (O_5,N_2958,N_2960);
and UO_6 (O_6,N_2945,N_2951);
and UO_7 (O_7,N_2962,N_2995);
nor UO_8 (O_8,N_2943,N_2983);
and UO_9 (O_9,N_2959,N_2974);
and UO_10 (O_10,N_2975,N_2941);
nor UO_11 (O_11,N_2986,N_2992);
and UO_12 (O_12,N_2982,N_2940);
nand UO_13 (O_13,N_2977,N_2947);
or UO_14 (O_14,N_2954,N_2979);
and UO_15 (O_15,N_2956,N_2948);
or UO_16 (O_16,N_2963,N_2953);
or UO_17 (O_17,N_2980,N_2993);
and UO_18 (O_18,N_2970,N_2981);
nand UO_19 (O_19,N_2957,N_2944);
or UO_20 (O_20,N_2988,N_2990);
and UO_21 (O_21,N_2994,N_2968);
or UO_22 (O_22,N_2942,N_2961);
and UO_23 (O_23,N_2964,N_2965);
nand UO_24 (O_24,N_2966,N_2955);
nand UO_25 (O_25,N_2989,N_2978);
nand UO_26 (O_26,N_2971,N_2987);
nand UO_27 (O_27,N_2996,N_2984);
nand UO_28 (O_28,N_2999,N_2985);
nand UO_29 (O_29,N_2998,N_2950);
nor UO_30 (O_30,N_2974,N_2944);
or UO_31 (O_31,N_2979,N_2955);
nor UO_32 (O_32,N_2992,N_2982);
nand UO_33 (O_33,N_2974,N_2988);
nand UO_34 (O_34,N_2943,N_2963);
nor UO_35 (O_35,N_2972,N_2950);
and UO_36 (O_36,N_2993,N_2978);
nor UO_37 (O_37,N_2977,N_2950);
and UO_38 (O_38,N_2956,N_2961);
nand UO_39 (O_39,N_2974,N_2983);
nor UO_40 (O_40,N_2967,N_2957);
nor UO_41 (O_41,N_2941,N_2962);
nand UO_42 (O_42,N_2949,N_2965);
or UO_43 (O_43,N_2988,N_2944);
and UO_44 (O_44,N_2957,N_2945);
or UO_45 (O_45,N_2960,N_2984);
nor UO_46 (O_46,N_2974,N_2977);
nor UO_47 (O_47,N_2963,N_2990);
nand UO_48 (O_48,N_2967,N_2974);
nand UO_49 (O_49,N_2949,N_2972);
nor UO_50 (O_50,N_2975,N_2979);
or UO_51 (O_51,N_2983,N_2990);
and UO_52 (O_52,N_2974,N_2960);
nor UO_53 (O_53,N_2954,N_2983);
nor UO_54 (O_54,N_2966,N_2940);
nor UO_55 (O_55,N_2981,N_2969);
nand UO_56 (O_56,N_2969,N_2943);
nand UO_57 (O_57,N_2941,N_2987);
or UO_58 (O_58,N_2969,N_2959);
nand UO_59 (O_59,N_2964,N_2959);
nor UO_60 (O_60,N_2991,N_2976);
and UO_61 (O_61,N_2986,N_2946);
nand UO_62 (O_62,N_2984,N_2949);
nand UO_63 (O_63,N_2979,N_2965);
nor UO_64 (O_64,N_2979,N_2984);
and UO_65 (O_65,N_2993,N_2989);
nor UO_66 (O_66,N_2948,N_2991);
or UO_67 (O_67,N_2975,N_2968);
nor UO_68 (O_68,N_2986,N_2948);
nor UO_69 (O_69,N_2945,N_2985);
and UO_70 (O_70,N_2996,N_2946);
or UO_71 (O_71,N_2966,N_2968);
nand UO_72 (O_72,N_2989,N_2992);
nand UO_73 (O_73,N_2996,N_2964);
nand UO_74 (O_74,N_2964,N_2972);
or UO_75 (O_75,N_2958,N_2969);
nand UO_76 (O_76,N_2988,N_2972);
or UO_77 (O_77,N_2974,N_2963);
nor UO_78 (O_78,N_2965,N_2974);
or UO_79 (O_79,N_2997,N_2989);
nand UO_80 (O_80,N_2943,N_2940);
and UO_81 (O_81,N_2979,N_2977);
or UO_82 (O_82,N_2968,N_2991);
or UO_83 (O_83,N_2995,N_2988);
or UO_84 (O_84,N_2947,N_2970);
nand UO_85 (O_85,N_2966,N_2992);
nor UO_86 (O_86,N_2981,N_2954);
nor UO_87 (O_87,N_2954,N_2949);
or UO_88 (O_88,N_2982,N_2973);
or UO_89 (O_89,N_2966,N_2976);
or UO_90 (O_90,N_2971,N_2995);
nor UO_91 (O_91,N_2979,N_2952);
nor UO_92 (O_92,N_2999,N_2998);
or UO_93 (O_93,N_2954,N_2959);
or UO_94 (O_94,N_2955,N_2990);
nand UO_95 (O_95,N_2980,N_2950);
nand UO_96 (O_96,N_2972,N_2995);
and UO_97 (O_97,N_2984,N_2957);
nand UO_98 (O_98,N_2980,N_2996);
or UO_99 (O_99,N_2979,N_2963);
or UO_100 (O_100,N_2966,N_2958);
nand UO_101 (O_101,N_2948,N_2947);
or UO_102 (O_102,N_2944,N_2993);
or UO_103 (O_103,N_2950,N_2947);
nand UO_104 (O_104,N_2957,N_2954);
nor UO_105 (O_105,N_2966,N_2951);
nor UO_106 (O_106,N_2963,N_2965);
nor UO_107 (O_107,N_2961,N_2978);
or UO_108 (O_108,N_2981,N_2989);
nand UO_109 (O_109,N_2958,N_2992);
or UO_110 (O_110,N_2988,N_2986);
and UO_111 (O_111,N_2992,N_2996);
and UO_112 (O_112,N_2948,N_2943);
and UO_113 (O_113,N_2967,N_2992);
or UO_114 (O_114,N_2946,N_2984);
nor UO_115 (O_115,N_2943,N_2991);
and UO_116 (O_116,N_2980,N_2942);
nor UO_117 (O_117,N_2940,N_2962);
or UO_118 (O_118,N_2985,N_2950);
and UO_119 (O_119,N_2994,N_2942);
and UO_120 (O_120,N_2975,N_2967);
nor UO_121 (O_121,N_2983,N_2971);
nor UO_122 (O_122,N_2959,N_2999);
nor UO_123 (O_123,N_2962,N_2994);
or UO_124 (O_124,N_2943,N_2971);
and UO_125 (O_125,N_2944,N_2975);
nand UO_126 (O_126,N_2960,N_2990);
nand UO_127 (O_127,N_2968,N_2981);
and UO_128 (O_128,N_2955,N_2959);
or UO_129 (O_129,N_2979,N_2993);
or UO_130 (O_130,N_2996,N_2955);
and UO_131 (O_131,N_2965,N_2992);
nor UO_132 (O_132,N_2955,N_2946);
nand UO_133 (O_133,N_2995,N_2989);
and UO_134 (O_134,N_2980,N_2961);
nor UO_135 (O_135,N_2979,N_2969);
or UO_136 (O_136,N_2993,N_2962);
nand UO_137 (O_137,N_2958,N_2997);
or UO_138 (O_138,N_2985,N_2990);
and UO_139 (O_139,N_2954,N_2962);
or UO_140 (O_140,N_2986,N_2972);
and UO_141 (O_141,N_2992,N_2970);
and UO_142 (O_142,N_2947,N_2958);
or UO_143 (O_143,N_2999,N_2955);
or UO_144 (O_144,N_2991,N_2996);
or UO_145 (O_145,N_2953,N_2959);
and UO_146 (O_146,N_2972,N_2943);
and UO_147 (O_147,N_2950,N_2941);
nand UO_148 (O_148,N_2968,N_2946);
and UO_149 (O_149,N_2947,N_2952);
and UO_150 (O_150,N_2986,N_2987);
or UO_151 (O_151,N_2944,N_2947);
or UO_152 (O_152,N_2990,N_2969);
and UO_153 (O_153,N_2988,N_2978);
nand UO_154 (O_154,N_2941,N_2991);
and UO_155 (O_155,N_2966,N_2978);
nor UO_156 (O_156,N_2966,N_2948);
and UO_157 (O_157,N_2987,N_2990);
nor UO_158 (O_158,N_2951,N_2971);
or UO_159 (O_159,N_2943,N_2982);
and UO_160 (O_160,N_2988,N_2960);
nor UO_161 (O_161,N_2992,N_2963);
nand UO_162 (O_162,N_2976,N_2951);
nand UO_163 (O_163,N_2977,N_2983);
nand UO_164 (O_164,N_2958,N_2980);
nand UO_165 (O_165,N_2988,N_2971);
or UO_166 (O_166,N_2976,N_2940);
nand UO_167 (O_167,N_2990,N_2993);
or UO_168 (O_168,N_2994,N_2995);
or UO_169 (O_169,N_2987,N_2964);
nor UO_170 (O_170,N_2990,N_2950);
and UO_171 (O_171,N_2961,N_2949);
nor UO_172 (O_172,N_2953,N_2994);
nor UO_173 (O_173,N_2983,N_2967);
and UO_174 (O_174,N_2943,N_2976);
and UO_175 (O_175,N_2963,N_2949);
or UO_176 (O_176,N_2987,N_2951);
nand UO_177 (O_177,N_2992,N_2997);
and UO_178 (O_178,N_2981,N_2945);
nand UO_179 (O_179,N_2974,N_2976);
and UO_180 (O_180,N_2960,N_2999);
nor UO_181 (O_181,N_2979,N_2992);
and UO_182 (O_182,N_2976,N_2975);
nor UO_183 (O_183,N_2992,N_2947);
nor UO_184 (O_184,N_2967,N_2945);
and UO_185 (O_185,N_2965,N_2968);
nand UO_186 (O_186,N_2943,N_2966);
nand UO_187 (O_187,N_2968,N_2997);
and UO_188 (O_188,N_2974,N_2940);
or UO_189 (O_189,N_2982,N_2998);
and UO_190 (O_190,N_2974,N_2998);
nand UO_191 (O_191,N_2960,N_2993);
or UO_192 (O_192,N_2948,N_2960);
nor UO_193 (O_193,N_2961,N_2983);
and UO_194 (O_194,N_2981,N_2966);
or UO_195 (O_195,N_2987,N_2968);
and UO_196 (O_196,N_2985,N_2988);
and UO_197 (O_197,N_2941,N_2942);
nor UO_198 (O_198,N_2951,N_2943);
nor UO_199 (O_199,N_2949,N_2942);
and UO_200 (O_200,N_2959,N_2967);
nor UO_201 (O_201,N_2962,N_2982);
and UO_202 (O_202,N_2950,N_2993);
or UO_203 (O_203,N_2958,N_2948);
or UO_204 (O_204,N_2984,N_2971);
nor UO_205 (O_205,N_2977,N_2998);
nor UO_206 (O_206,N_2981,N_2973);
nand UO_207 (O_207,N_2962,N_2956);
nand UO_208 (O_208,N_2952,N_2946);
nor UO_209 (O_209,N_2978,N_2940);
nand UO_210 (O_210,N_2976,N_2979);
or UO_211 (O_211,N_2946,N_2956);
nor UO_212 (O_212,N_2942,N_2967);
and UO_213 (O_213,N_2970,N_2961);
nor UO_214 (O_214,N_2942,N_2987);
and UO_215 (O_215,N_2981,N_2983);
and UO_216 (O_216,N_2989,N_2971);
and UO_217 (O_217,N_2977,N_2952);
nand UO_218 (O_218,N_2953,N_2986);
and UO_219 (O_219,N_2971,N_2967);
or UO_220 (O_220,N_2982,N_2946);
and UO_221 (O_221,N_2964,N_2956);
nand UO_222 (O_222,N_2943,N_2984);
or UO_223 (O_223,N_2974,N_2948);
nand UO_224 (O_224,N_2956,N_2995);
or UO_225 (O_225,N_2968,N_2954);
and UO_226 (O_226,N_2996,N_2986);
xnor UO_227 (O_227,N_2984,N_2976);
nor UO_228 (O_228,N_2972,N_2970);
nand UO_229 (O_229,N_2949,N_2993);
or UO_230 (O_230,N_2993,N_2955);
and UO_231 (O_231,N_2973,N_2968);
or UO_232 (O_232,N_2942,N_2977);
or UO_233 (O_233,N_2976,N_2986);
and UO_234 (O_234,N_2973,N_2966);
nor UO_235 (O_235,N_2953,N_2972);
nor UO_236 (O_236,N_2997,N_2981);
and UO_237 (O_237,N_2967,N_2962);
nor UO_238 (O_238,N_2984,N_2987);
nor UO_239 (O_239,N_2973,N_2948);
or UO_240 (O_240,N_2998,N_2948);
nor UO_241 (O_241,N_2973,N_2977);
nor UO_242 (O_242,N_2957,N_2960);
nand UO_243 (O_243,N_2959,N_2972);
nand UO_244 (O_244,N_2969,N_2998);
and UO_245 (O_245,N_2973,N_2944);
or UO_246 (O_246,N_2972,N_2981);
nand UO_247 (O_247,N_2973,N_2945);
and UO_248 (O_248,N_2944,N_2940);
nor UO_249 (O_249,N_2943,N_2946);
and UO_250 (O_250,N_2966,N_2967);
nand UO_251 (O_251,N_2974,N_2942);
nand UO_252 (O_252,N_2994,N_2963);
or UO_253 (O_253,N_2942,N_2986);
nor UO_254 (O_254,N_2955,N_2968);
nand UO_255 (O_255,N_2979,N_2974);
or UO_256 (O_256,N_2999,N_2958);
nor UO_257 (O_257,N_2966,N_2971);
nor UO_258 (O_258,N_2964,N_2994);
or UO_259 (O_259,N_2989,N_2986);
nand UO_260 (O_260,N_2943,N_2987);
and UO_261 (O_261,N_2965,N_2946);
nand UO_262 (O_262,N_2969,N_2978);
nor UO_263 (O_263,N_2974,N_2945);
or UO_264 (O_264,N_2940,N_2994);
nor UO_265 (O_265,N_2991,N_2988);
nor UO_266 (O_266,N_2963,N_2946);
or UO_267 (O_267,N_2991,N_2989);
or UO_268 (O_268,N_2982,N_2957);
nand UO_269 (O_269,N_2962,N_2984);
or UO_270 (O_270,N_2951,N_2980);
or UO_271 (O_271,N_2951,N_2950);
nor UO_272 (O_272,N_2968,N_2940);
nor UO_273 (O_273,N_2976,N_2983);
or UO_274 (O_274,N_2960,N_2940);
nand UO_275 (O_275,N_2987,N_2958);
nor UO_276 (O_276,N_2965,N_2975);
nor UO_277 (O_277,N_2970,N_2950);
and UO_278 (O_278,N_2950,N_2940);
xor UO_279 (O_279,N_2988,N_2984);
and UO_280 (O_280,N_2985,N_2978);
or UO_281 (O_281,N_2957,N_2981);
or UO_282 (O_282,N_2985,N_2998);
or UO_283 (O_283,N_2963,N_2940);
nand UO_284 (O_284,N_2946,N_2973);
and UO_285 (O_285,N_2942,N_2978);
nand UO_286 (O_286,N_2943,N_2994);
and UO_287 (O_287,N_2984,N_2982);
or UO_288 (O_288,N_2998,N_2952);
and UO_289 (O_289,N_2995,N_2966);
and UO_290 (O_290,N_2968,N_2976);
nor UO_291 (O_291,N_2940,N_2980);
nand UO_292 (O_292,N_2981,N_2977);
and UO_293 (O_293,N_2981,N_2993);
nand UO_294 (O_294,N_2981,N_2991);
and UO_295 (O_295,N_2975,N_2961);
and UO_296 (O_296,N_2991,N_2955);
or UO_297 (O_297,N_2967,N_2985);
or UO_298 (O_298,N_2956,N_2980);
nor UO_299 (O_299,N_2947,N_2960);
or UO_300 (O_300,N_2979,N_2981);
nor UO_301 (O_301,N_2973,N_2994);
nand UO_302 (O_302,N_2984,N_2995);
nor UO_303 (O_303,N_2994,N_2956);
nor UO_304 (O_304,N_2982,N_2945);
and UO_305 (O_305,N_2998,N_2992);
or UO_306 (O_306,N_2962,N_2998);
nand UO_307 (O_307,N_2967,N_2940);
and UO_308 (O_308,N_2950,N_2967);
or UO_309 (O_309,N_2950,N_2996);
or UO_310 (O_310,N_2944,N_2945);
and UO_311 (O_311,N_2948,N_2955);
nand UO_312 (O_312,N_2959,N_2996);
nor UO_313 (O_313,N_2989,N_2976);
nand UO_314 (O_314,N_2941,N_2990);
nand UO_315 (O_315,N_2982,N_2990);
nor UO_316 (O_316,N_2989,N_2984);
nand UO_317 (O_317,N_2964,N_2941);
nor UO_318 (O_318,N_2980,N_2946);
and UO_319 (O_319,N_2953,N_2942);
nand UO_320 (O_320,N_2973,N_2999);
nand UO_321 (O_321,N_2945,N_2965);
and UO_322 (O_322,N_2970,N_2995);
and UO_323 (O_323,N_2999,N_2995);
and UO_324 (O_324,N_2967,N_2989);
nor UO_325 (O_325,N_2991,N_2971);
xor UO_326 (O_326,N_2999,N_2953);
nor UO_327 (O_327,N_2986,N_2961);
or UO_328 (O_328,N_2957,N_2986);
nand UO_329 (O_329,N_2979,N_2960);
and UO_330 (O_330,N_2956,N_2952);
and UO_331 (O_331,N_2970,N_2999);
and UO_332 (O_332,N_2959,N_2982);
nand UO_333 (O_333,N_2987,N_2944);
and UO_334 (O_334,N_2997,N_2994);
and UO_335 (O_335,N_2968,N_2967);
xor UO_336 (O_336,N_2947,N_2969);
and UO_337 (O_337,N_2961,N_2952);
and UO_338 (O_338,N_2984,N_2985);
and UO_339 (O_339,N_2968,N_2947);
nand UO_340 (O_340,N_2940,N_2941);
nand UO_341 (O_341,N_2998,N_2994);
nand UO_342 (O_342,N_2946,N_2957);
nor UO_343 (O_343,N_2971,N_2985);
nand UO_344 (O_344,N_2998,N_2966);
and UO_345 (O_345,N_2949,N_2974);
nor UO_346 (O_346,N_2956,N_2990);
or UO_347 (O_347,N_2980,N_2952);
and UO_348 (O_348,N_2959,N_2976);
and UO_349 (O_349,N_2974,N_2994);
and UO_350 (O_350,N_2972,N_2996);
or UO_351 (O_351,N_2944,N_2946);
nand UO_352 (O_352,N_2946,N_2981);
nand UO_353 (O_353,N_2973,N_2983);
and UO_354 (O_354,N_2994,N_2959);
nor UO_355 (O_355,N_2949,N_2983);
or UO_356 (O_356,N_2940,N_2952);
and UO_357 (O_357,N_2974,N_2955);
or UO_358 (O_358,N_2989,N_2982);
nor UO_359 (O_359,N_2951,N_2994);
and UO_360 (O_360,N_2968,N_2996);
nand UO_361 (O_361,N_2993,N_2999);
and UO_362 (O_362,N_2978,N_2994);
or UO_363 (O_363,N_2984,N_2958);
nor UO_364 (O_364,N_2990,N_2972);
nand UO_365 (O_365,N_2948,N_2968);
or UO_366 (O_366,N_2953,N_2956);
or UO_367 (O_367,N_2941,N_2999);
or UO_368 (O_368,N_2984,N_2941);
nand UO_369 (O_369,N_2976,N_2960);
nor UO_370 (O_370,N_2992,N_2977);
or UO_371 (O_371,N_2995,N_2947);
nand UO_372 (O_372,N_2961,N_2996);
or UO_373 (O_373,N_2950,N_2982);
and UO_374 (O_374,N_2991,N_2966);
or UO_375 (O_375,N_2992,N_2941);
and UO_376 (O_376,N_2941,N_2954);
or UO_377 (O_377,N_2991,N_2975);
and UO_378 (O_378,N_2985,N_2974);
nand UO_379 (O_379,N_2995,N_2944);
nand UO_380 (O_380,N_2980,N_2948);
nor UO_381 (O_381,N_2952,N_2985);
nand UO_382 (O_382,N_2999,N_2987);
and UO_383 (O_383,N_2995,N_2961);
nand UO_384 (O_384,N_2999,N_2986);
or UO_385 (O_385,N_2963,N_2981);
nor UO_386 (O_386,N_2992,N_2984);
nor UO_387 (O_387,N_2970,N_2979);
and UO_388 (O_388,N_2941,N_2963);
and UO_389 (O_389,N_2942,N_2993);
nand UO_390 (O_390,N_2941,N_2957);
nand UO_391 (O_391,N_2990,N_2943);
nand UO_392 (O_392,N_2974,N_2992);
xnor UO_393 (O_393,N_2966,N_2945);
nor UO_394 (O_394,N_2957,N_2989);
and UO_395 (O_395,N_2957,N_2961);
or UO_396 (O_396,N_2959,N_2985);
nor UO_397 (O_397,N_2969,N_2963);
and UO_398 (O_398,N_2945,N_2964);
nand UO_399 (O_399,N_2969,N_2980);
nor UO_400 (O_400,N_2983,N_2962);
or UO_401 (O_401,N_2964,N_2992);
nand UO_402 (O_402,N_2979,N_2968);
or UO_403 (O_403,N_2960,N_2949);
and UO_404 (O_404,N_2992,N_2961);
nor UO_405 (O_405,N_2997,N_2988);
or UO_406 (O_406,N_2970,N_2975);
nor UO_407 (O_407,N_2948,N_2940);
nand UO_408 (O_408,N_2994,N_2949);
or UO_409 (O_409,N_2941,N_2949);
or UO_410 (O_410,N_2955,N_2992);
and UO_411 (O_411,N_2959,N_2948);
nand UO_412 (O_412,N_2945,N_2991);
nor UO_413 (O_413,N_2985,N_2961);
nand UO_414 (O_414,N_2989,N_2952);
nor UO_415 (O_415,N_2969,N_2973);
nor UO_416 (O_416,N_2969,N_2946);
nand UO_417 (O_417,N_2967,N_2977);
nand UO_418 (O_418,N_2957,N_2953);
nand UO_419 (O_419,N_2976,N_2973);
nand UO_420 (O_420,N_2958,N_2989);
and UO_421 (O_421,N_2947,N_2979);
nand UO_422 (O_422,N_2979,N_2966);
and UO_423 (O_423,N_2964,N_2943);
nor UO_424 (O_424,N_2996,N_2985);
nand UO_425 (O_425,N_2978,N_2996);
nand UO_426 (O_426,N_2996,N_2958);
or UO_427 (O_427,N_2974,N_2943);
nand UO_428 (O_428,N_2961,N_2998);
nand UO_429 (O_429,N_2962,N_2969);
or UO_430 (O_430,N_2978,N_2957);
nor UO_431 (O_431,N_2994,N_2941);
nor UO_432 (O_432,N_2998,N_2976);
nor UO_433 (O_433,N_2971,N_2999);
nand UO_434 (O_434,N_2973,N_2950);
or UO_435 (O_435,N_2972,N_2987);
or UO_436 (O_436,N_2972,N_2963);
nand UO_437 (O_437,N_2978,N_2971);
and UO_438 (O_438,N_2946,N_2949);
or UO_439 (O_439,N_2958,N_2991);
or UO_440 (O_440,N_2968,N_2949);
and UO_441 (O_441,N_2990,N_2984);
and UO_442 (O_442,N_2961,N_2990);
nand UO_443 (O_443,N_2982,N_2986);
and UO_444 (O_444,N_2949,N_2967);
nor UO_445 (O_445,N_2996,N_2995);
or UO_446 (O_446,N_2977,N_2968);
or UO_447 (O_447,N_2995,N_2943);
nor UO_448 (O_448,N_2985,N_2993);
and UO_449 (O_449,N_2946,N_2992);
xnor UO_450 (O_450,N_2953,N_2989);
nor UO_451 (O_451,N_2978,N_2998);
and UO_452 (O_452,N_2970,N_2943);
or UO_453 (O_453,N_2974,N_2947);
or UO_454 (O_454,N_2957,N_2965);
nand UO_455 (O_455,N_2950,N_2995);
or UO_456 (O_456,N_2961,N_2971);
and UO_457 (O_457,N_2944,N_2969);
or UO_458 (O_458,N_2978,N_2973);
or UO_459 (O_459,N_2975,N_2995);
and UO_460 (O_460,N_2978,N_2968);
and UO_461 (O_461,N_2945,N_2998);
nor UO_462 (O_462,N_2991,N_2973);
nor UO_463 (O_463,N_2945,N_2947);
and UO_464 (O_464,N_2995,N_2945);
nand UO_465 (O_465,N_2945,N_2999);
nand UO_466 (O_466,N_2986,N_2991);
and UO_467 (O_467,N_2982,N_2961);
and UO_468 (O_468,N_2956,N_2950);
and UO_469 (O_469,N_2966,N_2953);
and UO_470 (O_470,N_2945,N_2989);
or UO_471 (O_471,N_2942,N_2948);
or UO_472 (O_472,N_2972,N_2941);
nand UO_473 (O_473,N_2980,N_2943);
or UO_474 (O_474,N_2958,N_2985);
and UO_475 (O_475,N_2997,N_2969);
and UO_476 (O_476,N_2975,N_2946);
and UO_477 (O_477,N_2981,N_2976);
nand UO_478 (O_478,N_2960,N_2995);
or UO_479 (O_479,N_2956,N_2943);
nand UO_480 (O_480,N_2973,N_2997);
nor UO_481 (O_481,N_2970,N_2989);
nand UO_482 (O_482,N_2984,N_2951);
or UO_483 (O_483,N_2945,N_2992);
nor UO_484 (O_484,N_2981,N_2958);
or UO_485 (O_485,N_2983,N_2944);
nor UO_486 (O_486,N_2941,N_2968);
nand UO_487 (O_487,N_2992,N_2952);
nor UO_488 (O_488,N_2972,N_2945);
or UO_489 (O_489,N_2972,N_2966);
nand UO_490 (O_490,N_2985,N_2975);
xor UO_491 (O_491,N_2943,N_2996);
or UO_492 (O_492,N_2940,N_2949);
or UO_493 (O_493,N_2941,N_2966);
nor UO_494 (O_494,N_2993,N_2970);
or UO_495 (O_495,N_2962,N_2960);
nand UO_496 (O_496,N_2953,N_2958);
nor UO_497 (O_497,N_2956,N_2993);
and UO_498 (O_498,N_2993,N_2971);
and UO_499 (O_499,N_2999,N_2991);
endmodule