module basic_1500_15000_2000_5_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1269,In_883);
nor U1 (N_1,In_867,In_1295);
nand U2 (N_2,In_1199,In_54);
nor U3 (N_3,In_22,In_1244);
or U4 (N_4,In_1222,In_835);
or U5 (N_5,In_1322,In_485);
and U6 (N_6,In_1133,In_56);
nor U7 (N_7,In_7,In_875);
nand U8 (N_8,In_1487,In_28);
nor U9 (N_9,In_925,In_1006);
and U10 (N_10,In_193,In_1448);
nand U11 (N_11,In_598,In_824);
and U12 (N_12,In_618,In_1426);
and U13 (N_13,In_154,In_335);
and U14 (N_14,In_1052,In_1441);
nor U15 (N_15,In_669,In_146);
nand U16 (N_16,In_1039,In_434);
or U17 (N_17,In_1323,In_223);
nor U18 (N_18,In_619,In_164);
and U19 (N_19,In_869,In_15);
nand U20 (N_20,In_581,In_499);
or U21 (N_21,In_169,In_887);
and U22 (N_22,In_594,In_293);
and U23 (N_23,In_543,In_3);
nand U24 (N_24,In_1086,In_329);
or U25 (N_25,In_593,In_641);
or U26 (N_26,In_857,In_799);
nor U27 (N_27,In_988,In_989);
nand U28 (N_28,In_791,In_209);
and U29 (N_29,In_1012,In_916);
or U30 (N_30,In_936,In_100);
nor U31 (N_31,In_1210,In_592);
nor U32 (N_32,In_966,In_433);
nand U33 (N_33,In_938,In_905);
nor U34 (N_34,In_348,In_745);
nor U35 (N_35,In_773,In_1185);
nand U36 (N_36,In_275,In_1471);
nor U37 (N_37,In_784,In_698);
nor U38 (N_38,In_2,In_970);
xnor U39 (N_39,In_1241,In_334);
nand U40 (N_40,In_1394,In_397);
nor U41 (N_41,In_1071,In_555);
or U42 (N_42,In_113,In_1449);
nor U43 (N_43,In_1396,In_263);
nand U44 (N_44,In_688,In_554);
nand U45 (N_45,In_294,In_1499);
and U46 (N_46,In_70,In_468);
nor U47 (N_47,In_1351,In_1255);
and U48 (N_48,In_1137,In_336);
and U49 (N_49,In_1380,In_785);
or U50 (N_50,In_980,In_390);
nor U51 (N_51,In_347,In_179);
and U52 (N_52,In_261,In_591);
and U53 (N_53,In_1458,In_1000);
nand U54 (N_54,In_1319,In_231);
nand U55 (N_55,In_958,In_333);
or U56 (N_56,In_1250,In_354);
nand U57 (N_57,In_913,In_508);
nand U58 (N_58,In_1212,In_291);
nor U59 (N_59,In_38,In_901);
or U60 (N_60,In_77,In_675);
and U61 (N_61,In_1324,In_663);
nand U62 (N_62,In_166,In_821);
and U63 (N_63,In_626,In_622);
and U64 (N_64,In_1248,In_1034);
nand U65 (N_65,In_64,In_1390);
nor U66 (N_66,In_488,In_1329);
or U67 (N_67,In_1206,In_378);
nor U68 (N_68,In_1285,In_1371);
nand U69 (N_69,In_631,In_1013);
and U70 (N_70,In_1171,In_599);
xor U71 (N_71,In_415,In_221);
nor U72 (N_72,In_740,In_1294);
nand U73 (N_73,In_1454,In_476);
nand U74 (N_74,In_1313,In_1409);
and U75 (N_75,In_601,In_803);
nand U76 (N_76,In_86,In_1189);
nor U77 (N_77,In_426,In_888);
nand U78 (N_78,In_482,In_1433);
nor U79 (N_79,In_123,In_802);
or U80 (N_80,In_1003,In_1218);
and U81 (N_81,In_1138,In_1361);
nor U82 (N_82,In_98,In_1015);
and U83 (N_83,In_1498,In_705);
nand U84 (N_84,In_199,In_1427);
nand U85 (N_85,In_1221,In_501);
and U86 (N_86,In_246,In_122);
nor U87 (N_87,In_1372,In_1431);
and U88 (N_88,In_1419,In_300);
or U89 (N_89,In_420,In_232);
and U90 (N_90,In_227,In_1173);
nor U91 (N_91,In_578,In_854);
and U92 (N_92,In_1273,In_1050);
nor U93 (N_93,In_818,In_617);
nand U94 (N_94,In_837,In_142);
nand U95 (N_95,In_878,In_521);
or U96 (N_96,In_523,In_832);
nand U97 (N_97,In_1475,In_764);
nand U98 (N_98,In_345,In_1169);
and U99 (N_99,In_74,In_915);
and U100 (N_100,In_121,In_165);
and U101 (N_101,In_949,In_944);
and U102 (N_102,In_1280,In_1094);
nand U103 (N_103,In_406,In_519);
nand U104 (N_104,In_575,In_322);
or U105 (N_105,In_253,In_666);
nand U106 (N_106,In_349,In_537);
nand U107 (N_107,In_1192,In_1074);
nor U108 (N_108,In_877,In_224);
nand U109 (N_109,In_206,In_360);
nand U110 (N_110,In_1252,In_811);
nand U111 (N_111,In_961,In_1115);
nor U112 (N_112,In_50,In_481);
and U113 (N_113,In_1110,In_409);
nor U114 (N_114,In_1165,In_1155);
or U115 (N_115,In_82,In_67);
or U116 (N_116,In_1331,In_829);
and U117 (N_117,In_731,In_89);
nor U118 (N_118,In_1293,In_14);
nor U119 (N_119,In_385,In_690);
nor U120 (N_120,In_244,In_393);
and U121 (N_121,In_573,In_1384);
nor U122 (N_122,In_946,In_1335);
nand U123 (N_123,In_1057,In_1379);
or U124 (N_124,In_391,In_369);
nand U125 (N_125,In_107,In_110);
and U126 (N_126,In_1164,In_881);
and U127 (N_127,In_104,In_1166);
nand U128 (N_128,In_1044,In_1075);
nand U129 (N_129,In_967,In_1307);
xor U130 (N_130,In_282,In_724);
nand U131 (N_131,In_853,In_1183);
nand U132 (N_132,In_274,In_583);
xor U133 (N_133,In_342,In_845);
nor U134 (N_134,In_407,In_1438);
nand U135 (N_135,In_553,In_161);
and U136 (N_136,In_187,In_356);
and U137 (N_137,In_590,In_928);
nor U138 (N_138,In_569,In_1453);
or U139 (N_139,In_475,In_68);
nand U140 (N_140,In_295,In_1435);
nor U141 (N_141,In_712,In_339);
nand U142 (N_142,In_582,In_789);
nor U143 (N_143,In_1211,In_242);
or U144 (N_144,In_621,In_260);
nand U145 (N_145,In_305,In_262);
nor U146 (N_146,In_1456,In_115);
and U147 (N_147,In_504,In_1434);
nand U148 (N_148,In_126,In_235);
nand U149 (N_149,In_96,In_341);
and U150 (N_150,In_132,In_1200);
nor U151 (N_151,In_1108,In_167);
nand U152 (N_152,In_425,In_328);
xor U153 (N_153,In_754,In_536);
or U154 (N_154,In_463,In_1144);
nand U155 (N_155,In_408,In_384);
nand U156 (N_156,In_456,In_88);
and U157 (N_157,In_195,In_1385);
or U158 (N_158,In_93,In_823);
or U159 (N_159,In_302,In_664);
or U160 (N_160,In_672,In_1024);
nand U161 (N_161,In_494,In_924);
and U162 (N_162,In_171,In_612);
nor U163 (N_163,In_184,In_251);
nor U164 (N_164,In_1367,In_1151);
and U165 (N_165,In_95,In_984);
nor U166 (N_166,In_927,In_529);
nand U167 (N_167,In_674,In_911);
nor U168 (N_168,In_549,In_368);
nor U169 (N_169,In_1276,In_831);
and U170 (N_170,In_480,In_604);
and U171 (N_171,In_822,In_758);
or U172 (N_172,In_1261,In_752);
or U173 (N_173,In_284,In_280);
or U174 (N_174,In_114,In_816);
and U175 (N_175,In_140,In_388);
and U176 (N_176,In_863,In_846);
nand U177 (N_177,In_493,In_131);
nand U178 (N_178,In_1227,In_42);
nand U179 (N_179,In_891,In_646);
nand U180 (N_180,In_37,In_820);
xor U181 (N_181,In_1047,In_999);
nand U182 (N_182,In_239,In_185);
nand U183 (N_183,In_834,In_1135);
and U184 (N_184,In_254,In_212);
nor U185 (N_185,In_704,In_40);
nor U186 (N_186,In_1181,In_671);
nor U187 (N_187,In_807,In_1093);
or U188 (N_188,In_1021,In_511);
nand U189 (N_189,In_1387,In_1207);
and U190 (N_190,In_1466,In_895);
nor U191 (N_191,In_1179,In_661);
nor U192 (N_192,In_1298,In_948);
or U193 (N_193,In_323,In_57);
or U194 (N_194,In_325,In_781);
and U195 (N_195,In_365,In_80);
nand U196 (N_196,In_1123,In_1172);
nor U197 (N_197,In_484,In_782);
nand U198 (N_198,In_1083,In_1051);
and U199 (N_199,In_588,In_30);
xor U200 (N_200,In_1381,In_897);
nand U201 (N_201,In_1026,In_1481);
or U202 (N_202,In_196,In_547);
or U203 (N_203,In_910,In_1393);
nor U204 (N_204,In_1321,In_906);
nand U205 (N_205,In_440,In_733);
or U206 (N_206,In_1496,In_136);
nand U207 (N_207,In_205,In_163);
or U208 (N_208,In_699,In_902);
and U209 (N_209,In_252,In_686);
and U210 (N_210,In_116,In_934);
or U211 (N_211,In_1242,In_483);
or U212 (N_212,In_375,In_848);
and U213 (N_213,In_1405,In_85);
or U214 (N_214,In_978,In_1437);
and U215 (N_215,In_1160,In_1343);
and U216 (N_216,In_862,In_311);
or U217 (N_217,In_654,In_1220);
or U218 (N_218,In_1247,In_377);
nor U219 (N_219,In_1373,In_492);
nand U220 (N_220,In_792,In_1492);
nand U221 (N_221,In_1127,In_1283);
and U222 (N_222,In_880,In_531);
or U223 (N_223,In_35,In_505);
nand U224 (N_224,In_1476,In_540);
nand U225 (N_225,In_701,In_932);
and U226 (N_226,In_138,In_574);
and U227 (N_227,In_1272,In_296);
nand U228 (N_228,In_1326,In_1254);
nand U229 (N_229,In_361,In_1484);
and U230 (N_230,In_909,In_1215);
and U231 (N_231,In_744,In_662);
nand U232 (N_232,In_659,In_9);
nand U233 (N_233,In_1424,In_1100);
xnor U234 (N_234,In_614,In_1256);
and U235 (N_235,In_616,In_1359);
or U236 (N_236,In_315,In_1187);
nor U237 (N_237,In_422,In_903);
nor U238 (N_238,In_117,In_931);
nor U239 (N_239,In_145,In_213);
nand U240 (N_240,In_1461,In_387);
and U241 (N_241,In_49,In_1445);
or U242 (N_242,In_1062,In_552);
nand U243 (N_243,In_1099,In_1490);
or U244 (N_244,In_1447,In_746);
and U245 (N_245,In_33,In_797);
nand U246 (N_246,In_1091,In_429);
and U247 (N_247,In_873,In_147);
nor U248 (N_248,In_370,In_1286);
nand U249 (N_249,In_933,In_861);
and U250 (N_250,In_678,In_1300);
nor U251 (N_251,In_1344,In_525);
nor U252 (N_252,In_884,In_747);
nor U253 (N_253,In_860,In_279);
or U254 (N_254,In_995,In_1347);
or U255 (N_255,In_1129,In_65);
nor U256 (N_256,In_730,In_1180);
xnor U257 (N_257,In_776,In_1414);
and U258 (N_258,In_1284,In_1401);
nor U259 (N_259,In_798,In_542);
or U260 (N_260,In_1131,In_844);
and U261 (N_261,In_700,In_180);
nand U262 (N_262,In_450,In_75);
and U263 (N_263,In_84,In_697);
nor U264 (N_264,In_1463,In_177);
or U265 (N_265,In_608,In_1031);
and U266 (N_266,In_804,In_1443);
nand U267 (N_267,In_351,In_1305);
nor U268 (N_268,In_1375,In_689);
or U269 (N_269,In_265,In_577);
and U270 (N_270,In_108,In_1428);
and U271 (N_271,In_1098,In_1216);
and U272 (N_272,In_723,In_1146);
and U273 (N_273,In_1364,In_930);
and U274 (N_274,In_269,In_1362);
or U275 (N_275,In_1193,In_632);
or U276 (N_276,In_1067,In_1028);
and U277 (N_277,In_1400,In_418);
nand U278 (N_278,In_1469,In_973);
nor U279 (N_279,In_722,In_44);
nand U280 (N_280,In_1395,In_1310);
xnor U281 (N_281,In_1230,In_139);
or U282 (N_282,In_1337,In_445);
nor U283 (N_283,In_1336,In_273);
or U284 (N_284,In_864,In_1489);
and U285 (N_285,In_1494,In_994);
or U286 (N_286,In_696,In_448);
and U287 (N_287,In_320,In_120);
and U288 (N_288,In_653,In_10);
nor U289 (N_289,In_47,In_228);
nand U290 (N_290,In_1260,In_623);
nand U291 (N_291,In_1111,In_158);
or U292 (N_292,In_130,In_992);
nand U293 (N_293,In_1355,In_1332);
nor U294 (N_294,In_214,In_528);
nand U295 (N_295,In_585,In_477);
or U296 (N_296,In_951,In_935);
or U297 (N_297,In_278,In_1188);
nand U298 (N_298,In_976,In_1081);
nor U299 (N_299,In_1069,In_691);
nand U300 (N_300,In_457,In_996);
nand U301 (N_301,In_676,In_550);
nand U302 (N_302,In_306,In_1402);
and U303 (N_303,In_1114,In_371);
nand U304 (N_304,In_917,In_400);
nand U305 (N_305,In_1495,In_1366);
nor U306 (N_306,In_684,In_219);
nor U307 (N_307,In_124,In_486);
and U308 (N_308,In_413,In_1148);
and U309 (N_309,In_739,In_726);
and U310 (N_310,In_1061,In_292);
or U311 (N_311,In_685,In_1229);
or U312 (N_312,In_372,In_1035);
nand U313 (N_313,In_1368,In_1464);
nand U314 (N_314,In_204,In_1140);
nor U315 (N_315,In_90,In_1238);
nand U316 (N_316,In_506,In_17);
and U317 (N_317,In_1334,In_367);
nor U318 (N_318,In_979,In_299);
and U319 (N_319,In_1059,In_497);
nand U320 (N_320,In_896,In_959);
nor U321 (N_321,In_1142,In_827);
or U322 (N_322,In_937,In_637);
or U323 (N_323,In_383,In_101);
and U324 (N_324,In_725,In_1198);
nor U325 (N_325,In_419,In_756);
and U326 (N_326,In_133,In_940);
or U327 (N_327,In_62,In_514);
nor U328 (N_328,In_743,In_1446);
nor U329 (N_329,In_1297,In_1234);
nand U330 (N_330,In_836,In_1411);
and U331 (N_331,In_317,In_358);
or U332 (N_332,In_1124,In_668);
nor U333 (N_333,In_711,In_1485);
nor U334 (N_334,In_783,In_527);
or U335 (N_335,In_1262,In_424);
nor U336 (N_336,In_589,In_962);
nand U337 (N_337,In_83,In_211);
or U338 (N_338,In_355,In_1136);
or U339 (N_339,In_258,In_229);
nor U340 (N_340,In_1415,In_324);
nor U341 (N_341,In_283,In_1432);
nand U342 (N_342,In_469,In_713);
nor U343 (N_343,In_1048,In_314);
and U344 (N_344,In_1328,In_941);
nor U345 (N_345,In_1041,In_562);
or U346 (N_346,In_694,In_738);
nor U347 (N_347,In_777,In_210);
and U348 (N_348,In_330,In_1346);
nor U349 (N_349,In_148,In_718);
nor U350 (N_350,In_498,In_234);
or U351 (N_351,In_12,In_414);
nor U352 (N_352,In_503,In_1232);
nand U353 (N_353,In_1315,In_1259);
nor U354 (N_354,In_1491,In_1226);
nor U355 (N_355,In_868,In_45);
or U356 (N_356,In_629,In_1002);
or U357 (N_357,In_410,In_1042);
nor U358 (N_358,In_264,In_1444);
and U359 (N_359,In_183,In_1060);
or U360 (N_360,In_1376,In_1270);
and U361 (N_361,In_471,In_1406);
and U362 (N_362,In_735,In_1065);
and U363 (N_363,In_1420,In_765);
or U364 (N_364,In_1175,In_1090);
nor U365 (N_365,In_952,In_1350);
and U366 (N_366,In_702,In_1084);
nand U367 (N_367,In_97,In_1007);
and U368 (N_368,In_1416,In_1078);
nor U369 (N_369,In_660,In_36);
or U370 (N_370,In_1116,In_1479);
nor U371 (N_371,In_975,In_1309);
and U372 (N_372,In_99,In_1149);
and U373 (N_373,In_741,In_1388);
or U374 (N_374,In_1205,In_230);
nand U375 (N_375,In_796,In_1145);
and U376 (N_376,In_431,In_1243);
and U377 (N_377,In_26,In_865);
nand U378 (N_378,In_380,In_833);
nand U379 (N_379,In_1077,In_551);
nand U380 (N_380,In_805,In_399);
and U381 (N_381,In_137,In_257);
nor U382 (N_382,In_1055,In_401);
nand U383 (N_383,In_518,In_1287);
nor U384 (N_384,In_1195,In_808);
and U385 (N_385,In_1001,In_855);
nand U386 (N_386,In_1157,In_182);
or U387 (N_387,In_1455,In_1036);
and U388 (N_388,In_1143,In_268);
and U389 (N_389,In_708,In_1056);
nor U390 (N_390,In_1457,In_247);
and U391 (N_391,In_771,In_533);
nand U392 (N_392,In_1167,In_449);
and U393 (N_393,In_1472,In_879);
nor U394 (N_394,In_412,In_48);
nand U395 (N_395,In_289,In_1023);
and U396 (N_396,In_568,In_125);
nand U397 (N_397,In_715,In_1085);
nand U398 (N_398,In_404,In_770);
nand U399 (N_399,In_918,In_1153);
nor U400 (N_400,In_545,In_1352);
nand U401 (N_401,In_645,In_1089);
and U402 (N_402,In_1019,In_1080);
or U403 (N_403,In_59,In_395);
nand U404 (N_404,In_255,In_312);
nor U405 (N_405,In_1330,In_670);
and U406 (N_406,In_872,In_843);
nand U407 (N_407,In_21,In_60);
and U408 (N_408,In_597,In_673);
or U409 (N_409,In_198,In_814);
nand U410 (N_410,In_203,In_331);
or U411 (N_411,In_510,In_517);
nor U412 (N_412,In_579,In_319);
nor U413 (N_413,In_1049,In_1263);
and U414 (N_414,In_815,In_1082);
nand U415 (N_415,In_226,In_178);
or U416 (N_416,In_1308,In_584);
or U417 (N_417,In_892,In_627);
or U418 (N_418,In_301,In_1119);
nor U419 (N_419,In_972,In_478);
nand U420 (N_420,In_11,In_162);
nand U421 (N_421,In_611,In_1105);
and U422 (N_422,In_866,In_728);
and U423 (N_423,In_1468,In_1325);
and U424 (N_424,In_600,In_1004);
or U425 (N_425,In_859,In_403);
nor U426 (N_426,In_1407,In_1480);
nand U427 (N_427,In_382,In_141);
and U428 (N_428,In_516,In_29);
or U429 (N_429,In_1404,In_960);
and U430 (N_430,In_1070,In_1277);
or U431 (N_431,In_1374,In_774);
nor U432 (N_432,In_1271,In_462);
or U433 (N_433,In_1152,In_602);
and U434 (N_434,In_24,In_520);
nor U435 (N_435,In_1132,In_858);
and U436 (N_436,In_649,In_767);
and U437 (N_437,In_19,In_241);
nand U438 (N_438,In_1470,In_1306);
and U439 (N_439,In_1194,In_454);
nand U440 (N_440,In_1101,In_455);
and U441 (N_441,In_338,In_1303);
and U442 (N_442,In_248,In_1391);
or U443 (N_443,In_428,In_373);
or U444 (N_444,In_321,In_32);
and U445 (N_445,In_460,In_298);
nand U446 (N_446,In_706,In_716);
and U447 (N_447,In_1029,In_526);
nand U448 (N_448,In_1097,In_495);
and U449 (N_449,In_838,In_587);
and U450 (N_450,In_344,In_751);
nand U451 (N_451,In_216,In_559);
nor U452 (N_452,In_775,In_515);
nor U453 (N_453,In_1312,In_222);
or U454 (N_454,In_969,In_566);
nor U455 (N_455,In_558,In_633);
and U456 (N_456,In_1289,In_1473);
or U457 (N_457,In_532,In_1095);
nand U458 (N_458,In_0,In_172);
nor U459 (N_459,In_309,In_237);
nand U460 (N_460,In_806,In_544);
and U461 (N_461,In_652,In_290);
nand U462 (N_462,In_1282,In_1249);
or U463 (N_463,In_826,In_638);
nor U464 (N_464,In_1304,In_1073);
and U465 (N_465,In_1488,In_427);
nand U466 (N_466,In_1349,In_692);
nor U467 (N_467,In_386,In_1314);
and U468 (N_468,In_1421,In_755);
nand U469 (N_469,In_1239,In_452);
nand U470 (N_470,In_129,In_1122);
nand U471 (N_471,In_899,In_613);
xnor U472 (N_472,In_150,In_557);
nand U473 (N_473,In_467,In_956);
and U474 (N_474,In_1235,In_39);
xnor U475 (N_475,In_907,In_565);
nand U476 (N_476,In_453,In_1253);
and U477 (N_477,In_742,In_1369);
nand U478 (N_478,In_656,In_893);
nand U479 (N_479,In_856,In_363);
and U480 (N_480,In_636,In_190);
and U481 (N_481,In_990,In_1162);
nand U482 (N_482,In_1125,In_849);
or U483 (N_483,In_556,In_159);
nand U484 (N_484,In_1037,In_174);
nor U485 (N_485,In_1465,In_103);
nand U486 (N_486,In_233,In_761);
and U487 (N_487,In_939,In_1178);
and U488 (N_488,In_507,In_977);
and U489 (N_489,In_1202,In_1408);
nor U490 (N_490,In_1345,In_1267);
xor U491 (N_491,In_680,In_825);
nor U492 (N_492,In_795,In_446);
and U493 (N_493,In_55,In_625);
and U494 (N_494,In_762,In_1030);
nand U495 (N_495,In_1079,In_281);
or U496 (N_496,In_658,In_69);
and U497 (N_497,In_1112,In_522);
nand U498 (N_498,In_560,In_644);
nor U499 (N_499,In_191,In_46);
and U500 (N_500,In_197,In_719);
nor U501 (N_501,In_635,In_615);
nand U502 (N_502,In_679,In_1482);
or U503 (N_503,In_1186,In_398);
or U504 (N_504,In_71,In_303);
nand U505 (N_505,In_451,In_1474);
nor U506 (N_506,In_405,In_595);
and U507 (N_507,In_1225,In_1266);
or U508 (N_508,In_470,In_1291);
or U509 (N_509,In_530,In_1452);
and U510 (N_510,In_882,In_466);
and U511 (N_511,In_416,In_1333);
or U512 (N_512,In_667,In_548);
nor U513 (N_513,In_240,In_1104);
nand U514 (N_514,In_359,In_465);
and U515 (N_515,In_220,In_987);
nand U516 (N_516,In_357,In_1348);
and U517 (N_517,In_326,In_432);
nand U518 (N_518,In_1190,In_238);
or U519 (N_519,In_25,In_648);
and U520 (N_520,In_1054,In_1117);
nor U521 (N_521,In_1292,In_52);
or U522 (N_522,In_687,In_479);
or U523 (N_523,In_812,In_1360);
or U524 (N_524,In_1040,In_763);
nor U525 (N_525,In_1316,In_156);
and U526 (N_526,In_852,In_374);
nand U527 (N_527,In_778,In_1017);
nor U528 (N_528,In_58,In_986);
and U529 (N_529,In_693,In_1340);
nand U530 (N_530,In_102,In_707);
and U531 (N_531,In_474,In_1413);
nor U532 (N_532,In_630,In_842);
or U533 (N_533,In_1161,In_605);
and U534 (N_534,In_1422,In_1296);
and U535 (N_535,In_308,In_421);
nand U536 (N_536,In_423,In_1302);
or U537 (N_537,In_851,In_586);
or U538 (N_538,In_394,In_921);
nand U539 (N_539,In_717,In_1436);
nor U540 (N_540,In_974,In_218);
and U541 (N_541,In_639,In_955);
xnor U542 (N_542,In_1356,In_152);
nor U543 (N_543,In_160,In_1109);
nor U544 (N_544,In_41,In_118);
nor U545 (N_545,In_847,In_297);
or U546 (N_546,In_176,In_327);
or U547 (N_547,In_61,In_1182);
and U548 (N_548,In_1288,In_695);
nor U549 (N_549,In_997,In_1128);
and U550 (N_550,In_1442,In_8);
nor U551 (N_551,In_111,In_1354);
nand U552 (N_552,In_817,In_749);
nand U553 (N_553,In_1231,In_642);
nand U554 (N_554,In_491,In_1196);
or U555 (N_555,In_1009,In_1020);
nor U556 (N_556,In_106,In_1423);
or U557 (N_557,In_1478,In_1311);
and U558 (N_558,In_620,In_1320);
and U559 (N_559,In_993,In_524);
and U560 (N_560,In_801,In_874);
nor U561 (N_561,In_721,In_79);
or U562 (N_562,In_208,In_634);
or U563 (N_563,In_596,In_535);
nand U564 (N_564,In_541,In_43);
nor U565 (N_565,In_1043,In_1156);
or U566 (N_566,In_571,In_603);
nand U567 (N_567,In_1209,In_270);
or U568 (N_568,In_245,In_119);
nor U569 (N_569,In_1378,In_828);
or U570 (N_570,In_1197,In_157);
nor U571 (N_571,In_364,In_13);
nor U572 (N_572,In_1258,In_607);
nor U573 (N_573,In_1403,In_1);
and U574 (N_574,In_1102,In_1168);
and U575 (N_575,In_1058,In_1275);
or U576 (N_576,In_1365,In_1163);
and U577 (N_577,In_950,In_1451);
nand U578 (N_578,In_168,In_1107);
and U579 (N_579,In_800,In_1213);
nor U580 (N_580,In_1011,In_563);
nand U581 (N_581,In_982,In_175);
nor U582 (N_582,In_1016,In_362);
xor U583 (N_583,In_105,In_1045);
nor U584 (N_584,In_1363,In_1341);
and U585 (N_585,In_173,In_1066);
nand U586 (N_586,In_1439,In_1204);
xor U587 (N_587,In_1228,In_912);
or U588 (N_588,In_683,In_1223);
and U589 (N_589,In_650,In_63);
nor U590 (N_590,In_332,In_310);
nor U591 (N_591,In_128,In_1279);
and U592 (N_592,In_819,In_1224);
nand U593 (N_593,In_780,In_538);
and U594 (N_594,In_285,In_436);
or U595 (N_595,In_34,In_144);
nand U596 (N_596,In_734,In_813);
nand U597 (N_597,In_1008,In_983);
xnor U598 (N_598,In_1383,In_442);
nand U599 (N_599,In_1106,In_947);
or U600 (N_600,In_447,In_968);
nand U601 (N_601,In_1038,In_441);
nor U602 (N_602,In_1278,In_1025);
nand U603 (N_603,In_91,In_23);
and U604 (N_604,In_1072,In_886);
and U605 (N_605,In_1134,In_720);
and U606 (N_606,In_16,In_981);
nand U607 (N_607,In_710,In_243);
and U608 (N_608,In_1150,In_954);
or U609 (N_609,In_1005,In_92);
nand U610 (N_610,In_337,In_1068);
or U611 (N_611,In_443,In_1064);
and U612 (N_612,In_458,In_277);
or U613 (N_613,In_841,In_963);
nor U614 (N_614,In_760,In_271);
nor U615 (N_615,In_18,In_1177);
or U616 (N_616,In_1440,In_657);
nor U617 (N_617,In_1397,In_610);
nor U618 (N_618,In_1317,In_438);
nand U619 (N_619,In_922,In_1410);
and U620 (N_620,In_496,In_435);
nor U621 (N_621,In_489,In_509);
or U622 (N_622,In_76,In_1301);
nor U623 (N_623,In_215,In_53);
or U624 (N_624,In_766,In_757);
nor U625 (N_625,In_153,In_1268);
or U626 (N_626,In_1237,In_1327);
and U627 (N_627,In_87,In_748);
nand U628 (N_628,In_1339,In_31);
nand U629 (N_629,In_1233,In_1154);
nand U630 (N_630,In_1033,In_1096);
or U631 (N_631,In_1357,In_402);
nor U632 (N_632,In_1382,In_727);
nand U633 (N_633,In_272,In_376);
or U634 (N_634,In_1113,In_1417);
nand U635 (N_635,In_640,In_192);
nand U636 (N_636,In_1118,In_1398);
and U637 (N_637,In_1076,In_1486);
nand U638 (N_638,In_1170,In_628);
or U639 (N_639,In_1412,In_769);
or U640 (N_640,In_259,In_904);
nand U641 (N_641,In_1022,In_1264);
nor U642 (N_642,In_759,In_437);
nor U643 (N_643,In_236,In_267);
nand U644 (N_644,In_201,In_5);
or U645 (N_645,In_1208,In_1018);
and U646 (N_646,In_304,In_189);
nand U647 (N_647,In_151,In_66);
nand U648 (N_648,In_287,In_1418);
nand U649 (N_649,In_473,In_73);
nand U650 (N_650,In_225,In_965);
nand U651 (N_651,In_1184,In_1121);
and U652 (N_652,In_1450,In_643);
and U653 (N_653,In_170,In_112);
nand U654 (N_654,In_1088,In_1399);
or U655 (N_655,In_266,In_894);
and U656 (N_656,In_561,In_500);
nand U657 (N_657,In_459,In_1265);
or U658 (N_658,In_1203,In_1460);
nor U659 (N_659,In_72,In_1027);
and U660 (N_660,In_971,In_1274);
or U661 (N_661,In_1386,In_564);
or U662 (N_662,In_155,In_256);
nor U663 (N_663,In_786,In_839);
or U664 (N_664,In_1087,In_1147);
or U665 (N_665,In_889,In_1299);
nand U666 (N_666,In_1158,In_188);
nand U667 (N_667,In_127,In_1139);
and U668 (N_668,In_346,In_513);
nand U669 (N_669,In_4,In_809);
or U670 (N_670,In_714,In_651);
nor U671 (N_671,In_350,In_194);
nand U672 (N_672,In_1217,In_109);
and U673 (N_673,In_249,In_900);
and U674 (N_674,In_1462,In_1141);
nor U675 (N_675,In_461,In_709);
or U676 (N_676,In_1290,In_1201);
nor U677 (N_677,In_94,In_576);
nor U678 (N_678,In_366,In_20);
and U679 (N_679,In_1493,In_444);
nand U680 (N_680,In_1467,In_343);
nor U681 (N_681,In_472,In_953);
or U682 (N_682,In_181,In_957);
and U683 (N_683,In_250,In_840);
nor U684 (N_684,In_27,In_655);
and U685 (N_685,In_1358,In_1389);
nor U686 (N_686,In_81,In_307);
and U687 (N_687,In_1032,In_772);
or U688 (N_688,In_647,In_991);
nand U689 (N_689,In_1483,In_682);
nand U690 (N_690,In_464,In_736);
and U691 (N_691,In_353,In_539);
nand U692 (N_692,In_810,In_964);
and U693 (N_693,In_313,In_134);
nor U694 (N_694,In_787,In_1014);
or U695 (N_695,In_929,In_487);
nor U696 (N_696,In_502,In_830);
nand U697 (N_697,In_677,In_430);
nand U698 (N_698,In_919,In_512);
or U699 (N_699,In_1236,In_737);
or U700 (N_700,In_318,In_396);
and U701 (N_701,In_871,In_217);
and U702 (N_702,In_790,In_945);
nor U703 (N_703,In_779,In_943);
nor U704 (N_704,In_1053,In_316);
and U705 (N_705,In_567,In_1318);
nand U706 (N_706,In_876,In_920);
nand U707 (N_707,In_288,In_1214);
nand U708 (N_708,In_624,In_1281);
and U709 (N_709,In_890,In_143);
nand U710 (N_710,In_850,In_1219);
nor U711 (N_711,In_914,In_379);
and U712 (N_712,In_609,In_276);
nand U713 (N_713,In_1392,In_923);
and U714 (N_714,In_1338,In_6);
nor U715 (N_715,In_665,In_1459);
nand U716 (N_716,In_51,In_729);
and U717 (N_717,In_135,In_570);
or U718 (N_718,In_985,In_202);
and U719 (N_719,In_926,In_942);
or U720 (N_720,In_546,In_753);
nor U721 (N_721,In_534,In_200);
nand U722 (N_722,In_1370,In_207);
nand U723 (N_723,In_1497,In_1430);
and U724 (N_724,In_149,In_1377);
nand U725 (N_725,In_186,In_681);
nand U726 (N_726,In_78,In_1342);
and U727 (N_727,In_1174,In_788);
or U728 (N_728,In_606,In_703);
or U729 (N_729,In_1130,In_580);
and U730 (N_730,In_1257,In_389);
or U731 (N_731,In_750,In_1246);
or U732 (N_732,In_1425,In_1251);
or U733 (N_733,In_1429,In_417);
nand U734 (N_734,In_1159,In_794);
nor U735 (N_735,In_340,In_286);
and U736 (N_736,In_411,In_1477);
and U737 (N_737,In_1176,In_381);
nand U738 (N_738,In_392,In_490);
and U739 (N_739,In_793,In_1245);
and U740 (N_740,In_998,In_732);
and U741 (N_741,In_352,In_885);
nor U742 (N_742,In_870,In_1010);
nor U743 (N_743,In_1191,In_1046);
or U744 (N_744,In_768,In_908);
nor U745 (N_745,In_572,In_1063);
nand U746 (N_746,In_1353,In_439);
xnor U747 (N_747,In_1240,In_898);
nor U748 (N_748,In_1103,In_1120);
or U749 (N_749,In_1126,In_1092);
nor U750 (N_750,In_387,In_1266);
nor U751 (N_751,In_1303,In_1220);
and U752 (N_752,In_828,In_1467);
nor U753 (N_753,In_1431,In_265);
xor U754 (N_754,In_802,In_1122);
nand U755 (N_755,In_1196,In_1233);
and U756 (N_756,In_1374,In_422);
or U757 (N_757,In_1473,In_696);
and U758 (N_758,In_516,In_1360);
and U759 (N_759,In_786,In_340);
nand U760 (N_760,In_1060,In_307);
or U761 (N_761,In_1435,In_129);
or U762 (N_762,In_1178,In_1055);
or U763 (N_763,In_181,In_1047);
or U764 (N_764,In_604,In_1381);
and U765 (N_765,In_828,In_136);
nand U766 (N_766,In_1331,In_1231);
and U767 (N_767,In_418,In_83);
or U768 (N_768,In_1090,In_59);
nand U769 (N_769,In_657,In_397);
nand U770 (N_770,In_1249,In_1046);
xnor U771 (N_771,In_867,In_14);
and U772 (N_772,In_505,In_1440);
and U773 (N_773,In_150,In_683);
nor U774 (N_774,In_233,In_871);
nor U775 (N_775,In_1392,In_498);
and U776 (N_776,In_1324,In_118);
nor U777 (N_777,In_1190,In_718);
or U778 (N_778,In_745,In_1192);
or U779 (N_779,In_862,In_1053);
or U780 (N_780,In_526,In_1493);
or U781 (N_781,In_1271,In_528);
xor U782 (N_782,In_1097,In_25);
and U783 (N_783,In_932,In_9);
nand U784 (N_784,In_24,In_1263);
and U785 (N_785,In_813,In_5);
xor U786 (N_786,In_1401,In_675);
and U787 (N_787,In_924,In_481);
or U788 (N_788,In_280,In_1062);
or U789 (N_789,In_1180,In_168);
or U790 (N_790,In_1327,In_63);
and U791 (N_791,In_955,In_512);
nor U792 (N_792,In_1147,In_1380);
nor U793 (N_793,In_1289,In_859);
or U794 (N_794,In_325,In_1138);
nand U795 (N_795,In_1489,In_1319);
or U796 (N_796,In_1417,In_73);
or U797 (N_797,In_279,In_5);
nand U798 (N_798,In_408,In_346);
or U799 (N_799,In_340,In_1032);
nand U800 (N_800,In_1320,In_833);
nand U801 (N_801,In_626,In_1122);
or U802 (N_802,In_714,In_149);
nand U803 (N_803,In_1407,In_1259);
and U804 (N_804,In_1194,In_432);
and U805 (N_805,In_115,In_1259);
nor U806 (N_806,In_1150,In_92);
nor U807 (N_807,In_49,In_1007);
or U808 (N_808,In_1297,In_1089);
or U809 (N_809,In_1445,In_1209);
or U810 (N_810,In_625,In_384);
nor U811 (N_811,In_820,In_799);
or U812 (N_812,In_1229,In_433);
xor U813 (N_813,In_250,In_649);
nor U814 (N_814,In_1289,In_539);
nand U815 (N_815,In_29,In_646);
nand U816 (N_816,In_248,In_209);
or U817 (N_817,In_923,In_428);
and U818 (N_818,In_721,In_245);
nand U819 (N_819,In_538,In_574);
nor U820 (N_820,In_396,In_337);
nand U821 (N_821,In_478,In_961);
or U822 (N_822,In_1388,In_165);
xnor U823 (N_823,In_874,In_779);
nor U824 (N_824,In_1467,In_1409);
or U825 (N_825,In_958,In_1398);
or U826 (N_826,In_1231,In_1488);
nor U827 (N_827,In_148,In_757);
and U828 (N_828,In_1122,In_1408);
nor U829 (N_829,In_854,In_96);
or U830 (N_830,In_82,In_522);
or U831 (N_831,In_1360,In_993);
and U832 (N_832,In_192,In_149);
nand U833 (N_833,In_1026,In_91);
nor U834 (N_834,In_578,In_123);
nand U835 (N_835,In_646,In_450);
or U836 (N_836,In_873,In_329);
and U837 (N_837,In_1332,In_566);
nand U838 (N_838,In_1076,In_751);
nand U839 (N_839,In_590,In_273);
or U840 (N_840,In_1448,In_1407);
nand U841 (N_841,In_151,In_997);
nand U842 (N_842,In_415,In_239);
or U843 (N_843,In_413,In_1477);
and U844 (N_844,In_1433,In_1493);
and U845 (N_845,In_1257,In_270);
nor U846 (N_846,In_156,In_17);
or U847 (N_847,In_1391,In_886);
or U848 (N_848,In_1449,In_156);
and U849 (N_849,In_1253,In_1222);
or U850 (N_850,In_449,In_566);
nor U851 (N_851,In_545,In_683);
nor U852 (N_852,In_724,In_525);
or U853 (N_853,In_666,In_3);
nor U854 (N_854,In_656,In_639);
nand U855 (N_855,In_1208,In_185);
and U856 (N_856,In_115,In_1329);
or U857 (N_857,In_816,In_587);
xor U858 (N_858,In_3,In_388);
nand U859 (N_859,In_775,In_1105);
nand U860 (N_860,In_1026,In_95);
nand U861 (N_861,In_1281,In_0);
and U862 (N_862,In_878,In_43);
or U863 (N_863,In_570,In_1283);
and U864 (N_864,In_743,In_253);
nand U865 (N_865,In_500,In_67);
and U866 (N_866,In_1015,In_965);
and U867 (N_867,In_262,In_1394);
and U868 (N_868,In_948,In_135);
nor U869 (N_869,In_714,In_69);
nor U870 (N_870,In_1207,In_1184);
nor U871 (N_871,In_1236,In_264);
nand U872 (N_872,In_843,In_1013);
nor U873 (N_873,In_387,In_220);
or U874 (N_874,In_999,In_239);
or U875 (N_875,In_1465,In_172);
and U876 (N_876,In_153,In_994);
nor U877 (N_877,In_1493,In_270);
or U878 (N_878,In_985,In_771);
and U879 (N_879,In_1315,In_1053);
and U880 (N_880,In_1107,In_336);
nand U881 (N_881,In_11,In_784);
or U882 (N_882,In_288,In_577);
nand U883 (N_883,In_467,In_595);
and U884 (N_884,In_715,In_144);
or U885 (N_885,In_133,In_556);
and U886 (N_886,In_1274,In_121);
or U887 (N_887,In_753,In_1446);
nand U888 (N_888,In_1252,In_1285);
nand U889 (N_889,In_1236,In_167);
nor U890 (N_890,In_1068,In_1321);
nand U891 (N_891,In_607,In_1361);
nand U892 (N_892,In_1452,In_1481);
nand U893 (N_893,In_230,In_1230);
nand U894 (N_894,In_326,In_123);
or U895 (N_895,In_381,In_150);
nor U896 (N_896,In_922,In_937);
nand U897 (N_897,In_119,In_1366);
or U898 (N_898,In_987,In_202);
and U899 (N_899,In_317,In_721);
nand U900 (N_900,In_891,In_1234);
nand U901 (N_901,In_761,In_257);
or U902 (N_902,In_965,In_1285);
nand U903 (N_903,In_381,In_246);
nor U904 (N_904,In_914,In_555);
or U905 (N_905,In_311,In_638);
and U906 (N_906,In_1137,In_1363);
and U907 (N_907,In_762,In_195);
nor U908 (N_908,In_231,In_1458);
and U909 (N_909,In_0,In_888);
nand U910 (N_910,In_1369,In_1291);
and U911 (N_911,In_478,In_881);
nor U912 (N_912,In_1186,In_433);
or U913 (N_913,In_884,In_892);
and U914 (N_914,In_799,In_1200);
and U915 (N_915,In_144,In_478);
and U916 (N_916,In_1224,In_219);
and U917 (N_917,In_1265,In_1405);
nor U918 (N_918,In_376,In_691);
or U919 (N_919,In_42,In_834);
nor U920 (N_920,In_981,In_240);
and U921 (N_921,In_361,In_801);
nor U922 (N_922,In_1011,In_991);
nand U923 (N_923,In_1101,In_836);
xnor U924 (N_924,In_622,In_541);
or U925 (N_925,In_1389,In_177);
and U926 (N_926,In_86,In_605);
xor U927 (N_927,In_1345,In_1417);
nor U928 (N_928,In_1008,In_1336);
and U929 (N_929,In_1362,In_1182);
nor U930 (N_930,In_917,In_1491);
nand U931 (N_931,In_1383,In_124);
nor U932 (N_932,In_182,In_339);
nor U933 (N_933,In_10,In_1299);
nor U934 (N_934,In_640,In_1255);
nor U935 (N_935,In_389,In_853);
nor U936 (N_936,In_1186,In_445);
nand U937 (N_937,In_866,In_501);
nand U938 (N_938,In_945,In_98);
nor U939 (N_939,In_93,In_1125);
or U940 (N_940,In_1282,In_563);
nor U941 (N_941,In_373,In_151);
nand U942 (N_942,In_1354,In_1027);
or U943 (N_943,In_891,In_444);
nand U944 (N_944,In_1369,In_680);
and U945 (N_945,In_1198,In_296);
nand U946 (N_946,In_476,In_735);
or U947 (N_947,In_146,In_852);
or U948 (N_948,In_1154,In_545);
or U949 (N_949,In_1390,In_1371);
nand U950 (N_950,In_647,In_382);
and U951 (N_951,In_14,In_1302);
and U952 (N_952,In_875,In_232);
nand U953 (N_953,In_1370,In_904);
nand U954 (N_954,In_323,In_528);
xnor U955 (N_955,In_963,In_41);
or U956 (N_956,In_1301,In_114);
and U957 (N_957,In_1339,In_776);
or U958 (N_958,In_690,In_792);
or U959 (N_959,In_1103,In_501);
and U960 (N_960,In_1190,In_313);
or U961 (N_961,In_783,In_227);
and U962 (N_962,In_234,In_1469);
or U963 (N_963,In_1476,In_1096);
or U964 (N_964,In_1360,In_796);
and U965 (N_965,In_1466,In_1369);
nor U966 (N_966,In_1352,In_852);
nand U967 (N_967,In_1271,In_195);
or U968 (N_968,In_916,In_1093);
nor U969 (N_969,In_1026,In_585);
nand U970 (N_970,In_896,In_509);
or U971 (N_971,In_1272,In_1028);
and U972 (N_972,In_224,In_1211);
or U973 (N_973,In_510,In_1093);
nor U974 (N_974,In_128,In_1284);
and U975 (N_975,In_1123,In_175);
nor U976 (N_976,In_97,In_82);
nand U977 (N_977,In_426,In_772);
nand U978 (N_978,In_275,In_954);
nand U979 (N_979,In_110,In_1051);
or U980 (N_980,In_285,In_1360);
and U981 (N_981,In_685,In_11);
nand U982 (N_982,In_474,In_30);
and U983 (N_983,In_150,In_630);
and U984 (N_984,In_53,In_202);
or U985 (N_985,In_826,In_1493);
nand U986 (N_986,In_428,In_371);
nand U987 (N_987,In_70,In_894);
nand U988 (N_988,In_1142,In_1467);
and U989 (N_989,In_1071,In_349);
nor U990 (N_990,In_1486,In_230);
nor U991 (N_991,In_553,In_952);
or U992 (N_992,In_23,In_58);
nor U993 (N_993,In_293,In_139);
nor U994 (N_994,In_1191,In_1208);
or U995 (N_995,In_548,In_155);
or U996 (N_996,In_974,In_1369);
or U997 (N_997,In_161,In_490);
and U998 (N_998,In_389,In_476);
nor U999 (N_999,In_435,In_1396);
nor U1000 (N_1000,In_559,In_614);
or U1001 (N_1001,In_189,In_317);
nand U1002 (N_1002,In_475,In_211);
or U1003 (N_1003,In_371,In_95);
nor U1004 (N_1004,In_268,In_1184);
nor U1005 (N_1005,In_1486,In_1125);
and U1006 (N_1006,In_1201,In_786);
nor U1007 (N_1007,In_1018,In_1102);
and U1008 (N_1008,In_962,In_665);
and U1009 (N_1009,In_1285,In_1455);
nor U1010 (N_1010,In_32,In_1183);
nand U1011 (N_1011,In_570,In_242);
or U1012 (N_1012,In_555,In_887);
or U1013 (N_1013,In_253,In_1171);
nor U1014 (N_1014,In_71,In_1246);
or U1015 (N_1015,In_457,In_1224);
and U1016 (N_1016,In_702,In_1271);
or U1017 (N_1017,In_1162,In_653);
nand U1018 (N_1018,In_715,In_516);
nor U1019 (N_1019,In_1,In_52);
nor U1020 (N_1020,In_305,In_1381);
nor U1021 (N_1021,In_253,In_173);
and U1022 (N_1022,In_1001,In_433);
or U1023 (N_1023,In_1254,In_925);
or U1024 (N_1024,In_647,In_999);
nor U1025 (N_1025,In_557,In_728);
or U1026 (N_1026,In_1127,In_746);
and U1027 (N_1027,In_147,In_985);
or U1028 (N_1028,In_975,In_314);
or U1029 (N_1029,In_288,In_219);
nand U1030 (N_1030,In_1422,In_1157);
nand U1031 (N_1031,In_527,In_931);
and U1032 (N_1032,In_54,In_913);
nor U1033 (N_1033,In_87,In_1381);
and U1034 (N_1034,In_1194,In_17);
nor U1035 (N_1035,In_602,In_465);
nor U1036 (N_1036,In_1005,In_1003);
or U1037 (N_1037,In_1324,In_954);
nor U1038 (N_1038,In_782,In_1105);
and U1039 (N_1039,In_142,In_723);
or U1040 (N_1040,In_594,In_495);
or U1041 (N_1041,In_478,In_942);
and U1042 (N_1042,In_1004,In_298);
and U1043 (N_1043,In_767,In_1387);
nand U1044 (N_1044,In_1433,In_1150);
and U1045 (N_1045,In_437,In_77);
or U1046 (N_1046,In_339,In_1327);
and U1047 (N_1047,In_85,In_793);
and U1048 (N_1048,In_1326,In_281);
nand U1049 (N_1049,In_564,In_1437);
or U1050 (N_1050,In_99,In_1403);
and U1051 (N_1051,In_263,In_696);
and U1052 (N_1052,In_1280,In_129);
or U1053 (N_1053,In_690,In_178);
nor U1054 (N_1054,In_238,In_126);
nand U1055 (N_1055,In_832,In_713);
and U1056 (N_1056,In_453,In_543);
or U1057 (N_1057,In_414,In_1407);
and U1058 (N_1058,In_1296,In_598);
nor U1059 (N_1059,In_8,In_361);
nor U1060 (N_1060,In_199,In_603);
nand U1061 (N_1061,In_649,In_776);
or U1062 (N_1062,In_576,In_602);
nor U1063 (N_1063,In_202,In_1329);
or U1064 (N_1064,In_934,In_568);
or U1065 (N_1065,In_1157,In_830);
nand U1066 (N_1066,In_1035,In_1154);
and U1067 (N_1067,In_186,In_1345);
nand U1068 (N_1068,In_209,In_1030);
nand U1069 (N_1069,In_1453,In_743);
nor U1070 (N_1070,In_301,In_1111);
and U1071 (N_1071,In_1283,In_235);
and U1072 (N_1072,In_1254,In_326);
nand U1073 (N_1073,In_484,In_843);
or U1074 (N_1074,In_343,In_1481);
nand U1075 (N_1075,In_1499,In_872);
nor U1076 (N_1076,In_324,In_756);
nor U1077 (N_1077,In_1242,In_1187);
or U1078 (N_1078,In_621,In_384);
or U1079 (N_1079,In_472,In_737);
or U1080 (N_1080,In_805,In_932);
nor U1081 (N_1081,In_37,In_21);
nand U1082 (N_1082,In_893,In_965);
and U1083 (N_1083,In_1052,In_837);
nand U1084 (N_1084,In_550,In_382);
or U1085 (N_1085,In_1470,In_836);
or U1086 (N_1086,In_1403,In_812);
xor U1087 (N_1087,In_49,In_370);
or U1088 (N_1088,In_951,In_1219);
nand U1089 (N_1089,In_576,In_1307);
nand U1090 (N_1090,In_1226,In_198);
nand U1091 (N_1091,In_81,In_777);
nand U1092 (N_1092,In_496,In_704);
or U1093 (N_1093,In_757,In_117);
or U1094 (N_1094,In_1307,In_1329);
and U1095 (N_1095,In_1332,In_87);
and U1096 (N_1096,In_100,In_365);
nor U1097 (N_1097,In_673,In_211);
or U1098 (N_1098,In_1218,In_773);
nor U1099 (N_1099,In_967,In_407);
nand U1100 (N_1100,In_657,In_1420);
nor U1101 (N_1101,In_582,In_1147);
or U1102 (N_1102,In_85,In_1069);
and U1103 (N_1103,In_665,In_1367);
or U1104 (N_1104,In_536,In_115);
and U1105 (N_1105,In_972,In_284);
or U1106 (N_1106,In_1447,In_1405);
and U1107 (N_1107,In_29,In_1264);
or U1108 (N_1108,In_970,In_268);
and U1109 (N_1109,In_714,In_898);
nand U1110 (N_1110,In_74,In_633);
or U1111 (N_1111,In_1068,In_210);
and U1112 (N_1112,In_536,In_978);
and U1113 (N_1113,In_541,In_155);
nor U1114 (N_1114,In_164,In_258);
nand U1115 (N_1115,In_152,In_992);
nand U1116 (N_1116,In_1234,In_441);
and U1117 (N_1117,In_1033,In_165);
and U1118 (N_1118,In_1467,In_90);
nor U1119 (N_1119,In_105,In_1056);
nor U1120 (N_1120,In_747,In_1259);
or U1121 (N_1121,In_1488,In_336);
nand U1122 (N_1122,In_60,In_456);
nor U1123 (N_1123,In_976,In_1438);
nand U1124 (N_1124,In_889,In_315);
nand U1125 (N_1125,In_624,In_1046);
nand U1126 (N_1126,In_1480,In_670);
nor U1127 (N_1127,In_453,In_147);
nor U1128 (N_1128,In_284,In_663);
nand U1129 (N_1129,In_172,In_525);
nand U1130 (N_1130,In_717,In_522);
and U1131 (N_1131,In_1390,In_440);
nor U1132 (N_1132,In_1351,In_1444);
and U1133 (N_1133,In_293,In_128);
nor U1134 (N_1134,In_1257,In_428);
nand U1135 (N_1135,In_1024,In_128);
and U1136 (N_1136,In_501,In_1002);
or U1137 (N_1137,In_742,In_135);
nand U1138 (N_1138,In_431,In_936);
and U1139 (N_1139,In_225,In_610);
xor U1140 (N_1140,In_722,In_1243);
nor U1141 (N_1141,In_43,In_378);
or U1142 (N_1142,In_1036,In_91);
and U1143 (N_1143,In_1467,In_479);
nand U1144 (N_1144,In_85,In_168);
or U1145 (N_1145,In_485,In_167);
and U1146 (N_1146,In_1033,In_491);
and U1147 (N_1147,In_1123,In_1143);
and U1148 (N_1148,In_1030,In_1092);
nor U1149 (N_1149,In_1038,In_1137);
nand U1150 (N_1150,In_395,In_598);
nand U1151 (N_1151,In_206,In_1483);
and U1152 (N_1152,In_252,In_132);
or U1153 (N_1153,In_457,In_1230);
and U1154 (N_1154,In_219,In_1206);
nor U1155 (N_1155,In_767,In_753);
nor U1156 (N_1156,In_155,In_1199);
nor U1157 (N_1157,In_23,In_1018);
or U1158 (N_1158,In_1036,In_1169);
nor U1159 (N_1159,In_482,In_1125);
nor U1160 (N_1160,In_1087,In_1231);
or U1161 (N_1161,In_1030,In_68);
and U1162 (N_1162,In_1354,In_1000);
and U1163 (N_1163,In_1263,In_382);
xnor U1164 (N_1164,In_791,In_545);
or U1165 (N_1165,In_36,In_654);
nand U1166 (N_1166,In_618,In_1032);
nand U1167 (N_1167,In_1433,In_107);
and U1168 (N_1168,In_1261,In_999);
and U1169 (N_1169,In_410,In_960);
and U1170 (N_1170,In_705,In_233);
and U1171 (N_1171,In_849,In_1244);
nand U1172 (N_1172,In_1371,In_1243);
nand U1173 (N_1173,In_244,In_711);
nand U1174 (N_1174,In_1104,In_1212);
nand U1175 (N_1175,In_323,In_109);
and U1176 (N_1176,In_800,In_261);
nor U1177 (N_1177,In_1451,In_1046);
nand U1178 (N_1178,In_81,In_417);
and U1179 (N_1179,In_1268,In_619);
nor U1180 (N_1180,In_12,In_376);
nor U1181 (N_1181,In_973,In_497);
nand U1182 (N_1182,In_885,In_461);
nand U1183 (N_1183,In_753,In_1090);
nand U1184 (N_1184,In_1425,In_543);
or U1185 (N_1185,In_531,In_181);
or U1186 (N_1186,In_808,In_186);
nor U1187 (N_1187,In_51,In_320);
and U1188 (N_1188,In_1162,In_204);
nor U1189 (N_1189,In_859,In_986);
and U1190 (N_1190,In_1200,In_405);
nor U1191 (N_1191,In_500,In_489);
or U1192 (N_1192,In_24,In_187);
or U1193 (N_1193,In_1194,In_1152);
nand U1194 (N_1194,In_935,In_1370);
nand U1195 (N_1195,In_536,In_1492);
and U1196 (N_1196,In_668,In_1283);
or U1197 (N_1197,In_62,In_1029);
nand U1198 (N_1198,In_792,In_591);
and U1199 (N_1199,In_1217,In_1277);
or U1200 (N_1200,In_1037,In_789);
nand U1201 (N_1201,In_56,In_450);
nor U1202 (N_1202,In_227,In_47);
and U1203 (N_1203,In_1076,In_666);
or U1204 (N_1204,In_1184,In_706);
nor U1205 (N_1205,In_1357,In_765);
and U1206 (N_1206,In_1140,In_27);
and U1207 (N_1207,In_1279,In_1294);
nand U1208 (N_1208,In_1192,In_881);
and U1209 (N_1209,In_710,In_684);
nand U1210 (N_1210,In_1100,In_1053);
or U1211 (N_1211,In_191,In_1396);
and U1212 (N_1212,In_1431,In_1256);
or U1213 (N_1213,In_416,In_989);
nor U1214 (N_1214,In_1206,In_1205);
nor U1215 (N_1215,In_472,In_745);
or U1216 (N_1216,In_982,In_577);
and U1217 (N_1217,In_180,In_100);
and U1218 (N_1218,In_13,In_1224);
nor U1219 (N_1219,In_273,In_1114);
and U1220 (N_1220,In_561,In_744);
and U1221 (N_1221,In_1164,In_114);
nor U1222 (N_1222,In_640,In_122);
nand U1223 (N_1223,In_454,In_706);
and U1224 (N_1224,In_781,In_274);
nand U1225 (N_1225,In_1163,In_1248);
nor U1226 (N_1226,In_1364,In_1161);
nor U1227 (N_1227,In_776,In_317);
or U1228 (N_1228,In_78,In_788);
or U1229 (N_1229,In_1118,In_415);
nand U1230 (N_1230,In_985,In_1457);
or U1231 (N_1231,In_389,In_1012);
and U1232 (N_1232,In_1326,In_45);
and U1233 (N_1233,In_244,In_1417);
or U1234 (N_1234,In_82,In_1226);
nor U1235 (N_1235,In_1382,In_1232);
and U1236 (N_1236,In_556,In_180);
or U1237 (N_1237,In_643,In_538);
nor U1238 (N_1238,In_1172,In_1315);
or U1239 (N_1239,In_641,In_486);
nor U1240 (N_1240,In_1342,In_1432);
or U1241 (N_1241,In_1204,In_923);
and U1242 (N_1242,In_451,In_712);
and U1243 (N_1243,In_1088,In_342);
nand U1244 (N_1244,In_141,In_498);
nor U1245 (N_1245,In_773,In_222);
and U1246 (N_1246,In_1063,In_744);
nand U1247 (N_1247,In_532,In_34);
and U1248 (N_1248,In_213,In_1340);
nor U1249 (N_1249,In_553,In_1414);
nor U1250 (N_1250,In_915,In_1346);
or U1251 (N_1251,In_656,In_914);
or U1252 (N_1252,In_1171,In_920);
nand U1253 (N_1253,In_1469,In_231);
nand U1254 (N_1254,In_611,In_680);
nand U1255 (N_1255,In_140,In_123);
nand U1256 (N_1256,In_401,In_1216);
nand U1257 (N_1257,In_944,In_1043);
or U1258 (N_1258,In_1358,In_1497);
nand U1259 (N_1259,In_1288,In_948);
nand U1260 (N_1260,In_223,In_1187);
nor U1261 (N_1261,In_15,In_870);
nand U1262 (N_1262,In_993,In_665);
nand U1263 (N_1263,In_1261,In_581);
nor U1264 (N_1264,In_684,In_488);
and U1265 (N_1265,In_413,In_695);
and U1266 (N_1266,In_1014,In_168);
nor U1267 (N_1267,In_601,In_1327);
nor U1268 (N_1268,In_738,In_965);
and U1269 (N_1269,In_1273,In_1429);
and U1270 (N_1270,In_207,In_836);
and U1271 (N_1271,In_1170,In_971);
or U1272 (N_1272,In_877,In_1067);
and U1273 (N_1273,In_9,In_222);
nand U1274 (N_1274,In_274,In_1488);
and U1275 (N_1275,In_1108,In_984);
and U1276 (N_1276,In_846,In_457);
nor U1277 (N_1277,In_791,In_59);
and U1278 (N_1278,In_868,In_354);
and U1279 (N_1279,In_1253,In_44);
nor U1280 (N_1280,In_1176,In_322);
or U1281 (N_1281,In_24,In_1235);
or U1282 (N_1282,In_1053,In_980);
nand U1283 (N_1283,In_1254,In_455);
xor U1284 (N_1284,In_1423,In_1254);
or U1285 (N_1285,In_1360,In_432);
and U1286 (N_1286,In_489,In_1185);
and U1287 (N_1287,In_531,In_506);
nand U1288 (N_1288,In_1032,In_1474);
nand U1289 (N_1289,In_198,In_813);
and U1290 (N_1290,In_1470,In_1405);
and U1291 (N_1291,In_316,In_544);
nor U1292 (N_1292,In_278,In_137);
or U1293 (N_1293,In_433,In_1028);
nand U1294 (N_1294,In_771,In_544);
nor U1295 (N_1295,In_1220,In_157);
and U1296 (N_1296,In_1141,In_1386);
or U1297 (N_1297,In_946,In_1160);
or U1298 (N_1298,In_1082,In_841);
nor U1299 (N_1299,In_82,In_445);
nor U1300 (N_1300,In_546,In_572);
or U1301 (N_1301,In_8,In_510);
and U1302 (N_1302,In_93,In_1402);
or U1303 (N_1303,In_809,In_770);
and U1304 (N_1304,In_1469,In_15);
and U1305 (N_1305,In_1283,In_491);
and U1306 (N_1306,In_1348,In_330);
or U1307 (N_1307,In_273,In_434);
and U1308 (N_1308,In_1332,In_1112);
and U1309 (N_1309,In_1277,In_62);
or U1310 (N_1310,In_571,In_729);
nor U1311 (N_1311,In_1347,In_169);
and U1312 (N_1312,In_703,In_670);
or U1313 (N_1313,In_708,In_1109);
nand U1314 (N_1314,In_1492,In_182);
and U1315 (N_1315,In_652,In_367);
and U1316 (N_1316,In_17,In_25);
nand U1317 (N_1317,In_1443,In_449);
and U1318 (N_1318,In_1079,In_403);
and U1319 (N_1319,In_127,In_525);
and U1320 (N_1320,In_1139,In_1412);
or U1321 (N_1321,In_674,In_785);
or U1322 (N_1322,In_1241,In_1494);
and U1323 (N_1323,In_1331,In_458);
nor U1324 (N_1324,In_1369,In_1301);
nand U1325 (N_1325,In_1089,In_855);
or U1326 (N_1326,In_736,In_562);
or U1327 (N_1327,In_792,In_484);
xor U1328 (N_1328,In_237,In_1248);
and U1329 (N_1329,In_1275,In_760);
nor U1330 (N_1330,In_325,In_399);
nand U1331 (N_1331,In_1188,In_1058);
and U1332 (N_1332,In_323,In_814);
nand U1333 (N_1333,In_390,In_1027);
or U1334 (N_1334,In_435,In_344);
and U1335 (N_1335,In_938,In_1404);
nor U1336 (N_1336,In_105,In_4);
and U1337 (N_1337,In_467,In_37);
and U1338 (N_1338,In_434,In_1255);
and U1339 (N_1339,In_392,In_1089);
and U1340 (N_1340,In_239,In_1258);
nand U1341 (N_1341,In_925,In_198);
xnor U1342 (N_1342,In_349,In_276);
nand U1343 (N_1343,In_1371,In_609);
or U1344 (N_1344,In_756,In_100);
or U1345 (N_1345,In_673,In_771);
nand U1346 (N_1346,In_984,In_1420);
nor U1347 (N_1347,In_1111,In_1102);
and U1348 (N_1348,In_1229,In_846);
nor U1349 (N_1349,In_686,In_25);
xor U1350 (N_1350,In_1281,In_938);
and U1351 (N_1351,In_1289,In_402);
and U1352 (N_1352,In_840,In_682);
or U1353 (N_1353,In_351,In_621);
nand U1354 (N_1354,In_1377,In_462);
nand U1355 (N_1355,In_548,In_1191);
or U1356 (N_1356,In_1417,In_1147);
and U1357 (N_1357,In_769,In_581);
or U1358 (N_1358,In_937,In_300);
nor U1359 (N_1359,In_377,In_994);
and U1360 (N_1360,In_1158,In_364);
nor U1361 (N_1361,In_1075,In_638);
or U1362 (N_1362,In_1495,In_747);
nand U1363 (N_1363,In_846,In_1193);
and U1364 (N_1364,In_32,In_1468);
or U1365 (N_1365,In_625,In_1069);
nand U1366 (N_1366,In_1094,In_827);
nand U1367 (N_1367,In_305,In_52);
or U1368 (N_1368,In_989,In_417);
or U1369 (N_1369,In_160,In_1064);
nand U1370 (N_1370,In_792,In_1475);
nor U1371 (N_1371,In_1297,In_1332);
and U1372 (N_1372,In_675,In_876);
nor U1373 (N_1373,In_1320,In_361);
nor U1374 (N_1374,In_62,In_1207);
and U1375 (N_1375,In_201,In_598);
and U1376 (N_1376,In_1472,In_123);
or U1377 (N_1377,In_1311,In_463);
or U1378 (N_1378,In_216,In_538);
or U1379 (N_1379,In_163,In_1080);
nand U1380 (N_1380,In_151,In_841);
nand U1381 (N_1381,In_989,In_1175);
and U1382 (N_1382,In_1379,In_657);
nor U1383 (N_1383,In_761,In_118);
and U1384 (N_1384,In_598,In_1493);
nand U1385 (N_1385,In_357,In_476);
nand U1386 (N_1386,In_734,In_374);
and U1387 (N_1387,In_946,In_991);
or U1388 (N_1388,In_862,In_496);
and U1389 (N_1389,In_997,In_866);
and U1390 (N_1390,In_1470,In_718);
nor U1391 (N_1391,In_1262,In_476);
nor U1392 (N_1392,In_717,In_366);
nor U1393 (N_1393,In_1328,In_313);
and U1394 (N_1394,In_688,In_255);
or U1395 (N_1395,In_819,In_1196);
or U1396 (N_1396,In_61,In_989);
nand U1397 (N_1397,In_1390,In_61);
nor U1398 (N_1398,In_449,In_1156);
nand U1399 (N_1399,In_1113,In_698);
or U1400 (N_1400,In_689,In_52);
or U1401 (N_1401,In_1253,In_1012);
or U1402 (N_1402,In_1405,In_84);
or U1403 (N_1403,In_195,In_1238);
nor U1404 (N_1404,In_1351,In_244);
nand U1405 (N_1405,In_1194,In_1301);
and U1406 (N_1406,In_60,In_39);
nand U1407 (N_1407,In_853,In_1032);
or U1408 (N_1408,In_1052,In_25);
or U1409 (N_1409,In_1084,In_1081);
nor U1410 (N_1410,In_883,In_742);
and U1411 (N_1411,In_1306,In_1177);
nor U1412 (N_1412,In_810,In_1463);
nor U1413 (N_1413,In_649,In_301);
or U1414 (N_1414,In_743,In_1181);
nor U1415 (N_1415,In_1389,In_1496);
or U1416 (N_1416,In_493,In_885);
and U1417 (N_1417,In_1472,In_714);
and U1418 (N_1418,In_791,In_591);
or U1419 (N_1419,In_1143,In_790);
nand U1420 (N_1420,In_781,In_25);
or U1421 (N_1421,In_700,In_851);
and U1422 (N_1422,In_705,In_1398);
nor U1423 (N_1423,In_902,In_1050);
nor U1424 (N_1424,In_1230,In_1046);
nor U1425 (N_1425,In_999,In_1407);
and U1426 (N_1426,In_1407,In_106);
nor U1427 (N_1427,In_699,In_1145);
and U1428 (N_1428,In_1012,In_1);
nand U1429 (N_1429,In_1405,In_694);
nand U1430 (N_1430,In_1419,In_1382);
nand U1431 (N_1431,In_707,In_747);
nand U1432 (N_1432,In_544,In_970);
and U1433 (N_1433,In_192,In_1053);
nor U1434 (N_1434,In_121,In_68);
nand U1435 (N_1435,In_1090,In_1441);
nand U1436 (N_1436,In_642,In_499);
and U1437 (N_1437,In_576,In_1025);
nand U1438 (N_1438,In_414,In_1228);
and U1439 (N_1439,In_205,In_301);
nand U1440 (N_1440,In_1157,In_545);
nand U1441 (N_1441,In_1370,In_1251);
or U1442 (N_1442,In_480,In_1416);
or U1443 (N_1443,In_393,In_1497);
nor U1444 (N_1444,In_1,In_467);
or U1445 (N_1445,In_1036,In_1143);
nor U1446 (N_1446,In_1342,In_870);
nand U1447 (N_1447,In_553,In_865);
or U1448 (N_1448,In_504,In_1408);
nand U1449 (N_1449,In_503,In_1260);
nor U1450 (N_1450,In_900,In_271);
or U1451 (N_1451,In_1018,In_575);
nor U1452 (N_1452,In_1311,In_877);
and U1453 (N_1453,In_1042,In_31);
nor U1454 (N_1454,In_770,In_1306);
and U1455 (N_1455,In_672,In_1474);
nand U1456 (N_1456,In_33,In_732);
or U1457 (N_1457,In_123,In_352);
nor U1458 (N_1458,In_1206,In_615);
nor U1459 (N_1459,In_814,In_33);
or U1460 (N_1460,In_315,In_748);
and U1461 (N_1461,In_385,In_893);
and U1462 (N_1462,In_665,In_212);
nand U1463 (N_1463,In_1322,In_1063);
nor U1464 (N_1464,In_1174,In_1090);
nor U1465 (N_1465,In_1379,In_114);
nor U1466 (N_1466,In_109,In_95);
or U1467 (N_1467,In_129,In_961);
or U1468 (N_1468,In_209,In_964);
nand U1469 (N_1469,In_798,In_906);
nor U1470 (N_1470,In_1325,In_381);
nor U1471 (N_1471,In_297,In_90);
nor U1472 (N_1472,In_1354,In_1193);
or U1473 (N_1473,In_1361,In_183);
nand U1474 (N_1474,In_173,In_79);
or U1475 (N_1475,In_826,In_562);
and U1476 (N_1476,In_83,In_527);
nand U1477 (N_1477,In_368,In_74);
nand U1478 (N_1478,In_95,In_1347);
and U1479 (N_1479,In_1203,In_544);
nand U1480 (N_1480,In_1284,In_180);
nand U1481 (N_1481,In_861,In_1143);
or U1482 (N_1482,In_313,In_1137);
nand U1483 (N_1483,In_222,In_1040);
or U1484 (N_1484,In_675,In_1104);
nand U1485 (N_1485,In_1459,In_757);
nand U1486 (N_1486,In_788,In_124);
and U1487 (N_1487,In_646,In_1329);
or U1488 (N_1488,In_988,In_76);
or U1489 (N_1489,In_1164,In_877);
nand U1490 (N_1490,In_1472,In_1090);
and U1491 (N_1491,In_513,In_1257);
nand U1492 (N_1492,In_197,In_208);
or U1493 (N_1493,In_1010,In_540);
nand U1494 (N_1494,In_224,In_509);
and U1495 (N_1495,In_1308,In_167);
nor U1496 (N_1496,In_1111,In_445);
and U1497 (N_1497,In_1166,In_1496);
or U1498 (N_1498,In_1126,In_440);
nor U1499 (N_1499,In_1063,In_460);
and U1500 (N_1500,In_344,In_389);
nor U1501 (N_1501,In_1450,In_541);
nor U1502 (N_1502,In_869,In_1250);
xor U1503 (N_1503,In_1215,In_98);
or U1504 (N_1504,In_39,In_393);
and U1505 (N_1505,In_624,In_1251);
nand U1506 (N_1506,In_1109,In_412);
or U1507 (N_1507,In_540,In_951);
and U1508 (N_1508,In_487,In_276);
and U1509 (N_1509,In_1484,In_267);
and U1510 (N_1510,In_1001,In_659);
or U1511 (N_1511,In_1142,In_645);
xnor U1512 (N_1512,In_468,In_776);
and U1513 (N_1513,In_188,In_1145);
or U1514 (N_1514,In_670,In_784);
or U1515 (N_1515,In_1081,In_1191);
or U1516 (N_1516,In_954,In_391);
and U1517 (N_1517,In_153,In_174);
xor U1518 (N_1518,In_1229,In_1419);
or U1519 (N_1519,In_1169,In_131);
nor U1520 (N_1520,In_911,In_662);
or U1521 (N_1521,In_547,In_1372);
nor U1522 (N_1522,In_1275,In_559);
or U1523 (N_1523,In_277,In_34);
and U1524 (N_1524,In_1292,In_503);
nand U1525 (N_1525,In_1331,In_822);
nand U1526 (N_1526,In_989,In_947);
or U1527 (N_1527,In_532,In_403);
nor U1528 (N_1528,In_716,In_1457);
or U1529 (N_1529,In_1050,In_204);
or U1530 (N_1530,In_16,In_86);
and U1531 (N_1531,In_1384,In_259);
nand U1532 (N_1532,In_1336,In_1208);
nand U1533 (N_1533,In_797,In_231);
or U1534 (N_1534,In_291,In_592);
nand U1535 (N_1535,In_965,In_253);
nor U1536 (N_1536,In_1276,In_1200);
nor U1537 (N_1537,In_1400,In_1401);
nand U1538 (N_1538,In_847,In_1326);
nor U1539 (N_1539,In_268,In_256);
nand U1540 (N_1540,In_74,In_991);
nor U1541 (N_1541,In_637,In_1475);
or U1542 (N_1542,In_1474,In_629);
nor U1543 (N_1543,In_1081,In_1033);
nor U1544 (N_1544,In_1355,In_901);
and U1545 (N_1545,In_332,In_1476);
or U1546 (N_1546,In_1273,In_1319);
or U1547 (N_1547,In_445,In_835);
or U1548 (N_1548,In_677,In_1169);
nand U1549 (N_1549,In_1452,In_758);
nor U1550 (N_1550,In_1036,In_990);
nand U1551 (N_1551,In_603,In_106);
nor U1552 (N_1552,In_744,In_112);
nor U1553 (N_1553,In_1307,In_1081);
nor U1554 (N_1554,In_247,In_510);
nand U1555 (N_1555,In_558,In_480);
nor U1556 (N_1556,In_378,In_827);
or U1557 (N_1557,In_688,In_1487);
and U1558 (N_1558,In_279,In_227);
and U1559 (N_1559,In_445,In_821);
nand U1560 (N_1560,In_822,In_934);
and U1561 (N_1561,In_241,In_1128);
nor U1562 (N_1562,In_614,In_1331);
or U1563 (N_1563,In_926,In_727);
or U1564 (N_1564,In_249,In_1420);
nand U1565 (N_1565,In_1455,In_778);
nor U1566 (N_1566,In_660,In_467);
or U1567 (N_1567,In_1482,In_50);
nor U1568 (N_1568,In_467,In_522);
nand U1569 (N_1569,In_501,In_520);
nand U1570 (N_1570,In_1245,In_38);
or U1571 (N_1571,In_1400,In_167);
or U1572 (N_1572,In_307,In_918);
nor U1573 (N_1573,In_927,In_31);
and U1574 (N_1574,In_640,In_701);
and U1575 (N_1575,In_987,In_1343);
nor U1576 (N_1576,In_1489,In_1468);
or U1577 (N_1577,In_589,In_1188);
or U1578 (N_1578,In_400,In_1393);
nor U1579 (N_1579,In_440,In_411);
or U1580 (N_1580,In_55,In_345);
or U1581 (N_1581,In_310,In_176);
nor U1582 (N_1582,In_171,In_1151);
or U1583 (N_1583,In_514,In_1076);
nand U1584 (N_1584,In_617,In_73);
nand U1585 (N_1585,In_948,In_1408);
or U1586 (N_1586,In_148,In_1401);
or U1587 (N_1587,In_951,In_1308);
nand U1588 (N_1588,In_46,In_983);
or U1589 (N_1589,In_360,In_635);
nand U1590 (N_1590,In_339,In_246);
and U1591 (N_1591,In_524,In_487);
or U1592 (N_1592,In_1319,In_1053);
and U1593 (N_1593,In_642,In_1435);
nor U1594 (N_1594,In_1268,In_394);
or U1595 (N_1595,In_1060,In_485);
nor U1596 (N_1596,In_1190,In_685);
or U1597 (N_1597,In_1463,In_133);
nand U1598 (N_1598,In_1483,In_115);
nor U1599 (N_1599,In_1146,In_431);
or U1600 (N_1600,In_1070,In_947);
nor U1601 (N_1601,In_20,In_1384);
nor U1602 (N_1602,In_1231,In_539);
nor U1603 (N_1603,In_827,In_528);
and U1604 (N_1604,In_1170,In_746);
nand U1605 (N_1605,In_152,In_1091);
or U1606 (N_1606,In_562,In_929);
and U1607 (N_1607,In_1187,In_945);
and U1608 (N_1608,In_1171,In_1075);
and U1609 (N_1609,In_1011,In_385);
nor U1610 (N_1610,In_321,In_218);
and U1611 (N_1611,In_47,In_712);
nand U1612 (N_1612,In_1457,In_523);
nand U1613 (N_1613,In_212,In_318);
nand U1614 (N_1614,In_1167,In_730);
nand U1615 (N_1615,In_1175,In_901);
nand U1616 (N_1616,In_692,In_504);
and U1617 (N_1617,In_1146,In_161);
and U1618 (N_1618,In_1347,In_133);
nor U1619 (N_1619,In_21,In_107);
or U1620 (N_1620,In_526,In_247);
nor U1621 (N_1621,In_1291,In_1371);
nor U1622 (N_1622,In_174,In_126);
and U1623 (N_1623,In_1190,In_294);
nor U1624 (N_1624,In_394,In_1299);
nor U1625 (N_1625,In_472,In_1124);
and U1626 (N_1626,In_182,In_1451);
nand U1627 (N_1627,In_94,In_534);
or U1628 (N_1628,In_434,In_418);
nand U1629 (N_1629,In_230,In_1213);
and U1630 (N_1630,In_82,In_1210);
nor U1631 (N_1631,In_1134,In_1463);
or U1632 (N_1632,In_178,In_1086);
nor U1633 (N_1633,In_247,In_1443);
or U1634 (N_1634,In_388,In_69);
and U1635 (N_1635,In_456,In_1069);
nor U1636 (N_1636,In_554,In_1120);
and U1637 (N_1637,In_492,In_1190);
and U1638 (N_1638,In_325,In_573);
nor U1639 (N_1639,In_1292,In_1154);
nor U1640 (N_1640,In_11,In_1288);
or U1641 (N_1641,In_851,In_462);
nand U1642 (N_1642,In_917,In_65);
or U1643 (N_1643,In_1254,In_1493);
or U1644 (N_1644,In_316,In_1018);
or U1645 (N_1645,In_1201,In_43);
nand U1646 (N_1646,In_70,In_1451);
nand U1647 (N_1647,In_1273,In_339);
nor U1648 (N_1648,In_804,In_584);
nor U1649 (N_1649,In_1038,In_1023);
nand U1650 (N_1650,In_560,In_1354);
or U1651 (N_1651,In_1142,In_940);
nand U1652 (N_1652,In_95,In_551);
or U1653 (N_1653,In_605,In_618);
nand U1654 (N_1654,In_1056,In_299);
or U1655 (N_1655,In_873,In_952);
nor U1656 (N_1656,In_97,In_721);
and U1657 (N_1657,In_717,In_837);
nor U1658 (N_1658,In_1196,In_1322);
nor U1659 (N_1659,In_68,In_40);
nand U1660 (N_1660,In_315,In_1030);
and U1661 (N_1661,In_830,In_474);
nor U1662 (N_1662,In_640,In_1258);
nand U1663 (N_1663,In_664,In_39);
nand U1664 (N_1664,In_1379,In_41);
or U1665 (N_1665,In_1473,In_17);
or U1666 (N_1666,In_515,In_100);
nor U1667 (N_1667,In_1276,In_308);
nor U1668 (N_1668,In_101,In_1477);
nand U1669 (N_1669,In_1117,In_1307);
and U1670 (N_1670,In_1168,In_701);
and U1671 (N_1671,In_614,In_78);
and U1672 (N_1672,In_957,In_1285);
nand U1673 (N_1673,In_147,In_717);
or U1674 (N_1674,In_167,In_738);
or U1675 (N_1675,In_106,In_19);
nor U1676 (N_1676,In_952,In_1286);
nand U1677 (N_1677,In_1000,In_382);
and U1678 (N_1678,In_1075,In_906);
or U1679 (N_1679,In_1031,In_704);
nor U1680 (N_1680,In_757,In_1020);
and U1681 (N_1681,In_263,In_499);
nor U1682 (N_1682,In_702,In_17);
or U1683 (N_1683,In_529,In_1356);
nor U1684 (N_1684,In_1226,In_604);
nor U1685 (N_1685,In_1118,In_914);
nor U1686 (N_1686,In_1440,In_295);
and U1687 (N_1687,In_1197,In_1305);
or U1688 (N_1688,In_1202,In_478);
and U1689 (N_1689,In_992,In_1268);
and U1690 (N_1690,In_915,In_1015);
and U1691 (N_1691,In_324,In_1124);
or U1692 (N_1692,In_1280,In_1277);
or U1693 (N_1693,In_523,In_431);
nand U1694 (N_1694,In_590,In_527);
and U1695 (N_1695,In_1308,In_1099);
and U1696 (N_1696,In_349,In_1441);
nand U1697 (N_1697,In_130,In_1229);
nor U1698 (N_1698,In_1214,In_501);
nand U1699 (N_1699,In_954,In_1391);
or U1700 (N_1700,In_571,In_1217);
nand U1701 (N_1701,In_1183,In_1388);
nand U1702 (N_1702,In_789,In_781);
xnor U1703 (N_1703,In_39,In_794);
or U1704 (N_1704,In_907,In_413);
nand U1705 (N_1705,In_1004,In_513);
nand U1706 (N_1706,In_586,In_222);
nand U1707 (N_1707,In_1248,In_1037);
or U1708 (N_1708,In_303,In_1209);
and U1709 (N_1709,In_124,In_516);
xor U1710 (N_1710,In_58,In_409);
and U1711 (N_1711,In_890,In_686);
nor U1712 (N_1712,In_298,In_441);
and U1713 (N_1713,In_211,In_655);
or U1714 (N_1714,In_455,In_836);
or U1715 (N_1715,In_851,In_1372);
and U1716 (N_1716,In_573,In_1383);
nand U1717 (N_1717,In_1276,In_21);
nor U1718 (N_1718,In_915,In_374);
and U1719 (N_1719,In_1448,In_900);
nor U1720 (N_1720,In_629,In_923);
nor U1721 (N_1721,In_162,In_701);
nand U1722 (N_1722,In_1380,In_704);
or U1723 (N_1723,In_677,In_236);
nor U1724 (N_1724,In_780,In_736);
or U1725 (N_1725,In_297,In_825);
nand U1726 (N_1726,In_583,In_1313);
or U1727 (N_1727,In_589,In_1250);
xor U1728 (N_1728,In_1151,In_1386);
nand U1729 (N_1729,In_1162,In_1249);
nand U1730 (N_1730,In_769,In_181);
and U1731 (N_1731,In_613,In_379);
nor U1732 (N_1732,In_703,In_829);
nand U1733 (N_1733,In_27,In_836);
nand U1734 (N_1734,In_226,In_348);
nand U1735 (N_1735,In_1234,In_1490);
or U1736 (N_1736,In_61,In_369);
and U1737 (N_1737,In_851,In_154);
or U1738 (N_1738,In_1050,In_470);
nand U1739 (N_1739,In_1050,In_1177);
nor U1740 (N_1740,In_656,In_653);
nor U1741 (N_1741,In_477,In_592);
nor U1742 (N_1742,In_534,In_1080);
or U1743 (N_1743,In_177,In_1008);
and U1744 (N_1744,In_1150,In_277);
nand U1745 (N_1745,In_1082,In_87);
xor U1746 (N_1746,In_940,In_1066);
nand U1747 (N_1747,In_1053,In_41);
nand U1748 (N_1748,In_960,In_548);
nor U1749 (N_1749,In_1155,In_869);
and U1750 (N_1750,In_865,In_698);
and U1751 (N_1751,In_1213,In_847);
and U1752 (N_1752,In_1492,In_1484);
or U1753 (N_1753,In_1496,In_647);
and U1754 (N_1754,In_682,In_1446);
and U1755 (N_1755,In_1032,In_209);
and U1756 (N_1756,In_769,In_917);
and U1757 (N_1757,In_1075,In_1464);
or U1758 (N_1758,In_873,In_523);
or U1759 (N_1759,In_1006,In_517);
xnor U1760 (N_1760,In_1357,In_771);
xor U1761 (N_1761,In_168,In_419);
nor U1762 (N_1762,In_1407,In_1157);
nor U1763 (N_1763,In_918,In_1285);
or U1764 (N_1764,In_953,In_702);
and U1765 (N_1765,In_114,In_898);
nand U1766 (N_1766,In_1354,In_2);
nand U1767 (N_1767,In_1463,In_431);
nor U1768 (N_1768,In_635,In_495);
nand U1769 (N_1769,In_38,In_950);
nand U1770 (N_1770,In_522,In_432);
nand U1771 (N_1771,In_51,In_975);
nor U1772 (N_1772,In_740,In_84);
or U1773 (N_1773,In_1039,In_956);
and U1774 (N_1774,In_442,In_58);
nand U1775 (N_1775,In_1228,In_1451);
nand U1776 (N_1776,In_125,In_1334);
nand U1777 (N_1777,In_260,In_787);
nor U1778 (N_1778,In_907,In_293);
or U1779 (N_1779,In_184,In_682);
nor U1780 (N_1780,In_1090,In_966);
or U1781 (N_1781,In_1410,In_360);
nand U1782 (N_1782,In_544,In_1242);
or U1783 (N_1783,In_1272,In_1451);
and U1784 (N_1784,In_743,In_460);
or U1785 (N_1785,In_661,In_1316);
or U1786 (N_1786,In_448,In_1392);
nand U1787 (N_1787,In_501,In_1277);
nor U1788 (N_1788,In_137,In_1181);
and U1789 (N_1789,In_1032,In_962);
nor U1790 (N_1790,In_204,In_391);
or U1791 (N_1791,In_556,In_212);
and U1792 (N_1792,In_632,In_565);
nor U1793 (N_1793,In_12,In_1050);
and U1794 (N_1794,In_1344,In_654);
nand U1795 (N_1795,In_1455,In_167);
or U1796 (N_1796,In_1326,In_197);
and U1797 (N_1797,In_310,In_1085);
nor U1798 (N_1798,In_408,In_1281);
or U1799 (N_1799,In_909,In_724);
or U1800 (N_1800,In_478,In_518);
and U1801 (N_1801,In_773,In_1117);
and U1802 (N_1802,In_506,In_638);
or U1803 (N_1803,In_501,In_1151);
nor U1804 (N_1804,In_306,In_1251);
and U1805 (N_1805,In_1315,In_184);
nor U1806 (N_1806,In_1412,In_703);
nand U1807 (N_1807,In_1283,In_5);
nor U1808 (N_1808,In_1384,In_1271);
nand U1809 (N_1809,In_655,In_799);
or U1810 (N_1810,In_984,In_337);
or U1811 (N_1811,In_1178,In_1142);
or U1812 (N_1812,In_1245,In_1370);
nor U1813 (N_1813,In_977,In_179);
nand U1814 (N_1814,In_881,In_96);
or U1815 (N_1815,In_685,In_676);
xor U1816 (N_1816,In_574,In_800);
xor U1817 (N_1817,In_44,In_1371);
nor U1818 (N_1818,In_1368,In_1271);
or U1819 (N_1819,In_890,In_1365);
nand U1820 (N_1820,In_1189,In_1322);
or U1821 (N_1821,In_1323,In_800);
nor U1822 (N_1822,In_630,In_1290);
and U1823 (N_1823,In_660,In_1487);
nor U1824 (N_1824,In_1126,In_76);
and U1825 (N_1825,In_1348,In_1411);
and U1826 (N_1826,In_808,In_865);
or U1827 (N_1827,In_774,In_377);
and U1828 (N_1828,In_386,In_403);
nor U1829 (N_1829,In_1312,In_1163);
nand U1830 (N_1830,In_48,In_532);
or U1831 (N_1831,In_753,In_1356);
or U1832 (N_1832,In_1444,In_408);
nor U1833 (N_1833,In_560,In_650);
nor U1834 (N_1834,In_1101,In_1193);
nor U1835 (N_1835,In_1093,In_32);
and U1836 (N_1836,In_978,In_1038);
nor U1837 (N_1837,In_10,In_903);
and U1838 (N_1838,In_676,In_729);
and U1839 (N_1839,In_1281,In_161);
nand U1840 (N_1840,In_1435,In_785);
or U1841 (N_1841,In_84,In_1270);
nor U1842 (N_1842,In_1232,In_1422);
and U1843 (N_1843,In_1384,In_159);
and U1844 (N_1844,In_906,In_1400);
and U1845 (N_1845,In_667,In_190);
or U1846 (N_1846,In_519,In_1312);
or U1847 (N_1847,In_807,In_920);
nor U1848 (N_1848,In_1145,In_205);
or U1849 (N_1849,In_1108,In_1017);
nor U1850 (N_1850,In_691,In_1221);
or U1851 (N_1851,In_1055,In_342);
and U1852 (N_1852,In_806,In_982);
and U1853 (N_1853,In_848,In_1161);
nor U1854 (N_1854,In_969,In_976);
nor U1855 (N_1855,In_286,In_523);
and U1856 (N_1856,In_980,In_1423);
and U1857 (N_1857,In_992,In_1296);
and U1858 (N_1858,In_1104,In_188);
nand U1859 (N_1859,In_1402,In_1343);
and U1860 (N_1860,In_1107,In_461);
and U1861 (N_1861,In_261,In_1170);
or U1862 (N_1862,In_646,In_684);
or U1863 (N_1863,In_1465,In_1046);
and U1864 (N_1864,In_567,In_129);
nand U1865 (N_1865,In_211,In_689);
and U1866 (N_1866,In_1121,In_937);
nor U1867 (N_1867,In_1469,In_229);
nor U1868 (N_1868,In_993,In_920);
and U1869 (N_1869,In_1155,In_1053);
nand U1870 (N_1870,In_592,In_671);
xnor U1871 (N_1871,In_1019,In_1068);
and U1872 (N_1872,In_684,In_504);
nor U1873 (N_1873,In_1493,In_31);
or U1874 (N_1874,In_1320,In_781);
and U1875 (N_1875,In_997,In_308);
nor U1876 (N_1876,In_810,In_1428);
or U1877 (N_1877,In_709,In_970);
and U1878 (N_1878,In_439,In_630);
nand U1879 (N_1879,In_1496,In_1269);
nor U1880 (N_1880,In_728,In_154);
nand U1881 (N_1881,In_1309,In_818);
nand U1882 (N_1882,In_1401,In_452);
and U1883 (N_1883,In_476,In_842);
or U1884 (N_1884,In_1267,In_745);
and U1885 (N_1885,In_377,In_291);
nand U1886 (N_1886,In_943,In_56);
or U1887 (N_1887,In_1143,In_818);
nand U1888 (N_1888,In_706,In_3);
nand U1889 (N_1889,In_756,In_963);
or U1890 (N_1890,In_421,In_799);
nand U1891 (N_1891,In_1428,In_149);
nand U1892 (N_1892,In_1383,In_507);
nand U1893 (N_1893,In_1059,In_245);
nand U1894 (N_1894,In_1036,In_914);
nor U1895 (N_1895,In_1128,In_1058);
nand U1896 (N_1896,In_811,In_1166);
nor U1897 (N_1897,In_837,In_221);
or U1898 (N_1898,In_1332,In_1066);
nor U1899 (N_1899,In_1288,In_406);
and U1900 (N_1900,In_695,In_1452);
nand U1901 (N_1901,In_1383,In_181);
nor U1902 (N_1902,In_730,In_1497);
or U1903 (N_1903,In_943,In_1173);
or U1904 (N_1904,In_756,In_192);
or U1905 (N_1905,In_912,In_999);
and U1906 (N_1906,In_31,In_585);
or U1907 (N_1907,In_988,In_413);
nand U1908 (N_1908,In_884,In_397);
or U1909 (N_1909,In_925,In_842);
nand U1910 (N_1910,In_487,In_1490);
nand U1911 (N_1911,In_12,In_1344);
nand U1912 (N_1912,In_1173,In_1239);
nand U1913 (N_1913,In_1289,In_125);
xor U1914 (N_1914,In_1087,In_533);
and U1915 (N_1915,In_933,In_1429);
nor U1916 (N_1916,In_1221,In_1400);
and U1917 (N_1917,In_1180,In_192);
nand U1918 (N_1918,In_831,In_363);
and U1919 (N_1919,In_1281,In_555);
and U1920 (N_1920,In_1311,In_730);
or U1921 (N_1921,In_134,In_1450);
and U1922 (N_1922,In_662,In_1166);
nand U1923 (N_1923,In_1424,In_1496);
or U1924 (N_1924,In_1412,In_911);
nand U1925 (N_1925,In_1465,In_1445);
or U1926 (N_1926,In_605,In_1310);
and U1927 (N_1927,In_1190,In_549);
nand U1928 (N_1928,In_161,In_574);
nor U1929 (N_1929,In_89,In_1023);
and U1930 (N_1930,In_153,In_1336);
and U1931 (N_1931,In_773,In_680);
or U1932 (N_1932,In_1370,In_803);
or U1933 (N_1933,In_1277,In_375);
nor U1934 (N_1934,In_888,In_163);
and U1935 (N_1935,In_286,In_1393);
or U1936 (N_1936,In_199,In_526);
nor U1937 (N_1937,In_879,In_857);
and U1938 (N_1938,In_921,In_172);
nor U1939 (N_1939,In_160,In_1341);
nand U1940 (N_1940,In_1474,In_392);
nor U1941 (N_1941,In_1264,In_1268);
and U1942 (N_1942,In_1105,In_1241);
and U1943 (N_1943,In_500,In_563);
nand U1944 (N_1944,In_75,In_1428);
and U1945 (N_1945,In_1279,In_399);
or U1946 (N_1946,In_419,In_913);
and U1947 (N_1947,In_173,In_1269);
nor U1948 (N_1948,In_1380,In_956);
nand U1949 (N_1949,In_1181,In_325);
and U1950 (N_1950,In_1352,In_1437);
and U1951 (N_1951,In_933,In_1407);
nand U1952 (N_1952,In_117,In_132);
nand U1953 (N_1953,In_464,In_434);
nor U1954 (N_1954,In_253,In_637);
nand U1955 (N_1955,In_449,In_667);
and U1956 (N_1956,In_993,In_1041);
and U1957 (N_1957,In_827,In_435);
nor U1958 (N_1958,In_323,In_364);
nand U1959 (N_1959,In_1382,In_297);
or U1960 (N_1960,In_378,In_426);
and U1961 (N_1961,In_358,In_846);
and U1962 (N_1962,In_726,In_974);
nor U1963 (N_1963,In_878,In_1463);
nand U1964 (N_1964,In_477,In_739);
nand U1965 (N_1965,In_307,In_867);
and U1966 (N_1966,In_1145,In_174);
or U1967 (N_1967,In_1030,In_1271);
or U1968 (N_1968,In_1391,In_1414);
or U1969 (N_1969,In_1432,In_906);
nand U1970 (N_1970,In_1092,In_1166);
or U1971 (N_1971,In_129,In_1030);
nand U1972 (N_1972,In_152,In_1190);
nor U1973 (N_1973,In_1362,In_1449);
nor U1974 (N_1974,In_1374,In_797);
or U1975 (N_1975,In_16,In_437);
nor U1976 (N_1976,In_754,In_1452);
or U1977 (N_1977,In_757,In_581);
or U1978 (N_1978,In_988,In_65);
nor U1979 (N_1979,In_883,In_546);
and U1980 (N_1980,In_18,In_491);
xor U1981 (N_1981,In_342,In_1278);
nand U1982 (N_1982,In_1086,In_800);
nand U1983 (N_1983,In_453,In_484);
nor U1984 (N_1984,In_62,In_1240);
or U1985 (N_1985,In_785,In_47);
or U1986 (N_1986,In_561,In_47);
and U1987 (N_1987,In_135,In_71);
nor U1988 (N_1988,In_294,In_0);
and U1989 (N_1989,In_1188,In_939);
nand U1990 (N_1990,In_601,In_1334);
and U1991 (N_1991,In_1305,In_280);
and U1992 (N_1992,In_283,In_1284);
or U1993 (N_1993,In_1058,In_490);
nand U1994 (N_1994,In_706,In_1356);
nand U1995 (N_1995,In_1280,In_1235);
or U1996 (N_1996,In_851,In_341);
and U1997 (N_1997,In_82,In_1318);
nor U1998 (N_1998,In_76,In_2);
nor U1999 (N_1999,In_1148,In_1247);
and U2000 (N_2000,In_355,In_1144);
and U2001 (N_2001,In_480,In_880);
nor U2002 (N_2002,In_1101,In_796);
or U2003 (N_2003,In_151,In_196);
and U2004 (N_2004,In_522,In_890);
nand U2005 (N_2005,In_1123,In_1151);
or U2006 (N_2006,In_1296,In_313);
and U2007 (N_2007,In_1103,In_1169);
nand U2008 (N_2008,In_495,In_363);
and U2009 (N_2009,In_1190,In_943);
nand U2010 (N_2010,In_1320,In_405);
nor U2011 (N_2011,In_1052,In_990);
or U2012 (N_2012,In_1146,In_726);
and U2013 (N_2013,In_973,In_390);
nor U2014 (N_2014,In_515,In_541);
nor U2015 (N_2015,In_31,In_1145);
and U2016 (N_2016,In_1197,In_1291);
or U2017 (N_2017,In_38,In_1194);
and U2018 (N_2018,In_596,In_344);
or U2019 (N_2019,In_381,In_1194);
nand U2020 (N_2020,In_480,In_75);
and U2021 (N_2021,In_1366,In_1369);
nand U2022 (N_2022,In_1100,In_906);
nand U2023 (N_2023,In_279,In_1174);
nand U2024 (N_2024,In_566,In_791);
or U2025 (N_2025,In_141,In_456);
nor U2026 (N_2026,In_623,In_1318);
and U2027 (N_2027,In_722,In_604);
nor U2028 (N_2028,In_1020,In_244);
nand U2029 (N_2029,In_771,In_161);
nand U2030 (N_2030,In_876,In_267);
and U2031 (N_2031,In_1110,In_396);
or U2032 (N_2032,In_941,In_714);
nand U2033 (N_2033,In_836,In_82);
nor U2034 (N_2034,In_301,In_344);
nand U2035 (N_2035,In_584,In_1204);
or U2036 (N_2036,In_753,In_322);
or U2037 (N_2037,In_387,In_1220);
or U2038 (N_2038,In_144,In_1493);
or U2039 (N_2039,In_1469,In_386);
or U2040 (N_2040,In_1343,In_433);
and U2041 (N_2041,In_1101,In_434);
and U2042 (N_2042,In_474,In_497);
nand U2043 (N_2043,In_834,In_702);
nor U2044 (N_2044,In_1447,In_1032);
or U2045 (N_2045,In_1321,In_371);
and U2046 (N_2046,In_733,In_1257);
and U2047 (N_2047,In_266,In_436);
nor U2048 (N_2048,In_1002,In_1173);
and U2049 (N_2049,In_1135,In_511);
and U2050 (N_2050,In_1474,In_1341);
and U2051 (N_2051,In_798,In_201);
nor U2052 (N_2052,In_1019,In_1361);
nor U2053 (N_2053,In_853,In_307);
nor U2054 (N_2054,In_1122,In_885);
nand U2055 (N_2055,In_534,In_1150);
or U2056 (N_2056,In_1234,In_229);
or U2057 (N_2057,In_1284,In_826);
xnor U2058 (N_2058,In_416,In_112);
or U2059 (N_2059,In_578,In_865);
nand U2060 (N_2060,In_941,In_354);
nor U2061 (N_2061,In_1400,In_1231);
nor U2062 (N_2062,In_1119,In_1277);
and U2063 (N_2063,In_1083,In_260);
nor U2064 (N_2064,In_1487,In_382);
nand U2065 (N_2065,In_903,In_820);
and U2066 (N_2066,In_312,In_1353);
or U2067 (N_2067,In_283,In_413);
nor U2068 (N_2068,In_396,In_1101);
nand U2069 (N_2069,In_787,In_406);
nor U2070 (N_2070,In_622,In_750);
nand U2071 (N_2071,In_246,In_1028);
and U2072 (N_2072,In_202,In_871);
and U2073 (N_2073,In_925,In_1114);
nand U2074 (N_2074,In_548,In_764);
and U2075 (N_2075,In_962,In_778);
or U2076 (N_2076,In_99,In_158);
nor U2077 (N_2077,In_387,In_864);
and U2078 (N_2078,In_125,In_844);
or U2079 (N_2079,In_51,In_315);
or U2080 (N_2080,In_1032,In_318);
or U2081 (N_2081,In_406,In_120);
and U2082 (N_2082,In_1063,In_1499);
or U2083 (N_2083,In_46,In_988);
nor U2084 (N_2084,In_561,In_783);
nor U2085 (N_2085,In_1031,In_474);
nor U2086 (N_2086,In_879,In_413);
or U2087 (N_2087,In_340,In_609);
or U2088 (N_2088,In_813,In_644);
nand U2089 (N_2089,In_771,In_1037);
nor U2090 (N_2090,In_810,In_97);
xnor U2091 (N_2091,In_1241,In_1204);
nor U2092 (N_2092,In_45,In_1357);
nor U2093 (N_2093,In_216,In_1441);
or U2094 (N_2094,In_925,In_1341);
nor U2095 (N_2095,In_127,In_914);
or U2096 (N_2096,In_1050,In_411);
nand U2097 (N_2097,In_1499,In_1241);
or U2098 (N_2098,In_82,In_298);
nor U2099 (N_2099,In_177,In_717);
nand U2100 (N_2100,In_338,In_37);
nand U2101 (N_2101,In_128,In_807);
nand U2102 (N_2102,In_629,In_727);
nor U2103 (N_2103,In_35,In_89);
nor U2104 (N_2104,In_233,In_900);
and U2105 (N_2105,In_468,In_1256);
or U2106 (N_2106,In_1077,In_326);
or U2107 (N_2107,In_1484,In_230);
and U2108 (N_2108,In_774,In_563);
nand U2109 (N_2109,In_1409,In_1375);
and U2110 (N_2110,In_945,In_179);
nor U2111 (N_2111,In_1066,In_108);
nand U2112 (N_2112,In_1419,In_1047);
nor U2113 (N_2113,In_450,In_1136);
and U2114 (N_2114,In_188,In_546);
nand U2115 (N_2115,In_1143,In_482);
or U2116 (N_2116,In_935,In_217);
and U2117 (N_2117,In_578,In_1060);
and U2118 (N_2118,In_899,In_785);
and U2119 (N_2119,In_304,In_421);
nand U2120 (N_2120,In_1077,In_70);
nor U2121 (N_2121,In_600,In_747);
nand U2122 (N_2122,In_467,In_1456);
nand U2123 (N_2123,In_1456,In_669);
nand U2124 (N_2124,In_864,In_824);
nor U2125 (N_2125,In_334,In_578);
nor U2126 (N_2126,In_920,In_230);
nor U2127 (N_2127,In_1230,In_465);
and U2128 (N_2128,In_1268,In_1135);
nand U2129 (N_2129,In_1313,In_1179);
and U2130 (N_2130,In_1373,In_1004);
nor U2131 (N_2131,In_912,In_1480);
nand U2132 (N_2132,In_1483,In_767);
and U2133 (N_2133,In_100,In_530);
nor U2134 (N_2134,In_188,In_313);
nor U2135 (N_2135,In_654,In_72);
nor U2136 (N_2136,In_291,In_158);
and U2137 (N_2137,In_123,In_1479);
nor U2138 (N_2138,In_802,In_260);
and U2139 (N_2139,In_202,In_1181);
nand U2140 (N_2140,In_95,In_1175);
nor U2141 (N_2141,In_279,In_700);
nor U2142 (N_2142,In_1110,In_1431);
and U2143 (N_2143,In_946,In_333);
or U2144 (N_2144,In_1232,In_51);
or U2145 (N_2145,In_419,In_1287);
nor U2146 (N_2146,In_828,In_119);
or U2147 (N_2147,In_893,In_525);
nand U2148 (N_2148,In_947,In_941);
nor U2149 (N_2149,In_519,In_657);
and U2150 (N_2150,In_123,In_136);
or U2151 (N_2151,In_391,In_885);
nor U2152 (N_2152,In_922,In_1409);
nor U2153 (N_2153,In_144,In_1377);
and U2154 (N_2154,In_216,In_99);
and U2155 (N_2155,In_603,In_1125);
nand U2156 (N_2156,In_57,In_896);
and U2157 (N_2157,In_337,In_1490);
or U2158 (N_2158,In_868,In_421);
and U2159 (N_2159,In_661,In_1030);
or U2160 (N_2160,In_933,In_162);
or U2161 (N_2161,In_806,In_1156);
or U2162 (N_2162,In_931,In_1448);
nand U2163 (N_2163,In_1331,In_1214);
nand U2164 (N_2164,In_365,In_1354);
and U2165 (N_2165,In_1316,In_136);
and U2166 (N_2166,In_801,In_169);
and U2167 (N_2167,In_1204,In_501);
nor U2168 (N_2168,In_1145,In_551);
and U2169 (N_2169,In_75,In_424);
nand U2170 (N_2170,In_960,In_10);
nand U2171 (N_2171,In_501,In_1279);
nor U2172 (N_2172,In_99,In_915);
or U2173 (N_2173,In_323,In_1473);
nor U2174 (N_2174,In_132,In_213);
nor U2175 (N_2175,In_346,In_51);
or U2176 (N_2176,In_114,In_907);
nor U2177 (N_2177,In_377,In_807);
or U2178 (N_2178,In_111,In_718);
or U2179 (N_2179,In_1296,In_441);
nand U2180 (N_2180,In_1,In_101);
or U2181 (N_2181,In_990,In_1011);
or U2182 (N_2182,In_332,In_1115);
or U2183 (N_2183,In_858,In_118);
nor U2184 (N_2184,In_913,In_70);
and U2185 (N_2185,In_1018,In_864);
nor U2186 (N_2186,In_1235,In_814);
or U2187 (N_2187,In_1438,In_1050);
nor U2188 (N_2188,In_989,In_647);
nor U2189 (N_2189,In_1263,In_835);
nor U2190 (N_2190,In_785,In_915);
and U2191 (N_2191,In_485,In_763);
and U2192 (N_2192,In_61,In_354);
or U2193 (N_2193,In_47,In_404);
nand U2194 (N_2194,In_344,In_454);
nor U2195 (N_2195,In_605,In_1232);
nor U2196 (N_2196,In_1477,In_885);
nand U2197 (N_2197,In_676,In_608);
nand U2198 (N_2198,In_696,In_1240);
and U2199 (N_2199,In_1079,In_520);
nand U2200 (N_2200,In_1031,In_285);
nor U2201 (N_2201,In_1160,In_1155);
and U2202 (N_2202,In_726,In_83);
nor U2203 (N_2203,In_1008,In_919);
xnor U2204 (N_2204,In_812,In_200);
and U2205 (N_2205,In_1493,In_828);
nand U2206 (N_2206,In_684,In_120);
nor U2207 (N_2207,In_357,In_134);
nor U2208 (N_2208,In_1169,In_630);
nor U2209 (N_2209,In_534,In_377);
and U2210 (N_2210,In_1175,In_753);
or U2211 (N_2211,In_580,In_369);
nand U2212 (N_2212,In_119,In_1084);
nand U2213 (N_2213,In_387,In_1044);
nand U2214 (N_2214,In_169,In_120);
or U2215 (N_2215,In_794,In_800);
nor U2216 (N_2216,In_1390,In_654);
nand U2217 (N_2217,In_946,In_1309);
and U2218 (N_2218,In_699,In_1442);
and U2219 (N_2219,In_58,In_1286);
nand U2220 (N_2220,In_980,In_118);
nor U2221 (N_2221,In_197,In_1254);
nor U2222 (N_2222,In_1035,In_968);
and U2223 (N_2223,In_1187,In_1175);
and U2224 (N_2224,In_641,In_1238);
nor U2225 (N_2225,In_1294,In_741);
nand U2226 (N_2226,In_534,In_1234);
nor U2227 (N_2227,In_390,In_849);
and U2228 (N_2228,In_1458,In_1007);
or U2229 (N_2229,In_1495,In_280);
or U2230 (N_2230,In_446,In_1317);
nand U2231 (N_2231,In_356,In_418);
and U2232 (N_2232,In_810,In_219);
or U2233 (N_2233,In_151,In_1335);
or U2234 (N_2234,In_963,In_533);
nor U2235 (N_2235,In_310,In_1478);
nor U2236 (N_2236,In_973,In_752);
or U2237 (N_2237,In_687,In_879);
or U2238 (N_2238,In_1424,In_1191);
nor U2239 (N_2239,In_997,In_453);
nor U2240 (N_2240,In_593,In_663);
or U2241 (N_2241,In_412,In_538);
nand U2242 (N_2242,In_1113,In_963);
nor U2243 (N_2243,In_499,In_996);
nand U2244 (N_2244,In_1053,In_732);
nand U2245 (N_2245,In_41,In_976);
and U2246 (N_2246,In_829,In_359);
nand U2247 (N_2247,In_682,In_1422);
nand U2248 (N_2248,In_255,In_523);
nand U2249 (N_2249,In_655,In_635);
or U2250 (N_2250,In_1027,In_790);
and U2251 (N_2251,In_736,In_626);
nor U2252 (N_2252,In_639,In_817);
or U2253 (N_2253,In_1443,In_1217);
nor U2254 (N_2254,In_762,In_456);
and U2255 (N_2255,In_147,In_250);
and U2256 (N_2256,In_903,In_173);
nor U2257 (N_2257,In_1423,In_1413);
and U2258 (N_2258,In_939,In_1398);
and U2259 (N_2259,In_1306,In_612);
nand U2260 (N_2260,In_109,In_1329);
or U2261 (N_2261,In_1255,In_522);
or U2262 (N_2262,In_40,In_482);
nand U2263 (N_2263,In_998,In_1330);
or U2264 (N_2264,In_353,In_621);
nand U2265 (N_2265,In_638,In_300);
nor U2266 (N_2266,In_1275,In_1397);
nor U2267 (N_2267,In_284,In_1469);
nor U2268 (N_2268,In_18,In_1136);
nand U2269 (N_2269,In_1175,In_790);
or U2270 (N_2270,In_778,In_2);
or U2271 (N_2271,In_1177,In_1279);
nor U2272 (N_2272,In_395,In_830);
and U2273 (N_2273,In_1038,In_126);
and U2274 (N_2274,In_792,In_555);
nand U2275 (N_2275,In_227,In_508);
nor U2276 (N_2276,In_649,In_402);
or U2277 (N_2277,In_1313,In_1200);
nand U2278 (N_2278,In_49,In_988);
xnor U2279 (N_2279,In_319,In_1332);
nor U2280 (N_2280,In_564,In_91);
and U2281 (N_2281,In_807,In_1036);
and U2282 (N_2282,In_1480,In_726);
or U2283 (N_2283,In_287,In_506);
or U2284 (N_2284,In_135,In_951);
and U2285 (N_2285,In_171,In_1338);
nor U2286 (N_2286,In_401,In_810);
nand U2287 (N_2287,In_1030,In_255);
nand U2288 (N_2288,In_345,In_1026);
or U2289 (N_2289,In_1191,In_1139);
or U2290 (N_2290,In_1041,In_698);
nor U2291 (N_2291,In_698,In_50);
and U2292 (N_2292,In_73,In_1315);
nand U2293 (N_2293,In_1163,In_665);
nor U2294 (N_2294,In_129,In_82);
and U2295 (N_2295,In_1260,In_499);
nand U2296 (N_2296,In_1093,In_108);
nand U2297 (N_2297,In_0,In_1488);
nand U2298 (N_2298,In_697,In_1467);
nand U2299 (N_2299,In_93,In_716);
nand U2300 (N_2300,In_631,In_1243);
nand U2301 (N_2301,In_144,In_41);
and U2302 (N_2302,In_698,In_1419);
nand U2303 (N_2303,In_1125,In_928);
nor U2304 (N_2304,In_1084,In_912);
and U2305 (N_2305,In_1245,In_1253);
nor U2306 (N_2306,In_441,In_152);
nor U2307 (N_2307,In_825,In_704);
nand U2308 (N_2308,In_1190,In_407);
nor U2309 (N_2309,In_119,In_702);
nor U2310 (N_2310,In_317,In_34);
and U2311 (N_2311,In_1269,In_736);
and U2312 (N_2312,In_1410,In_906);
nor U2313 (N_2313,In_1367,In_632);
nand U2314 (N_2314,In_1027,In_553);
nor U2315 (N_2315,In_196,In_154);
or U2316 (N_2316,In_407,In_418);
and U2317 (N_2317,In_714,In_860);
or U2318 (N_2318,In_206,In_227);
and U2319 (N_2319,In_938,In_174);
nor U2320 (N_2320,In_1151,In_1261);
nand U2321 (N_2321,In_609,In_547);
or U2322 (N_2322,In_497,In_1414);
and U2323 (N_2323,In_798,In_1479);
and U2324 (N_2324,In_305,In_1188);
xor U2325 (N_2325,In_169,In_362);
and U2326 (N_2326,In_578,In_458);
nor U2327 (N_2327,In_1406,In_218);
or U2328 (N_2328,In_164,In_102);
nor U2329 (N_2329,In_1214,In_926);
or U2330 (N_2330,In_1169,In_1040);
nand U2331 (N_2331,In_1261,In_768);
and U2332 (N_2332,In_950,In_773);
nor U2333 (N_2333,In_762,In_1143);
nor U2334 (N_2334,In_687,In_1436);
or U2335 (N_2335,In_1182,In_1020);
and U2336 (N_2336,In_390,In_767);
nand U2337 (N_2337,In_876,In_316);
and U2338 (N_2338,In_1004,In_120);
and U2339 (N_2339,In_899,In_606);
and U2340 (N_2340,In_556,In_312);
nand U2341 (N_2341,In_141,In_1391);
nand U2342 (N_2342,In_273,In_157);
or U2343 (N_2343,In_1139,In_809);
nand U2344 (N_2344,In_846,In_616);
or U2345 (N_2345,In_1037,In_659);
nand U2346 (N_2346,In_356,In_714);
and U2347 (N_2347,In_826,In_1456);
nand U2348 (N_2348,In_1006,In_475);
and U2349 (N_2349,In_983,In_234);
and U2350 (N_2350,In_712,In_1383);
or U2351 (N_2351,In_1414,In_1474);
nor U2352 (N_2352,In_1327,In_1154);
nand U2353 (N_2353,In_1426,In_123);
and U2354 (N_2354,In_643,In_1331);
nand U2355 (N_2355,In_1141,In_764);
nand U2356 (N_2356,In_207,In_161);
nor U2357 (N_2357,In_1177,In_725);
nor U2358 (N_2358,In_361,In_980);
and U2359 (N_2359,In_668,In_358);
nand U2360 (N_2360,In_434,In_1380);
nand U2361 (N_2361,In_695,In_591);
and U2362 (N_2362,In_440,In_1469);
or U2363 (N_2363,In_653,In_1433);
nand U2364 (N_2364,In_328,In_129);
nand U2365 (N_2365,In_1,In_1298);
or U2366 (N_2366,In_555,In_7);
nand U2367 (N_2367,In_658,In_335);
nand U2368 (N_2368,In_875,In_240);
or U2369 (N_2369,In_1155,In_1129);
and U2370 (N_2370,In_489,In_585);
and U2371 (N_2371,In_1146,In_938);
and U2372 (N_2372,In_1104,In_718);
and U2373 (N_2373,In_1156,In_1348);
nor U2374 (N_2374,In_343,In_500);
nor U2375 (N_2375,In_1072,In_932);
nand U2376 (N_2376,In_942,In_1040);
or U2377 (N_2377,In_820,In_1038);
nand U2378 (N_2378,In_116,In_759);
or U2379 (N_2379,In_1270,In_275);
nand U2380 (N_2380,In_731,In_1242);
nor U2381 (N_2381,In_81,In_271);
nand U2382 (N_2382,In_434,In_369);
and U2383 (N_2383,In_682,In_458);
and U2384 (N_2384,In_553,In_1376);
nand U2385 (N_2385,In_928,In_1135);
nor U2386 (N_2386,In_568,In_1313);
or U2387 (N_2387,In_19,In_473);
and U2388 (N_2388,In_1267,In_1230);
nand U2389 (N_2389,In_130,In_16);
nand U2390 (N_2390,In_942,In_1271);
nand U2391 (N_2391,In_1463,In_590);
or U2392 (N_2392,In_1155,In_14);
nor U2393 (N_2393,In_281,In_1067);
and U2394 (N_2394,In_930,In_180);
nand U2395 (N_2395,In_28,In_1316);
or U2396 (N_2396,In_266,In_101);
xnor U2397 (N_2397,In_760,In_947);
nor U2398 (N_2398,In_240,In_788);
nand U2399 (N_2399,In_724,In_839);
or U2400 (N_2400,In_1195,In_253);
or U2401 (N_2401,In_1190,In_373);
nor U2402 (N_2402,In_1063,In_1339);
or U2403 (N_2403,In_377,In_530);
or U2404 (N_2404,In_594,In_1350);
nor U2405 (N_2405,In_437,In_111);
and U2406 (N_2406,In_667,In_934);
and U2407 (N_2407,In_969,In_389);
and U2408 (N_2408,In_1174,In_851);
or U2409 (N_2409,In_824,In_486);
or U2410 (N_2410,In_585,In_717);
or U2411 (N_2411,In_890,In_1228);
or U2412 (N_2412,In_425,In_837);
nand U2413 (N_2413,In_948,In_1243);
and U2414 (N_2414,In_264,In_502);
nor U2415 (N_2415,In_701,In_179);
nor U2416 (N_2416,In_882,In_265);
nor U2417 (N_2417,In_1038,In_920);
nand U2418 (N_2418,In_1146,In_893);
nor U2419 (N_2419,In_97,In_777);
nor U2420 (N_2420,In_330,In_925);
nor U2421 (N_2421,In_468,In_748);
and U2422 (N_2422,In_1284,In_622);
or U2423 (N_2423,In_926,In_1372);
and U2424 (N_2424,In_486,In_1213);
and U2425 (N_2425,In_1447,In_126);
nor U2426 (N_2426,In_757,In_1192);
nor U2427 (N_2427,In_37,In_208);
nand U2428 (N_2428,In_237,In_1192);
nand U2429 (N_2429,In_865,In_764);
nand U2430 (N_2430,In_273,In_1063);
or U2431 (N_2431,In_56,In_545);
and U2432 (N_2432,In_433,In_390);
nand U2433 (N_2433,In_463,In_324);
or U2434 (N_2434,In_1058,In_153);
and U2435 (N_2435,In_511,In_638);
nand U2436 (N_2436,In_308,In_449);
nor U2437 (N_2437,In_403,In_3);
and U2438 (N_2438,In_126,In_1134);
nor U2439 (N_2439,In_492,In_942);
nor U2440 (N_2440,In_962,In_547);
nor U2441 (N_2441,In_606,In_1257);
nand U2442 (N_2442,In_765,In_399);
nor U2443 (N_2443,In_982,In_99);
nand U2444 (N_2444,In_1469,In_411);
and U2445 (N_2445,In_1253,In_1310);
and U2446 (N_2446,In_1331,In_170);
or U2447 (N_2447,In_1329,In_668);
nor U2448 (N_2448,In_227,In_619);
xor U2449 (N_2449,In_1050,In_1463);
and U2450 (N_2450,In_228,In_646);
nand U2451 (N_2451,In_176,In_56);
or U2452 (N_2452,In_234,In_1367);
nand U2453 (N_2453,In_860,In_280);
nand U2454 (N_2454,In_1338,In_1041);
and U2455 (N_2455,In_40,In_547);
nand U2456 (N_2456,In_191,In_333);
nor U2457 (N_2457,In_641,In_687);
and U2458 (N_2458,In_222,In_1211);
nand U2459 (N_2459,In_308,In_1178);
or U2460 (N_2460,In_659,In_1266);
nor U2461 (N_2461,In_1097,In_83);
nand U2462 (N_2462,In_1437,In_1289);
nor U2463 (N_2463,In_1172,In_573);
or U2464 (N_2464,In_382,In_459);
nor U2465 (N_2465,In_192,In_1247);
nor U2466 (N_2466,In_1366,In_1456);
nand U2467 (N_2467,In_585,In_668);
nand U2468 (N_2468,In_492,In_654);
nor U2469 (N_2469,In_162,In_149);
and U2470 (N_2470,In_1362,In_348);
nand U2471 (N_2471,In_722,In_417);
or U2472 (N_2472,In_1072,In_1227);
nand U2473 (N_2473,In_405,In_383);
nand U2474 (N_2474,In_349,In_657);
and U2475 (N_2475,In_1055,In_93);
or U2476 (N_2476,In_104,In_134);
or U2477 (N_2477,In_300,In_1249);
and U2478 (N_2478,In_397,In_1345);
nand U2479 (N_2479,In_19,In_462);
or U2480 (N_2480,In_3,In_1176);
nor U2481 (N_2481,In_762,In_941);
or U2482 (N_2482,In_32,In_1240);
and U2483 (N_2483,In_924,In_298);
nor U2484 (N_2484,In_1008,In_14);
nor U2485 (N_2485,In_696,In_409);
and U2486 (N_2486,In_1018,In_1311);
nor U2487 (N_2487,In_631,In_484);
nand U2488 (N_2488,In_1068,In_101);
nor U2489 (N_2489,In_984,In_1043);
nand U2490 (N_2490,In_934,In_53);
and U2491 (N_2491,In_58,In_47);
nor U2492 (N_2492,In_1408,In_995);
nor U2493 (N_2493,In_1415,In_1027);
or U2494 (N_2494,In_1431,In_821);
and U2495 (N_2495,In_328,In_489);
or U2496 (N_2496,In_1241,In_1464);
or U2497 (N_2497,In_1354,In_1112);
or U2498 (N_2498,In_1299,In_1067);
or U2499 (N_2499,In_95,In_126);
nand U2500 (N_2500,In_662,In_416);
nor U2501 (N_2501,In_142,In_113);
or U2502 (N_2502,In_1351,In_215);
or U2503 (N_2503,In_858,In_1181);
and U2504 (N_2504,In_1260,In_164);
or U2505 (N_2505,In_568,In_253);
nor U2506 (N_2506,In_129,In_240);
nand U2507 (N_2507,In_1302,In_853);
nor U2508 (N_2508,In_566,In_170);
and U2509 (N_2509,In_1407,In_1158);
nor U2510 (N_2510,In_410,In_1351);
nor U2511 (N_2511,In_925,In_1215);
nor U2512 (N_2512,In_246,In_1298);
and U2513 (N_2513,In_639,In_1211);
nor U2514 (N_2514,In_764,In_428);
nand U2515 (N_2515,In_891,In_511);
or U2516 (N_2516,In_122,In_1341);
or U2517 (N_2517,In_84,In_264);
nor U2518 (N_2518,In_977,In_1200);
nand U2519 (N_2519,In_464,In_1389);
nor U2520 (N_2520,In_1141,In_94);
nor U2521 (N_2521,In_1264,In_1066);
nor U2522 (N_2522,In_715,In_784);
nand U2523 (N_2523,In_990,In_494);
or U2524 (N_2524,In_1480,In_26);
and U2525 (N_2525,In_734,In_565);
nor U2526 (N_2526,In_870,In_339);
nor U2527 (N_2527,In_1072,In_445);
or U2528 (N_2528,In_1155,In_1418);
nand U2529 (N_2529,In_253,In_156);
or U2530 (N_2530,In_18,In_970);
nand U2531 (N_2531,In_1014,In_810);
and U2532 (N_2532,In_43,In_733);
xnor U2533 (N_2533,In_321,In_102);
nand U2534 (N_2534,In_1010,In_796);
nand U2535 (N_2535,In_1407,In_31);
nand U2536 (N_2536,In_1214,In_1301);
and U2537 (N_2537,In_279,In_720);
nor U2538 (N_2538,In_634,In_1282);
nor U2539 (N_2539,In_1051,In_1305);
nor U2540 (N_2540,In_1499,In_111);
nor U2541 (N_2541,In_1093,In_238);
or U2542 (N_2542,In_300,In_931);
or U2543 (N_2543,In_1118,In_586);
or U2544 (N_2544,In_1436,In_281);
or U2545 (N_2545,In_1440,In_1406);
and U2546 (N_2546,In_248,In_967);
nand U2547 (N_2547,In_1042,In_905);
and U2548 (N_2548,In_1089,In_1290);
nor U2549 (N_2549,In_1337,In_208);
nand U2550 (N_2550,In_200,In_584);
or U2551 (N_2551,In_779,In_457);
nand U2552 (N_2552,In_795,In_1331);
or U2553 (N_2553,In_1220,In_1157);
or U2554 (N_2554,In_1164,In_198);
and U2555 (N_2555,In_576,In_1086);
nor U2556 (N_2556,In_999,In_1295);
and U2557 (N_2557,In_1419,In_1094);
or U2558 (N_2558,In_238,In_1472);
nand U2559 (N_2559,In_660,In_504);
or U2560 (N_2560,In_1280,In_692);
xnor U2561 (N_2561,In_1474,In_167);
nand U2562 (N_2562,In_1212,In_1155);
nor U2563 (N_2563,In_1034,In_381);
nand U2564 (N_2564,In_121,In_473);
and U2565 (N_2565,In_1148,In_48);
nor U2566 (N_2566,In_1405,In_1291);
and U2567 (N_2567,In_757,In_745);
nor U2568 (N_2568,In_782,In_571);
nor U2569 (N_2569,In_396,In_919);
or U2570 (N_2570,In_651,In_658);
nand U2571 (N_2571,In_1125,In_1157);
nor U2572 (N_2572,In_37,In_79);
nand U2573 (N_2573,In_874,In_162);
or U2574 (N_2574,In_613,In_707);
and U2575 (N_2575,In_1063,In_260);
nand U2576 (N_2576,In_1004,In_1365);
and U2577 (N_2577,In_1192,In_817);
and U2578 (N_2578,In_311,In_781);
nor U2579 (N_2579,In_795,In_533);
nor U2580 (N_2580,In_848,In_76);
nand U2581 (N_2581,In_1170,In_1010);
or U2582 (N_2582,In_1318,In_1176);
or U2583 (N_2583,In_755,In_1036);
nand U2584 (N_2584,In_1278,In_166);
nand U2585 (N_2585,In_767,In_1098);
nor U2586 (N_2586,In_1040,In_779);
and U2587 (N_2587,In_1241,In_271);
nor U2588 (N_2588,In_618,In_1358);
and U2589 (N_2589,In_594,In_1157);
nor U2590 (N_2590,In_714,In_816);
nor U2591 (N_2591,In_6,In_626);
nor U2592 (N_2592,In_816,In_147);
or U2593 (N_2593,In_11,In_35);
and U2594 (N_2594,In_107,In_903);
or U2595 (N_2595,In_904,In_906);
nor U2596 (N_2596,In_1107,In_350);
or U2597 (N_2597,In_1178,In_490);
nor U2598 (N_2598,In_861,In_111);
or U2599 (N_2599,In_1178,In_1433);
or U2600 (N_2600,In_359,In_753);
nand U2601 (N_2601,In_1042,In_198);
or U2602 (N_2602,In_15,In_645);
or U2603 (N_2603,In_797,In_615);
nand U2604 (N_2604,In_399,In_1235);
or U2605 (N_2605,In_1234,In_156);
nor U2606 (N_2606,In_920,In_1123);
and U2607 (N_2607,In_650,In_260);
nand U2608 (N_2608,In_537,In_826);
and U2609 (N_2609,In_1113,In_382);
nand U2610 (N_2610,In_510,In_82);
nand U2611 (N_2611,In_1324,In_1408);
nand U2612 (N_2612,In_1327,In_726);
or U2613 (N_2613,In_771,In_351);
nand U2614 (N_2614,In_740,In_440);
nor U2615 (N_2615,In_1200,In_1409);
nand U2616 (N_2616,In_523,In_1179);
nor U2617 (N_2617,In_621,In_332);
or U2618 (N_2618,In_516,In_712);
and U2619 (N_2619,In_120,In_644);
nor U2620 (N_2620,In_690,In_1188);
and U2621 (N_2621,In_466,In_1142);
or U2622 (N_2622,In_622,In_1117);
nor U2623 (N_2623,In_46,In_1102);
nand U2624 (N_2624,In_355,In_725);
nor U2625 (N_2625,In_1024,In_797);
and U2626 (N_2626,In_901,In_1007);
xnor U2627 (N_2627,In_355,In_1042);
and U2628 (N_2628,In_1147,In_1260);
and U2629 (N_2629,In_886,In_1050);
nand U2630 (N_2630,In_1088,In_1116);
and U2631 (N_2631,In_621,In_773);
and U2632 (N_2632,In_898,In_839);
or U2633 (N_2633,In_471,In_528);
and U2634 (N_2634,In_159,In_1314);
or U2635 (N_2635,In_985,In_161);
nand U2636 (N_2636,In_868,In_1116);
nand U2637 (N_2637,In_1212,In_794);
nor U2638 (N_2638,In_1221,In_627);
nor U2639 (N_2639,In_984,In_925);
nor U2640 (N_2640,In_1195,In_810);
or U2641 (N_2641,In_940,In_405);
and U2642 (N_2642,In_460,In_95);
nor U2643 (N_2643,In_697,In_1048);
nand U2644 (N_2644,In_186,In_976);
nand U2645 (N_2645,In_1196,In_488);
nor U2646 (N_2646,In_900,In_877);
or U2647 (N_2647,In_301,In_1315);
and U2648 (N_2648,In_1108,In_566);
nor U2649 (N_2649,In_656,In_628);
nand U2650 (N_2650,In_1242,In_196);
or U2651 (N_2651,In_549,In_12);
and U2652 (N_2652,In_1320,In_182);
nor U2653 (N_2653,In_683,In_689);
and U2654 (N_2654,In_1166,In_1469);
and U2655 (N_2655,In_174,In_1177);
nand U2656 (N_2656,In_70,In_1198);
nor U2657 (N_2657,In_604,In_848);
nor U2658 (N_2658,In_617,In_1214);
and U2659 (N_2659,In_1068,In_1145);
nor U2660 (N_2660,In_1485,In_780);
and U2661 (N_2661,In_1457,In_693);
and U2662 (N_2662,In_1218,In_1040);
nor U2663 (N_2663,In_516,In_166);
nor U2664 (N_2664,In_1169,In_1153);
nor U2665 (N_2665,In_634,In_253);
nor U2666 (N_2666,In_290,In_610);
nand U2667 (N_2667,In_589,In_664);
or U2668 (N_2668,In_228,In_1210);
or U2669 (N_2669,In_188,In_1147);
or U2670 (N_2670,In_1304,In_384);
or U2671 (N_2671,In_1474,In_656);
or U2672 (N_2672,In_916,In_1030);
nand U2673 (N_2673,In_1306,In_1430);
or U2674 (N_2674,In_757,In_186);
or U2675 (N_2675,In_451,In_1183);
or U2676 (N_2676,In_562,In_896);
nor U2677 (N_2677,In_955,In_1091);
and U2678 (N_2678,In_958,In_487);
nand U2679 (N_2679,In_516,In_298);
and U2680 (N_2680,In_343,In_1301);
nand U2681 (N_2681,In_1045,In_177);
nand U2682 (N_2682,In_77,In_1143);
and U2683 (N_2683,In_841,In_353);
or U2684 (N_2684,In_1232,In_1237);
nor U2685 (N_2685,In_621,In_336);
and U2686 (N_2686,In_1023,In_124);
and U2687 (N_2687,In_493,In_349);
nand U2688 (N_2688,In_392,In_1188);
or U2689 (N_2689,In_730,In_93);
nand U2690 (N_2690,In_136,In_642);
nor U2691 (N_2691,In_143,In_487);
nor U2692 (N_2692,In_350,In_184);
nand U2693 (N_2693,In_390,In_921);
or U2694 (N_2694,In_1434,In_1019);
or U2695 (N_2695,In_161,In_828);
nand U2696 (N_2696,In_769,In_736);
or U2697 (N_2697,In_944,In_87);
or U2698 (N_2698,In_491,In_372);
or U2699 (N_2699,In_159,In_755);
nor U2700 (N_2700,In_697,In_571);
nor U2701 (N_2701,In_250,In_115);
or U2702 (N_2702,In_1397,In_451);
or U2703 (N_2703,In_1405,In_860);
nor U2704 (N_2704,In_446,In_863);
nand U2705 (N_2705,In_753,In_1007);
nor U2706 (N_2706,In_1082,In_1486);
or U2707 (N_2707,In_899,In_1182);
nor U2708 (N_2708,In_1168,In_103);
nand U2709 (N_2709,In_1080,In_1260);
or U2710 (N_2710,In_1055,In_1256);
or U2711 (N_2711,In_648,In_1053);
nand U2712 (N_2712,In_594,In_413);
nand U2713 (N_2713,In_761,In_1461);
and U2714 (N_2714,In_561,In_112);
or U2715 (N_2715,In_1287,In_1485);
nor U2716 (N_2716,In_593,In_580);
nor U2717 (N_2717,In_796,In_694);
or U2718 (N_2718,In_632,In_769);
or U2719 (N_2719,In_1093,In_1362);
nor U2720 (N_2720,In_1327,In_264);
xnor U2721 (N_2721,In_382,In_822);
nand U2722 (N_2722,In_286,In_578);
or U2723 (N_2723,In_869,In_557);
and U2724 (N_2724,In_316,In_255);
and U2725 (N_2725,In_1409,In_356);
or U2726 (N_2726,In_1124,In_55);
nor U2727 (N_2727,In_502,In_283);
nand U2728 (N_2728,In_690,In_474);
or U2729 (N_2729,In_286,In_1008);
or U2730 (N_2730,In_961,In_76);
nand U2731 (N_2731,In_740,In_1373);
and U2732 (N_2732,In_446,In_268);
nor U2733 (N_2733,In_58,In_331);
nand U2734 (N_2734,In_1270,In_1462);
nand U2735 (N_2735,In_57,In_181);
or U2736 (N_2736,In_593,In_1138);
nand U2737 (N_2737,In_1394,In_1482);
nor U2738 (N_2738,In_1105,In_777);
and U2739 (N_2739,In_208,In_1049);
nor U2740 (N_2740,In_1100,In_305);
or U2741 (N_2741,In_238,In_1246);
or U2742 (N_2742,In_1495,In_1341);
nor U2743 (N_2743,In_1189,In_401);
and U2744 (N_2744,In_105,In_1389);
and U2745 (N_2745,In_13,In_408);
nor U2746 (N_2746,In_62,In_1007);
nor U2747 (N_2747,In_68,In_1045);
or U2748 (N_2748,In_567,In_503);
and U2749 (N_2749,In_1406,In_21);
nand U2750 (N_2750,In_1327,In_747);
nand U2751 (N_2751,In_1286,In_211);
or U2752 (N_2752,In_1143,In_63);
and U2753 (N_2753,In_1471,In_1156);
and U2754 (N_2754,In_268,In_601);
nand U2755 (N_2755,In_1161,In_1012);
and U2756 (N_2756,In_258,In_325);
nor U2757 (N_2757,In_525,In_695);
nand U2758 (N_2758,In_382,In_702);
nor U2759 (N_2759,In_752,In_89);
nor U2760 (N_2760,In_538,In_1140);
or U2761 (N_2761,In_363,In_259);
nor U2762 (N_2762,In_303,In_1079);
nand U2763 (N_2763,In_843,In_1440);
nor U2764 (N_2764,In_441,In_632);
nand U2765 (N_2765,In_43,In_772);
nor U2766 (N_2766,In_743,In_1004);
nor U2767 (N_2767,In_360,In_337);
and U2768 (N_2768,In_1307,In_1279);
nor U2769 (N_2769,In_229,In_395);
nor U2770 (N_2770,In_143,In_178);
or U2771 (N_2771,In_297,In_300);
or U2772 (N_2772,In_685,In_867);
nand U2773 (N_2773,In_768,In_512);
nor U2774 (N_2774,In_1321,In_311);
or U2775 (N_2775,In_801,In_1448);
and U2776 (N_2776,In_20,In_48);
and U2777 (N_2777,In_130,In_837);
and U2778 (N_2778,In_1479,In_394);
nor U2779 (N_2779,In_851,In_824);
and U2780 (N_2780,In_704,In_1192);
and U2781 (N_2781,In_1070,In_158);
or U2782 (N_2782,In_307,In_462);
and U2783 (N_2783,In_1451,In_795);
nor U2784 (N_2784,In_744,In_1333);
or U2785 (N_2785,In_1030,In_513);
and U2786 (N_2786,In_135,In_1466);
xnor U2787 (N_2787,In_811,In_280);
or U2788 (N_2788,In_1422,In_296);
or U2789 (N_2789,In_1202,In_1411);
and U2790 (N_2790,In_1085,In_483);
nor U2791 (N_2791,In_1452,In_384);
nor U2792 (N_2792,In_253,In_11);
nand U2793 (N_2793,In_182,In_422);
nor U2794 (N_2794,In_639,In_1191);
nand U2795 (N_2795,In_772,In_3);
and U2796 (N_2796,In_582,In_755);
nor U2797 (N_2797,In_1190,In_740);
nor U2798 (N_2798,In_331,In_1347);
and U2799 (N_2799,In_122,In_624);
nand U2800 (N_2800,In_698,In_451);
or U2801 (N_2801,In_509,In_398);
and U2802 (N_2802,In_172,In_1191);
nand U2803 (N_2803,In_393,In_1020);
nand U2804 (N_2804,In_97,In_1095);
nand U2805 (N_2805,In_1044,In_832);
and U2806 (N_2806,In_156,In_1324);
nor U2807 (N_2807,In_832,In_1287);
or U2808 (N_2808,In_1326,In_1420);
nand U2809 (N_2809,In_850,In_1128);
or U2810 (N_2810,In_512,In_1093);
nor U2811 (N_2811,In_925,In_284);
nor U2812 (N_2812,In_1044,In_545);
nor U2813 (N_2813,In_411,In_696);
nand U2814 (N_2814,In_852,In_800);
nor U2815 (N_2815,In_832,In_433);
and U2816 (N_2816,In_1104,In_586);
or U2817 (N_2817,In_650,In_591);
xnor U2818 (N_2818,In_822,In_454);
and U2819 (N_2819,In_744,In_28);
nand U2820 (N_2820,In_127,In_724);
nor U2821 (N_2821,In_1186,In_602);
and U2822 (N_2822,In_1457,In_1210);
and U2823 (N_2823,In_897,In_1089);
or U2824 (N_2824,In_117,In_1498);
and U2825 (N_2825,In_204,In_175);
nor U2826 (N_2826,In_986,In_72);
nor U2827 (N_2827,In_529,In_995);
and U2828 (N_2828,In_186,In_738);
or U2829 (N_2829,In_870,In_645);
and U2830 (N_2830,In_1216,In_15);
and U2831 (N_2831,In_1231,In_583);
or U2832 (N_2832,In_639,In_519);
and U2833 (N_2833,In_1153,In_479);
nor U2834 (N_2834,In_1408,In_670);
or U2835 (N_2835,In_1025,In_1009);
nand U2836 (N_2836,In_792,In_782);
or U2837 (N_2837,In_1377,In_1172);
and U2838 (N_2838,In_879,In_1338);
nor U2839 (N_2839,In_1403,In_363);
and U2840 (N_2840,In_933,In_117);
nor U2841 (N_2841,In_760,In_662);
or U2842 (N_2842,In_36,In_1385);
and U2843 (N_2843,In_730,In_818);
nand U2844 (N_2844,In_487,In_82);
or U2845 (N_2845,In_788,In_774);
nor U2846 (N_2846,In_732,In_933);
nor U2847 (N_2847,In_850,In_1226);
nor U2848 (N_2848,In_1091,In_842);
nor U2849 (N_2849,In_217,In_492);
nand U2850 (N_2850,In_812,In_664);
or U2851 (N_2851,In_774,In_1385);
nand U2852 (N_2852,In_468,In_842);
nand U2853 (N_2853,In_1001,In_247);
and U2854 (N_2854,In_700,In_522);
nand U2855 (N_2855,In_240,In_914);
or U2856 (N_2856,In_938,In_550);
and U2857 (N_2857,In_1408,In_1365);
nand U2858 (N_2858,In_828,In_1017);
and U2859 (N_2859,In_588,In_1213);
nand U2860 (N_2860,In_1205,In_830);
or U2861 (N_2861,In_863,In_896);
or U2862 (N_2862,In_1313,In_622);
nand U2863 (N_2863,In_293,In_968);
nand U2864 (N_2864,In_967,In_470);
nor U2865 (N_2865,In_454,In_1224);
or U2866 (N_2866,In_512,In_820);
or U2867 (N_2867,In_1382,In_899);
nor U2868 (N_2868,In_1062,In_1104);
nand U2869 (N_2869,In_505,In_811);
nor U2870 (N_2870,In_1140,In_195);
nor U2871 (N_2871,In_812,In_1243);
or U2872 (N_2872,In_1196,In_885);
nand U2873 (N_2873,In_651,In_1216);
nor U2874 (N_2874,In_99,In_205);
or U2875 (N_2875,In_365,In_926);
nand U2876 (N_2876,In_562,In_454);
nor U2877 (N_2877,In_1060,In_1169);
or U2878 (N_2878,In_428,In_1480);
and U2879 (N_2879,In_551,In_1216);
and U2880 (N_2880,In_1417,In_889);
nand U2881 (N_2881,In_1203,In_1116);
or U2882 (N_2882,In_215,In_767);
and U2883 (N_2883,In_1065,In_367);
and U2884 (N_2884,In_922,In_493);
and U2885 (N_2885,In_859,In_499);
and U2886 (N_2886,In_449,In_464);
nor U2887 (N_2887,In_1102,In_574);
nand U2888 (N_2888,In_1141,In_756);
and U2889 (N_2889,In_934,In_573);
or U2890 (N_2890,In_601,In_549);
and U2891 (N_2891,In_580,In_573);
and U2892 (N_2892,In_621,In_980);
and U2893 (N_2893,In_718,In_613);
nor U2894 (N_2894,In_1300,In_162);
nor U2895 (N_2895,In_130,In_181);
or U2896 (N_2896,In_676,In_436);
nor U2897 (N_2897,In_895,In_31);
nand U2898 (N_2898,In_1155,In_955);
nor U2899 (N_2899,In_174,In_691);
nor U2900 (N_2900,In_1167,In_689);
or U2901 (N_2901,In_715,In_1123);
nand U2902 (N_2902,In_1086,In_856);
nor U2903 (N_2903,In_491,In_138);
or U2904 (N_2904,In_840,In_124);
and U2905 (N_2905,In_838,In_704);
nand U2906 (N_2906,In_383,In_1096);
or U2907 (N_2907,In_1068,In_651);
and U2908 (N_2908,In_803,In_1439);
and U2909 (N_2909,In_1233,In_897);
and U2910 (N_2910,In_1205,In_1131);
nand U2911 (N_2911,In_731,In_1406);
or U2912 (N_2912,In_797,In_1145);
nand U2913 (N_2913,In_1254,In_549);
or U2914 (N_2914,In_1416,In_1466);
nor U2915 (N_2915,In_1134,In_988);
and U2916 (N_2916,In_1320,In_941);
and U2917 (N_2917,In_527,In_973);
or U2918 (N_2918,In_368,In_602);
or U2919 (N_2919,In_791,In_701);
and U2920 (N_2920,In_884,In_208);
nor U2921 (N_2921,In_846,In_1067);
nand U2922 (N_2922,In_297,In_942);
nor U2923 (N_2923,In_583,In_873);
and U2924 (N_2924,In_1357,In_286);
nor U2925 (N_2925,In_355,In_126);
or U2926 (N_2926,In_585,In_1364);
or U2927 (N_2927,In_99,In_1188);
and U2928 (N_2928,In_350,In_844);
nand U2929 (N_2929,In_1098,In_411);
or U2930 (N_2930,In_427,In_1486);
and U2931 (N_2931,In_539,In_234);
and U2932 (N_2932,In_352,In_1354);
or U2933 (N_2933,In_777,In_1020);
nor U2934 (N_2934,In_1278,In_1004);
and U2935 (N_2935,In_1435,In_1253);
nand U2936 (N_2936,In_699,In_685);
nor U2937 (N_2937,In_990,In_451);
or U2938 (N_2938,In_136,In_106);
or U2939 (N_2939,In_732,In_997);
and U2940 (N_2940,In_855,In_1319);
xnor U2941 (N_2941,In_1413,In_1475);
or U2942 (N_2942,In_1299,In_586);
nor U2943 (N_2943,In_871,In_1256);
nor U2944 (N_2944,In_195,In_1392);
and U2945 (N_2945,In_1260,In_578);
or U2946 (N_2946,In_753,In_713);
or U2947 (N_2947,In_1245,In_1329);
nand U2948 (N_2948,In_148,In_1079);
and U2949 (N_2949,In_1167,In_536);
nand U2950 (N_2950,In_1453,In_411);
nor U2951 (N_2951,In_687,In_668);
and U2952 (N_2952,In_793,In_913);
or U2953 (N_2953,In_43,In_1226);
nor U2954 (N_2954,In_852,In_75);
and U2955 (N_2955,In_1112,In_965);
and U2956 (N_2956,In_1435,In_40);
and U2957 (N_2957,In_1331,In_412);
and U2958 (N_2958,In_470,In_159);
nand U2959 (N_2959,In_1234,In_356);
and U2960 (N_2960,In_1072,In_760);
and U2961 (N_2961,In_497,In_346);
nand U2962 (N_2962,In_1462,In_451);
and U2963 (N_2963,In_248,In_1337);
nand U2964 (N_2964,In_813,In_1013);
and U2965 (N_2965,In_1064,In_253);
and U2966 (N_2966,In_254,In_1034);
nor U2967 (N_2967,In_1146,In_1350);
or U2968 (N_2968,In_270,In_593);
and U2969 (N_2969,In_37,In_1296);
or U2970 (N_2970,In_712,In_433);
or U2971 (N_2971,In_393,In_66);
nor U2972 (N_2972,In_1169,In_221);
or U2973 (N_2973,In_721,In_555);
and U2974 (N_2974,In_41,In_455);
nor U2975 (N_2975,In_380,In_1155);
nand U2976 (N_2976,In_734,In_130);
or U2977 (N_2977,In_1048,In_890);
or U2978 (N_2978,In_555,In_114);
and U2979 (N_2979,In_1156,In_1076);
and U2980 (N_2980,In_1178,In_975);
or U2981 (N_2981,In_273,In_260);
and U2982 (N_2982,In_226,In_405);
nand U2983 (N_2983,In_2,In_811);
nand U2984 (N_2984,In_844,In_1145);
or U2985 (N_2985,In_100,In_424);
and U2986 (N_2986,In_1111,In_798);
nand U2987 (N_2987,In_919,In_406);
nand U2988 (N_2988,In_437,In_345);
or U2989 (N_2989,In_661,In_1201);
nor U2990 (N_2990,In_713,In_488);
nand U2991 (N_2991,In_384,In_1179);
nand U2992 (N_2992,In_872,In_1138);
nor U2993 (N_2993,In_780,In_1067);
nor U2994 (N_2994,In_856,In_432);
or U2995 (N_2995,In_739,In_1148);
nor U2996 (N_2996,In_1311,In_421);
nor U2997 (N_2997,In_1214,In_584);
and U2998 (N_2998,In_302,In_402);
nand U2999 (N_2999,In_704,In_919);
nand U3000 (N_3000,N_1804,N_1941);
xor U3001 (N_3001,N_2367,N_1011);
nand U3002 (N_3002,N_1797,N_2627);
nor U3003 (N_3003,N_2827,N_307);
or U3004 (N_3004,N_258,N_2767);
nor U3005 (N_3005,N_1544,N_2849);
nand U3006 (N_3006,N_1819,N_728);
and U3007 (N_3007,N_1141,N_1813);
nand U3008 (N_3008,N_2904,N_1402);
nand U3009 (N_3009,N_773,N_2118);
nand U3010 (N_3010,N_1571,N_1555);
or U3011 (N_3011,N_2829,N_1421);
nand U3012 (N_3012,N_1768,N_856);
nand U3013 (N_3013,N_1683,N_2355);
nor U3014 (N_3014,N_2582,N_2747);
nor U3015 (N_3015,N_336,N_2759);
or U3016 (N_3016,N_786,N_1973);
nor U3017 (N_3017,N_2839,N_2104);
and U3018 (N_3018,N_1496,N_2326);
or U3019 (N_3019,N_2570,N_2841);
and U3020 (N_3020,N_2261,N_2229);
or U3021 (N_3021,N_1291,N_1138);
and U3022 (N_3022,N_1734,N_2497);
nor U3023 (N_3023,N_2212,N_2375);
nand U3024 (N_3024,N_606,N_790);
nand U3025 (N_3025,N_957,N_1023);
nor U3026 (N_3026,N_1371,N_2821);
nand U3027 (N_3027,N_2672,N_253);
nand U3028 (N_3028,N_919,N_1602);
or U3029 (N_3029,N_1261,N_2132);
nand U3030 (N_3030,N_2708,N_2650);
and U3031 (N_3031,N_1244,N_2880);
nor U3032 (N_3032,N_2310,N_2499);
nor U3033 (N_3033,N_1993,N_114);
nor U3034 (N_3034,N_941,N_690);
nand U3035 (N_3035,N_635,N_886);
and U3036 (N_3036,N_842,N_1039);
nand U3037 (N_3037,N_371,N_460);
nor U3038 (N_3038,N_2577,N_399);
or U3039 (N_3039,N_2642,N_303);
or U3040 (N_3040,N_1445,N_1056);
nand U3041 (N_3041,N_2282,N_2308);
or U3042 (N_3042,N_16,N_580);
nand U3043 (N_3043,N_2381,N_392);
or U3044 (N_3044,N_1466,N_1652);
or U3045 (N_3045,N_48,N_722);
nand U3046 (N_3046,N_747,N_202);
nor U3047 (N_3047,N_1034,N_2750);
nand U3048 (N_3048,N_1902,N_1213);
or U3049 (N_3049,N_1552,N_1562);
nand U3050 (N_3050,N_697,N_1416);
and U3051 (N_3051,N_1324,N_311);
nand U3052 (N_3052,N_1367,N_933);
nor U3053 (N_3053,N_2875,N_2848);
nand U3054 (N_3054,N_907,N_1438);
nor U3055 (N_3055,N_2241,N_1137);
or U3056 (N_3056,N_2438,N_1358);
and U3057 (N_3057,N_1300,N_2309);
or U3058 (N_3058,N_2193,N_1456);
and U3059 (N_3059,N_242,N_1986);
or U3060 (N_3060,N_818,N_1968);
and U3061 (N_3061,N_776,N_2316);
nand U3062 (N_3062,N_1014,N_1925);
and U3063 (N_3063,N_2624,N_2909);
or U3064 (N_3064,N_2536,N_1432);
nand U3065 (N_3065,N_2518,N_2723);
nand U3066 (N_3066,N_2244,N_270);
or U3067 (N_3067,N_2539,N_463);
nor U3068 (N_3068,N_596,N_1999);
or U3069 (N_3069,N_548,N_2973);
or U3070 (N_3070,N_1297,N_2288);
xnor U3071 (N_3071,N_2145,N_372);
nand U3072 (N_3072,N_2083,N_444);
or U3073 (N_3073,N_837,N_2558);
nand U3074 (N_3074,N_2034,N_19);
or U3075 (N_3075,N_479,N_508);
nor U3076 (N_3076,N_2555,N_1911);
and U3077 (N_3077,N_874,N_2891);
nand U3078 (N_3078,N_1543,N_288);
nand U3079 (N_3079,N_1210,N_1946);
nand U3080 (N_3080,N_1910,N_1181);
nor U3081 (N_3081,N_2311,N_1994);
nor U3082 (N_3082,N_2784,N_2760);
nand U3083 (N_3083,N_1679,N_404);
nor U3084 (N_3084,N_601,N_589);
and U3085 (N_3085,N_1712,N_2632);
and U3086 (N_3086,N_939,N_2325);
or U3087 (N_3087,N_86,N_1092);
or U3088 (N_3088,N_2961,N_2005);
nand U3089 (N_3089,N_1388,N_1448);
nor U3090 (N_3090,N_2385,N_1059);
or U3091 (N_3091,N_2575,N_588);
or U3092 (N_3092,N_1954,N_2303);
nand U3093 (N_3093,N_2836,N_2087);
nand U3094 (N_3094,N_1126,N_2060);
nand U3095 (N_3095,N_2078,N_2675);
nand U3096 (N_3096,N_1006,N_2562);
and U3097 (N_3097,N_2520,N_2307);
and U3098 (N_3098,N_1451,N_1807);
nand U3099 (N_3099,N_2274,N_1969);
or U3100 (N_3100,N_2948,N_687);
nand U3101 (N_3101,N_2994,N_2787);
nor U3102 (N_3102,N_96,N_2894);
and U3103 (N_3103,N_1614,N_1470);
and U3104 (N_3104,N_1714,N_1403);
nor U3105 (N_3105,N_2015,N_1453);
nor U3106 (N_3106,N_781,N_1333);
and U3107 (N_3107,N_1391,N_2055);
and U3108 (N_3108,N_1121,N_1425);
nand U3109 (N_3109,N_2442,N_844);
and U3110 (N_3110,N_1334,N_2062);
nor U3111 (N_3111,N_2801,N_969);
and U3112 (N_3112,N_2924,N_1338);
nand U3113 (N_3113,N_2548,N_1839);
and U3114 (N_3114,N_1695,N_1878);
nor U3115 (N_3115,N_2870,N_2168);
or U3116 (N_3116,N_797,N_1662);
nor U3117 (N_3117,N_1017,N_488);
nor U3118 (N_3118,N_2815,N_1145);
or U3119 (N_3119,N_1251,N_2342);
and U3120 (N_3120,N_988,N_2082);
and U3121 (N_3121,N_1109,N_2323);
nand U3122 (N_3122,N_1701,N_843);
nand U3123 (N_3123,N_2987,N_2211);
nand U3124 (N_3124,N_2895,N_2446);
and U3125 (N_3125,N_953,N_1236);
and U3126 (N_3126,N_1361,N_1444);
or U3127 (N_3127,N_1579,N_1962);
nand U3128 (N_3128,N_2882,N_1634);
xor U3129 (N_3129,N_252,N_2175);
nand U3130 (N_3130,N_2450,N_1755);
nor U3131 (N_3131,N_986,N_1147);
nand U3132 (N_3132,N_1206,N_1215);
nand U3133 (N_3133,N_1085,N_1200);
or U3134 (N_3134,N_2187,N_1867);
or U3135 (N_3135,N_2739,N_1676);
nand U3136 (N_3136,N_2532,N_2661);
nor U3137 (N_3137,N_2471,N_1142);
and U3138 (N_3138,N_2741,N_2724);
and U3139 (N_3139,N_1276,N_1531);
and U3140 (N_3140,N_1103,N_2706);
and U3141 (N_3141,N_902,N_956);
and U3142 (N_3142,N_334,N_1664);
and U3143 (N_3143,N_1742,N_1033);
and U3144 (N_3144,N_1196,N_1952);
and U3145 (N_3145,N_474,N_1417);
or U3146 (N_3146,N_1263,N_2028);
or U3147 (N_3147,N_2235,N_2863);
nand U3148 (N_3148,N_1616,N_1754);
nor U3149 (N_3149,N_891,N_2406);
and U3150 (N_3150,N_195,N_881);
and U3151 (N_3151,N_2547,N_1331);
and U3152 (N_3152,N_2596,N_1524);
nand U3153 (N_3153,N_2720,N_350);
or U3154 (N_3154,N_1259,N_2778);
xor U3155 (N_3155,N_299,N_5);
and U3156 (N_3156,N_2253,N_435);
and U3157 (N_3157,N_2692,N_2172);
nor U3158 (N_3158,N_2958,N_1098);
or U3159 (N_3159,N_2588,N_87);
nand U3160 (N_3160,N_771,N_1390);
nand U3161 (N_3161,N_2594,N_2379);
and U3162 (N_3162,N_1897,N_1711);
or U3163 (N_3163,N_897,N_2368);
xnor U3164 (N_3164,N_2484,N_1239);
or U3165 (N_3165,N_591,N_2862);
and U3166 (N_3166,N_794,N_414);
nor U3167 (N_3167,N_1314,N_2736);
and U3168 (N_3168,N_379,N_851);
or U3169 (N_3169,N_424,N_1406);
nor U3170 (N_3170,N_678,N_2176);
nand U3171 (N_3171,N_1180,N_155);
or U3172 (N_3172,N_1189,N_181);
or U3173 (N_3173,N_1904,N_2737);
or U3174 (N_3174,N_332,N_623);
and U3175 (N_3175,N_1736,N_2744);
nor U3176 (N_3176,N_485,N_1356);
nand U3177 (N_3177,N_137,N_70);
nand U3178 (N_3178,N_2731,N_654);
or U3179 (N_3179,N_216,N_1503);
nor U3180 (N_3180,N_1975,N_38);
nand U3181 (N_3181,N_2441,N_621);
or U3182 (N_3182,N_396,N_339);
or U3183 (N_3183,N_1942,N_4);
nor U3184 (N_3184,N_2237,N_1928);
nand U3185 (N_3185,N_22,N_849);
nand U3186 (N_3186,N_207,N_324);
or U3187 (N_3187,N_639,N_1667);
nand U3188 (N_3188,N_2873,N_2592);
nand U3189 (N_3189,N_2398,N_1895);
and U3190 (N_3190,N_867,N_602);
or U3191 (N_3191,N_1534,N_21);
or U3192 (N_3192,N_2141,N_2581);
nand U3193 (N_3193,N_520,N_511);
and U3194 (N_3194,N_43,N_373);
nand U3195 (N_3195,N_173,N_2860);
nand U3196 (N_3196,N_600,N_2722);
and U3197 (N_3197,N_1468,N_276);
and U3198 (N_3198,N_2792,N_2170);
and U3199 (N_3199,N_2197,N_132);
nor U3200 (N_3200,N_2046,N_2437);
nor U3201 (N_3201,N_1112,N_2667);
and U3202 (N_3202,N_2640,N_1328);
or U3203 (N_3203,N_0,N_1685);
and U3204 (N_3204,N_186,N_2324);
xnor U3205 (N_3205,N_1963,N_920);
and U3206 (N_3206,N_2139,N_1364);
nand U3207 (N_3207,N_198,N_2267);
nor U3208 (N_3208,N_2803,N_145);
or U3209 (N_3209,N_2469,N_2299);
nand U3210 (N_3210,N_1646,N_2344);
and U3211 (N_3211,N_121,N_1709);
nand U3212 (N_3212,N_971,N_572);
nor U3213 (N_3213,N_934,N_734);
and U3214 (N_3214,N_1791,N_1829);
nand U3215 (N_3215,N_323,N_1723);
and U3216 (N_3216,N_2550,N_605);
and U3217 (N_3217,N_2298,N_1788);
or U3218 (N_3218,N_2492,N_1392);
or U3219 (N_3219,N_1221,N_598);
nor U3220 (N_3220,N_2430,N_1461);
or U3221 (N_3221,N_177,N_2833);
nand U3222 (N_3222,N_88,N_1855);
nand U3223 (N_3223,N_2579,N_1158);
nor U3224 (N_3224,N_221,N_80);
nor U3225 (N_3225,N_1281,N_2522);
or U3226 (N_3226,N_1865,N_2766);
or U3227 (N_3227,N_812,N_1735);
nand U3228 (N_3228,N_889,N_1572);
nand U3229 (N_3229,N_468,N_2589);
nor U3230 (N_3230,N_2352,N_2651);
and U3231 (N_3231,N_2854,N_1386);
or U3232 (N_3232,N_65,N_1738);
and U3233 (N_3233,N_487,N_2847);
nor U3234 (N_3234,N_866,N_397);
or U3235 (N_3235,N_2341,N_142);
nor U3236 (N_3236,N_1615,N_2729);
and U3237 (N_3237,N_2630,N_2656);
nand U3238 (N_3238,N_2066,N_1009);
nand U3239 (N_3239,N_1107,N_811);
nand U3240 (N_3240,N_293,N_1192);
or U3241 (N_3241,N_73,N_394);
or U3242 (N_3242,N_2531,N_1316);
and U3243 (N_3243,N_1363,N_2916);
xnor U3244 (N_3244,N_1677,N_657);
xor U3245 (N_3245,N_213,N_2923);
nand U3246 (N_3246,N_2752,N_1506);
nor U3247 (N_3247,N_2049,N_1686);
or U3248 (N_3248,N_1163,N_633);
and U3249 (N_3249,N_2151,N_532);
and U3250 (N_3250,N_854,N_1258);
nand U3251 (N_3251,N_829,N_1832);
nand U3252 (N_3252,N_237,N_1565);
or U3253 (N_3253,N_449,N_2043);
nor U3254 (N_3254,N_523,N_2042);
or U3255 (N_3255,N_2888,N_2611);
nand U3256 (N_3256,N_1280,N_69);
nand U3257 (N_3257,N_1597,N_1341);
or U3258 (N_3258,N_1015,N_1117);
nor U3259 (N_3259,N_2421,N_536);
or U3260 (N_3260,N_15,N_2514);
nor U3261 (N_3261,N_617,N_2972);
nor U3262 (N_3262,N_774,N_2200);
or U3263 (N_3263,N_2691,N_501);
nor U3264 (N_3264,N_1640,N_164);
and U3265 (N_3265,N_1326,N_3);
or U3266 (N_3266,N_451,N_2655);
nand U3267 (N_3267,N_2440,N_1607);
or U3268 (N_3268,N_302,N_1576);
nand U3269 (N_3269,N_2432,N_101);
or U3270 (N_3270,N_1294,N_2559);
or U3271 (N_3271,N_665,N_354);
or U3272 (N_3272,N_835,N_1970);
and U3273 (N_3273,N_2830,N_567);
or U3274 (N_3274,N_2802,N_1484);
nand U3275 (N_3275,N_1332,N_2563);
and U3276 (N_3276,N_402,N_1810);
nor U3277 (N_3277,N_923,N_2992);
and U3278 (N_3278,N_2807,N_1439);
and U3279 (N_3279,N_461,N_1250);
and U3280 (N_3280,N_1449,N_2707);
nand U3281 (N_3281,N_1757,N_808);
or U3282 (N_3282,N_2897,N_2333);
and U3283 (N_3283,N_2872,N_767);
and U3284 (N_3284,N_1146,N_1493);
and U3285 (N_3285,N_1004,N_2881);
and U3286 (N_3286,N_499,N_1474);
nand U3287 (N_3287,N_1826,N_2728);
nand U3288 (N_3288,N_2865,N_766);
or U3289 (N_3289,N_13,N_2063);
and U3290 (N_3290,N_405,N_1477);
or U3291 (N_3291,N_2601,N_1708);
or U3292 (N_3292,N_83,N_1778);
or U3293 (N_3293,N_709,N_421);
or U3294 (N_3294,N_2826,N_2297);
nor U3295 (N_3295,N_860,N_2521);
and U3296 (N_3296,N_973,N_356);
nor U3297 (N_3297,N_319,N_892);
nand U3298 (N_3298,N_2657,N_1);
and U3299 (N_3299,N_1834,N_1564);
and U3300 (N_3300,N_2733,N_1949);
and U3301 (N_3301,N_2052,N_2387);
or U3302 (N_3302,N_1990,N_282);
and U3303 (N_3303,N_2604,N_1266);
or U3304 (N_3304,N_1434,N_1007);
nor U3305 (N_3305,N_1995,N_2705);
nor U3306 (N_3306,N_2101,N_2491);
and U3307 (N_3307,N_315,N_440);
nor U3308 (N_3308,N_2753,N_93);
or U3309 (N_3309,N_1610,N_1197);
and U3310 (N_3310,N_2250,N_441);
nor U3311 (N_3311,N_2969,N_925);
nor U3312 (N_3312,N_2302,N_400);
nor U3313 (N_3313,N_2340,N_2209);
or U3314 (N_3314,N_248,N_870);
and U3315 (N_3315,N_732,N_2931);
and U3316 (N_3316,N_1773,N_1859);
and U3317 (N_3317,N_2294,N_1162);
nand U3318 (N_3318,N_1177,N_954);
nand U3319 (N_3319,N_158,N_62);
nor U3320 (N_3320,N_984,N_498);
nand U3321 (N_3321,N_1872,N_1921);
nand U3322 (N_3322,N_267,N_2996);
nor U3323 (N_3323,N_2852,N_427);
nor U3324 (N_3324,N_2029,N_1959);
and U3325 (N_3325,N_1852,N_586);
or U3326 (N_3326,N_510,N_582);
and U3327 (N_3327,N_916,N_1526);
nor U3328 (N_3328,N_91,N_2265);
nand U3329 (N_3329,N_668,N_2735);
or U3330 (N_3330,N_317,N_702);
nand U3331 (N_3331,N_1856,N_1527);
or U3332 (N_3332,N_587,N_2730);
or U3333 (N_3333,N_2415,N_557);
nor U3334 (N_3334,N_2781,N_1613);
nand U3335 (N_3335,N_2813,N_2293);
nor U3336 (N_3336,N_2444,N_661);
or U3337 (N_3337,N_68,N_1900);
nand U3338 (N_3338,N_862,N_117);
nor U3339 (N_3339,N_1149,N_219);
or U3340 (N_3340,N_1397,N_1948);
or U3341 (N_3341,N_2757,N_140);
and U3342 (N_3342,N_2384,N_2866);
nand U3343 (N_3343,N_2050,N_272);
and U3344 (N_3344,N_1937,N_2107);
or U3345 (N_3345,N_1249,N_286);
and U3346 (N_3346,N_955,N_991);
nand U3347 (N_3347,N_2892,N_977);
nor U3348 (N_3348,N_1716,N_1498);
or U3349 (N_3349,N_1557,N_1270);
nand U3350 (N_3350,N_2185,N_431);
nand U3351 (N_3351,N_749,N_1310);
nor U3352 (N_3352,N_1411,N_692);
and U3353 (N_3353,N_1520,N_1471);
or U3354 (N_3354,N_1026,N_470);
nor U3355 (N_3355,N_2633,N_249);
and U3356 (N_3356,N_1751,N_2806);
and U3357 (N_3357,N_2037,N_2603);
nand U3358 (N_3358,N_935,N_348);
and U3359 (N_3359,N_1670,N_2997);
and U3360 (N_3360,N_1956,N_800);
nand U3361 (N_3361,N_644,N_1288);
nand U3362 (N_3362,N_2424,N_660);
or U3363 (N_3363,N_2966,N_693);
or U3364 (N_3364,N_1871,N_2179);
nor U3365 (N_3365,N_1873,N_1737);
and U3366 (N_3366,N_200,N_2800);
nand U3367 (N_3367,N_318,N_1337);
or U3368 (N_3368,N_2779,N_1671);
nor U3369 (N_3369,N_585,N_231);
or U3370 (N_3370,N_187,N_1187);
and U3371 (N_3371,N_2144,N_1118);
or U3372 (N_3372,N_2869,N_2004);
nand U3373 (N_3373,N_1972,N_1611);
or U3374 (N_3374,N_1508,N_2554);
xnor U3375 (N_3375,N_574,N_741);
or U3376 (N_3376,N_570,N_1798);
nand U3377 (N_3377,N_465,N_2071);
nor U3378 (N_3378,N_2980,N_107);
and U3379 (N_3379,N_1849,N_2912);
nor U3380 (N_3380,N_278,N_2478);
nor U3381 (N_3381,N_215,N_1499);
nor U3382 (N_3382,N_2528,N_1379);
or U3383 (N_3383,N_848,N_2962);
or U3384 (N_3384,N_552,N_1581);
nor U3385 (N_3385,N_1978,N_1626);
nor U3386 (N_3386,N_1786,N_2067);
and U3387 (N_3387,N_24,N_1374);
nand U3388 (N_3388,N_1580,N_2164);
and U3389 (N_3389,N_445,N_1772);
nand U3390 (N_3390,N_30,N_352);
nand U3391 (N_3391,N_2669,N_1428);
nor U3392 (N_3392,N_1269,N_736);
nand U3393 (N_3393,N_130,N_1167);
nor U3394 (N_3394,N_172,N_2534);
and U3395 (N_3395,N_1024,N_2116);
nor U3396 (N_3396,N_1600,N_2845);
and U3397 (N_3397,N_1050,N_1702);
nand U3398 (N_3398,N_224,N_2496);
or U3399 (N_3399,N_2190,N_2191);
or U3400 (N_3400,N_2758,N_1784);
nand U3401 (N_3401,N_1424,N_937);
nor U3402 (N_3402,N_2631,N_1894);
nand U3403 (N_3403,N_1035,N_2954);
nor U3404 (N_3404,N_2089,N_1431);
nor U3405 (N_3405,N_1715,N_2161);
nand U3406 (N_3406,N_2339,N_2889);
nor U3407 (N_3407,N_2449,N_430);
or U3408 (N_3408,N_491,N_559);
and U3409 (N_3409,N_2405,N_1143);
nor U3410 (N_3410,N_1789,N_1814);
and U3411 (N_3411,N_375,N_1020);
nor U3412 (N_3412,N_2156,N_456);
and U3413 (N_3413,N_1522,N_2468);
nor U3414 (N_3414,N_2743,N_2018);
or U3415 (N_3415,N_929,N_2016);
and U3416 (N_3416,N_1380,N_2138);
or U3417 (N_3417,N_711,N_551);
or U3418 (N_3418,N_2347,N_545);
and U3419 (N_3419,N_2649,N_2192);
nand U3420 (N_3420,N_1642,N_2218);
nor U3421 (N_3421,N_351,N_2359);
nand U3422 (N_3422,N_139,N_2686);
and U3423 (N_3423,N_201,N_2431);
or U3424 (N_3424,N_154,N_255);
nor U3425 (N_3425,N_2354,N_2003);
and U3426 (N_3426,N_921,N_1512);
nand U3427 (N_3427,N_1212,N_2);
and U3428 (N_3428,N_1663,N_964);
and U3429 (N_3429,N_1822,N_761);
and U3430 (N_3430,N_2552,N_1689);
nor U3431 (N_3431,N_2755,N_1229);
and U3432 (N_3432,N_772,N_2930);
nand U3433 (N_3433,N_129,N_1160);
or U3434 (N_3434,N_368,N_2915);
and U3435 (N_3435,N_787,N_824);
or U3436 (N_3436,N_648,N_2628);
nor U3437 (N_3437,N_2305,N_1560);
or U3438 (N_3438,N_2762,N_1880);
or U3439 (N_3439,N_967,N_1489);
and U3440 (N_3440,N_2328,N_2911);
or U3441 (N_3441,N_157,N_2266);
nor U3442 (N_3442,N_1286,N_719);
or U3443 (N_3443,N_1985,N_2740);
nand U3444 (N_3444,N_2986,N_1760);
nand U3445 (N_3445,N_847,N_2843);
nor U3446 (N_3446,N_46,N_2998);
nor U3447 (N_3447,N_1981,N_2751);
nand U3448 (N_3448,N_2887,N_806);
or U3449 (N_3449,N_1152,N_1843);
and U3450 (N_3450,N_2634,N_578);
nand U3451 (N_3451,N_1623,N_316);
and U3452 (N_3452,N_1185,N_417);
or U3453 (N_3453,N_320,N_553);
and U3454 (N_3454,N_1809,N_656);
and U3455 (N_3455,N_1070,N_1119);
nor U3456 (N_3456,N_529,N_1290);
or U3457 (N_3457,N_2685,N_85);
or U3458 (N_3458,N_1365,N_390);
or U3459 (N_3459,N_575,N_2702);
and U3460 (N_3460,N_533,N_1964);
nor U3461 (N_3461,N_1758,N_2689);
and U3462 (N_3462,N_2117,N_2977);
nand U3463 (N_3463,N_974,N_2745);
nand U3464 (N_3464,N_1785,N_555);
nor U3465 (N_3465,N_2360,N_2959);
xnor U3466 (N_3466,N_2402,N_539);
nand U3467 (N_3467,N_2734,N_1087);
nand U3468 (N_3468,N_698,N_2975);
nand U3469 (N_3469,N_2590,N_2726);
nor U3470 (N_3470,N_1150,N_2622);
nor U3471 (N_3471,N_2597,N_1874);
nor U3472 (N_3472,N_489,N_484);
nand U3473 (N_3473,N_29,N_238);
and U3474 (N_3474,N_344,N_667);
or U3475 (N_3475,N_1818,N_915);
or U3476 (N_3476,N_357,N_2495);
nor U3477 (N_3477,N_810,N_2804);
or U3478 (N_3478,N_1277,N_128);
and U3479 (N_3479,N_949,N_1165);
and U3480 (N_3480,N_611,N_31);
xor U3481 (N_3481,N_2228,N_1260);
and U3482 (N_3482,N_2465,N_2782);
or U3483 (N_3483,N_314,N_443);
nor U3484 (N_3484,N_863,N_740);
nor U3485 (N_3485,N_1605,N_494);
and U3486 (N_3486,N_2527,N_642);
nand U3487 (N_3487,N_1114,N_2128);
nor U3488 (N_3488,N_2537,N_197);
nand U3489 (N_3489,N_1621,N_718);
nand U3490 (N_3490,N_2814,N_903);
nor U3491 (N_3491,N_377,N_1120);
or U3492 (N_3492,N_1031,N_161);
nor U3493 (N_3493,N_2868,N_1123);
nand U3494 (N_3494,N_1974,N_2719);
nor U3495 (N_3495,N_212,N_2697);
nor U3496 (N_3496,N_1648,N_2572);
nand U3497 (N_3497,N_1336,N_2125);
and U3498 (N_3498,N_170,N_2797);
nand U3499 (N_3499,N_1222,N_1319);
and U3500 (N_3500,N_1209,N_2893);
or U3501 (N_3501,N_1838,N_2607);
nor U3502 (N_3502,N_1528,N_2971);
nor U3503 (N_3503,N_2248,N_691);
nor U3504 (N_3504,N_2223,N_229);
and U3505 (N_3505,N_1226,N_614);
or U3506 (N_3506,N_1530,N_1651);
nor U3507 (N_3507,N_2383,N_2131);
or U3508 (N_3508,N_2350,N_569);
and U3509 (N_3509,N_1776,N_852);
or U3510 (N_3510,N_2490,N_176);
and U3511 (N_3511,N_45,N_2382);
and U3512 (N_3512,N_2525,N_2059);
nand U3513 (N_3513,N_655,N_1110);
nand U3514 (N_3514,N_1061,N_2903);
nand U3515 (N_3515,N_2024,N_2487);
or U3516 (N_3516,N_1780,N_688);
and U3517 (N_3517,N_2798,N_2370);
and U3518 (N_3518,N_1960,N_680);
or U3519 (N_3519,N_2045,N_2819);
nand U3520 (N_3520,N_653,N_2162);
nor U3521 (N_3521,N_2785,N_2203);
or U3522 (N_3522,N_2306,N_2252);
and U3523 (N_3523,N_777,N_2940);
nand U3524 (N_3524,N_2098,N_42);
or U3525 (N_3525,N_2166,N_2304);
nor U3526 (N_3526,N_832,N_1984);
nor U3527 (N_3527,N_483,N_1179);
xnor U3528 (N_3528,N_1546,N_261);
and U3529 (N_3529,N_751,N_1279);
and U3530 (N_3530,N_2153,N_813);
and U3531 (N_3531,N_151,N_946);
nand U3532 (N_3532,N_2716,N_2748);
or U3533 (N_3533,N_770,N_1299);
nand U3534 (N_3534,N_839,N_2789);
or U3535 (N_3535,N_1746,N_1824);
or U3536 (N_3536,N_289,N_2953);
nor U3537 (N_3537,N_2113,N_757);
and U3538 (N_3538,N_1548,N_2428);
nand U3539 (N_3539,N_541,N_1054);
nor U3540 (N_3540,N_1161,N_1745);
or U3541 (N_3541,N_2985,N_960);
or U3542 (N_3542,N_2565,N_2772);
nand U3543 (N_3543,N_2538,N_226);
nor U3544 (N_3544,N_1140,N_1485);
or U3545 (N_3545,N_2617,N_8);
nand U3546 (N_3546,N_1382,N_1647);
nor U3547 (N_3547,N_1377,N_1016);
or U3548 (N_3548,N_1684,N_2600);
or U3549 (N_3549,N_2680,N_1883);
and U3550 (N_3550,N_715,N_2378);
nand U3551 (N_3551,N_1488,N_1099);
or U3552 (N_3552,N_2717,N_1877);
or U3553 (N_3553,N_1944,N_1084);
nand U3554 (N_3554,N_1398,N_266);
or U3555 (N_3555,N_883,N_1455);
or U3556 (N_3556,N_2074,N_707);
nor U3557 (N_3557,N_2917,N_47);
nor U3558 (N_3558,N_2557,N_95);
and U3559 (N_3559,N_855,N_1131);
nor U3560 (N_3560,N_1182,N_183);
and U3561 (N_3561,N_244,N_296);
nor U3562 (N_3562,N_2913,N_819);
or U3563 (N_3563,N_2455,N_2900);
nor U3564 (N_3564,N_2380,N_1917);
nand U3565 (N_3565,N_133,N_1096);
nor U3566 (N_3566,N_1979,N_2859);
nor U3567 (N_3567,N_2837,N_401);
or U3568 (N_3568,N_1452,N_2287);
nand U3569 (N_3569,N_958,N_178);
or U3570 (N_3570,N_2436,N_795);
nand U3571 (N_3571,N_223,N_1047);
or U3572 (N_3572,N_1203,N_663);
nor U3573 (N_3573,N_1139,N_876);
nand U3574 (N_3574,N_2505,N_2115);
and U3575 (N_3575,N_534,N_428);
and U3576 (N_3576,N_674,N_1368);
or U3577 (N_3577,N_1036,N_917);
nand U3578 (N_3578,N_525,N_169);
nand U3579 (N_3579,N_2974,N_2535);
or U3580 (N_3580,N_2693,N_2317);
nand U3581 (N_3581,N_1583,N_2159);
and U3582 (N_3582,N_1346,N_1312);
and U3583 (N_3583,N_2277,N_1174);
or U3584 (N_3584,N_2593,N_597);
or U3585 (N_3585,N_234,N_560);
and U3586 (N_3586,N_2206,N_2754);
nand U3587 (N_3587,N_1081,N_126);
nor U3588 (N_3588,N_2182,N_1966);
and U3589 (N_3589,N_1835,N_2599);
nand U3590 (N_3590,N_2613,N_2770);
nand U3591 (N_3591,N_2701,N_2944);
or U3592 (N_3592,N_84,N_645);
or U3593 (N_3593,N_1350,N_12);
or U3594 (N_3594,N_2205,N_2439);
and U3595 (N_3595,N_2510,N_884);
nand U3596 (N_3596,N_846,N_2319);
nor U3597 (N_3597,N_2541,N_2158);
nand U3598 (N_3598,N_664,N_2929);
or U3599 (N_3599,N_2279,N_2371);
nor U3600 (N_3600,N_1062,N_815);
or U3601 (N_3601,N_2566,N_1915);
nand U3602 (N_3602,N_1408,N_981);
or U3603 (N_3603,N_1321,N_2687);
and U3604 (N_3604,N_2818,N_2610);
and U3605 (N_3605,N_1068,N_2756);
or U3606 (N_3606,N_341,N_845);
and U3607 (N_3607,N_1644,N_454);
and U3608 (N_3608,N_2173,N_1638);
nand U3609 (N_3609,N_2982,N_1658);
nand U3610 (N_3610,N_64,N_230);
and U3611 (N_3611,N_144,N_1933);
nor U3612 (N_3612,N_2918,N_2318);
and U3613 (N_3613,N_1055,N_2102);
and U3614 (N_3614,N_232,N_1044);
nor U3615 (N_3615,N_1327,N_1436);
and U3616 (N_3616,N_1690,N_1752);
nand U3617 (N_3617,N_947,N_1858);
or U3618 (N_3618,N_1559,N_1584);
nand U3619 (N_3619,N_637,N_1799);
and U3620 (N_3620,N_1577,N_134);
or U3621 (N_3621,N_1609,N_28);
or U3622 (N_3622,N_163,N_2264);
or U3623 (N_3623,N_1665,N_793);
nand U3624 (N_3624,N_1899,N_1262);
nor U3625 (N_3625,N_993,N_2453);
nor U3626 (N_3626,N_60,N_2199);
or U3627 (N_3627,N_1385,N_2092);
nor U3628 (N_3628,N_2242,N_149);
and U3629 (N_3629,N_1935,N_2216);
nand U3630 (N_3630,N_1636,N_1650);
and U3631 (N_3631,N_2896,N_2967);
or U3632 (N_3632,N_2636,N_1396);
nand U3633 (N_3633,N_983,N_2952);
nor U3634 (N_3634,N_828,N_1256);
nand U3635 (N_3635,N_2585,N_2470);
nand U3636 (N_3636,N_2411,N_1443);
nand U3637 (N_3637,N_1298,N_74);
and U3638 (N_3638,N_1514,N_2844);
or U3639 (N_3639,N_2676,N_873);
nor U3640 (N_3640,N_679,N_2433);
xor U3641 (N_3641,N_1971,N_2713);
nor U3642 (N_3642,N_189,N_1082);
xor U3643 (N_3643,N_730,N_2659);
or U3644 (N_3644,N_2910,N_2703);
nand U3645 (N_3645,N_486,N_1292);
nor U3646 (N_3646,N_2425,N_1558);
nor U3647 (N_3647,N_807,N_2479);
nand U3648 (N_3648,N_2885,N_2993);
or U3649 (N_3649,N_609,N_634);
nand U3650 (N_3650,N_1657,N_995);
and U3651 (N_3651,N_549,N_2991);
and U3652 (N_3652,N_1048,N_1487);
and U3653 (N_3653,N_2937,N_658);
nor U3654 (N_3654,N_1344,N_2409);
nand U3655 (N_3655,N_1569,N_1483);
nor U3656 (N_3656,N_447,N_1501);
nand U3657 (N_3657,N_1028,N_513);
nand U3658 (N_3658,N_1698,N_931);
nand U3659 (N_3659,N_522,N_98);
nand U3660 (N_3660,N_938,N_1617);
nor U3661 (N_3661,N_206,N_416);
nand U3662 (N_3662,N_2561,N_1729);
or U3663 (N_3663,N_975,N_558);
and U3664 (N_3664,N_1914,N_1705);
or U3665 (N_3665,N_759,N_1549);
nor U3666 (N_3666,N_285,N_2452);
nand U3667 (N_3667,N_6,N_1673);
or U3668 (N_3668,N_1171,N_2808);
nand U3669 (N_3669,N_2926,N_821);
nand U3670 (N_3670,N_566,N_1248);
nand U3671 (N_3671,N_274,N_335);
nand U3672 (N_3672,N_2738,N_2867);
xor U3673 (N_3673,N_1076,N_300);
and U3674 (N_3674,N_407,N_1604);
nor U3675 (N_3675,N_2513,N_214);
nor U3676 (N_3676,N_2461,N_1481);
nor U3677 (N_3677,N_950,N_1101);
or U3678 (N_3678,N_49,N_1500);
nand U3679 (N_3679,N_2677,N_2472);
nor U3680 (N_3680,N_725,N_564);
nand U3681 (N_3681,N_2774,N_321);
or U3682 (N_3682,N_2070,N_275);
and U3683 (N_3683,N_895,N_433);
and U3684 (N_3684,N_1864,N_801);
or U3685 (N_3685,N_612,N_481);
nand U3686 (N_3686,N_409,N_387);
nand U3687 (N_3687,N_573,N_263);
nand U3688 (N_3688,N_738,N_1366);
nor U3689 (N_3689,N_1717,N_2167);
or U3690 (N_3690,N_325,N_864);
or U3691 (N_3691,N_1870,N_1653);
and U3692 (N_3692,N_1243,N_2908);
and U3693 (N_3693,N_378,N_1151);
nor U3694 (N_3694,N_2445,N_713);
or U3695 (N_3695,N_446,N_890);
nand U3696 (N_3696,N_217,N_2508);
nand U3697 (N_3697,N_2517,N_1929);
nand U3698 (N_3698,N_2823,N_987);
nor U3699 (N_3699,N_75,N_438);
nand U3700 (N_3700,N_1214,N_432);
nand U3701 (N_3701,N_2155,N_2856);
nand U3702 (N_3702,N_1507,N_2286);
xnor U3703 (N_3703,N_1509,N_2811);
nor U3704 (N_3704,N_53,N_301);
or U3705 (N_3705,N_2777,N_2956);
nor U3706 (N_3706,N_677,N_768);
and U3707 (N_3707,N_391,N_442);
or U3708 (N_3708,N_2876,N_23);
or U3709 (N_3709,N_2048,N_670);
nor U3710 (N_3710,N_2690,N_742);
nor U3711 (N_3711,N_1790,N_2320);
nand U3712 (N_3712,N_415,N_1726);
and U3713 (N_3713,N_1223,N_472);
and U3714 (N_3714,N_904,N_2553);
or U3715 (N_3715,N_1775,N_1885);
and U3716 (N_3716,N_1342,N_2389);
or U3717 (N_3717,N_518,N_2506);
nor U3718 (N_3718,N_1596,N_1907);
or U3719 (N_3719,N_2256,N_2204);
nor U3720 (N_3720,N_1733,N_35);
xnor U3721 (N_3721,N_148,N_1064);
nand U3722 (N_3722,N_2044,N_2725);
nand U3723 (N_3723,N_419,N_999);
nor U3724 (N_3724,N_168,N_458);
nand U3725 (N_3725,N_1144,N_1598);
and U3726 (N_3726,N_826,N_2143);
or U3727 (N_3727,N_1924,N_1517);
or U3728 (N_3728,N_1624,N_343);
or U3729 (N_3729,N_1802,N_1265);
nand U3730 (N_3730,N_1713,N_1043);
nand U3731 (N_3731,N_240,N_2871);
nor U3732 (N_3732,N_827,N_188);
or U3733 (N_3733,N_2919,N_1491);
nand U3734 (N_3734,N_452,N_705);
nand U3735 (N_3735,N_2400,N_2369);
and U3736 (N_3736,N_604,N_1127);
or U3737 (N_3737,N_1010,N_2095);
or U3738 (N_3738,N_853,N_1351);
and U3739 (N_3739,N_1282,N_2221);
nand U3740 (N_3740,N_1207,N_2855);
nor U3741 (N_3741,N_1926,N_1052);
or U3742 (N_3742,N_1619,N_1739);
nor U3743 (N_3743,N_14,N_733);
and U3744 (N_3744,N_2120,N_56);
or U3745 (N_3745,N_1817,N_783);
and U3746 (N_3746,N_227,N_1862);
nand U3747 (N_3747,N_500,N_1821);
nor U3748 (N_3748,N_72,N_1513);
nor U3749 (N_3749,N_1612,N_834);
nand U3750 (N_3750,N_1857,N_2451);
and U3751 (N_3751,N_54,N_2335);
or U3752 (N_3752,N_517,N_210);
nand U3753 (N_3753,N_649,N_1108);
nor U3754 (N_3754,N_882,N_2002);
nor U3755 (N_3755,N_1720,N_712);
nor U3756 (N_3756,N_2031,N_1480);
and U3757 (N_3757,N_2077,N_2851);
nand U3758 (N_3758,N_2435,N_1232);
or U3759 (N_3759,N_2011,N_77);
and U3760 (N_3760,N_708,N_7);
nor U3761 (N_3761,N_2502,N_1037);
nor U3762 (N_3762,N_1154,N_1442);
nand U3763 (N_3763,N_1000,N_2960);
nor U3764 (N_3764,N_2681,N_1191);
nor U3765 (N_3765,N_2549,N_2764);
and U3766 (N_3766,N_2949,N_2017);
and U3767 (N_3767,N_2619,N_1422);
nor U3768 (N_3768,N_2300,N_1947);
nor U3769 (N_3769,N_2296,N_1586);
nand U3770 (N_3770,N_961,N_2260);
or U3771 (N_3771,N_1796,N_1782);
or U3772 (N_3772,N_2477,N_1285);
or U3773 (N_3773,N_2671,N_1876);
nand U3774 (N_3774,N_71,N_310);
or U3775 (N_3775,N_1905,N_50);
and U3776 (N_3776,N_36,N_1842);
and U3777 (N_3777,N_2065,N_1175);
nand U3778 (N_3778,N_2732,N_1058);
or U3779 (N_3779,N_2979,N_2058);
nor U3780 (N_3780,N_1375,N_1518);
nor U3781 (N_3781,N_1811,N_1497);
and U3782 (N_3782,N_1322,N_2606);
nor U3783 (N_3783,N_2219,N_1992);
or U3784 (N_3784,N_682,N_1343);
and U3785 (N_3785,N_666,N_647);
or U3786 (N_3786,N_167,N_1951);
and U3787 (N_3787,N_1756,N_1204);
or U3788 (N_3788,N_1631,N_367);
nor U3789 (N_3789,N_2858,N_1831);
nand U3790 (N_3790,N_1732,N_1875);
nor U3791 (N_3791,N_901,N_2920);
or U3792 (N_3792,N_2051,N_2482);
nand U3793 (N_3793,N_2417,N_1094);
and U3794 (N_3794,N_2112,N_594);
nor U3795 (N_3795,N_1458,N_942);
nor U3796 (N_3796,N_2616,N_2652);
and U3797 (N_3797,N_2614,N_1998);
and U3798 (N_3798,N_1601,N_519);
nor U3799 (N_3799,N_2883,N_1257);
and U3800 (N_3800,N_2181,N_347);
nand U3801 (N_3801,N_1812,N_506);
and U3802 (N_3802,N_82,N_436);
nand U3803 (N_3803,N_865,N_2399);
or U3804 (N_3804,N_652,N_714);
or U3805 (N_3805,N_1413,N_208);
or U3806 (N_3806,N_1886,N_147);
nand U3807 (N_3807,N_2314,N_116);
and U3808 (N_3808,N_2794,N_1660);
or U3809 (N_3809,N_469,N_2401);
nor U3810 (N_3810,N_2220,N_124);
nand U3811 (N_3811,N_982,N_99);
nand U3812 (N_3812,N_222,N_1655);
nand U3813 (N_3813,N_2476,N_294);
and U3814 (N_3814,N_561,N_2023);
nand U3815 (N_3815,N_1628,N_290);
or U3816 (N_3816,N_1414,N_1389);
nor U3817 (N_3817,N_2999,N_630);
nand U3818 (N_3818,N_322,N_1427);
nor U3819 (N_3819,N_2864,N_1030);
nand U3820 (N_3820,N_595,N_1252);
nand U3821 (N_3821,N_1889,N_1563);
and U3822 (N_3822,N_218,N_620);
or U3823 (N_3823,N_2013,N_2620);
nand U3824 (N_3824,N_2322,N_2578);
or U3825 (N_3825,N_2571,N_2457);
nand U3826 (N_3826,N_2208,N_2103);
nor U3827 (N_3827,N_646,N_1410);
and U3828 (N_3828,N_2573,N_2025);
nor U3829 (N_3829,N_980,N_872);
nor U3830 (N_3830,N_1965,N_1318);
or U3831 (N_3831,N_1240,N_2776);
or U3832 (N_3832,N_1633,N_1482);
nor U3833 (N_3833,N_1860,N_1306);
and U3834 (N_3834,N_123,N_2090);
nand U3835 (N_3835,N_1659,N_1955);
nor U3836 (N_3836,N_809,N_1731);
and U3837 (N_3837,N_2595,N_192);
and U3838 (N_3838,N_1106,N_1846);
nor U3839 (N_3839,N_112,N_1095);
nor U3840 (N_3840,N_2488,N_2775);
or U3841 (N_3841,N_127,N_1950);
nor U3842 (N_3842,N_2938,N_1393);
or U3843 (N_3843,N_1594,N_1065);
and U3844 (N_3844,N_1057,N_2460);
nor U3845 (N_3845,N_779,N_857);
nor U3846 (N_3846,N_804,N_2788);
or U3847 (N_3847,N_1588,N_2019);
nor U3848 (N_3848,N_2812,N_1186);
or U3849 (N_3849,N_1125,N_2810);
and U3850 (N_3850,N_2222,N_1097);
and U3851 (N_3851,N_778,N_788);
nand U3852 (N_3852,N_55,N_333);
and U3853 (N_3853,N_1961,N_724);
nand U3854 (N_3854,N_2964,N_2336);
nor U3855 (N_3855,N_641,N_2721);
nand U3856 (N_3856,N_2662,N_1582);
or U3857 (N_3857,N_756,N_1930);
and U3858 (N_3858,N_1032,N_2928);
or U3859 (N_3859,N_1884,N_1370);
or U3860 (N_3860,N_2947,N_726);
or U3861 (N_3861,N_477,N_2567);
or U3862 (N_3862,N_482,N_1122);
nand U3863 (N_3863,N_2643,N_2524);
or U3864 (N_3864,N_425,N_875);
and U3865 (N_3865,N_1828,N_2429);
nand U3866 (N_3866,N_502,N_2574);
nor U3867 (N_3867,N_1678,N_2366);
or U3868 (N_3868,N_2503,N_1237);
and U3869 (N_3869,N_2331,N_2981);
nor U3870 (N_3870,N_2825,N_1075);
nor U3871 (N_3871,N_2699,N_2365);
nand U3872 (N_3872,N_2329,N_2334);
nor U3873 (N_3873,N_1246,N_2180);
and U3874 (N_3874,N_191,N_1932);
or U3875 (N_3875,N_1132,N_2345);
nand U3876 (N_3876,N_1661,N_2273);
nor U3877 (N_3877,N_1589,N_706);
and U3878 (N_3878,N_1077,N_2965);
or U3879 (N_3879,N_662,N_1561);
nor U3880 (N_3880,N_1792,N_366);
nand U3881 (N_3881,N_2134,N_1625);
nand U3882 (N_3882,N_2414,N_2214);
nand U3883 (N_3883,N_2094,N_2022);
or U3884 (N_3884,N_618,N_1093);
nand U3885 (N_3885,N_327,N_426);
nor U3886 (N_3886,N_264,N_1774);
and U3887 (N_3887,N_1347,N_1510);
or U3888 (N_3888,N_2925,N_1128);
nand U3889 (N_3889,N_1523,N_2100);
or U3890 (N_3890,N_2799,N_2832);
xor U3891 (N_3891,N_1707,N_2395);
nor U3892 (N_3892,N_729,N_2000);
or U3893 (N_3893,N_1918,N_78);
nand U3894 (N_3894,N_2413,N_2084);
nor U3895 (N_3895,N_2765,N_1072);
nor U3896 (N_3896,N_1536,N_496);
or U3897 (N_3897,N_1194,N_493);
nor U3898 (N_3898,N_543,N_220);
and U3899 (N_3899,N_2647,N_2249);
and U3900 (N_3900,N_1848,N_780);
nor U3901 (N_3901,N_480,N_2140);
nand U3902 (N_3902,N_1532,N_2394);
or U3903 (N_3903,N_1515,N_535);
nor U3904 (N_3904,N_1195,N_2861);
and U3905 (N_3905,N_2263,N_2709);
nor U3906 (N_3906,N_1400,N_516);
and U3907 (N_3907,N_2041,N_2093);
nand U3908 (N_3908,N_686,N_1271);
nand U3909 (N_3909,N_948,N_1632);
nand U3910 (N_3910,N_2280,N_2227);
nor U3911 (N_3911,N_2466,N_1021);
nor U3912 (N_3912,N_1301,N_792);
and U3913 (N_3913,N_1490,N_546);
and U3914 (N_3914,N_1492,N_789);
and U3915 (N_3915,N_2262,N_423);
xor U3916 (N_3916,N_1309,N_1018);
nor U3917 (N_3917,N_640,N_976);
or U3918 (N_3918,N_174,N_361);
nor U3919 (N_3919,N_295,N_1267);
nand U3920 (N_3920,N_2990,N_265);
and U3921 (N_3921,N_2276,N_2448);
nor U3922 (N_3922,N_2612,N_388);
and U3923 (N_3923,N_2668,N_2010);
and U3924 (N_3924,N_1228,N_273);
nand U3925 (N_3925,N_1861,N_743);
and U3926 (N_3926,N_20,N_2251);
nor U3927 (N_3927,N_2905,N_739);
or U3928 (N_3928,N_2129,N_1387);
nor U3929 (N_3929,N_2637,N_590);
and U3930 (N_3930,N_1801,N_1725);
nor U3931 (N_3931,N_673,N_262);
and U3932 (N_3932,N_2608,N_2073);
nand U3933 (N_3933,N_2922,N_2943);
nor U3934 (N_3934,N_403,N_18);
or U3935 (N_3935,N_2312,N_2560);
nand U3936 (N_3936,N_1225,N_1457);
nand U3937 (N_3937,N_2284,N_1866);
or U3938 (N_3938,N_283,N_2635);
nor U3939 (N_3939,N_737,N_2511);
or U3940 (N_3940,N_823,N_753);
and U3941 (N_3941,N_577,N_1296);
nor U3942 (N_3942,N_2225,N_2351);
or U3943 (N_3943,N_1803,N_1741);
and U3944 (N_3944,N_2257,N_643);
nor U3945 (N_3945,N_389,N_2348);
and U3946 (N_3946,N_2523,N_1666);
and U3947 (N_3947,N_943,N_858);
nand U3948 (N_3948,N_2749,N_2178);
nor U3949 (N_3949,N_681,N_1383);
and U3950 (N_3950,N_1762,N_2035);
or U3951 (N_3951,N_1606,N_79);
or U3952 (N_3952,N_259,N_136);
nor U3953 (N_3953,N_2850,N_1551);
nand U3954 (N_3954,N_113,N_225);
nand U3955 (N_3955,N_571,N_2121);
nor U3956 (N_3956,N_2485,N_2254);
nor U3957 (N_3957,N_2332,N_1643);
nand U3958 (N_3958,N_1478,N_1511);
nor U3959 (N_3959,N_1129,N_2822);
or U3960 (N_3960,N_2877,N_17);
or U3961 (N_3961,N_2064,N_696);
or U3962 (N_3962,N_2978,N_239);
or U3963 (N_3963,N_2467,N_2270);
or U3964 (N_3964,N_2878,N_2088);
and U3965 (N_3965,N_2626,N_1674);
or U3966 (N_3966,N_2337,N_930);
nor U3967 (N_3967,N_526,N_2816);
or U3968 (N_3968,N_2551,N_2447);
xnor U3969 (N_3969,N_1234,N_406);
or U3970 (N_3970,N_328,N_1502);
nand U3971 (N_3971,N_2684,N_2475);
nor U3972 (N_3972,N_1836,N_326);
and U3973 (N_3973,N_1447,N_672);
nand U3974 (N_3974,N_926,N_1696);
or U3975 (N_3975,N_342,N_650);
and U3976 (N_3976,N_385,N_1302);
and U3977 (N_3977,N_2516,N_2160);
nor U3978 (N_3978,N_281,N_1041);
or U3979 (N_3979,N_1887,N_2970);
and U3980 (N_3980,N_1429,N_297);
nand U3981 (N_3981,N_2408,N_721);
nor U3982 (N_3982,N_358,N_1293);
nor U3983 (N_3983,N_997,N_1881);
and U3984 (N_3984,N_1592,N_2504);
and U3985 (N_3985,N_1157,N_861);
or U3986 (N_3986,N_723,N_184);
nor U3987 (N_3987,N_1704,N_1080);
or U3988 (N_3988,N_579,N_2110);
nand U3989 (N_3989,N_1808,N_1888);
nor U3990 (N_3990,N_2519,N_2097);
nand U3991 (N_3991,N_473,N_1345);
nor U3992 (N_3992,N_1989,N_748);
and U3993 (N_3993,N_763,N_2796);
or U3994 (N_3994,N_1272,N_2480);
or U3995 (N_3995,N_1777,N_44);
and U3996 (N_3996,N_540,N_1845);
nand U3997 (N_3997,N_1996,N_1198);
or U3998 (N_3998,N_2137,N_689);
nor U3999 (N_3999,N_2183,N_2780);
xnor U4000 (N_4000,N_850,N_1460);
or U4001 (N_4001,N_2963,N_2927);
and U4002 (N_4002,N_1469,N_251);
nand U4003 (N_4003,N_2422,N_1538);
and U4004 (N_4004,N_1710,N_1083);
nor U4005 (N_4005,N_2462,N_1476);
nor U4006 (N_4006,N_67,N_1202);
and U4007 (N_4007,N_2295,N_2941);
nand U4008 (N_4008,N_1654,N_2007);
and U4009 (N_4009,N_1467,N_1193);
or U4010 (N_4010,N_305,N_1574);
or U4011 (N_4011,N_2638,N_2358);
or U4012 (N_4012,N_1892,N_2119);
and U4013 (N_4013,N_108,N_1218);
nand U4014 (N_4014,N_2169,N_365);
nor U4015 (N_4015,N_816,N_345);
nor U4016 (N_4016,N_2454,N_1423);
and U4017 (N_4017,N_1340,N_731);
and U4018 (N_4018,N_1486,N_2188);
nand U4019 (N_4019,N_1854,N_374);
nand U4020 (N_4020,N_2838,N_2146);
or U4021 (N_4021,N_913,N_1850);
and U4022 (N_4022,N_1693,N_906);
nor U4023 (N_4023,N_2111,N_2272);
nor U4024 (N_4024,N_968,N_165);
nand U4025 (N_4025,N_2040,N_833);
nor U4026 (N_4026,N_2085,N_254);
and U4027 (N_4027,N_2598,N_1242);
or U4028 (N_4028,N_2194,N_1539);
and U4029 (N_4029,N_1407,N_1384);
nand U4030 (N_4030,N_166,N_1172);
and U4031 (N_4031,N_490,N_466);
nor U4032 (N_4032,N_1833,N_476);
nand U4033 (N_4033,N_236,N_1373);
nand U4034 (N_4034,N_1148,N_2509);
nor U4035 (N_4035,N_966,N_716);
or U4036 (N_4036,N_360,N_1934);
or U4037 (N_4037,N_2968,N_1620);
or U4038 (N_4038,N_2416,N_798);
or U4039 (N_4039,N_1357,N_1957);
or U4040 (N_4040,N_2275,N_1903);
or U4041 (N_4041,N_885,N_2489);
nand U4042 (N_4042,N_2698,N_841);
and U4043 (N_4043,N_2127,N_2079);
or U4044 (N_4044,N_1308,N_1100);
and U4045 (N_4045,N_2840,N_2727);
and U4046 (N_4046,N_2377,N_1718);
nand U4047 (N_4047,N_41,N_143);
nand U4048 (N_4048,N_1254,N_2820);
and U4049 (N_4049,N_1003,N_1837);
nand U4050 (N_4050,N_1627,N_313);
or U4051 (N_4051,N_1630,N_629);
and U4052 (N_4052,N_2412,N_1208);
and U4053 (N_4053,N_1369,N_2824);
nor U4054 (N_4054,N_2147,N_504);
and U4055 (N_4055,N_1019,N_1890);
nand U4056 (N_4056,N_2623,N_10);
nor U4057 (N_4057,N_1073,N_2290);
nor U4058 (N_4058,N_1815,N_1622);
and U4059 (N_4059,N_2618,N_1013);
nor U4060 (N_4060,N_700,N_455);
nand U4061 (N_4061,N_1494,N_531);
or U4062 (N_4062,N_2258,N_972);
and U4063 (N_4063,N_1415,N_2742);
or U4064 (N_4064,N_1323,N_39);
or U4065 (N_4065,N_1295,N_2790);
and U4066 (N_4066,N_2817,N_33);
nand U4067 (N_4067,N_329,N_1464);
nor U4068 (N_4068,N_422,N_497);
nor U4069 (N_4069,N_1090,N_785);
and U4070 (N_4070,N_2884,N_235);
or U4071 (N_4071,N_512,N_2246);
nand U4072 (N_4072,N_298,N_2463);
nor U4073 (N_4073,N_1220,N_27);
and U4074 (N_4074,N_1916,N_1635);
nor U4075 (N_4075,N_1287,N_1395);
nand U4076 (N_4076,N_1991,N_699);
and U4077 (N_4077,N_1656,N_1472);
xnor U4078 (N_4078,N_1231,N_791);
nor U4079 (N_4079,N_727,N_2243);
xor U4080 (N_4080,N_2343,N_2795);
nand U4081 (N_4081,N_185,N_2150);
or U4082 (N_4082,N_1102,N_2934);
nor U4083 (N_4083,N_256,N_156);
nand U4084 (N_4084,N_1027,N_537);
nand U4085 (N_4085,N_2586,N_1069);
or U4086 (N_4086,N_2715,N_1575);
and U4087 (N_4087,N_381,N_1420);
or U4088 (N_4088,N_1183,N_1091);
and U4089 (N_4089,N_81,N_1982);
nand U4090 (N_4090,N_1553,N_1853);
nor U4091 (N_4091,N_171,N_1317);
nand U4092 (N_4092,N_2349,N_1519);
and U4093 (N_4093,N_805,N_2989);
nand U4094 (N_4094,N_475,N_1426);
nand U4095 (N_4095,N_26,N_1320);
nand U4096 (N_4096,N_125,N_271);
and U4097 (N_4097,N_1067,N_2545);
or U4098 (N_4098,N_2769,N_814);
and U4099 (N_4099,N_1541,N_978);
or U4100 (N_4100,N_2393,N_568);
and U4101 (N_4101,N_162,N_576);
nand U4102 (N_4102,N_131,N_695);
nor U4103 (N_4103,N_2109,N_1669);
nand U4104 (N_4104,N_160,N_1002);
nor U4105 (N_4105,N_625,N_2292);
nand U4106 (N_4106,N_1053,N_448);
and U4107 (N_4107,N_2983,N_2874);
nor U4108 (N_4108,N_565,N_1931);
and U4109 (N_4109,N_970,N_1074);
or U4110 (N_4110,N_1694,N_120);
nor U4111 (N_4111,N_1078,N_243);
nor U4112 (N_4112,N_1475,N_2364);
and U4113 (N_4113,N_2163,N_1800);
and U4114 (N_4114,N_703,N_386);
and U4115 (N_4115,N_1794,N_2486);
or U4116 (N_4116,N_58,N_418);
or U4117 (N_4117,N_2047,N_1763);
nor U4118 (N_4118,N_636,N_2584);
and U4119 (N_4119,N_887,N_1463);
nor U4120 (N_4120,N_2068,N_2665);
and U4121 (N_4121,N_2507,N_1354);
nor U4122 (N_4122,N_1164,N_2081);
nor U4123 (N_4123,N_745,N_2886);
or U4124 (N_4124,N_2846,N_752);
and U4125 (N_4125,N_122,N_1159);
nor U4126 (N_4126,N_312,N_878);
or U4127 (N_4127,N_11,N_76);
nor U4128 (N_4128,N_1750,N_104);
nor U4129 (N_4129,N_1608,N_1042);
nor U4130 (N_4130,N_899,N_2230);
and U4131 (N_4131,N_615,N_100);
nand U4132 (N_4132,N_277,N_1692);
nand U4133 (N_4133,N_2404,N_1116);
nand U4134 (N_4134,N_593,N_1976);
and U4135 (N_4135,N_1029,N_1136);
nand U4136 (N_4136,N_1891,N_2038);
nor U4137 (N_4137,N_1190,N_2696);
or U4138 (N_4138,N_119,N_2056);
or U4139 (N_4139,N_951,N_2621);
nor U4140 (N_4140,N_284,N_1537);
nand U4141 (N_4141,N_1233,N_291);
nand U4142 (N_4142,N_2240,N_492);
nor U4143 (N_4143,N_2791,N_2936);
nand U4144 (N_4144,N_363,N_985);
or U4145 (N_4145,N_1639,N_701);
nand U4146 (N_4146,N_2285,N_1542);
nand U4147 (N_4147,N_1437,N_1987);
or U4148 (N_4148,N_2032,N_2512);
and U4149 (N_4149,N_1005,N_268);
and U4150 (N_4150,N_1219,N_2670);
or U4151 (N_4151,N_1591,N_2133);
nor U4152 (N_4152,N_2210,N_1001);
and U4153 (N_4153,N_2646,N_994);
and U4154 (N_4154,N_1188,N_1205);
nand U4155 (N_4155,N_1681,N_204);
or U4156 (N_4156,N_2653,N_584);
or U4157 (N_4157,N_2174,N_2809);
or U4158 (N_4158,N_179,N_2291);
and U4159 (N_4159,N_359,N_2939);
nor U4160 (N_4160,N_1329,N_241);
or U4161 (N_4161,N_1869,N_260);
or U4162 (N_4162,N_2529,N_66);
and U4163 (N_4163,N_2255,N_2202);
nor U4164 (N_4164,N_2148,N_97);
nand U4165 (N_4165,N_908,N_507);
or U4166 (N_4166,N_1893,N_2746);
or U4167 (N_4167,N_2184,N_1008);
nand U4168 (N_4168,N_1779,N_515);
nand U4169 (N_4169,N_1170,N_894);
and U4170 (N_4170,N_784,N_2278);
nor U4171 (N_4171,N_599,N_626);
nand U4172 (N_4172,N_1401,N_94);
and U4173 (N_4173,N_1253,N_1820);
nand U4174 (N_4174,N_1923,N_2126);
nor U4175 (N_4175,N_105,N_1945);
nand U4176 (N_4176,N_1394,N_1372);
or U4177 (N_4177,N_1533,N_2501);
nor U4178 (N_4178,N_1706,N_1958);
or U4179 (N_4179,N_304,N_106);
and U4180 (N_4180,N_1724,N_1089);
nor U4181 (N_4181,N_2907,N_246);
nor U4182 (N_4182,N_607,N_802);
or U4183 (N_4183,N_2644,N_2427);
or U4184 (N_4184,N_1264,N_2459);
and U4185 (N_4185,N_1521,N_2786);
and U4186 (N_4186,N_2682,N_2654);
or U4187 (N_4187,N_193,N_180);
nor U4188 (N_4188,N_150,N_2935);
nand U4189 (N_4189,N_2615,N_37);
and U4190 (N_4190,N_2231,N_2443);
or U4191 (N_4191,N_90,N_1540);
and U4192 (N_4192,N_562,N_1086);
or U4193 (N_4193,N_2526,N_2039);
and U4194 (N_4194,N_671,N_1504);
nand U4195 (N_4195,N_613,N_2315);
or U4196 (N_4196,N_395,N_464);
or U4197 (N_4197,N_471,N_831);
or U4198 (N_4198,N_63,N_1303);
or U4199 (N_4199,N_182,N_2195);
or U4200 (N_4200,N_1844,N_1404);
and U4201 (N_4201,N_292,N_1134);
or U4202 (N_4202,N_1721,N_1446);
nor U4203 (N_4203,N_918,N_1066);
or U4204 (N_4204,N_619,N_1133);
or U4205 (N_4205,N_676,N_1997);
and U4206 (N_4206,N_2494,N_979);
or U4207 (N_4207,N_102,N_2327);
or U4208 (N_4208,N_2591,N_1908);
or U4209 (N_4209,N_2648,N_1920);
nand U4210 (N_4210,N_2080,N_2711);
nor U4211 (N_4211,N_898,N_2245);
nand U4212 (N_4212,N_755,N_1783);
nor U4213 (N_4213,N_1359,N_2207);
or U4214 (N_4214,N_880,N_556);
and U4215 (N_4215,N_1550,N_2396);
nand U4216 (N_4216,N_659,N_1238);
and U4217 (N_4217,N_1830,N_1983);
and U4218 (N_4218,N_1217,N_1289);
nor U4219 (N_4219,N_530,N_2543);
nand U4220 (N_4220,N_1435,N_1283);
or U4221 (N_4221,N_382,N_211);
nand U4222 (N_4222,N_1740,N_2556);
and U4223 (N_4223,N_1759,N_2828);
nand U4224 (N_4224,N_1587,N_803);
or U4225 (N_4225,N_2515,N_459);
and U4226 (N_4226,N_462,N_720);
nor U4227 (N_4227,N_2014,N_2374);
or U4228 (N_4228,N_1547,N_1703);
or U4229 (N_4229,N_2857,N_2123);
nor U4230 (N_4230,N_1173,N_2124);
nor U4231 (N_4231,N_2076,N_1573);
or U4232 (N_4232,N_2921,N_1227);
or U4233 (N_4233,N_859,N_2664);
nand U4234 (N_4234,N_2694,N_527);
nor U4235 (N_4235,N_2006,N_1355);
nor U4236 (N_4236,N_1730,N_838);
and U4237 (N_4237,N_2346,N_760);
nor U4238 (N_4238,N_2135,N_2012);
nand U4239 (N_4239,N_1381,N_384);
nor U4240 (N_4240,N_2033,N_190);
or U4241 (N_4241,N_1433,N_840);
nand U4242 (N_4242,N_1936,N_2238);
nor U4243 (N_4243,N_2761,N_1418);
or U4244 (N_4244,N_2338,N_2281);
or U4245 (N_4245,N_2625,N_353);
nor U4246 (N_4246,N_685,N_2793);
nor U4247 (N_4247,N_1590,N_2239);
and U4248 (N_4248,N_822,N_398);
and U4249 (N_4249,N_1980,N_457);
or U4250 (N_4250,N_1749,N_437);
or U4251 (N_4251,N_1863,N_2714);
and U4252 (N_4252,N_1851,N_331);
nand U4253 (N_4253,N_627,N_355);
nor U4254 (N_4254,N_1771,N_1953);
and U4255 (N_4255,N_2641,N_1769);
nand U4256 (N_4256,N_478,N_879);
and U4257 (N_4257,N_2362,N_111);
nor U4258 (N_4258,N_369,N_1535);
or U4259 (N_4259,N_1040,N_228);
nand U4260 (N_4260,N_628,N_2957);
nand U4261 (N_4261,N_1352,N_2269);
and U4262 (N_4262,N_1570,N_544);
and U4263 (N_4263,N_554,N_817);
nand U4264 (N_4264,N_2569,N_1753);
or U4265 (N_4265,N_1672,N_309);
nand U4266 (N_4266,N_2899,N_34);
and U4267 (N_4267,N_2356,N_675);
nand U4268 (N_4268,N_2530,N_2390);
and U4269 (N_4269,N_412,N_2157);
and U4270 (N_4270,N_1025,N_2313);
and U4271 (N_4271,N_159,N_825);
and U4272 (N_4272,N_1770,N_550);
and U4273 (N_4273,N_2105,N_2950);
or U4274 (N_4274,N_2456,N_1049);
and U4275 (N_4275,N_453,N_888);
nor U4276 (N_4276,N_2008,N_2988);
and U4277 (N_4277,N_2061,N_1744);
nand U4278 (N_4278,N_944,N_1599);
and U4279 (N_4279,N_370,N_524);
nand U4280 (N_4280,N_1459,N_1554);
and U4281 (N_4281,N_509,N_413);
or U4282 (N_4282,N_2583,N_2026);
and U4283 (N_4283,N_1938,N_279);
and U4284 (N_4284,N_338,N_1727);
or U4285 (N_4285,N_247,N_135);
nor U4286 (N_4286,N_393,N_9);
nand U4287 (N_4287,N_1637,N_1430);
nand U4288 (N_4288,N_2933,N_1787);
nor U4289 (N_4289,N_2130,N_1748);
nor U4290 (N_4290,N_754,N_346);
and U4291 (N_4291,N_990,N_1767);
and U4292 (N_4292,N_1728,N_2036);
nand U4293 (N_4293,N_59,N_2481);
and U4294 (N_4294,N_2587,N_710);
nand U4295 (N_4295,N_2403,N_1311);
and U4296 (N_4296,N_434,N_203);
and U4297 (N_4297,N_1284,N_2673);
nand U4298 (N_4298,N_2945,N_1278);
nand U4299 (N_4299,N_2388,N_1268);
nand U4300 (N_4300,N_2666,N_1166);
nor U4301 (N_4301,N_1922,N_871);
nand U4302 (N_4302,N_1585,N_1567);
or U4303 (N_4303,N_376,N_199);
and U4304 (N_4304,N_2386,N_2645);
and U4305 (N_4305,N_830,N_2096);
nand U4306 (N_4306,N_2695,N_952);
nor U4307 (N_4307,N_2984,N_1330);
nor U4308 (N_4308,N_1827,N_2283);
nand U4309 (N_4309,N_2544,N_735);
nor U4310 (N_4310,N_1988,N_1168);
and U4311 (N_4311,N_2835,N_1629);
or U4312 (N_4312,N_2688,N_337);
nand U4313 (N_4313,N_2473,N_138);
and U4314 (N_4314,N_1201,N_965);
and U4315 (N_4315,N_782,N_2658);
and U4316 (N_4316,N_1105,N_2189);
or U4317 (N_4317,N_514,N_932);
nor U4318 (N_4318,N_1805,N_1038);
and U4319 (N_4319,N_2426,N_799);
nand U4320 (N_4320,N_2683,N_1071);
or U4321 (N_4321,N_1224,N_2853);
or U4322 (N_4322,N_1315,N_2233);
nor U4323 (N_4323,N_911,N_306);
nand U4324 (N_4324,N_1680,N_2165);
nand U4325 (N_4325,N_362,N_1211);
and U4326 (N_4326,N_52,N_2142);
nand U4327 (N_4327,N_1841,N_2771);
or U4328 (N_4328,N_2149,N_2321);
and U4329 (N_4329,N_2942,N_1556);
or U4330 (N_4330,N_89,N_61);
and U4331 (N_4331,N_538,N_1568);
nand U4332 (N_4332,N_1130,N_364);
nand U4333 (N_4333,N_2533,N_1566);
or U4334 (N_4334,N_936,N_2154);
nor U4335 (N_4335,N_622,N_1943);
and U4336 (N_4336,N_1376,N_1241);
and U4337 (N_4337,N_1440,N_2906);
nor U4338 (N_4338,N_910,N_1761);
nor U4339 (N_4339,N_631,N_581);
and U4340 (N_4340,N_758,N_2901);
xor U4341 (N_4341,N_1153,N_257);
xor U4342 (N_4342,N_1155,N_1305);
nand U4343 (N_4343,N_420,N_1699);
and U4344 (N_4344,N_945,N_1764);
or U4345 (N_4345,N_2391,N_2392);
and U4346 (N_4346,N_1063,N_1896);
and U4347 (N_4347,N_547,N_2196);
or U4348 (N_4348,N_521,N_280);
xor U4349 (N_4349,N_1847,N_2268);
or U4350 (N_4350,N_1505,N_2030);
and U4351 (N_4351,N_196,N_1906);
nor U4352 (N_4352,N_2072,N_1882);
or U4353 (N_4353,N_1325,N_2106);
xor U4354 (N_4354,N_2660,N_2493);
or U4355 (N_4355,N_1940,N_287);
nor U4356 (N_4356,N_2247,N_2783);
or U4357 (N_4357,N_762,N_2602);
nand U4358 (N_4358,N_2879,N_2678);
nand U4359 (N_4359,N_1719,N_1668);
or U4360 (N_4360,N_2700,N_1697);
nor U4361 (N_4361,N_2932,N_563);
and U4362 (N_4362,N_2679,N_1156);
or U4363 (N_4363,N_940,N_924);
or U4364 (N_4364,N_2418,N_912);
and U4365 (N_4365,N_1967,N_2027);
or U4366 (N_4366,N_2419,N_57);
nor U4367 (N_4367,N_450,N_2773);
nor U4368 (N_4368,N_909,N_380);
nor U4369 (N_4369,N_2605,N_1335);
and U4370 (N_4370,N_2234,N_2363);
xor U4371 (N_4371,N_1176,N_1245);
or U4372 (N_4372,N_2674,N_439);
nor U4373 (N_4373,N_2136,N_2464);
or U4374 (N_4374,N_2224,N_1641);
or U4375 (N_4375,N_1275,N_1529);
or U4376 (N_4376,N_1313,N_1795);
nor U4377 (N_4377,N_1088,N_1399);
nor U4378 (N_4378,N_2301,N_2236);
nor U4379 (N_4379,N_2376,N_2171);
nand U4380 (N_4380,N_2353,N_1022);
or U4381 (N_4381,N_1675,N_1104);
and U4382 (N_4382,N_1274,N_2226);
or U4383 (N_4383,N_2152,N_1691);
or U4384 (N_4384,N_1793,N_141);
nand U4385 (N_4385,N_2069,N_1307);
nand U4386 (N_4386,N_608,N_2372);
or U4387 (N_4387,N_2842,N_505);
or U4388 (N_4388,N_1649,N_153);
nand U4389 (N_4389,N_250,N_2122);
nand U4390 (N_4390,N_349,N_2086);
or U4391 (N_4391,N_2540,N_2232);
xnor U4392 (N_4392,N_2054,N_684);
and U4393 (N_4393,N_651,N_2001);
or U4394 (N_4394,N_1912,N_2217);
nand U4395 (N_4395,N_2330,N_624);
nand U4396 (N_4396,N_764,N_92);
or U4397 (N_4397,N_1113,N_616);
and U4398 (N_4398,N_1682,N_1060);
and U4399 (N_4399,N_1348,N_2834);
or U4400 (N_4400,N_2099,N_1273);
or U4401 (N_4401,N_2955,N_1409);
nor U4402 (N_4402,N_2474,N_900);
or U4403 (N_4403,N_2629,N_1235);
nand U4404 (N_4404,N_1473,N_528);
nand U4405 (N_4405,N_1349,N_959);
nor U4406 (N_4406,N_2021,N_1722);
and U4407 (N_4407,N_410,N_109);
nor U4408 (N_4408,N_1454,N_1247);
and U4409 (N_4409,N_1766,N_32);
and U4410 (N_4410,N_495,N_25);
and U4411 (N_4411,N_1545,N_1495);
nor U4412 (N_4412,N_896,N_2357);
and U4413 (N_4413,N_205,N_2898);
nor U4414 (N_4414,N_2407,N_2420);
nor U4415 (N_4415,N_103,N_1747);
nor U4416 (N_4416,N_2057,N_928);
nor U4417 (N_4417,N_893,N_1012);
nand U4418 (N_4418,N_411,N_1412);
nor U4419 (N_4419,N_765,N_383);
nor U4420 (N_4420,N_1743,N_175);
and U4421 (N_4421,N_2271,N_542);
nand U4422 (N_4422,N_683,N_963);
or U4423 (N_4423,N_1901,N_2108);
and U4424 (N_4424,N_1045,N_836);
and U4425 (N_4425,N_1479,N_2075);
or U4426 (N_4426,N_1111,N_2114);
nand U4427 (N_4427,N_1645,N_1595);
and U4428 (N_4428,N_2914,N_2712);
and U4429 (N_4429,N_429,N_744);
xor U4430 (N_4430,N_194,N_51);
and U4431 (N_4431,N_1051,N_2500);
or U4432 (N_4432,N_1898,N_1184);
or U4433 (N_4433,N_1765,N_992);
and U4434 (N_4434,N_1977,N_2423);
nand U4435 (N_4435,N_796,N_2483);
nor U4436 (N_4436,N_1360,N_603);
nor U4437 (N_4437,N_1700,N_2951);
nand U4438 (N_4438,N_2718,N_1169);
nor U4439 (N_4439,N_269,N_1816);
and U4440 (N_4440,N_914,N_638);
nor U4441 (N_4441,N_905,N_1578);
nand U4442 (N_4442,N_330,N_2946);
nor U4443 (N_4443,N_2639,N_110);
or U4444 (N_4444,N_2186,N_1405);
xor U4445 (N_4445,N_927,N_115);
or U4446 (N_4446,N_2498,N_2213);
nor U4447 (N_4447,N_233,N_1304);
nand U4448 (N_4448,N_750,N_1688);
nor U4449 (N_4449,N_769,N_717);
or U4450 (N_4450,N_2373,N_2434);
nand U4451 (N_4451,N_118,N_503);
and U4452 (N_4452,N_2564,N_1135);
and U4453 (N_4453,N_2902,N_2091);
nor U4454 (N_4454,N_2995,N_998);
nor U4455 (N_4455,N_694,N_1919);
nand U4456 (N_4456,N_1124,N_2546);
nand U4457 (N_4457,N_1618,N_2289);
nor U4458 (N_4458,N_2020,N_2053);
nand U4459 (N_4459,N_2831,N_1339);
and U4460 (N_4460,N_2710,N_1462);
and U4461 (N_4461,N_583,N_1516);
and U4462 (N_4462,N_2568,N_1046);
and U4463 (N_4463,N_2361,N_1216);
and U4464 (N_4464,N_2768,N_1840);
nor U4465 (N_4465,N_922,N_2259);
or U4466 (N_4466,N_1825,N_2976);
nand U4467 (N_4467,N_820,N_1450);
xor U4468 (N_4468,N_40,N_2397);
and U4469 (N_4469,N_2580,N_996);
and U4470 (N_4470,N_775,N_1879);
or U4471 (N_4471,N_467,N_2763);
and U4472 (N_4472,N_869,N_1909);
nor U4473 (N_4473,N_1927,N_146);
nand U4474 (N_4474,N_408,N_1465);
nand U4475 (N_4475,N_1913,N_704);
and U4476 (N_4476,N_1178,N_2576);
nand U4477 (N_4477,N_868,N_1230);
nand U4478 (N_4478,N_1419,N_610);
nor U4479 (N_4479,N_209,N_1823);
nor U4480 (N_4480,N_746,N_1353);
or U4481 (N_4481,N_962,N_2704);
nand U4482 (N_4482,N_632,N_1255);
or U4483 (N_4483,N_2542,N_152);
nand U4484 (N_4484,N_1687,N_2201);
and U4485 (N_4485,N_989,N_1939);
or U4486 (N_4486,N_1441,N_2198);
nor U4487 (N_4487,N_1868,N_1362);
and U4488 (N_4488,N_2215,N_245);
nand U4489 (N_4489,N_1378,N_2410);
and U4490 (N_4490,N_2609,N_669);
nor U4491 (N_4491,N_592,N_1806);
or U4492 (N_4492,N_1525,N_2177);
nand U4493 (N_4493,N_2663,N_340);
and U4494 (N_4494,N_1079,N_308);
nand U4495 (N_4495,N_2458,N_1115);
and U4496 (N_4496,N_2890,N_2805);
and U4497 (N_4497,N_2009,N_1199);
or U4498 (N_4498,N_877,N_1593);
or U4499 (N_4499,N_1603,N_1781);
or U4500 (N_4500,N_1549,N_243);
nand U4501 (N_4501,N_1437,N_247);
or U4502 (N_4502,N_604,N_1795);
nand U4503 (N_4503,N_2046,N_27);
and U4504 (N_4504,N_1948,N_1074);
nor U4505 (N_4505,N_2689,N_1367);
nor U4506 (N_4506,N_33,N_793);
nor U4507 (N_4507,N_2661,N_769);
nor U4508 (N_4508,N_2723,N_314);
and U4509 (N_4509,N_2645,N_1963);
nor U4510 (N_4510,N_2377,N_1806);
nor U4511 (N_4511,N_116,N_31);
nor U4512 (N_4512,N_1802,N_1890);
nand U4513 (N_4513,N_1364,N_232);
and U4514 (N_4514,N_2280,N_1739);
or U4515 (N_4515,N_1027,N_181);
nor U4516 (N_4516,N_1956,N_655);
xor U4517 (N_4517,N_1410,N_654);
and U4518 (N_4518,N_1578,N_54);
nand U4519 (N_4519,N_1316,N_32);
or U4520 (N_4520,N_783,N_1077);
xnor U4521 (N_4521,N_2093,N_2358);
or U4522 (N_4522,N_1824,N_2332);
or U4523 (N_4523,N_2164,N_2847);
or U4524 (N_4524,N_1331,N_2323);
nand U4525 (N_4525,N_2078,N_480);
nand U4526 (N_4526,N_347,N_1662);
or U4527 (N_4527,N_1414,N_1391);
and U4528 (N_4528,N_1848,N_2149);
nand U4529 (N_4529,N_374,N_2356);
nor U4530 (N_4530,N_2218,N_62);
or U4531 (N_4531,N_2139,N_1047);
nand U4532 (N_4532,N_2816,N_1326);
nor U4533 (N_4533,N_602,N_2308);
or U4534 (N_4534,N_1365,N_778);
nand U4535 (N_4535,N_2129,N_2745);
or U4536 (N_4536,N_2566,N_678);
nor U4537 (N_4537,N_197,N_2659);
and U4538 (N_4538,N_2474,N_1584);
nand U4539 (N_4539,N_152,N_2531);
nand U4540 (N_4540,N_2763,N_543);
nor U4541 (N_4541,N_2964,N_633);
and U4542 (N_4542,N_167,N_1883);
nor U4543 (N_4543,N_46,N_1006);
or U4544 (N_4544,N_2904,N_931);
nand U4545 (N_4545,N_210,N_1103);
nor U4546 (N_4546,N_1879,N_894);
and U4547 (N_4547,N_748,N_832);
or U4548 (N_4548,N_2365,N_575);
nand U4549 (N_4549,N_666,N_208);
nand U4550 (N_4550,N_650,N_500);
nand U4551 (N_4551,N_1441,N_584);
nand U4552 (N_4552,N_610,N_1663);
nand U4553 (N_4553,N_1042,N_956);
or U4554 (N_4554,N_1844,N_91);
and U4555 (N_4555,N_1987,N_2517);
and U4556 (N_4556,N_445,N_2354);
and U4557 (N_4557,N_2487,N_2462);
nor U4558 (N_4558,N_157,N_397);
nand U4559 (N_4559,N_983,N_817);
xnor U4560 (N_4560,N_42,N_2025);
and U4561 (N_4561,N_310,N_1049);
nand U4562 (N_4562,N_1820,N_2472);
nand U4563 (N_4563,N_963,N_1623);
nand U4564 (N_4564,N_2806,N_2229);
or U4565 (N_4565,N_76,N_1972);
or U4566 (N_4566,N_1013,N_811);
nand U4567 (N_4567,N_1683,N_512);
nand U4568 (N_4568,N_989,N_2480);
nand U4569 (N_4569,N_681,N_1635);
nand U4570 (N_4570,N_586,N_863);
or U4571 (N_4571,N_1256,N_2889);
nor U4572 (N_4572,N_1715,N_852);
and U4573 (N_4573,N_1579,N_1212);
nand U4574 (N_4574,N_400,N_47);
and U4575 (N_4575,N_789,N_216);
or U4576 (N_4576,N_478,N_737);
and U4577 (N_4577,N_2938,N_1761);
and U4578 (N_4578,N_807,N_84);
and U4579 (N_4579,N_382,N_219);
nor U4580 (N_4580,N_1719,N_1318);
nor U4581 (N_4581,N_2514,N_2137);
xnor U4582 (N_4582,N_2338,N_1113);
nand U4583 (N_4583,N_1657,N_792);
and U4584 (N_4584,N_2056,N_334);
and U4585 (N_4585,N_2164,N_2994);
nand U4586 (N_4586,N_1746,N_459);
nand U4587 (N_4587,N_608,N_199);
and U4588 (N_4588,N_931,N_1656);
nor U4589 (N_4589,N_2846,N_87);
nor U4590 (N_4590,N_2874,N_321);
nor U4591 (N_4591,N_1968,N_2535);
nor U4592 (N_4592,N_1341,N_1355);
nor U4593 (N_4593,N_2640,N_2090);
and U4594 (N_4594,N_2184,N_1823);
or U4595 (N_4595,N_284,N_1275);
or U4596 (N_4596,N_219,N_82);
and U4597 (N_4597,N_141,N_1228);
nor U4598 (N_4598,N_1398,N_392);
or U4599 (N_4599,N_612,N_1435);
nand U4600 (N_4600,N_2549,N_417);
nand U4601 (N_4601,N_1793,N_908);
nor U4602 (N_4602,N_1837,N_1143);
or U4603 (N_4603,N_1761,N_1972);
nand U4604 (N_4604,N_2062,N_2335);
and U4605 (N_4605,N_1632,N_80);
nand U4606 (N_4606,N_2059,N_891);
and U4607 (N_4607,N_2386,N_659);
or U4608 (N_4608,N_1312,N_1658);
or U4609 (N_4609,N_1867,N_2919);
or U4610 (N_4610,N_1924,N_570);
nand U4611 (N_4611,N_2552,N_842);
and U4612 (N_4612,N_1645,N_309);
and U4613 (N_4613,N_699,N_2504);
nor U4614 (N_4614,N_2069,N_1806);
and U4615 (N_4615,N_1892,N_1692);
nor U4616 (N_4616,N_2805,N_2806);
nor U4617 (N_4617,N_2517,N_2468);
or U4618 (N_4618,N_559,N_2987);
and U4619 (N_4619,N_607,N_2700);
nor U4620 (N_4620,N_2417,N_2302);
nand U4621 (N_4621,N_2783,N_2316);
and U4622 (N_4622,N_192,N_64);
and U4623 (N_4623,N_2749,N_2189);
or U4624 (N_4624,N_2743,N_1297);
and U4625 (N_4625,N_707,N_2317);
or U4626 (N_4626,N_2972,N_2520);
nand U4627 (N_4627,N_443,N_2813);
nor U4628 (N_4628,N_296,N_56);
nor U4629 (N_4629,N_1333,N_31);
or U4630 (N_4630,N_1357,N_2512);
nand U4631 (N_4631,N_543,N_2658);
or U4632 (N_4632,N_167,N_1171);
and U4633 (N_4633,N_599,N_2557);
and U4634 (N_4634,N_638,N_1582);
nor U4635 (N_4635,N_1717,N_1727);
and U4636 (N_4636,N_1337,N_1057);
nand U4637 (N_4637,N_1279,N_902);
or U4638 (N_4638,N_2369,N_1583);
and U4639 (N_4639,N_1973,N_2025);
nand U4640 (N_4640,N_996,N_2927);
and U4641 (N_4641,N_2780,N_1980);
nand U4642 (N_4642,N_500,N_1592);
nor U4643 (N_4643,N_2490,N_2981);
and U4644 (N_4644,N_2026,N_1040);
nand U4645 (N_4645,N_2191,N_2781);
and U4646 (N_4646,N_2492,N_1081);
and U4647 (N_4647,N_33,N_1827);
and U4648 (N_4648,N_1396,N_220);
or U4649 (N_4649,N_2554,N_1409);
nor U4650 (N_4650,N_2219,N_1001);
and U4651 (N_4651,N_1920,N_1159);
and U4652 (N_4652,N_515,N_1688);
nor U4653 (N_4653,N_813,N_1365);
or U4654 (N_4654,N_2396,N_2683);
or U4655 (N_4655,N_2947,N_1936);
or U4656 (N_4656,N_314,N_63);
nand U4657 (N_4657,N_2328,N_61);
and U4658 (N_4658,N_434,N_1371);
nor U4659 (N_4659,N_690,N_371);
nor U4660 (N_4660,N_74,N_2755);
nor U4661 (N_4661,N_1581,N_1360);
or U4662 (N_4662,N_369,N_681);
or U4663 (N_4663,N_2192,N_104);
or U4664 (N_4664,N_508,N_1855);
nor U4665 (N_4665,N_131,N_1719);
nor U4666 (N_4666,N_2960,N_1700);
nand U4667 (N_4667,N_823,N_1952);
or U4668 (N_4668,N_2323,N_2445);
nand U4669 (N_4669,N_701,N_1340);
nor U4670 (N_4670,N_2455,N_543);
nand U4671 (N_4671,N_2817,N_636);
nor U4672 (N_4672,N_1027,N_2661);
nor U4673 (N_4673,N_1087,N_1605);
and U4674 (N_4674,N_574,N_1709);
or U4675 (N_4675,N_2886,N_1285);
nand U4676 (N_4676,N_1049,N_1807);
and U4677 (N_4677,N_2862,N_1821);
nand U4678 (N_4678,N_1804,N_1952);
or U4679 (N_4679,N_2991,N_1392);
or U4680 (N_4680,N_1516,N_2626);
nand U4681 (N_4681,N_2628,N_2973);
or U4682 (N_4682,N_140,N_2566);
nor U4683 (N_4683,N_943,N_960);
nand U4684 (N_4684,N_2583,N_2746);
nand U4685 (N_4685,N_2245,N_2757);
and U4686 (N_4686,N_2745,N_430);
and U4687 (N_4687,N_1620,N_2567);
nand U4688 (N_4688,N_1809,N_1078);
and U4689 (N_4689,N_3,N_334);
nor U4690 (N_4690,N_49,N_1666);
or U4691 (N_4691,N_1039,N_1816);
and U4692 (N_4692,N_2741,N_2644);
or U4693 (N_4693,N_2794,N_573);
or U4694 (N_4694,N_2604,N_2333);
or U4695 (N_4695,N_1196,N_2335);
and U4696 (N_4696,N_738,N_2532);
nand U4697 (N_4697,N_1733,N_2353);
or U4698 (N_4698,N_1256,N_2112);
nor U4699 (N_4699,N_207,N_1548);
or U4700 (N_4700,N_2371,N_1581);
and U4701 (N_4701,N_825,N_1470);
or U4702 (N_4702,N_1238,N_2337);
and U4703 (N_4703,N_766,N_1858);
or U4704 (N_4704,N_1099,N_1472);
and U4705 (N_4705,N_1980,N_2702);
or U4706 (N_4706,N_1833,N_1416);
or U4707 (N_4707,N_718,N_1225);
nand U4708 (N_4708,N_1009,N_1422);
and U4709 (N_4709,N_1868,N_683);
or U4710 (N_4710,N_1212,N_924);
and U4711 (N_4711,N_349,N_2349);
or U4712 (N_4712,N_1612,N_51);
nor U4713 (N_4713,N_1229,N_276);
and U4714 (N_4714,N_570,N_1318);
and U4715 (N_4715,N_2708,N_2389);
and U4716 (N_4716,N_2616,N_373);
or U4717 (N_4717,N_2951,N_2174);
and U4718 (N_4718,N_626,N_1825);
nand U4719 (N_4719,N_978,N_1552);
xor U4720 (N_4720,N_460,N_2686);
or U4721 (N_4721,N_443,N_2980);
and U4722 (N_4722,N_96,N_500);
nor U4723 (N_4723,N_723,N_865);
or U4724 (N_4724,N_2085,N_2518);
and U4725 (N_4725,N_612,N_7);
and U4726 (N_4726,N_1698,N_41);
or U4727 (N_4727,N_2490,N_744);
nor U4728 (N_4728,N_2618,N_2072);
or U4729 (N_4729,N_1243,N_493);
nand U4730 (N_4730,N_618,N_1183);
and U4731 (N_4731,N_1736,N_2099);
and U4732 (N_4732,N_1416,N_1508);
nor U4733 (N_4733,N_2191,N_617);
nand U4734 (N_4734,N_1447,N_183);
and U4735 (N_4735,N_1026,N_1415);
and U4736 (N_4736,N_2857,N_2348);
and U4737 (N_4737,N_654,N_1857);
or U4738 (N_4738,N_2301,N_2414);
nor U4739 (N_4739,N_1795,N_214);
or U4740 (N_4740,N_317,N_1917);
or U4741 (N_4741,N_1062,N_275);
and U4742 (N_4742,N_2506,N_2896);
and U4743 (N_4743,N_2823,N_1771);
nand U4744 (N_4744,N_210,N_1035);
nor U4745 (N_4745,N_2802,N_1812);
and U4746 (N_4746,N_1886,N_1281);
nand U4747 (N_4747,N_1398,N_2455);
nand U4748 (N_4748,N_1963,N_178);
or U4749 (N_4749,N_2987,N_832);
nand U4750 (N_4750,N_2609,N_472);
nand U4751 (N_4751,N_2907,N_1801);
or U4752 (N_4752,N_1873,N_364);
and U4753 (N_4753,N_899,N_1461);
nand U4754 (N_4754,N_1920,N_2615);
nand U4755 (N_4755,N_109,N_1713);
and U4756 (N_4756,N_1660,N_2574);
nand U4757 (N_4757,N_2369,N_350);
and U4758 (N_4758,N_825,N_2717);
and U4759 (N_4759,N_2671,N_2053);
or U4760 (N_4760,N_225,N_2221);
or U4761 (N_4761,N_466,N_2609);
xor U4762 (N_4762,N_804,N_1356);
nor U4763 (N_4763,N_483,N_646);
or U4764 (N_4764,N_1441,N_1219);
and U4765 (N_4765,N_378,N_1073);
nand U4766 (N_4766,N_2630,N_97);
or U4767 (N_4767,N_2966,N_1302);
nand U4768 (N_4768,N_2900,N_2332);
nand U4769 (N_4769,N_787,N_190);
and U4770 (N_4770,N_300,N_1701);
nor U4771 (N_4771,N_2494,N_1494);
nand U4772 (N_4772,N_2939,N_1293);
nand U4773 (N_4773,N_2084,N_230);
nand U4774 (N_4774,N_1061,N_2576);
nand U4775 (N_4775,N_690,N_2370);
and U4776 (N_4776,N_1817,N_924);
and U4777 (N_4777,N_939,N_2881);
and U4778 (N_4778,N_805,N_1345);
or U4779 (N_4779,N_2743,N_1857);
nand U4780 (N_4780,N_2633,N_134);
nand U4781 (N_4781,N_1685,N_1065);
nand U4782 (N_4782,N_2075,N_1785);
and U4783 (N_4783,N_802,N_281);
nand U4784 (N_4784,N_1864,N_2430);
or U4785 (N_4785,N_1798,N_700);
xor U4786 (N_4786,N_2321,N_119);
and U4787 (N_4787,N_708,N_2998);
or U4788 (N_4788,N_1974,N_142);
nand U4789 (N_4789,N_426,N_1879);
nand U4790 (N_4790,N_62,N_227);
nor U4791 (N_4791,N_2985,N_1008);
nand U4792 (N_4792,N_2573,N_916);
nand U4793 (N_4793,N_1766,N_2819);
xor U4794 (N_4794,N_2389,N_1773);
nor U4795 (N_4795,N_1993,N_855);
nand U4796 (N_4796,N_251,N_2270);
and U4797 (N_4797,N_2862,N_2914);
nor U4798 (N_4798,N_2150,N_2877);
nor U4799 (N_4799,N_1629,N_396);
nor U4800 (N_4800,N_1419,N_1392);
nand U4801 (N_4801,N_1183,N_1591);
and U4802 (N_4802,N_2056,N_824);
nor U4803 (N_4803,N_2738,N_1706);
nor U4804 (N_4804,N_966,N_2333);
nor U4805 (N_4805,N_193,N_2347);
and U4806 (N_4806,N_2326,N_324);
nand U4807 (N_4807,N_1591,N_2029);
and U4808 (N_4808,N_561,N_2767);
or U4809 (N_4809,N_2012,N_2397);
nor U4810 (N_4810,N_2554,N_1841);
nor U4811 (N_4811,N_1516,N_1798);
or U4812 (N_4812,N_1083,N_336);
and U4813 (N_4813,N_2814,N_1362);
nand U4814 (N_4814,N_296,N_2789);
nor U4815 (N_4815,N_286,N_2244);
nand U4816 (N_4816,N_1188,N_787);
and U4817 (N_4817,N_1267,N_1160);
or U4818 (N_4818,N_1620,N_250);
nand U4819 (N_4819,N_2892,N_430);
and U4820 (N_4820,N_2988,N_2031);
or U4821 (N_4821,N_630,N_1656);
and U4822 (N_4822,N_2928,N_573);
nor U4823 (N_4823,N_991,N_186);
nor U4824 (N_4824,N_1402,N_2451);
or U4825 (N_4825,N_2702,N_1606);
and U4826 (N_4826,N_1745,N_1039);
or U4827 (N_4827,N_133,N_749);
or U4828 (N_4828,N_2559,N_2132);
or U4829 (N_4829,N_1682,N_2162);
nor U4830 (N_4830,N_407,N_1256);
nor U4831 (N_4831,N_1888,N_1697);
nor U4832 (N_4832,N_161,N_490);
or U4833 (N_4833,N_2985,N_1678);
and U4834 (N_4834,N_1552,N_1116);
or U4835 (N_4835,N_548,N_1268);
and U4836 (N_4836,N_2224,N_2884);
nand U4837 (N_4837,N_364,N_37);
or U4838 (N_4838,N_1012,N_2798);
nand U4839 (N_4839,N_1805,N_1621);
nand U4840 (N_4840,N_1104,N_454);
nor U4841 (N_4841,N_1096,N_2227);
nor U4842 (N_4842,N_2753,N_1314);
xor U4843 (N_4843,N_1429,N_683);
nor U4844 (N_4844,N_1298,N_2431);
nand U4845 (N_4845,N_2798,N_2858);
nor U4846 (N_4846,N_1535,N_483);
or U4847 (N_4847,N_1625,N_847);
nor U4848 (N_4848,N_1937,N_2896);
nand U4849 (N_4849,N_1082,N_39);
or U4850 (N_4850,N_1045,N_1372);
nand U4851 (N_4851,N_715,N_2526);
and U4852 (N_4852,N_1023,N_547);
nand U4853 (N_4853,N_1967,N_903);
nor U4854 (N_4854,N_1598,N_1124);
or U4855 (N_4855,N_1820,N_1299);
nor U4856 (N_4856,N_949,N_1539);
and U4857 (N_4857,N_13,N_2102);
or U4858 (N_4858,N_1758,N_1548);
or U4859 (N_4859,N_1835,N_2510);
and U4860 (N_4860,N_2761,N_1523);
nand U4861 (N_4861,N_1651,N_2148);
xnor U4862 (N_4862,N_2704,N_2894);
and U4863 (N_4863,N_2708,N_1567);
or U4864 (N_4864,N_1320,N_1827);
or U4865 (N_4865,N_2225,N_233);
or U4866 (N_4866,N_180,N_817);
nand U4867 (N_4867,N_2365,N_220);
nor U4868 (N_4868,N_2805,N_2306);
and U4869 (N_4869,N_1945,N_2170);
nand U4870 (N_4870,N_1157,N_1875);
nor U4871 (N_4871,N_2925,N_1038);
nor U4872 (N_4872,N_991,N_1682);
and U4873 (N_4873,N_2486,N_1842);
nand U4874 (N_4874,N_2044,N_2304);
and U4875 (N_4875,N_1134,N_1441);
nand U4876 (N_4876,N_1009,N_113);
or U4877 (N_4877,N_2373,N_279);
and U4878 (N_4878,N_2805,N_1017);
nor U4879 (N_4879,N_2225,N_1578);
nor U4880 (N_4880,N_2865,N_387);
and U4881 (N_4881,N_1359,N_1665);
nand U4882 (N_4882,N_128,N_1097);
nor U4883 (N_4883,N_2723,N_1444);
nand U4884 (N_4884,N_2101,N_1183);
nand U4885 (N_4885,N_2856,N_543);
nand U4886 (N_4886,N_2494,N_1792);
or U4887 (N_4887,N_1974,N_1211);
or U4888 (N_4888,N_1642,N_1989);
and U4889 (N_4889,N_2887,N_1239);
or U4890 (N_4890,N_8,N_2732);
nor U4891 (N_4891,N_43,N_650);
or U4892 (N_4892,N_2671,N_2084);
or U4893 (N_4893,N_1512,N_2030);
or U4894 (N_4894,N_924,N_2475);
nor U4895 (N_4895,N_1759,N_2028);
or U4896 (N_4896,N_1297,N_58);
nor U4897 (N_4897,N_2285,N_2836);
and U4898 (N_4898,N_1466,N_151);
nor U4899 (N_4899,N_2407,N_2259);
or U4900 (N_4900,N_1137,N_2949);
nor U4901 (N_4901,N_2573,N_405);
nor U4902 (N_4902,N_1187,N_2338);
or U4903 (N_4903,N_815,N_2107);
nor U4904 (N_4904,N_506,N_1092);
and U4905 (N_4905,N_293,N_644);
nand U4906 (N_4906,N_527,N_2922);
nand U4907 (N_4907,N_1541,N_2956);
and U4908 (N_4908,N_1586,N_541);
and U4909 (N_4909,N_1056,N_2353);
and U4910 (N_4910,N_1721,N_1892);
and U4911 (N_4911,N_601,N_593);
or U4912 (N_4912,N_834,N_2408);
nand U4913 (N_4913,N_979,N_731);
nand U4914 (N_4914,N_867,N_2624);
nor U4915 (N_4915,N_2986,N_1847);
nor U4916 (N_4916,N_1799,N_542);
nand U4917 (N_4917,N_754,N_727);
or U4918 (N_4918,N_2067,N_153);
nor U4919 (N_4919,N_816,N_1051);
nor U4920 (N_4920,N_2105,N_1771);
nand U4921 (N_4921,N_1904,N_250);
and U4922 (N_4922,N_1616,N_348);
nand U4923 (N_4923,N_823,N_2512);
and U4924 (N_4924,N_720,N_2977);
and U4925 (N_4925,N_1235,N_771);
and U4926 (N_4926,N_2187,N_1332);
nand U4927 (N_4927,N_1034,N_2725);
or U4928 (N_4928,N_2761,N_2094);
nor U4929 (N_4929,N_2822,N_581);
nand U4930 (N_4930,N_2740,N_166);
and U4931 (N_4931,N_1022,N_1004);
nand U4932 (N_4932,N_668,N_1581);
xnor U4933 (N_4933,N_2776,N_2878);
nor U4934 (N_4934,N_2930,N_1482);
nor U4935 (N_4935,N_450,N_910);
and U4936 (N_4936,N_2507,N_2982);
nand U4937 (N_4937,N_900,N_641);
nor U4938 (N_4938,N_2638,N_16);
and U4939 (N_4939,N_1084,N_832);
or U4940 (N_4940,N_1594,N_1994);
nand U4941 (N_4941,N_642,N_1213);
or U4942 (N_4942,N_2544,N_1707);
nand U4943 (N_4943,N_846,N_1215);
nor U4944 (N_4944,N_1233,N_2598);
and U4945 (N_4945,N_1855,N_1873);
nand U4946 (N_4946,N_678,N_2513);
xnor U4947 (N_4947,N_2245,N_2587);
or U4948 (N_4948,N_390,N_125);
nor U4949 (N_4949,N_1305,N_8);
nand U4950 (N_4950,N_744,N_284);
nand U4951 (N_4951,N_1670,N_396);
or U4952 (N_4952,N_1719,N_2910);
nand U4953 (N_4953,N_2803,N_503);
nor U4954 (N_4954,N_271,N_1901);
or U4955 (N_4955,N_1382,N_2735);
nand U4956 (N_4956,N_568,N_2365);
nand U4957 (N_4957,N_1050,N_2957);
nand U4958 (N_4958,N_119,N_616);
or U4959 (N_4959,N_2441,N_2537);
and U4960 (N_4960,N_2658,N_462);
and U4961 (N_4961,N_332,N_1017);
nand U4962 (N_4962,N_750,N_1401);
or U4963 (N_4963,N_52,N_2741);
or U4964 (N_4964,N_1896,N_2989);
nand U4965 (N_4965,N_1936,N_2787);
or U4966 (N_4966,N_1139,N_604);
and U4967 (N_4967,N_659,N_2605);
or U4968 (N_4968,N_2336,N_1319);
nor U4969 (N_4969,N_2296,N_1229);
nor U4970 (N_4970,N_2573,N_235);
and U4971 (N_4971,N_1771,N_224);
nor U4972 (N_4972,N_1921,N_2214);
or U4973 (N_4973,N_1795,N_642);
nand U4974 (N_4974,N_982,N_2027);
or U4975 (N_4975,N_2402,N_2079);
nor U4976 (N_4976,N_2577,N_2002);
and U4977 (N_4977,N_1511,N_2238);
and U4978 (N_4978,N_926,N_1646);
nor U4979 (N_4979,N_423,N_1271);
and U4980 (N_4980,N_2861,N_436);
or U4981 (N_4981,N_1788,N_541);
or U4982 (N_4982,N_2322,N_1226);
nand U4983 (N_4983,N_1524,N_53);
nand U4984 (N_4984,N_897,N_2844);
nand U4985 (N_4985,N_2950,N_637);
or U4986 (N_4986,N_349,N_2390);
and U4987 (N_4987,N_2624,N_2830);
and U4988 (N_4988,N_2907,N_2629);
nand U4989 (N_4989,N_1835,N_2154);
nor U4990 (N_4990,N_2744,N_686);
and U4991 (N_4991,N_2437,N_1002);
xnor U4992 (N_4992,N_498,N_1643);
or U4993 (N_4993,N_2482,N_1689);
nand U4994 (N_4994,N_1265,N_611);
or U4995 (N_4995,N_1592,N_527);
or U4996 (N_4996,N_222,N_2701);
and U4997 (N_4997,N_292,N_1254);
or U4998 (N_4998,N_1101,N_1738);
and U4999 (N_4999,N_285,N_497);
or U5000 (N_5000,N_2124,N_1393);
or U5001 (N_5001,N_1843,N_2082);
or U5002 (N_5002,N_2616,N_1522);
or U5003 (N_5003,N_832,N_897);
or U5004 (N_5004,N_1833,N_848);
or U5005 (N_5005,N_1593,N_305);
nor U5006 (N_5006,N_416,N_404);
nand U5007 (N_5007,N_668,N_2475);
or U5008 (N_5008,N_1251,N_1199);
or U5009 (N_5009,N_611,N_1686);
nand U5010 (N_5010,N_2895,N_1789);
or U5011 (N_5011,N_1617,N_974);
nand U5012 (N_5012,N_121,N_637);
nand U5013 (N_5013,N_2578,N_978);
nor U5014 (N_5014,N_2633,N_1767);
or U5015 (N_5015,N_2706,N_2769);
nand U5016 (N_5016,N_2742,N_1934);
nand U5017 (N_5017,N_1811,N_463);
or U5018 (N_5018,N_1319,N_698);
or U5019 (N_5019,N_514,N_2031);
or U5020 (N_5020,N_1535,N_2512);
and U5021 (N_5021,N_1016,N_925);
and U5022 (N_5022,N_1875,N_1335);
and U5023 (N_5023,N_1860,N_202);
or U5024 (N_5024,N_2581,N_1462);
nand U5025 (N_5025,N_2286,N_1428);
nand U5026 (N_5026,N_614,N_2366);
or U5027 (N_5027,N_1008,N_1784);
nand U5028 (N_5028,N_2351,N_756);
and U5029 (N_5029,N_1499,N_1730);
or U5030 (N_5030,N_2741,N_1131);
and U5031 (N_5031,N_1941,N_2247);
or U5032 (N_5032,N_2754,N_1383);
or U5033 (N_5033,N_1823,N_658);
and U5034 (N_5034,N_2701,N_2155);
nand U5035 (N_5035,N_1615,N_1193);
and U5036 (N_5036,N_1655,N_568);
xor U5037 (N_5037,N_997,N_616);
and U5038 (N_5038,N_1715,N_2613);
nor U5039 (N_5039,N_1589,N_1220);
nand U5040 (N_5040,N_1859,N_166);
and U5041 (N_5041,N_2893,N_1290);
and U5042 (N_5042,N_1702,N_1454);
nand U5043 (N_5043,N_2458,N_521);
nor U5044 (N_5044,N_2968,N_2987);
and U5045 (N_5045,N_2820,N_1762);
or U5046 (N_5046,N_51,N_2947);
and U5047 (N_5047,N_545,N_782);
and U5048 (N_5048,N_2206,N_1907);
nand U5049 (N_5049,N_1751,N_391);
or U5050 (N_5050,N_906,N_1735);
or U5051 (N_5051,N_2709,N_1863);
and U5052 (N_5052,N_299,N_2853);
or U5053 (N_5053,N_359,N_1142);
and U5054 (N_5054,N_502,N_2729);
nor U5055 (N_5055,N_2288,N_715);
and U5056 (N_5056,N_542,N_290);
or U5057 (N_5057,N_1536,N_106);
or U5058 (N_5058,N_1440,N_2743);
nor U5059 (N_5059,N_958,N_2338);
nand U5060 (N_5060,N_1614,N_1834);
nand U5061 (N_5061,N_2714,N_2070);
or U5062 (N_5062,N_1188,N_1385);
or U5063 (N_5063,N_117,N_1589);
or U5064 (N_5064,N_2569,N_1117);
and U5065 (N_5065,N_1971,N_2055);
nor U5066 (N_5066,N_2567,N_199);
or U5067 (N_5067,N_1147,N_2703);
nor U5068 (N_5068,N_2595,N_189);
nand U5069 (N_5069,N_1499,N_277);
and U5070 (N_5070,N_1744,N_1895);
nor U5071 (N_5071,N_1721,N_576);
nor U5072 (N_5072,N_2545,N_2823);
nor U5073 (N_5073,N_460,N_1758);
or U5074 (N_5074,N_1414,N_1630);
nor U5075 (N_5075,N_2885,N_2460);
or U5076 (N_5076,N_1824,N_1992);
or U5077 (N_5077,N_2200,N_2525);
or U5078 (N_5078,N_758,N_830);
and U5079 (N_5079,N_2940,N_2570);
or U5080 (N_5080,N_2534,N_2572);
xnor U5081 (N_5081,N_1844,N_1266);
and U5082 (N_5082,N_1799,N_1780);
and U5083 (N_5083,N_2187,N_43);
nor U5084 (N_5084,N_371,N_2637);
or U5085 (N_5085,N_238,N_1465);
or U5086 (N_5086,N_2209,N_1085);
or U5087 (N_5087,N_1946,N_1464);
and U5088 (N_5088,N_1126,N_1890);
nand U5089 (N_5089,N_824,N_1342);
nor U5090 (N_5090,N_993,N_2355);
nor U5091 (N_5091,N_2203,N_1770);
and U5092 (N_5092,N_944,N_2553);
and U5093 (N_5093,N_2768,N_2467);
and U5094 (N_5094,N_412,N_2878);
or U5095 (N_5095,N_2502,N_2983);
and U5096 (N_5096,N_1829,N_2199);
nand U5097 (N_5097,N_421,N_2653);
or U5098 (N_5098,N_1890,N_1421);
nor U5099 (N_5099,N_2870,N_1698);
or U5100 (N_5100,N_2464,N_1520);
nand U5101 (N_5101,N_491,N_2585);
and U5102 (N_5102,N_2291,N_1061);
nor U5103 (N_5103,N_605,N_248);
nand U5104 (N_5104,N_1609,N_2493);
nand U5105 (N_5105,N_1352,N_469);
nor U5106 (N_5106,N_1721,N_2662);
nand U5107 (N_5107,N_547,N_372);
or U5108 (N_5108,N_1111,N_1447);
or U5109 (N_5109,N_1546,N_58);
and U5110 (N_5110,N_1215,N_20);
nor U5111 (N_5111,N_1540,N_2864);
nor U5112 (N_5112,N_379,N_2626);
nor U5113 (N_5113,N_2313,N_2544);
xnor U5114 (N_5114,N_2038,N_2499);
nor U5115 (N_5115,N_357,N_2319);
or U5116 (N_5116,N_372,N_946);
nand U5117 (N_5117,N_1188,N_2755);
nor U5118 (N_5118,N_1918,N_1050);
or U5119 (N_5119,N_2982,N_1748);
nand U5120 (N_5120,N_2643,N_470);
and U5121 (N_5121,N_2616,N_2865);
nand U5122 (N_5122,N_549,N_1399);
nor U5123 (N_5123,N_754,N_2674);
nor U5124 (N_5124,N_556,N_1590);
nand U5125 (N_5125,N_406,N_2445);
nor U5126 (N_5126,N_1187,N_2172);
nand U5127 (N_5127,N_1095,N_2283);
or U5128 (N_5128,N_400,N_2044);
or U5129 (N_5129,N_2113,N_2698);
xor U5130 (N_5130,N_2610,N_2504);
and U5131 (N_5131,N_494,N_2144);
nand U5132 (N_5132,N_2401,N_1430);
nor U5133 (N_5133,N_2781,N_2239);
or U5134 (N_5134,N_2495,N_890);
nor U5135 (N_5135,N_1447,N_412);
nand U5136 (N_5136,N_1309,N_1210);
and U5137 (N_5137,N_2990,N_2863);
or U5138 (N_5138,N_758,N_1768);
nand U5139 (N_5139,N_1571,N_321);
nand U5140 (N_5140,N_143,N_1036);
and U5141 (N_5141,N_2409,N_42);
and U5142 (N_5142,N_2171,N_1928);
and U5143 (N_5143,N_897,N_1613);
nand U5144 (N_5144,N_301,N_2573);
or U5145 (N_5145,N_604,N_2793);
nand U5146 (N_5146,N_2711,N_431);
or U5147 (N_5147,N_2369,N_292);
or U5148 (N_5148,N_625,N_1569);
nor U5149 (N_5149,N_839,N_1272);
nand U5150 (N_5150,N_1471,N_46);
nor U5151 (N_5151,N_1113,N_2186);
nand U5152 (N_5152,N_2697,N_2449);
or U5153 (N_5153,N_1147,N_760);
and U5154 (N_5154,N_1302,N_183);
or U5155 (N_5155,N_713,N_1974);
or U5156 (N_5156,N_1247,N_748);
or U5157 (N_5157,N_780,N_1955);
nor U5158 (N_5158,N_222,N_2188);
nand U5159 (N_5159,N_1159,N_2104);
or U5160 (N_5160,N_2121,N_2501);
nor U5161 (N_5161,N_1734,N_1694);
nand U5162 (N_5162,N_790,N_920);
and U5163 (N_5163,N_21,N_2342);
or U5164 (N_5164,N_1708,N_373);
or U5165 (N_5165,N_1767,N_2185);
and U5166 (N_5166,N_2247,N_506);
nand U5167 (N_5167,N_2171,N_2409);
or U5168 (N_5168,N_2576,N_2763);
nor U5169 (N_5169,N_2000,N_270);
xor U5170 (N_5170,N_2118,N_1430);
and U5171 (N_5171,N_2770,N_75);
nand U5172 (N_5172,N_2707,N_140);
and U5173 (N_5173,N_2881,N_339);
nor U5174 (N_5174,N_1359,N_870);
or U5175 (N_5175,N_2055,N_316);
and U5176 (N_5176,N_1079,N_1690);
and U5177 (N_5177,N_723,N_579);
nor U5178 (N_5178,N_159,N_367);
xor U5179 (N_5179,N_1214,N_2870);
or U5180 (N_5180,N_850,N_1688);
nand U5181 (N_5181,N_1649,N_239);
and U5182 (N_5182,N_112,N_1370);
or U5183 (N_5183,N_2603,N_1607);
nor U5184 (N_5184,N_1109,N_755);
and U5185 (N_5185,N_1084,N_2207);
nor U5186 (N_5186,N_1306,N_1881);
nor U5187 (N_5187,N_636,N_2896);
nand U5188 (N_5188,N_2164,N_923);
and U5189 (N_5189,N_1139,N_2645);
and U5190 (N_5190,N_2640,N_1283);
nand U5191 (N_5191,N_445,N_1233);
or U5192 (N_5192,N_423,N_903);
nand U5193 (N_5193,N_1159,N_607);
and U5194 (N_5194,N_67,N_2795);
nor U5195 (N_5195,N_2399,N_1347);
nand U5196 (N_5196,N_2025,N_1761);
nor U5197 (N_5197,N_1737,N_513);
nor U5198 (N_5198,N_2810,N_24);
nor U5199 (N_5199,N_1578,N_40);
nor U5200 (N_5200,N_776,N_699);
or U5201 (N_5201,N_1904,N_1366);
and U5202 (N_5202,N_1358,N_2430);
or U5203 (N_5203,N_460,N_2789);
nand U5204 (N_5204,N_85,N_1979);
or U5205 (N_5205,N_2316,N_511);
nand U5206 (N_5206,N_2691,N_1600);
nor U5207 (N_5207,N_1585,N_1867);
or U5208 (N_5208,N_683,N_717);
and U5209 (N_5209,N_1206,N_2495);
nand U5210 (N_5210,N_2361,N_1289);
nand U5211 (N_5211,N_2408,N_327);
nand U5212 (N_5212,N_2536,N_873);
nor U5213 (N_5213,N_2638,N_2632);
nand U5214 (N_5214,N_985,N_2212);
nor U5215 (N_5215,N_1100,N_626);
nor U5216 (N_5216,N_482,N_2980);
nor U5217 (N_5217,N_2739,N_704);
xor U5218 (N_5218,N_1370,N_1850);
nand U5219 (N_5219,N_1922,N_608);
and U5220 (N_5220,N_1829,N_846);
nand U5221 (N_5221,N_1457,N_506);
nor U5222 (N_5222,N_2505,N_2397);
nand U5223 (N_5223,N_2164,N_911);
nand U5224 (N_5224,N_2530,N_1446);
or U5225 (N_5225,N_928,N_510);
and U5226 (N_5226,N_1460,N_1696);
nor U5227 (N_5227,N_138,N_2019);
nor U5228 (N_5228,N_2830,N_1583);
or U5229 (N_5229,N_397,N_942);
nor U5230 (N_5230,N_2017,N_2628);
and U5231 (N_5231,N_2542,N_2887);
nand U5232 (N_5232,N_366,N_2074);
and U5233 (N_5233,N_2987,N_1992);
or U5234 (N_5234,N_429,N_1605);
or U5235 (N_5235,N_742,N_2362);
and U5236 (N_5236,N_688,N_269);
or U5237 (N_5237,N_1276,N_2742);
and U5238 (N_5238,N_1600,N_275);
nand U5239 (N_5239,N_1601,N_121);
and U5240 (N_5240,N_2344,N_136);
or U5241 (N_5241,N_2581,N_2270);
or U5242 (N_5242,N_1380,N_1776);
nor U5243 (N_5243,N_2425,N_2062);
nand U5244 (N_5244,N_1046,N_603);
nand U5245 (N_5245,N_2144,N_1172);
or U5246 (N_5246,N_2902,N_473);
or U5247 (N_5247,N_2408,N_288);
and U5248 (N_5248,N_600,N_181);
or U5249 (N_5249,N_2019,N_60);
or U5250 (N_5250,N_1965,N_63);
and U5251 (N_5251,N_2156,N_824);
or U5252 (N_5252,N_1150,N_110);
nand U5253 (N_5253,N_2705,N_2485);
nor U5254 (N_5254,N_1849,N_1416);
or U5255 (N_5255,N_122,N_2525);
nor U5256 (N_5256,N_1796,N_2679);
nor U5257 (N_5257,N_2563,N_625);
nand U5258 (N_5258,N_2111,N_1798);
nor U5259 (N_5259,N_53,N_2228);
or U5260 (N_5260,N_1837,N_2587);
and U5261 (N_5261,N_2369,N_788);
and U5262 (N_5262,N_614,N_1006);
and U5263 (N_5263,N_1200,N_95);
or U5264 (N_5264,N_410,N_1964);
or U5265 (N_5265,N_1325,N_2978);
or U5266 (N_5266,N_2672,N_742);
nand U5267 (N_5267,N_215,N_782);
or U5268 (N_5268,N_162,N_1238);
nand U5269 (N_5269,N_895,N_649);
nand U5270 (N_5270,N_218,N_242);
nor U5271 (N_5271,N_881,N_310);
nand U5272 (N_5272,N_1953,N_2221);
nand U5273 (N_5273,N_738,N_2942);
nand U5274 (N_5274,N_134,N_980);
nor U5275 (N_5275,N_2336,N_308);
nand U5276 (N_5276,N_1003,N_56);
nand U5277 (N_5277,N_2749,N_338);
nor U5278 (N_5278,N_2380,N_2246);
nand U5279 (N_5279,N_1230,N_879);
nor U5280 (N_5280,N_933,N_1328);
and U5281 (N_5281,N_1463,N_2006);
and U5282 (N_5282,N_887,N_2519);
nor U5283 (N_5283,N_575,N_1941);
or U5284 (N_5284,N_453,N_1646);
or U5285 (N_5285,N_2995,N_2489);
and U5286 (N_5286,N_2132,N_2245);
nand U5287 (N_5287,N_2584,N_2077);
and U5288 (N_5288,N_2062,N_1247);
nand U5289 (N_5289,N_668,N_1059);
xnor U5290 (N_5290,N_205,N_400);
and U5291 (N_5291,N_2366,N_2898);
nor U5292 (N_5292,N_2488,N_1190);
nor U5293 (N_5293,N_1684,N_504);
nand U5294 (N_5294,N_2721,N_973);
nand U5295 (N_5295,N_2425,N_2561);
or U5296 (N_5296,N_1976,N_2546);
nand U5297 (N_5297,N_1366,N_2508);
and U5298 (N_5298,N_1884,N_1393);
or U5299 (N_5299,N_736,N_1572);
and U5300 (N_5300,N_2987,N_2790);
or U5301 (N_5301,N_2134,N_2517);
nor U5302 (N_5302,N_10,N_2078);
nand U5303 (N_5303,N_804,N_903);
nand U5304 (N_5304,N_564,N_2858);
and U5305 (N_5305,N_672,N_1673);
or U5306 (N_5306,N_2971,N_1110);
or U5307 (N_5307,N_973,N_2519);
or U5308 (N_5308,N_1337,N_119);
xnor U5309 (N_5309,N_1396,N_245);
or U5310 (N_5310,N_507,N_780);
and U5311 (N_5311,N_2357,N_644);
and U5312 (N_5312,N_2981,N_705);
and U5313 (N_5313,N_58,N_1481);
nand U5314 (N_5314,N_373,N_580);
nor U5315 (N_5315,N_1130,N_2550);
or U5316 (N_5316,N_2172,N_2892);
nand U5317 (N_5317,N_1508,N_2506);
or U5318 (N_5318,N_551,N_2222);
nor U5319 (N_5319,N_2484,N_2216);
and U5320 (N_5320,N_2175,N_585);
xor U5321 (N_5321,N_1449,N_1564);
or U5322 (N_5322,N_2022,N_2688);
nand U5323 (N_5323,N_2261,N_919);
and U5324 (N_5324,N_2511,N_2010);
and U5325 (N_5325,N_170,N_580);
nand U5326 (N_5326,N_1835,N_2803);
nor U5327 (N_5327,N_2857,N_2301);
nor U5328 (N_5328,N_2020,N_1837);
and U5329 (N_5329,N_2933,N_1509);
nand U5330 (N_5330,N_1721,N_642);
and U5331 (N_5331,N_2666,N_344);
nand U5332 (N_5332,N_2412,N_2370);
nor U5333 (N_5333,N_2425,N_1527);
nor U5334 (N_5334,N_1700,N_1507);
and U5335 (N_5335,N_1658,N_2034);
nand U5336 (N_5336,N_793,N_2821);
or U5337 (N_5337,N_320,N_2314);
nand U5338 (N_5338,N_517,N_2337);
and U5339 (N_5339,N_1532,N_1792);
or U5340 (N_5340,N_1518,N_1207);
nor U5341 (N_5341,N_1365,N_2472);
or U5342 (N_5342,N_176,N_1107);
xor U5343 (N_5343,N_458,N_2658);
or U5344 (N_5344,N_1241,N_2054);
nor U5345 (N_5345,N_58,N_1083);
nand U5346 (N_5346,N_1075,N_1334);
nor U5347 (N_5347,N_2973,N_196);
nand U5348 (N_5348,N_1086,N_2563);
nor U5349 (N_5349,N_2321,N_1861);
nor U5350 (N_5350,N_1932,N_1752);
and U5351 (N_5351,N_457,N_1473);
nand U5352 (N_5352,N_1249,N_135);
and U5353 (N_5353,N_122,N_1735);
and U5354 (N_5354,N_856,N_1344);
nor U5355 (N_5355,N_1117,N_2918);
nand U5356 (N_5356,N_304,N_2672);
nor U5357 (N_5357,N_2741,N_1448);
nor U5358 (N_5358,N_321,N_2649);
and U5359 (N_5359,N_447,N_2431);
and U5360 (N_5360,N_275,N_2439);
nor U5361 (N_5361,N_2601,N_1719);
nand U5362 (N_5362,N_2607,N_1981);
and U5363 (N_5363,N_1985,N_2196);
nor U5364 (N_5364,N_2153,N_2546);
or U5365 (N_5365,N_844,N_336);
or U5366 (N_5366,N_567,N_2445);
nand U5367 (N_5367,N_1246,N_651);
nor U5368 (N_5368,N_2385,N_1462);
and U5369 (N_5369,N_1010,N_1642);
nor U5370 (N_5370,N_1235,N_816);
nand U5371 (N_5371,N_89,N_2450);
nor U5372 (N_5372,N_578,N_2920);
nand U5373 (N_5373,N_1146,N_1105);
nor U5374 (N_5374,N_2717,N_2559);
or U5375 (N_5375,N_763,N_2191);
nand U5376 (N_5376,N_1487,N_1514);
nor U5377 (N_5377,N_287,N_617);
nand U5378 (N_5378,N_2911,N_1399);
and U5379 (N_5379,N_2950,N_877);
nand U5380 (N_5380,N_2575,N_544);
nor U5381 (N_5381,N_1775,N_57);
or U5382 (N_5382,N_950,N_8);
and U5383 (N_5383,N_858,N_2745);
or U5384 (N_5384,N_2420,N_712);
nand U5385 (N_5385,N_2109,N_422);
nor U5386 (N_5386,N_2063,N_1299);
and U5387 (N_5387,N_2187,N_2119);
nand U5388 (N_5388,N_420,N_2771);
or U5389 (N_5389,N_1350,N_1184);
and U5390 (N_5390,N_2317,N_993);
or U5391 (N_5391,N_1717,N_2443);
or U5392 (N_5392,N_699,N_541);
nor U5393 (N_5393,N_2950,N_927);
nand U5394 (N_5394,N_2503,N_1569);
nor U5395 (N_5395,N_2962,N_2024);
and U5396 (N_5396,N_1446,N_2252);
nor U5397 (N_5397,N_2251,N_1223);
nand U5398 (N_5398,N_1397,N_1264);
or U5399 (N_5399,N_1364,N_661);
nor U5400 (N_5400,N_2945,N_2368);
nor U5401 (N_5401,N_1924,N_2228);
nor U5402 (N_5402,N_2410,N_2158);
nand U5403 (N_5403,N_879,N_311);
and U5404 (N_5404,N_2789,N_283);
and U5405 (N_5405,N_1265,N_816);
or U5406 (N_5406,N_257,N_2130);
nor U5407 (N_5407,N_825,N_1038);
nand U5408 (N_5408,N_633,N_1373);
nor U5409 (N_5409,N_102,N_1687);
nor U5410 (N_5410,N_1070,N_734);
and U5411 (N_5411,N_2141,N_2108);
nand U5412 (N_5412,N_297,N_2075);
or U5413 (N_5413,N_1289,N_1955);
nor U5414 (N_5414,N_510,N_1984);
and U5415 (N_5415,N_438,N_782);
or U5416 (N_5416,N_1251,N_1911);
nand U5417 (N_5417,N_2275,N_732);
xor U5418 (N_5418,N_2135,N_2492);
or U5419 (N_5419,N_2042,N_1446);
xor U5420 (N_5420,N_352,N_2123);
and U5421 (N_5421,N_2336,N_1949);
nand U5422 (N_5422,N_1856,N_2031);
or U5423 (N_5423,N_449,N_516);
nand U5424 (N_5424,N_1628,N_1037);
nand U5425 (N_5425,N_1556,N_2091);
nor U5426 (N_5426,N_800,N_1368);
and U5427 (N_5427,N_1314,N_1377);
nor U5428 (N_5428,N_2716,N_448);
or U5429 (N_5429,N_910,N_2336);
nor U5430 (N_5430,N_2669,N_1916);
and U5431 (N_5431,N_2127,N_2857);
nor U5432 (N_5432,N_2625,N_36);
and U5433 (N_5433,N_488,N_1882);
nor U5434 (N_5434,N_1663,N_1888);
and U5435 (N_5435,N_178,N_1135);
and U5436 (N_5436,N_2813,N_2292);
and U5437 (N_5437,N_1515,N_352);
nor U5438 (N_5438,N_174,N_2669);
and U5439 (N_5439,N_652,N_2679);
and U5440 (N_5440,N_571,N_63);
or U5441 (N_5441,N_1831,N_825);
and U5442 (N_5442,N_1106,N_1418);
or U5443 (N_5443,N_163,N_1169);
nor U5444 (N_5444,N_175,N_2677);
nand U5445 (N_5445,N_1901,N_2834);
and U5446 (N_5446,N_1030,N_2656);
nor U5447 (N_5447,N_2971,N_1355);
nor U5448 (N_5448,N_459,N_131);
nor U5449 (N_5449,N_1872,N_1481);
nand U5450 (N_5450,N_1501,N_2115);
nand U5451 (N_5451,N_2576,N_1258);
or U5452 (N_5452,N_1108,N_1776);
or U5453 (N_5453,N_239,N_584);
and U5454 (N_5454,N_1534,N_2934);
nor U5455 (N_5455,N_320,N_2086);
and U5456 (N_5456,N_1561,N_2366);
or U5457 (N_5457,N_2869,N_235);
nand U5458 (N_5458,N_889,N_2154);
and U5459 (N_5459,N_480,N_2442);
nand U5460 (N_5460,N_1462,N_2608);
or U5461 (N_5461,N_1354,N_2373);
nand U5462 (N_5462,N_2211,N_1647);
nand U5463 (N_5463,N_2997,N_1835);
or U5464 (N_5464,N_2384,N_123);
and U5465 (N_5465,N_2985,N_422);
nand U5466 (N_5466,N_600,N_2204);
or U5467 (N_5467,N_996,N_222);
and U5468 (N_5468,N_1427,N_824);
or U5469 (N_5469,N_1878,N_57);
nand U5470 (N_5470,N_1983,N_1511);
nor U5471 (N_5471,N_2313,N_1062);
nand U5472 (N_5472,N_296,N_1648);
nor U5473 (N_5473,N_258,N_1366);
or U5474 (N_5474,N_1950,N_893);
nor U5475 (N_5475,N_389,N_1976);
or U5476 (N_5476,N_642,N_1665);
xnor U5477 (N_5477,N_2342,N_1492);
nor U5478 (N_5478,N_1330,N_240);
nor U5479 (N_5479,N_723,N_2363);
nand U5480 (N_5480,N_762,N_1273);
and U5481 (N_5481,N_1174,N_158);
or U5482 (N_5482,N_2801,N_2177);
or U5483 (N_5483,N_1698,N_339);
or U5484 (N_5484,N_2092,N_709);
nand U5485 (N_5485,N_81,N_122);
or U5486 (N_5486,N_2374,N_2510);
nand U5487 (N_5487,N_1585,N_1392);
nand U5488 (N_5488,N_2032,N_197);
and U5489 (N_5489,N_2550,N_2119);
or U5490 (N_5490,N_2250,N_223);
nor U5491 (N_5491,N_1214,N_538);
and U5492 (N_5492,N_2483,N_2013);
nand U5493 (N_5493,N_2623,N_140);
and U5494 (N_5494,N_412,N_1377);
xnor U5495 (N_5495,N_2588,N_1467);
and U5496 (N_5496,N_1770,N_1654);
and U5497 (N_5497,N_2793,N_1852);
and U5498 (N_5498,N_104,N_885);
or U5499 (N_5499,N_290,N_2487);
or U5500 (N_5500,N_961,N_144);
nand U5501 (N_5501,N_1424,N_275);
nor U5502 (N_5502,N_2260,N_451);
and U5503 (N_5503,N_2789,N_389);
nor U5504 (N_5504,N_855,N_1061);
or U5505 (N_5505,N_1251,N_1436);
nand U5506 (N_5506,N_1771,N_566);
nand U5507 (N_5507,N_2388,N_518);
nor U5508 (N_5508,N_2421,N_1963);
and U5509 (N_5509,N_334,N_1355);
nand U5510 (N_5510,N_867,N_1398);
nand U5511 (N_5511,N_278,N_534);
nor U5512 (N_5512,N_2426,N_881);
and U5513 (N_5513,N_2358,N_550);
nand U5514 (N_5514,N_1376,N_2915);
and U5515 (N_5515,N_979,N_1506);
and U5516 (N_5516,N_1350,N_2546);
or U5517 (N_5517,N_344,N_2396);
or U5518 (N_5518,N_302,N_1166);
nor U5519 (N_5519,N_993,N_2838);
or U5520 (N_5520,N_1664,N_2035);
nand U5521 (N_5521,N_1782,N_2000);
nor U5522 (N_5522,N_1830,N_2637);
or U5523 (N_5523,N_2889,N_863);
nor U5524 (N_5524,N_942,N_1813);
and U5525 (N_5525,N_2121,N_308);
nor U5526 (N_5526,N_817,N_919);
nand U5527 (N_5527,N_2256,N_1794);
and U5528 (N_5528,N_1445,N_921);
and U5529 (N_5529,N_2345,N_48);
nand U5530 (N_5530,N_1218,N_143);
and U5531 (N_5531,N_33,N_2418);
nand U5532 (N_5532,N_2248,N_1890);
nor U5533 (N_5533,N_451,N_2065);
or U5534 (N_5534,N_0,N_939);
or U5535 (N_5535,N_1097,N_874);
nor U5536 (N_5536,N_493,N_2212);
nand U5537 (N_5537,N_519,N_981);
or U5538 (N_5538,N_1956,N_152);
or U5539 (N_5539,N_2294,N_708);
nand U5540 (N_5540,N_243,N_515);
and U5541 (N_5541,N_570,N_2852);
nor U5542 (N_5542,N_2835,N_2585);
nand U5543 (N_5543,N_569,N_2960);
nand U5544 (N_5544,N_1936,N_1743);
or U5545 (N_5545,N_1545,N_1926);
nor U5546 (N_5546,N_1981,N_1005);
nand U5547 (N_5547,N_1650,N_2958);
nand U5548 (N_5548,N_1333,N_2463);
nand U5549 (N_5549,N_1144,N_809);
xnor U5550 (N_5550,N_2690,N_1893);
nand U5551 (N_5551,N_1145,N_2013);
and U5552 (N_5552,N_939,N_844);
or U5553 (N_5553,N_1910,N_1759);
and U5554 (N_5554,N_1172,N_1859);
nand U5555 (N_5555,N_2526,N_1834);
or U5556 (N_5556,N_185,N_375);
or U5557 (N_5557,N_163,N_2337);
nor U5558 (N_5558,N_1123,N_2700);
nand U5559 (N_5559,N_2517,N_2100);
nand U5560 (N_5560,N_287,N_2115);
nand U5561 (N_5561,N_574,N_67);
nand U5562 (N_5562,N_634,N_1961);
nand U5563 (N_5563,N_522,N_1254);
nor U5564 (N_5564,N_2838,N_657);
or U5565 (N_5565,N_2613,N_2731);
or U5566 (N_5566,N_1110,N_2588);
nand U5567 (N_5567,N_1973,N_1794);
and U5568 (N_5568,N_2565,N_1165);
xnor U5569 (N_5569,N_422,N_842);
and U5570 (N_5570,N_1118,N_8);
nand U5571 (N_5571,N_56,N_252);
and U5572 (N_5572,N_154,N_688);
or U5573 (N_5573,N_1340,N_2022);
or U5574 (N_5574,N_1731,N_198);
nand U5575 (N_5575,N_923,N_347);
or U5576 (N_5576,N_153,N_1953);
or U5577 (N_5577,N_1207,N_899);
nor U5578 (N_5578,N_1808,N_130);
xnor U5579 (N_5579,N_4,N_2767);
and U5580 (N_5580,N_2269,N_223);
nand U5581 (N_5581,N_337,N_1679);
or U5582 (N_5582,N_325,N_1679);
xor U5583 (N_5583,N_111,N_2972);
nand U5584 (N_5584,N_2649,N_2315);
nor U5585 (N_5585,N_1458,N_243);
nor U5586 (N_5586,N_1124,N_1894);
nand U5587 (N_5587,N_2152,N_1839);
and U5588 (N_5588,N_1525,N_522);
nor U5589 (N_5589,N_713,N_2234);
or U5590 (N_5590,N_2898,N_2655);
or U5591 (N_5591,N_1349,N_1234);
nand U5592 (N_5592,N_144,N_1582);
or U5593 (N_5593,N_2654,N_1797);
and U5594 (N_5594,N_2138,N_1774);
nor U5595 (N_5595,N_287,N_2813);
nand U5596 (N_5596,N_1559,N_1123);
nand U5597 (N_5597,N_1357,N_71);
or U5598 (N_5598,N_1856,N_2558);
or U5599 (N_5599,N_2464,N_353);
nand U5600 (N_5600,N_1491,N_1315);
nand U5601 (N_5601,N_1571,N_165);
and U5602 (N_5602,N_1830,N_127);
or U5603 (N_5603,N_2051,N_2323);
and U5604 (N_5604,N_677,N_665);
nor U5605 (N_5605,N_2978,N_981);
nand U5606 (N_5606,N_2309,N_1669);
nor U5607 (N_5607,N_2079,N_2762);
nor U5608 (N_5608,N_502,N_2596);
and U5609 (N_5609,N_2294,N_2232);
nand U5610 (N_5610,N_294,N_2148);
nor U5611 (N_5611,N_1080,N_1789);
nor U5612 (N_5612,N_2086,N_2474);
or U5613 (N_5613,N_1473,N_658);
nand U5614 (N_5614,N_1157,N_1371);
nor U5615 (N_5615,N_2899,N_1998);
nor U5616 (N_5616,N_2750,N_2479);
and U5617 (N_5617,N_334,N_1146);
and U5618 (N_5618,N_1813,N_445);
nand U5619 (N_5619,N_124,N_87);
and U5620 (N_5620,N_724,N_510);
nor U5621 (N_5621,N_210,N_527);
nand U5622 (N_5622,N_55,N_604);
or U5623 (N_5623,N_2118,N_1566);
nor U5624 (N_5624,N_1009,N_2992);
nand U5625 (N_5625,N_552,N_1265);
or U5626 (N_5626,N_1261,N_456);
nand U5627 (N_5627,N_419,N_1817);
nand U5628 (N_5628,N_352,N_2485);
nand U5629 (N_5629,N_2682,N_860);
or U5630 (N_5630,N_2877,N_988);
or U5631 (N_5631,N_2775,N_1618);
nand U5632 (N_5632,N_1687,N_260);
nand U5633 (N_5633,N_672,N_2964);
nand U5634 (N_5634,N_850,N_401);
nor U5635 (N_5635,N_1303,N_670);
nor U5636 (N_5636,N_1402,N_393);
nor U5637 (N_5637,N_1917,N_392);
or U5638 (N_5638,N_942,N_1198);
and U5639 (N_5639,N_1558,N_896);
nand U5640 (N_5640,N_2030,N_840);
nor U5641 (N_5641,N_231,N_2151);
nand U5642 (N_5642,N_1967,N_698);
and U5643 (N_5643,N_1082,N_2333);
and U5644 (N_5644,N_664,N_472);
nand U5645 (N_5645,N_1985,N_2157);
or U5646 (N_5646,N_861,N_2325);
nor U5647 (N_5647,N_2922,N_2157);
or U5648 (N_5648,N_52,N_1493);
or U5649 (N_5649,N_1661,N_1060);
nor U5650 (N_5650,N_473,N_878);
nand U5651 (N_5651,N_1907,N_331);
nand U5652 (N_5652,N_1061,N_2668);
and U5653 (N_5653,N_2113,N_2633);
nand U5654 (N_5654,N_495,N_2479);
nand U5655 (N_5655,N_1828,N_269);
nor U5656 (N_5656,N_1985,N_2232);
or U5657 (N_5657,N_1057,N_1134);
nand U5658 (N_5658,N_2231,N_2531);
or U5659 (N_5659,N_1816,N_2603);
nor U5660 (N_5660,N_307,N_650);
or U5661 (N_5661,N_905,N_2487);
nor U5662 (N_5662,N_1333,N_2286);
and U5663 (N_5663,N_1340,N_348);
or U5664 (N_5664,N_540,N_1860);
nor U5665 (N_5665,N_1897,N_1855);
nand U5666 (N_5666,N_1593,N_1165);
and U5667 (N_5667,N_2962,N_1874);
nor U5668 (N_5668,N_899,N_683);
and U5669 (N_5669,N_1115,N_865);
or U5670 (N_5670,N_1258,N_1173);
nand U5671 (N_5671,N_2808,N_2332);
nor U5672 (N_5672,N_916,N_1386);
nor U5673 (N_5673,N_1354,N_955);
nand U5674 (N_5674,N_2168,N_1760);
nor U5675 (N_5675,N_1168,N_1932);
and U5676 (N_5676,N_1210,N_1246);
and U5677 (N_5677,N_1242,N_1384);
nor U5678 (N_5678,N_977,N_836);
or U5679 (N_5679,N_1448,N_2988);
nor U5680 (N_5680,N_494,N_1552);
and U5681 (N_5681,N_1892,N_1656);
nor U5682 (N_5682,N_981,N_1109);
or U5683 (N_5683,N_1801,N_292);
and U5684 (N_5684,N_224,N_379);
nand U5685 (N_5685,N_581,N_2782);
nor U5686 (N_5686,N_305,N_1922);
or U5687 (N_5687,N_2094,N_1073);
and U5688 (N_5688,N_2127,N_2242);
nand U5689 (N_5689,N_437,N_1059);
nand U5690 (N_5690,N_57,N_289);
nand U5691 (N_5691,N_2274,N_582);
nor U5692 (N_5692,N_1117,N_2219);
or U5693 (N_5693,N_2070,N_631);
and U5694 (N_5694,N_2814,N_2078);
nand U5695 (N_5695,N_1317,N_2099);
xor U5696 (N_5696,N_1152,N_1682);
nor U5697 (N_5697,N_87,N_286);
nor U5698 (N_5698,N_1625,N_1527);
or U5699 (N_5699,N_331,N_1822);
nand U5700 (N_5700,N_1910,N_1514);
or U5701 (N_5701,N_2854,N_688);
or U5702 (N_5702,N_2079,N_1161);
nor U5703 (N_5703,N_2303,N_1286);
and U5704 (N_5704,N_1083,N_659);
nand U5705 (N_5705,N_1820,N_2920);
or U5706 (N_5706,N_2995,N_442);
or U5707 (N_5707,N_266,N_2935);
nor U5708 (N_5708,N_820,N_493);
nor U5709 (N_5709,N_275,N_120);
nor U5710 (N_5710,N_866,N_2802);
nand U5711 (N_5711,N_349,N_2128);
or U5712 (N_5712,N_1824,N_343);
nand U5713 (N_5713,N_2403,N_274);
and U5714 (N_5714,N_1852,N_2828);
nand U5715 (N_5715,N_52,N_994);
nand U5716 (N_5716,N_311,N_719);
nand U5717 (N_5717,N_1310,N_830);
or U5718 (N_5718,N_2331,N_329);
or U5719 (N_5719,N_1806,N_2882);
nor U5720 (N_5720,N_846,N_1619);
nand U5721 (N_5721,N_2481,N_24);
or U5722 (N_5722,N_1439,N_911);
nor U5723 (N_5723,N_2750,N_2843);
nand U5724 (N_5724,N_2875,N_2913);
and U5725 (N_5725,N_1625,N_1059);
nor U5726 (N_5726,N_1473,N_178);
or U5727 (N_5727,N_338,N_2072);
or U5728 (N_5728,N_1526,N_2117);
nor U5729 (N_5729,N_455,N_2893);
or U5730 (N_5730,N_2056,N_2011);
and U5731 (N_5731,N_2795,N_1271);
or U5732 (N_5732,N_184,N_654);
nand U5733 (N_5733,N_2775,N_308);
and U5734 (N_5734,N_937,N_532);
nand U5735 (N_5735,N_763,N_1197);
nor U5736 (N_5736,N_1257,N_2017);
or U5737 (N_5737,N_167,N_138);
nor U5738 (N_5738,N_1597,N_2112);
and U5739 (N_5739,N_2740,N_209);
nand U5740 (N_5740,N_1524,N_241);
nor U5741 (N_5741,N_2438,N_2329);
or U5742 (N_5742,N_1876,N_2699);
and U5743 (N_5743,N_88,N_1481);
nand U5744 (N_5744,N_1203,N_2269);
nor U5745 (N_5745,N_801,N_1980);
nor U5746 (N_5746,N_383,N_2876);
nand U5747 (N_5747,N_1215,N_1526);
or U5748 (N_5748,N_2820,N_2606);
or U5749 (N_5749,N_2756,N_720);
nor U5750 (N_5750,N_2719,N_2615);
nand U5751 (N_5751,N_750,N_1070);
nor U5752 (N_5752,N_1018,N_2612);
or U5753 (N_5753,N_232,N_1289);
nor U5754 (N_5754,N_2778,N_1082);
or U5755 (N_5755,N_2911,N_2592);
or U5756 (N_5756,N_1189,N_2189);
nand U5757 (N_5757,N_2560,N_1271);
and U5758 (N_5758,N_1470,N_311);
and U5759 (N_5759,N_1928,N_830);
and U5760 (N_5760,N_1854,N_1951);
and U5761 (N_5761,N_2121,N_594);
and U5762 (N_5762,N_2954,N_2450);
nand U5763 (N_5763,N_97,N_1793);
and U5764 (N_5764,N_1537,N_413);
and U5765 (N_5765,N_2763,N_2250);
and U5766 (N_5766,N_304,N_2966);
or U5767 (N_5767,N_219,N_65);
nand U5768 (N_5768,N_704,N_1001);
and U5769 (N_5769,N_57,N_2006);
and U5770 (N_5770,N_307,N_1754);
nand U5771 (N_5771,N_2067,N_849);
or U5772 (N_5772,N_1050,N_2290);
nor U5773 (N_5773,N_1858,N_1414);
nand U5774 (N_5774,N_2598,N_2549);
and U5775 (N_5775,N_2915,N_1719);
and U5776 (N_5776,N_1714,N_1158);
or U5777 (N_5777,N_2242,N_2995);
nor U5778 (N_5778,N_2452,N_1657);
and U5779 (N_5779,N_942,N_756);
nor U5780 (N_5780,N_2118,N_101);
nor U5781 (N_5781,N_554,N_2312);
nand U5782 (N_5782,N_476,N_465);
or U5783 (N_5783,N_2403,N_1279);
or U5784 (N_5784,N_577,N_2534);
nor U5785 (N_5785,N_1996,N_1154);
or U5786 (N_5786,N_2041,N_729);
nor U5787 (N_5787,N_1570,N_756);
and U5788 (N_5788,N_2831,N_556);
and U5789 (N_5789,N_189,N_2649);
and U5790 (N_5790,N_262,N_2539);
nand U5791 (N_5791,N_472,N_2496);
nor U5792 (N_5792,N_1184,N_47);
nor U5793 (N_5793,N_1418,N_309);
and U5794 (N_5794,N_1898,N_2002);
or U5795 (N_5795,N_428,N_727);
and U5796 (N_5796,N_1608,N_2995);
nand U5797 (N_5797,N_2302,N_2941);
nor U5798 (N_5798,N_2699,N_342);
nor U5799 (N_5799,N_588,N_386);
nand U5800 (N_5800,N_2077,N_1127);
or U5801 (N_5801,N_1807,N_1454);
nand U5802 (N_5802,N_461,N_1305);
nor U5803 (N_5803,N_2907,N_2932);
nor U5804 (N_5804,N_1768,N_2341);
and U5805 (N_5805,N_1761,N_2598);
and U5806 (N_5806,N_1474,N_816);
nand U5807 (N_5807,N_2516,N_2676);
or U5808 (N_5808,N_1542,N_356);
nand U5809 (N_5809,N_591,N_1722);
or U5810 (N_5810,N_2226,N_1242);
or U5811 (N_5811,N_2374,N_2181);
and U5812 (N_5812,N_1208,N_96);
nor U5813 (N_5813,N_1008,N_811);
and U5814 (N_5814,N_974,N_1092);
or U5815 (N_5815,N_1148,N_2289);
and U5816 (N_5816,N_240,N_2060);
and U5817 (N_5817,N_315,N_1087);
nand U5818 (N_5818,N_521,N_96);
and U5819 (N_5819,N_1567,N_1701);
or U5820 (N_5820,N_906,N_2630);
nor U5821 (N_5821,N_1383,N_2124);
or U5822 (N_5822,N_681,N_1176);
or U5823 (N_5823,N_548,N_2542);
nand U5824 (N_5824,N_2177,N_509);
nand U5825 (N_5825,N_1917,N_1451);
nor U5826 (N_5826,N_2803,N_2921);
or U5827 (N_5827,N_1268,N_2021);
xor U5828 (N_5828,N_1465,N_1709);
or U5829 (N_5829,N_2842,N_2895);
nor U5830 (N_5830,N_580,N_1587);
nor U5831 (N_5831,N_1498,N_1455);
nand U5832 (N_5832,N_758,N_238);
and U5833 (N_5833,N_1323,N_516);
nor U5834 (N_5834,N_1602,N_516);
nor U5835 (N_5835,N_437,N_2494);
or U5836 (N_5836,N_1923,N_2108);
nor U5837 (N_5837,N_2583,N_2997);
nand U5838 (N_5838,N_1106,N_784);
and U5839 (N_5839,N_1561,N_557);
nor U5840 (N_5840,N_2526,N_1757);
or U5841 (N_5841,N_2342,N_2995);
or U5842 (N_5842,N_1486,N_1820);
nor U5843 (N_5843,N_1319,N_2975);
nor U5844 (N_5844,N_1722,N_1231);
nand U5845 (N_5845,N_932,N_2868);
nand U5846 (N_5846,N_782,N_690);
nor U5847 (N_5847,N_420,N_2677);
or U5848 (N_5848,N_431,N_1261);
nand U5849 (N_5849,N_799,N_2534);
nor U5850 (N_5850,N_2285,N_1617);
and U5851 (N_5851,N_1281,N_2);
or U5852 (N_5852,N_1145,N_1455);
and U5853 (N_5853,N_2126,N_314);
nand U5854 (N_5854,N_1600,N_722);
nor U5855 (N_5855,N_2228,N_2747);
and U5856 (N_5856,N_348,N_829);
nor U5857 (N_5857,N_782,N_689);
nor U5858 (N_5858,N_866,N_275);
or U5859 (N_5859,N_264,N_1022);
or U5860 (N_5860,N_1400,N_630);
and U5861 (N_5861,N_1497,N_1506);
nor U5862 (N_5862,N_1278,N_1236);
or U5863 (N_5863,N_32,N_2202);
or U5864 (N_5864,N_1033,N_272);
nand U5865 (N_5865,N_2595,N_302);
or U5866 (N_5866,N_2958,N_879);
nor U5867 (N_5867,N_725,N_2489);
nor U5868 (N_5868,N_1272,N_518);
or U5869 (N_5869,N_2853,N_2069);
nor U5870 (N_5870,N_2517,N_2155);
nor U5871 (N_5871,N_2325,N_2062);
and U5872 (N_5872,N_267,N_1785);
nor U5873 (N_5873,N_1785,N_662);
nand U5874 (N_5874,N_1733,N_436);
and U5875 (N_5875,N_1115,N_1040);
and U5876 (N_5876,N_545,N_2277);
nor U5877 (N_5877,N_609,N_1411);
nand U5878 (N_5878,N_1909,N_1324);
nand U5879 (N_5879,N_240,N_1510);
nor U5880 (N_5880,N_355,N_1865);
or U5881 (N_5881,N_2525,N_1434);
and U5882 (N_5882,N_2371,N_1065);
nor U5883 (N_5883,N_339,N_1269);
or U5884 (N_5884,N_2209,N_2047);
nand U5885 (N_5885,N_1548,N_2145);
nand U5886 (N_5886,N_1994,N_124);
or U5887 (N_5887,N_2049,N_89);
nand U5888 (N_5888,N_618,N_1241);
nand U5889 (N_5889,N_1089,N_1623);
or U5890 (N_5890,N_219,N_731);
or U5891 (N_5891,N_419,N_357);
or U5892 (N_5892,N_2833,N_2303);
or U5893 (N_5893,N_1868,N_2677);
or U5894 (N_5894,N_2812,N_2684);
and U5895 (N_5895,N_1471,N_2338);
nor U5896 (N_5896,N_1808,N_2497);
and U5897 (N_5897,N_1600,N_645);
and U5898 (N_5898,N_1806,N_118);
nor U5899 (N_5899,N_2569,N_2882);
and U5900 (N_5900,N_535,N_973);
nor U5901 (N_5901,N_1317,N_2530);
nor U5902 (N_5902,N_1708,N_2881);
nor U5903 (N_5903,N_2582,N_1044);
or U5904 (N_5904,N_14,N_230);
nor U5905 (N_5905,N_2897,N_478);
nor U5906 (N_5906,N_1885,N_954);
nor U5907 (N_5907,N_2949,N_2315);
nor U5908 (N_5908,N_1635,N_1563);
and U5909 (N_5909,N_1184,N_1188);
nand U5910 (N_5910,N_2883,N_843);
nor U5911 (N_5911,N_550,N_412);
or U5912 (N_5912,N_545,N_594);
nand U5913 (N_5913,N_1813,N_1152);
nand U5914 (N_5914,N_2263,N_250);
or U5915 (N_5915,N_2452,N_1470);
nor U5916 (N_5916,N_2050,N_2102);
nor U5917 (N_5917,N_972,N_2515);
and U5918 (N_5918,N_1757,N_1055);
and U5919 (N_5919,N_2247,N_2724);
nand U5920 (N_5920,N_1239,N_2545);
nor U5921 (N_5921,N_2593,N_1083);
or U5922 (N_5922,N_2713,N_2225);
or U5923 (N_5923,N_430,N_2938);
or U5924 (N_5924,N_238,N_1184);
nand U5925 (N_5925,N_304,N_699);
nor U5926 (N_5926,N_51,N_1768);
or U5927 (N_5927,N_2890,N_699);
and U5928 (N_5928,N_2418,N_209);
nand U5929 (N_5929,N_151,N_1734);
or U5930 (N_5930,N_2555,N_1080);
nor U5931 (N_5931,N_91,N_2303);
nor U5932 (N_5932,N_2781,N_1238);
or U5933 (N_5933,N_509,N_903);
and U5934 (N_5934,N_983,N_546);
nor U5935 (N_5935,N_1333,N_2594);
nor U5936 (N_5936,N_1642,N_2644);
nand U5937 (N_5937,N_1592,N_2471);
and U5938 (N_5938,N_1089,N_555);
nand U5939 (N_5939,N_1668,N_2057);
and U5940 (N_5940,N_934,N_2980);
or U5941 (N_5941,N_793,N_1989);
nor U5942 (N_5942,N_1849,N_2151);
nand U5943 (N_5943,N_568,N_1206);
nand U5944 (N_5944,N_2528,N_2187);
or U5945 (N_5945,N_264,N_2721);
and U5946 (N_5946,N_1663,N_2449);
nand U5947 (N_5947,N_2361,N_378);
nand U5948 (N_5948,N_2592,N_2076);
nor U5949 (N_5949,N_1785,N_288);
and U5950 (N_5950,N_2030,N_2768);
and U5951 (N_5951,N_1658,N_2537);
nand U5952 (N_5952,N_2244,N_2921);
and U5953 (N_5953,N_1211,N_1216);
or U5954 (N_5954,N_1970,N_2636);
and U5955 (N_5955,N_1602,N_2954);
nand U5956 (N_5956,N_927,N_2329);
nor U5957 (N_5957,N_193,N_797);
nand U5958 (N_5958,N_2295,N_1008);
nor U5959 (N_5959,N_2401,N_1420);
or U5960 (N_5960,N_1667,N_2227);
or U5961 (N_5961,N_464,N_1204);
or U5962 (N_5962,N_25,N_498);
or U5963 (N_5963,N_129,N_636);
nand U5964 (N_5964,N_335,N_714);
or U5965 (N_5965,N_2406,N_2603);
nor U5966 (N_5966,N_1695,N_1850);
nand U5967 (N_5967,N_1315,N_272);
and U5968 (N_5968,N_2587,N_1940);
or U5969 (N_5969,N_2491,N_1082);
or U5970 (N_5970,N_1484,N_2612);
and U5971 (N_5971,N_1864,N_906);
or U5972 (N_5972,N_2209,N_2360);
or U5973 (N_5973,N_101,N_1489);
or U5974 (N_5974,N_345,N_2619);
or U5975 (N_5975,N_1245,N_267);
and U5976 (N_5976,N_2659,N_2682);
or U5977 (N_5977,N_1946,N_586);
nor U5978 (N_5978,N_753,N_47);
nor U5979 (N_5979,N_1329,N_593);
nor U5980 (N_5980,N_2607,N_193);
nor U5981 (N_5981,N_398,N_2289);
or U5982 (N_5982,N_1911,N_1044);
nor U5983 (N_5983,N_953,N_1818);
nor U5984 (N_5984,N_2255,N_32);
or U5985 (N_5985,N_544,N_2990);
nor U5986 (N_5986,N_603,N_1256);
nand U5987 (N_5987,N_2686,N_641);
nor U5988 (N_5988,N_572,N_123);
or U5989 (N_5989,N_2983,N_34);
and U5990 (N_5990,N_2963,N_978);
and U5991 (N_5991,N_1816,N_1147);
nand U5992 (N_5992,N_2705,N_2565);
xnor U5993 (N_5993,N_2471,N_744);
nand U5994 (N_5994,N_499,N_542);
nor U5995 (N_5995,N_2554,N_2261);
nor U5996 (N_5996,N_777,N_1742);
nand U5997 (N_5997,N_2139,N_2353);
nor U5998 (N_5998,N_675,N_1350);
nor U5999 (N_5999,N_387,N_421);
nor U6000 (N_6000,N_5795,N_5906);
or U6001 (N_6001,N_3744,N_3723);
nor U6002 (N_6002,N_5585,N_4856);
and U6003 (N_6003,N_5817,N_3748);
and U6004 (N_6004,N_5498,N_5901);
and U6005 (N_6005,N_3722,N_3648);
nand U6006 (N_6006,N_4809,N_3965);
or U6007 (N_6007,N_3104,N_3398);
nand U6008 (N_6008,N_4750,N_3186);
nand U6009 (N_6009,N_4067,N_3565);
and U6010 (N_6010,N_3263,N_3576);
nand U6011 (N_6011,N_5350,N_5614);
or U6012 (N_6012,N_3456,N_5996);
nand U6013 (N_6013,N_5912,N_4507);
and U6014 (N_6014,N_3006,N_3168);
and U6015 (N_6015,N_5482,N_4563);
or U6016 (N_6016,N_5290,N_4373);
nand U6017 (N_6017,N_4588,N_3608);
and U6018 (N_6018,N_5608,N_4354);
or U6019 (N_6019,N_4817,N_4480);
nand U6020 (N_6020,N_5777,N_5063);
nor U6021 (N_6021,N_3108,N_3626);
nor U6022 (N_6022,N_3789,N_4719);
and U6023 (N_6023,N_4850,N_3474);
nand U6024 (N_6024,N_4463,N_5926);
nor U6025 (N_6025,N_3176,N_5533);
and U6026 (N_6026,N_3933,N_4431);
or U6027 (N_6027,N_3316,N_5379);
or U6028 (N_6028,N_3547,N_4397);
nand U6029 (N_6029,N_3686,N_4937);
nand U6030 (N_6030,N_3348,N_3553);
nor U6031 (N_6031,N_5723,N_3486);
or U6032 (N_6032,N_4299,N_5489);
nor U6033 (N_6033,N_4611,N_5786);
nand U6034 (N_6034,N_5376,N_4529);
nand U6035 (N_6035,N_3107,N_4016);
nand U6036 (N_6036,N_3241,N_4590);
and U6037 (N_6037,N_4302,N_4743);
or U6038 (N_6038,N_4316,N_3950);
nor U6039 (N_6039,N_4601,N_3335);
and U6040 (N_6040,N_4199,N_5472);
nor U6041 (N_6041,N_3084,N_3853);
or U6042 (N_6042,N_3217,N_4591);
nand U6043 (N_6043,N_4481,N_3513);
nor U6044 (N_6044,N_3393,N_3767);
or U6045 (N_6045,N_4886,N_4244);
nand U6046 (N_6046,N_4757,N_3735);
and U6047 (N_6047,N_5479,N_4716);
or U6048 (N_6048,N_5011,N_4685);
or U6049 (N_6049,N_4806,N_3362);
nor U6050 (N_6050,N_3167,N_4721);
and U6051 (N_6051,N_5109,N_5270);
nand U6052 (N_6052,N_4863,N_4043);
or U6053 (N_6053,N_3187,N_3886);
nor U6054 (N_6054,N_5341,N_3394);
nor U6055 (N_6055,N_5949,N_3544);
nor U6056 (N_6056,N_5371,N_5712);
and U6057 (N_6057,N_3321,N_5726);
nor U6058 (N_6058,N_3026,N_4267);
nand U6059 (N_6059,N_5496,N_4028);
nor U6060 (N_6060,N_5149,N_3232);
or U6061 (N_6061,N_3034,N_3437);
nor U6062 (N_6062,N_3236,N_4147);
nor U6063 (N_6063,N_5237,N_5984);
nand U6064 (N_6064,N_4892,N_5210);
and U6065 (N_6065,N_3360,N_3438);
or U6066 (N_6066,N_3048,N_5054);
and U6067 (N_6067,N_5071,N_4361);
nor U6068 (N_6068,N_4714,N_4889);
nor U6069 (N_6069,N_5811,N_5846);
or U6070 (N_6070,N_3624,N_4428);
and U6071 (N_6071,N_5158,N_5528);
nand U6072 (N_6072,N_4207,N_4745);
nand U6073 (N_6073,N_5782,N_3039);
nor U6074 (N_6074,N_5240,N_5464);
or U6075 (N_6075,N_5890,N_5781);
and U6076 (N_6076,N_5447,N_5577);
nand U6077 (N_6077,N_5667,N_4639);
nor U6078 (N_6078,N_3949,N_3032);
or U6079 (N_6079,N_3075,N_5920);
nand U6080 (N_6080,N_4795,N_3505);
or U6081 (N_6081,N_5431,N_4787);
nand U6082 (N_6082,N_3813,N_5282);
or U6083 (N_6083,N_4180,N_3778);
or U6084 (N_6084,N_5275,N_3925);
or U6085 (N_6085,N_3552,N_3707);
nand U6086 (N_6086,N_4421,N_4926);
nor U6087 (N_6087,N_5862,N_5609);
and U6088 (N_6088,N_3826,N_4116);
nand U6089 (N_6089,N_4951,N_4363);
or U6090 (N_6090,N_4675,N_3694);
nor U6091 (N_6091,N_4625,N_4018);
or U6092 (N_6092,N_5245,N_5174);
nand U6093 (N_6093,N_4818,N_5799);
nor U6094 (N_6094,N_3257,N_4642);
nor U6095 (N_6095,N_4621,N_5132);
and U6096 (N_6096,N_5491,N_4240);
and U6097 (N_6097,N_4755,N_3643);
or U6098 (N_6098,N_4712,N_4236);
or U6099 (N_6099,N_5775,N_4358);
or U6100 (N_6100,N_5870,N_5448);
or U6101 (N_6101,N_5874,N_3568);
and U6102 (N_6102,N_3312,N_4989);
nand U6103 (N_6103,N_3504,N_3916);
and U6104 (N_6104,N_3889,N_5702);
xnor U6105 (N_6105,N_4437,N_3237);
nand U6106 (N_6106,N_3213,N_5902);
nor U6107 (N_6107,N_5087,N_5815);
nor U6108 (N_6108,N_3426,N_4350);
and U6109 (N_6109,N_3894,N_5160);
nor U6110 (N_6110,N_4532,N_3387);
and U6111 (N_6111,N_4950,N_4980);
or U6112 (N_6112,N_5114,N_5737);
and U6113 (N_6113,N_4117,N_4624);
xor U6114 (N_6114,N_5007,N_4972);
nand U6115 (N_6115,N_4545,N_4938);
nand U6116 (N_6116,N_4276,N_4749);
and U6117 (N_6117,N_3253,N_3013);
or U6118 (N_6118,N_4238,N_4053);
or U6119 (N_6119,N_4086,N_3961);
nor U6120 (N_6120,N_3753,N_4837);
nor U6121 (N_6121,N_3842,N_3841);
and U6122 (N_6122,N_5622,N_5875);
nor U6123 (N_6123,N_5192,N_5218);
and U6124 (N_6124,N_3984,N_4357);
or U6125 (N_6125,N_4660,N_5857);
or U6126 (N_6126,N_5956,N_4943);
or U6127 (N_6127,N_3855,N_5567);
or U6128 (N_6128,N_3058,N_5497);
and U6129 (N_6129,N_3132,N_3097);
and U6130 (N_6130,N_4620,N_3715);
and U6131 (N_6131,N_5717,N_5280);
or U6132 (N_6132,N_3745,N_5238);
or U6133 (N_6133,N_4371,N_4157);
nor U6134 (N_6134,N_3710,N_4499);
nor U6135 (N_6135,N_5823,N_5801);
nor U6136 (N_6136,N_3867,N_5829);
and U6137 (N_6137,N_3462,N_3849);
or U6138 (N_6138,N_5190,N_3077);
or U6139 (N_6139,N_5584,N_3687);
nor U6140 (N_6140,N_3602,N_3177);
and U6141 (N_6141,N_3935,N_5592);
nand U6142 (N_6142,N_4115,N_5826);
nor U6143 (N_6143,N_4403,N_5961);
nor U6144 (N_6144,N_3846,N_3772);
or U6145 (N_6145,N_3421,N_3963);
and U6146 (N_6146,N_3378,N_5761);
nor U6147 (N_6147,N_5661,N_3164);
nor U6148 (N_6148,N_3470,N_3671);
or U6149 (N_6149,N_3133,N_5217);
nor U6150 (N_6150,N_4544,N_5408);
nand U6151 (N_6151,N_5285,N_5928);
or U6152 (N_6152,N_4342,N_3004);
nor U6153 (N_6153,N_3999,N_3681);
or U6154 (N_6154,N_5587,N_4074);
and U6155 (N_6155,N_5014,N_5615);
or U6156 (N_6156,N_5611,N_4287);
nor U6157 (N_6157,N_5539,N_5220);
nand U6158 (N_6158,N_3952,N_4643);
nor U6159 (N_6159,N_4002,N_4145);
nor U6160 (N_6160,N_5105,N_3159);
and U6161 (N_6161,N_3319,N_3498);
nor U6162 (N_6162,N_5636,N_3756);
nor U6163 (N_6163,N_5517,N_5876);
nand U6164 (N_6164,N_5886,N_3981);
and U6165 (N_6165,N_5720,N_5982);
and U6166 (N_6166,N_4406,N_3340);
nor U6167 (N_6167,N_4435,N_5260);
nor U6168 (N_6168,N_5714,N_4670);
nand U6169 (N_6169,N_5230,N_4770);
nand U6170 (N_6170,N_3808,N_4124);
nand U6171 (N_6171,N_4022,N_5674);
and U6172 (N_6172,N_3342,N_5677);
nor U6173 (N_6173,N_5945,N_5239);
or U6174 (N_6174,N_4033,N_4232);
nor U6175 (N_6175,N_4652,N_3871);
nand U6176 (N_6176,N_3721,N_4498);
and U6177 (N_6177,N_5589,N_3765);
or U6178 (N_6178,N_5803,N_3351);
and U6179 (N_6179,N_4303,N_5368);
or U6180 (N_6180,N_5575,N_3969);
xnor U6181 (N_6181,N_4132,N_3863);
nor U6182 (N_6182,N_5625,N_3233);
or U6183 (N_6183,N_4204,N_5925);
nor U6184 (N_6184,N_3011,N_5839);
nand U6185 (N_6185,N_5568,N_4667);
nand U6186 (N_6186,N_5933,N_4317);
nor U6187 (N_6187,N_5663,N_5731);
nand U6188 (N_6188,N_4993,N_3230);
nor U6189 (N_6189,N_4726,N_4095);
nor U6190 (N_6190,N_5166,N_5018);
and U6191 (N_6191,N_4899,N_4493);
nor U6192 (N_6192,N_4253,N_3339);
nor U6193 (N_6193,N_5868,N_5969);
nand U6194 (N_6194,N_4091,N_5035);
nor U6195 (N_6195,N_5012,N_5346);
nor U6196 (N_6196,N_3771,N_5740);
nand U6197 (N_6197,N_5778,N_3429);
or U6198 (N_6198,N_4212,N_5459);
nor U6199 (N_6199,N_5798,N_5983);
or U6200 (N_6200,N_5534,N_3243);
or U6201 (N_6201,N_4554,N_4125);
or U6202 (N_6202,N_5721,N_4870);
nor U6203 (N_6203,N_5200,N_5168);
nand U6204 (N_6204,N_4995,N_4780);
nand U6205 (N_6205,N_3953,N_4008);
nor U6206 (N_6206,N_4559,N_5177);
and U6207 (N_6207,N_4045,N_5957);
nand U6208 (N_6208,N_5655,N_5435);
and U6209 (N_6209,N_5793,N_4737);
or U6210 (N_6210,N_4884,N_4882);
nand U6211 (N_6211,N_4496,N_5686);
nand U6212 (N_6212,N_4164,N_5252);
and U6213 (N_6213,N_5223,N_5896);
nand U6214 (N_6214,N_3661,N_4484);
nor U6215 (N_6215,N_3079,N_4548);
and U6216 (N_6216,N_3215,N_3884);
and U6217 (N_6217,N_5658,N_4669);
nor U6218 (N_6218,N_3258,N_5649);
nand U6219 (N_6219,N_5405,N_4665);
nor U6220 (N_6220,N_3860,N_5576);
nand U6221 (N_6221,N_5402,N_3030);
nand U6222 (N_6222,N_3008,N_5856);
nor U6223 (N_6223,N_5020,N_5488);
and U6224 (N_6224,N_5578,N_5774);
or U6225 (N_6225,N_3918,N_5049);
or U6226 (N_6226,N_3412,N_5932);
or U6227 (N_6227,N_3046,N_3928);
or U6228 (N_6228,N_3469,N_4701);
nor U6229 (N_6229,N_4869,N_3214);
and U6230 (N_6230,N_5470,N_4345);
nor U6231 (N_6231,N_4285,N_3388);
and U6232 (N_6232,N_3146,N_5347);
nor U6233 (N_6233,N_4275,N_5443);
or U6234 (N_6234,N_4891,N_3502);
and U6235 (N_6235,N_5162,N_4202);
nand U6236 (N_6236,N_3290,N_3171);
nor U6237 (N_6237,N_5530,N_4622);
or U6238 (N_6238,N_4800,N_4222);
nand U6239 (N_6239,N_4860,N_3773);
nor U6240 (N_6240,N_4509,N_3158);
and U6241 (N_6241,N_4450,N_4593);
and U6242 (N_6242,N_5469,N_5026);
and U6243 (N_6243,N_5808,N_5526);
and U6244 (N_6244,N_5255,N_4245);
nand U6245 (N_6245,N_3838,N_5022);
and U6246 (N_6246,N_5329,N_5088);
nand U6247 (N_6247,N_4468,N_3788);
and U6248 (N_6248,N_3797,N_4184);
or U6249 (N_6249,N_3955,N_4042);
and U6250 (N_6250,N_3248,N_4278);
nand U6251 (N_6251,N_4602,N_5999);
nor U6252 (N_6252,N_3210,N_4374);
nor U6253 (N_6253,N_4341,N_4930);
or U6254 (N_6254,N_3810,N_4235);
and U6255 (N_6255,N_5827,N_3044);
nor U6256 (N_6256,N_4816,N_4143);
nand U6257 (N_6257,N_5452,N_3052);
nor U6258 (N_6258,N_5084,N_5072);
or U6259 (N_6259,N_3637,N_3542);
and U6260 (N_6260,N_4713,N_5784);
nor U6261 (N_6261,N_4748,N_4650);
nand U6262 (N_6262,N_3834,N_3267);
nor U6263 (N_6263,N_4206,N_3635);
or U6264 (N_6264,N_4901,N_3571);
nor U6265 (N_6265,N_4195,N_5785);
nand U6266 (N_6266,N_4141,N_4488);
nand U6267 (N_6267,N_4252,N_3518);
and U6268 (N_6268,N_4512,N_5748);
and U6269 (N_6269,N_3559,N_3795);
and U6270 (N_6270,N_4518,N_3835);
or U6271 (N_6271,N_5085,N_5715);
nor U6272 (N_6272,N_4596,N_3774);
or U6273 (N_6273,N_3154,N_3366);
nor U6274 (N_6274,N_3997,N_5525);
nor U6275 (N_6275,N_4013,N_4183);
nor U6276 (N_6276,N_4872,N_4606);
nand U6277 (N_6277,N_4990,N_4689);
nand U6278 (N_6278,N_4348,N_5788);
or U6279 (N_6279,N_5481,N_3747);
or U6280 (N_6280,N_3049,N_5582);
or U6281 (N_6281,N_5753,N_3225);
or U6282 (N_6282,N_4017,N_3464);
nor U6283 (N_6283,N_3787,N_4858);
and U6284 (N_6284,N_5716,N_4516);
nor U6285 (N_6285,N_4107,N_3382);
nor U6286 (N_6286,N_3716,N_5633);
nor U6287 (N_6287,N_5898,N_3951);
nor U6288 (N_6288,N_3100,N_4375);
and U6289 (N_6289,N_4706,N_4440);
and U6290 (N_6290,N_5380,N_4490);
and U6291 (N_6291,N_3799,N_3990);
and U6292 (N_6292,N_5466,N_3252);
nand U6293 (N_6293,N_4328,N_4466);
nand U6294 (N_6294,N_3208,N_5449);
nor U6295 (N_6295,N_5334,N_5473);
nor U6296 (N_6296,N_4411,N_4129);
nor U6297 (N_6297,N_5410,N_5416);
and U6298 (N_6298,N_3452,N_4945);
nand U6299 (N_6299,N_4925,N_5694);
nor U6300 (N_6300,N_3289,N_3482);
nor U6301 (N_6301,N_4366,N_5978);
or U6302 (N_6302,N_4740,N_3440);
and U6303 (N_6303,N_4137,N_4283);
nand U6304 (N_6304,N_4400,N_3831);
nand U6305 (N_6305,N_5216,N_4582);
or U6306 (N_6306,N_4981,N_3384);
and U6307 (N_6307,N_3015,N_4258);
and U6308 (N_6308,N_4911,N_5994);
or U6309 (N_6309,N_4325,N_5535);
nor U6310 (N_6310,N_4900,N_3690);
and U6311 (N_6311,N_3807,N_4152);
nand U6312 (N_6312,N_3515,N_3657);
or U6313 (N_6313,N_4613,N_4955);
and U6314 (N_6314,N_3524,N_3848);
nand U6315 (N_6315,N_3455,N_5882);
nor U6316 (N_6316,N_3446,N_4326);
or U6317 (N_6317,N_4991,N_4081);
or U6318 (N_6318,N_3124,N_4176);
nand U6319 (N_6319,N_3895,N_4920);
and U6320 (N_6320,N_4021,N_4208);
nand U6321 (N_6321,N_3299,N_5976);
or U6322 (N_6322,N_4452,N_3212);
or U6323 (N_6323,N_4815,N_4163);
nand U6324 (N_6324,N_3574,N_5554);
nor U6325 (N_6325,N_3535,N_3862);
nor U6326 (N_6326,N_3956,N_5215);
nand U6327 (N_6327,N_4055,N_4982);
or U6328 (N_6328,N_3493,N_5383);
nor U6329 (N_6329,N_3960,N_5821);
or U6330 (N_6330,N_5648,N_4142);
or U6331 (N_6331,N_4395,N_5809);
or U6332 (N_6332,N_4457,N_4629);
and U6333 (N_6333,N_3979,N_3577);
nor U6334 (N_6334,N_4793,N_3078);
nor U6335 (N_6335,N_5092,N_4465);
and U6336 (N_6336,N_3536,N_5706);
or U6337 (N_6337,N_5373,N_3817);
nor U6338 (N_6338,N_5860,N_5056);
nand U6339 (N_6339,N_5779,N_3226);
nor U6340 (N_6340,N_4974,N_5900);
nor U6341 (N_6341,N_5362,N_5852);
or U6342 (N_6342,N_3254,N_4835);
nor U6343 (N_6343,N_5427,N_3231);
or U6344 (N_6344,N_4487,N_4075);
or U6345 (N_6345,N_4730,N_4715);
and U6346 (N_6346,N_4257,N_3785);
nand U6347 (N_6347,N_3709,N_3009);
or U6348 (N_6348,N_4663,N_4517);
or U6349 (N_6349,N_4690,N_4420);
nand U6350 (N_6350,N_4194,N_5915);
or U6351 (N_6351,N_5083,N_4814);
nor U6352 (N_6352,N_5231,N_5492);
nor U6353 (N_6353,N_4523,N_5244);
nor U6354 (N_6354,N_5221,N_5951);
nor U6355 (N_6355,N_4094,N_4369);
nor U6356 (N_6356,N_5283,N_5598);
nand U6357 (N_6357,N_3373,N_4648);
or U6358 (N_6358,N_3472,N_5760);
and U6359 (N_6359,N_4557,N_4359);
xor U6360 (N_6360,N_5509,N_3644);
nor U6361 (N_6361,N_4272,N_3037);
nor U6362 (N_6362,N_4140,N_3940);
nand U6363 (N_6363,N_5082,N_5000);
nor U6364 (N_6364,N_3454,N_4578);
nand U6365 (N_6365,N_4992,N_5523);
nand U6366 (N_6366,N_3076,N_3409);
and U6367 (N_6367,N_5420,N_5848);
xor U6368 (N_6368,N_5503,N_4134);
nor U6369 (N_6369,N_4378,N_5502);
and U6370 (N_6370,N_5964,N_5513);
nand U6371 (N_6371,N_4030,N_3594);
and U6372 (N_6372,N_4682,N_5058);
nand U6373 (N_6373,N_5551,N_3488);
and U6374 (N_6374,N_5391,N_3139);
and U6375 (N_6375,N_4246,N_3395);
nor U6376 (N_6376,N_5165,N_5224);
and U6377 (N_6377,N_3777,N_3972);
nor U6378 (N_6378,N_3677,N_4310);
nor U6379 (N_6379,N_5264,N_5745);
or U6380 (N_6380,N_3255,N_5594);
or U6381 (N_6381,N_3297,N_4553);
nand U6382 (N_6382,N_5953,N_5262);
nor U6383 (N_6383,N_4438,N_3062);
and U6384 (N_6384,N_4692,N_4315);
nand U6385 (N_6385,N_4751,N_5243);
and U6386 (N_6386,N_5791,N_4429);
or U6387 (N_6387,N_4187,N_4828);
nor U6388 (N_6388,N_4177,N_4402);
nand U6389 (N_6389,N_5671,N_3377);
nor U6390 (N_6390,N_5693,N_5429);
nor U6391 (N_6391,N_5261,N_4513);
nor U6392 (N_6392,N_3822,N_5424);
nand U6393 (N_6393,N_4932,N_5382);
or U6394 (N_6394,N_3095,N_5922);
xor U6395 (N_6395,N_5642,N_4447);
nand U6396 (N_6396,N_5604,N_5769);
or U6397 (N_6397,N_3560,N_4076);
and U6398 (N_6398,N_5581,N_3349);
nand U6399 (N_6399,N_5540,N_4736);
nor U6400 (N_6400,N_3134,N_4691);
and U6401 (N_6401,N_5102,N_3761);
and U6402 (N_6402,N_3223,N_4004);
and U6403 (N_6403,N_4112,N_5550);
and U6404 (N_6404,N_5757,N_4158);
nand U6405 (N_6405,N_4636,N_3156);
or U6406 (N_6406,N_4201,N_4603);
or U6407 (N_6407,N_5790,N_3216);
and U6408 (N_6408,N_5400,N_3010);
nand U6409 (N_6409,N_4464,N_5352);
and U6410 (N_6410,N_4168,N_4467);
nand U6411 (N_6411,N_3404,N_4864);
nor U6412 (N_6412,N_5374,N_4247);
nand U6413 (N_6413,N_5947,N_4502);
nor U6414 (N_6414,N_5254,N_3368);
nand U6415 (N_6415,N_3879,N_4680);
nand U6416 (N_6416,N_4600,N_3851);
or U6417 (N_6417,N_5699,N_4426);
nand U6418 (N_6418,N_3613,N_4475);
and U6419 (N_6419,N_5032,N_3196);
nor U6420 (N_6420,N_3794,N_4093);
and U6421 (N_6421,N_3408,N_3000);
nand U6422 (N_6422,N_4471,N_5954);
nor U6423 (N_6423,N_3859,N_4922);
nand U6424 (N_6424,N_4641,N_5475);
nor U6425 (N_6425,N_3054,N_5337);
nand U6426 (N_6426,N_5314,N_5330);
nor U6427 (N_6427,N_5751,N_3380);
nand U6428 (N_6428,N_5653,N_3012);
nor U6429 (N_6429,N_5421,N_4010);
nand U6430 (N_6430,N_3638,N_5486);
or U6431 (N_6431,N_4005,N_3971);
nand U6432 (N_6432,N_3750,N_5871);
and U6433 (N_6433,N_3523,N_3125);
nor U6434 (N_6434,N_3307,N_5847);
and U6435 (N_6435,N_3458,N_4581);
nor U6436 (N_6436,N_4966,N_3857);
or U6437 (N_6437,N_3682,N_5457);
and U6438 (N_6438,N_4226,N_4949);
or U6439 (N_6439,N_5806,N_4329);
and U6440 (N_6440,N_5484,N_5364);
nor U6441 (N_6441,N_5172,N_5855);
and U6442 (N_6442,N_3658,N_5718);
nand U6443 (N_6443,N_4758,N_3617);
and U6444 (N_6444,N_3966,N_5003);
and U6445 (N_6445,N_5370,N_4580);
nor U6446 (N_6446,N_4617,N_4827);
nor U6447 (N_6447,N_5746,N_3890);
or U6448 (N_6448,N_3946,N_3138);
and U6449 (N_6449,N_3419,N_4696);
nor U6450 (N_6450,N_5097,N_5041);
or U6451 (N_6451,N_4893,N_3094);
and U6452 (N_6452,N_3942,N_4027);
xnor U6453 (N_6453,N_5090,N_3934);
or U6454 (N_6454,N_3620,N_3228);
and U6455 (N_6455,N_4063,N_3092);
nor U6456 (N_6456,N_4673,N_3313);
or U6457 (N_6457,N_4847,N_3578);
or U6458 (N_6458,N_4791,N_3113);
nand U6459 (N_6459,N_4928,N_3194);
nor U6460 (N_6460,N_4967,N_5300);
nor U6461 (N_6461,N_5924,N_4254);
or U6462 (N_6462,N_5242,N_3072);
nor U6463 (N_6463,N_5415,N_3873);
nor U6464 (N_6464,N_5378,N_5394);
nand U6465 (N_6465,N_4106,N_4947);
nand U6466 (N_6466,N_4768,N_5134);
or U6467 (N_6467,N_5197,N_3271);
and U6468 (N_6468,N_3431,N_3291);
and U6469 (N_6469,N_3910,N_4969);
or U6470 (N_6470,N_5294,N_3222);
nand U6471 (N_6471,N_4890,N_4156);
nor U6472 (N_6472,N_4085,N_5468);
nor U6473 (N_6473,N_5770,N_3318);
or U6474 (N_6474,N_3840,N_5112);
and U6475 (N_6475,N_3800,N_5814);
and U6476 (N_6476,N_5738,N_5837);
or U6477 (N_6477,N_5311,N_4078);
nand U6478 (N_6478,N_5091,N_5247);
xor U6479 (N_6479,N_4698,N_3606);
or U6480 (N_6480,N_5646,N_4666);
nor U6481 (N_6481,N_3927,N_5086);
and U6482 (N_6482,N_4702,N_3902);
or U6483 (N_6483,N_5796,N_5529);
and U6484 (N_6484,N_5708,N_3325);
or U6485 (N_6485,N_3737,N_5810);
nor U6486 (N_6486,N_3468,N_5624);
nor U6487 (N_6487,N_4668,N_4126);
nor U6488 (N_6488,N_4561,N_4656);
nor U6489 (N_6489,N_3533,N_4771);
or U6490 (N_6490,N_4623,N_4089);
or U6491 (N_6491,N_4057,N_5545);
nor U6492 (N_6492,N_3850,N_5600);
nor U6493 (N_6493,N_5516,N_4574);
nand U6494 (N_6494,N_5253,N_4775);
nor U6495 (N_6495,N_4555,N_3896);
nor U6496 (N_6496,N_3926,N_4229);
nand U6497 (N_6497,N_3150,N_3988);
nand U6498 (N_6498,N_4006,N_4594);
or U6499 (N_6499,N_5357,N_5617);
nand U6500 (N_6500,N_5683,N_5246);
nand U6501 (N_6501,N_3945,N_5025);
or U6502 (N_6502,N_3603,N_3982);
nor U6503 (N_6503,N_3604,N_5336);
or U6504 (N_6504,N_4300,N_3181);
nand U6505 (N_6505,N_5580,N_5015);
or U6506 (N_6506,N_3203,N_4760);
nand U6507 (N_6507,N_5755,N_3369);
or U6508 (N_6508,N_5818,N_5844);
and U6509 (N_6509,N_5107,N_3182);
nand U6510 (N_6510,N_5507,N_3310);
and U6511 (N_6511,N_5752,N_4489);
nand U6512 (N_6512,N_3425,N_4710);
nor U6513 (N_6513,N_4695,N_3976);
nand U6514 (N_6514,N_3475,N_4798);
nand U6515 (N_6515,N_3106,N_4384);
and U6516 (N_6516,N_5916,N_5910);
nor U6517 (N_6517,N_5395,N_4764);
nor U6518 (N_6518,N_3740,N_5004);
nand U6519 (N_6519,N_5414,N_3135);
and U6520 (N_6520,N_4248,N_5866);
or U6521 (N_6521,N_5017,N_4694);
and U6522 (N_6522,N_5317,N_4224);
and U6523 (N_6523,N_3112,N_4821);
and U6524 (N_6524,N_4776,N_4878);
nand U6525 (N_6525,N_3580,N_3487);
nand U6526 (N_6526,N_3047,N_5560);
nor U6527 (N_6527,N_3645,N_3344);
or U6528 (N_6528,N_3557,N_4699);
nand U6529 (N_6529,N_3759,N_4994);
xnor U6530 (N_6530,N_3123,N_4973);
or U6531 (N_6531,N_3651,N_4918);
nand U6532 (N_6532,N_3017,N_5859);
nor U6533 (N_6533,N_3676,N_4451);
nand U6534 (N_6534,N_4802,N_4136);
nand U6535 (N_6535,N_3760,N_3973);
and U6536 (N_6536,N_3165,N_5040);
or U6537 (N_6537,N_5583,N_4414);
and U6538 (N_6538,N_3987,N_5064);
nand U6539 (N_6539,N_3068,N_5967);
nand U6540 (N_6540,N_5772,N_3038);
nor U6541 (N_6541,N_5519,N_3619);
nor U6542 (N_6542,N_5601,N_4873);
nand U6543 (N_6543,N_3207,N_5226);
or U6544 (N_6544,N_3962,N_5023);
and U6545 (N_6545,N_3101,N_3828);
or U6546 (N_6546,N_5764,N_3292);
nor U6547 (N_6547,N_3764,N_3714);
and U6548 (N_6548,N_3306,N_5180);
nor U6549 (N_6549,N_5236,N_3596);
nand U6550 (N_6550,N_3691,N_4346);
or U6551 (N_6551,N_4933,N_4340);
or U6552 (N_6552,N_5403,N_5749);
nand U6553 (N_6553,N_3711,N_4627);
nor U6554 (N_6554,N_4923,N_3457);
nand U6555 (N_6555,N_3647,N_3669);
or U6556 (N_6556,N_3051,N_3330);
nand U6557 (N_6557,N_5101,N_3983);
and U6558 (N_6558,N_3649,N_5315);
or U6559 (N_6559,N_4778,N_5309);
and U6560 (N_6560,N_4836,N_5044);
or U6561 (N_6561,N_4659,N_5303);
nor U6562 (N_6562,N_3566,N_3116);
nor U6563 (N_6563,N_4413,N_4999);
nand U6564 (N_6564,N_3027,N_4306);
nor U6565 (N_6565,N_3202,N_4753);
nand U6566 (N_6566,N_3998,N_3405);
nand U6567 (N_6567,N_4854,N_3259);
xor U6568 (N_6568,N_5418,N_4959);
and U6569 (N_6569,N_5623,N_4568);
nor U6570 (N_6570,N_4182,N_5842);
and U6571 (N_6571,N_5854,N_3358);
and U6572 (N_6572,N_3121,N_3147);
or U6573 (N_6573,N_3195,N_4839);
or U6574 (N_6574,N_4330,N_5590);
or U6575 (N_6575,N_4961,N_4508);
nand U6576 (N_6576,N_5835,N_3695);
or U6577 (N_6577,N_5335,N_5019);
xnor U6578 (N_6578,N_3256,N_3205);
or U6579 (N_6579,N_4876,N_5096);
or U6580 (N_6580,N_3720,N_3876);
nor U6581 (N_6581,N_5679,N_3250);
or U6582 (N_6582,N_4233,N_4963);
nor U6583 (N_6583,N_5390,N_5505);
or U6584 (N_6584,N_4472,N_3583);
and U6585 (N_6585,N_5323,N_3726);
and U6586 (N_6586,N_3684,N_5207);
nand U6587 (N_6587,N_4853,N_3569);
and U6588 (N_6588,N_4040,N_4479);
or U6589 (N_6589,N_4934,N_4409);
nor U6590 (N_6590,N_5353,N_5662);
nand U6591 (N_6591,N_4765,N_4219);
nand U6592 (N_6592,N_5425,N_3821);
nand U6593 (N_6593,N_4410,N_5256);
nor U6594 (N_6594,N_4797,N_3743);
and U6595 (N_6595,N_3907,N_4801);
nand U6596 (N_6596,N_5666,N_3120);
or U6597 (N_6597,N_4250,N_3572);
nor U6598 (N_6598,N_3598,N_3540);
nor U6599 (N_6599,N_4511,N_3184);
nand U6600 (N_6600,N_5989,N_4756);
and U6601 (N_6601,N_4014,N_4610);
nand U6602 (N_6602,N_4392,N_3439);
or U6603 (N_6603,N_5241,N_3467);
nor U6604 (N_6604,N_4144,N_4108);
or U6605 (N_6605,N_3609,N_5709);
and U6606 (N_6606,N_3162,N_5965);
or U6607 (N_6607,N_3149,N_5794);
nor U6608 (N_6608,N_5897,N_3266);
nor U6609 (N_6609,N_3126,N_4181);
or U6610 (N_6610,N_3801,N_4062);
or U6611 (N_6611,N_5036,N_4486);
nor U6612 (N_6612,N_4658,N_3623);
or U6613 (N_6613,N_4333,N_5150);
and U6614 (N_6614,N_4564,N_4054);
and U6615 (N_6615,N_4349,N_5657);
or U6616 (N_6616,N_4209,N_4294);
and U6617 (N_6617,N_5068,N_3844);
nor U6618 (N_6618,N_3242,N_5828);
nor U6619 (N_6619,N_5127,N_5327);
nand U6620 (N_6620,N_4987,N_5816);
nor U6621 (N_6621,N_4996,N_3970);
nand U6622 (N_6622,N_3734,N_5997);
and U6623 (N_6623,N_5387,N_5125);
nand U6624 (N_6624,N_4412,N_5650);
and U6625 (N_6625,N_4543,N_5504);
nand U6626 (N_6626,N_5621,N_4709);
nor U6627 (N_6627,N_4521,N_5428);
nand U6628 (N_6628,N_4880,N_5389);
and U6629 (N_6629,N_3911,N_3875);
or U6630 (N_6630,N_5973,N_4065);
nor U6631 (N_6631,N_3527,N_4200);
nand U6632 (N_6632,N_4441,N_5266);
or U6633 (N_6633,N_3667,N_5461);
nand U6634 (N_6634,N_3031,N_4038);
and U6635 (N_6635,N_5038,N_3520);
nand U6636 (N_6636,N_4874,N_5603);
nand U6637 (N_6637,N_5152,N_5183);
and U6638 (N_6638,N_3442,N_3153);
nand U6639 (N_6639,N_3868,N_5100);
and U6640 (N_6640,N_4225,N_3433);
nor U6641 (N_6641,N_3538,N_3727);
and U6642 (N_6642,N_3061,N_3353);
or U6643 (N_6643,N_4483,N_5628);
nand U6644 (N_6644,N_3087,N_3296);
and U6645 (N_6645,N_4677,N_5184);
nand U6646 (N_6646,N_3328,N_3696);
or U6647 (N_6647,N_3444,N_5463);
and U6648 (N_6648,N_4540,N_5538);
or U6649 (N_6649,N_3803,N_3836);
nand U6650 (N_6650,N_3085,N_5211);
nand U6651 (N_6651,N_3646,N_4968);
and U6652 (N_6652,N_4717,N_5372);
nor U6653 (N_6653,N_4295,N_5208);
nand U6654 (N_6654,N_5295,N_5313);
or U6655 (N_6655,N_5832,N_5135);
or U6656 (N_6656,N_3268,N_3589);
or U6657 (N_6657,N_3561,N_5681);
or U6658 (N_6658,N_3705,N_3346);
nand U6659 (N_6659,N_4192,N_3118);
and U6660 (N_6660,N_5542,N_3303);
and U6661 (N_6661,N_3443,N_5700);
and U6662 (N_6662,N_4971,N_5074);
and U6663 (N_6663,N_3347,N_3595);
and U6664 (N_6664,N_4855,N_4178);
nand U6665 (N_6665,N_4867,N_3627);
and U6666 (N_6666,N_3675,N_3664);
nor U6667 (N_6667,N_3854,N_5771);
nand U6668 (N_6668,N_4166,N_3521);
and U6669 (N_6669,N_5863,N_5830);
and U6670 (N_6670,N_5122,N_4784);
and U6671 (N_6671,N_4179,N_3930);
nand U6672 (N_6672,N_3270,N_5154);
or U6673 (N_6673,N_4585,N_5462);
or U6674 (N_6674,N_3418,N_5729);
nor U6675 (N_6675,N_5432,N_4804);
or U6676 (N_6676,N_4820,N_5506);
or U6677 (N_6677,N_3337,N_4227);
nand U6678 (N_6678,N_4887,N_3142);
and U6679 (N_6679,N_4957,N_4597);
nor U6680 (N_6680,N_4482,N_3516);
and U6681 (N_6681,N_5203,N_4007);
and U6682 (N_6682,N_5892,N_4851);
and U6683 (N_6683,N_4866,N_3179);
xnor U6684 (N_6684,N_5952,N_5413);
nor U6685 (N_6685,N_3731,N_5985);
nor U6686 (N_6686,N_4048,N_4927);
nor U6687 (N_6687,N_5942,N_4576);
nor U6688 (N_6688,N_5865,N_5053);
nand U6689 (N_6689,N_4777,N_3370);
and U6690 (N_6690,N_4915,N_3461);
nand U6691 (N_6691,N_4034,N_4595);
and U6692 (N_6692,N_3057,N_5687);
nand U6693 (N_6693,N_5307,N_4845);
nand U6694 (N_6694,N_4370,N_3385);
nand U6695 (N_6695,N_5296,N_3338);
and U6696 (N_6696,N_4683,N_3003);
or U6697 (N_6697,N_5094,N_5170);
and U6698 (N_6698,N_5804,N_4237);
or U6699 (N_6699,N_3436,N_5128);
or U6700 (N_6700,N_5146,N_5055);
nand U6701 (N_6701,N_5116,N_4343);
or U6702 (N_6702,N_3417,N_4243);
nand U6703 (N_6703,N_4738,N_5393);
and U6704 (N_6704,N_3847,N_5607);
nand U6705 (N_6705,N_5284,N_4842);
and U6706 (N_6706,N_3447,N_4687);
nor U6707 (N_6707,N_4912,N_5016);
nand U6708 (N_6708,N_5783,N_4314);
nor U6709 (N_6709,N_4427,N_4807);
or U6710 (N_6710,N_4088,N_3898);
and U6711 (N_6711,N_5297,N_3173);
nand U6712 (N_6712,N_3775,N_4919);
nand U6713 (N_6713,N_5986,N_4504);
or U6714 (N_6714,N_5792,N_5634);
nand U6715 (N_6715,N_5549,N_5175);
and U6716 (N_6716,N_5196,N_5045);
or U6717 (N_6717,N_4139,N_3415);
or U6718 (N_6718,N_4386,N_3453);
and U6719 (N_6719,N_5312,N_5747);
or U6720 (N_6720,N_5703,N_3539);
and U6721 (N_6721,N_3301,N_5291);
nor U6722 (N_6722,N_3279,N_4979);
nand U6723 (N_6723,N_5487,N_3110);
and U6724 (N_6724,N_5917,N_4584);
nand U6725 (N_6725,N_3309,N_4998);
and U6726 (N_6726,N_3776,N_3152);
and U6727 (N_6727,N_3416,N_4256);
nor U6728 (N_6728,N_4097,N_3315);
and U6729 (N_6729,N_5873,N_5093);
nor U6730 (N_6730,N_5490,N_5198);
nor U6731 (N_6731,N_5618,N_3490);
nand U6732 (N_6732,N_5209,N_4883);
xor U6733 (N_6733,N_3506,N_4041);
xor U6734 (N_6734,N_3631,N_5722);
and U6735 (N_6735,N_3280,N_5298);
or U6736 (N_6736,N_3151,N_3674);
nor U6737 (N_6737,N_4565,N_3365);
and U6738 (N_6738,N_3234,N_4644);
nand U6739 (N_6739,N_3276,N_4001);
or U6740 (N_6740,N_4259,N_5050);
nor U6741 (N_6741,N_3702,N_4822);
or U6742 (N_6742,N_3912,N_4834);
nand U6743 (N_6743,N_3712,N_3996);
nand U6744 (N_6744,N_5822,N_5501);
nand U6745 (N_6745,N_4515,N_4154);
nand U6746 (N_6746,N_3700,N_3169);
or U6747 (N_6747,N_5652,N_5117);
nor U6748 (N_6748,N_3680,N_4609);
nor U6749 (N_6749,N_3249,N_5073);
nor U6750 (N_6750,N_4153,N_3074);
nor U6751 (N_6751,N_5186,N_4734);
or U6752 (N_6752,N_4841,N_3913);
and U6753 (N_6753,N_4895,N_3102);
nand U6754 (N_6754,N_5909,N_3209);
nand U6755 (N_6755,N_5735,N_4657);
or U6756 (N_6756,N_3837,N_5914);
nand U6757 (N_6757,N_5939,N_5845);
nor U6758 (N_6758,N_3128,N_4510);
and U6759 (N_6759,N_5111,N_5365);
and U6760 (N_6760,N_4684,N_5684);
nor U6761 (N_6761,N_5310,N_5493);
or U6762 (N_6762,N_4266,N_4339);
nand U6763 (N_6763,N_3809,N_4731);
nor U6764 (N_6764,N_4324,N_4525);
nor U6765 (N_6765,N_3188,N_5610);
and U6766 (N_6766,N_4264,N_5696);
nor U6767 (N_6767,N_3567,N_3549);
xor U6768 (N_6768,N_4478,N_3494);
or U6769 (N_6769,N_3944,N_5713);
nor U6770 (N_6770,N_5320,N_3080);
and U6771 (N_6771,N_4304,N_3086);
xnor U6772 (N_6772,N_3802,N_5267);
nand U6773 (N_6773,N_5557,N_5682);
nor U6774 (N_6774,N_3144,N_5227);
and U6775 (N_6775,N_3632,N_3820);
and U6776 (N_6776,N_4262,N_5750);
nor U6777 (N_6777,N_4211,N_4448);
and U6778 (N_6778,N_5477,N_3227);
and U6779 (N_6779,N_4607,N_3141);
or U6780 (N_6780,N_4046,N_3478);
and U6781 (N_6781,N_4551,N_5437);
nor U6782 (N_6782,N_3220,N_5358);
nand U6783 (N_6783,N_3939,N_3678);
or U6784 (N_6784,N_5511,N_4197);
and U6785 (N_6785,N_3304,N_4728);
nand U6786 (N_6786,N_4338,N_4746);
nand U6787 (N_6787,N_5744,N_5654);
and U6788 (N_6788,N_4382,N_4619);
and U6789 (N_6789,N_4297,N_5759);
nand U6790 (N_6790,N_4879,N_3670);
and U6791 (N_6791,N_3109,N_4032);
nand U6792 (N_6792,N_5272,N_5273);
nor U6793 (N_6793,N_3389,N_5911);
nor U6794 (N_6794,N_3450,N_3466);
and U6795 (N_6795,N_5458,N_5339);
nor U6796 (N_6796,N_5991,N_5946);
nand U6797 (N_6797,N_5189,N_4355);
nand U6798 (N_6798,N_5042,N_3754);
and U6799 (N_6799,N_5222,N_5292);
and U6800 (N_6800,N_5668,N_4781);
or U6801 (N_6801,N_5375,N_3947);
nor U6802 (N_6802,N_3798,N_4009);
or U6803 (N_6803,N_5248,N_3622);
and U6804 (N_6804,N_5979,N_3978);
or U6805 (N_6805,N_5021,N_5066);
and U6806 (N_6806,N_5558,N_5727);
nand U6807 (N_6807,N_3065,N_5235);
and U6808 (N_6808,N_4251,N_3096);
or U6809 (N_6809,N_3193,N_5299);
nand U6810 (N_6810,N_5454,N_5841);
nand U6811 (N_6811,N_4024,N_4105);
nor U6812 (N_6812,N_3751,N_4724);
nor U6813 (N_6813,N_3201,N_3974);
nand U6814 (N_6814,N_5331,N_4575);
and U6815 (N_6815,N_5034,N_3780);
or U6816 (N_6816,N_5635,N_3558);
and U6817 (N_6817,N_5510,N_4073);
nand U6818 (N_6818,N_3053,N_4196);
or U6819 (N_6819,N_3285,N_4436);
or U6820 (N_6820,N_3035,N_5411);
and U6821 (N_6821,N_3239,N_5301);
nor U6822 (N_6822,N_5213,N_4492);
nand U6823 (N_6823,N_3359,N_3041);
nand U6824 (N_6824,N_3273,N_4174);
or U6825 (N_6825,N_3564,N_3229);
nor U6826 (N_6826,N_5319,N_5591);
nor U6827 (N_6827,N_5031,N_5069);
nor U6828 (N_6828,N_5923,N_4390);
nor U6829 (N_6829,N_5548,N_5690);
and U6830 (N_6830,N_4394,N_3356);
nor U6831 (N_6831,N_4353,N_4231);
or U6832 (N_6832,N_3345,N_4894);
nor U6833 (N_6833,N_4960,N_3445);
nor U6834 (N_6834,N_5179,N_4172);
nor U6835 (N_6835,N_4221,N_3355);
nor U6836 (N_6836,N_5104,N_3878);
or U6837 (N_6837,N_5234,N_3763);
nor U6838 (N_6838,N_4096,N_5518);
nand U6839 (N_6839,N_3397,N_3379);
or U6840 (N_6840,N_3891,N_5404);
or U6841 (N_6841,N_4069,N_5768);
xor U6842 (N_6842,N_3305,N_5872);
nand U6843 (N_6843,N_4917,N_5439);
or U6844 (N_6844,N_5173,N_5360);
nor U6845 (N_6845,N_4123,N_3762);
and U6846 (N_6846,N_5569,N_3070);
nand U6847 (N_6847,N_3324,N_3314);
and U6848 (N_6848,N_4070,N_3964);
nor U6849 (N_6849,N_4598,N_3874);
or U6850 (N_6850,N_3204,N_5889);
or U6851 (N_6851,N_3901,N_4941);
or U6852 (N_6852,N_5195,N_3931);
or U6853 (N_6853,N_5471,N_3697);
nand U6854 (N_6854,N_3614,N_4445);
nor U6855 (N_6855,N_5995,N_3423);
or U6856 (N_6856,N_5521,N_3489);
nand U6857 (N_6857,N_3779,N_4026);
and U6858 (N_6858,N_4442,N_5825);
or U6859 (N_6859,N_3640,N_3655);
and U6860 (N_6860,N_4171,N_4351);
nor U6861 (N_6861,N_5397,N_3600);
nand U6862 (N_6862,N_3332,N_4039);
and U6863 (N_6863,N_3050,N_5763);
or U6864 (N_6864,N_5233,N_5321);
or U6865 (N_6865,N_5877,N_5955);
xor U6866 (N_6866,N_5159,N_3654);
nand U6867 (N_6867,N_5271,N_4773);
and U6868 (N_6868,N_4399,N_3190);
nand U6869 (N_6869,N_5377,N_3792);
nand U6870 (N_6870,N_4742,N_5919);
nand U6871 (N_6871,N_5316,N_5325);
nand U6872 (N_6872,N_5126,N_3766);
and U6873 (N_6873,N_4470,N_4396);
and U6874 (N_6874,N_4799,N_4111);
nor U6875 (N_6875,N_5787,N_3793);
and U6876 (N_6876,N_4430,N_4092);
nand U6877 (N_6877,N_5451,N_4100);
nand U6878 (N_6878,N_5199,N_5990);
nand U6879 (N_6879,N_3390,N_4906);
nand U6880 (N_6880,N_4012,N_5941);
nand U6881 (N_6881,N_5051,N_5453);
or U6882 (N_6882,N_3904,N_3829);
nor U6883 (N_6883,N_4970,N_3510);
nor U6884 (N_6884,N_5563,N_4634);
and U6885 (N_6885,N_5802,N_3191);
nand U6886 (N_6886,N_5520,N_4120);
nor U6887 (N_6887,N_4331,N_4458);
nor U6888 (N_6888,N_4454,N_4948);
nor U6889 (N_6889,N_5711,N_3752);
and U6890 (N_6890,N_4567,N_3260);
nand U6891 (N_6891,N_4615,N_4676);
and U6892 (N_6892,N_3556,N_3414);
nor U6893 (N_6893,N_4954,N_3601);
or U6894 (N_6894,N_4646,N_5143);
nor U6895 (N_6895,N_4049,N_4398);
nor U6896 (N_6896,N_4569,N_5355);
and U6897 (N_6897,N_5514,N_5742);
nand U6898 (N_6898,N_3591,N_3530);
and U6899 (N_6899,N_5422,N_3200);
or U6900 (N_6900,N_4189,N_3742);
and U6901 (N_6901,N_3511,N_4560);
and U6902 (N_6902,N_3845,N_4772);
nor U6903 (N_6903,N_4577,N_3736);
nor U6904 (N_6904,N_5369,N_3548);
or U6905 (N_6905,N_4635,N_4352);
nor U6906 (N_6906,N_4064,N_4347);
or U6907 (N_6907,N_3924,N_5602);
nor U6908 (N_6908,N_3679,N_3579);
and U6909 (N_6909,N_4035,N_5620);
nor U6910 (N_6910,N_5640,N_3781);
or U6911 (N_6911,N_3514,N_3713);
nor U6912 (N_6912,N_3391,N_3546);
nor U6913 (N_6913,N_3430,N_3371);
xor U6914 (N_6914,N_4763,N_4503);
nand U6915 (N_6915,N_4662,N_4628);
nor U6916 (N_6916,N_3016,N_4290);
nor U6917 (N_6917,N_4379,N_5899);
and U6918 (N_6918,N_3865,N_5263);
or U6919 (N_6919,N_5258,N_4727);
nor U6920 (N_6920,N_4832,N_3206);
nor U6921 (N_6921,N_5185,N_3495);
nor U6922 (N_6922,N_3732,N_5543);
or U6923 (N_6923,N_5851,N_5412);
nand U6924 (N_6924,N_3435,N_4146);
xnor U6925 (N_6925,N_5571,N_3352);
or U6926 (N_6926,N_4418,N_4313);
or U6927 (N_6927,N_3020,N_5278);
nor U6928 (N_6928,N_5758,N_4587);
or U6929 (N_6929,N_4681,N_4997);
and U6930 (N_6930,N_4277,N_4831);
xor U6931 (N_6931,N_3018,N_5903);
and U6932 (N_6932,N_3512,N_4808);
nand U6933 (N_6933,N_3336,N_3861);
and U6934 (N_6934,N_3899,N_4896);
or U6935 (N_6935,N_5766,N_5188);
or U6936 (N_6936,N_3432,N_4273);
and U6937 (N_6937,N_3381,N_4630);
nand U6938 (N_6938,N_3915,N_4813);
and U6939 (N_6939,N_4985,N_3738);
nand U6940 (N_6940,N_4288,N_3967);
and U6941 (N_6941,N_3791,N_4099);
and U6942 (N_6942,N_4579,N_4762);
and U6943 (N_6943,N_5354,N_5547);
nor U6944 (N_6944,N_5118,N_5884);
nand U6945 (N_6945,N_3718,N_4372);
nand U6946 (N_6946,N_3954,N_4393);
nor U6947 (N_6947,N_3919,N_4083);
and U6948 (N_6948,N_4223,N_5065);
and U6949 (N_6949,N_4618,N_5356);
nor U6950 (N_6950,N_5115,N_5958);
or U6951 (N_6951,N_5921,N_3022);
and U6952 (N_6952,N_4520,N_5524);
nor U6953 (N_6953,N_3042,N_5833);
nand U6954 (N_6954,N_3501,N_4434);
and U6955 (N_6955,N_5287,N_3334);
and U6956 (N_6956,N_4902,N_3685);
nor U6957 (N_6957,N_3588,N_3326);
and U6958 (N_6958,N_4519,N_5559);
nand U6959 (N_6959,N_5975,N_4589);
and U6960 (N_6960,N_5008,N_3823);
nand U6961 (N_6961,N_4811,N_3991);
xor U6962 (N_6962,N_4327,N_3562);
nand U6963 (N_6963,N_4538,N_3730);
nor U6964 (N_6964,N_3093,N_4029);
or U6965 (N_6965,N_5800,N_5689);
nor U6966 (N_6966,N_5137,N_3114);
nor U6967 (N_6967,N_3806,N_3517);
nand U6968 (N_6968,N_3363,N_5417);
nand U6969 (N_6969,N_5813,N_3693);
or U6970 (N_6970,N_4052,N_4360);
nor U6971 (N_6971,N_5660,N_3819);
and U6972 (N_6972,N_5324,N_4401);
nor U6973 (N_6973,N_4051,N_4066);
nand U6974 (N_6974,N_3434,N_4356);
or U6975 (N_6975,N_3033,N_5030);
nor U6976 (N_6976,N_5384,N_4826);
nor U6977 (N_6977,N_4131,N_4186);
or U6978 (N_6978,N_5037,N_3872);
nor U6979 (N_6979,N_5943,N_4861);
nor U6980 (N_6980,N_5555,N_5695);
nand U6981 (N_6981,N_4364,N_5359);
nand U6982 (N_6982,N_5478,N_4311);
or U6983 (N_6983,N_4819,N_3375);
and U6984 (N_6984,N_5572,N_4058);
or U6985 (N_6985,N_3247,N_4782);
xor U6986 (N_6986,N_5441,N_5776);
or U6987 (N_6987,N_4417,N_3465);
or U6988 (N_6988,N_5156,N_5419);
and U6989 (N_6989,N_3900,N_3218);
and U6990 (N_6990,N_3367,N_4640);
or U6991 (N_6991,N_5322,N_3839);
nor U6992 (N_6992,N_5269,N_3877);
nor U6993 (N_6993,N_4103,N_4110);
nor U6994 (N_6994,N_4151,N_3350);
nand U6995 (N_6995,N_5887,N_4261);
or U6996 (N_6996,N_4647,N_3909);
nand U6997 (N_6997,N_4485,N_3719);
or U6998 (N_6998,N_5274,N_5512);
nand U6999 (N_6999,N_3587,N_4649);
nor U7000 (N_7000,N_4514,N_5206);
and U7001 (N_7001,N_3060,N_4293);
or U7002 (N_7002,N_3025,N_4976);
nand U7003 (N_7003,N_5992,N_4794);
nand U7004 (N_7004,N_3628,N_5333);
and U7005 (N_7005,N_4783,N_5632);
nand U7006 (N_7006,N_3399,N_5386);
nor U7007 (N_7007,N_5138,N_4986);
and U7008 (N_7008,N_3522,N_4217);
and U7009 (N_7009,N_5052,N_4305);
nor U7010 (N_7010,N_4693,N_3914);
and U7011 (N_7011,N_4905,N_4079);
nor U7012 (N_7012,N_5931,N_5698);
or U7013 (N_7013,N_4859,N_4852);
nand U7014 (N_7014,N_4788,N_4505);
nor U7015 (N_7015,N_3610,N_3311);
or U7016 (N_7016,N_5219,N_5225);
or U7017 (N_7017,N_3534,N_3269);
and U7018 (N_7018,N_5039,N_3029);
nand U7019 (N_7019,N_5697,N_4903);
nand U7020 (N_7020,N_3881,N_3480);
nor U7021 (N_7021,N_4671,N_5710);
or U7022 (N_7022,N_5728,N_5893);
and U7023 (N_7023,N_4368,N_4334);
or U7024 (N_7024,N_4249,N_5161);
nand U7025 (N_7025,N_3975,N_5789);
nand U7026 (N_7026,N_4558,N_3758);
nor U7027 (N_7027,N_5201,N_3653);
and U7028 (N_7028,N_5527,N_3288);
nor U7029 (N_7029,N_3917,N_5927);
nor U7030 (N_7030,N_3717,N_3361);
nor U7031 (N_7031,N_4138,N_3485);
nand U7032 (N_7032,N_4205,N_5907);
nor U7033 (N_7033,N_5145,N_4688);
and U7034 (N_7034,N_4215,N_5259);
and U7035 (N_7035,N_5361,N_5605);
or U7036 (N_7036,N_4723,N_4830);
or U7037 (N_7037,N_5250,N_3261);
nor U7038 (N_7038,N_4881,N_3545);
or U7039 (N_7039,N_4704,N_5880);
or U7040 (N_7040,N_3441,N_5665);
nand U7041 (N_7041,N_4664,N_5878);
nor U7042 (N_7042,N_5399,N_4432);
and U7043 (N_7043,N_3725,N_3724);
nor U7044 (N_7044,N_5881,N_3570);
nor U7045 (N_7045,N_3551,N_3175);
and U7046 (N_7046,N_4633,N_5741);
nand U7047 (N_7047,N_5599,N_5306);
nand U7048 (N_7048,N_3883,N_5345);
nand U7049 (N_7049,N_4023,N_4733);
or U7050 (N_7050,N_4015,N_3383);
nor U7051 (N_7051,N_5398,N_4605);
nor U7052 (N_7052,N_4119,N_3043);
nor U7053 (N_7053,N_5627,N_4050);
and U7054 (N_7054,N_4255,N_4234);
nand U7055 (N_7055,N_3959,N_3088);
and U7056 (N_7056,N_4708,N_3985);
and U7057 (N_7057,N_4188,N_3659);
nand U7058 (N_7058,N_5205,N_4460);
and U7059 (N_7059,N_3235,N_4495);
nand U7060 (N_7060,N_3199,N_3612);
nand U7061 (N_7061,N_4265,N_5651);
or U7062 (N_7062,N_5739,N_3908);
or U7063 (N_7063,N_3563,N_3786);
nand U7064 (N_7064,N_5819,N_4082);
or U7065 (N_7065,N_4857,N_3341);
or U7066 (N_7066,N_5688,N_3059);
nand U7067 (N_7067,N_5998,N_3322);
and U7068 (N_7068,N_3770,N_5456);
nand U7069 (N_7069,N_4122,N_4292);
and U7070 (N_7070,N_3286,N_5656);
nor U7071 (N_7071,N_3019,N_3157);
or U7072 (N_7072,N_5009,N_3636);
and U7073 (N_7073,N_5780,N_4964);
and U7074 (N_7074,N_3211,N_3262);
nor U7075 (N_7075,N_4810,N_3427);
or U7076 (N_7076,N_3790,N_3056);
nand U7077 (N_7077,N_5467,N_5977);
and U7078 (N_7078,N_3172,N_5106);
and U7079 (N_7079,N_4844,N_3221);
nor U7080 (N_7080,N_4829,N_4722);
or U7081 (N_7081,N_5597,N_5136);
or U7082 (N_7082,N_4838,N_5385);
or U7083 (N_7083,N_4846,N_3663);
nand U7084 (N_7084,N_3308,N_4104);
nand U7085 (N_7085,N_5980,N_5057);
xor U7086 (N_7086,N_5754,N_4921);
or U7087 (N_7087,N_4868,N_4534);
and U7088 (N_7088,N_4239,N_3597);
and U7089 (N_7089,N_4672,N_3980);
nand U7090 (N_7090,N_3634,N_3994);
nor U7091 (N_7091,N_3923,N_3449);
or U7092 (N_7092,N_3396,N_4645);
nor U7093 (N_7093,N_5332,N_5685);
nor U7094 (N_7094,N_4220,N_3708);
nor U7095 (N_7095,N_4216,N_5349);
and U7096 (N_7096,N_5445,N_4935);
or U7097 (N_7097,N_5913,N_5048);
and U7098 (N_7098,N_4573,N_3298);
or U7099 (N_7099,N_3986,N_5010);
nor U7100 (N_7100,N_3130,N_3411);
nand U7101 (N_7101,N_3673,N_3818);
or U7102 (N_7102,N_3001,N_3701);
and U7103 (N_7103,N_3103,N_4072);
nor U7104 (N_7104,N_4433,N_5797);
nor U7105 (N_7105,N_3024,N_3473);
and U7106 (N_7106,N_4367,N_4865);
and U7107 (N_7107,N_4133,N_3880);
nor U7108 (N_7108,N_4703,N_3968);
nand U7109 (N_7109,N_4446,N_4185);
and U7110 (N_7110,N_5564,N_5164);
or U7111 (N_7111,N_3672,N_5864);
or U7112 (N_7112,N_4908,N_5444);
nor U7113 (N_7113,N_3040,N_5672);
nand U7114 (N_7114,N_3413,N_4165);
and U7115 (N_7115,N_3064,N_3650);
or U7116 (N_7116,N_4461,N_3402);
or U7117 (N_7117,N_3995,N_5005);
and U7118 (N_7118,N_3989,N_4825);
nor U7119 (N_7119,N_3903,N_5147);
or U7120 (N_7120,N_4061,N_5756);
nor U7121 (N_7121,N_5767,N_4269);
and U7122 (N_7122,N_4155,N_5151);
nor U7123 (N_7123,N_4497,N_5773);
nand U7124 (N_7124,N_3036,N_4218);
nor U7125 (N_7125,N_5725,N_5340);
or U7126 (N_7126,N_3492,N_4477);
or U7127 (N_7127,N_5631,N_5480);
and U7128 (N_7128,N_5455,N_4939);
or U7129 (N_7129,N_3272,N_5613);
nand U7130 (N_7130,N_3573,N_4779);
and U7131 (N_7131,N_4946,N_3825);
or U7132 (N_7132,N_3448,N_5843);
and U7133 (N_7133,N_3784,N_5446);
nor U7134 (N_7134,N_5423,N_4213);
or U7135 (N_7135,N_5027,N_3073);
and U7136 (N_7136,N_4469,N_3083);
nor U7137 (N_7137,N_5120,N_3582);
nand U7138 (N_7138,N_3586,N_5148);
nor U7139 (N_7139,N_3277,N_5119);
nor U7140 (N_7140,N_3615,N_3198);
or U7141 (N_7141,N_3641,N_5123);
and U7142 (N_7142,N_4387,N_3706);
nor U7143 (N_7143,N_5281,N_3014);
nand U7144 (N_7144,N_5474,N_4871);
or U7145 (N_7145,N_3769,N_4975);
nor U7146 (N_7146,N_5080,N_5396);
nor U7147 (N_7147,N_4501,N_4036);
nor U7148 (N_7148,N_4910,N_4550);
nor U7149 (N_7149,N_3481,N_5204);
nand U7150 (N_7150,N_5265,N_4556);
nor U7151 (N_7151,N_3621,N_3704);
and U7152 (N_7152,N_3893,N_3526);
and U7153 (N_7153,N_4444,N_3922);
and U7154 (N_7154,N_5879,N_3459);
and U7155 (N_7155,N_5573,N_5971);
or U7156 (N_7156,N_5108,N_5647);
or U7157 (N_7157,N_3300,N_5113);
and U7158 (N_7158,N_4674,N_4711);
and U7159 (N_7159,N_3625,N_3629);
or U7160 (N_7160,N_4759,N_5812);
or U7161 (N_7161,N_3554,N_4230);
or U7162 (N_7162,N_3665,N_5110);
nor U7163 (N_7163,N_5743,N_3136);
and U7164 (N_7164,N_3816,N_5433);
xor U7165 (N_7165,N_5719,N_4769);
or U7166 (N_7166,N_3140,N_4546);
nand U7167 (N_7167,N_4415,N_3509);
nand U7168 (N_7168,N_3815,N_3219);
nor U7169 (N_7169,N_4391,N_3098);
and U7170 (N_7170,N_4385,N_3246);
and U7171 (N_7171,N_4637,N_4833);
nor U7172 (N_7172,N_3581,N_4506);
or U7173 (N_7173,N_4774,N_4592);
and U7174 (N_7174,N_3630,N_5202);
nor U7175 (N_7175,N_4913,N_4080);
nand U7176 (N_7176,N_3392,N_3178);
or U7177 (N_7177,N_3189,N_5169);
nor U7178 (N_7178,N_3386,N_4380);
nand U7179 (N_7179,N_4494,N_3451);
xor U7180 (N_7180,N_5544,N_4068);
nor U7181 (N_7181,N_3002,N_5318);
nor U7182 (N_7182,N_4228,N_3028);
or U7183 (N_7183,N_4127,N_5409);
nand U7184 (N_7184,N_4885,N_3729);
nand U7185 (N_7185,N_3357,N_5130);
nor U7186 (N_7186,N_4898,N_5836);
or U7187 (N_7187,N_4586,N_4322);
nand U7188 (N_7188,N_3376,N_4336);
or U7189 (N_7189,N_3920,N_4309);
and U7190 (N_7190,N_4344,N_5908);
nor U7191 (N_7191,N_5326,N_5619);
or U7192 (N_7192,N_3782,N_3275);
nor U7193 (N_7193,N_5701,N_3856);
or U7194 (N_7194,N_5579,N_5099);
or U7195 (N_7195,N_4614,N_3499);
nor U7196 (N_7196,N_3111,N_5302);
nand U7197 (N_7197,N_4752,N_5144);
nand U7198 (N_7198,N_5029,N_4455);
or U7199 (N_7199,N_3733,N_4953);
nand U7200 (N_7200,N_3528,N_4000);
nor U7201 (N_7201,N_5279,N_4805);
nor U7202 (N_7202,N_5734,N_3887);
or U7203 (N_7203,N_3703,N_5500);
nand U7204 (N_7204,N_4323,N_3282);
nor U7205 (N_7205,N_5556,N_4459);
or U7206 (N_7206,N_5171,N_5434);
or U7207 (N_7207,N_4381,N_4632);
nand U7208 (N_7208,N_5495,N_4425);
nand U7209 (N_7209,N_5343,N_4599);
or U7210 (N_7210,N_4848,N_5328);
and U7211 (N_7211,N_4552,N_4170);
or U7212 (N_7212,N_4419,N_4707);
or U7213 (N_7213,N_3131,N_4408);
nor U7214 (N_7214,N_3166,N_5124);
nand U7215 (N_7215,N_3639,N_4978);
and U7216 (N_7216,N_4280,N_4616);
nor U7217 (N_7217,N_3082,N_5251);
nor U7218 (N_7218,N_4404,N_3407);
or U7219 (N_7219,N_4533,N_5935);
nor U7220 (N_7220,N_4084,N_5407);
nor U7221 (N_7221,N_5293,N_5078);
nor U7222 (N_7222,N_5494,N_5178);
and U7223 (N_7223,N_4977,N_5392);
or U7224 (N_7224,N_5163,N_3948);
or U7225 (N_7225,N_3500,N_3921);
or U7226 (N_7226,N_5157,N_3420);
nor U7227 (N_7227,N_3741,N_4697);
nand U7228 (N_7228,N_5981,N_4274);
nand U7229 (N_7229,N_5595,N_4929);
and U7230 (N_7230,N_5142,N_4956);
nor U7231 (N_7231,N_4862,N_4160);
nand U7232 (N_7232,N_4549,N_4135);
nand U7233 (N_7233,N_3843,N_3023);
nand U7234 (N_7234,N_4321,N_3401);
or U7235 (N_7235,N_5348,N_5043);
or U7236 (N_7236,N_4289,N_5678);
nor U7237 (N_7237,N_5586,N_5515);
and U7238 (N_7238,N_5670,N_3585);
or U7239 (N_7239,N_4526,N_5805);
or U7240 (N_7240,N_4952,N_4803);
nand U7241 (N_7241,N_5062,N_4263);
or U7242 (N_7242,N_4984,N_3905);
nor U7243 (N_7243,N_4651,N_5289);
nand U7244 (N_7244,N_4796,N_3869);
or U7245 (N_7245,N_3864,N_4761);
nor U7246 (N_7246,N_4608,N_3105);
or U7247 (N_7247,N_3329,N_3692);
nor U7248 (N_7248,N_3327,N_5574);
nor U7249 (N_7249,N_5193,N_5930);
or U7250 (N_7250,N_4888,N_4118);
or U7251 (N_7251,N_3555,N_3320);
or U7252 (N_7252,N_5944,N_5936);
nor U7253 (N_7253,N_3668,N_3089);
nand U7254 (N_7254,N_4307,N_5089);
nand U7255 (N_7255,N_4940,N_5561);
or U7256 (N_7256,N_3463,N_3055);
and U7257 (N_7257,N_5344,N_5733);
and U7258 (N_7258,N_4101,N_5616);
or U7259 (N_7259,N_3005,N_4789);
and U7260 (N_7260,N_5305,N_5940);
nor U7261 (N_7261,N_5904,N_3611);
or U7262 (N_7262,N_3185,N_3148);
nand U7263 (N_7263,N_4570,N_5508);
and U7264 (N_7264,N_3652,N_4916);
or U7265 (N_7265,N_3768,N_4150);
or U7266 (N_7266,N_3264,N_4113);
nand U7267 (N_7267,N_5869,N_5187);
and U7268 (N_7268,N_5061,N_4161);
or U7269 (N_7269,N_3827,N_5366);
nor U7270 (N_7270,N_5047,N_5765);
and U7271 (N_7271,N_3531,N_4766);
nand U7272 (N_7272,N_4003,N_4102);
xnor U7273 (N_7273,N_4931,N_4566);
and U7274 (N_7274,N_5553,N_3071);
and U7275 (N_7275,N_5541,N_3066);
nor U7276 (N_7276,N_4296,N_4942);
nand U7277 (N_7277,N_4260,N_3333);
or U7278 (N_7278,N_4528,N_4109);
nand U7279 (N_7279,N_4291,N_4090);
and U7280 (N_7280,N_5388,N_3858);
nor U7281 (N_7281,N_5891,N_5566);
or U7282 (N_7282,N_5596,N_5905);
and U7283 (N_7283,N_4524,N_3529);
or U7284 (N_7284,N_3888,N_4407);
nor U7285 (N_7285,N_4443,N_5006);
nor U7286 (N_7286,N_5191,N_5692);
nor U7287 (N_7287,N_5532,N_3605);
nand U7288 (N_7288,N_3543,N_5212);
and U7289 (N_7289,N_5033,N_4877);
nand U7290 (N_7290,N_4193,N_4128);
nor U7291 (N_7291,N_5970,N_5476);
and U7292 (N_7292,N_3943,N_4203);
nand U7293 (N_7293,N_3666,N_5895);
xor U7294 (N_7294,N_5351,N_5853);
and U7295 (N_7295,N_3633,N_5001);
nor U7296 (N_7296,N_3119,N_5831);
nand U7297 (N_7297,N_3115,N_3163);
nand U7298 (N_7298,N_3491,N_5629);
nand U7299 (N_7299,N_3081,N_5705);
nand U7300 (N_7300,N_5673,N_5081);
or U7301 (N_7301,N_4025,N_4767);
or U7302 (N_7302,N_5304,N_4914);
and U7303 (N_7303,N_4572,N_4654);
or U7304 (N_7304,N_5277,N_5762);
and U7305 (N_7305,N_3616,N_4098);
or U7306 (N_7306,N_3484,N_5129);
nand U7307 (N_7307,N_5641,N_5680);
nand U7308 (N_7308,N_4604,N_3410);
nor U7309 (N_7309,N_4718,N_5531);
nand U7310 (N_7310,N_5121,N_4377);
or U7311 (N_7311,N_4319,N_5079);
or U7312 (N_7312,N_3403,N_5861);
nand U7313 (N_7313,N_4653,N_5367);
nor U7314 (N_7314,N_3424,N_5644);
nand U7315 (N_7315,N_3476,N_3323);
nand U7316 (N_7316,N_4790,N_5363);
nand U7317 (N_7317,N_4383,N_4149);
nor U7318 (N_7318,N_3045,N_5257);
or U7319 (N_7319,N_4453,N_4958);
and U7320 (N_7320,N_5155,N_5133);
or U7321 (N_7321,N_4019,N_5849);
nor U7322 (N_7322,N_3155,N_4167);
nand U7323 (N_7323,N_5131,N_5704);
or U7324 (N_7324,N_3689,N_3091);
nand U7325 (N_7325,N_3343,N_3929);
and U7326 (N_7326,N_4547,N_5436);
and U7327 (N_7327,N_3607,N_3532);
and U7328 (N_7328,N_3977,N_5963);
nor U7329 (N_7329,N_4562,N_4424);
and U7330 (N_7330,N_3656,N_4121);
nor U7331 (N_7331,N_4159,N_4530);
nor U7332 (N_7332,N_5338,N_5676);
or U7333 (N_7333,N_3477,N_5167);
and U7334 (N_7334,N_3906,N_3069);
nor U7335 (N_7335,N_4527,N_5522);
or U7336 (N_7336,N_5588,N_3958);
nand U7337 (N_7337,N_3428,N_5807);
and U7338 (N_7338,N_4060,N_3238);
or U7339 (N_7339,N_5834,N_3728);
nor U7340 (N_7340,N_3174,N_5707);
nor U7341 (N_7341,N_5308,N_3796);
or U7342 (N_7342,N_4449,N_5499);
nor U7343 (N_7343,N_3143,N_4725);
and U7344 (N_7344,N_4754,N_5938);
xnor U7345 (N_7345,N_4522,N_3183);
nand U7346 (N_7346,N_5028,N_5637);
nor U7347 (N_7347,N_5867,N_3897);
or U7348 (N_7348,N_4271,N_4175);
or U7349 (N_7349,N_3519,N_4298);
or U7350 (N_7350,N_3746,N_5929);
or U7351 (N_7351,N_5046,N_3936);
nor U7352 (N_7352,N_3739,N_3508);
nand U7353 (N_7353,N_4849,N_5732);
xnor U7354 (N_7354,N_4741,N_4537);
or U7355 (N_7355,N_5934,N_5249);
nand U7356 (N_7356,N_3804,N_4130);
and U7357 (N_7357,N_3007,N_5987);
nand U7358 (N_7358,N_5013,N_4011);
nand U7359 (N_7359,N_5430,N_5214);
nor U7360 (N_7360,N_5153,N_5824);
nor U7361 (N_7361,N_4612,N_3525);
nand U7362 (N_7362,N_4476,N_3145);
and U7363 (N_7363,N_5630,N_4539);
nand U7364 (N_7364,N_5342,N_5691);
nand U7365 (N_7365,N_3137,N_3882);
nand U7366 (N_7366,N_4071,N_5103);
nand U7367 (N_7367,N_3870,N_4473);
nand U7368 (N_7368,N_5950,N_4439);
nand U7369 (N_7369,N_4337,N_5736);
nor U7370 (N_7370,N_3294,N_3941);
nand U7371 (N_7371,N_3584,N_4700);
nor U7372 (N_7372,N_3284,N_4747);
nor U7373 (N_7373,N_5988,N_3660);
nand U7374 (N_7374,N_4279,N_4281);
or U7375 (N_7375,N_5438,N_4389);
and U7376 (N_7376,N_3590,N_3749);
nand U7377 (N_7377,N_4583,N_3287);
and U7378 (N_7378,N_4875,N_4571);
and U7379 (N_7379,N_3833,N_4729);
nand U7380 (N_7380,N_3317,N_5095);
nand U7381 (N_7381,N_3170,N_5643);
nor U7382 (N_7382,N_3832,N_5406);
nand U7383 (N_7383,N_4214,N_3683);
or U7384 (N_7384,N_5565,N_5228);
nor U7385 (N_7385,N_3460,N_3274);
nor U7386 (N_7386,N_3244,N_3699);
nor U7387 (N_7387,N_5937,N_5060);
or U7388 (N_7388,N_5664,N_4148);
nand U7389 (N_7389,N_3331,N_4422);
nor U7390 (N_7390,N_3496,N_4720);
nand U7391 (N_7391,N_3245,N_3541);
nand U7392 (N_7392,N_3830,N_5537);
nand U7393 (N_7393,N_4824,N_5288);
or U7394 (N_7394,N_4786,N_3192);
nand U7395 (N_7395,N_3992,N_4679);
and U7396 (N_7396,N_3302,N_4983);
and U7397 (N_7397,N_5229,N_4944);
nand U7398 (N_7398,N_5612,N_4655);
or U7399 (N_7399,N_4044,N_5959);
or U7400 (N_7400,N_3892,N_5639);
nor U7401 (N_7401,N_5450,N_4732);
or U7402 (N_7402,N_4631,N_5141);
nor U7403 (N_7403,N_4907,N_5442);
or U7404 (N_7404,N_3293,N_4190);
or U7405 (N_7405,N_5730,N_5440);
nor U7406 (N_7406,N_5888,N_3812);
or U7407 (N_7407,N_3805,N_3364);
and U7408 (N_7408,N_3021,N_5993);
and U7409 (N_7409,N_3599,N_5286);
and U7410 (N_7410,N_4210,N_3471);
nand U7411 (N_7411,N_3374,N_3063);
or U7412 (N_7412,N_3224,N_4335);
nand U7413 (N_7413,N_5858,N_4405);
or U7414 (N_7414,N_4376,N_5024);
and U7415 (N_7415,N_4474,N_5606);
or U7416 (N_7416,N_4840,N_4785);
or U7417 (N_7417,N_5381,N_4792);
nand U7418 (N_7418,N_4268,N_5659);
nand U7419 (N_7419,N_5968,N_4365);
nand U7420 (N_7420,N_3885,N_5485);
nor U7421 (N_7421,N_4318,N_5645);
and U7422 (N_7422,N_4241,N_4924);
or U7423 (N_7423,N_5268,N_3281);
nand U7424 (N_7424,N_3251,N_4191);
and U7425 (N_7425,N_3422,N_4739);
nor U7426 (N_7426,N_5838,N_4491);
and U7427 (N_7427,N_5960,N_5460);
and U7428 (N_7428,N_3483,N_3283);
or U7429 (N_7429,N_3160,N_4320);
nand U7430 (N_7430,N_4897,N_5176);
and U7431 (N_7431,N_3783,N_3811);
and U7432 (N_7432,N_3662,N_4416);
nand U7433 (N_7433,N_4077,N_5181);
nor U7434 (N_7434,N_4362,N_3755);
or U7435 (N_7435,N_5075,N_5724);
nand U7436 (N_7436,N_5426,N_5638);
or U7437 (N_7437,N_4962,N_5232);
nor U7438 (N_7438,N_3099,N_5894);
nor U7439 (N_7439,N_5465,N_4308);
nand U7440 (N_7440,N_5002,N_4114);
nor U7441 (N_7441,N_3618,N_3117);
or U7442 (N_7442,N_4286,N_3757);
nand U7443 (N_7443,N_4087,N_5276);
nor U7444 (N_7444,N_4169,N_5070);
or U7445 (N_7445,N_3593,N_5962);
nor U7446 (N_7446,N_5059,N_4456);
or U7447 (N_7447,N_3507,N_3372);
or U7448 (N_7448,N_4686,N_3406);
nand U7449 (N_7449,N_5840,N_4056);
nor U7450 (N_7450,N_4535,N_4388);
or U7451 (N_7451,N_5552,N_3180);
nand U7452 (N_7452,N_3479,N_5675);
xor U7453 (N_7453,N_3592,N_4162);
nand U7454 (N_7454,N_4909,N_5562);
nor U7455 (N_7455,N_4031,N_3240);
nand U7456 (N_7456,N_5401,N_5669);
nand U7457 (N_7457,N_3127,N_3265);
or U7458 (N_7458,N_3550,N_4843);
nor U7459 (N_7459,N_3122,N_4462);
and U7460 (N_7460,N_5483,N_3938);
nand U7461 (N_7461,N_4198,N_5140);
or U7462 (N_7462,N_4735,N_5966);
and U7463 (N_7463,N_5182,N_3090);
and U7464 (N_7464,N_3497,N_3161);
or U7465 (N_7465,N_4301,N_4744);
nand U7466 (N_7466,N_3400,N_4284);
nand U7467 (N_7467,N_5194,N_3698);
nor U7468 (N_7468,N_4626,N_3295);
and U7469 (N_7469,N_5139,N_5850);
or U7470 (N_7470,N_3937,N_4661);
or U7471 (N_7471,N_3503,N_5972);
or U7472 (N_7472,N_5593,N_5098);
and U7473 (N_7473,N_4812,N_4965);
and U7474 (N_7474,N_3852,N_3824);
nor U7475 (N_7475,N_4270,N_4705);
and U7476 (N_7476,N_4500,N_5974);
nor U7477 (N_7477,N_3278,N_5885);
nand U7478 (N_7478,N_5570,N_3957);
or U7479 (N_7479,N_3537,N_5067);
and U7480 (N_7480,N_4059,N_4173);
nand U7481 (N_7481,N_4823,N_5076);
and U7482 (N_7482,N_5626,N_3575);
nor U7483 (N_7483,N_4541,N_4904);
and U7484 (N_7484,N_3197,N_3354);
and U7485 (N_7485,N_5820,N_4282);
nor U7486 (N_7486,N_4242,N_3932);
or U7487 (N_7487,N_4678,N_4047);
and U7488 (N_7488,N_4936,N_3866);
and U7489 (N_7489,N_5546,N_4423);
and U7490 (N_7490,N_4531,N_3814);
and U7491 (N_7491,N_3993,N_5536);
or U7492 (N_7492,N_4988,N_5948);
nand U7493 (N_7493,N_3067,N_4638);
or U7494 (N_7494,N_4536,N_3642);
nor U7495 (N_7495,N_3129,N_4037);
and U7496 (N_7496,N_4312,N_5077);
or U7497 (N_7497,N_4020,N_5918);
nand U7498 (N_7498,N_3688,N_4542);
nor U7499 (N_7499,N_4332,N_5883);
and U7500 (N_7500,N_4749,N_4556);
or U7501 (N_7501,N_4391,N_5810);
nor U7502 (N_7502,N_3741,N_4281);
or U7503 (N_7503,N_4082,N_3612);
nand U7504 (N_7504,N_4027,N_5481);
nand U7505 (N_7505,N_4303,N_3265);
and U7506 (N_7506,N_5744,N_4587);
or U7507 (N_7507,N_3776,N_4310);
and U7508 (N_7508,N_4479,N_3310);
nand U7509 (N_7509,N_5587,N_4704);
and U7510 (N_7510,N_3942,N_4188);
nand U7511 (N_7511,N_5086,N_5406);
nor U7512 (N_7512,N_3316,N_5983);
nor U7513 (N_7513,N_3460,N_5695);
xor U7514 (N_7514,N_3988,N_3440);
and U7515 (N_7515,N_3250,N_3880);
and U7516 (N_7516,N_5376,N_5732);
or U7517 (N_7517,N_5577,N_3185);
or U7518 (N_7518,N_5148,N_5994);
nand U7519 (N_7519,N_4853,N_4200);
or U7520 (N_7520,N_5559,N_3039);
or U7521 (N_7521,N_4171,N_5506);
nand U7522 (N_7522,N_4307,N_5467);
nand U7523 (N_7523,N_5253,N_4097);
nand U7524 (N_7524,N_3284,N_4952);
nand U7525 (N_7525,N_4906,N_4625);
or U7526 (N_7526,N_3922,N_4566);
xnor U7527 (N_7527,N_5977,N_5786);
nand U7528 (N_7528,N_5171,N_4169);
and U7529 (N_7529,N_4939,N_3169);
nor U7530 (N_7530,N_3699,N_4953);
nor U7531 (N_7531,N_4832,N_4970);
xor U7532 (N_7532,N_3671,N_5259);
nand U7533 (N_7533,N_5225,N_4833);
or U7534 (N_7534,N_3563,N_4719);
nand U7535 (N_7535,N_5949,N_5877);
nor U7536 (N_7536,N_4954,N_3939);
and U7537 (N_7537,N_4354,N_3036);
nand U7538 (N_7538,N_3923,N_3742);
nand U7539 (N_7539,N_4736,N_3914);
or U7540 (N_7540,N_3323,N_4944);
or U7541 (N_7541,N_3082,N_3070);
nor U7542 (N_7542,N_4105,N_5956);
nor U7543 (N_7543,N_5540,N_5139);
xor U7544 (N_7544,N_4166,N_5199);
and U7545 (N_7545,N_4650,N_3696);
nand U7546 (N_7546,N_4757,N_4330);
nand U7547 (N_7547,N_3382,N_5202);
nand U7548 (N_7548,N_3246,N_5631);
nand U7549 (N_7549,N_5414,N_3004);
nand U7550 (N_7550,N_5524,N_3311);
and U7551 (N_7551,N_4664,N_4648);
nand U7552 (N_7552,N_3098,N_5469);
or U7553 (N_7553,N_4254,N_5650);
or U7554 (N_7554,N_5622,N_5056);
nor U7555 (N_7555,N_5379,N_5542);
or U7556 (N_7556,N_4332,N_3015);
nor U7557 (N_7557,N_4354,N_4821);
nand U7558 (N_7558,N_3407,N_4492);
or U7559 (N_7559,N_4944,N_3161);
nand U7560 (N_7560,N_3607,N_4699);
and U7561 (N_7561,N_3346,N_3184);
nand U7562 (N_7562,N_3145,N_5599);
nand U7563 (N_7563,N_5747,N_4523);
nand U7564 (N_7564,N_3588,N_4859);
nand U7565 (N_7565,N_4819,N_4945);
or U7566 (N_7566,N_5036,N_3726);
nand U7567 (N_7567,N_3696,N_5734);
nand U7568 (N_7568,N_5283,N_4222);
or U7569 (N_7569,N_5222,N_5079);
and U7570 (N_7570,N_5581,N_4135);
or U7571 (N_7571,N_4786,N_3014);
nor U7572 (N_7572,N_5022,N_3393);
nand U7573 (N_7573,N_3194,N_4310);
nor U7574 (N_7574,N_5531,N_3294);
xnor U7575 (N_7575,N_5061,N_5982);
nand U7576 (N_7576,N_5397,N_3916);
or U7577 (N_7577,N_5832,N_5200);
or U7578 (N_7578,N_5365,N_4149);
nor U7579 (N_7579,N_3851,N_5107);
or U7580 (N_7580,N_5709,N_3247);
nand U7581 (N_7581,N_3383,N_3211);
nor U7582 (N_7582,N_3711,N_5391);
and U7583 (N_7583,N_4657,N_3485);
or U7584 (N_7584,N_5289,N_3038);
nand U7585 (N_7585,N_3755,N_3560);
or U7586 (N_7586,N_4575,N_3262);
and U7587 (N_7587,N_5941,N_5504);
and U7588 (N_7588,N_5957,N_5831);
nand U7589 (N_7589,N_3941,N_4706);
or U7590 (N_7590,N_3518,N_4285);
or U7591 (N_7591,N_5222,N_5045);
nor U7592 (N_7592,N_3423,N_5209);
nor U7593 (N_7593,N_5045,N_5932);
nor U7594 (N_7594,N_4243,N_4461);
nor U7595 (N_7595,N_5471,N_3645);
nand U7596 (N_7596,N_3594,N_4911);
and U7597 (N_7597,N_5414,N_4579);
nand U7598 (N_7598,N_4862,N_4046);
and U7599 (N_7599,N_4101,N_3432);
nor U7600 (N_7600,N_3840,N_5456);
nand U7601 (N_7601,N_3197,N_5556);
or U7602 (N_7602,N_4614,N_3008);
nor U7603 (N_7603,N_3300,N_3084);
and U7604 (N_7604,N_3791,N_3694);
or U7605 (N_7605,N_5113,N_5353);
xor U7606 (N_7606,N_5359,N_3698);
nor U7607 (N_7607,N_3958,N_5777);
and U7608 (N_7608,N_5285,N_4021);
and U7609 (N_7609,N_5751,N_5556);
nor U7610 (N_7610,N_3567,N_4569);
nor U7611 (N_7611,N_5132,N_4078);
or U7612 (N_7612,N_5960,N_5559);
nand U7613 (N_7613,N_4641,N_4223);
or U7614 (N_7614,N_3327,N_3929);
nand U7615 (N_7615,N_4260,N_3435);
nand U7616 (N_7616,N_3071,N_3364);
nand U7617 (N_7617,N_4215,N_5858);
or U7618 (N_7618,N_5417,N_3151);
or U7619 (N_7619,N_5288,N_3434);
nor U7620 (N_7620,N_3190,N_5089);
nor U7621 (N_7621,N_3157,N_3146);
nand U7622 (N_7622,N_5427,N_5616);
nand U7623 (N_7623,N_4500,N_5006);
xor U7624 (N_7624,N_3750,N_4744);
and U7625 (N_7625,N_5617,N_3307);
nand U7626 (N_7626,N_4460,N_4963);
and U7627 (N_7627,N_3763,N_5691);
or U7628 (N_7628,N_3520,N_4289);
or U7629 (N_7629,N_3018,N_5045);
and U7630 (N_7630,N_3008,N_3117);
nand U7631 (N_7631,N_3223,N_4366);
and U7632 (N_7632,N_5149,N_5755);
nor U7633 (N_7633,N_3705,N_3624);
or U7634 (N_7634,N_3809,N_3939);
nand U7635 (N_7635,N_5674,N_5126);
or U7636 (N_7636,N_5480,N_3364);
nor U7637 (N_7637,N_3547,N_3947);
nand U7638 (N_7638,N_5588,N_4925);
or U7639 (N_7639,N_5945,N_5181);
or U7640 (N_7640,N_3454,N_5516);
or U7641 (N_7641,N_3546,N_5577);
or U7642 (N_7642,N_4671,N_3443);
nor U7643 (N_7643,N_5067,N_3620);
and U7644 (N_7644,N_5802,N_4894);
nor U7645 (N_7645,N_5869,N_4491);
and U7646 (N_7646,N_5999,N_3597);
and U7647 (N_7647,N_4874,N_4814);
nor U7648 (N_7648,N_4708,N_5466);
and U7649 (N_7649,N_5162,N_4750);
nand U7650 (N_7650,N_5193,N_5212);
nand U7651 (N_7651,N_3820,N_4765);
nand U7652 (N_7652,N_4898,N_5988);
and U7653 (N_7653,N_3939,N_3512);
nor U7654 (N_7654,N_5294,N_5117);
and U7655 (N_7655,N_3267,N_3058);
nor U7656 (N_7656,N_3665,N_3065);
nand U7657 (N_7657,N_5051,N_3253);
or U7658 (N_7658,N_3761,N_3541);
nor U7659 (N_7659,N_4984,N_5250);
and U7660 (N_7660,N_5364,N_4515);
and U7661 (N_7661,N_4270,N_3045);
and U7662 (N_7662,N_5349,N_4115);
or U7663 (N_7663,N_5650,N_3938);
nand U7664 (N_7664,N_5442,N_5847);
nand U7665 (N_7665,N_4028,N_4295);
or U7666 (N_7666,N_5237,N_3403);
or U7667 (N_7667,N_4441,N_4282);
or U7668 (N_7668,N_4424,N_3496);
and U7669 (N_7669,N_3219,N_4963);
nor U7670 (N_7670,N_3122,N_3726);
nor U7671 (N_7671,N_5480,N_3771);
and U7672 (N_7672,N_5944,N_3960);
nor U7673 (N_7673,N_4294,N_5267);
and U7674 (N_7674,N_5851,N_3607);
nand U7675 (N_7675,N_3161,N_4380);
nand U7676 (N_7676,N_3634,N_5422);
or U7677 (N_7677,N_3033,N_4412);
nor U7678 (N_7678,N_5764,N_4451);
or U7679 (N_7679,N_4124,N_3192);
nand U7680 (N_7680,N_4404,N_4688);
and U7681 (N_7681,N_3675,N_3989);
and U7682 (N_7682,N_4851,N_5813);
nand U7683 (N_7683,N_4713,N_4901);
nor U7684 (N_7684,N_4323,N_5581);
or U7685 (N_7685,N_4131,N_4776);
nand U7686 (N_7686,N_5432,N_5356);
and U7687 (N_7687,N_4163,N_4687);
nor U7688 (N_7688,N_3434,N_3178);
nor U7689 (N_7689,N_3274,N_5696);
nand U7690 (N_7690,N_4921,N_4428);
and U7691 (N_7691,N_3383,N_5482);
nand U7692 (N_7692,N_4268,N_5455);
or U7693 (N_7693,N_4418,N_4301);
or U7694 (N_7694,N_3202,N_3437);
nor U7695 (N_7695,N_3973,N_5276);
or U7696 (N_7696,N_3212,N_4215);
or U7697 (N_7697,N_4258,N_4460);
and U7698 (N_7698,N_3580,N_3419);
nor U7699 (N_7699,N_4387,N_4161);
nor U7700 (N_7700,N_3882,N_3711);
or U7701 (N_7701,N_4313,N_3040);
nor U7702 (N_7702,N_3798,N_4147);
nor U7703 (N_7703,N_4365,N_5474);
nand U7704 (N_7704,N_3241,N_5186);
and U7705 (N_7705,N_4340,N_3161);
and U7706 (N_7706,N_3078,N_5632);
nor U7707 (N_7707,N_5813,N_5753);
nand U7708 (N_7708,N_5712,N_4421);
and U7709 (N_7709,N_4022,N_5681);
nand U7710 (N_7710,N_3671,N_4611);
nand U7711 (N_7711,N_3275,N_3625);
nand U7712 (N_7712,N_3709,N_5956);
or U7713 (N_7713,N_4684,N_5582);
nand U7714 (N_7714,N_5215,N_5703);
or U7715 (N_7715,N_3464,N_5182);
and U7716 (N_7716,N_3245,N_5388);
xor U7717 (N_7717,N_4183,N_4972);
nor U7718 (N_7718,N_4910,N_4968);
nand U7719 (N_7719,N_5052,N_5785);
and U7720 (N_7720,N_4128,N_3536);
and U7721 (N_7721,N_3090,N_4704);
nor U7722 (N_7722,N_5892,N_4688);
nor U7723 (N_7723,N_3976,N_4096);
nor U7724 (N_7724,N_4196,N_5350);
nand U7725 (N_7725,N_4303,N_4492);
or U7726 (N_7726,N_5017,N_3315);
and U7727 (N_7727,N_4478,N_5375);
nand U7728 (N_7728,N_4381,N_4489);
or U7729 (N_7729,N_5010,N_3355);
nand U7730 (N_7730,N_4536,N_5260);
or U7731 (N_7731,N_5583,N_5668);
nor U7732 (N_7732,N_3916,N_3944);
or U7733 (N_7733,N_4690,N_5035);
nand U7734 (N_7734,N_4436,N_4531);
and U7735 (N_7735,N_3815,N_5668);
and U7736 (N_7736,N_5802,N_5047);
or U7737 (N_7737,N_3079,N_5107);
and U7738 (N_7738,N_5745,N_4673);
nand U7739 (N_7739,N_4958,N_5715);
nand U7740 (N_7740,N_4207,N_3060);
and U7741 (N_7741,N_5968,N_4904);
or U7742 (N_7742,N_5059,N_3320);
nor U7743 (N_7743,N_5076,N_4915);
nor U7744 (N_7744,N_5823,N_5711);
or U7745 (N_7745,N_3167,N_5620);
nand U7746 (N_7746,N_3792,N_4330);
nor U7747 (N_7747,N_5055,N_3743);
xor U7748 (N_7748,N_3256,N_3157);
or U7749 (N_7749,N_4278,N_5417);
nor U7750 (N_7750,N_4418,N_5664);
and U7751 (N_7751,N_3375,N_5188);
nor U7752 (N_7752,N_5889,N_3401);
nand U7753 (N_7753,N_3376,N_3205);
or U7754 (N_7754,N_5588,N_3310);
nand U7755 (N_7755,N_4613,N_3615);
nand U7756 (N_7756,N_5053,N_3772);
nor U7757 (N_7757,N_4996,N_4413);
or U7758 (N_7758,N_4027,N_4769);
or U7759 (N_7759,N_5647,N_4566);
nor U7760 (N_7760,N_3662,N_5861);
nand U7761 (N_7761,N_5076,N_3153);
nand U7762 (N_7762,N_3417,N_5551);
nor U7763 (N_7763,N_3043,N_4994);
and U7764 (N_7764,N_4419,N_5417);
nand U7765 (N_7765,N_5106,N_4804);
nand U7766 (N_7766,N_5972,N_3210);
or U7767 (N_7767,N_4729,N_3102);
and U7768 (N_7768,N_3552,N_4332);
and U7769 (N_7769,N_3526,N_4141);
nand U7770 (N_7770,N_3626,N_5360);
or U7771 (N_7771,N_4852,N_4164);
nor U7772 (N_7772,N_3728,N_3968);
or U7773 (N_7773,N_3997,N_4729);
or U7774 (N_7774,N_3126,N_5408);
nor U7775 (N_7775,N_4713,N_3253);
nand U7776 (N_7776,N_3259,N_4837);
nor U7777 (N_7777,N_5407,N_5217);
nand U7778 (N_7778,N_3739,N_4186);
nor U7779 (N_7779,N_4339,N_3122);
or U7780 (N_7780,N_5431,N_5912);
or U7781 (N_7781,N_5164,N_3677);
nor U7782 (N_7782,N_5509,N_3327);
and U7783 (N_7783,N_5251,N_3540);
nor U7784 (N_7784,N_3386,N_5935);
or U7785 (N_7785,N_4188,N_4737);
or U7786 (N_7786,N_4891,N_5324);
or U7787 (N_7787,N_3904,N_4612);
nor U7788 (N_7788,N_3058,N_4667);
nand U7789 (N_7789,N_4419,N_4260);
nor U7790 (N_7790,N_3721,N_4771);
and U7791 (N_7791,N_4142,N_4910);
nand U7792 (N_7792,N_4922,N_3626);
nor U7793 (N_7793,N_4337,N_4352);
nor U7794 (N_7794,N_4185,N_3954);
xor U7795 (N_7795,N_4709,N_5902);
or U7796 (N_7796,N_4355,N_5371);
nor U7797 (N_7797,N_3839,N_5120);
and U7798 (N_7798,N_4052,N_4891);
xnor U7799 (N_7799,N_4259,N_4385);
or U7800 (N_7800,N_4349,N_3481);
nand U7801 (N_7801,N_4011,N_3684);
and U7802 (N_7802,N_3260,N_5585);
or U7803 (N_7803,N_4859,N_3030);
or U7804 (N_7804,N_4102,N_5516);
nor U7805 (N_7805,N_5397,N_4428);
nand U7806 (N_7806,N_5001,N_5268);
and U7807 (N_7807,N_4921,N_4108);
xor U7808 (N_7808,N_3679,N_4674);
nand U7809 (N_7809,N_4997,N_5306);
nor U7810 (N_7810,N_4371,N_4139);
nor U7811 (N_7811,N_3327,N_5458);
nand U7812 (N_7812,N_5566,N_3193);
nand U7813 (N_7813,N_4540,N_4211);
or U7814 (N_7814,N_4640,N_3373);
or U7815 (N_7815,N_5446,N_4793);
or U7816 (N_7816,N_4103,N_3232);
or U7817 (N_7817,N_4546,N_5519);
nor U7818 (N_7818,N_4000,N_4220);
and U7819 (N_7819,N_5014,N_3641);
and U7820 (N_7820,N_4286,N_4375);
and U7821 (N_7821,N_5788,N_5028);
or U7822 (N_7822,N_5296,N_3678);
nor U7823 (N_7823,N_5965,N_4840);
and U7824 (N_7824,N_5155,N_5822);
nor U7825 (N_7825,N_4492,N_3310);
or U7826 (N_7826,N_3429,N_3265);
nand U7827 (N_7827,N_5975,N_3111);
nand U7828 (N_7828,N_4146,N_5313);
nor U7829 (N_7829,N_4573,N_5395);
nor U7830 (N_7830,N_5192,N_3463);
nand U7831 (N_7831,N_5943,N_5135);
or U7832 (N_7832,N_5724,N_4583);
nand U7833 (N_7833,N_4287,N_3477);
nor U7834 (N_7834,N_5311,N_3622);
nand U7835 (N_7835,N_5860,N_4812);
or U7836 (N_7836,N_3459,N_3600);
and U7837 (N_7837,N_5561,N_3190);
or U7838 (N_7838,N_3562,N_3162);
nand U7839 (N_7839,N_5504,N_4378);
or U7840 (N_7840,N_3756,N_5487);
nand U7841 (N_7841,N_4884,N_3194);
nand U7842 (N_7842,N_5238,N_5075);
nor U7843 (N_7843,N_3293,N_5378);
nand U7844 (N_7844,N_5125,N_3726);
xnor U7845 (N_7845,N_4118,N_4351);
nand U7846 (N_7846,N_4096,N_3061);
nor U7847 (N_7847,N_4279,N_4626);
nor U7848 (N_7848,N_4694,N_5768);
nand U7849 (N_7849,N_3821,N_3778);
nand U7850 (N_7850,N_4475,N_5948);
or U7851 (N_7851,N_4370,N_5921);
nand U7852 (N_7852,N_3237,N_3637);
nor U7853 (N_7853,N_3302,N_4878);
and U7854 (N_7854,N_5029,N_5001);
or U7855 (N_7855,N_3057,N_4015);
or U7856 (N_7856,N_3106,N_4116);
nor U7857 (N_7857,N_4502,N_4196);
or U7858 (N_7858,N_3986,N_5361);
or U7859 (N_7859,N_5918,N_4466);
nor U7860 (N_7860,N_5530,N_5564);
nor U7861 (N_7861,N_5859,N_5009);
or U7862 (N_7862,N_5284,N_3156);
nor U7863 (N_7863,N_4232,N_5226);
or U7864 (N_7864,N_3147,N_3694);
nor U7865 (N_7865,N_3094,N_4933);
nor U7866 (N_7866,N_5440,N_3484);
nand U7867 (N_7867,N_3927,N_5499);
nand U7868 (N_7868,N_3314,N_4419);
nand U7869 (N_7869,N_4351,N_5750);
and U7870 (N_7870,N_3355,N_4279);
nor U7871 (N_7871,N_5516,N_4571);
and U7872 (N_7872,N_5577,N_5661);
or U7873 (N_7873,N_3963,N_5981);
nand U7874 (N_7874,N_3915,N_5162);
nand U7875 (N_7875,N_4695,N_4070);
nor U7876 (N_7876,N_3136,N_4594);
and U7877 (N_7877,N_3651,N_4168);
or U7878 (N_7878,N_5314,N_3314);
and U7879 (N_7879,N_4366,N_5674);
and U7880 (N_7880,N_3953,N_4152);
nand U7881 (N_7881,N_5470,N_5673);
nand U7882 (N_7882,N_4104,N_3131);
and U7883 (N_7883,N_4358,N_4422);
xor U7884 (N_7884,N_5893,N_5328);
or U7885 (N_7885,N_5745,N_5500);
or U7886 (N_7886,N_4809,N_4974);
or U7887 (N_7887,N_4880,N_3671);
nand U7888 (N_7888,N_5402,N_3609);
nand U7889 (N_7889,N_3916,N_3051);
nor U7890 (N_7890,N_3159,N_3811);
nand U7891 (N_7891,N_5059,N_3096);
xor U7892 (N_7892,N_5868,N_5314);
nor U7893 (N_7893,N_3534,N_4820);
nor U7894 (N_7894,N_4382,N_3539);
and U7895 (N_7895,N_3180,N_4782);
or U7896 (N_7896,N_3490,N_4582);
nand U7897 (N_7897,N_5247,N_4265);
and U7898 (N_7898,N_3148,N_3583);
and U7899 (N_7899,N_3921,N_4709);
and U7900 (N_7900,N_5848,N_4807);
or U7901 (N_7901,N_4645,N_4048);
and U7902 (N_7902,N_5661,N_4665);
nor U7903 (N_7903,N_4675,N_5909);
or U7904 (N_7904,N_3049,N_4172);
nand U7905 (N_7905,N_4234,N_4029);
nand U7906 (N_7906,N_4247,N_5147);
nor U7907 (N_7907,N_3691,N_4459);
or U7908 (N_7908,N_4234,N_3102);
nand U7909 (N_7909,N_4911,N_3547);
nand U7910 (N_7910,N_3549,N_5837);
and U7911 (N_7911,N_4703,N_4371);
nand U7912 (N_7912,N_3651,N_4262);
and U7913 (N_7913,N_3085,N_4596);
or U7914 (N_7914,N_4282,N_5630);
xnor U7915 (N_7915,N_5924,N_5444);
nand U7916 (N_7916,N_4272,N_3489);
or U7917 (N_7917,N_4165,N_4209);
nand U7918 (N_7918,N_4493,N_5247);
and U7919 (N_7919,N_4668,N_5354);
nor U7920 (N_7920,N_3216,N_5245);
nor U7921 (N_7921,N_3120,N_5628);
nand U7922 (N_7922,N_3557,N_5457);
nand U7923 (N_7923,N_4993,N_4001);
and U7924 (N_7924,N_4604,N_5765);
or U7925 (N_7925,N_4821,N_5094);
nand U7926 (N_7926,N_3778,N_4484);
nand U7927 (N_7927,N_3107,N_3726);
or U7928 (N_7928,N_3123,N_3048);
nor U7929 (N_7929,N_3010,N_5118);
and U7930 (N_7930,N_3666,N_3902);
nand U7931 (N_7931,N_5293,N_5393);
or U7932 (N_7932,N_5403,N_5966);
and U7933 (N_7933,N_4672,N_4958);
nand U7934 (N_7934,N_5592,N_4200);
nand U7935 (N_7935,N_4965,N_5277);
or U7936 (N_7936,N_3539,N_5230);
nor U7937 (N_7937,N_5385,N_4518);
and U7938 (N_7938,N_4795,N_4183);
or U7939 (N_7939,N_4439,N_3139);
or U7940 (N_7940,N_4311,N_5722);
nand U7941 (N_7941,N_4550,N_4299);
nand U7942 (N_7942,N_3624,N_5595);
nand U7943 (N_7943,N_5084,N_3801);
nand U7944 (N_7944,N_3343,N_4979);
or U7945 (N_7945,N_4163,N_3614);
or U7946 (N_7946,N_5513,N_5193);
nand U7947 (N_7947,N_5191,N_3460);
and U7948 (N_7948,N_3086,N_5253);
nor U7949 (N_7949,N_4147,N_5024);
or U7950 (N_7950,N_4191,N_5794);
nand U7951 (N_7951,N_5820,N_3611);
nor U7952 (N_7952,N_4713,N_4768);
nand U7953 (N_7953,N_5197,N_4685);
or U7954 (N_7954,N_5633,N_5645);
or U7955 (N_7955,N_5984,N_5060);
or U7956 (N_7956,N_5672,N_5217);
nor U7957 (N_7957,N_5584,N_3280);
nor U7958 (N_7958,N_3828,N_4784);
or U7959 (N_7959,N_5085,N_3490);
or U7960 (N_7960,N_4013,N_5501);
nand U7961 (N_7961,N_4856,N_4815);
or U7962 (N_7962,N_4230,N_5344);
nor U7963 (N_7963,N_3196,N_3758);
or U7964 (N_7964,N_3287,N_3488);
nand U7965 (N_7965,N_4073,N_5540);
or U7966 (N_7966,N_3688,N_5817);
nor U7967 (N_7967,N_4617,N_5891);
and U7968 (N_7968,N_3699,N_4029);
or U7969 (N_7969,N_3942,N_4860);
or U7970 (N_7970,N_3993,N_3983);
nor U7971 (N_7971,N_4020,N_5009);
or U7972 (N_7972,N_4194,N_3387);
nor U7973 (N_7973,N_3272,N_5785);
nor U7974 (N_7974,N_3475,N_5349);
and U7975 (N_7975,N_3880,N_5977);
or U7976 (N_7976,N_3690,N_5029);
nor U7977 (N_7977,N_5317,N_4440);
nand U7978 (N_7978,N_4923,N_3669);
and U7979 (N_7979,N_4183,N_3954);
or U7980 (N_7980,N_4462,N_3222);
nand U7981 (N_7981,N_3272,N_4743);
or U7982 (N_7982,N_5029,N_4697);
nor U7983 (N_7983,N_3090,N_5718);
nand U7984 (N_7984,N_4747,N_3426);
and U7985 (N_7985,N_3128,N_4826);
nand U7986 (N_7986,N_5055,N_4011);
nor U7987 (N_7987,N_5959,N_3149);
or U7988 (N_7988,N_5855,N_5599);
and U7989 (N_7989,N_3079,N_3270);
and U7990 (N_7990,N_5532,N_5918);
or U7991 (N_7991,N_5144,N_4978);
nand U7992 (N_7992,N_4245,N_3137);
and U7993 (N_7993,N_3480,N_5068);
or U7994 (N_7994,N_3940,N_4132);
nand U7995 (N_7995,N_3508,N_5866);
nor U7996 (N_7996,N_5724,N_4787);
nand U7997 (N_7997,N_4780,N_5992);
nand U7998 (N_7998,N_4060,N_3643);
and U7999 (N_7999,N_5088,N_4224);
nand U8000 (N_8000,N_4240,N_5895);
and U8001 (N_8001,N_3488,N_5427);
and U8002 (N_8002,N_3644,N_4200);
or U8003 (N_8003,N_4193,N_4599);
nor U8004 (N_8004,N_5664,N_5297);
and U8005 (N_8005,N_4965,N_3685);
nand U8006 (N_8006,N_4219,N_3612);
or U8007 (N_8007,N_5300,N_3988);
nor U8008 (N_8008,N_5984,N_4602);
nand U8009 (N_8009,N_5523,N_4409);
nand U8010 (N_8010,N_5389,N_4882);
nand U8011 (N_8011,N_4077,N_3476);
or U8012 (N_8012,N_4922,N_3435);
xor U8013 (N_8013,N_3643,N_3990);
nand U8014 (N_8014,N_5822,N_5387);
nor U8015 (N_8015,N_5224,N_4355);
nor U8016 (N_8016,N_5876,N_5163);
or U8017 (N_8017,N_3300,N_5030);
nand U8018 (N_8018,N_4108,N_5259);
and U8019 (N_8019,N_4306,N_5079);
nand U8020 (N_8020,N_3490,N_3129);
or U8021 (N_8021,N_3512,N_3238);
nand U8022 (N_8022,N_3122,N_5171);
and U8023 (N_8023,N_4254,N_3151);
or U8024 (N_8024,N_4494,N_4136);
nor U8025 (N_8025,N_5936,N_3762);
and U8026 (N_8026,N_3978,N_5709);
and U8027 (N_8027,N_4958,N_3458);
nand U8028 (N_8028,N_4996,N_4548);
nand U8029 (N_8029,N_5631,N_5374);
nor U8030 (N_8030,N_3917,N_4137);
nand U8031 (N_8031,N_3967,N_4923);
nand U8032 (N_8032,N_3298,N_3087);
and U8033 (N_8033,N_4484,N_3571);
or U8034 (N_8034,N_5938,N_5453);
xor U8035 (N_8035,N_5353,N_3326);
nor U8036 (N_8036,N_3196,N_5043);
or U8037 (N_8037,N_4231,N_4894);
and U8038 (N_8038,N_3401,N_4401);
and U8039 (N_8039,N_4392,N_5331);
or U8040 (N_8040,N_4768,N_4532);
and U8041 (N_8041,N_4020,N_3648);
and U8042 (N_8042,N_4468,N_3231);
or U8043 (N_8043,N_4406,N_3660);
nor U8044 (N_8044,N_3927,N_4214);
and U8045 (N_8045,N_5507,N_5076);
nor U8046 (N_8046,N_4970,N_3757);
nor U8047 (N_8047,N_4461,N_4447);
and U8048 (N_8048,N_5493,N_4707);
and U8049 (N_8049,N_3597,N_5087);
nor U8050 (N_8050,N_4430,N_5845);
nor U8051 (N_8051,N_5689,N_4854);
and U8052 (N_8052,N_5135,N_4053);
and U8053 (N_8053,N_4376,N_5619);
nand U8054 (N_8054,N_4336,N_5354);
nor U8055 (N_8055,N_5890,N_3070);
and U8056 (N_8056,N_3857,N_4757);
or U8057 (N_8057,N_5093,N_3737);
nor U8058 (N_8058,N_4781,N_3693);
nor U8059 (N_8059,N_4414,N_4945);
or U8060 (N_8060,N_3671,N_4789);
nor U8061 (N_8061,N_4726,N_3979);
and U8062 (N_8062,N_5154,N_4130);
nor U8063 (N_8063,N_5266,N_3197);
nor U8064 (N_8064,N_3122,N_4357);
and U8065 (N_8065,N_4878,N_3335);
nor U8066 (N_8066,N_4396,N_5614);
nor U8067 (N_8067,N_5340,N_3686);
or U8068 (N_8068,N_5285,N_3915);
and U8069 (N_8069,N_3254,N_3565);
nand U8070 (N_8070,N_5465,N_5096);
and U8071 (N_8071,N_4279,N_3859);
and U8072 (N_8072,N_5337,N_4124);
nor U8073 (N_8073,N_3090,N_4292);
and U8074 (N_8074,N_5994,N_4357);
and U8075 (N_8075,N_5703,N_3284);
nor U8076 (N_8076,N_5972,N_4871);
or U8077 (N_8077,N_3278,N_3783);
nand U8078 (N_8078,N_4139,N_4735);
nor U8079 (N_8079,N_5066,N_3330);
nor U8080 (N_8080,N_3421,N_5394);
nand U8081 (N_8081,N_4082,N_4944);
nor U8082 (N_8082,N_4910,N_5980);
nand U8083 (N_8083,N_4273,N_4776);
and U8084 (N_8084,N_5694,N_3316);
and U8085 (N_8085,N_5614,N_3110);
nor U8086 (N_8086,N_3106,N_5035);
nand U8087 (N_8087,N_5969,N_5676);
nand U8088 (N_8088,N_4797,N_5962);
or U8089 (N_8089,N_4886,N_3713);
nor U8090 (N_8090,N_4818,N_4173);
and U8091 (N_8091,N_5906,N_3389);
nand U8092 (N_8092,N_4128,N_4003);
nand U8093 (N_8093,N_4841,N_3078);
nor U8094 (N_8094,N_5275,N_4565);
nand U8095 (N_8095,N_4715,N_3619);
or U8096 (N_8096,N_4046,N_3187);
or U8097 (N_8097,N_3173,N_5138);
nand U8098 (N_8098,N_4072,N_3510);
and U8099 (N_8099,N_3391,N_3625);
nor U8100 (N_8100,N_4772,N_4511);
nand U8101 (N_8101,N_3521,N_5285);
nor U8102 (N_8102,N_3573,N_3508);
nand U8103 (N_8103,N_3068,N_3991);
nand U8104 (N_8104,N_3460,N_3177);
nand U8105 (N_8105,N_5001,N_3337);
and U8106 (N_8106,N_4292,N_5596);
nor U8107 (N_8107,N_3971,N_3299);
nand U8108 (N_8108,N_4556,N_5854);
or U8109 (N_8109,N_3821,N_3631);
or U8110 (N_8110,N_4605,N_4335);
nand U8111 (N_8111,N_5986,N_4212);
xor U8112 (N_8112,N_4458,N_3335);
or U8113 (N_8113,N_5640,N_4101);
or U8114 (N_8114,N_3660,N_4959);
nand U8115 (N_8115,N_5693,N_3597);
and U8116 (N_8116,N_4109,N_3045);
or U8117 (N_8117,N_5493,N_3712);
nor U8118 (N_8118,N_3852,N_4030);
nor U8119 (N_8119,N_4094,N_3918);
or U8120 (N_8120,N_5850,N_5003);
nand U8121 (N_8121,N_4055,N_3024);
nand U8122 (N_8122,N_4594,N_5754);
or U8123 (N_8123,N_4219,N_3349);
or U8124 (N_8124,N_4764,N_4266);
and U8125 (N_8125,N_4390,N_5870);
nor U8126 (N_8126,N_4445,N_4126);
and U8127 (N_8127,N_4920,N_5773);
or U8128 (N_8128,N_5394,N_5663);
nor U8129 (N_8129,N_3070,N_4126);
and U8130 (N_8130,N_5787,N_4844);
nor U8131 (N_8131,N_5775,N_4009);
and U8132 (N_8132,N_4715,N_3884);
and U8133 (N_8133,N_5939,N_5150);
nand U8134 (N_8134,N_4133,N_4599);
nor U8135 (N_8135,N_3309,N_5224);
and U8136 (N_8136,N_4666,N_5215);
nand U8137 (N_8137,N_4456,N_4118);
and U8138 (N_8138,N_4242,N_5428);
or U8139 (N_8139,N_3507,N_5679);
nand U8140 (N_8140,N_3013,N_3906);
or U8141 (N_8141,N_4567,N_3948);
nor U8142 (N_8142,N_5512,N_3780);
nor U8143 (N_8143,N_3115,N_3471);
nand U8144 (N_8144,N_5974,N_3235);
nand U8145 (N_8145,N_4161,N_4780);
or U8146 (N_8146,N_3083,N_3021);
nand U8147 (N_8147,N_5541,N_4930);
nor U8148 (N_8148,N_3493,N_3134);
and U8149 (N_8149,N_4351,N_3513);
or U8150 (N_8150,N_3260,N_4422);
nor U8151 (N_8151,N_3832,N_5654);
and U8152 (N_8152,N_3831,N_4176);
or U8153 (N_8153,N_3800,N_4907);
or U8154 (N_8154,N_3133,N_5625);
nand U8155 (N_8155,N_5928,N_3548);
and U8156 (N_8156,N_4919,N_5546);
or U8157 (N_8157,N_5647,N_4976);
nand U8158 (N_8158,N_4732,N_5049);
xnor U8159 (N_8159,N_4768,N_4114);
or U8160 (N_8160,N_4878,N_5886);
or U8161 (N_8161,N_5494,N_5285);
nor U8162 (N_8162,N_3556,N_3509);
nor U8163 (N_8163,N_5619,N_5593);
or U8164 (N_8164,N_4132,N_3689);
nor U8165 (N_8165,N_4994,N_4667);
nor U8166 (N_8166,N_3466,N_4416);
nor U8167 (N_8167,N_5390,N_4348);
or U8168 (N_8168,N_5016,N_5380);
and U8169 (N_8169,N_5605,N_3961);
and U8170 (N_8170,N_3030,N_3950);
or U8171 (N_8171,N_5285,N_5236);
and U8172 (N_8172,N_4339,N_5184);
or U8173 (N_8173,N_4835,N_5781);
or U8174 (N_8174,N_5116,N_5632);
nor U8175 (N_8175,N_3280,N_5925);
nor U8176 (N_8176,N_3288,N_3505);
nor U8177 (N_8177,N_3417,N_4766);
or U8178 (N_8178,N_5214,N_3119);
or U8179 (N_8179,N_3603,N_4535);
nand U8180 (N_8180,N_5941,N_3361);
nand U8181 (N_8181,N_5920,N_5875);
nand U8182 (N_8182,N_3728,N_3897);
nor U8183 (N_8183,N_5487,N_4992);
and U8184 (N_8184,N_3123,N_5173);
or U8185 (N_8185,N_5977,N_4111);
nand U8186 (N_8186,N_4804,N_3414);
and U8187 (N_8187,N_4956,N_5170);
and U8188 (N_8188,N_4726,N_5223);
nor U8189 (N_8189,N_4255,N_4638);
nor U8190 (N_8190,N_3825,N_4337);
nor U8191 (N_8191,N_5276,N_3223);
nand U8192 (N_8192,N_5984,N_4847);
or U8193 (N_8193,N_4022,N_3862);
nand U8194 (N_8194,N_3709,N_5913);
nand U8195 (N_8195,N_3670,N_4821);
or U8196 (N_8196,N_5225,N_5206);
nand U8197 (N_8197,N_3116,N_3642);
nor U8198 (N_8198,N_5490,N_3907);
or U8199 (N_8199,N_4621,N_3277);
and U8200 (N_8200,N_5734,N_5934);
and U8201 (N_8201,N_4442,N_5408);
or U8202 (N_8202,N_3961,N_3900);
nor U8203 (N_8203,N_4732,N_4942);
and U8204 (N_8204,N_3790,N_4393);
nand U8205 (N_8205,N_3121,N_5635);
or U8206 (N_8206,N_3461,N_4128);
nand U8207 (N_8207,N_3422,N_3284);
and U8208 (N_8208,N_4668,N_5964);
nor U8209 (N_8209,N_4129,N_4402);
nor U8210 (N_8210,N_5708,N_3374);
nand U8211 (N_8211,N_3322,N_4033);
nor U8212 (N_8212,N_3906,N_4361);
or U8213 (N_8213,N_5757,N_4312);
nor U8214 (N_8214,N_4344,N_4687);
nor U8215 (N_8215,N_3268,N_3110);
or U8216 (N_8216,N_5430,N_4450);
xnor U8217 (N_8217,N_5724,N_5097);
nor U8218 (N_8218,N_4049,N_3028);
nand U8219 (N_8219,N_3355,N_3113);
and U8220 (N_8220,N_3001,N_4517);
and U8221 (N_8221,N_3301,N_4376);
or U8222 (N_8222,N_5479,N_4222);
nor U8223 (N_8223,N_3313,N_5296);
nand U8224 (N_8224,N_5187,N_5899);
and U8225 (N_8225,N_4688,N_4815);
nor U8226 (N_8226,N_4407,N_3953);
and U8227 (N_8227,N_4892,N_5152);
nand U8228 (N_8228,N_4163,N_3936);
nor U8229 (N_8229,N_4023,N_4006);
nor U8230 (N_8230,N_3663,N_4441);
or U8231 (N_8231,N_3698,N_3483);
nor U8232 (N_8232,N_4198,N_3943);
and U8233 (N_8233,N_4423,N_5896);
nor U8234 (N_8234,N_5750,N_4996);
and U8235 (N_8235,N_3881,N_4883);
nand U8236 (N_8236,N_5164,N_4436);
and U8237 (N_8237,N_4911,N_4184);
and U8238 (N_8238,N_5872,N_4748);
or U8239 (N_8239,N_4382,N_3384);
and U8240 (N_8240,N_3065,N_4088);
nor U8241 (N_8241,N_3188,N_4973);
nor U8242 (N_8242,N_5839,N_3181);
xor U8243 (N_8243,N_4076,N_5206);
or U8244 (N_8244,N_3503,N_5295);
nand U8245 (N_8245,N_3260,N_5067);
nor U8246 (N_8246,N_3324,N_3744);
nand U8247 (N_8247,N_4753,N_3722);
and U8248 (N_8248,N_3498,N_5015);
and U8249 (N_8249,N_5068,N_4957);
nor U8250 (N_8250,N_4377,N_5390);
nand U8251 (N_8251,N_3147,N_5536);
and U8252 (N_8252,N_3108,N_5884);
nor U8253 (N_8253,N_5275,N_4378);
nand U8254 (N_8254,N_3063,N_3401);
or U8255 (N_8255,N_4067,N_4057);
nor U8256 (N_8256,N_5296,N_5598);
nand U8257 (N_8257,N_3098,N_3759);
and U8258 (N_8258,N_4754,N_3951);
and U8259 (N_8259,N_4247,N_4262);
and U8260 (N_8260,N_5093,N_5702);
or U8261 (N_8261,N_3650,N_3301);
nor U8262 (N_8262,N_5746,N_4367);
and U8263 (N_8263,N_3385,N_4250);
nand U8264 (N_8264,N_3441,N_4236);
nand U8265 (N_8265,N_3064,N_5458);
nand U8266 (N_8266,N_3066,N_4421);
nor U8267 (N_8267,N_5784,N_4133);
nand U8268 (N_8268,N_3929,N_4065);
and U8269 (N_8269,N_4686,N_5157);
or U8270 (N_8270,N_3222,N_3036);
or U8271 (N_8271,N_4556,N_4758);
nor U8272 (N_8272,N_3410,N_3127);
nand U8273 (N_8273,N_3919,N_4726);
and U8274 (N_8274,N_3091,N_5560);
nor U8275 (N_8275,N_5473,N_3420);
and U8276 (N_8276,N_5422,N_4416);
nand U8277 (N_8277,N_3623,N_3108);
and U8278 (N_8278,N_5575,N_4782);
and U8279 (N_8279,N_5307,N_3871);
and U8280 (N_8280,N_5114,N_4993);
and U8281 (N_8281,N_5475,N_4957);
nand U8282 (N_8282,N_4463,N_5076);
and U8283 (N_8283,N_5283,N_3118);
nor U8284 (N_8284,N_5933,N_5822);
nand U8285 (N_8285,N_4954,N_3484);
nor U8286 (N_8286,N_4457,N_4289);
nor U8287 (N_8287,N_5274,N_3779);
nor U8288 (N_8288,N_3796,N_5082);
and U8289 (N_8289,N_5523,N_3781);
or U8290 (N_8290,N_3568,N_5019);
or U8291 (N_8291,N_4001,N_3434);
or U8292 (N_8292,N_4568,N_5772);
nand U8293 (N_8293,N_4043,N_4162);
nand U8294 (N_8294,N_4864,N_5576);
or U8295 (N_8295,N_5218,N_5358);
nand U8296 (N_8296,N_5266,N_3582);
nor U8297 (N_8297,N_3166,N_4160);
and U8298 (N_8298,N_4210,N_5868);
nor U8299 (N_8299,N_4733,N_3256);
nand U8300 (N_8300,N_5859,N_5018);
or U8301 (N_8301,N_4866,N_3004);
nand U8302 (N_8302,N_5202,N_5605);
or U8303 (N_8303,N_3841,N_3060);
and U8304 (N_8304,N_5249,N_3751);
or U8305 (N_8305,N_3371,N_4675);
or U8306 (N_8306,N_4427,N_4587);
and U8307 (N_8307,N_5183,N_3986);
nand U8308 (N_8308,N_5130,N_3059);
nand U8309 (N_8309,N_5232,N_4849);
and U8310 (N_8310,N_5915,N_5759);
nor U8311 (N_8311,N_3977,N_3097);
nand U8312 (N_8312,N_5892,N_4501);
nand U8313 (N_8313,N_3767,N_4330);
nand U8314 (N_8314,N_4765,N_4075);
nand U8315 (N_8315,N_4309,N_5104);
nor U8316 (N_8316,N_5124,N_5708);
nand U8317 (N_8317,N_3745,N_5024);
nand U8318 (N_8318,N_4686,N_3742);
or U8319 (N_8319,N_5187,N_3998);
nor U8320 (N_8320,N_5443,N_4674);
and U8321 (N_8321,N_4526,N_3812);
and U8322 (N_8322,N_3242,N_5276);
nor U8323 (N_8323,N_4398,N_4483);
nor U8324 (N_8324,N_3719,N_5000);
and U8325 (N_8325,N_3608,N_5558);
and U8326 (N_8326,N_5512,N_5901);
nor U8327 (N_8327,N_4738,N_5967);
or U8328 (N_8328,N_3040,N_5760);
nand U8329 (N_8329,N_3557,N_4873);
nor U8330 (N_8330,N_4294,N_5353);
and U8331 (N_8331,N_4277,N_3882);
and U8332 (N_8332,N_3344,N_4328);
or U8333 (N_8333,N_4722,N_4310);
or U8334 (N_8334,N_5382,N_5311);
nand U8335 (N_8335,N_5929,N_4169);
or U8336 (N_8336,N_4092,N_3612);
and U8337 (N_8337,N_4694,N_4670);
nor U8338 (N_8338,N_3628,N_5486);
or U8339 (N_8339,N_5726,N_4374);
nand U8340 (N_8340,N_4762,N_3706);
or U8341 (N_8341,N_4529,N_3445);
and U8342 (N_8342,N_4433,N_5558);
nand U8343 (N_8343,N_3859,N_3077);
and U8344 (N_8344,N_4611,N_5764);
nand U8345 (N_8345,N_4976,N_4352);
nand U8346 (N_8346,N_3638,N_5016);
nor U8347 (N_8347,N_5217,N_5774);
nand U8348 (N_8348,N_4117,N_3659);
nor U8349 (N_8349,N_5933,N_4667);
nor U8350 (N_8350,N_3460,N_4754);
nor U8351 (N_8351,N_4546,N_4242);
nand U8352 (N_8352,N_4773,N_4352);
or U8353 (N_8353,N_4710,N_3750);
and U8354 (N_8354,N_4563,N_4080);
or U8355 (N_8355,N_5300,N_3366);
nor U8356 (N_8356,N_4524,N_5260);
and U8357 (N_8357,N_5617,N_5235);
and U8358 (N_8358,N_3459,N_3210);
nor U8359 (N_8359,N_3668,N_4218);
or U8360 (N_8360,N_3950,N_4287);
and U8361 (N_8361,N_5856,N_4610);
and U8362 (N_8362,N_3682,N_5279);
or U8363 (N_8363,N_3519,N_5497);
nor U8364 (N_8364,N_5946,N_5067);
and U8365 (N_8365,N_4239,N_4875);
and U8366 (N_8366,N_3631,N_3294);
nand U8367 (N_8367,N_3154,N_3958);
and U8368 (N_8368,N_5785,N_3022);
nand U8369 (N_8369,N_4828,N_4314);
and U8370 (N_8370,N_3358,N_3617);
and U8371 (N_8371,N_4384,N_3980);
nand U8372 (N_8372,N_3599,N_3242);
or U8373 (N_8373,N_3391,N_4051);
or U8374 (N_8374,N_3684,N_5630);
nand U8375 (N_8375,N_5313,N_4539);
or U8376 (N_8376,N_3900,N_4668);
nor U8377 (N_8377,N_5705,N_5006);
nor U8378 (N_8378,N_3346,N_5405);
nand U8379 (N_8379,N_4515,N_4514);
or U8380 (N_8380,N_4255,N_5495);
and U8381 (N_8381,N_3433,N_4485);
nand U8382 (N_8382,N_4547,N_4463);
nor U8383 (N_8383,N_3474,N_5635);
and U8384 (N_8384,N_4178,N_5443);
and U8385 (N_8385,N_3584,N_3611);
or U8386 (N_8386,N_4582,N_5352);
nor U8387 (N_8387,N_4186,N_5166);
nand U8388 (N_8388,N_3873,N_3715);
or U8389 (N_8389,N_3136,N_4217);
nor U8390 (N_8390,N_5741,N_5935);
nor U8391 (N_8391,N_5589,N_3684);
nand U8392 (N_8392,N_3569,N_4103);
and U8393 (N_8393,N_3512,N_3063);
nand U8394 (N_8394,N_4037,N_5268);
nor U8395 (N_8395,N_4204,N_4501);
nand U8396 (N_8396,N_5087,N_5431);
or U8397 (N_8397,N_4435,N_3730);
nand U8398 (N_8398,N_4093,N_3671);
and U8399 (N_8399,N_3304,N_5758);
and U8400 (N_8400,N_4300,N_3996);
nor U8401 (N_8401,N_3793,N_4846);
nor U8402 (N_8402,N_4696,N_5080);
and U8403 (N_8403,N_4426,N_5540);
nor U8404 (N_8404,N_3082,N_4461);
nor U8405 (N_8405,N_3902,N_5877);
nor U8406 (N_8406,N_3146,N_3363);
or U8407 (N_8407,N_4383,N_4745);
nand U8408 (N_8408,N_3308,N_4215);
nand U8409 (N_8409,N_5322,N_4934);
nand U8410 (N_8410,N_5982,N_5989);
nor U8411 (N_8411,N_4504,N_4631);
xnor U8412 (N_8412,N_3822,N_5602);
and U8413 (N_8413,N_4665,N_4709);
or U8414 (N_8414,N_4706,N_5038);
nand U8415 (N_8415,N_4750,N_5385);
and U8416 (N_8416,N_4579,N_3263);
and U8417 (N_8417,N_3613,N_5873);
and U8418 (N_8418,N_3262,N_4774);
or U8419 (N_8419,N_5058,N_5105);
or U8420 (N_8420,N_5661,N_3467);
nand U8421 (N_8421,N_4890,N_3914);
nor U8422 (N_8422,N_3158,N_5159);
or U8423 (N_8423,N_4432,N_3779);
and U8424 (N_8424,N_3024,N_5411);
nor U8425 (N_8425,N_5434,N_5081);
nand U8426 (N_8426,N_3216,N_4187);
or U8427 (N_8427,N_4230,N_3234);
and U8428 (N_8428,N_4633,N_3412);
or U8429 (N_8429,N_5604,N_4950);
or U8430 (N_8430,N_4303,N_4705);
and U8431 (N_8431,N_4608,N_4999);
and U8432 (N_8432,N_5393,N_5574);
nor U8433 (N_8433,N_5391,N_5789);
or U8434 (N_8434,N_3973,N_3719);
or U8435 (N_8435,N_3326,N_4920);
nor U8436 (N_8436,N_4636,N_4439);
or U8437 (N_8437,N_3534,N_5931);
or U8438 (N_8438,N_3513,N_5777);
nand U8439 (N_8439,N_3950,N_5328);
and U8440 (N_8440,N_4628,N_5046);
or U8441 (N_8441,N_4485,N_3277);
and U8442 (N_8442,N_5010,N_3301);
nand U8443 (N_8443,N_3410,N_3719);
and U8444 (N_8444,N_5741,N_3607);
or U8445 (N_8445,N_5099,N_4171);
nor U8446 (N_8446,N_3959,N_3228);
or U8447 (N_8447,N_5032,N_5732);
nor U8448 (N_8448,N_4996,N_3872);
nand U8449 (N_8449,N_3921,N_5063);
nor U8450 (N_8450,N_5428,N_4663);
nand U8451 (N_8451,N_3728,N_5377);
or U8452 (N_8452,N_5141,N_5329);
and U8453 (N_8453,N_5035,N_3766);
and U8454 (N_8454,N_4597,N_4461);
nor U8455 (N_8455,N_4436,N_3525);
or U8456 (N_8456,N_3549,N_4815);
nor U8457 (N_8457,N_4997,N_3246);
or U8458 (N_8458,N_3226,N_4647);
or U8459 (N_8459,N_3405,N_5914);
nand U8460 (N_8460,N_5868,N_3675);
or U8461 (N_8461,N_4198,N_5155);
or U8462 (N_8462,N_4681,N_3176);
or U8463 (N_8463,N_5008,N_3208);
and U8464 (N_8464,N_3667,N_4904);
nand U8465 (N_8465,N_5583,N_4142);
nand U8466 (N_8466,N_5389,N_3503);
or U8467 (N_8467,N_3929,N_5379);
nor U8468 (N_8468,N_4631,N_3206);
nand U8469 (N_8469,N_5142,N_4833);
or U8470 (N_8470,N_4282,N_4668);
xnor U8471 (N_8471,N_4416,N_4624);
and U8472 (N_8472,N_5829,N_4117);
nand U8473 (N_8473,N_4827,N_4490);
and U8474 (N_8474,N_4762,N_4888);
or U8475 (N_8475,N_4580,N_5513);
nor U8476 (N_8476,N_5284,N_3142);
and U8477 (N_8477,N_3059,N_4051);
nor U8478 (N_8478,N_4495,N_4404);
or U8479 (N_8479,N_4233,N_3300);
or U8480 (N_8480,N_4150,N_4544);
nand U8481 (N_8481,N_4038,N_5446);
xor U8482 (N_8482,N_3368,N_4347);
nor U8483 (N_8483,N_3896,N_4111);
or U8484 (N_8484,N_4260,N_5678);
or U8485 (N_8485,N_5332,N_5631);
and U8486 (N_8486,N_3277,N_5662);
nand U8487 (N_8487,N_3209,N_3336);
or U8488 (N_8488,N_3911,N_5491);
xor U8489 (N_8489,N_5109,N_5685);
xnor U8490 (N_8490,N_5479,N_4707);
or U8491 (N_8491,N_3118,N_3936);
nand U8492 (N_8492,N_5749,N_5228);
nand U8493 (N_8493,N_5482,N_5352);
nand U8494 (N_8494,N_3844,N_5431);
nor U8495 (N_8495,N_4914,N_3156);
nor U8496 (N_8496,N_5721,N_5362);
nor U8497 (N_8497,N_4433,N_4240);
nand U8498 (N_8498,N_3829,N_3530);
or U8499 (N_8499,N_4545,N_4558);
nor U8500 (N_8500,N_4550,N_3016);
or U8501 (N_8501,N_4387,N_4185);
nand U8502 (N_8502,N_5318,N_4438);
nand U8503 (N_8503,N_4415,N_4252);
nand U8504 (N_8504,N_3485,N_5265);
nand U8505 (N_8505,N_4534,N_5947);
or U8506 (N_8506,N_5518,N_5820);
or U8507 (N_8507,N_3051,N_5362);
or U8508 (N_8508,N_3718,N_5608);
nor U8509 (N_8509,N_4206,N_5196);
nand U8510 (N_8510,N_4653,N_4713);
nand U8511 (N_8511,N_3632,N_5886);
or U8512 (N_8512,N_5369,N_5403);
nor U8513 (N_8513,N_4041,N_4182);
nand U8514 (N_8514,N_5856,N_5366);
nand U8515 (N_8515,N_5071,N_3984);
nor U8516 (N_8516,N_4816,N_5591);
nor U8517 (N_8517,N_5574,N_5668);
nand U8518 (N_8518,N_5319,N_4334);
nand U8519 (N_8519,N_3834,N_3027);
nor U8520 (N_8520,N_5089,N_5914);
nor U8521 (N_8521,N_5381,N_4690);
or U8522 (N_8522,N_3275,N_4180);
nand U8523 (N_8523,N_3935,N_4745);
nor U8524 (N_8524,N_5876,N_4420);
xnor U8525 (N_8525,N_4685,N_3344);
nand U8526 (N_8526,N_4049,N_3640);
or U8527 (N_8527,N_5384,N_3265);
nor U8528 (N_8528,N_4274,N_4964);
and U8529 (N_8529,N_3063,N_4397);
nor U8530 (N_8530,N_3129,N_3082);
nor U8531 (N_8531,N_4884,N_3754);
nor U8532 (N_8532,N_3727,N_3951);
nor U8533 (N_8533,N_3771,N_5464);
nand U8534 (N_8534,N_5114,N_3413);
nor U8535 (N_8535,N_5556,N_5215);
nor U8536 (N_8536,N_3929,N_5580);
nand U8537 (N_8537,N_3092,N_3510);
and U8538 (N_8538,N_5743,N_4620);
or U8539 (N_8539,N_5275,N_5518);
nor U8540 (N_8540,N_5311,N_4513);
nand U8541 (N_8541,N_4470,N_4607);
nand U8542 (N_8542,N_4992,N_3429);
nand U8543 (N_8543,N_3378,N_5315);
or U8544 (N_8544,N_5634,N_4339);
nor U8545 (N_8545,N_3215,N_4073);
or U8546 (N_8546,N_5549,N_3657);
nor U8547 (N_8547,N_5124,N_5298);
nand U8548 (N_8548,N_5519,N_5052);
nor U8549 (N_8549,N_4664,N_4692);
nand U8550 (N_8550,N_5755,N_5695);
or U8551 (N_8551,N_5482,N_5619);
nand U8552 (N_8552,N_3576,N_3533);
or U8553 (N_8553,N_5390,N_4496);
or U8554 (N_8554,N_3493,N_3983);
nor U8555 (N_8555,N_5508,N_3437);
nor U8556 (N_8556,N_3471,N_3333);
nor U8557 (N_8557,N_3380,N_4580);
or U8558 (N_8558,N_4141,N_5176);
and U8559 (N_8559,N_5676,N_5001);
nor U8560 (N_8560,N_3350,N_5824);
nor U8561 (N_8561,N_5786,N_5983);
or U8562 (N_8562,N_4968,N_3834);
and U8563 (N_8563,N_4366,N_3626);
and U8564 (N_8564,N_3135,N_4806);
nor U8565 (N_8565,N_5334,N_3013);
nand U8566 (N_8566,N_4102,N_5300);
nand U8567 (N_8567,N_5011,N_3945);
nand U8568 (N_8568,N_4108,N_3536);
or U8569 (N_8569,N_5457,N_5472);
nand U8570 (N_8570,N_5093,N_5574);
nand U8571 (N_8571,N_3816,N_5208);
nand U8572 (N_8572,N_4222,N_4826);
and U8573 (N_8573,N_5201,N_5809);
and U8574 (N_8574,N_4940,N_3090);
nand U8575 (N_8575,N_5408,N_5981);
nand U8576 (N_8576,N_4235,N_4947);
and U8577 (N_8577,N_3184,N_4618);
or U8578 (N_8578,N_4482,N_3229);
nor U8579 (N_8579,N_5111,N_5745);
and U8580 (N_8580,N_3417,N_5448);
and U8581 (N_8581,N_3540,N_5451);
nor U8582 (N_8582,N_5749,N_4810);
nand U8583 (N_8583,N_5139,N_4768);
nor U8584 (N_8584,N_5756,N_3933);
nand U8585 (N_8585,N_4950,N_5709);
nand U8586 (N_8586,N_5119,N_3412);
and U8587 (N_8587,N_5612,N_4489);
and U8588 (N_8588,N_5248,N_3181);
nand U8589 (N_8589,N_3496,N_3070);
and U8590 (N_8590,N_5796,N_3648);
nand U8591 (N_8591,N_3461,N_5599);
nand U8592 (N_8592,N_4155,N_3923);
and U8593 (N_8593,N_3461,N_3255);
and U8594 (N_8594,N_5265,N_5135);
and U8595 (N_8595,N_3467,N_4117);
and U8596 (N_8596,N_3616,N_3240);
or U8597 (N_8597,N_4695,N_4597);
nor U8598 (N_8598,N_3340,N_3569);
nor U8599 (N_8599,N_3658,N_5973);
or U8600 (N_8600,N_4428,N_5234);
nand U8601 (N_8601,N_3982,N_3748);
or U8602 (N_8602,N_5112,N_5756);
nor U8603 (N_8603,N_5935,N_5315);
and U8604 (N_8604,N_3360,N_4612);
nor U8605 (N_8605,N_3128,N_3325);
nand U8606 (N_8606,N_3445,N_4578);
and U8607 (N_8607,N_5136,N_4642);
nor U8608 (N_8608,N_5906,N_4810);
nor U8609 (N_8609,N_3311,N_5665);
nand U8610 (N_8610,N_5434,N_4300);
or U8611 (N_8611,N_4482,N_5539);
nand U8612 (N_8612,N_5756,N_3086);
nor U8613 (N_8613,N_5162,N_5575);
nand U8614 (N_8614,N_4108,N_5063);
or U8615 (N_8615,N_4484,N_5515);
or U8616 (N_8616,N_5622,N_3290);
or U8617 (N_8617,N_4572,N_3915);
or U8618 (N_8618,N_5805,N_4870);
nor U8619 (N_8619,N_5413,N_4020);
nand U8620 (N_8620,N_4275,N_3132);
or U8621 (N_8621,N_5093,N_3443);
nor U8622 (N_8622,N_4399,N_3071);
nor U8623 (N_8623,N_4491,N_3158);
xnor U8624 (N_8624,N_5858,N_4336);
nor U8625 (N_8625,N_3456,N_3030);
or U8626 (N_8626,N_5874,N_4868);
nand U8627 (N_8627,N_3653,N_3812);
nand U8628 (N_8628,N_4868,N_5241);
nand U8629 (N_8629,N_3908,N_4607);
nand U8630 (N_8630,N_3216,N_5471);
or U8631 (N_8631,N_4918,N_4666);
and U8632 (N_8632,N_5416,N_5547);
xor U8633 (N_8633,N_4113,N_3559);
nor U8634 (N_8634,N_5089,N_3438);
nand U8635 (N_8635,N_3070,N_4388);
or U8636 (N_8636,N_4701,N_4654);
nand U8637 (N_8637,N_3204,N_5385);
or U8638 (N_8638,N_3271,N_4948);
nor U8639 (N_8639,N_3693,N_3866);
and U8640 (N_8640,N_3442,N_5326);
and U8641 (N_8641,N_4422,N_5681);
nor U8642 (N_8642,N_4994,N_4765);
and U8643 (N_8643,N_5124,N_4580);
and U8644 (N_8644,N_3184,N_4600);
nand U8645 (N_8645,N_3452,N_5919);
or U8646 (N_8646,N_3802,N_3940);
and U8647 (N_8647,N_4436,N_5604);
or U8648 (N_8648,N_3694,N_5027);
nand U8649 (N_8649,N_5224,N_5003);
nand U8650 (N_8650,N_4342,N_3950);
or U8651 (N_8651,N_3214,N_4581);
or U8652 (N_8652,N_3119,N_5398);
and U8653 (N_8653,N_3864,N_4499);
nand U8654 (N_8654,N_3220,N_3450);
or U8655 (N_8655,N_5588,N_4753);
nand U8656 (N_8656,N_5377,N_5392);
nor U8657 (N_8657,N_4103,N_3052);
or U8658 (N_8658,N_4790,N_4780);
and U8659 (N_8659,N_5426,N_5619);
nand U8660 (N_8660,N_3339,N_4980);
and U8661 (N_8661,N_5701,N_3619);
nor U8662 (N_8662,N_3353,N_4714);
and U8663 (N_8663,N_4398,N_4896);
nand U8664 (N_8664,N_4102,N_5130);
nor U8665 (N_8665,N_4975,N_3745);
nor U8666 (N_8666,N_5393,N_5788);
nand U8667 (N_8667,N_4579,N_4606);
and U8668 (N_8668,N_4314,N_5971);
nand U8669 (N_8669,N_3946,N_5566);
nand U8670 (N_8670,N_3916,N_3065);
nor U8671 (N_8671,N_3827,N_5132);
and U8672 (N_8672,N_4577,N_3467);
and U8673 (N_8673,N_4053,N_5547);
and U8674 (N_8674,N_4973,N_4544);
nor U8675 (N_8675,N_5569,N_4111);
and U8676 (N_8676,N_5235,N_3301);
and U8677 (N_8677,N_4277,N_3857);
nor U8678 (N_8678,N_4623,N_5032);
or U8679 (N_8679,N_5291,N_3304);
or U8680 (N_8680,N_5163,N_3456);
and U8681 (N_8681,N_5978,N_3670);
and U8682 (N_8682,N_5990,N_4496);
nand U8683 (N_8683,N_3824,N_5499);
and U8684 (N_8684,N_4588,N_3354);
or U8685 (N_8685,N_3775,N_5537);
or U8686 (N_8686,N_4154,N_3157);
nor U8687 (N_8687,N_3981,N_4117);
and U8688 (N_8688,N_5300,N_5016);
nand U8689 (N_8689,N_4825,N_5408);
and U8690 (N_8690,N_3587,N_3128);
or U8691 (N_8691,N_4527,N_3292);
nand U8692 (N_8692,N_5353,N_4289);
nand U8693 (N_8693,N_4391,N_5981);
nand U8694 (N_8694,N_5967,N_5020);
nor U8695 (N_8695,N_3985,N_4924);
nor U8696 (N_8696,N_3726,N_4993);
nor U8697 (N_8697,N_3236,N_3103);
nor U8698 (N_8698,N_3349,N_3079);
and U8699 (N_8699,N_3661,N_4247);
or U8700 (N_8700,N_4996,N_3259);
or U8701 (N_8701,N_4775,N_3287);
and U8702 (N_8702,N_3204,N_4290);
nand U8703 (N_8703,N_5025,N_3289);
nand U8704 (N_8704,N_4753,N_4425);
nor U8705 (N_8705,N_4780,N_5289);
or U8706 (N_8706,N_5040,N_3038);
or U8707 (N_8707,N_5091,N_5900);
nor U8708 (N_8708,N_4680,N_5321);
and U8709 (N_8709,N_5039,N_5645);
and U8710 (N_8710,N_5174,N_3985);
or U8711 (N_8711,N_4787,N_4451);
nor U8712 (N_8712,N_5356,N_5854);
nor U8713 (N_8713,N_5554,N_5435);
or U8714 (N_8714,N_3115,N_3383);
xor U8715 (N_8715,N_3911,N_4815);
and U8716 (N_8716,N_4520,N_4949);
nor U8717 (N_8717,N_5371,N_4795);
or U8718 (N_8718,N_4377,N_3068);
or U8719 (N_8719,N_3068,N_5981);
and U8720 (N_8720,N_3356,N_5350);
and U8721 (N_8721,N_4405,N_4136);
and U8722 (N_8722,N_5188,N_5849);
or U8723 (N_8723,N_4796,N_5368);
nand U8724 (N_8724,N_4173,N_4470);
nand U8725 (N_8725,N_3062,N_5453);
or U8726 (N_8726,N_4083,N_3285);
and U8727 (N_8727,N_3072,N_5872);
and U8728 (N_8728,N_3703,N_4274);
and U8729 (N_8729,N_3391,N_5115);
and U8730 (N_8730,N_5127,N_4736);
nor U8731 (N_8731,N_4387,N_3931);
and U8732 (N_8732,N_3834,N_4230);
and U8733 (N_8733,N_3238,N_4345);
and U8734 (N_8734,N_5676,N_3270);
nand U8735 (N_8735,N_4446,N_5277);
nor U8736 (N_8736,N_3155,N_3761);
nor U8737 (N_8737,N_3685,N_4649);
or U8738 (N_8738,N_5046,N_4327);
nor U8739 (N_8739,N_4080,N_3649);
or U8740 (N_8740,N_3405,N_3684);
nand U8741 (N_8741,N_5200,N_3607);
nor U8742 (N_8742,N_4936,N_5255);
nand U8743 (N_8743,N_3103,N_5262);
nor U8744 (N_8744,N_4935,N_3751);
or U8745 (N_8745,N_3449,N_4548);
nor U8746 (N_8746,N_3111,N_4435);
nor U8747 (N_8747,N_5085,N_5009);
or U8748 (N_8748,N_4517,N_5610);
nor U8749 (N_8749,N_5939,N_5333);
and U8750 (N_8750,N_4085,N_5530);
and U8751 (N_8751,N_3833,N_4753);
nand U8752 (N_8752,N_5870,N_4869);
nand U8753 (N_8753,N_3611,N_5142);
or U8754 (N_8754,N_5211,N_4197);
or U8755 (N_8755,N_3168,N_5628);
nor U8756 (N_8756,N_4945,N_3459);
and U8757 (N_8757,N_4490,N_4130);
and U8758 (N_8758,N_5757,N_5394);
nand U8759 (N_8759,N_5367,N_5768);
nor U8760 (N_8760,N_5666,N_3786);
nor U8761 (N_8761,N_5867,N_3951);
nor U8762 (N_8762,N_5394,N_5932);
nand U8763 (N_8763,N_5965,N_3023);
nor U8764 (N_8764,N_5036,N_3804);
nor U8765 (N_8765,N_5449,N_4852);
nand U8766 (N_8766,N_4220,N_4142);
and U8767 (N_8767,N_5765,N_5863);
and U8768 (N_8768,N_3824,N_5788);
or U8769 (N_8769,N_3524,N_5241);
and U8770 (N_8770,N_3725,N_3826);
nor U8771 (N_8771,N_3182,N_4423);
or U8772 (N_8772,N_4665,N_4967);
nand U8773 (N_8773,N_5979,N_4722);
or U8774 (N_8774,N_3792,N_5395);
nand U8775 (N_8775,N_5295,N_5131);
or U8776 (N_8776,N_3960,N_4128);
nor U8777 (N_8777,N_4304,N_5298);
and U8778 (N_8778,N_4478,N_3522);
nor U8779 (N_8779,N_3045,N_3496);
nand U8780 (N_8780,N_3178,N_4972);
or U8781 (N_8781,N_3890,N_5718);
and U8782 (N_8782,N_4528,N_3771);
nand U8783 (N_8783,N_4513,N_4098);
nand U8784 (N_8784,N_5126,N_3210);
nand U8785 (N_8785,N_5145,N_5352);
nor U8786 (N_8786,N_4589,N_5705);
and U8787 (N_8787,N_3402,N_5453);
nand U8788 (N_8788,N_5656,N_5446);
nor U8789 (N_8789,N_4682,N_4192);
or U8790 (N_8790,N_4667,N_5141);
or U8791 (N_8791,N_4253,N_5237);
or U8792 (N_8792,N_5416,N_3883);
nand U8793 (N_8793,N_5658,N_5451);
and U8794 (N_8794,N_5371,N_5183);
or U8795 (N_8795,N_3508,N_3235);
or U8796 (N_8796,N_5199,N_3978);
and U8797 (N_8797,N_4706,N_3178);
and U8798 (N_8798,N_3323,N_3274);
and U8799 (N_8799,N_4620,N_5732);
nand U8800 (N_8800,N_4200,N_4342);
and U8801 (N_8801,N_3341,N_5337);
nor U8802 (N_8802,N_3316,N_3477);
nand U8803 (N_8803,N_5466,N_3037);
and U8804 (N_8804,N_4997,N_5669);
and U8805 (N_8805,N_4490,N_5816);
nand U8806 (N_8806,N_5215,N_4314);
and U8807 (N_8807,N_4707,N_5736);
and U8808 (N_8808,N_5900,N_4878);
nand U8809 (N_8809,N_4621,N_4751);
nor U8810 (N_8810,N_5982,N_5675);
nor U8811 (N_8811,N_3143,N_4114);
nor U8812 (N_8812,N_5507,N_5804);
or U8813 (N_8813,N_4745,N_3522);
nor U8814 (N_8814,N_3117,N_5280);
or U8815 (N_8815,N_4341,N_5010);
nand U8816 (N_8816,N_3064,N_4827);
or U8817 (N_8817,N_5565,N_5515);
or U8818 (N_8818,N_4762,N_5933);
and U8819 (N_8819,N_3709,N_3163);
nand U8820 (N_8820,N_4839,N_5309);
and U8821 (N_8821,N_3874,N_5441);
and U8822 (N_8822,N_3842,N_5771);
or U8823 (N_8823,N_3608,N_4995);
and U8824 (N_8824,N_5826,N_4340);
nor U8825 (N_8825,N_3518,N_5915);
and U8826 (N_8826,N_3078,N_3969);
nand U8827 (N_8827,N_4360,N_4625);
nand U8828 (N_8828,N_3823,N_5313);
nor U8829 (N_8829,N_5312,N_5901);
nand U8830 (N_8830,N_4852,N_3065);
nor U8831 (N_8831,N_3154,N_3074);
or U8832 (N_8832,N_4792,N_4840);
nand U8833 (N_8833,N_5864,N_3579);
nor U8834 (N_8834,N_5934,N_5814);
nand U8835 (N_8835,N_4520,N_5435);
or U8836 (N_8836,N_3799,N_3597);
or U8837 (N_8837,N_5730,N_5066);
or U8838 (N_8838,N_5301,N_3996);
nand U8839 (N_8839,N_5927,N_5653);
and U8840 (N_8840,N_5853,N_3633);
nor U8841 (N_8841,N_5508,N_5240);
or U8842 (N_8842,N_3973,N_5784);
or U8843 (N_8843,N_5260,N_5227);
nand U8844 (N_8844,N_3292,N_3749);
nand U8845 (N_8845,N_4160,N_5080);
or U8846 (N_8846,N_3806,N_3140);
or U8847 (N_8847,N_5047,N_5018);
or U8848 (N_8848,N_4956,N_5479);
and U8849 (N_8849,N_4216,N_5350);
and U8850 (N_8850,N_5821,N_4910);
and U8851 (N_8851,N_3504,N_5908);
or U8852 (N_8852,N_4224,N_5178);
or U8853 (N_8853,N_5391,N_3150);
nand U8854 (N_8854,N_3132,N_3941);
and U8855 (N_8855,N_5959,N_5886);
xnor U8856 (N_8856,N_5845,N_4791);
and U8857 (N_8857,N_4597,N_3604);
or U8858 (N_8858,N_4699,N_5654);
nor U8859 (N_8859,N_3153,N_4159);
nand U8860 (N_8860,N_3910,N_4710);
nand U8861 (N_8861,N_5614,N_5001);
nor U8862 (N_8862,N_3472,N_4859);
nor U8863 (N_8863,N_3305,N_4830);
and U8864 (N_8864,N_4427,N_3619);
nand U8865 (N_8865,N_5966,N_5212);
nor U8866 (N_8866,N_4661,N_5954);
nand U8867 (N_8867,N_3905,N_4599);
nor U8868 (N_8868,N_4427,N_4364);
nand U8869 (N_8869,N_3744,N_4719);
nor U8870 (N_8870,N_3775,N_3246);
or U8871 (N_8871,N_4852,N_5034);
nand U8872 (N_8872,N_3328,N_3198);
or U8873 (N_8873,N_5289,N_3453);
or U8874 (N_8874,N_5270,N_5356);
or U8875 (N_8875,N_5372,N_5277);
or U8876 (N_8876,N_5428,N_4177);
nand U8877 (N_8877,N_4719,N_5799);
or U8878 (N_8878,N_3553,N_4596);
nand U8879 (N_8879,N_4889,N_5028);
nor U8880 (N_8880,N_5574,N_4036);
and U8881 (N_8881,N_5254,N_3526);
nor U8882 (N_8882,N_5901,N_3880);
or U8883 (N_8883,N_5973,N_3655);
and U8884 (N_8884,N_4041,N_3976);
and U8885 (N_8885,N_5251,N_3815);
or U8886 (N_8886,N_4067,N_3140);
or U8887 (N_8887,N_4742,N_3762);
and U8888 (N_8888,N_3114,N_4060);
nor U8889 (N_8889,N_4550,N_5249);
or U8890 (N_8890,N_5222,N_4891);
or U8891 (N_8891,N_5613,N_4337);
nand U8892 (N_8892,N_3962,N_3762);
nor U8893 (N_8893,N_4482,N_5730);
nor U8894 (N_8894,N_4479,N_5825);
nor U8895 (N_8895,N_4723,N_4278);
nor U8896 (N_8896,N_5133,N_3773);
and U8897 (N_8897,N_3330,N_3349);
or U8898 (N_8898,N_5952,N_4822);
and U8899 (N_8899,N_4453,N_4603);
nor U8900 (N_8900,N_5632,N_4685);
or U8901 (N_8901,N_3979,N_4601);
or U8902 (N_8902,N_5746,N_4007);
and U8903 (N_8903,N_4070,N_5049);
nand U8904 (N_8904,N_5673,N_3856);
nand U8905 (N_8905,N_4654,N_5653);
nor U8906 (N_8906,N_3113,N_5129);
nand U8907 (N_8907,N_5684,N_5170);
nor U8908 (N_8908,N_5788,N_3823);
nor U8909 (N_8909,N_3617,N_3969);
nor U8910 (N_8910,N_3234,N_5625);
or U8911 (N_8911,N_3334,N_4503);
nor U8912 (N_8912,N_5186,N_4081);
nor U8913 (N_8913,N_3509,N_4879);
nor U8914 (N_8914,N_5284,N_4518);
and U8915 (N_8915,N_4396,N_4777);
or U8916 (N_8916,N_3535,N_5728);
and U8917 (N_8917,N_4094,N_4399);
and U8918 (N_8918,N_4192,N_4459);
nor U8919 (N_8919,N_5581,N_3860);
or U8920 (N_8920,N_5831,N_4874);
and U8921 (N_8921,N_3370,N_3161);
nor U8922 (N_8922,N_5626,N_5729);
or U8923 (N_8923,N_3670,N_3868);
nand U8924 (N_8924,N_3530,N_5566);
nor U8925 (N_8925,N_4121,N_5928);
and U8926 (N_8926,N_5109,N_4801);
nor U8927 (N_8927,N_5169,N_4107);
nand U8928 (N_8928,N_5806,N_3231);
and U8929 (N_8929,N_3155,N_4805);
and U8930 (N_8930,N_4077,N_5456);
or U8931 (N_8931,N_5113,N_4062);
nand U8932 (N_8932,N_4257,N_5776);
and U8933 (N_8933,N_3814,N_4432);
nand U8934 (N_8934,N_5885,N_5116);
nand U8935 (N_8935,N_5494,N_5545);
xor U8936 (N_8936,N_4988,N_3156);
nand U8937 (N_8937,N_3662,N_4374);
or U8938 (N_8938,N_5883,N_4675);
nand U8939 (N_8939,N_3495,N_3157);
and U8940 (N_8940,N_5306,N_5113);
nand U8941 (N_8941,N_5288,N_5043);
nand U8942 (N_8942,N_3901,N_5902);
nand U8943 (N_8943,N_4866,N_5942);
or U8944 (N_8944,N_5960,N_5808);
nor U8945 (N_8945,N_3462,N_4522);
nand U8946 (N_8946,N_4021,N_4946);
nand U8947 (N_8947,N_5533,N_4972);
or U8948 (N_8948,N_4862,N_3525);
or U8949 (N_8949,N_5229,N_5379);
and U8950 (N_8950,N_5711,N_3830);
and U8951 (N_8951,N_4745,N_3599);
and U8952 (N_8952,N_3564,N_3255);
or U8953 (N_8953,N_5752,N_3790);
and U8954 (N_8954,N_3002,N_3308);
nor U8955 (N_8955,N_5519,N_4610);
or U8956 (N_8956,N_5058,N_3013);
xnor U8957 (N_8957,N_3591,N_4084);
nand U8958 (N_8958,N_4935,N_5976);
or U8959 (N_8959,N_3482,N_3183);
and U8960 (N_8960,N_4397,N_3648);
nor U8961 (N_8961,N_5219,N_5062);
nor U8962 (N_8962,N_4118,N_5080);
nand U8963 (N_8963,N_4663,N_4680);
and U8964 (N_8964,N_4544,N_4867);
nand U8965 (N_8965,N_3161,N_5771);
nor U8966 (N_8966,N_3029,N_4860);
nand U8967 (N_8967,N_3015,N_4919);
nor U8968 (N_8968,N_4405,N_5653);
and U8969 (N_8969,N_4178,N_3865);
nand U8970 (N_8970,N_4217,N_3493);
nand U8971 (N_8971,N_4971,N_3602);
nand U8972 (N_8972,N_4543,N_5616);
xnor U8973 (N_8973,N_4827,N_3857);
and U8974 (N_8974,N_4658,N_3260);
and U8975 (N_8975,N_5908,N_3294);
or U8976 (N_8976,N_4186,N_5264);
nor U8977 (N_8977,N_4000,N_3783);
nor U8978 (N_8978,N_3520,N_3071);
and U8979 (N_8979,N_4684,N_3422);
nor U8980 (N_8980,N_3211,N_3190);
nand U8981 (N_8981,N_5448,N_5967);
or U8982 (N_8982,N_5372,N_4624);
nand U8983 (N_8983,N_4075,N_4243);
or U8984 (N_8984,N_4519,N_5707);
or U8985 (N_8985,N_3113,N_3945);
or U8986 (N_8986,N_4859,N_3656);
or U8987 (N_8987,N_3693,N_5044);
nor U8988 (N_8988,N_4174,N_5696);
and U8989 (N_8989,N_5152,N_5097);
and U8990 (N_8990,N_3421,N_3982);
and U8991 (N_8991,N_4382,N_3459);
nand U8992 (N_8992,N_5764,N_3906);
or U8993 (N_8993,N_3305,N_5535);
or U8994 (N_8994,N_5245,N_5121);
nand U8995 (N_8995,N_3258,N_3220);
or U8996 (N_8996,N_5145,N_4967);
or U8997 (N_8997,N_3459,N_3285);
nand U8998 (N_8998,N_5367,N_4185);
and U8999 (N_8999,N_5538,N_5627);
and U9000 (N_9000,N_6010,N_6620);
nand U9001 (N_9001,N_8100,N_8770);
nand U9002 (N_9002,N_6684,N_8850);
and U9003 (N_9003,N_7190,N_6405);
nor U9004 (N_9004,N_8160,N_7400);
and U9005 (N_9005,N_7563,N_7506);
and U9006 (N_9006,N_7691,N_8460);
or U9007 (N_9007,N_8335,N_6993);
and U9008 (N_9008,N_6446,N_8824);
and U9009 (N_9009,N_7107,N_7581);
nand U9010 (N_9010,N_7282,N_6631);
nor U9011 (N_9011,N_6347,N_7233);
or U9012 (N_9012,N_6423,N_7343);
nand U9013 (N_9013,N_8813,N_6653);
or U9014 (N_9014,N_6475,N_6361);
nor U9015 (N_9015,N_7673,N_6056);
or U9016 (N_9016,N_7876,N_7933);
nand U9017 (N_9017,N_8282,N_7812);
and U9018 (N_9018,N_8585,N_8587);
or U9019 (N_9019,N_8801,N_7366);
or U9020 (N_9020,N_7165,N_7304);
or U9021 (N_9021,N_8441,N_8336);
nand U9022 (N_9022,N_7106,N_7639);
or U9023 (N_9023,N_8731,N_7333);
nor U9024 (N_9024,N_7450,N_8911);
and U9025 (N_9025,N_8118,N_7924);
nor U9026 (N_9026,N_8330,N_6990);
nor U9027 (N_9027,N_6739,N_7986);
nand U9028 (N_9028,N_8463,N_6542);
or U9029 (N_9029,N_6401,N_6395);
nor U9030 (N_9030,N_7605,N_8649);
nand U9031 (N_9031,N_6590,N_8570);
or U9032 (N_9032,N_8740,N_6089);
nand U9033 (N_9033,N_7626,N_7432);
nor U9034 (N_9034,N_6218,N_7861);
or U9035 (N_9035,N_6978,N_8200);
nand U9036 (N_9036,N_7126,N_6678);
and U9037 (N_9037,N_6384,N_7698);
and U9038 (N_9038,N_8959,N_7655);
and U9039 (N_9039,N_8063,N_8853);
and U9040 (N_9040,N_6176,N_8241);
nor U9041 (N_9041,N_6037,N_7497);
and U9042 (N_9042,N_7813,N_7397);
nand U9043 (N_9043,N_8641,N_8148);
nor U9044 (N_9044,N_7839,N_8970);
nor U9045 (N_9045,N_8298,N_6961);
nand U9046 (N_9046,N_7988,N_7641);
nor U9047 (N_9047,N_7765,N_7015);
nand U9048 (N_9048,N_6874,N_8104);
or U9049 (N_9049,N_6035,N_6459);
nor U9050 (N_9050,N_7380,N_7582);
nand U9051 (N_9051,N_8738,N_7818);
or U9052 (N_9052,N_8779,N_7970);
nor U9053 (N_9053,N_8943,N_6626);
and U9054 (N_9054,N_7887,N_7284);
nor U9055 (N_9055,N_8202,N_7259);
and U9056 (N_9056,N_7586,N_7437);
and U9057 (N_9057,N_8851,N_8924);
and U9058 (N_9058,N_6718,N_6344);
xor U9059 (N_9059,N_7489,N_8765);
or U9060 (N_9060,N_7923,N_7434);
nor U9061 (N_9061,N_7822,N_7474);
or U9062 (N_9062,N_8101,N_8605);
or U9063 (N_9063,N_6400,N_6505);
nand U9064 (N_9064,N_6354,N_7393);
nor U9065 (N_9065,N_6920,N_7324);
nor U9066 (N_9066,N_8533,N_8664);
nor U9067 (N_9067,N_7151,N_6875);
or U9068 (N_9068,N_7102,N_6638);
and U9069 (N_9069,N_6301,N_7121);
nand U9070 (N_9070,N_8354,N_7961);
nand U9071 (N_9071,N_8239,N_8192);
and U9072 (N_9072,N_6655,N_6440);
and U9073 (N_9073,N_8651,N_7774);
or U9074 (N_9074,N_7242,N_6456);
or U9075 (N_9075,N_6078,N_8543);
or U9076 (N_9076,N_6223,N_8506);
nand U9077 (N_9077,N_7695,N_7300);
nor U9078 (N_9078,N_7569,N_8012);
or U9079 (N_9079,N_8385,N_6801);
nand U9080 (N_9080,N_6532,N_6750);
nand U9081 (N_9081,N_8075,N_8000);
or U9082 (N_9082,N_8464,N_8279);
nand U9083 (N_9083,N_8107,N_6868);
or U9084 (N_9084,N_8375,N_6022);
nor U9085 (N_9085,N_8793,N_6646);
nand U9086 (N_9086,N_8629,N_8870);
or U9087 (N_9087,N_7409,N_6018);
and U9088 (N_9088,N_7128,N_7926);
or U9089 (N_9089,N_8842,N_7120);
or U9090 (N_9090,N_7355,N_6283);
nand U9091 (N_9091,N_6890,N_7723);
nand U9092 (N_9092,N_8359,N_6691);
and U9093 (N_9093,N_7195,N_7711);
nand U9094 (N_9094,N_8799,N_7184);
or U9095 (N_9095,N_6666,N_8652);
nand U9096 (N_9096,N_7344,N_6489);
or U9097 (N_9097,N_7656,N_6723);
and U9098 (N_9098,N_8611,N_8519);
nor U9099 (N_9099,N_6327,N_7199);
or U9100 (N_9100,N_6997,N_8412);
nor U9101 (N_9101,N_7020,N_8708);
and U9102 (N_9102,N_8630,N_6892);
nor U9103 (N_9103,N_7441,N_6178);
and U9104 (N_9104,N_6225,N_7252);
and U9105 (N_9105,N_6445,N_8676);
and U9106 (N_9106,N_8092,N_8727);
and U9107 (N_9107,N_6659,N_7328);
nand U9108 (N_9108,N_8673,N_6586);
and U9109 (N_9109,N_7447,N_6469);
and U9110 (N_9110,N_8219,N_7023);
and U9111 (N_9111,N_7049,N_6944);
nor U9112 (N_9112,N_7918,N_7636);
or U9113 (N_9113,N_8584,N_6396);
nor U9114 (N_9114,N_7222,N_7751);
or U9115 (N_9115,N_7521,N_8531);
or U9116 (N_9116,N_7978,N_7171);
nand U9117 (N_9117,N_8030,N_6486);
and U9118 (N_9118,N_6434,N_6724);
and U9119 (N_9119,N_8480,N_8961);
and U9120 (N_9120,N_7584,N_8302);
or U9121 (N_9121,N_6166,N_7935);
nand U9122 (N_9122,N_8348,N_7492);
and U9123 (N_9123,N_8536,N_6209);
or U9124 (N_9124,N_6113,N_6851);
and U9125 (N_9125,N_6317,N_8266);
nor U9126 (N_9126,N_7330,N_8149);
nand U9127 (N_9127,N_7231,N_6118);
and U9128 (N_9128,N_6135,N_8973);
nand U9129 (N_9129,N_7541,N_7485);
or U9130 (N_9130,N_8129,N_6714);
and U9131 (N_9131,N_7824,N_8036);
or U9132 (N_9132,N_7356,N_7276);
and U9133 (N_9133,N_6557,N_7227);
and U9134 (N_9134,N_7285,N_7281);
nand U9135 (N_9135,N_7709,N_8748);
nor U9136 (N_9136,N_8841,N_7033);
nor U9137 (N_9137,N_8600,N_8314);
nor U9138 (N_9138,N_7214,N_8556);
nor U9139 (N_9139,N_8142,N_8168);
or U9140 (N_9140,N_8274,N_7863);
or U9141 (N_9141,N_6364,N_6329);
nor U9142 (N_9142,N_8918,N_6378);
nor U9143 (N_9143,N_8618,N_8325);
nor U9144 (N_9144,N_7189,N_8544);
nor U9145 (N_9145,N_8019,N_7209);
nand U9146 (N_9146,N_8729,N_8095);
or U9147 (N_9147,N_8828,N_7613);
nand U9148 (N_9148,N_8420,N_7994);
and U9149 (N_9149,N_6270,N_8322);
and U9150 (N_9150,N_7144,N_8760);
and U9151 (N_9151,N_7286,N_7414);
and U9152 (N_9152,N_8426,N_7725);
nor U9153 (N_9153,N_8462,N_6133);
nand U9154 (N_9154,N_6121,N_6312);
nor U9155 (N_9155,N_7311,N_8331);
nor U9156 (N_9156,N_7538,N_7159);
nand U9157 (N_9157,N_6200,N_7325);
or U9158 (N_9158,N_7309,N_6161);
nor U9159 (N_9159,N_6951,N_6970);
nand U9160 (N_9160,N_7481,N_8317);
nor U9161 (N_9161,N_6972,N_8127);
and U9162 (N_9162,N_8508,N_6611);
nor U9163 (N_9163,N_6231,N_8007);
nor U9164 (N_9164,N_6303,N_8589);
nand U9165 (N_9165,N_7827,N_6389);
or U9166 (N_9166,N_6485,N_7158);
and U9167 (N_9167,N_6214,N_8747);
nand U9168 (N_9168,N_8419,N_7053);
and U9169 (N_9169,N_7891,N_7118);
nand U9170 (N_9170,N_6612,N_7999);
or U9171 (N_9171,N_8830,N_6262);
and U9172 (N_9172,N_7490,N_8437);
or U9173 (N_9173,N_7044,N_8262);
and U9174 (N_9174,N_6044,N_7019);
nand U9175 (N_9175,N_7235,N_8137);
and U9176 (N_9176,N_6331,N_7901);
and U9177 (N_9177,N_7200,N_8287);
nand U9178 (N_9178,N_8915,N_6585);
nand U9179 (N_9179,N_7660,N_8203);
nand U9180 (N_9180,N_6449,N_7833);
or U9181 (N_9181,N_7098,N_8761);
and U9182 (N_9182,N_6786,N_8675);
nor U9183 (N_9183,N_8581,N_6987);
nor U9184 (N_9184,N_6358,N_7726);
nand U9185 (N_9185,N_7795,N_6922);
nor U9186 (N_9186,N_7853,N_7975);
nand U9187 (N_9187,N_6735,N_7805);
and U9188 (N_9188,N_6315,N_8020);
nor U9189 (N_9189,N_7801,N_7456);
nand U9190 (N_9190,N_6151,N_7676);
and U9191 (N_9191,N_6550,N_6241);
nand U9192 (N_9192,N_6840,N_6265);
and U9193 (N_9193,N_7410,N_8739);
or U9194 (N_9194,N_8424,N_6424);
and U9195 (N_9195,N_7472,N_7576);
and U9196 (N_9196,N_7722,N_6249);
or U9197 (N_9197,N_8763,N_7316);
or U9198 (N_9198,N_6066,N_6212);
or U9199 (N_9199,N_8667,N_8947);
nor U9200 (N_9200,N_7368,N_6776);
or U9201 (N_9201,N_8491,N_7154);
nand U9202 (N_9202,N_8212,N_7848);
nor U9203 (N_9203,N_7954,N_7059);
or U9204 (N_9204,N_6994,N_7750);
nand U9205 (N_9205,N_7479,N_7577);
or U9206 (N_9206,N_6180,N_8159);
and U9207 (N_9207,N_7606,N_7076);
nand U9208 (N_9208,N_6957,N_8762);
nand U9209 (N_9209,N_8364,N_8068);
or U9210 (N_9210,N_6269,N_7303);
or U9211 (N_9211,N_6919,N_7379);
or U9212 (N_9212,N_8473,N_6592);
and U9213 (N_9213,N_7788,N_7082);
nand U9214 (N_9214,N_8048,N_7369);
or U9215 (N_9215,N_7160,N_8646);
or U9216 (N_9216,N_8874,N_7706);
nand U9217 (N_9217,N_6103,N_8610);
and U9218 (N_9218,N_6722,N_6802);
and U9219 (N_9219,N_7790,N_7141);
and U9220 (N_9220,N_7864,N_6268);
nand U9221 (N_9221,N_6837,N_6895);
nand U9222 (N_9222,N_8808,N_8757);
nand U9223 (N_9223,N_6237,N_7390);
nor U9224 (N_9224,N_8032,N_7599);
nand U9225 (N_9225,N_6584,N_8848);
and U9226 (N_9226,N_7939,N_6527);
or U9227 (N_9227,N_8522,N_8714);
nor U9228 (N_9228,N_7216,N_6810);
and U9229 (N_9229,N_8777,N_8690);
nor U9230 (N_9230,N_7405,N_6232);
or U9231 (N_9231,N_6379,N_7283);
nand U9232 (N_9232,N_7928,N_6322);
or U9233 (N_9233,N_7520,N_6179);
nor U9234 (N_9234,N_7399,N_8070);
and U9235 (N_9235,N_8328,N_7731);
and U9236 (N_9236,N_7712,N_7187);
nand U9237 (N_9237,N_6906,N_8498);
nor U9238 (N_9238,N_6478,N_6539);
nand U9239 (N_9239,N_8838,N_7984);
nand U9240 (N_9240,N_7539,N_7564);
nand U9241 (N_9241,N_6187,N_6336);
or U9242 (N_9242,N_8832,N_7218);
nor U9243 (N_9243,N_8146,N_7512);
and U9244 (N_9244,N_6497,N_6554);
or U9245 (N_9245,N_8607,N_8505);
nor U9246 (N_9246,N_8422,N_6762);
nand U9247 (N_9247,N_8246,N_8694);
nor U9248 (N_9248,N_8827,N_7460);
nor U9249 (N_9249,N_8242,N_6233);
or U9250 (N_9250,N_6097,N_7873);
and U9251 (N_9251,N_7640,N_6383);
and U9252 (N_9252,N_8861,N_8493);
nor U9253 (N_9253,N_8091,N_6641);
nor U9254 (N_9254,N_7769,N_7557);
or U9255 (N_9255,N_7888,N_8257);
nand U9256 (N_9256,N_7401,N_7845);
and U9257 (N_9257,N_6615,N_8488);
nand U9258 (N_9258,N_8016,N_8178);
nor U9259 (N_9259,N_8632,N_7775);
or U9260 (N_9260,N_8253,N_6228);
or U9261 (N_9261,N_7406,N_7302);
or U9262 (N_9262,N_8014,N_8555);
xor U9263 (N_9263,N_6912,N_7882);
nor U9264 (N_9264,N_6453,N_7271);
and U9265 (N_9265,N_6227,N_8660);
nand U9266 (N_9266,N_6467,N_7088);
and U9267 (N_9267,N_6516,N_6885);
or U9268 (N_9268,N_6551,N_6660);
or U9269 (N_9269,N_8988,N_8197);
nor U9270 (N_9270,N_8711,N_7364);
nor U9271 (N_9271,N_8971,N_8450);
nand U9272 (N_9272,N_8005,N_6192);
nand U9273 (N_9273,N_7560,N_7558);
nor U9274 (N_9274,N_8472,N_6328);
nand U9275 (N_9275,N_6864,N_6145);
and U9276 (N_9276,N_6063,N_8256);
and U9277 (N_9277,N_8414,N_8477);
or U9278 (N_9278,N_8042,N_8678);
xnor U9279 (N_9279,N_8749,N_7256);
or U9280 (N_9280,N_6075,N_6777);
or U9281 (N_9281,N_8873,N_8656);
and U9282 (N_9282,N_6706,N_8897);
nor U9283 (N_9283,N_6877,N_7219);
nor U9284 (N_9284,N_8164,N_8550);
nand U9285 (N_9285,N_7186,N_8367);
and U9286 (N_9286,N_6363,N_7395);
or U9287 (N_9287,N_7001,N_7335);
or U9288 (N_9288,N_6578,N_6980);
and U9289 (N_9289,N_8310,N_6435);
nor U9290 (N_9290,N_7646,N_6355);
and U9291 (N_9291,N_8677,N_7056);
nand U9292 (N_9292,N_7573,N_7346);
and U9293 (N_9293,N_6515,N_6402);
nor U9294 (N_9294,N_7525,N_7163);
and U9295 (N_9295,N_6753,N_8475);
or U9296 (N_9296,N_8914,N_8225);
and U9297 (N_9297,N_8735,N_8237);
nor U9298 (N_9298,N_8297,N_6211);
or U9299 (N_9299,N_8388,N_8431);
or U9300 (N_9300,N_7772,N_8776);
or U9301 (N_9301,N_7119,N_6153);
nand U9302 (N_9302,N_8213,N_6887);
nor U9303 (N_9303,N_7721,N_7846);
nand U9304 (N_9304,N_6052,N_6308);
nand U9305 (N_9305,N_8980,N_8248);
xnor U9306 (N_9306,N_6084,N_7062);
and U9307 (N_9307,N_6282,N_7137);
nand U9308 (N_9308,N_7315,N_8175);
nand U9309 (N_9309,N_7111,N_6642);
nand U9310 (N_9310,N_7927,N_7890);
nand U9311 (N_9311,N_7357,N_8347);
and U9312 (N_9312,N_6791,N_8109);
or U9313 (N_9313,N_8376,N_7530);
nor U9314 (N_9314,N_7168,N_7246);
nand U9315 (N_9315,N_7420,N_6736);
nor U9316 (N_9316,N_7900,N_7844);
and U9317 (N_9317,N_6900,N_7650);
nor U9318 (N_9318,N_7327,N_7819);
or U9319 (N_9319,N_7592,N_6464);
nand U9320 (N_9320,N_7943,N_8767);
and U9321 (N_9321,N_8295,N_6155);
nand U9322 (N_9322,N_6427,N_6108);
nor U9323 (N_9323,N_7510,N_6130);
or U9324 (N_9324,N_7310,N_7229);
and U9325 (N_9325,N_6512,N_8560);
nor U9326 (N_9326,N_6725,N_8534);
or U9327 (N_9327,N_6356,N_6841);
and U9328 (N_9328,N_7828,N_7081);
or U9329 (N_9329,N_6280,N_7247);
or U9330 (N_9330,N_8957,N_8083);
nor U9331 (N_9331,N_6125,N_6186);
nor U9332 (N_9332,N_8936,N_7260);
and U9333 (N_9333,N_8901,N_6468);
or U9334 (N_9334,N_7261,N_8571);
and U9335 (N_9335,N_8120,N_6934);
nor U9336 (N_9336,N_6996,N_7419);
and U9337 (N_9337,N_6968,N_8954);
nor U9338 (N_9338,N_6815,N_8133);
and U9339 (N_9339,N_6945,N_7947);
nand U9340 (N_9340,N_7297,N_8114);
nor U9341 (N_9341,N_7683,N_7708);
and U9342 (N_9342,N_6021,N_7099);
nor U9343 (N_9343,N_6937,N_7796);
nand U9344 (N_9344,N_8602,N_6558);
nand U9345 (N_9345,N_6398,N_7880);
xor U9346 (N_9346,N_7294,N_6134);
nor U9347 (N_9347,N_8964,N_7299);
nand U9348 (N_9348,N_8965,N_7425);
and U9349 (N_9349,N_8486,N_7508);
and U9350 (N_9350,N_7135,N_8717);
nor U9351 (N_9351,N_7152,N_6335);
nand U9352 (N_9352,N_6392,N_7729);
or U9353 (N_9353,N_6829,N_6704);
or U9354 (N_9354,N_7161,N_6414);
nor U9355 (N_9355,N_7651,N_8408);
nor U9356 (N_9356,N_6323,N_8963);
and U9357 (N_9357,N_7625,N_7074);
nor U9358 (N_9358,N_6368,N_7264);
nor U9359 (N_9359,N_6658,N_8126);
and U9360 (N_9360,N_6340,N_8878);
nor U9361 (N_9361,N_8028,N_7741);
or U9362 (N_9362,N_8860,N_8902);
nor U9363 (N_9363,N_6733,N_8260);
and U9364 (N_9364,N_8448,N_7453);
nor U9365 (N_9365,N_8162,N_6962);
or U9366 (N_9366,N_6928,N_6524);
nand U9367 (N_9367,N_8590,N_8184);
or U9368 (N_9368,N_6275,N_7945);
nor U9369 (N_9369,N_6817,N_8945);
nor U9370 (N_9370,N_7411,N_7753);
or U9371 (N_9371,N_6047,N_7457);
and U9372 (N_9372,N_7480,N_8134);
nor U9373 (N_9373,N_8350,N_7179);
and U9374 (N_9374,N_8796,N_7644);
nor U9375 (N_9375,N_8542,N_7793);
nand U9376 (N_9376,N_6501,N_8045);
and U9377 (N_9377,N_7546,N_6170);
and U9378 (N_9378,N_6734,N_6309);
nand U9379 (N_9379,N_8051,N_8983);
nor U9380 (N_9380,N_7013,N_7280);
and U9381 (N_9381,N_7667,N_8825);
nand U9382 (N_9382,N_8829,N_6544);
and U9383 (N_9383,N_7045,N_7570);
nand U9384 (N_9384,N_7178,N_7779);
and U9385 (N_9385,N_8292,N_8831);
and U9386 (N_9386,N_8946,N_6796);
or U9387 (N_9387,N_6599,N_6955);
and U9388 (N_9388,N_8593,N_8374);
or U9389 (N_9389,N_8352,N_8261);
and U9390 (N_9390,N_6152,N_6117);
xnor U9391 (N_9391,N_8709,N_7980);
xnor U9392 (N_9392,N_7471,N_8906);
nand U9393 (N_9393,N_7476,N_8156);
and U9394 (N_9394,N_6519,N_6958);
nor U9395 (N_9395,N_6305,N_8236);
nand U9396 (N_9396,N_8461,N_7814);
and U9397 (N_9397,N_6393,N_7465);
nand U9398 (N_9398,N_7338,N_8913);
nor U9399 (N_9399,N_8620,N_6844);
and U9400 (N_9400,N_7898,N_7604);
nand U9401 (N_9401,N_6253,N_8222);
and U9402 (N_9402,N_6029,N_6698);
nand U9403 (N_9403,N_7549,N_7792);
and U9404 (N_9404,N_7830,N_7206);
and U9405 (N_9405,N_8147,N_6112);
or U9406 (N_9406,N_8639,N_7534);
and U9407 (N_9407,N_7413,N_7136);
and U9408 (N_9408,N_8953,N_8784);
and U9409 (N_9409,N_7872,N_6013);
xor U9410 (N_9410,N_6897,N_8840);
nor U9411 (N_9411,N_7782,N_7204);
or U9412 (N_9412,N_6605,N_6004);
and U9413 (N_9413,N_7621,N_6616);
nand U9414 (N_9414,N_7585,N_8423);
or U9415 (N_9415,N_7298,N_8806);
nor U9416 (N_9416,N_8859,N_8663);
nand U9417 (N_9417,N_7825,N_8938);
nand U9418 (N_9418,N_8500,N_6346);
nor U9419 (N_9419,N_7421,N_8898);
nand U9420 (N_9420,N_7951,N_8903);
nand U9421 (N_9421,N_8465,N_6737);
nor U9422 (N_9422,N_7087,N_8856);
or U9423 (N_9423,N_8254,N_7942);
nand U9424 (N_9424,N_8135,N_7679);
nand U9425 (N_9425,N_8532,N_8153);
or U9426 (N_9426,N_7503,N_8528);
nand U9427 (N_9427,N_8283,N_8190);
nor U9428 (N_9428,N_8251,N_8659);
nand U9429 (N_9429,N_7452,N_6109);
nand U9430 (N_9430,N_6000,N_7245);
or U9431 (N_9431,N_6549,N_6861);
nor U9432 (N_9432,N_7267,N_6741);
and U9433 (N_9433,N_6795,N_8545);
nor U9434 (N_9434,N_7365,N_8792);
nor U9435 (N_9435,N_8710,N_7682);
and U9436 (N_9436,N_6421,N_6416);
nor U9437 (N_9437,N_8205,N_7720);
and U9438 (N_9438,N_7856,N_6778);
and U9439 (N_9439,N_7496,N_7095);
nor U9440 (N_9440,N_7342,N_7645);
or U9441 (N_9441,N_8598,N_6410);
and U9442 (N_9442,N_7865,N_6483);
and U9443 (N_9443,N_7759,N_6633);
nor U9444 (N_9444,N_6831,N_8785);
or U9445 (N_9445,N_8379,N_6098);
nor U9446 (N_9446,N_6479,N_6183);
and U9447 (N_9447,N_6482,N_7685);
nand U9448 (N_9448,N_8929,N_6255);
or U9449 (N_9449,N_7170,N_6832);
and U9450 (N_9450,N_8301,N_6950);
nand U9451 (N_9451,N_7791,N_6163);
and U9452 (N_9452,N_6530,N_8235);
nand U9453 (N_9453,N_6419,N_7616);
or U9454 (N_9454,N_6277,N_6732);
or U9455 (N_9455,N_7764,N_7551);
nand U9456 (N_9456,N_6731,N_7628);
nand U9457 (N_9457,N_7883,N_8391);
xnor U9458 (N_9458,N_8113,N_7296);
and U9459 (N_9459,N_7114,N_7067);
and U9460 (N_9460,N_6805,N_8382);
or U9461 (N_9461,N_8997,N_7132);
and U9462 (N_9462,N_8182,N_6476);
nand U9463 (N_9463,N_6362,N_8323);
and U9464 (N_9464,N_8769,N_7312);
nor U9465 (N_9465,N_7835,N_7279);
and U9466 (N_9466,N_8716,N_7587);
and U9467 (N_9467,N_8557,N_8619);
and U9468 (N_9468,N_7993,N_8691);
nor U9469 (N_9469,N_7717,N_7478);
or U9470 (N_9470,N_8278,N_8567);
nor U9471 (N_9471,N_7666,N_8196);
nand U9472 (N_9472,N_6701,N_7373);
nor U9473 (N_9473,N_8204,N_8128);
or U9474 (N_9474,N_8504,N_7174);
nand U9475 (N_9475,N_6325,N_6792);
nand U9476 (N_9476,N_6999,N_6694);
or U9477 (N_9477,N_7700,N_8002);
nand U9478 (N_9478,N_8920,N_8642);
nand U9479 (N_9479,N_8208,N_6054);
or U9480 (N_9480,N_7248,N_8948);
nor U9481 (N_9481,N_6065,N_7042);
nand U9482 (N_9482,N_6789,N_7439);
nand U9483 (N_9483,N_6717,N_6046);
and U9484 (N_9484,N_6597,N_6058);
nand U9485 (N_9485,N_8723,N_6905);
nand U9486 (N_9486,N_6956,N_6746);
or U9487 (N_9487,N_7799,N_7398);
nor U9488 (N_9488,N_6690,N_8327);
nor U9489 (N_9489,N_8839,N_7418);
or U9490 (N_9490,N_6806,N_6634);
and U9491 (N_9491,N_7351,N_6728);
nor U9492 (N_9492,N_8201,N_8568);
nand U9493 (N_9493,N_8791,N_7009);
and U9494 (N_9494,N_8866,N_6657);
nand U9495 (N_9495,N_6193,N_6727);
or U9496 (N_9496,N_6219,N_8687);
nor U9497 (N_9497,N_6106,N_7167);
and U9498 (N_9498,N_6859,N_6008);
and U9499 (N_9499,N_6122,N_6374);
and U9500 (N_9500,N_7331,N_6337);
nor U9501 (N_9501,N_8170,N_7547);
or U9502 (N_9502,N_8277,N_8199);
nand U9503 (N_9503,N_8746,N_7208);
and U9504 (N_9504,N_8577,N_8181);
nor U9505 (N_9505,N_7877,N_8362);
nor U9506 (N_9506,N_6663,N_8966);
or U9507 (N_9507,N_8023,N_7983);
nor U9508 (N_9508,N_8734,N_7652);
nor U9509 (N_9509,N_7874,N_8549);
nand U9510 (N_9510,N_7967,N_7972);
or U9511 (N_9511,N_8112,N_6100);
nand U9512 (N_9512,N_7024,N_7384);
nor U9513 (N_9513,N_7739,N_7579);
and U9514 (N_9514,N_7070,N_6165);
or U9515 (N_9515,N_7803,N_7672);
xor U9516 (N_9516,N_6502,N_8077);
nand U9517 (N_9517,N_8291,N_8141);
or U9518 (N_9518,N_8061,N_8919);
nand U9519 (N_9519,N_7594,N_6441);
nor U9520 (N_9520,N_7462,N_8221);
or U9521 (N_9521,N_7913,N_7958);
or U9522 (N_9522,N_8693,N_6935);
and U9523 (N_9523,N_8010,N_6466);
or U9524 (N_9524,N_7046,N_6050);
nand U9525 (N_9525,N_7662,N_6229);
nand U9526 (N_9526,N_7854,N_8115);
nor U9527 (N_9527,N_8290,N_8227);
nand U9528 (N_9528,N_6992,N_8518);
and U9529 (N_9529,N_6099,N_7507);
nor U9530 (N_9530,N_6986,N_8099);
nor U9531 (N_9531,N_6438,N_7386);
and U9532 (N_9532,N_8737,N_7806);
and U9533 (N_9533,N_6751,N_6238);
and U9534 (N_9534,N_8270,N_7292);
nor U9535 (N_9535,N_6692,N_6856);
nor U9536 (N_9536,N_7155,N_8650);
or U9537 (N_9537,N_6821,N_6738);
or U9538 (N_9538,N_6509,N_6302);
or U9539 (N_9539,N_8858,N_7925);
nand U9540 (N_9540,N_8993,N_6017);
nand U9541 (N_9541,N_6357,N_6748);
nand U9542 (N_9542,N_7860,N_7275);
nand U9543 (N_9543,N_8284,N_6824);
nand U9544 (N_9544,N_8978,N_8977);
nor U9545 (N_9545,N_7878,N_7934);
or U9546 (N_9546,N_7562,N_7408);
nand U9547 (N_9547,N_6600,N_8643);
nor U9548 (N_9548,N_8495,N_8854);
or U9549 (N_9549,N_7424,N_7635);
and U9550 (N_9550,N_6839,N_6548);
and U9551 (N_9551,N_8218,N_7536);
or U9552 (N_9552,N_8941,N_7502);
nand U9553 (N_9553,N_7664,N_8249);
or U9554 (N_9554,N_8683,N_8794);
and U9555 (N_9555,N_6290,N_7445);
nor U9556 (N_9556,N_8670,N_8108);
and U9557 (N_9557,N_7113,N_8718);
or U9558 (N_9558,N_8833,N_8198);
and U9559 (N_9559,N_6371,N_6858);
nand U9560 (N_9560,N_6375,N_8443);
or U9561 (N_9561,N_8054,N_6068);
or U9562 (N_9562,N_8052,N_6598);
or U9563 (N_9563,N_7583,N_7797);
nor U9564 (N_9564,N_7843,N_8349);
nor U9565 (N_9565,N_8381,N_8612);
nor U9566 (N_9566,N_7244,N_6552);
and U9567 (N_9567,N_8622,N_7704);
or U9568 (N_9568,N_6070,N_6568);
nor U9569 (N_9569,N_7193,N_6319);
nand U9570 (N_9570,N_6291,N_8836);
or U9571 (N_9571,N_8377,N_6266);
nor U9572 (N_9572,N_6158,N_6581);
nand U9573 (N_9573,N_6577,N_7198);
and U9574 (N_9574,N_8719,N_6849);
and U9575 (N_9575,N_7498,N_7182);
or U9576 (N_9576,N_8214,N_7851);
nor U9577 (N_9577,N_8053,N_6349);
and U9578 (N_9578,N_6760,N_6043);
or U9579 (N_9579,N_8880,N_6074);
nand U9580 (N_9580,N_6391,N_6721);
nor U9581 (N_9581,N_7277,N_6332);
nand U9582 (N_9582,N_7960,N_7162);
nor U9583 (N_9583,N_8435,N_7871);
xor U9584 (N_9584,N_7225,N_7763);
and U9585 (N_9585,N_6205,N_6142);
nor U9586 (N_9586,N_7973,N_6518);
and U9587 (N_9587,N_8855,N_7719);
and U9588 (N_9588,N_8985,N_8684);
or U9589 (N_9589,N_6168,N_6556);
nand U9590 (N_9590,N_7869,N_8682);
or U9591 (N_9591,N_8986,N_6490);
or U9592 (N_9592,N_8318,N_6009);
or U9593 (N_9593,N_6898,N_8043);
or U9594 (N_9594,N_8787,N_8165);
nor U9595 (N_9595,N_6442,N_6785);
nor U9596 (N_9596,N_6793,N_8937);
or U9597 (N_9597,N_8636,N_6132);
nor U9598 (N_9598,N_8172,N_6073);
or U9599 (N_9599,N_6822,N_6886);
or U9600 (N_9600,N_6111,N_6139);
xnor U9601 (N_9601,N_7509,N_8163);
nor U9602 (N_9602,N_7896,N_6865);
and U9603 (N_9603,N_7029,N_6930);
and U9604 (N_9604,N_6235,N_6720);
and U9605 (N_9605,N_6259,N_7981);
or U9606 (N_9606,N_7491,N_6069);
or U9607 (N_9607,N_7744,N_6463);
nand U9608 (N_9608,N_8846,N_7254);
nand U9609 (N_9609,N_6545,N_8469);
and U9610 (N_9610,N_7964,N_6670);
nor U9611 (N_9611,N_7962,N_7817);
or U9612 (N_9612,N_6669,N_7468);
nand U9613 (N_9613,N_8276,N_6879);
nor U9614 (N_9614,N_6667,N_6496);
and U9615 (N_9615,N_7713,N_6093);
nand U9616 (N_9616,N_7987,N_7207);
nand U9617 (N_9617,N_7417,N_7362);
and U9618 (N_9618,N_6217,N_8195);
and U9619 (N_9619,N_8247,N_7429);
nor U9620 (N_9620,N_7443,N_6215);
nand U9621 (N_9621,N_8013,N_8783);
nor U9622 (N_9622,N_6546,N_7270);
or U9623 (N_9623,N_8805,N_8586);
or U9624 (N_9624,N_7084,N_8098);
or U9625 (N_9625,N_6116,N_6896);
and U9626 (N_9626,N_6036,N_6494);
or U9627 (N_9627,N_7879,N_6366);
or U9628 (N_9628,N_8125,N_6039);
and U9629 (N_9629,N_8837,N_8096);
or U9630 (N_9630,N_7638,N_8515);
nand U9631 (N_9631,N_8883,N_6474);
and U9632 (N_9632,N_7117,N_8501);
nand U9633 (N_9633,N_8228,N_7077);
xnor U9634 (N_9634,N_8753,N_8551);
and U9635 (N_9635,N_8921,N_8174);
and U9636 (N_9636,N_8686,N_7370);
nand U9637 (N_9637,N_6601,N_8759);
and U9638 (N_9638,N_6430,N_6250);
nand U9639 (N_9639,N_8666,N_8427);
and U9640 (N_9640,N_6324,N_7350);
or U9641 (N_9641,N_7832,N_7665);
nor U9642 (N_9642,N_6081,N_6201);
nand U9643 (N_9643,N_7959,N_6610);
and U9644 (N_9644,N_6110,N_6529);
nand U9645 (N_9645,N_8105,N_8516);
or U9646 (N_9646,N_6848,N_8627);
and U9647 (N_9647,N_6889,N_8722);
or U9648 (N_9648,N_6451,N_8378);
and U9649 (N_9649,N_8080,N_7018);
nand U9650 (N_9650,N_6630,N_8458);
nor U9651 (N_9651,N_6436,N_8699);
or U9652 (N_9652,N_6120,N_8299);
nor U9653 (N_9653,N_8972,N_6621);
or U9654 (N_9654,N_7278,N_7301);
or U9655 (N_9655,N_7430,N_8417);
nor U9656 (N_9656,N_7730,N_7505);
and U9657 (N_9657,N_7483,N_6462);
nor U9658 (N_9658,N_8741,N_7929);
and U9659 (N_9659,N_6816,N_6560);
nor U9660 (N_9660,N_6297,N_6665);
nand U9661 (N_9661,N_8591,N_8442);
and U9662 (N_9662,N_7705,N_6051);
nor U9663 (N_9663,N_7372,N_7404);
and U9664 (N_9664,N_8345,N_7212);
nand U9665 (N_9665,N_7561,N_8554);
nor U9666 (N_9666,N_6812,N_6107);
or U9667 (N_9667,N_7976,N_6353);
xnor U9668 (N_9668,N_7979,N_8967);
and U9669 (N_9669,N_6273,N_8672);
or U9670 (N_9670,N_8730,N_6272);
nand U9671 (N_9671,N_6729,N_8703);
or U9672 (N_9672,N_7532,N_7752);
nor U9673 (N_9673,N_6064,N_7367);
and U9674 (N_9674,N_8403,N_8782);
or U9675 (N_9675,N_8707,N_7501);
nand U9676 (N_9676,N_8807,N_7798);
nor U9677 (N_9677,N_7684,N_8539);
or U9678 (N_9678,N_7363,N_7523);
or U9679 (N_9679,N_8040,N_8333);
or U9680 (N_9680,N_6471,N_6863);
nor U9681 (N_9681,N_6860,N_7057);
nand U9682 (N_9682,N_7093,N_8090);
nor U9683 (N_9683,N_6244,N_7268);
and U9684 (N_9684,N_7771,N_7620);
and U9685 (N_9685,N_8312,N_7052);
nand U9686 (N_9686,N_7540,N_6716);
nor U9687 (N_9687,N_8363,N_7122);
nor U9688 (N_9688,N_6876,N_6939);
nand U9689 (N_9689,N_6783,N_8188);
nor U9690 (N_9690,N_8017,N_6705);
nor U9691 (N_9691,N_8059,N_6564);
and U9692 (N_9692,N_7157,N_7670);
and U9693 (N_9693,N_7230,N_8244);
nand U9694 (N_9694,N_6662,N_6715);
or U9695 (N_9695,N_7668,N_6007);
nand U9696 (N_9696,N_7321,N_7897);
or U9697 (N_9697,N_6182,N_6917);
or U9698 (N_9698,N_7176,N_7036);
or U9699 (N_9699,N_8527,N_6974);
or U9700 (N_9700,N_6020,N_6596);
nand U9701 (N_9701,N_6418,N_8987);
nor U9702 (N_9702,N_8546,N_8595);
and U9703 (N_9703,N_6891,N_6213);
or U9704 (N_9704,N_6799,N_8538);
or U9705 (N_9705,N_6087,N_8255);
nor U9706 (N_9706,N_6147,N_6406);
or U9707 (N_9707,N_6632,N_8613);
nand U9708 (N_9708,N_7808,N_7051);
and U9709 (N_9709,N_6888,N_7156);
nor U9710 (N_9710,N_7780,N_8339);
nand U9711 (N_9711,N_6311,N_8313);
nor U9712 (N_9712,N_8006,N_8608);
or U9713 (N_9713,N_6454,N_8233);
nor U9714 (N_9714,N_7781,N_7050);
nand U9715 (N_9715,N_7580,N_6077);
nand U9716 (N_9716,N_7747,N_7458);
nor U9717 (N_9717,N_6604,N_8922);
and U9718 (N_9718,N_8823,N_6903);
and U9719 (N_9719,N_6710,N_7513);
and U9720 (N_9720,N_6730,N_7047);
and U9721 (N_9721,N_8822,N_7391);
nor U9722 (N_9722,N_8386,N_8304);
or U9723 (N_9723,N_6012,N_6061);
or U9724 (N_9724,N_7965,N_7575);
nand U9725 (N_9725,N_8790,N_8240);
or U9726 (N_9726,N_6673,N_6288);
nor U9727 (N_9727,N_8238,N_6541);
or U9728 (N_9728,N_7007,N_6342);
and U9729 (N_9729,N_6742,N_7694);
nor U9730 (N_9730,N_6932,N_7908);
nand U9731 (N_9731,N_7089,N_7461);
or U9732 (N_9732,N_6834,N_6144);
and U9733 (N_9733,N_8698,N_8418);
nor U9734 (N_9734,N_7738,N_7319);
nand U9735 (N_9735,N_8575,N_7041);
and U9736 (N_9736,N_6510,N_8803);
nor U9737 (N_9737,N_8102,N_6159);
nor U9738 (N_9738,N_7669,N_7306);
or U9739 (N_9739,N_7895,N_8750);
nand U9740 (N_9740,N_6126,N_8306);
nor U9741 (N_9741,N_8136,N_8628);
and U9742 (N_9742,N_8576,N_6651);
nor U9743 (N_9743,N_6038,N_8402);
or U9744 (N_9744,N_6579,N_6076);
nand U9745 (N_9745,N_6027,N_6914);
nand U9746 (N_9746,N_7787,N_7946);
or U9747 (N_9747,N_6026,N_8434);
and U9748 (N_9748,N_8191,N_6867);
nand U9749 (N_9749,N_6664,N_6572);
nand U9750 (N_9750,N_8647,N_8724);
nand U9751 (N_9751,N_7693,N_8018);
nor U9752 (N_9752,N_6367,N_7675);
nand U9753 (N_9753,N_7953,N_7710);
and U9754 (N_9754,N_8523,N_8056);
or U9755 (N_9755,N_8513,N_7516);
or U9756 (N_9756,N_8079,N_7349);
or U9757 (N_9757,N_6775,N_6033);
or U9758 (N_9758,N_8788,N_8024);
nor U9759 (N_9759,N_6257,N_6031);
nand U9760 (N_9760,N_8078,N_6908);
nand U9761 (N_9761,N_7515,N_8668);
nand U9762 (N_9762,N_7097,N_6382);
and U9763 (N_9763,N_7522,N_7906);
and U9764 (N_9764,N_6360,N_7555);
and U9765 (N_9765,N_8867,N_8132);
xnor U9766 (N_9766,N_8989,N_7446);
or U9767 (N_9767,N_6003,N_8521);
nand U9768 (N_9768,N_6940,N_6190);
nand U9769 (N_9769,N_6455,N_8826);
nor U9770 (N_9770,N_8293,N_8494);
and U9771 (N_9771,N_6412,N_6758);
and U9772 (N_9772,N_8143,N_7326);
or U9773 (N_9773,N_8625,N_6096);
and U9774 (N_9774,N_6060,N_7086);
nor U9775 (N_9775,N_8578,N_7153);
nor U9776 (N_9776,N_8934,N_8895);
and U9777 (N_9777,N_6439,N_6473);
or U9778 (N_9778,N_6744,N_6656);
and U9779 (N_9779,N_6189,N_7542);
and U9780 (N_9780,N_8046,N_8702);
nand U9781 (N_9781,N_6500,N_7841);
and U9782 (N_9782,N_8250,N_8887);
nand U9783 (N_9783,N_6866,N_6433);
nor U9784 (N_9784,N_8615,N_7094);
or U9785 (N_9785,N_8396,N_7632);
or U9786 (N_9786,N_8211,N_7482);
or U9787 (N_9787,N_8992,N_8525);
nor U9788 (N_9788,N_7893,N_7996);
nand U9789 (N_9789,N_7228,N_6306);
nand U9790 (N_9790,N_8569,N_7008);
or U9791 (N_9791,N_8234,N_8062);
nand U9792 (N_9792,N_8093,N_8975);
nand U9793 (N_9793,N_7085,N_8692);
nor U9794 (N_9794,N_6915,N_6652);
or U9795 (N_9795,N_6504,N_6570);
and U9796 (N_9796,N_6294,N_6526);
nor U9797 (N_9797,N_8994,N_8082);
nor U9798 (N_9798,N_7941,N_7716);
or U9799 (N_9799,N_7003,N_8366);
or U9800 (N_9800,N_6697,N_8907);
and U9801 (N_9801,N_6521,N_7595);
and U9802 (N_9802,N_7078,N_7714);
nor U9803 (N_9803,N_7014,N_8065);
or U9804 (N_9804,N_8187,N_6623);
xor U9805 (N_9805,N_6310,N_8144);
and U9806 (N_9806,N_6470,N_6603);
or U9807 (N_9807,N_8021,N_6771);
or U9808 (N_9808,N_8637,N_7287);
and U9809 (N_9809,N_8818,N_7777);
nor U9810 (N_9810,N_6624,N_8439);
nor U9811 (N_9811,N_7026,N_6828);
or U9812 (N_9812,N_7907,N_7464);
and U9813 (N_9813,N_8609,N_7140);
nor U9814 (N_9814,N_8232,N_7403);
and U9815 (N_9815,N_6749,N_6499);
nand U9816 (N_9816,N_8654,N_7428);
nand U9817 (N_9817,N_8035,N_7096);
nor U9818 (N_9818,N_8074,N_7305);
nor U9819 (N_9819,N_8326,N_7347);
nand U9820 (N_9820,N_8995,N_6574);
or U9821 (N_9821,N_7360,N_8927);
nor U9822 (N_9822,N_7511,N_8089);
nand U9823 (N_9823,N_6713,N_6565);
or U9824 (N_9824,N_6894,N_6627);
nand U9825 (N_9825,N_8031,N_7131);
nor U9826 (N_9826,N_8008,N_6933);
and U9827 (N_9827,N_6636,N_6818);
and U9828 (N_9828,N_7699,N_6674);
nor U9829 (N_9829,N_6661,N_7091);
or U9830 (N_9830,N_7688,N_8140);
nor U9831 (N_9831,N_6101,N_8588);
nor U9832 (N_9832,N_8106,N_8721);
nand U9833 (N_9833,N_6843,N_7185);
nand U9834 (N_9834,N_8857,N_8321);
nor U9835 (N_9835,N_6083,N_6137);
nor U9836 (N_9836,N_6048,N_7240);
nor U9837 (N_9837,N_7022,N_8455);
nor U9838 (N_9838,N_8932,N_6514);
xnor U9839 (N_9839,N_8490,N_6823);
nor U9840 (N_9840,N_8511,N_7147);
nor U9841 (N_9841,N_6184,N_6005);
nand U9842 (N_9842,N_8220,N_6407);
and U9843 (N_9843,N_6292,N_6588);
and U9844 (N_9844,N_7703,N_6880);
nor U9845 (N_9845,N_7633,N_8389);
and U9846 (N_9846,N_6747,N_6756);
nor U9847 (N_9847,N_8520,N_6913);
xnor U9848 (N_9848,N_8514,N_8496);
nor U9849 (N_9849,N_7810,N_7030);
or U9850 (N_9850,N_6787,N_8680);
and U9851 (N_9851,N_7909,N_6321);
nand U9852 (N_9852,N_8003,N_8621);
and U9853 (N_9853,N_8038,N_7197);
and U9854 (N_9854,N_7886,N_8705);
nor U9855 (N_9855,N_6872,N_8122);
and U9856 (N_9856,N_7715,N_7455);
xnor U9857 (N_9857,N_7232,N_7188);
and U9858 (N_9858,N_8479,N_8026);
and U9859 (N_9859,N_6491,N_6320);
nand U9860 (N_9860,N_8541,N_8928);
nand U9861 (N_9861,N_6014,N_6567);
nand U9862 (N_9862,N_7394,N_6278);
or U9863 (N_9863,N_8180,N_7533);
or U9864 (N_9864,N_6025,N_6991);
nand U9865 (N_9865,N_8130,N_6893);
nand U9866 (N_9866,N_8474,N_6369);
or U9867 (N_9867,N_8193,N_6884);
nand U9868 (N_9868,N_8645,N_7902);
and U9869 (N_9869,N_7768,N_8351);
or U9870 (N_9870,N_7090,N_6587);
or U9871 (N_9871,N_8267,N_6589);
or U9872 (N_9872,N_6709,N_7011);
or U9873 (N_9873,N_8701,N_7473);
nor U9874 (N_9874,N_6904,N_6878);
nor U9875 (N_9875,N_6975,N_8073);
or U9876 (N_9876,N_7221,N_6220);
or U9877 (N_9877,N_8644,N_8344);
nand U9878 (N_9878,N_7527,N_8072);
nand U9879 (N_9879,N_7037,N_8275);
and U9880 (N_9880,N_8558,N_7821);
or U9881 (N_9881,N_7892,N_6830);
nor U9882 (N_9882,N_8923,N_7940);
or U9883 (N_9883,N_7493,N_6687);
nor U9884 (N_9884,N_6927,N_7265);
nand U9885 (N_9885,N_8355,N_8969);
nand U9886 (N_9886,N_8071,N_7133);
or U9887 (N_9887,N_6045,N_6966);
and U9888 (N_9888,N_7005,N_8662);
nand U9889 (N_9889,N_6767,N_8653);
nand U9890 (N_9890,N_8380,N_7484);
nor U9891 (N_9891,N_6431,N_7323);
nor U9892 (N_9892,N_8999,N_8847);
nand U9893 (N_9893,N_6377,N_8272);
nand U9894 (N_9894,N_6617,N_7177);
or U9895 (N_9895,N_7396,N_6520);
nand U9896 (N_9896,N_7637,N_6417);
nor U9897 (N_9897,N_8599,N_6755);
nor U9898 (N_9898,N_7467,N_7387);
and U9899 (N_9899,N_7448,N_8802);
or U9900 (N_9900,N_7035,N_6985);
nand U9901 (N_9901,N_8027,N_8280);
nor U9902 (N_9902,N_8361,N_7758);
or U9903 (N_9903,N_8121,N_6350);
or U9904 (N_9904,N_8268,N_7250);
nand U9905 (N_9905,N_8171,N_7032);
nor U9906 (N_9906,N_7064,N_6857);
and U9907 (N_9907,N_8535,N_8981);
nor U9908 (N_9908,N_7903,N_7631);
and U9909 (N_9909,N_8626,N_6129);
or U9910 (N_9910,N_7995,N_8503);
and U9911 (N_9911,N_6256,N_6681);
nand U9912 (N_9912,N_7172,N_6640);
and U9913 (N_9913,N_6973,N_7931);
nor U9914 (N_9914,N_8764,N_7028);
or U9915 (N_9915,N_7488,N_7966);
or U9916 (N_9916,N_8088,N_8037);
nor U9917 (N_9917,N_8893,N_7702);
nand U9918 (N_9918,N_6923,N_7870);
and U9919 (N_9919,N_6450,N_8562);
nand U9920 (N_9920,N_8616,N_8273);
nor U9921 (N_9921,N_6759,N_6964);
nor U9922 (N_9922,N_8715,N_8720);
nor U9923 (N_9923,N_6537,N_6618);
nor U9924 (N_9924,N_8768,N_6719);
nor U9925 (N_9925,N_8795,N_7332);
or U9926 (N_9926,N_6929,N_8566);
nand U9927 (N_9927,N_6080,N_8916);
and U9928 (N_9928,N_7381,N_7371);
nand U9929 (N_9929,N_7567,N_7069);
nor U9930 (N_9930,N_7063,N_8706);
nand U9931 (N_9931,N_7422,N_8755);
nand U9932 (N_9932,N_6172,N_6943);
and U9933 (N_9933,N_6138,N_6365);
or U9934 (N_9934,N_7991,N_7495);
or U9935 (N_9935,N_7006,N_7211);
and U9936 (N_9936,N_8561,N_8157);
and U9937 (N_9937,N_6757,N_7025);
or U9938 (N_9938,N_8565,N_7377);
and U9939 (N_9939,N_6946,N_6862);
nand U9940 (N_9940,N_7615,N_6267);
nor U9941 (N_9941,N_8428,N_7736);
nor U9942 (N_9942,N_7838,N_8635);
or U9943 (N_9943,N_6199,N_7339);
nand U9944 (N_9944,N_8564,N_6969);
nor U9945 (N_9945,N_8781,N_6484);
nand U9946 (N_9946,N_8001,N_6788);
nor U9947 (N_9947,N_8440,N_7109);
or U9948 (N_9948,N_8390,N_6575);
or U9949 (N_9949,N_6006,N_6194);
nand U9950 (N_9950,N_6836,N_8674);
nand U9951 (N_9951,N_7689,N_7215);
nor U9952 (N_9952,N_7115,N_8917);
and U9953 (N_9953,N_8392,N_7194);
nor U9954 (N_9954,N_6164,N_6094);
and U9955 (N_9955,N_6171,N_6281);
or U9956 (N_9956,N_7080,N_8679);
nor U9957 (N_9957,N_7653,N_6488);
nor U9958 (N_9958,N_6234,N_6207);
or U9959 (N_9959,N_8736,N_8811);
or U9960 (N_9960,N_7657,N_6260);
nor U9961 (N_9961,N_7610,N_6779);
and U9962 (N_9962,N_7735,N_7234);
nor U9963 (N_9963,N_8582,N_6300);
nor U9964 (N_9964,N_8695,N_6188);
or U9965 (N_9965,N_7680,N_8353);
nor U9966 (N_9966,N_8329,N_6146);
nor U9967 (N_9967,N_7142,N_8231);
or U9968 (N_9968,N_6053,N_6162);
nor U9969 (N_9969,N_6765,N_7857);
nand U9970 (N_9970,N_7884,N_8343);
and U9971 (N_9971,N_7374,N_7950);
and U9972 (N_9972,N_6899,N_8732);
nand U9973 (N_9973,N_6429,N_8456);
nor U9974 (N_9974,N_7504,N_6248);
and U9975 (N_9975,N_8956,N_7647);
nand U9976 (N_9976,N_8185,N_7815);
nand U9977 (N_9977,N_7811,N_6593);
nand U9978 (N_9978,N_8263,N_8905);
or U9979 (N_9979,N_7936,N_8069);
nand U9980 (N_9980,N_6809,N_6425);
nand U9981 (N_9981,N_8151,N_7257);
nor U9982 (N_9982,N_7002,N_7341);
and U9983 (N_9983,N_6015,N_8844);
nand U9984 (N_9984,N_6989,N_6049);
nor U9985 (N_9985,N_6645,N_6334);
nor U9986 (N_9986,N_6675,N_7110);
or U9987 (N_9987,N_6761,N_6534);
or U9988 (N_9988,N_8935,N_8933);
and U9989 (N_9989,N_6938,N_6206);
xnor U9990 (N_9990,N_6740,N_6062);
and U9991 (N_9991,N_8940,N_8119);
or U9992 (N_9992,N_7762,N_8530);
or U9993 (N_9993,N_6203,N_6870);
or U9994 (N_9994,N_7989,N_6814);
nand U9995 (N_9995,N_6293,N_7746);
nor U9996 (N_9996,N_6561,N_8872);
nand U9997 (N_9997,N_8572,N_8909);
nor U9998 (N_9998,N_7910,N_6827);
or U9999 (N_9999,N_7322,N_8207);
or U10000 (N_10000,N_7487,N_7974);
nor U10001 (N_10001,N_7922,N_8453);
or U10002 (N_10002,N_7912,N_7238);
or U10003 (N_10003,N_7955,N_6167);
or U10004 (N_10004,N_6030,N_8055);
and U10005 (N_10005,N_7642,N_8033);
and U10006 (N_10006,N_7494,N_6523);
or U10007 (N_10007,N_8004,N_7358);
and U10008 (N_10008,N_8452,N_6648);
and U10009 (N_10009,N_7938,N_8712);
or U10010 (N_10010,N_6954,N_6088);
and U10011 (N_10011,N_8540,N_8743);
and U10012 (N_10012,N_8294,N_8131);
and U10013 (N_10013,N_8183,N_7992);
nor U10014 (N_10014,N_6298,N_8815);
or U10015 (N_10015,N_8265,N_7291);
xnor U10016 (N_10016,N_8766,N_7624);
and U10017 (N_10017,N_6835,N_7100);
or U10018 (N_10018,N_6602,N_8696);
and U10019 (N_10019,N_6647,N_7834);
and U10020 (N_10020,N_6811,N_7911);
and U10021 (N_10021,N_7957,N_8259);
nand U10022 (N_10022,N_8689,N_7500);
xor U10023 (N_10023,N_6079,N_8713);
nand U10024 (N_10024,N_8489,N_8481);
and U10025 (N_10025,N_7202,N_7038);
nor U10026 (N_10026,N_7842,N_6123);
and U10027 (N_10027,N_7674,N_8145);
and U10028 (N_10028,N_8338,N_8022);
and U10029 (N_10029,N_7031,N_8960);
nor U10030 (N_10030,N_7255,N_7802);
or U10031 (N_10031,N_7071,N_8773);
nor U10032 (N_10032,N_8583,N_6072);
nor U10033 (N_10033,N_7969,N_8483);
nor U10034 (N_10034,N_6381,N_7535);
and U10035 (N_10035,N_7866,N_7916);
and U10036 (N_10036,N_6808,N_6703);
nor U10037 (N_10037,N_8057,N_8368);
or U10038 (N_10038,N_8733,N_8681);
and U10039 (N_10039,N_6745,N_6873);
nand U10040 (N_10040,N_8404,N_7778);
nand U10041 (N_10041,N_7392,N_7004);
and U10042 (N_10042,N_8308,N_8401);
or U10043 (N_10043,N_8410,N_7449);
nor U10044 (N_10044,N_6525,N_6882);
nor U10045 (N_10045,N_6639,N_6543);
nor U10046 (N_10046,N_7166,N_6115);
and U10047 (N_10047,N_8413,N_6654);
nor U10048 (N_10048,N_6650,N_6492);
or U10049 (N_10049,N_7251,N_6608);
nand U10050 (N_10050,N_6842,N_8797);
nor U10051 (N_10051,N_8438,N_6285);
and U10052 (N_10052,N_7748,N_8816);
and U10053 (N_10053,N_8976,N_7034);
nor U10054 (N_10054,N_8215,N_6128);
nand U10055 (N_10055,N_8601,N_8800);
and U10056 (N_10056,N_6230,N_7000);
nor U10057 (N_10057,N_6854,N_8315);
or U10058 (N_10058,N_8123,N_8789);
nor U10059 (N_10059,N_6770,N_7431);
and U10060 (N_10060,N_8161,N_6804);
nand U10061 (N_10061,N_8210,N_8809);
nor U10062 (N_10062,N_8507,N_8476);
nand U10063 (N_10063,N_6845,N_8487);
or U10064 (N_10064,N_6702,N_6372);
nor U10065 (N_10065,N_6067,N_8086);
nand U10066 (N_10066,N_6924,N_8320);
nor U10067 (N_10067,N_6941,N_6846);
nor U10068 (N_10068,N_7129,N_8342);
nand U10069 (N_10069,N_8958,N_6911);
and U10070 (N_10070,N_8597,N_8869);
or U10071 (N_10071,N_7678,N_8819);
nor U10072 (N_10072,N_7337,N_7894);
nand U10073 (N_10073,N_7619,N_6339);
and U10074 (N_10074,N_7027,N_7737);
nor U10075 (N_10075,N_6011,N_6318);
nand U10076 (N_10076,N_8049,N_7314);
nor U10077 (N_10077,N_8974,N_7728);
and U10078 (N_10078,N_8296,N_8155);
nand U10079 (N_10079,N_8775,N_8243);
nor U10080 (N_10080,N_6685,N_8449);
nor U10081 (N_10081,N_7249,N_8688);
or U10082 (N_10082,N_8497,N_8025);
or U10083 (N_10083,N_8925,N_6819);
nor U10084 (N_10084,N_6376,N_8305);
nand U10085 (N_10085,N_6826,N_8526);
and U10086 (N_10086,N_8400,N_6124);
nand U10087 (N_10087,N_7727,N_6258);
nand U10088 (N_10088,N_7630,N_8176);
nand U10089 (N_10089,N_6531,N_6784);
and U10090 (N_10090,N_7426,N_8300);
and U10091 (N_10091,N_6984,N_6221);
nor U10092 (N_10092,N_7320,N_8875);
and U10093 (N_10093,N_6995,N_6825);
and U10094 (N_10094,N_7127,N_6313);
and U10095 (N_10095,N_6982,N_7293);
or U10096 (N_10096,N_8648,N_7754);
or U10097 (N_10097,N_7210,N_6448);
nor U10098 (N_10098,N_6447,N_6437);
and U10099 (N_10099,N_8728,N_7648);
or U10100 (N_10100,N_7862,N_7150);
nor U10101 (N_10101,N_7840,N_6409);
nand U10102 (N_10102,N_7308,N_8116);
nand U10103 (N_10103,N_7968,N_7574);
or U10104 (N_10104,N_6023,N_7145);
nand U10105 (N_10105,N_7952,N_8812);
xnor U10106 (N_10106,N_6040,N_7442);
and U10107 (N_10107,N_6465,N_7318);
or U10108 (N_10108,N_7345,N_6803);
xor U10109 (N_10109,N_7944,N_8217);
and U10110 (N_10110,N_6573,N_6743);
nand U10111 (N_10111,N_6511,N_8150);
or U10112 (N_10112,N_7990,N_6677);
nor U10113 (N_10113,N_8087,N_8863);
nand U10114 (N_10114,N_7459,N_6580);
nand U10115 (N_10115,N_6239,N_6963);
nand U10116 (N_10116,N_8604,N_6797);
nand U10117 (N_10117,N_8559,N_6752);
and U10118 (N_10118,N_8912,N_8614);
or U10119 (N_10119,N_6082,N_7932);
or U10120 (N_10120,N_8942,N_8084);
nor U10121 (N_10121,N_6855,N_8754);
nor U10122 (N_10122,N_8446,N_8982);
nor U10123 (N_10123,N_7690,N_7545);
nand U10124 (N_10124,N_7092,N_6769);
or U10125 (N_10125,N_8657,N_8962);
or U10126 (N_10126,N_7733,N_6028);
and U10127 (N_10127,N_8360,N_6901);
nand U10128 (N_10128,N_6576,N_7734);
nand U10129 (N_10129,N_6700,N_7800);
or U10130 (N_10130,N_7463,N_6635);
nand U10131 (N_10131,N_6457,N_7451);
xor U10132 (N_10132,N_8047,N_6949);
or U10133 (N_10133,N_7677,N_6119);
nor U10134 (N_10134,N_6024,N_7614);
nand U10135 (N_10135,N_8886,N_8603);
or U10136 (N_10136,N_7724,N_7205);
nor U10137 (N_10137,N_6763,N_6041);
nand U10138 (N_10138,N_6493,N_8179);
and U10139 (N_10139,N_6095,N_6296);
and U10140 (N_10140,N_6790,N_7273);
and U10141 (N_10141,N_8640,N_6528);
nand U10142 (N_10142,N_8415,N_8447);
or U10143 (N_10143,N_7164,N_6348);
or U10144 (N_10144,N_7956,N_6415);
or U10145 (N_10145,N_7982,N_6341);
or U10146 (N_10146,N_8394,N_6413);
and U10147 (N_10147,N_7217,N_6981);
nand U10148 (N_10148,N_6345,N_8617);
and U10149 (N_10149,N_7048,N_7192);
nand U10150 (N_10150,N_8665,N_6246);
and U10151 (N_10151,N_6408,N_8771);
and U10152 (N_10152,N_7340,N_8484);
or U10153 (N_10153,N_8138,N_6953);
nor U10154 (N_10154,N_6614,N_6090);
or U10155 (N_10155,N_7203,N_8634);
nor U10156 (N_10156,N_7262,N_8356);
or U10157 (N_10157,N_7075,N_6330);
nand U10158 (N_10158,N_6979,N_6533);
nor U10159 (N_10159,N_6370,N_6196);
nor U10160 (N_10160,N_8810,N_8406);
or U10161 (N_10161,N_8303,N_7125);
and U10162 (N_10162,N_6071,N_7073);
nand U10163 (N_10163,N_7600,N_8758);
nand U10164 (N_10164,N_6385,N_7123);
or U10165 (N_10165,N_6708,N_6764);
xnor U10166 (N_10166,N_8756,N_7440);
nor U10167 (N_10167,N_7831,N_8574);
or U10168 (N_10168,N_7544,N_8177);
and U10169 (N_10169,N_8411,N_8186);
and U10170 (N_10170,N_8209,N_6279);
and U10171 (N_10171,N_6352,N_6243);
nor U10172 (N_10172,N_7359,N_8194);
and U10173 (N_10173,N_8009,N_8467);
nor U10174 (N_10174,N_8704,N_7526);
nand U10175 (N_10175,N_7761,N_6173);
or U10176 (N_10176,N_6925,N_6668);
nand U10177 (N_10177,N_6177,N_6918);
nor U10178 (N_10178,N_7593,N_8899);
and U10179 (N_10179,N_8742,N_8393);
and U10180 (N_10180,N_8466,N_7881);
nor U10181 (N_10181,N_8216,N_6916);
nor U10182 (N_10182,N_7823,N_8655);
nand U10183 (N_10183,N_7977,N_8804);
and U10184 (N_10184,N_8432,N_8384);
or U10185 (N_10185,N_6403,N_7499);
and U10186 (N_10186,N_8269,N_7058);
and U10187 (N_10187,N_8889,N_7565);
or U10188 (N_10188,N_7837,N_6967);
nor U10189 (N_10189,N_7829,N_7971);
nand U10190 (N_10190,N_7921,N_7718);
nand U10191 (N_10191,N_8206,N_7435);
and U10192 (N_10192,N_8094,N_8596);
or U10193 (N_10193,N_8189,N_7416);
and U10194 (N_10194,N_6261,N_6452);
nor U10195 (N_10195,N_6390,N_6032);
or U10196 (N_10196,N_6798,N_7617);
or U10197 (N_10197,N_6774,N_7313);
or U10198 (N_10198,N_8502,N_8968);
and U10199 (N_10199,N_7687,N_6559);
nand U10200 (N_10200,N_6091,N_7571);
nor U10201 (N_10201,N_8468,N_8882);
nand U10202 (N_10202,N_7354,N_7904);
nor U10203 (N_10203,N_8669,N_7143);
and U10204 (N_10204,N_7609,N_7732);
nor U10205 (N_10205,N_8369,N_7985);
nand U10206 (N_10206,N_8383,N_6271);
nand U10207 (N_10207,N_6712,N_7169);
and U10208 (N_10208,N_7590,N_8594);
nand U10209 (N_10209,N_6148,N_7072);
nor U10210 (N_10210,N_8845,N_7589);
nor U10211 (N_10211,N_6948,N_7634);
nor U10212 (N_10212,N_7612,N_7378);
nor U10213 (N_10213,N_7611,N_8271);
and U10214 (N_10214,N_6114,N_7820);
nand U10215 (N_10215,N_8926,N_6420);
nor U10216 (N_10216,N_6883,N_6936);
nand U10217 (N_10217,N_6625,N_8879);
or U10218 (N_10218,N_8371,N_8311);
or U10219 (N_10219,N_6224,N_7043);
nand U10220 (N_10220,N_8332,N_7686);
nand U10221 (N_10221,N_7017,N_6387);
and U10222 (N_10222,N_6343,N_6998);
nor U10223 (N_10223,N_8226,N_7191);
nand U10224 (N_10224,N_8725,N_7183);
or U10225 (N_10225,N_7290,N_6140);
nor U10226 (N_10226,N_8041,N_7213);
nand U10227 (N_10227,N_6143,N_7130);
or U10228 (N_10228,N_6326,N_8835);
and U10229 (N_10229,N_6853,N_7237);
nor U10230 (N_10230,N_7949,N_6977);
nor U10231 (N_10231,N_6571,N_6477);
nand U10232 (N_10232,N_8436,N_7289);
or U10233 (N_10233,N_8990,N_6380);
nand U10234 (N_10234,N_7836,N_6495);
nor U10235 (N_10235,N_6696,N_6016);
nand U10236 (N_10236,N_8798,N_7353);
nand U10237 (N_10237,N_6251,N_7295);
or U10238 (N_10238,N_8224,N_8537);
nand U10239 (N_10239,N_6536,N_6562);
and U10240 (N_10240,N_6522,N_6594);
or U10241 (N_10241,N_7783,N_6820);
nand U10242 (N_10242,N_7477,N_7742);
or U10243 (N_10243,N_7475,N_7789);
and U10244 (N_10244,N_6386,N_7794);
and U10245 (N_10245,N_7847,N_6606);
or U10246 (N_10246,N_6607,N_8429);
and U10247 (N_10247,N_7173,N_6085);
or U10248 (N_10248,N_8772,N_6699);
and U10249 (N_10249,N_6643,N_7361);
nor U10250 (N_10250,N_6264,N_7849);
nor U10251 (N_10251,N_8229,N_7376);
and U10252 (N_10252,N_8552,N_6942);
nor U10253 (N_10253,N_6289,N_6104);
and U10254 (N_10254,N_8563,N_7068);
nand U10255 (N_10255,N_8471,N_6683);
and U10256 (N_10256,N_6781,N_6092);
nor U10257 (N_10257,N_6609,N_8117);
and U10258 (N_10258,N_7329,N_8373);
nand U10259 (N_10259,N_8786,N_8814);
and U10260 (N_10260,N_7917,N_6195);
nor U10261 (N_10261,N_8671,N_8820);
and U10262 (N_10262,N_6503,N_7899);
nor U10263 (N_10263,N_7658,N_7175);
and U10264 (N_10264,N_8852,N_8316);
nand U10265 (N_10265,N_8700,N_7756);
or U10266 (N_10266,N_7486,N_6216);
or U10267 (N_10267,N_7550,N_8890);
or U10268 (N_10268,N_6034,N_8979);
or U10269 (N_10269,N_8076,N_8931);
nor U10270 (N_10270,N_7743,N_6773);
nor U10271 (N_10271,N_8862,N_6245);
or U10272 (N_10272,N_8950,N_8307);
or U10273 (N_10273,N_8864,N_6553);
and U10274 (N_10274,N_6686,N_7124);
or U10275 (N_10275,N_7889,N_6185);
nor U10276 (N_10276,N_8894,N_7444);
or U10277 (N_10277,N_7553,N_6432);
and U10278 (N_10278,N_7627,N_7021);
or U10279 (N_10279,N_8744,N_7514);
nor U10280 (N_10280,N_6569,N_8370);
nand U10281 (N_10281,N_8060,N_6869);
and U10282 (N_10282,N_8154,N_6689);
or U10283 (N_10283,N_6613,N_8067);
or U10284 (N_10284,N_7963,N_6460);
nand U10285 (N_10285,N_7852,N_8745);
xnor U10286 (N_10286,N_8685,N_7223);
nand U10287 (N_10287,N_7201,N_6287);
nand U10288 (N_10288,N_6782,N_8029);
or U10289 (N_10289,N_8553,N_6902);
nand U10290 (N_10290,N_6517,N_7543);
nand U10291 (N_10291,N_8892,N_8286);
nand U10292 (N_10292,N_8421,N_8821);
and U10293 (N_10293,N_8623,N_8492);
and U10294 (N_10294,N_6274,N_6286);
nand U10295 (N_10295,N_7598,N_6057);
and U10296 (N_10296,N_6688,N_8944);
nand U10297 (N_10297,N_8173,N_7867);
nand U10298 (N_10298,N_8955,N_8478);
nand U10299 (N_10299,N_8780,N_7766);
or U10300 (N_10300,N_7809,N_7998);
nand U10301 (N_10301,N_6059,N_6411);
nor U10302 (N_10302,N_8050,N_7552);
nor U10303 (N_10303,N_7760,N_7607);
nand U10304 (N_10304,N_8340,N_6555);
xnor U10305 (N_10305,N_6254,N_7454);
and U10306 (N_10306,N_7423,N_6794);
nand U10307 (N_10307,N_7083,N_8015);
or U10308 (N_10308,N_7274,N_7826);
or U10309 (N_10309,N_7701,N_8365);
nand U10310 (N_10310,N_6154,N_7243);
nor U10311 (N_10311,N_8896,N_6508);
nor U10312 (N_10312,N_7622,N_6222);
nand U10313 (N_10313,N_7065,N_6443);
nand U10314 (N_10314,N_7755,N_8904);
and U10315 (N_10315,N_7915,N_7334);
nor U10316 (N_10316,N_6461,N_7696);
and U10317 (N_10317,N_8834,N_8416);
and U10318 (N_10318,N_8592,N_6210);
and U10319 (N_10319,N_6247,N_6160);
or U10320 (N_10320,N_6671,N_6240);
or U10321 (N_10321,N_7643,N_8843);
and U10322 (N_10322,N_7226,N_6169);
nor U10323 (N_10323,N_8726,N_8877);
nor U10324 (N_10324,N_6881,N_8580);
and U10325 (N_10325,N_6619,N_7383);
and U10326 (N_10326,N_6628,N_7601);
and U10327 (N_10327,N_7804,N_8011);
nor U10328 (N_10328,N_8252,N_6404);
nor U10329 (N_10329,N_6226,N_6388);
nand U10330 (N_10330,N_8524,N_8334);
nor U10331 (N_10331,N_6850,N_8579);
nor U10332 (N_10332,N_7116,N_6481);
nor U10333 (N_10333,N_7740,N_7180);
or U10334 (N_10334,N_8509,N_7263);
nor U10335 (N_10335,N_7578,N_6295);
nand U10336 (N_10336,N_8871,N_7785);
and U10337 (N_10337,N_6582,N_7608);
nand U10338 (N_10338,N_8405,N_8139);
nor U10339 (N_10339,N_7531,N_7770);
and U10340 (N_10340,N_7266,N_7382);
nor U10341 (N_10341,N_7745,N_7066);
nand U10342 (N_10342,N_8996,N_8281);
and U10343 (N_10343,N_6422,N_6242);
nand U10344 (N_10344,N_7697,N_7149);
nor U10345 (N_10345,N_8482,N_6754);
nand U10346 (N_10346,N_8658,N_7919);
nor U10347 (N_10347,N_7948,N_6487);
nor U10348 (N_10348,N_7554,N_6637);
nor U10349 (N_10349,N_6540,N_7105);
nand U10350 (N_10350,N_7597,N_7352);
and U10351 (N_10351,N_8930,N_8908);
nor U10352 (N_10352,N_6695,N_7671);
or U10353 (N_10353,N_6394,N_6513);
or U10354 (N_10354,N_8398,N_7524);
or U10355 (N_10355,N_7389,N_8885);
or U10356 (N_10356,N_8573,N_8425);
nor U10357 (N_10357,N_7054,N_7239);
nand U10358 (N_10358,N_6472,N_8289);
nand U10359 (N_10359,N_8081,N_8358);
nor U10360 (N_10360,N_6156,N_6157);
and U10361 (N_10361,N_8357,N_7773);
and U10362 (N_10362,N_8258,N_8661);
nand U10363 (N_10363,N_7146,N_8058);
nor U10364 (N_10364,N_7850,N_7914);
nor U10365 (N_10365,N_7427,N_8433);
and U10366 (N_10366,N_7040,N_6175);
or U10367 (N_10367,N_6591,N_6359);
or U10368 (N_10368,N_7572,N_6959);
and U10369 (N_10369,N_7588,N_8888);
and U10370 (N_10370,N_6768,N_6338);
and U10371 (N_10371,N_8529,N_7776);
nand U10372 (N_10372,N_7108,N_7937);
nand U10373 (N_10373,N_6105,N_7629);
nor U10374 (N_10374,N_8085,N_8778);
nor U10375 (N_10375,N_6807,N_7307);
and U10376 (N_10376,N_7288,N_6780);
nand U10377 (N_10377,N_8097,N_7517);
or U10378 (N_10378,N_8285,N_7749);
nand U10379 (N_10379,N_8697,N_8499);
and U10380 (N_10380,N_7623,N_6314);
nand U10381 (N_10381,N_8638,N_8849);
nor U10382 (N_10382,N_6299,N_7104);
xnor U10383 (N_10383,N_7385,N_8939);
or U10384 (N_10384,N_6909,N_6252);
or U10385 (N_10385,N_7786,N_7692);
or U10386 (N_10386,N_6595,N_6150);
and U10387 (N_10387,N_7930,N_6426);
or U10388 (N_10388,N_7039,N_7519);
or U10389 (N_10389,N_7112,N_7548);
nand U10390 (N_10390,N_6766,N_6711);
nand U10391 (N_10391,N_8409,N_8457);
nor U10392 (N_10392,N_6679,N_6498);
nand U10393 (N_10393,N_6284,N_8454);
nand U10394 (N_10394,N_7659,N_8167);
and U10395 (N_10395,N_8288,N_8624);
nor U10396 (N_10396,N_6197,N_7103);
nor U10397 (N_10397,N_6141,N_7566);
nand U10398 (N_10398,N_6910,N_6174);
and U10399 (N_10399,N_8900,N_8324);
nor U10400 (N_10400,N_6676,N_8152);
nand U10401 (N_10401,N_6672,N_6693);
and U10402 (N_10402,N_8633,N_7253);
and U10403 (N_10403,N_7220,N_6535);
or U10404 (N_10404,N_6800,N_8949);
and U10405 (N_10405,N_7407,N_6852);
or U10406 (N_10406,N_8517,N_7241);
nor U10407 (N_10407,N_8444,N_7663);
and U10408 (N_10408,N_8547,N_8951);
nand U10409 (N_10409,N_7603,N_7618);
and U10410 (N_10410,N_6707,N_7859);
nor U10411 (N_10411,N_6019,N_6847);
and U10412 (N_10412,N_6772,N_6198);
nor U10413 (N_10413,N_6149,N_6307);
nand U10414 (N_10414,N_7905,N_8399);
and U10415 (N_10415,N_8991,N_6351);
nand U10416 (N_10416,N_8230,N_8485);
nand U10417 (N_10417,N_7375,N_7061);
or U10418 (N_10418,N_7602,N_7649);
nand U10419 (N_10419,N_6871,N_7518);
nor U10420 (N_10420,N_7868,N_8124);
nor U10421 (N_10421,N_7012,N_8309);
and U10422 (N_10422,N_8387,N_7920);
nor U10423 (N_10423,N_8264,N_7568);
nor U10424 (N_10424,N_8774,N_8223);
and U10425 (N_10425,N_7816,N_7596);
and U10426 (N_10426,N_6907,N_7139);
nand U10427 (N_10427,N_6988,N_8111);
and U10428 (N_10428,N_7317,N_6960);
nand U10429 (N_10429,N_7055,N_6506);
nand U10430 (N_10430,N_7138,N_6131);
or U10431 (N_10431,N_7060,N_8044);
nand U10432 (N_10432,N_6926,N_7767);
nor U10433 (N_10433,N_7010,N_7858);
and U10434 (N_10434,N_6236,N_8459);
nor U10435 (N_10435,N_6202,N_6263);
nor U10436 (N_10436,N_6538,N_7224);
nor U10437 (N_10437,N_6947,N_6181);
or U10438 (N_10438,N_7402,N_8372);
nor U10439 (N_10439,N_6931,N_7016);
or U10440 (N_10440,N_7466,N_8817);
or U10441 (N_10441,N_7757,N_8397);
and U10442 (N_10442,N_7707,N_8512);
nand U10443 (N_10443,N_8751,N_8430);
nor U10444 (N_10444,N_8341,N_6566);
nand U10445 (N_10445,N_8876,N_6399);
nor U10446 (N_10446,N_6001,N_6304);
or U10447 (N_10447,N_7997,N_6204);
or U10448 (N_10448,N_8868,N_7556);
nand U10449 (N_10449,N_6276,N_7236);
or U10450 (N_10450,N_8110,N_7336);
nor U10451 (N_10451,N_6316,N_7101);
nand U10452 (N_10452,N_6726,N_7272);
or U10453 (N_10453,N_6042,N_6563);
nand U10454 (N_10454,N_6813,N_6649);
nor U10455 (N_10455,N_8606,N_6507);
nand U10456 (N_10456,N_8066,N_7079);
or U10457 (N_10457,N_7855,N_6458);
nor U10458 (N_10458,N_6102,N_8395);
nor U10459 (N_10459,N_7412,N_7654);
nor U10460 (N_10460,N_8158,N_8470);
or U10461 (N_10461,N_7885,N_6444);
or U10462 (N_10462,N_6838,N_6208);
nand U10463 (N_10463,N_8881,N_6682);
and U10464 (N_10464,N_8039,N_8865);
nor U10465 (N_10465,N_8445,N_6397);
nor U10466 (N_10466,N_7258,N_6373);
or U10467 (N_10467,N_6976,N_8451);
or U10468 (N_10468,N_8034,N_7348);
nor U10469 (N_10469,N_8407,N_8998);
or U10470 (N_10470,N_7148,N_6127);
or U10471 (N_10471,N_6622,N_6983);
and U10472 (N_10472,N_8064,N_8103);
or U10473 (N_10473,N_7269,N_6644);
and U10474 (N_10474,N_7537,N_7529);
nor U10475 (N_10475,N_8548,N_7436);
or U10476 (N_10476,N_7807,N_6002);
or U10477 (N_10477,N_6952,N_8910);
and U10478 (N_10478,N_6428,N_7196);
xor U10479 (N_10479,N_8952,N_6547);
nand U10480 (N_10480,N_7438,N_7388);
nor U10481 (N_10481,N_6480,N_8346);
nor U10482 (N_10482,N_6086,N_8752);
or U10483 (N_10483,N_7528,N_7415);
nand U10484 (N_10484,N_8891,N_7661);
nand U10485 (N_10485,N_6629,N_6191);
or U10486 (N_10486,N_6971,N_7784);
or U10487 (N_10487,N_7591,N_6680);
nor U10488 (N_10488,N_6833,N_7559);
nor U10489 (N_10489,N_7181,N_7681);
nor U10490 (N_10490,N_8319,N_7875);
or U10491 (N_10491,N_8510,N_6333);
and U10492 (N_10492,N_6055,N_7433);
or U10493 (N_10493,N_6921,N_8984);
nor U10494 (N_10494,N_8631,N_7470);
nor U10495 (N_10495,N_6136,N_8169);
and U10496 (N_10496,N_6965,N_7469);
nor U10497 (N_10497,N_8884,N_7134);
and U10498 (N_10498,N_8337,N_8245);
and U10499 (N_10499,N_6583,N_8166);
or U10500 (N_10500,N_6113,N_8411);
or U10501 (N_10501,N_6081,N_6385);
nand U10502 (N_10502,N_6126,N_6435);
and U10503 (N_10503,N_6225,N_6084);
nand U10504 (N_10504,N_6413,N_6432);
nand U10505 (N_10505,N_6290,N_8828);
and U10506 (N_10506,N_8511,N_7236);
nor U10507 (N_10507,N_7500,N_6577);
nor U10508 (N_10508,N_6003,N_8106);
nand U10509 (N_10509,N_8583,N_8219);
nor U10510 (N_10510,N_6919,N_6761);
or U10511 (N_10511,N_7370,N_6435);
nor U10512 (N_10512,N_7880,N_8140);
nor U10513 (N_10513,N_7745,N_7346);
or U10514 (N_10514,N_6695,N_7904);
nor U10515 (N_10515,N_7069,N_7427);
or U10516 (N_10516,N_6682,N_8742);
or U10517 (N_10517,N_8309,N_8635);
or U10518 (N_10518,N_6819,N_8463);
and U10519 (N_10519,N_6664,N_8204);
nand U10520 (N_10520,N_8676,N_6862);
and U10521 (N_10521,N_8366,N_7775);
xor U10522 (N_10522,N_8056,N_7629);
nand U10523 (N_10523,N_6914,N_6236);
nor U10524 (N_10524,N_8136,N_6497);
or U10525 (N_10525,N_7643,N_6050);
nor U10526 (N_10526,N_8787,N_8816);
nand U10527 (N_10527,N_8570,N_8865);
and U10528 (N_10528,N_8578,N_6396);
and U10529 (N_10529,N_6820,N_8849);
nand U10530 (N_10530,N_8641,N_6375);
nor U10531 (N_10531,N_8632,N_6488);
or U10532 (N_10532,N_8723,N_8752);
xnor U10533 (N_10533,N_6110,N_6142);
and U10534 (N_10534,N_6734,N_8844);
nor U10535 (N_10535,N_8367,N_8028);
nand U10536 (N_10536,N_7732,N_8169);
nand U10537 (N_10537,N_6757,N_6680);
and U10538 (N_10538,N_7038,N_8794);
and U10539 (N_10539,N_8893,N_7750);
and U10540 (N_10540,N_8150,N_8960);
nand U10541 (N_10541,N_8662,N_8952);
or U10542 (N_10542,N_6739,N_8316);
and U10543 (N_10543,N_7091,N_7359);
or U10544 (N_10544,N_6359,N_7127);
and U10545 (N_10545,N_7604,N_7193);
and U10546 (N_10546,N_8829,N_8791);
and U10547 (N_10547,N_6676,N_6554);
nand U10548 (N_10548,N_8773,N_8981);
or U10549 (N_10549,N_8488,N_7696);
or U10550 (N_10550,N_7732,N_8766);
nand U10551 (N_10551,N_7712,N_7098);
nor U10552 (N_10552,N_8087,N_6157);
nor U10553 (N_10553,N_8095,N_8165);
nor U10554 (N_10554,N_6470,N_8905);
and U10555 (N_10555,N_6944,N_7500);
nor U10556 (N_10556,N_7886,N_7574);
or U10557 (N_10557,N_8886,N_6865);
nand U10558 (N_10558,N_6713,N_8667);
nand U10559 (N_10559,N_8652,N_7965);
and U10560 (N_10560,N_7788,N_6837);
nor U10561 (N_10561,N_7877,N_6779);
nand U10562 (N_10562,N_8822,N_8659);
and U10563 (N_10563,N_8062,N_8728);
or U10564 (N_10564,N_8301,N_8607);
nand U10565 (N_10565,N_7616,N_6873);
and U10566 (N_10566,N_8468,N_7922);
nor U10567 (N_10567,N_8575,N_8618);
nor U10568 (N_10568,N_7934,N_6873);
and U10569 (N_10569,N_7734,N_7208);
nand U10570 (N_10570,N_8744,N_6573);
nand U10571 (N_10571,N_8706,N_8110);
nand U10572 (N_10572,N_8478,N_7035);
and U10573 (N_10573,N_8960,N_8745);
or U10574 (N_10574,N_6368,N_6992);
nor U10575 (N_10575,N_8164,N_6885);
or U10576 (N_10576,N_7629,N_7887);
nand U10577 (N_10577,N_8737,N_6666);
nor U10578 (N_10578,N_8744,N_8702);
or U10579 (N_10579,N_7241,N_7650);
nor U10580 (N_10580,N_6538,N_7917);
and U10581 (N_10581,N_6665,N_6880);
or U10582 (N_10582,N_7102,N_8736);
and U10583 (N_10583,N_6832,N_6037);
nor U10584 (N_10584,N_8972,N_8579);
and U10585 (N_10585,N_7728,N_6334);
or U10586 (N_10586,N_8913,N_7537);
nor U10587 (N_10587,N_6966,N_7142);
nor U10588 (N_10588,N_8895,N_6924);
nand U10589 (N_10589,N_7744,N_8156);
nor U10590 (N_10590,N_7620,N_8657);
nand U10591 (N_10591,N_8617,N_7798);
nor U10592 (N_10592,N_8434,N_8658);
nor U10593 (N_10593,N_6811,N_8731);
nand U10594 (N_10594,N_7116,N_6835);
nor U10595 (N_10595,N_8022,N_6963);
nand U10596 (N_10596,N_7720,N_8565);
or U10597 (N_10597,N_8842,N_7122);
and U10598 (N_10598,N_6482,N_6788);
and U10599 (N_10599,N_7902,N_7439);
nand U10600 (N_10600,N_7505,N_7099);
nand U10601 (N_10601,N_6508,N_8642);
or U10602 (N_10602,N_8082,N_7187);
nor U10603 (N_10603,N_7227,N_6693);
nor U10604 (N_10604,N_6157,N_6285);
and U10605 (N_10605,N_8365,N_6758);
nand U10606 (N_10606,N_8485,N_6211);
and U10607 (N_10607,N_8981,N_8640);
or U10608 (N_10608,N_7477,N_7303);
nor U10609 (N_10609,N_6062,N_7905);
or U10610 (N_10610,N_6929,N_6271);
nor U10611 (N_10611,N_6788,N_7782);
nand U10612 (N_10612,N_7394,N_6113);
nor U10613 (N_10613,N_6885,N_7996);
or U10614 (N_10614,N_7470,N_6384);
and U10615 (N_10615,N_7131,N_7683);
nand U10616 (N_10616,N_6402,N_8091);
or U10617 (N_10617,N_6565,N_6515);
or U10618 (N_10618,N_8164,N_7390);
nand U10619 (N_10619,N_8982,N_8760);
nor U10620 (N_10620,N_7923,N_8136);
or U10621 (N_10621,N_6280,N_7019);
and U10622 (N_10622,N_8862,N_7381);
nor U10623 (N_10623,N_6956,N_6957);
or U10624 (N_10624,N_7132,N_6628);
nand U10625 (N_10625,N_7403,N_6432);
nor U10626 (N_10626,N_7217,N_7872);
nand U10627 (N_10627,N_7900,N_6620);
nand U10628 (N_10628,N_7924,N_7657);
and U10629 (N_10629,N_8036,N_7771);
nor U10630 (N_10630,N_6813,N_7152);
nand U10631 (N_10631,N_6099,N_6043);
nor U10632 (N_10632,N_7667,N_8129);
nand U10633 (N_10633,N_6561,N_6488);
nor U10634 (N_10634,N_6214,N_7357);
nor U10635 (N_10635,N_8854,N_8681);
nor U10636 (N_10636,N_8905,N_6767);
xor U10637 (N_10637,N_8004,N_6673);
nor U10638 (N_10638,N_6804,N_8936);
and U10639 (N_10639,N_8419,N_6470);
and U10640 (N_10640,N_8859,N_7621);
and U10641 (N_10641,N_8245,N_6146);
nand U10642 (N_10642,N_6087,N_8458);
nand U10643 (N_10643,N_8665,N_6610);
or U10644 (N_10644,N_8654,N_8928);
or U10645 (N_10645,N_7875,N_6914);
nand U10646 (N_10646,N_7766,N_6077);
nor U10647 (N_10647,N_8272,N_7531);
and U10648 (N_10648,N_6363,N_8130);
and U10649 (N_10649,N_8368,N_7771);
nor U10650 (N_10650,N_7625,N_8421);
nand U10651 (N_10651,N_7277,N_8128);
and U10652 (N_10652,N_6704,N_6462);
xor U10653 (N_10653,N_6945,N_7560);
or U10654 (N_10654,N_8536,N_6447);
nand U10655 (N_10655,N_8679,N_6851);
nor U10656 (N_10656,N_8265,N_7209);
nand U10657 (N_10657,N_6496,N_7291);
nor U10658 (N_10658,N_6196,N_7243);
and U10659 (N_10659,N_8716,N_6275);
and U10660 (N_10660,N_7513,N_7957);
nand U10661 (N_10661,N_7340,N_8215);
nand U10662 (N_10662,N_6508,N_6208);
and U10663 (N_10663,N_6418,N_7489);
or U10664 (N_10664,N_6983,N_7908);
and U10665 (N_10665,N_7264,N_7192);
and U10666 (N_10666,N_8280,N_6007);
and U10667 (N_10667,N_8397,N_8972);
nor U10668 (N_10668,N_7839,N_7831);
and U10669 (N_10669,N_7436,N_6561);
and U10670 (N_10670,N_8260,N_7824);
and U10671 (N_10671,N_7943,N_8147);
nand U10672 (N_10672,N_6838,N_8643);
nor U10673 (N_10673,N_7595,N_6439);
or U10674 (N_10674,N_8232,N_6018);
and U10675 (N_10675,N_7396,N_6100);
nor U10676 (N_10676,N_7945,N_7207);
or U10677 (N_10677,N_8235,N_6017);
and U10678 (N_10678,N_6708,N_6253);
or U10679 (N_10679,N_7840,N_7277);
nor U10680 (N_10680,N_8877,N_6907);
or U10681 (N_10681,N_8574,N_6979);
or U10682 (N_10682,N_8536,N_8743);
nand U10683 (N_10683,N_7521,N_7869);
nor U10684 (N_10684,N_8197,N_8628);
and U10685 (N_10685,N_7890,N_8116);
and U10686 (N_10686,N_6161,N_6328);
nor U10687 (N_10687,N_6361,N_6603);
nor U10688 (N_10688,N_6375,N_7825);
nor U10689 (N_10689,N_8548,N_7974);
nor U10690 (N_10690,N_6139,N_8198);
and U10691 (N_10691,N_6322,N_8358);
and U10692 (N_10692,N_8390,N_8164);
nor U10693 (N_10693,N_6527,N_6364);
or U10694 (N_10694,N_6919,N_7002);
or U10695 (N_10695,N_8403,N_6949);
or U10696 (N_10696,N_6775,N_6478);
nor U10697 (N_10697,N_6139,N_8552);
nor U10698 (N_10698,N_7945,N_6367);
or U10699 (N_10699,N_7370,N_6720);
nand U10700 (N_10700,N_8153,N_7795);
nand U10701 (N_10701,N_6214,N_8238);
nor U10702 (N_10702,N_8151,N_8395);
and U10703 (N_10703,N_6468,N_7017);
or U10704 (N_10704,N_6486,N_6314);
xor U10705 (N_10705,N_8304,N_6114);
and U10706 (N_10706,N_6371,N_6524);
and U10707 (N_10707,N_6357,N_8509);
nand U10708 (N_10708,N_7563,N_8585);
or U10709 (N_10709,N_7350,N_7169);
nor U10710 (N_10710,N_6888,N_8148);
nor U10711 (N_10711,N_8795,N_7217);
nor U10712 (N_10712,N_8207,N_7127);
nor U10713 (N_10713,N_8155,N_6726);
and U10714 (N_10714,N_6136,N_8871);
or U10715 (N_10715,N_6656,N_7129);
xor U10716 (N_10716,N_8732,N_8686);
and U10717 (N_10717,N_8440,N_6161);
and U10718 (N_10718,N_6034,N_7641);
xor U10719 (N_10719,N_6611,N_8227);
and U10720 (N_10720,N_6788,N_6714);
nor U10721 (N_10721,N_6117,N_7643);
and U10722 (N_10722,N_8908,N_7977);
nor U10723 (N_10723,N_8669,N_8195);
nor U10724 (N_10724,N_8865,N_6303);
nand U10725 (N_10725,N_6068,N_7644);
or U10726 (N_10726,N_6579,N_8930);
and U10727 (N_10727,N_7690,N_6566);
or U10728 (N_10728,N_7867,N_8464);
or U10729 (N_10729,N_8810,N_6508);
nor U10730 (N_10730,N_6960,N_8492);
and U10731 (N_10731,N_8742,N_8103);
and U10732 (N_10732,N_8089,N_6341);
nand U10733 (N_10733,N_7078,N_8854);
nand U10734 (N_10734,N_8381,N_6722);
and U10735 (N_10735,N_8474,N_8436);
or U10736 (N_10736,N_6715,N_8019);
or U10737 (N_10737,N_6974,N_8900);
nand U10738 (N_10738,N_8132,N_6353);
and U10739 (N_10739,N_7342,N_8000);
and U10740 (N_10740,N_6691,N_8431);
nand U10741 (N_10741,N_7862,N_6533);
or U10742 (N_10742,N_8245,N_7965);
xor U10743 (N_10743,N_6344,N_7978);
nand U10744 (N_10744,N_8396,N_7468);
or U10745 (N_10745,N_6283,N_7485);
or U10746 (N_10746,N_8059,N_6646);
and U10747 (N_10747,N_6965,N_6068);
or U10748 (N_10748,N_7303,N_8216);
or U10749 (N_10749,N_6277,N_8746);
nor U10750 (N_10750,N_6579,N_6947);
nor U10751 (N_10751,N_7140,N_8903);
and U10752 (N_10752,N_6216,N_7604);
nand U10753 (N_10753,N_6311,N_8415);
nand U10754 (N_10754,N_6054,N_7620);
nand U10755 (N_10755,N_6142,N_7941);
nor U10756 (N_10756,N_8390,N_6738);
and U10757 (N_10757,N_6859,N_6778);
and U10758 (N_10758,N_6040,N_6838);
nand U10759 (N_10759,N_8225,N_7934);
nor U10760 (N_10760,N_8561,N_8615);
nor U10761 (N_10761,N_6967,N_8711);
nand U10762 (N_10762,N_6014,N_7015);
or U10763 (N_10763,N_6285,N_6155);
nand U10764 (N_10764,N_6064,N_8850);
nand U10765 (N_10765,N_8322,N_6795);
and U10766 (N_10766,N_7807,N_7489);
nand U10767 (N_10767,N_6585,N_6972);
nor U10768 (N_10768,N_7304,N_8797);
nand U10769 (N_10769,N_7099,N_7870);
or U10770 (N_10770,N_7043,N_7120);
nand U10771 (N_10771,N_8056,N_7329);
nor U10772 (N_10772,N_8972,N_8679);
nor U10773 (N_10773,N_8997,N_8445);
xor U10774 (N_10774,N_7772,N_6530);
or U10775 (N_10775,N_7484,N_8957);
or U10776 (N_10776,N_8447,N_6148);
nor U10777 (N_10777,N_7278,N_6657);
nand U10778 (N_10778,N_6772,N_8420);
and U10779 (N_10779,N_6118,N_6011);
nand U10780 (N_10780,N_8710,N_6717);
or U10781 (N_10781,N_6868,N_7970);
nor U10782 (N_10782,N_8696,N_8699);
or U10783 (N_10783,N_8024,N_6100);
and U10784 (N_10784,N_6918,N_6943);
nor U10785 (N_10785,N_8711,N_6980);
or U10786 (N_10786,N_7799,N_8575);
or U10787 (N_10787,N_7990,N_7383);
or U10788 (N_10788,N_8582,N_7751);
nand U10789 (N_10789,N_7875,N_7167);
nor U10790 (N_10790,N_7656,N_7253);
nand U10791 (N_10791,N_7000,N_6960);
and U10792 (N_10792,N_7858,N_6604);
nor U10793 (N_10793,N_8364,N_7254);
or U10794 (N_10794,N_6484,N_6186);
nor U10795 (N_10795,N_8725,N_8068);
or U10796 (N_10796,N_6536,N_7695);
nor U10797 (N_10797,N_8154,N_8020);
or U10798 (N_10798,N_7044,N_6711);
nand U10799 (N_10799,N_8570,N_7220);
and U10800 (N_10800,N_8927,N_8619);
nand U10801 (N_10801,N_6906,N_6988);
nand U10802 (N_10802,N_7596,N_8190);
nand U10803 (N_10803,N_7714,N_7376);
nand U10804 (N_10804,N_7592,N_7106);
and U10805 (N_10805,N_6820,N_7552);
or U10806 (N_10806,N_8504,N_6871);
nor U10807 (N_10807,N_6745,N_8778);
and U10808 (N_10808,N_7411,N_7298);
and U10809 (N_10809,N_8103,N_6180);
nand U10810 (N_10810,N_8826,N_7261);
or U10811 (N_10811,N_7397,N_7803);
or U10812 (N_10812,N_6677,N_6139);
nor U10813 (N_10813,N_7297,N_6835);
or U10814 (N_10814,N_6388,N_7092);
nand U10815 (N_10815,N_6729,N_6405);
nand U10816 (N_10816,N_7244,N_8048);
and U10817 (N_10817,N_6410,N_8029);
or U10818 (N_10818,N_7386,N_7446);
nor U10819 (N_10819,N_6493,N_8026);
and U10820 (N_10820,N_6768,N_6545);
or U10821 (N_10821,N_7605,N_6979);
or U10822 (N_10822,N_7952,N_8619);
nor U10823 (N_10823,N_6741,N_6530);
or U10824 (N_10824,N_6194,N_6607);
nor U10825 (N_10825,N_7857,N_8583);
and U10826 (N_10826,N_8550,N_6633);
or U10827 (N_10827,N_7511,N_6964);
nor U10828 (N_10828,N_7406,N_6247);
nor U10829 (N_10829,N_8245,N_7379);
or U10830 (N_10830,N_7911,N_6239);
nand U10831 (N_10831,N_8470,N_6072);
nand U10832 (N_10832,N_8317,N_6961);
nor U10833 (N_10833,N_8788,N_7410);
nand U10834 (N_10834,N_8063,N_6638);
and U10835 (N_10835,N_6406,N_8493);
nor U10836 (N_10836,N_8844,N_6163);
nand U10837 (N_10837,N_8949,N_6009);
or U10838 (N_10838,N_6856,N_6194);
and U10839 (N_10839,N_7870,N_7033);
or U10840 (N_10840,N_8769,N_8930);
nor U10841 (N_10841,N_8915,N_8881);
and U10842 (N_10842,N_7267,N_8104);
or U10843 (N_10843,N_8943,N_7600);
or U10844 (N_10844,N_6295,N_8443);
nand U10845 (N_10845,N_7322,N_6523);
nand U10846 (N_10846,N_7279,N_7661);
xnor U10847 (N_10847,N_6159,N_7357);
nand U10848 (N_10848,N_6655,N_7044);
and U10849 (N_10849,N_8816,N_7276);
nor U10850 (N_10850,N_8479,N_6973);
nor U10851 (N_10851,N_8355,N_8416);
nor U10852 (N_10852,N_7740,N_6832);
nand U10853 (N_10853,N_8224,N_7052);
nor U10854 (N_10854,N_7606,N_8386);
and U10855 (N_10855,N_8153,N_6772);
and U10856 (N_10856,N_7473,N_7140);
nand U10857 (N_10857,N_7346,N_7327);
and U10858 (N_10858,N_7189,N_7907);
nor U10859 (N_10859,N_7506,N_7257);
or U10860 (N_10860,N_7392,N_6269);
nand U10861 (N_10861,N_6230,N_6729);
and U10862 (N_10862,N_6881,N_6033);
nand U10863 (N_10863,N_6894,N_8112);
and U10864 (N_10864,N_7096,N_6351);
or U10865 (N_10865,N_8518,N_7300);
and U10866 (N_10866,N_7482,N_8961);
and U10867 (N_10867,N_6650,N_7039);
and U10868 (N_10868,N_8889,N_8946);
or U10869 (N_10869,N_6932,N_6447);
or U10870 (N_10870,N_8132,N_6939);
nand U10871 (N_10871,N_6325,N_6728);
and U10872 (N_10872,N_6196,N_6853);
and U10873 (N_10873,N_7792,N_7539);
and U10874 (N_10874,N_7761,N_8864);
or U10875 (N_10875,N_7742,N_7612);
nor U10876 (N_10876,N_7470,N_6463);
and U10877 (N_10877,N_8888,N_7890);
xor U10878 (N_10878,N_6009,N_6131);
nand U10879 (N_10879,N_8723,N_6543);
or U10880 (N_10880,N_8773,N_6405);
or U10881 (N_10881,N_8318,N_6221);
nand U10882 (N_10882,N_8722,N_6447);
and U10883 (N_10883,N_8271,N_6078);
nor U10884 (N_10884,N_6960,N_6446);
or U10885 (N_10885,N_6737,N_8365);
and U10886 (N_10886,N_8269,N_6510);
and U10887 (N_10887,N_6234,N_7449);
and U10888 (N_10888,N_7242,N_7785);
nand U10889 (N_10889,N_6853,N_7799);
and U10890 (N_10890,N_7625,N_7296);
or U10891 (N_10891,N_7384,N_6050);
nor U10892 (N_10892,N_6088,N_6361);
nand U10893 (N_10893,N_8376,N_8872);
or U10894 (N_10894,N_6208,N_7775);
and U10895 (N_10895,N_7105,N_6079);
nand U10896 (N_10896,N_7459,N_8323);
or U10897 (N_10897,N_8113,N_8204);
and U10898 (N_10898,N_8320,N_6688);
and U10899 (N_10899,N_8876,N_8919);
and U10900 (N_10900,N_8655,N_8857);
or U10901 (N_10901,N_6128,N_7753);
or U10902 (N_10902,N_8400,N_8262);
or U10903 (N_10903,N_6886,N_7353);
and U10904 (N_10904,N_7478,N_7484);
nor U10905 (N_10905,N_6172,N_8213);
nand U10906 (N_10906,N_7123,N_7658);
or U10907 (N_10907,N_6642,N_6955);
nor U10908 (N_10908,N_7887,N_8332);
or U10909 (N_10909,N_6706,N_6826);
nor U10910 (N_10910,N_8444,N_7436);
nor U10911 (N_10911,N_6384,N_6361);
or U10912 (N_10912,N_7786,N_6834);
or U10913 (N_10913,N_6027,N_6454);
nand U10914 (N_10914,N_8437,N_6101);
or U10915 (N_10915,N_8489,N_7543);
or U10916 (N_10916,N_8089,N_7491);
nand U10917 (N_10917,N_6712,N_6553);
and U10918 (N_10918,N_7491,N_8570);
or U10919 (N_10919,N_7321,N_8571);
or U10920 (N_10920,N_8564,N_8378);
nand U10921 (N_10921,N_6206,N_7625);
nor U10922 (N_10922,N_6724,N_7338);
nand U10923 (N_10923,N_6211,N_6214);
and U10924 (N_10924,N_6567,N_6559);
and U10925 (N_10925,N_6343,N_7819);
nand U10926 (N_10926,N_8009,N_8710);
nand U10927 (N_10927,N_8887,N_8169);
and U10928 (N_10928,N_6542,N_7243);
or U10929 (N_10929,N_6605,N_7557);
or U10930 (N_10930,N_7792,N_7735);
and U10931 (N_10931,N_8121,N_7618);
and U10932 (N_10932,N_7251,N_8772);
and U10933 (N_10933,N_8716,N_6517);
nor U10934 (N_10934,N_8009,N_7604);
and U10935 (N_10935,N_7148,N_7476);
or U10936 (N_10936,N_8514,N_6631);
nand U10937 (N_10937,N_7743,N_8832);
or U10938 (N_10938,N_8155,N_8521);
nor U10939 (N_10939,N_7806,N_7312);
nand U10940 (N_10940,N_7331,N_8718);
or U10941 (N_10941,N_6653,N_8036);
nor U10942 (N_10942,N_6825,N_6853);
nand U10943 (N_10943,N_8884,N_8987);
or U10944 (N_10944,N_6429,N_6042);
or U10945 (N_10945,N_7543,N_7423);
and U10946 (N_10946,N_6017,N_6469);
nor U10947 (N_10947,N_8254,N_6883);
nand U10948 (N_10948,N_7467,N_8200);
or U10949 (N_10949,N_8298,N_8244);
nand U10950 (N_10950,N_8305,N_6089);
nor U10951 (N_10951,N_8391,N_7182);
nand U10952 (N_10952,N_8431,N_8176);
and U10953 (N_10953,N_7993,N_6580);
and U10954 (N_10954,N_6523,N_6153);
and U10955 (N_10955,N_7898,N_8070);
or U10956 (N_10956,N_8260,N_8227);
or U10957 (N_10957,N_7176,N_7617);
and U10958 (N_10958,N_7838,N_8186);
or U10959 (N_10959,N_8386,N_7902);
or U10960 (N_10960,N_6903,N_8806);
nand U10961 (N_10961,N_6959,N_7432);
nor U10962 (N_10962,N_8465,N_8890);
or U10963 (N_10963,N_6528,N_7367);
or U10964 (N_10964,N_6962,N_6936);
nor U10965 (N_10965,N_7277,N_7807);
nor U10966 (N_10966,N_8018,N_7997);
nor U10967 (N_10967,N_7108,N_6664);
and U10968 (N_10968,N_6094,N_8041);
nand U10969 (N_10969,N_7331,N_8993);
or U10970 (N_10970,N_8986,N_7752);
or U10971 (N_10971,N_8619,N_8810);
nor U10972 (N_10972,N_6747,N_7559);
and U10973 (N_10973,N_6954,N_7029);
nor U10974 (N_10974,N_6597,N_8319);
nand U10975 (N_10975,N_8000,N_8472);
xor U10976 (N_10976,N_7193,N_8532);
and U10977 (N_10977,N_8536,N_8703);
and U10978 (N_10978,N_8967,N_8167);
and U10979 (N_10979,N_8826,N_6820);
nor U10980 (N_10980,N_6869,N_7458);
and U10981 (N_10981,N_8253,N_6852);
nand U10982 (N_10982,N_7726,N_8244);
and U10983 (N_10983,N_6852,N_8774);
or U10984 (N_10984,N_8180,N_8858);
nand U10985 (N_10985,N_8204,N_8925);
nor U10986 (N_10986,N_7916,N_8260);
nor U10987 (N_10987,N_7879,N_8260);
nor U10988 (N_10988,N_6539,N_6448);
or U10989 (N_10989,N_7341,N_7162);
and U10990 (N_10990,N_7034,N_7013);
or U10991 (N_10991,N_7144,N_6537);
and U10992 (N_10992,N_7776,N_8555);
nor U10993 (N_10993,N_8249,N_8995);
nor U10994 (N_10994,N_6441,N_7415);
or U10995 (N_10995,N_7538,N_8572);
nor U10996 (N_10996,N_8641,N_7051);
nor U10997 (N_10997,N_7300,N_7167);
and U10998 (N_10998,N_8576,N_6636);
nand U10999 (N_10999,N_7282,N_7152);
or U11000 (N_11000,N_6089,N_7211);
and U11001 (N_11001,N_6223,N_6087);
nor U11002 (N_11002,N_7044,N_7271);
or U11003 (N_11003,N_6336,N_6442);
or U11004 (N_11004,N_8547,N_8959);
or U11005 (N_11005,N_7269,N_8524);
or U11006 (N_11006,N_7087,N_6105);
nand U11007 (N_11007,N_8207,N_6518);
or U11008 (N_11008,N_8613,N_8919);
and U11009 (N_11009,N_6172,N_6209);
nor U11010 (N_11010,N_7120,N_7809);
nand U11011 (N_11011,N_6714,N_8877);
and U11012 (N_11012,N_8609,N_7823);
xor U11013 (N_11013,N_8368,N_7579);
nor U11014 (N_11014,N_7491,N_8163);
nand U11015 (N_11015,N_8703,N_7817);
or U11016 (N_11016,N_8825,N_7391);
nand U11017 (N_11017,N_7558,N_8331);
or U11018 (N_11018,N_7730,N_8241);
nor U11019 (N_11019,N_6655,N_7139);
and U11020 (N_11020,N_6439,N_6075);
and U11021 (N_11021,N_6255,N_7473);
or U11022 (N_11022,N_8249,N_7255);
or U11023 (N_11023,N_7814,N_8436);
nand U11024 (N_11024,N_7001,N_8862);
nand U11025 (N_11025,N_7041,N_8822);
nand U11026 (N_11026,N_7355,N_7072);
nor U11027 (N_11027,N_6835,N_8235);
xnor U11028 (N_11028,N_6720,N_7563);
or U11029 (N_11029,N_8277,N_6127);
nand U11030 (N_11030,N_6767,N_8360);
nor U11031 (N_11031,N_8124,N_7980);
nand U11032 (N_11032,N_7237,N_7468);
and U11033 (N_11033,N_6737,N_7311);
nor U11034 (N_11034,N_8011,N_8791);
and U11035 (N_11035,N_7526,N_8665);
and U11036 (N_11036,N_8720,N_7421);
nor U11037 (N_11037,N_6139,N_7016);
nor U11038 (N_11038,N_8752,N_8312);
nor U11039 (N_11039,N_8483,N_6399);
nor U11040 (N_11040,N_6865,N_8633);
nor U11041 (N_11041,N_6248,N_6719);
nor U11042 (N_11042,N_6335,N_6861);
and U11043 (N_11043,N_7524,N_7113);
nand U11044 (N_11044,N_6787,N_6166);
nor U11045 (N_11045,N_8370,N_6020);
xor U11046 (N_11046,N_8683,N_7472);
nor U11047 (N_11047,N_8218,N_7934);
xnor U11048 (N_11048,N_7105,N_8770);
and U11049 (N_11049,N_7481,N_7360);
nand U11050 (N_11050,N_7574,N_8944);
or U11051 (N_11051,N_8070,N_6439);
nor U11052 (N_11052,N_6907,N_6212);
or U11053 (N_11053,N_6328,N_7606);
nor U11054 (N_11054,N_8198,N_6282);
nor U11055 (N_11055,N_8916,N_6259);
nand U11056 (N_11056,N_8205,N_7033);
nand U11057 (N_11057,N_6756,N_7872);
and U11058 (N_11058,N_6989,N_7783);
nor U11059 (N_11059,N_7888,N_8173);
and U11060 (N_11060,N_6265,N_6945);
nor U11061 (N_11061,N_8734,N_7600);
nor U11062 (N_11062,N_6366,N_6545);
and U11063 (N_11063,N_7625,N_6559);
nor U11064 (N_11064,N_8940,N_7496);
nand U11065 (N_11065,N_7518,N_7288);
or U11066 (N_11066,N_7590,N_7747);
nor U11067 (N_11067,N_7822,N_8878);
or U11068 (N_11068,N_7295,N_7144);
nand U11069 (N_11069,N_8955,N_7706);
and U11070 (N_11070,N_8973,N_6943);
nor U11071 (N_11071,N_8089,N_6207);
or U11072 (N_11072,N_6747,N_7581);
nand U11073 (N_11073,N_8148,N_6461);
nor U11074 (N_11074,N_6250,N_7239);
nor U11075 (N_11075,N_6922,N_6881);
or U11076 (N_11076,N_7025,N_7950);
or U11077 (N_11077,N_8943,N_7248);
and U11078 (N_11078,N_6399,N_7521);
nor U11079 (N_11079,N_7426,N_7948);
nand U11080 (N_11080,N_6318,N_8530);
and U11081 (N_11081,N_7092,N_6275);
and U11082 (N_11082,N_8908,N_7681);
and U11083 (N_11083,N_7273,N_6907);
nand U11084 (N_11084,N_8476,N_6485);
and U11085 (N_11085,N_8137,N_6064);
nand U11086 (N_11086,N_8317,N_8055);
nor U11087 (N_11087,N_7688,N_6877);
nor U11088 (N_11088,N_7961,N_8594);
and U11089 (N_11089,N_7408,N_7759);
or U11090 (N_11090,N_6716,N_6417);
nor U11091 (N_11091,N_8705,N_6442);
and U11092 (N_11092,N_8298,N_6055);
nor U11093 (N_11093,N_8072,N_8669);
or U11094 (N_11094,N_6126,N_8699);
and U11095 (N_11095,N_6074,N_6237);
nand U11096 (N_11096,N_6880,N_8082);
and U11097 (N_11097,N_8023,N_8471);
or U11098 (N_11098,N_6275,N_8464);
nand U11099 (N_11099,N_8015,N_6246);
nand U11100 (N_11100,N_7733,N_6554);
or U11101 (N_11101,N_6776,N_8733);
nand U11102 (N_11102,N_7203,N_7406);
nand U11103 (N_11103,N_8591,N_8413);
nor U11104 (N_11104,N_8624,N_7289);
nand U11105 (N_11105,N_8874,N_7469);
nor U11106 (N_11106,N_8493,N_8003);
and U11107 (N_11107,N_7636,N_8808);
or U11108 (N_11108,N_6199,N_6341);
or U11109 (N_11109,N_6445,N_6570);
and U11110 (N_11110,N_6581,N_8868);
and U11111 (N_11111,N_7883,N_7330);
and U11112 (N_11112,N_7675,N_7686);
and U11113 (N_11113,N_7814,N_7987);
or U11114 (N_11114,N_7883,N_6837);
nor U11115 (N_11115,N_7627,N_7000);
nand U11116 (N_11116,N_8427,N_6894);
nor U11117 (N_11117,N_6429,N_7721);
nand U11118 (N_11118,N_6536,N_6059);
nor U11119 (N_11119,N_6041,N_6270);
nor U11120 (N_11120,N_8064,N_6896);
and U11121 (N_11121,N_6053,N_7762);
nor U11122 (N_11122,N_8381,N_6998);
or U11123 (N_11123,N_6624,N_8258);
and U11124 (N_11124,N_8541,N_7353);
nand U11125 (N_11125,N_7114,N_8191);
or U11126 (N_11126,N_6702,N_8907);
or U11127 (N_11127,N_6384,N_6095);
or U11128 (N_11128,N_8189,N_7958);
nor U11129 (N_11129,N_8644,N_7798);
nor U11130 (N_11130,N_8952,N_7657);
nand U11131 (N_11131,N_7579,N_6799);
nand U11132 (N_11132,N_7563,N_8636);
nand U11133 (N_11133,N_7566,N_7419);
nor U11134 (N_11134,N_7784,N_7753);
and U11135 (N_11135,N_8512,N_8399);
nor U11136 (N_11136,N_8865,N_7359);
nor U11137 (N_11137,N_8877,N_6810);
and U11138 (N_11138,N_8468,N_8570);
or U11139 (N_11139,N_8895,N_6352);
nor U11140 (N_11140,N_6738,N_7659);
nand U11141 (N_11141,N_6695,N_7348);
or U11142 (N_11142,N_6401,N_7759);
nor U11143 (N_11143,N_7069,N_8569);
nor U11144 (N_11144,N_7078,N_8391);
nor U11145 (N_11145,N_8837,N_6669);
and U11146 (N_11146,N_7388,N_8626);
and U11147 (N_11147,N_8473,N_6614);
and U11148 (N_11148,N_6010,N_7816);
xnor U11149 (N_11149,N_8757,N_6748);
nand U11150 (N_11150,N_7467,N_8531);
xnor U11151 (N_11151,N_8279,N_8506);
nor U11152 (N_11152,N_7451,N_8845);
or U11153 (N_11153,N_8293,N_6858);
nor U11154 (N_11154,N_8167,N_6006);
nand U11155 (N_11155,N_6069,N_6701);
or U11156 (N_11156,N_6056,N_7907);
nand U11157 (N_11157,N_6215,N_8582);
nor U11158 (N_11158,N_8554,N_7605);
nand U11159 (N_11159,N_8867,N_8772);
nor U11160 (N_11160,N_8129,N_8320);
nand U11161 (N_11161,N_8028,N_6633);
nand U11162 (N_11162,N_8869,N_8196);
and U11163 (N_11163,N_8643,N_8974);
nand U11164 (N_11164,N_7937,N_6898);
and U11165 (N_11165,N_6729,N_7672);
and U11166 (N_11166,N_6575,N_7103);
and U11167 (N_11167,N_8677,N_6189);
or U11168 (N_11168,N_7392,N_6348);
or U11169 (N_11169,N_7723,N_7534);
and U11170 (N_11170,N_7048,N_6908);
nand U11171 (N_11171,N_6907,N_7830);
and U11172 (N_11172,N_8587,N_6134);
nor U11173 (N_11173,N_6166,N_6675);
nor U11174 (N_11174,N_8818,N_6129);
nand U11175 (N_11175,N_6235,N_8030);
or U11176 (N_11176,N_8129,N_7292);
and U11177 (N_11177,N_8529,N_8180);
or U11178 (N_11178,N_6687,N_8871);
nor U11179 (N_11179,N_7065,N_8411);
or U11180 (N_11180,N_7563,N_7634);
nand U11181 (N_11181,N_8918,N_8880);
nor U11182 (N_11182,N_8809,N_6996);
nand U11183 (N_11183,N_6244,N_7098);
or U11184 (N_11184,N_6302,N_8058);
nor U11185 (N_11185,N_8133,N_8271);
nor U11186 (N_11186,N_6327,N_7432);
nor U11187 (N_11187,N_6304,N_8312);
and U11188 (N_11188,N_7142,N_7130);
or U11189 (N_11189,N_6890,N_6216);
or U11190 (N_11190,N_6245,N_6374);
or U11191 (N_11191,N_8464,N_8710);
nor U11192 (N_11192,N_8237,N_6346);
and U11193 (N_11193,N_8696,N_7412);
or U11194 (N_11194,N_8649,N_6373);
or U11195 (N_11195,N_7332,N_8423);
nor U11196 (N_11196,N_8231,N_7495);
and U11197 (N_11197,N_7837,N_6975);
nand U11198 (N_11198,N_7470,N_8110);
nor U11199 (N_11199,N_7282,N_7561);
nand U11200 (N_11200,N_8976,N_7638);
nand U11201 (N_11201,N_8804,N_8027);
or U11202 (N_11202,N_8434,N_7783);
and U11203 (N_11203,N_7828,N_6216);
nand U11204 (N_11204,N_8962,N_6722);
or U11205 (N_11205,N_7199,N_8585);
and U11206 (N_11206,N_8309,N_7976);
nand U11207 (N_11207,N_8549,N_8703);
nand U11208 (N_11208,N_6173,N_7809);
nor U11209 (N_11209,N_7384,N_8601);
nand U11210 (N_11210,N_6615,N_6868);
nor U11211 (N_11211,N_6595,N_8787);
nor U11212 (N_11212,N_7336,N_7640);
nor U11213 (N_11213,N_8153,N_6889);
and U11214 (N_11214,N_7193,N_8837);
or U11215 (N_11215,N_6640,N_7575);
or U11216 (N_11216,N_7663,N_8471);
and U11217 (N_11217,N_6236,N_7619);
nor U11218 (N_11218,N_7845,N_7505);
or U11219 (N_11219,N_6485,N_8455);
xnor U11220 (N_11220,N_8790,N_7859);
and U11221 (N_11221,N_6567,N_6678);
nor U11222 (N_11222,N_8497,N_6979);
and U11223 (N_11223,N_8276,N_6269);
nor U11224 (N_11224,N_8710,N_6701);
nor U11225 (N_11225,N_8953,N_7640);
and U11226 (N_11226,N_6205,N_7838);
nand U11227 (N_11227,N_8663,N_8341);
nand U11228 (N_11228,N_7284,N_7346);
nor U11229 (N_11229,N_8558,N_7283);
and U11230 (N_11230,N_7135,N_8168);
nor U11231 (N_11231,N_8349,N_7290);
nor U11232 (N_11232,N_7794,N_7945);
and U11233 (N_11233,N_7907,N_6133);
nor U11234 (N_11234,N_8927,N_7073);
xnor U11235 (N_11235,N_6553,N_8009);
and U11236 (N_11236,N_8353,N_8942);
nor U11237 (N_11237,N_7985,N_7101);
and U11238 (N_11238,N_7007,N_7853);
nor U11239 (N_11239,N_7399,N_8536);
and U11240 (N_11240,N_7548,N_7995);
nor U11241 (N_11241,N_7461,N_8295);
or U11242 (N_11242,N_6558,N_8013);
nor U11243 (N_11243,N_8153,N_7779);
or U11244 (N_11244,N_6791,N_6178);
nand U11245 (N_11245,N_8773,N_7987);
xor U11246 (N_11246,N_8658,N_7582);
nor U11247 (N_11247,N_7876,N_6566);
and U11248 (N_11248,N_7150,N_6007);
or U11249 (N_11249,N_8280,N_6973);
or U11250 (N_11250,N_7667,N_6323);
nand U11251 (N_11251,N_8941,N_7033);
and U11252 (N_11252,N_7650,N_6219);
or U11253 (N_11253,N_6195,N_6685);
nand U11254 (N_11254,N_8853,N_8032);
or U11255 (N_11255,N_7833,N_6071);
or U11256 (N_11256,N_7820,N_8073);
nor U11257 (N_11257,N_8291,N_6516);
and U11258 (N_11258,N_8367,N_8306);
nand U11259 (N_11259,N_8150,N_6886);
or U11260 (N_11260,N_6982,N_6938);
nand U11261 (N_11261,N_8211,N_7674);
nor U11262 (N_11262,N_6044,N_8648);
nor U11263 (N_11263,N_6302,N_7578);
nor U11264 (N_11264,N_7019,N_7822);
nand U11265 (N_11265,N_7979,N_6265);
nor U11266 (N_11266,N_6211,N_8440);
and U11267 (N_11267,N_6981,N_6201);
or U11268 (N_11268,N_6215,N_8632);
nor U11269 (N_11269,N_8049,N_8228);
nor U11270 (N_11270,N_8697,N_7914);
nand U11271 (N_11271,N_7000,N_7369);
nand U11272 (N_11272,N_7818,N_7441);
and U11273 (N_11273,N_8015,N_6534);
xor U11274 (N_11274,N_8106,N_8066);
or U11275 (N_11275,N_8073,N_8009);
nor U11276 (N_11276,N_8367,N_6763);
and U11277 (N_11277,N_8597,N_8119);
or U11278 (N_11278,N_8211,N_6661);
and U11279 (N_11279,N_7691,N_8990);
and U11280 (N_11280,N_8339,N_8917);
or U11281 (N_11281,N_8543,N_8155);
or U11282 (N_11282,N_7560,N_7561);
nand U11283 (N_11283,N_8778,N_8422);
nand U11284 (N_11284,N_8102,N_6441);
nand U11285 (N_11285,N_6698,N_6746);
nand U11286 (N_11286,N_7210,N_7770);
or U11287 (N_11287,N_8670,N_6887);
nor U11288 (N_11288,N_8025,N_8604);
and U11289 (N_11289,N_6528,N_7237);
or U11290 (N_11290,N_6087,N_6382);
nand U11291 (N_11291,N_6563,N_6312);
nor U11292 (N_11292,N_8062,N_6336);
and U11293 (N_11293,N_7925,N_7841);
and U11294 (N_11294,N_8590,N_7836);
nand U11295 (N_11295,N_7856,N_6756);
nor U11296 (N_11296,N_6628,N_6118);
nor U11297 (N_11297,N_6395,N_6436);
and U11298 (N_11298,N_7069,N_8851);
and U11299 (N_11299,N_8443,N_8848);
nand U11300 (N_11300,N_8155,N_7767);
nor U11301 (N_11301,N_7020,N_8211);
and U11302 (N_11302,N_8948,N_8755);
and U11303 (N_11303,N_8986,N_8679);
and U11304 (N_11304,N_8712,N_6821);
nand U11305 (N_11305,N_6061,N_6568);
nor U11306 (N_11306,N_7761,N_7887);
nor U11307 (N_11307,N_6288,N_7869);
and U11308 (N_11308,N_7558,N_7528);
or U11309 (N_11309,N_8290,N_6239);
and U11310 (N_11310,N_6522,N_8222);
nor U11311 (N_11311,N_8703,N_6103);
or U11312 (N_11312,N_8720,N_7584);
and U11313 (N_11313,N_6907,N_7113);
nor U11314 (N_11314,N_8557,N_6139);
nand U11315 (N_11315,N_8589,N_6575);
nand U11316 (N_11316,N_7353,N_6116);
nor U11317 (N_11317,N_7559,N_7256);
or U11318 (N_11318,N_8234,N_8531);
and U11319 (N_11319,N_7703,N_7811);
and U11320 (N_11320,N_8757,N_7699);
nand U11321 (N_11321,N_6245,N_6259);
and U11322 (N_11322,N_7103,N_6861);
nor U11323 (N_11323,N_8917,N_6441);
nand U11324 (N_11324,N_6107,N_7072);
nor U11325 (N_11325,N_8088,N_8562);
nand U11326 (N_11326,N_6646,N_7692);
nand U11327 (N_11327,N_8115,N_8499);
nor U11328 (N_11328,N_7917,N_7598);
nor U11329 (N_11329,N_6453,N_6800);
and U11330 (N_11330,N_6248,N_7459);
nor U11331 (N_11331,N_8551,N_7235);
and U11332 (N_11332,N_8299,N_8461);
or U11333 (N_11333,N_7624,N_6976);
and U11334 (N_11334,N_8595,N_7748);
and U11335 (N_11335,N_6879,N_6355);
nand U11336 (N_11336,N_7134,N_8474);
or U11337 (N_11337,N_7479,N_7485);
and U11338 (N_11338,N_8457,N_6366);
nor U11339 (N_11339,N_7060,N_6909);
or U11340 (N_11340,N_6015,N_6800);
nand U11341 (N_11341,N_7286,N_8739);
and U11342 (N_11342,N_8269,N_8981);
xor U11343 (N_11343,N_6374,N_8823);
nor U11344 (N_11344,N_7045,N_7922);
nor U11345 (N_11345,N_8712,N_6026);
nand U11346 (N_11346,N_8305,N_8476);
nor U11347 (N_11347,N_8885,N_8180);
nand U11348 (N_11348,N_8036,N_8503);
nand U11349 (N_11349,N_7180,N_7234);
and U11350 (N_11350,N_6678,N_8868);
nor U11351 (N_11351,N_8865,N_6335);
nor U11352 (N_11352,N_6996,N_6927);
or U11353 (N_11353,N_8317,N_6169);
nand U11354 (N_11354,N_6547,N_6035);
or U11355 (N_11355,N_8135,N_7921);
nor U11356 (N_11356,N_6361,N_8578);
and U11357 (N_11357,N_8465,N_6270);
or U11358 (N_11358,N_8988,N_6345);
nand U11359 (N_11359,N_6870,N_8278);
or U11360 (N_11360,N_6638,N_8095);
or U11361 (N_11361,N_8642,N_8197);
and U11362 (N_11362,N_8980,N_8038);
and U11363 (N_11363,N_6063,N_8269);
nand U11364 (N_11364,N_6444,N_6808);
xor U11365 (N_11365,N_6387,N_6328);
nand U11366 (N_11366,N_7915,N_8414);
or U11367 (N_11367,N_6723,N_7035);
or U11368 (N_11368,N_8275,N_8721);
nor U11369 (N_11369,N_6690,N_7398);
xor U11370 (N_11370,N_8125,N_6112);
nand U11371 (N_11371,N_7415,N_6507);
nor U11372 (N_11372,N_8823,N_8489);
nand U11373 (N_11373,N_8614,N_7460);
nand U11374 (N_11374,N_7604,N_7508);
nand U11375 (N_11375,N_8735,N_7696);
or U11376 (N_11376,N_6701,N_8786);
xor U11377 (N_11377,N_8247,N_8338);
nor U11378 (N_11378,N_7742,N_6434);
and U11379 (N_11379,N_8027,N_8241);
nand U11380 (N_11380,N_6445,N_6268);
or U11381 (N_11381,N_7210,N_8458);
and U11382 (N_11382,N_7491,N_8152);
and U11383 (N_11383,N_8547,N_6535);
or U11384 (N_11384,N_6026,N_8632);
nand U11385 (N_11385,N_8586,N_8508);
nor U11386 (N_11386,N_7742,N_8474);
xor U11387 (N_11387,N_7007,N_8704);
and U11388 (N_11388,N_8017,N_7535);
or U11389 (N_11389,N_8586,N_8612);
nor U11390 (N_11390,N_8240,N_6888);
and U11391 (N_11391,N_7269,N_8044);
and U11392 (N_11392,N_8805,N_7948);
and U11393 (N_11393,N_7153,N_6677);
or U11394 (N_11394,N_8800,N_7893);
and U11395 (N_11395,N_8674,N_7967);
nand U11396 (N_11396,N_6020,N_6056);
nand U11397 (N_11397,N_7222,N_7446);
and U11398 (N_11398,N_8681,N_7013);
nand U11399 (N_11399,N_7976,N_6968);
nand U11400 (N_11400,N_8242,N_6661);
or U11401 (N_11401,N_8579,N_8383);
and U11402 (N_11402,N_6513,N_6148);
or U11403 (N_11403,N_6654,N_7979);
and U11404 (N_11404,N_8210,N_7531);
nand U11405 (N_11405,N_6178,N_6348);
nor U11406 (N_11406,N_8369,N_8977);
nor U11407 (N_11407,N_8408,N_8923);
and U11408 (N_11408,N_6354,N_8461);
or U11409 (N_11409,N_6240,N_7077);
nand U11410 (N_11410,N_6064,N_8941);
and U11411 (N_11411,N_6961,N_7447);
nor U11412 (N_11412,N_7776,N_6953);
and U11413 (N_11413,N_7410,N_7699);
and U11414 (N_11414,N_7786,N_7428);
nor U11415 (N_11415,N_7477,N_6521);
and U11416 (N_11416,N_6059,N_6655);
or U11417 (N_11417,N_6209,N_7778);
nand U11418 (N_11418,N_6573,N_6770);
nor U11419 (N_11419,N_8890,N_8165);
and U11420 (N_11420,N_6726,N_6908);
nor U11421 (N_11421,N_8467,N_7696);
nor U11422 (N_11422,N_6619,N_7575);
nor U11423 (N_11423,N_6068,N_6031);
and U11424 (N_11424,N_6286,N_8179);
or U11425 (N_11425,N_8663,N_6414);
nor U11426 (N_11426,N_8256,N_6997);
nor U11427 (N_11427,N_7322,N_6231);
nand U11428 (N_11428,N_8753,N_6989);
or U11429 (N_11429,N_8591,N_7668);
and U11430 (N_11430,N_8941,N_7695);
nor U11431 (N_11431,N_8067,N_6729);
nand U11432 (N_11432,N_8028,N_6596);
nor U11433 (N_11433,N_7641,N_6748);
nor U11434 (N_11434,N_6579,N_8421);
or U11435 (N_11435,N_6816,N_7525);
nor U11436 (N_11436,N_7128,N_6731);
nand U11437 (N_11437,N_6700,N_7084);
and U11438 (N_11438,N_8036,N_6228);
and U11439 (N_11439,N_8952,N_8145);
nor U11440 (N_11440,N_7617,N_8209);
and U11441 (N_11441,N_6459,N_8889);
nor U11442 (N_11442,N_8714,N_8896);
and U11443 (N_11443,N_6037,N_6954);
and U11444 (N_11444,N_7977,N_8310);
xnor U11445 (N_11445,N_6272,N_8518);
and U11446 (N_11446,N_8655,N_6597);
nor U11447 (N_11447,N_7941,N_8130);
xor U11448 (N_11448,N_7115,N_7768);
and U11449 (N_11449,N_7248,N_8463);
nor U11450 (N_11450,N_8981,N_6362);
nor U11451 (N_11451,N_7406,N_6272);
nand U11452 (N_11452,N_6787,N_6583);
nand U11453 (N_11453,N_7916,N_6467);
nand U11454 (N_11454,N_6283,N_7578);
and U11455 (N_11455,N_6069,N_7433);
or U11456 (N_11456,N_8676,N_8011);
or U11457 (N_11457,N_7033,N_7039);
and U11458 (N_11458,N_8561,N_6150);
or U11459 (N_11459,N_6637,N_8432);
and U11460 (N_11460,N_8172,N_8933);
and U11461 (N_11461,N_6397,N_6764);
nand U11462 (N_11462,N_7043,N_7776);
and U11463 (N_11463,N_8137,N_6455);
nor U11464 (N_11464,N_7154,N_6130);
or U11465 (N_11465,N_6947,N_6773);
nand U11466 (N_11466,N_8746,N_8362);
nor U11467 (N_11467,N_6421,N_8419);
nor U11468 (N_11468,N_8590,N_8094);
nand U11469 (N_11469,N_7352,N_7915);
nor U11470 (N_11470,N_8235,N_6709);
or U11471 (N_11471,N_8685,N_6140);
or U11472 (N_11472,N_6884,N_7634);
nand U11473 (N_11473,N_6621,N_8843);
and U11474 (N_11474,N_7768,N_8671);
or U11475 (N_11475,N_7435,N_8918);
or U11476 (N_11476,N_8453,N_6897);
or U11477 (N_11477,N_8654,N_7081);
nand U11478 (N_11478,N_7837,N_7999);
nand U11479 (N_11479,N_8505,N_6735);
nor U11480 (N_11480,N_8032,N_7921);
nor U11481 (N_11481,N_7657,N_7579);
or U11482 (N_11482,N_6500,N_8893);
and U11483 (N_11483,N_7296,N_6058);
and U11484 (N_11484,N_6096,N_6615);
or U11485 (N_11485,N_7615,N_8040);
nand U11486 (N_11486,N_6899,N_7099);
nand U11487 (N_11487,N_8022,N_6057);
nand U11488 (N_11488,N_6512,N_6102);
nor U11489 (N_11489,N_7863,N_6835);
nand U11490 (N_11490,N_8786,N_7077);
nand U11491 (N_11491,N_6347,N_6323);
nand U11492 (N_11492,N_8115,N_6224);
nand U11493 (N_11493,N_7250,N_6334);
nor U11494 (N_11494,N_6668,N_6142);
nor U11495 (N_11495,N_6286,N_7103);
or U11496 (N_11496,N_7190,N_7702);
and U11497 (N_11497,N_8536,N_7568);
or U11498 (N_11498,N_8728,N_7347);
xnor U11499 (N_11499,N_8386,N_6104);
or U11500 (N_11500,N_8978,N_6055);
nand U11501 (N_11501,N_7975,N_6605);
and U11502 (N_11502,N_7404,N_6895);
nand U11503 (N_11503,N_6469,N_8551);
and U11504 (N_11504,N_8644,N_7655);
or U11505 (N_11505,N_6975,N_6563);
nor U11506 (N_11506,N_6180,N_7239);
or U11507 (N_11507,N_6641,N_7272);
nand U11508 (N_11508,N_7284,N_7910);
and U11509 (N_11509,N_8970,N_7103);
nand U11510 (N_11510,N_6502,N_8995);
or U11511 (N_11511,N_8942,N_6120);
nor U11512 (N_11512,N_7722,N_7921);
nand U11513 (N_11513,N_6624,N_8997);
and U11514 (N_11514,N_6489,N_7858);
or U11515 (N_11515,N_6844,N_6608);
nor U11516 (N_11516,N_8846,N_6752);
nand U11517 (N_11517,N_8630,N_7417);
or U11518 (N_11518,N_6842,N_6536);
and U11519 (N_11519,N_6756,N_8506);
nand U11520 (N_11520,N_6929,N_8842);
or U11521 (N_11521,N_6336,N_6786);
nand U11522 (N_11522,N_8972,N_7813);
or U11523 (N_11523,N_7481,N_7497);
and U11524 (N_11524,N_8782,N_6100);
or U11525 (N_11525,N_7608,N_6838);
or U11526 (N_11526,N_6294,N_6206);
and U11527 (N_11527,N_6507,N_8037);
and U11528 (N_11528,N_8021,N_6466);
nand U11529 (N_11529,N_6421,N_8038);
nor U11530 (N_11530,N_6137,N_8586);
or U11531 (N_11531,N_8096,N_6413);
nor U11532 (N_11532,N_7252,N_8684);
and U11533 (N_11533,N_8294,N_8182);
or U11534 (N_11534,N_7250,N_8237);
or U11535 (N_11535,N_6497,N_8609);
nand U11536 (N_11536,N_8307,N_7583);
or U11537 (N_11537,N_6904,N_6548);
xnor U11538 (N_11538,N_7567,N_8215);
nand U11539 (N_11539,N_7789,N_7777);
xnor U11540 (N_11540,N_7122,N_6743);
nor U11541 (N_11541,N_6129,N_8287);
and U11542 (N_11542,N_7504,N_8757);
nor U11543 (N_11543,N_6981,N_6319);
nor U11544 (N_11544,N_7831,N_6238);
and U11545 (N_11545,N_8954,N_6438);
nor U11546 (N_11546,N_8564,N_7348);
nor U11547 (N_11547,N_7372,N_8513);
and U11548 (N_11548,N_8173,N_7830);
nor U11549 (N_11549,N_7799,N_6546);
nor U11550 (N_11550,N_6892,N_7136);
nand U11551 (N_11551,N_8233,N_6700);
nand U11552 (N_11552,N_8680,N_7287);
or U11553 (N_11553,N_7657,N_7890);
or U11554 (N_11554,N_8759,N_7113);
nor U11555 (N_11555,N_6126,N_6465);
and U11556 (N_11556,N_6669,N_6644);
and U11557 (N_11557,N_6301,N_8277);
or U11558 (N_11558,N_7192,N_7923);
nand U11559 (N_11559,N_7873,N_7550);
or U11560 (N_11560,N_7477,N_6929);
and U11561 (N_11561,N_6271,N_8804);
and U11562 (N_11562,N_6580,N_8834);
or U11563 (N_11563,N_6793,N_6629);
and U11564 (N_11564,N_6584,N_8232);
or U11565 (N_11565,N_7371,N_6813);
nand U11566 (N_11566,N_6926,N_6499);
nor U11567 (N_11567,N_8878,N_8734);
and U11568 (N_11568,N_7726,N_6290);
nand U11569 (N_11569,N_6284,N_6448);
nor U11570 (N_11570,N_8228,N_6465);
nand U11571 (N_11571,N_6029,N_7341);
nand U11572 (N_11572,N_8443,N_6165);
or U11573 (N_11573,N_8391,N_7207);
xor U11574 (N_11574,N_7885,N_7225);
or U11575 (N_11575,N_8150,N_6953);
nor U11576 (N_11576,N_6300,N_6968);
and U11577 (N_11577,N_6823,N_8120);
nand U11578 (N_11578,N_7444,N_8257);
and U11579 (N_11579,N_6890,N_7858);
or U11580 (N_11580,N_6950,N_8541);
nor U11581 (N_11581,N_8447,N_6446);
nand U11582 (N_11582,N_8790,N_6175);
nand U11583 (N_11583,N_7657,N_8159);
or U11584 (N_11584,N_7612,N_8559);
or U11585 (N_11585,N_6881,N_6397);
or U11586 (N_11586,N_8460,N_6852);
nand U11587 (N_11587,N_6734,N_7672);
or U11588 (N_11588,N_8364,N_7611);
or U11589 (N_11589,N_7996,N_8829);
and U11590 (N_11590,N_6094,N_8249);
or U11591 (N_11591,N_8937,N_6778);
or U11592 (N_11592,N_7259,N_8466);
and U11593 (N_11593,N_6929,N_7578);
nand U11594 (N_11594,N_7648,N_6740);
or U11595 (N_11595,N_7296,N_6016);
and U11596 (N_11596,N_6795,N_7646);
and U11597 (N_11597,N_6515,N_6299);
nor U11598 (N_11598,N_6653,N_6922);
or U11599 (N_11599,N_7722,N_8722);
and U11600 (N_11600,N_7715,N_6269);
nor U11601 (N_11601,N_7165,N_7525);
nand U11602 (N_11602,N_7004,N_6289);
or U11603 (N_11603,N_7762,N_7598);
and U11604 (N_11604,N_6449,N_8121);
nand U11605 (N_11605,N_7547,N_7420);
or U11606 (N_11606,N_8235,N_7435);
and U11607 (N_11607,N_8171,N_6655);
nor U11608 (N_11608,N_7097,N_7126);
and U11609 (N_11609,N_6577,N_7662);
and U11610 (N_11610,N_8514,N_7411);
nand U11611 (N_11611,N_8561,N_8212);
and U11612 (N_11612,N_8346,N_8455);
and U11613 (N_11613,N_7818,N_6396);
and U11614 (N_11614,N_6521,N_6327);
or U11615 (N_11615,N_7892,N_6852);
or U11616 (N_11616,N_8671,N_7306);
nand U11617 (N_11617,N_6107,N_8115);
nand U11618 (N_11618,N_8525,N_8251);
or U11619 (N_11619,N_8122,N_8134);
or U11620 (N_11620,N_6380,N_8811);
nor U11621 (N_11621,N_6994,N_8021);
or U11622 (N_11622,N_8535,N_6410);
or U11623 (N_11623,N_8175,N_8941);
and U11624 (N_11624,N_7099,N_6752);
or U11625 (N_11625,N_7609,N_8257);
nor U11626 (N_11626,N_7554,N_7482);
or U11627 (N_11627,N_6881,N_6487);
nand U11628 (N_11628,N_7150,N_8715);
nand U11629 (N_11629,N_8429,N_6434);
and U11630 (N_11630,N_6856,N_8525);
nor U11631 (N_11631,N_6493,N_7275);
or U11632 (N_11632,N_7926,N_8146);
nor U11633 (N_11633,N_7275,N_6141);
and U11634 (N_11634,N_6902,N_7837);
or U11635 (N_11635,N_6509,N_6282);
nor U11636 (N_11636,N_6587,N_8503);
or U11637 (N_11637,N_7584,N_6460);
nand U11638 (N_11638,N_7426,N_7348);
or U11639 (N_11639,N_8006,N_6861);
nor U11640 (N_11640,N_8994,N_7264);
nand U11641 (N_11641,N_6559,N_7261);
nand U11642 (N_11642,N_6358,N_8583);
or U11643 (N_11643,N_8920,N_6653);
nor U11644 (N_11644,N_6509,N_7087);
and U11645 (N_11645,N_7268,N_7235);
and U11646 (N_11646,N_7403,N_8781);
or U11647 (N_11647,N_8953,N_6277);
nand U11648 (N_11648,N_7969,N_6890);
nand U11649 (N_11649,N_7571,N_8960);
and U11650 (N_11650,N_7450,N_7330);
nor U11651 (N_11651,N_8763,N_8975);
nand U11652 (N_11652,N_6018,N_8545);
or U11653 (N_11653,N_7436,N_7033);
or U11654 (N_11654,N_8899,N_8168);
nor U11655 (N_11655,N_6100,N_6014);
or U11656 (N_11656,N_8118,N_7653);
nand U11657 (N_11657,N_8307,N_8302);
nor U11658 (N_11658,N_6880,N_7782);
nand U11659 (N_11659,N_7748,N_8478);
and U11660 (N_11660,N_6795,N_6963);
nand U11661 (N_11661,N_6055,N_7794);
nor U11662 (N_11662,N_6577,N_8660);
nand U11663 (N_11663,N_8576,N_7797);
and U11664 (N_11664,N_6030,N_6304);
nor U11665 (N_11665,N_7674,N_8549);
and U11666 (N_11666,N_7018,N_6467);
or U11667 (N_11667,N_7531,N_8285);
and U11668 (N_11668,N_6375,N_6495);
and U11669 (N_11669,N_7520,N_7115);
nand U11670 (N_11670,N_7718,N_8145);
nand U11671 (N_11671,N_8915,N_8947);
nand U11672 (N_11672,N_7811,N_7077);
nand U11673 (N_11673,N_7040,N_8546);
or U11674 (N_11674,N_7026,N_6922);
nand U11675 (N_11675,N_7563,N_7242);
nor U11676 (N_11676,N_6755,N_6987);
nor U11677 (N_11677,N_7863,N_6834);
or U11678 (N_11678,N_8587,N_6103);
nor U11679 (N_11679,N_7357,N_8758);
or U11680 (N_11680,N_8392,N_7944);
nor U11681 (N_11681,N_6958,N_6889);
and U11682 (N_11682,N_6207,N_7126);
nor U11683 (N_11683,N_6976,N_7839);
and U11684 (N_11684,N_7329,N_8703);
nor U11685 (N_11685,N_8233,N_6289);
nor U11686 (N_11686,N_7466,N_8089);
or U11687 (N_11687,N_8952,N_7350);
nor U11688 (N_11688,N_7446,N_7379);
nand U11689 (N_11689,N_7114,N_6064);
nand U11690 (N_11690,N_7773,N_6583);
xnor U11691 (N_11691,N_6392,N_7090);
nand U11692 (N_11692,N_7123,N_8112);
and U11693 (N_11693,N_6181,N_7620);
nor U11694 (N_11694,N_6750,N_7002);
nand U11695 (N_11695,N_7984,N_6757);
or U11696 (N_11696,N_8423,N_8343);
nor U11697 (N_11697,N_7061,N_7487);
and U11698 (N_11698,N_7969,N_8016);
nand U11699 (N_11699,N_7298,N_7874);
nand U11700 (N_11700,N_7998,N_8602);
and U11701 (N_11701,N_7841,N_8221);
and U11702 (N_11702,N_8410,N_7844);
nor U11703 (N_11703,N_6758,N_7503);
or U11704 (N_11704,N_8863,N_8236);
nor U11705 (N_11705,N_7190,N_8087);
or U11706 (N_11706,N_7658,N_8952);
nor U11707 (N_11707,N_6455,N_7559);
and U11708 (N_11708,N_7117,N_8274);
and U11709 (N_11709,N_7298,N_7943);
nor U11710 (N_11710,N_6596,N_6448);
or U11711 (N_11711,N_7686,N_6033);
nor U11712 (N_11712,N_6565,N_8331);
and U11713 (N_11713,N_7296,N_6533);
nor U11714 (N_11714,N_7130,N_8317);
nor U11715 (N_11715,N_8089,N_8342);
nor U11716 (N_11716,N_7391,N_7086);
nor U11717 (N_11717,N_8924,N_8866);
nor U11718 (N_11718,N_7727,N_7501);
nor U11719 (N_11719,N_6971,N_6351);
nor U11720 (N_11720,N_7673,N_7177);
or U11721 (N_11721,N_6441,N_7774);
and U11722 (N_11722,N_8110,N_7150);
nand U11723 (N_11723,N_8010,N_7971);
nand U11724 (N_11724,N_6625,N_7409);
nor U11725 (N_11725,N_7721,N_7198);
nand U11726 (N_11726,N_6811,N_7105);
and U11727 (N_11727,N_8577,N_6813);
or U11728 (N_11728,N_8413,N_6395);
or U11729 (N_11729,N_6639,N_8298);
and U11730 (N_11730,N_7274,N_7567);
nor U11731 (N_11731,N_7896,N_7323);
nand U11732 (N_11732,N_6028,N_7055);
nor U11733 (N_11733,N_6333,N_6798);
nor U11734 (N_11734,N_6716,N_7323);
nand U11735 (N_11735,N_6200,N_8027);
nand U11736 (N_11736,N_8904,N_6816);
or U11737 (N_11737,N_7610,N_8307);
and U11738 (N_11738,N_7262,N_8038);
nand U11739 (N_11739,N_8860,N_6711);
nand U11740 (N_11740,N_7461,N_8083);
nand U11741 (N_11741,N_7528,N_6204);
and U11742 (N_11742,N_7775,N_7361);
and U11743 (N_11743,N_6278,N_6740);
and U11744 (N_11744,N_8946,N_8382);
or U11745 (N_11745,N_6677,N_7780);
and U11746 (N_11746,N_6052,N_7594);
and U11747 (N_11747,N_6671,N_6864);
nor U11748 (N_11748,N_6694,N_6704);
nor U11749 (N_11749,N_6449,N_8964);
nor U11750 (N_11750,N_6359,N_8418);
nor U11751 (N_11751,N_8290,N_8669);
and U11752 (N_11752,N_8749,N_6413);
nand U11753 (N_11753,N_7993,N_7684);
and U11754 (N_11754,N_6425,N_7697);
or U11755 (N_11755,N_7691,N_6523);
and U11756 (N_11756,N_8344,N_7715);
or U11757 (N_11757,N_7013,N_7065);
and U11758 (N_11758,N_8060,N_6045);
nor U11759 (N_11759,N_6850,N_7751);
xnor U11760 (N_11760,N_6485,N_7040);
nand U11761 (N_11761,N_7852,N_8127);
nand U11762 (N_11762,N_7847,N_6080);
and U11763 (N_11763,N_7737,N_8094);
nand U11764 (N_11764,N_8268,N_7146);
or U11765 (N_11765,N_6667,N_8748);
nand U11766 (N_11766,N_6927,N_8096);
xor U11767 (N_11767,N_7273,N_7277);
nand U11768 (N_11768,N_8903,N_8136);
and U11769 (N_11769,N_8358,N_8085);
nand U11770 (N_11770,N_8513,N_6702);
nand U11771 (N_11771,N_6645,N_6359);
xor U11772 (N_11772,N_8358,N_8859);
and U11773 (N_11773,N_8353,N_6218);
nor U11774 (N_11774,N_8020,N_7799);
nor U11775 (N_11775,N_6683,N_7368);
nor U11776 (N_11776,N_6353,N_6570);
and U11777 (N_11777,N_7227,N_6953);
and U11778 (N_11778,N_8748,N_8087);
nand U11779 (N_11779,N_6678,N_7849);
or U11780 (N_11780,N_6867,N_7974);
nor U11781 (N_11781,N_7086,N_8345);
and U11782 (N_11782,N_7750,N_7334);
or U11783 (N_11783,N_7354,N_8006);
or U11784 (N_11784,N_7188,N_6280);
nand U11785 (N_11785,N_7695,N_8045);
nand U11786 (N_11786,N_6352,N_6877);
xnor U11787 (N_11787,N_8348,N_6874);
and U11788 (N_11788,N_8114,N_7723);
nor U11789 (N_11789,N_8871,N_8295);
nand U11790 (N_11790,N_6640,N_7722);
and U11791 (N_11791,N_7384,N_6532);
and U11792 (N_11792,N_8157,N_6172);
and U11793 (N_11793,N_8696,N_7339);
nand U11794 (N_11794,N_6896,N_8724);
or U11795 (N_11795,N_6758,N_8969);
nand U11796 (N_11796,N_8268,N_8612);
or U11797 (N_11797,N_7239,N_7236);
nor U11798 (N_11798,N_7679,N_7153);
nor U11799 (N_11799,N_7715,N_6545);
or U11800 (N_11800,N_6217,N_8855);
and U11801 (N_11801,N_6612,N_7948);
or U11802 (N_11802,N_6517,N_8450);
and U11803 (N_11803,N_7991,N_7702);
nor U11804 (N_11804,N_6378,N_8657);
or U11805 (N_11805,N_6202,N_6455);
nand U11806 (N_11806,N_7881,N_7587);
nand U11807 (N_11807,N_6431,N_7067);
nor U11808 (N_11808,N_8255,N_7333);
nand U11809 (N_11809,N_7271,N_7883);
and U11810 (N_11810,N_8402,N_6723);
or U11811 (N_11811,N_6332,N_8707);
nand U11812 (N_11812,N_7641,N_8735);
nand U11813 (N_11813,N_6830,N_8743);
and U11814 (N_11814,N_8107,N_7397);
nand U11815 (N_11815,N_7365,N_7684);
nor U11816 (N_11816,N_7607,N_6675);
or U11817 (N_11817,N_8965,N_6684);
nand U11818 (N_11818,N_8066,N_7307);
nand U11819 (N_11819,N_6961,N_7484);
nor U11820 (N_11820,N_6898,N_7949);
or U11821 (N_11821,N_8978,N_7670);
or U11822 (N_11822,N_7078,N_7047);
or U11823 (N_11823,N_6789,N_7490);
and U11824 (N_11824,N_7376,N_7771);
or U11825 (N_11825,N_8428,N_6399);
nand U11826 (N_11826,N_6965,N_6340);
or U11827 (N_11827,N_7539,N_7967);
or U11828 (N_11828,N_8760,N_6272);
nand U11829 (N_11829,N_8603,N_8704);
nand U11830 (N_11830,N_6427,N_6070);
or U11831 (N_11831,N_8108,N_8401);
and U11832 (N_11832,N_8835,N_7195);
or U11833 (N_11833,N_8501,N_7525);
nor U11834 (N_11834,N_7986,N_7560);
nand U11835 (N_11835,N_7016,N_7231);
and U11836 (N_11836,N_6781,N_7303);
and U11837 (N_11837,N_8665,N_8297);
nor U11838 (N_11838,N_6357,N_8303);
nand U11839 (N_11839,N_6775,N_6944);
nand U11840 (N_11840,N_6186,N_8084);
nand U11841 (N_11841,N_7643,N_7600);
nor U11842 (N_11842,N_7657,N_8914);
or U11843 (N_11843,N_6288,N_7966);
or U11844 (N_11844,N_6145,N_7551);
nor U11845 (N_11845,N_7491,N_6369);
and U11846 (N_11846,N_7382,N_6816);
nor U11847 (N_11847,N_7507,N_6936);
or U11848 (N_11848,N_7787,N_8665);
nor U11849 (N_11849,N_7775,N_7052);
nand U11850 (N_11850,N_8779,N_8641);
or U11851 (N_11851,N_7428,N_7206);
nor U11852 (N_11852,N_7790,N_8498);
nand U11853 (N_11853,N_8580,N_6002);
nor U11854 (N_11854,N_8735,N_6180);
nor U11855 (N_11855,N_8122,N_8177);
nand U11856 (N_11856,N_7481,N_6666);
and U11857 (N_11857,N_6801,N_7687);
nor U11858 (N_11858,N_6339,N_7270);
and U11859 (N_11859,N_6193,N_8153);
and U11860 (N_11860,N_6664,N_8295);
or U11861 (N_11861,N_8033,N_8230);
and U11862 (N_11862,N_7651,N_6650);
nor U11863 (N_11863,N_7466,N_6896);
and U11864 (N_11864,N_7589,N_8204);
nand U11865 (N_11865,N_7732,N_8422);
nand U11866 (N_11866,N_7396,N_7003);
nor U11867 (N_11867,N_7871,N_6030);
nand U11868 (N_11868,N_7557,N_8985);
nand U11869 (N_11869,N_7655,N_7133);
nor U11870 (N_11870,N_6470,N_8121);
nand U11871 (N_11871,N_6143,N_8717);
nand U11872 (N_11872,N_7416,N_6079);
nor U11873 (N_11873,N_8218,N_8729);
xnor U11874 (N_11874,N_6786,N_7351);
xnor U11875 (N_11875,N_7124,N_8543);
and U11876 (N_11876,N_8462,N_7373);
nand U11877 (N_11877,N_6467,N_7000);
or U11878 (N_11878,N_8484,N_7033);
and U11879 (N_11879,N_6815,N_8429);
nand U11880 (N_11880,N_7298,N_6606);
xnor U11881 (N_11881,N_8680,N_7375);
nor U11882 (N_11882,N_7242,N_6884);
or U11883 (N_11883,N_6081,N_6055);
nand U11884 (N_11884,N_6745,N_7164);
nor U11885 (N_11885,N_6662,N_6074);
and U11886 (N_11886,N_7299,N_6303);
and U11887 (N_11887,N_8617,N_6750);
and U11888 (N_11888,N_8810,N_8388);
or U11889 (N_11889,N_8857,N_6144);
nor U11890 (N_11890,N_7897,N_6353);
nor U11891 (N_11891,N_7254,N_8997);
or U11892 (N_11892,N_8341,N_8137);
or U11893 (N_11893,N_6077,N_8577);
and U11894 (N_11894,N_6403,N_7289);
and U11895 (N_11895,N_6490,N_6060);
and U11896 (N_11896,N_7412,N_8875);
and U11897 (N_11897,N_7671,N_6872);
nand U11898 (N_11898,N_8426,N_7324);
or U11899 (N_11899,N_6215,N_7336);
or U11900 (N_11900,N_8455,N_8649);
nand U11901 (N_11901,N_8585,N_8912);
nand U11902 (N_11902,N_6789,N_7011);
and U11903 (N_11903,N_7139,N_6949);
nor U11904 (N_11904,N_6971,N_8688);
or U11905 (N_11905,N_8263,N_6104);
nor U11906 (N_11906,N_7050,N_6069);
nor U11907 (N_11907,N_7225,N_8431);
nor U11908 (N_11908,N_6749,N_6794);
nand U11909 (N_11909,N_8565,N_6993);
nor U11910 (N_11910,N_7847,N_7369);
or U11911 (N_11911,N_6278,N_8593);
and U11912 (N_11912,N_8234,N_7840);
nor U11913 (N_11913,N_7063,N_6354);
or U11914 (N_11914,N_6747,N_6509);
and U11915 (N_11915,N_8347,N_7697);
and U11916 (N_11916,N_7072,N_6351);
nor U11917 (N_11917,N_6632,N_7745);
nor U11918 (N_11918,N_7919,N_6684);
and U11919 (N_11919,N_6513,N_7957);
and U11920 (N_11920,N_6527,N_8860);
or U11921 (N_11921,N_7371,N_7377);
and U11922 (N_11922,N_6847,N_6072);
and U11923 (N_11923,N_6420,N_8929);
and U11924 (N_11924,N_6428,N_6207);
nand U11925 (N_11925,N_8601,N_8239);
nor U11926 (N_11926,N_7825,N_6336);
nor U11927 (N_11927,N_7798,N_6651);
and U11928 (N_11928,N_6789,N_7728);
nand U11929 (N_11929,N_8987,N_6841);
nand U11930 (N_11930,N_6174,N_7025);
nand U11931 (N_11931,N_8391,N_7264);
and U11932 (N_11932,N_7565,N_6951);
and U11933 (N_11933,N_8806,N_7992);
and U11934 (N_11934,N_6343,N_7771);
or U11935 (N_11935,N_7896,N_8210);
nand U11936 (N_11936,N_8774,N_7168);
nand U11937 (N_11937,N_6515,N_7546);
and U11938 (N_11938,N_8947,N_6451);
nor U11939 (N_11939,N_8393,N_6797);
nor U11940 (N_11940,N_8252,N_6047);
nand U11941 (N_11941,N_7818,N_8511);
nor U11942 (N_11942,N_6431,N_6705);
and U11943 (N_11943,N_8544,N_6774);
nor U11944 (N_11944,N_7483,N_6889);
and U11945 (N_11945,N_7767,N_8768);
or U11946 (N_11946,N_7119,N_7781);
or U11947 (N_11947,N_7230,N_7326);
or U11948 (N_11948,N_7011,N_7467);
nand U11949 (N_11949,N_7363,N_7654);
nor U11950 (N_11950,N_6291,N_7389);
or U11951 (N_11951,N_6898,N_7169);
nor U11952 (N_11952,N_6724,N_6325);
or U11953 (N_11953,N_7917,N_6656);
and U11954 (N_11954,N_7345,N_7078);
or U11955 (N_11955,N_7611,N_6754);
or U11956 (N_11956,N_7108,N_8587);
nor U11957 (N_11957,N_7157,N_8378);
and U11958 (N_11958,N_7352,N_8153);
or U11959 (N_11959,N_6616,N_8423);
or U11960 (N_11960,N_8209,N_8784);
and U11961 (N_11961,N_8582,N_7509);
nand U11962 (N_11962,N_6907,N_8560);
and U11963 (N_11963,N_7547,N_7930);
nor U11964 (N_11964,N_7085,N_7475);
and U11965 (N_11965,N_8481,N_8597);
nand U11966 (N_11966,N_6288,N_6003);
or U11967 (N_11967,N_6404,N_6762);
or U11968 (N_11968,N_8176,N_7182);
nor U11969 (N_11969,N_6127,N_7708);
xnor U11970 (N_11970,N_7136,N_6648);
nand U11971 (N_11971,N_8256,N_6123);
nand U11972 (N_11972,N_7469,N_8201);
nor U11973 (N_11973,N_8826,N_6819);
nor U11974 (N_11974,N_7215,N_6083);
nand U11975 (N_11975,N_6977,N_6800);
nor U11976 (N_11976,N_6203,N_6496);
nand U11977 (N_11977,N_8015,N_8386);
nor U11978 (N_11978,N_7387,N_7076);
or U11979 (N_11979,N_7650,N_6360);
nor U11980 (N_11980,N_8113,N_7713);
nand U11981 (N_11981,N_8984,N_7107);
or U11982 (N_11982,N_6942,N_8564);
nor U11983 (N_11983,N_8735,N_6205);
nor U11984 (N_11984,N_6532,N_7779);
nor U11985 (N_11985,N_7491,N_6187);
nor U11986 (N_11986,N_6594,N_6169);
nand U11987 (N_11987,N_7432,N_6272);
nand U11988 (N_11988,N_6074,N_6605);
nor U11989 (N_11989,N_8089,N_7328);
nand U11990 (N_11990,N_8891,N_6388);
and U11991 (N_11991,N_6822,N_6169);
or U11992 (N_11992,N_7185,N_8425);
xnor U11993 (N_11993,N_6125,N_8443);
nand U11994 (N_11994,N_7136,N_6382);
and U11995 (N_11995,N_8206,N_7029);
nor U11996 (N_11996,N_6110,N_7357);
or U11997 (N_11997,N_6687,N_6609);
nor U11998 (N_11998,N_6294,N_7314);
and U11999 (N_11999,N_8294,N_8106);
or U12000 (N_12000,N_10441,N_9509);
nand U12001 (N_12001,N_10945,N_10506);
nor U12002 (N_12002,N_10776,N_9840);
and U12003 (N_12003,N_10458,N_9845);
nor U12004 (N_12004,N_11896,N_11073);
or U12005 (N_12005,N_11215,N_10371);
and U12006 (N_12006,N_11994,N_9388);
and U12007 (N_12007,N_11977,N_9265);
nand U12008 (N_12008,N_9135,N_11616);
or U12009 (N_12009,N_11317,N_10723);
nor U12010 (N_12010,N_9182,N_11097);
nor U12011 (N_12011,N_9128,N_10327);
or U12012 (N_12012,N_9444,N_10392);
and U12013 (N_12013,N_11422,N_9919);
and U12014 (N_12014,N_11483,N_10321);
nand U12015 (N_12015,N_9007,N_9886);
and U12016 (N_12016,N_10678,N_11840);
and U12017 (N_12017,N_10164,N_9391);
nor U12018 (N_12018,N_11057,N_9584);
and U12019 (N_12019,N_10648,N_10501);
nand U12020 (N_12020,N_11711,N_9168);
nand U12021 (N_12021,N_10140,N_11550);
or U12022 (N_12022,N_9697,N_11839);
nand U12023 (N_12023,N_9652,N_10829);
nand U12024 (N_12024,N_11131,N_9839);
nand U12025 (N_12025,N_11918,N_11635);
or U12026 (N_12026,N_11868,N_9914);
nor U12027 (N_12027,N_11944,N_11698);
nand U12028 (N_12028,N_9183,N_11360);
nor U12029 (N_12029,N_9267,N_10621);
nand U12030 (N_12030,N_10922,N_11556);
nor U12031 (N_12031,N_10571,N_10969);
nor U12032 (N_12032,N_10080,N_10467);
nor U12033 (N_12033,N_11740,N_9010);
nand U12034 (N_12034,N_9131,N_10985);
and U12035 (N_12035,N_9789,N_9989);
or U12036 (N_12036,N_10335,N_10070);
and U12037 (N_12037,N_9113,N_9687);
and U12038 (N_12038,N_10499,N_9816);
or U12039 (N_12039,N_9931,N_11794);
or U12040 (N_12040,N_9881,N_10149);
nand U12041 (N_12041,N_11436,N_10572);
nor U12042 (N_12042,N_10803,N_10048);
nand U12043 (N_12043,N_9598,N_10737);
nand U12044 (N_12044,N_10575,N_9617);
nand U12045 (N_12045,N_11569,N_10645);
nand U12046 (N_12046,N_9074,N_10624);
and U12047 (N_12047,N_9222,N_11820);
and U12048 (N_12048,N_11674,N_9136);
nor U12049 (N_12049,N_11899,N_11156);
or U12050 (N_12050,N_11661,N_10225);
or U12051 (N_12051,N_9485,N_9775);
or U12052 (N_12052,N_11161,N_9525);
nor U12053 (N_12053,N_9063,N_11295);
and U12054 (N_12054,N_10010,N_10868);
nor U12055 (N_12055,N_11330,N_11885);
nand U12056 (N_12056,N_9167,N_10366);
or U12057 (N_12057,N_11645,N_9984);
and U12058 (N_12058,N_10958,N_10461);
or U12059 (N_12059,N_10451,N_9982);
nor U12060 (N_12060,N_11888,N_11694);
or U12061 (N_12061,N_10325,N_10090);
and U12062 (N_12062,N_10518,N_9745);
and U12063 (N_12063,N_11157,N_9466);
nor U12064 (N_12064,N_9472,N_10794);
and U12065 (N_12065,N_11838,N_11408);
or U12066 (N_12066,N_9512,N_11591);
nand U12067 (N_12067,N_9766,N_9952);
nand U12068 (N_12068,N_11276,N_11233);
nor U12069 (N_12069,N_11389,N_10888);
and U12070 (N_12070,N_9702,N_10897);
or U12071 (N_12071,N_11493,N_10283);
or U12072 (N_12072,N_9254,N_11512);
and U12073 (N_12073,N_10084,N_10522);
and U12074 (N_12074,N_11029,N_11334);
nand U12075 (N_12075,N_11614,N_9126);
nor U12076 (N_12076,N_10857,N_11874);
or U12077 (N_12077,N_9056,N_10736);
nand U12078 (N_12078,N_10491,N_10513);
nand U12079 (N_12079,N_10312,N_9871);
or U12080 (N_12080,N_10788,N_11311);
nor U12081 (N_12081,N_9944,N_10960);
or U12082 (N_12082,N_9383,N_10374);
or U12083 (N_12083,N_10432,N_9636);
and U12084 (N_12084,N_11639,N_9635);
and U12085 (N_12085,N_10060,N_11078);
or U12086 (N_12086,N_9451,N_11609);
and U12087 (N_12087,N_9703,N_10347);
and U12088 (N_12088,N_10121,N_10019);
and U12089 (N_12089,N_10183,N_9505);
or U12090 (N_12090,N_9731,N_11087);
nor U12091 (N_12091,N_11842,N_10578);
nor U12092 (N_12092,N_11858,N_11049);
or U12093 (N_12093,N_10005,N_11160);
and U12094 (N_12094,N_10502,N_11691);
and U12095 (N_12095,N_11789,N_11118);
nand U12096 (N_12096,N_10714,N_11807);
and U12097 (N_12097,N_10505,N_11419);
nand U12098 (N_12098,N_10343,N_10870);
nand U12099 (N_12099,N_9061,N_9329);
or U12100 (N_12100,N_9318,N_11343);
nor U12101 (N_12101,N_11172,N_9541);
or U12102 (N_12102,N_9399,N_10229);
nor U12103 (N_12103,N_11997,N_11416);
or U12104 (N_12104,N_10285,N_11222);
or U12105 (N_12105,N_10134,N_11564);
nor U12106 (N_12106,N_11460,N_10342);
nor U12107 (N_12107,N_11745,N_9744);
nand U12108 (N_12108,N_11504,N_10802);
or U12109 (N_12109,N_9592,N_9022);
or U12110 (N_12110,N_11017,N_10246);
and U12111 (N_12111,N_9250,N_10628);
nor U12112 (N_12112,N_11916,N_10963);
nand U12113 (N_12113,N_11604,N_11749);
nand U12114 (N_12114,N_10365,N_10083);
or U12115 (N_12115,N_9749,N_11035);
or U12116 (N_12116,N_10983,N_9033);
nand U12117 (N_12117,N_9282,N_9410);
nand U12118 (N_12118,N_11407,N_9682);
and U12119 (N_12119,N_11865,N_11795);
nor U12120 (N_12120,N_11379,N_9849);
nand U12121 (N_12121,N_11574,N_11266);
nor U12122 (N_12122,N_11421,N_11747);
or U12123 (N_12123,N_10034,N_11475);
nand U12124 (N_12124,N_9715,N_10287);
nor U12125 (N_12125,N_11655,N_11909);
nand U12126 (N_12126,N_9530,N_11299);
and U12127 (N_12127,N_10784,N_9279);
nand U12128 (N_12128,N_11592,N_11787);
and U12129 (N_12129,N_11692,N_11968);
nor U12130 (N_12130,N_9284,N_9760);
and U12131 (N_12131,N_10667,N_11052);
and U12132 (N_12132,N_11353,N_10742);
nor U12133 (N_12133,N_10962,N_11641);
or U12134 (N_12134,N_11991,N_9418);
nand U12135 (N_12135,N_9387,N_11522);
or U12136 (N_12136,N_10176,N_11294);
and U12137 (N_12137,N_9686,N_11676);
or U12138 (N_12138,N_9629,N_11092);
and U12139 (N_12139,N_10031,N_10185);
and U12140 (N_12140,N_11174,N_11077);
or U12141 (N_12141,N_9903,N_10546);
or U12142 (N_12142,N_10727,N_9213);
and U12143 (N_12143,N_9493,N_11859);
nor U12144 (N_12144,N_9967,N_9085);
nor U12145 (N_12145,N_10486,N_10063);
or U12146 (N_12146,N_10406,N_11385);
nor U12147 (N_12147,N_9558,N_11646);
nand U12148 (N_12148,N_11381,N_10977);
and U12149 (N_12149,N_11523,N_11467);
nand U12150 (N_12150,N_9920,N_9091);
nand U12151 (N_12151,N_9726,N_11201);
or U12152 (N_12152,N_11628,N_10047);
and U12153 (N_12153,N_10733,N_11098);
and U12154 (N_12154,N_9513,N_11702);
nand U12155 (N_12155,N_10195,N_10033);
and U12156 (N_12156,N_9564,N_11457);
nor U12157 (N_12157,N_10497,N_9405);
nor U12158 (N_12158,N_11496,N_10867);
nor U12159 (N_12159,N_9298,N_10315);
nor U12160 (N_12160,N_9211,N_9407);
nor U12161 (N_12161,N_10940,N_9151);
and U12162 (N_12162,N_11399,N_11230);
nor U12163 (N_12163,N_10167,N_9495);
and U12164 (N_12164,N_11338,N_10680);
nor U12165 (N_12165,N_10565,N_9794);
nor U12166 (N_12166,N_11666,N_11454);
or U12167 (N_12167,N_10878,N_10649);
and U12168 (N_12168,N_9619,N_11244);
and U12169 (N_12169,N_9909,N_9833);
nor U12170 (N_12170,N_10475,N_9315);
nand U12171 (N_12171,N_11573,N_10282);
and U12172 (N_12172,N_9662,N_11113);
xnor U12173 (N_12173,N_9140,N_10222);
or U12174 (N_12174,N_11624,N_10636);
or U12175 (N_12175,N_9752,N_9452);
nor U12176 (N_12176,N_9311,N_9396);
nor U12177 (N_12177,N_9049,N_10384);
nor U12178 (N_12178,N_10671,N_9884);
and U12179 (N_12179,N_11216,N_9779);
nor U12180 (N_12180,N_11985,N_10120);
nor U12181 (N_12181,N_10852,N_11486);
nand U12182 (N_12182,N_9175,N_11713);
and U12183 (N_12183,N_10494,N_10937);
or U12184 (N_12184,N_9027,N_9976);
nor U12185 (N_12185,N_11701,N_9861);
and U12186 (N_12186,N_10712,N_9954);
and U12187 (N_12187,N_11709,N_10541);
and U12188 (N_12188,N_11786,N_10240);
nand U12189 (N_12189,N_9973,N_10482);
or U12190 (N_12190,N_10827,N_9440);
nor U12191 (N_12191,N_9520,N_10400);
nor U12192 (N_12192,N_11423,N_11028);
and U12193 (N_12193,N_10331,N_10859);
nand U12194 (N_12194,N_10604,N_11283);
and U12195 (N_12195,N_11860,N_10472);
nand U12196 (N_12196,N_11171,N_10840);
nor U12197 (N_12197,N_11324,N_11750);
and U12198 (N_12198,N_9005,N_9004);
nor U12199 (N_12199,N_10007,N_9947);
or U12200 (N_12200,N_9785,N_10532);
or U12201 (N_12201,N_9278,N_9568);
nor U12202 (N_12202,N_11779,N_11083);
nand U12203 (N_12203,N_10068,N_11339);
nor U12204 (N_12204,N_10387,N_11207);
nor U12205 (N_12205,N_10261,N_10825);
nand U12206 (N_12206,N_9623,N_10207);
nor U12207 (N_12207,N_10540,N_10975);
nor U12208 (N_12208,N_11047,N_11341);
or U12209 (N_12209,N_9776,N_11870);
and U12210 (N_12210,N_10114,N_11933);
nand U12211 (N_12211,N_11211,N_9087);
nand U12212 (N_12212,N_9368,N_9292);
nand U12213 (N_12213,N_10364,N_10037);
nor U12214 (N_12214,N_9783,N_10013);
nor U12215 (N_12215,N_10533,N_10317);
and U12216 (N_12216,N_11151,N_9372);
nor U12217 (N_12217,N_11945,N_11042);
or U12218 (N_12218,N_10961,N_9707);
or U12219 (N_12219,N_11760,N_11878);
and U12220 (N_12220,N_10179,N_10218);
or U12221 (N_12221,N_10526,N_10035);
and U12222 (N_12222,N_10110,N_11549);
or U12223 (N_12223,N_10214,N_11815);
nand U12224 (N_12224,N_11154,N_10308);
or U12225 (N_12225,N_11068,N_9806);
nor U12226 (N_12226,N_11956,N_9469);
or U12227 (N_12227,N_9264,N_10855);
nand U12228 (N_12228,N_10421,N_9646);
or U12229 (N_12229,N_9661,N_9412);
and U12230 (N_12230,N_11588,N_11146);
nor U12231 (N_12231,N_10698,N_9538);
nand U12232 (N_12232,N_9274,N_9384);
nor U12233 (N_12233,N_9216,N_11800);
and U12234 (N_12234,N_11148,N_10171);
or U12235 (N_12235,N_10136,N_10147);
and U12236 (N_12236,N_11951,N_9842);
nor U12237 (N_12237,N_11371,N_11848);
and U12238 (N_12238,N_9351,N_9563);
or U12239 (N_12239,N_9470,N_9255);
or U12240 (N_12240,N_9637,N_10133);
and U12241 (N_12241,N_9890,N_9263);
or U12242 (N_12242,N_9089,N_9753);
nor U12243 (N_12243,N_11272,N_11468);
and U12244 (N_12244,N_10675,N_10633);
and U12245 (N_12245,N_10202,N_9559);
and U12246 (N_12246,N_11386,N_11947);
nor U12247 (N_12247,N_10560,N_10326);
and U12248 (N_12248,N_10403,N_10423);
nand U12249 (N_12249,N_9041,N_9077);
nand U12250 (N_12250,N_10724,N_11829);
nand U12251 (N_12251,N_11852,N_10228);
or U12252 (N_12252,N_10641,N_9432);
nand U12253 (N_12253,N_10883,N_11817);
and U12254 (N_12254,N_9992,N_9281);
nand U12255 (N_12255,N_11167,N_11026);
and U12256 (N_12256,N_11595,N_11741);
and U12257 (N_12257,N_9097,N_9373);
nor U12258 (N_12258,N_9215,N_9577);
and U12259 (N_12259,N_9709,N_9117);
or U12260 (N_12260,N_10128,N_11372);
and U12261 (N_12261,N_11875,N_10844);
or U12262 (N_12262,N_10212,N_9523);
nor U12263 (N_12263,N_11206,N_10188);
nor U12264 (N_12264,N_9024,N_11186);
or U12265 (N_12265,N_9247,N_10334);
nand U12266 (N_12266,N_11724,N_11632);
or U12267 (N_12267,N_10757,N_10354);
nand U12268 (N_12268,N_11182,N_9376);
and U12269 (N_12269,N_11205,N_9681);
nor U12270 (N_12270,N_10933,N_10989);
and U12271 (N_12271,N_9916,N_11965);
nand U12272 (N_12272,N_11476,N_11623);
nand U12273 (N_12273,N_11919,N_10694);
nand U12274 (N_12274,N_10337,N_9361);
and U12275 (N_12275,N_9851,N_10748);
and U12276 (N_12276,N_9150,N_11554);
nand U12277 (N_12277,N_11445,N_11722);
and U12278 (N_12278,N_10391,N_9964);
or U12279 (N_12279,N_11889,N_9310);
nand U12280 (N_12280,N_10024,N_10011);
and U12281 (N_12281,N_10169,N_11469);
and U12282 (N_12282,N_10655,N_11364);
nand U12283 (N_12283,N_9060,N_9632);
nand U12284 (N_12284,N_10320,N_10425);
nand U12285 (N_12285,N_9484,N_10510);
nor U12286 (N_12286,N_11253,N_9521);
nor U12287 (N_12287,N_10701,N_9290);
nor U12288 (N_12288,N_11718,N_10886);
and U12289 (N_12289,N_10660,N_9319);
and U12290 (N_12290,N_10992,N_11424);
nor U12291 (N_12291,N_11432,N_11040);
nor U12292 (N_12292,N_11366,N_10367);
nor U12293 (N_12293,N_10890,N_9116);
and U12294 (N_12294,N_10064,N_9506);
nand U12295 (N_12295,N_10664,N_11545);
nor U12296 (N_12296,N_10098,N_11365);
and U12297 (N_12297,N_11477,N_11547);
nor U12298 (N_12298,N_9957,N_9447);
nor U12299 (N_12299,N_9908,N_10725);
and U12300 (N_12300,N_9489,N_10235);
and U12301 (N_12301,N_11001,N_10487);
nand U12302 (N_12302,N_10789,N_11524);
nand U12303 (N_12303,N_11448,N_9999);
nand U12304 (N_12304,N_11530,N_9557);
nor U12305 (N_12305,N_9295,N_10920);
nand U12306 (N_12306,N_9531,N_11672);
or U12307 (N_12307,N_11344,N_9542);
and U12308 (N_12308,N_9346,N_11122);
or U12309 (N_12309,N_9631,N_10051);
nor U12310 (N_12310,N_11950,N_9322);
nand U12311 (N_12311,N_9019,N_9669);
nand U12312 (N_12312,N_10613,N_10914);
nand U12313 (N_12313,N_11952,N_9575);
nand U12314 (N_12314,N_10081,N_10659);
and U12315 (N_12315,N_9585,N_9481);
and U12316 (N_12316,N_10155,N_9743);
nor U12317 (N_12317,N_10061,N_9016);
and U12318 (N_12318,N_9343,N_9667);
and U12319 (N_12319,N_11904,N_10215);
and U12320 (N_12320,N_10602,N_10462);
and U12321 (N_12321,N_9369,N_10708);
or U12322 (N_12322,N_9475,N_9959);
or U12323 (N_12323,N_9257,N_11696);
nor U12324 (N_12324,N_11697,N_9694);
or U12325 (N_12325,N_11836,N_9364);
and U12326 (N_12326,N_10153,N_10818);
and U12327 (N_12327,N_11426,N_10144);
nand U12328 (N_12328,N_9756,N_10180);
or U12329 (N_12329,N_9122,N_11850);
and U12330 (N_12330,N_10590,N_9430);
and U12331 (N_12331,N_9386,N_11136);
nand U12332 (N_12332,N_10699,N_9483);
nand U12333 (N_12333,N_11518,N_10549);
nor U12334 (N_12334,N_11914,N_9170);
and U12335 (N_12335,N_11585,N_11030);
or U12336 (N_12336,N_10516,N_9306);
nand U12337 (N_12337,N_10231,N_10785);
nor U12338 (N_12338,N_9738,N_9428);
and U12339 (N_12339,N_10639,N_10769);
nand U12340 (N_12340,N_10311,N_10453);
nor U12341 (N_12341,N_10952,N_10580);
or U12342 (N_12342,N_10772,N_10836);
and U12343 (N_12343,N_10187,N_11046);
or U12344 (N_12344,N_10924,N_10653);
nand U12345 (N_12345,N_9961,N_11369);
nand U12346 (N_12346,N_11450,N_11743);
nor U12347 (N_12347,N_11902,N_10971);
nor U12348 (N_12348,N_10129,N_11231);
xnor U12349 (N_12349,N_9394,N_11346);
nand U12350 (N_12350,N_10091,N_9268);
or U12351 (N_12351,N_9486,N_9494);
nand U12352 (N_12352,N_9032,N_11123);
nand U12353 (N_12353,N_10608,N_11248);
or U12354 (N_12354,N_10774,N_10126);
nor U12355 (N_12355,N_10324,N_10730);
or U12356 (N_12356,N_11022,N_11106);
nand U12357 (N_12357,N_9784,N_10143);
or U12358 (N_12358,N_9181,N_9101);
nand U12359 (N_12359,N_11663,N_11758);
and U12360 (N_12360,N_9260,N_10361);
and U12361 (N_12361,N_9514,N_10348);
nand U12362 (N_12362,N_11528,N_11915);
or U12363 (N_12363,N_11152,N_10761);
and U12364 (N_12364,N_10766,N_10564);
nand U12365 (N_12365,N_11742,N_11855);
and U12366 (N_12366,N_11159,N_11018);
nand U12367 (N_12367,N_11390,N_10490);
and U12368 (N_12368,N_9972,N_11451);
or U12369 (N_12369,N_9649,N_11459);
nand U12370 (N_12370,N_10747,N_9271);
nand U12371 (N_12371,N_10074,N_9663);
xor U12372 (N_12372,N_9915,N_10591);
and U12373 (N_12373,N_9859,N_11349);
or U12374 (N_12374,N_9630,N_11594);
or U12375 (N_12375,N_9664,N_11605);
nand U12376 (N_12376,N_9273,N_10805);
nor U12377 (N_12377,N_10270,N_10227);
and U12378 (N_12378,N_10473,N_9297);
and U12379 (N_12379,N_9765,N_10431);
nor U12380 (N_12380,N_11084,N_10359);
nand U12381 (N_12381,N_9843,N_11656);
and U12382 (N_12382,N_10955,N_11826);
and U12383 (N_12383,N_11138,N_9611);
xor U12384 (N_12384,N_9650,N_9820);
nand U12385 (N_12385,N_11567,N_11246);
nand U12386 (N_12386,N_10899,N_11150);
nor U12387 (N_12387,N_10456,N_11622);
or U12388 (N_12388,N_10615,N_10731);
and U12389 (N_12389,N_11831,N_9622);
and U12390 (N_12390,N_9473,N_11680);
nand U12391 (N_12391,N_11586,N_10071);
nand U12392 (N_12392,N_11617,N_10452);
xor U12393 (N_12393,N_11402,N_9836);
and U12394 (N_12394,N_11514,N_10589);
nor U12395 (N_12395,N_9404,N_11214);
and U12396 (N_12396,N_9971,N_11380);
or U12397 (N_12397,N_11897,N_9696);
or U12398 (N_12398,N_11089,N_11577);
nor U12399 (N_12399,N_10630,N_11086);
and U12400 (N_12400,N_10078,N_11983);
nor U12401 (N_12401,N_10843,N_11576);
nand U12402 (N_12402,N_9479,N_9353);
nand U12403 (N_12403,N_9038,N_10224);
nand U12404 (N_12404,N_11431,N_10740);
nand U12405 (N_12405,N_9827,N_11583);
and U12406 (N_12406,N_11273,N_10601);
nand U12407 (N_12407,N_10220,N_9928);
nand U12408 (N_12408,N_9933,N_11044);
and U12409 (N_12409,N_9535,N_10131);
and U12410 (N_12410,N_11433,N_10934);
nand U12411 (N_12411,N_10323,N_11218);
and U12412 (N_12412,N_10523,N_10003);
nor U12413 (N_12413,N_9892,N_9571);
xor U12414 (N_12414,N_11793,N_9189);
or U12415 (N_12415,N_10640,N_11797);
nand U12416 (N_12416,N_9922,N_10865);
or U12417 (N_12417,N_11927,N_10854);
nor U12418 (N_12418,N_9730,N_10721);
nand U12419 (N_12419,N_9862,N_10583);
or U12420 (N_12420,N_11562,N_11551);
and U12421 (N_12421,N_10662,N_10539);
xnor U12422 (N_12422,N_9224,N_9453);
or U12423 (N_12423,N_11863,N_11447);
and U12424 (N_12424,N_11715,N_10014);
and U12425 (N_12425,N_10792,N_9732);
or U12426 (N_12426,N_10587,N_10293);
nand U12427 (N_12427,N_11686,N_9621);
nand U12428 (N_12428,N_10668,N_9251);
or U12429 (N_12429,N_10935,N_10237);
nor U12430 (N_12430,N_9478,N_11900);
nand U12431 (N_12431,N_10072,N_11305);
nand U12432 (N_12432,N_11382,N_11401);
or U12433 (N_12433,N_9461,N_9114);
nor U12434 (N_12434,N_9397,N_10446);
or U12435 (N_12435,N_11166,N_9258);
and U12436 (N_12436,N_11315,N_10562);
or U12437 (N_12437,N_11307,N_10422);
and U12438 (N_12438,N_10631,N_11727);
nand U12439 (N_12439,N_10350,N_11880);
and U12440 (N_12440,N_11892,N_9201);
or U12441 (N_12441,N_11144,N_11285);
nor U12442 (N_12442,N_11578,N_9230);
nand U12443 (N_12443,N_9171,N_11356);
nor U12444 (N_12444,N_9786,N_11190);
or U12445 (N_12445,N_9507,N_9269);
nand U12446 (N_12446,N_11261,N_9819);
nand U12447 (N_12447,N_10388,N_11337);
and U12448 (N_12448,N_10500,N_11168);
or U12449 (N_12449,N_9291,N_11263);
nor U12450 (N_12450,N_10450,N_11103);
or U12451 (N_12451,N_9625,N_11194);
or U12452 (N_12452,N_11240,N_10980);
nand U12453 (N_12453,N_9550,N_9082);
and U12454 (N_12454,N_9727,N_10535);
nor U12455 (N_12455,N_9203,N_11809);
or U12456 (N_12456,N_9482,N_11081);
xor U12457 (N_12457,N_11212,N_10125);
nand U12458 (N_12458,N_10162,N_9145);
and U12459 (N_12459,N_9398,N_10874);
and U12460 (N_12460,N_11465,N_9148);
or U12461 (N_12461,N_11660,N_10412);
nand U12462 (N_12462,N_9729,N_11634);
nor U12463 (N_12463,N_9582,N_9093);
nor U12464 (N_12464,N_10846,N_11129);
nor U12465 (N_12465,N_9672,N_10052);
nand U12466 (N_12466,N_11277,N_9380);
and U12467 (N_12467,N_9001,N_11926);
or U12468 (N_12468,N_9831,N_11041);
and U12469 (N_12469,N_11293,N_10069);
or U12470 (N_12470,N_9031,N_11120);
nand U12471 (N_12471,N_9718,N_9324);
nand U12472 (N_12472,N_10612,N_9503);
or U12473 (N_12473,N_9830,N_10988);
nand U12474 (N_12474,N_11967,N_9763);
nor U12475 (N_12475,N_9445,N_10611);
or U12476 (N_12476,N_9228,N_10213);
nand U12477 (N_12477,N_11730,N_10566);
nor U12478 (N_12478,N_11598,N_10307);
nand U12479 (N_12479,N_11388,N_11280);
nor U12480 (N_12480,N_11841,N_10279);
nand U12481 (N_12481,N_10370,N_11670);
xor U12482 (N_12482,N_11746,N_9543);
nor U12483 (N_12483,N_10086,N_9790);
nor U12484 (N_12484,N_11505,N_10161);
and U12485 (N_12485,N_10408,N_9416);
and U12486 (N_12486,N_11529,N_11688);
nand U12487 (N_12487,N_11024,N_11845);
nor U12488 (N_12488,N_10625,N_11267);
nor U12489 (N_12489,N_11527,N_9529);
nand U12490 (N_12490,N_11544,N_10004);
nor U12491 (N_12491,N_9837,N_11125);
nand U12492 (N_12492,N_10809,N_11657);
or U12493 (N_12493,N_11568,N_10349);
nor U12494 (N_12494,N_9722,N_10481);
or U12495 (N_12495,N_9515,N_9302);
nor U12496 (N_12496,N_11056,N_9460);
or U12497 (N_12497,N_11905,N_10206);
and U12498 (N_12498,N_9210,N_9985);
or U12499 (N_12499,N_11378,N_9614);
and U12500 (N_12500,N_9601,N_10561);
nand U12501 (N_12501,N_9246,N_9860);
nand U12502 (N_12502,N_10907,N_9803);
and U12503 (N_12503,N_9534,N_11607);
nor U12504 (N_12504,N_9668,N_9173);
or U12505 (N_12505,N_11893,N_10923);
and U12506 (N_12506,N_10563,N_11415);
nor U12507 (N_12507,N_10638,N_11964);
or U12508 (N_12508,N_10118,N_10036);
and U12509 (N_12509,N_11683,N_9127);
nand U12510 (N_12510,N_10309,N_10586);
nor U12511 (N_12511,N_11020,N_11109);
and U12512 (N_12512,N_9174,N_10108);
and U12513 (N_12513,N_11289,N_11239);
or U12514 (N_12514,N_9457,N_11034);
nand U12515 (N_12515,N_11269,N_10008);
nor U12516 (N_12516,N_10767,N_9873);
and U12517 (N_12517,N_9051,N_10864);
nor U12518 (N_12518,N_11287,N_11478);
and U12519 (N_12519,N_9366,N_9504);
nand U12520 (N_12520,N_11517,N_9880);
nand U12521 (N_12521,N_11636,N_9132);
or U12522 (N_12522,N_11335,N_9708);
and U12523 (N_12523,N_9390,N_9645);
xor U12524 (N_12524,N_9105,N_10635);
and U12525 (N_12525,N_9937,N_11492);
nand U12526 (N_12526,N_10763,N_10913);
or U12527 (N_12527,N_10389,N_10877);
or U12528 (N_12528,N_9047,N_11648);
or U12529 (N_12529,N_9517,N_9782);
nor U12530 (N_12530,N_9234,N_10966);
or U12531 (N_12531,N_10023,N_10170);
and U12532 (N_12532,N_11488,N_9675);
xor U12533 (N_12533,N_9095,N_11310);
xor U12534 (N_12534,N_11179,N_9000);
and U12535 (N_12535,N_11145,N_10697);
and U12536 (N_12536,N_9912,N_9239);
nand U12537 (N_12537,N_9141,N_10651);
nor U12538 (N_12538,N_11254,N_11198);
nor U12539 (N_12539,N_10970,N_11699);
or U12540 (N_12540,N_10558,N_11400);
or U12541 (N_12541,N_9639,N_9283);
or U12542 (N_12542,N_11185,N_9294);
and U12543 (N_12543,N_9879,N_11535);
nand U12544 (N_12544,N_9583,N_11351);
nor U12545 (N_12545,N_10281,N_10470);
or U12546 (N_12546,N_9968,N_11099);
nor U12547 (N_12547,N_10407,N_11191);
or U12548 (N_12548,N_11355,N_10375);
and U12549 (N_12549,N_10726,N_11425);
nor U12550 (N_12550,N_10948,N_9356);
and U12551 (N_12551,N_10909,N_9003);
and U12552 (N_12552,N_11251,N_9423);
or U12553 (N_12553,N_10305,N_10820);
or U12554 (N_12554,N_10076,N_9307);
nor U12555 (N_12555,N_10369,N_11873);
or U12556 (N_12556,N_11543,N_9613);
or U12557 (N_12557,N_10410,N_10976);
nand U12558 (N_12558,N_10816,N_10592);
nor U12559 (N_12559,N_9433,N_11930);
nor U12560 (N_12560,N_11345,N_11911);
or U12561 (N_12561,N_10255,N_10087);
or U12562 (N_12562,N_10559,N_9878);
and U12563 (N_12563,N_9719,N_11940);
nand U12564 (N_12564,N_9088,N_11043);
nor U12565 (N_12565,N_9690,N_10530);
or U12566 (N_12566,N_9325,N_9487);
and U12567 (N_12567,N_10099,N_11590);
or U12568 (N_12568,N_11681,N_9169);
nor U12569 (N_12569,N_9233,N_10900);
nor U12570 (N_12570,N_9855,N_11558);
nand U12571 (N_12571,N_10780,N_10607);
nand U12572 (N_12572,N_10509,N_9802);
or U12573 (N_12573,N_11479,N_11466);
and U12574 (N_12574,N_11966,N_11347);
or U12575 (N_12575,N_10594,N_11005);
or U12576 (N_12576,N_9628,N_9146);
nand U12577 (N_12577,N_11497,N_9219);
nor U12578 (N_12578,N_11960,N_11328);
or U12579 (N_12579,N_11819,N_11177);
and U12580 (N_12580,N_9987,N_10845);
nand U12581 (N_12581,N_10765,N_11252);
nand U12582 (N_12582,N_10947,N_11771);
nand U12583 (N_12583,N_10584,N_10550);
nor U12584 (N_12584,N_10496,N_11935);
or U12585 (N_12585,N_10393,N_9020);
and U12586 (N_12586,N_11255,N_10463);
nor U12587 (N_12587,N_10267,N_9997);
or U12588 (N_12588,N_10191,N_10538);
nor U12589 (N_12589,N_9133,N_11112);
nor U12590 (N_12590,N_10504,N_10710);
nor U12591 (N_12591,N_11602,N_10706);
nand U12592 (N_12592,N_9025,N_10015);
xnor U12593 (N_12593,N_10092,N_9917);
nor U12594 (N_12594,N_10531,N_9787);
nor U12595 (N_12595,N_10148,N_11612);
and U12596 (N_12596,N_11553,N_11766);
and U12597 (N_12597,N_10663,N_11223);
nand U12598 (N_12598,N_10771,N_11397);
and U12599 (N_12599,N_10783,N_10995);
or U12600 (N_12600,N_10097,N_9305);
nor U12601 (N_12601,N_9597,N_10703);
nand U12602 (N_12602,N_9287,N_9442);
and U12603 (N_12603,N_11290,N_9238);
and U12604 (N_12604,N_9034,N_10079);
and U12605 (N_12605,N_11003,N_9017);
or U12606 (N_12606,N_11652,N_11704);
nand U12607 (N_12607,N_10986,N_10095);
or U12608 (N_12608,N_9897,N_10860);
nand U12609 (N_12609,N_10186,N_10908);
nand U12610 (N_12610,N_10953,N_9648);
and U12611 (N_12611,N_11782,N_9710);
or U12612 (N_12612,N_10629,N_11059);
and U12613 (N_12613,N_9064,N_11832);
nor U12614 (N_12614,N_10145,N_9562);
or U12615 (N_12615,N_10260,N_11708);
or U12616 (N_12616,N_10764,N_9317);
and U12617 (N_12617,N_9981,N_10753);
nor U12618 (N_12618,N_11521,N_11257);
xor U12619 (N_12619,N_10398,N_10042);
nor U12620 (N_12620,N_11620,N_10000);
or U12621 (N_12621,N_11494,N_9735);
or U12622 (N_12622,N_11487,N_11716);
and U12623 (N_12623,N_9808,N_11326);
nand U12624 (N_12624,N_9098,N_9924);
and U12625 (N_12625,N_9698,N_10112);
nand U12626 (N_12626,N_10380,N_10959);
or U12627 (N_12627,N_10248,N_9759);
and U12628 (N_12628,N_11931,N_11474);
nand U12629 (N_12629,N_11226,N_10344);
nor U12630 (N_12630,N_9907,N_11955);
nand U12631 (N_12631,N_10073,N_11471);
nor U12632 (N_12632,N_10009,N_9414);
and U12633 (N_12633,N_11582,N_11565);
and U12634 (N_12634,N_11165,N_9092);
and U12635 (N_12635,N_10268,N_11358);
xnor U12636 (N_12636,N_9545,N_9153);
and U12637 (N_12637,N_11606,N_10738);
or U12638 (N_12638,N_10249,N_11164);
and U12639 (N_12639,N_10198,N_11321);
or U12640 (N_12640,N_11835,N_10043);
or U12641 (N_12641,N_10791,N_9377);
nor U12642 (N_12642,N_9026,N_10379);
or U12643 (N_12643,N_10288,N_9330);
and U12644 (N_12644,N_10386,N_10096);
and U12645 (N_12645,N_10142,N_9904);
and U12646 (N_12646,N_11116,N_11629);
nor U12647 (N_12647,N_9081,N_10360);
or U12648 (N_12648,N_9159,N_10987);
nor U12649 (N_12649,N_10626,N_10259);
and U12650 (N_12650,N_11532,N_11303);
nor U12651 (N_12651,N_10906,N_9161);
and U12652 (N_12652,N_9272,N_11943);
and U12653 (N_12653,N_9657,N_9023);
nand U12654 (N_12654,N_10221,N_9328);
nor U12655 (N_12655,N_10290,N_9491);
or U12656 (N_12656,N_11108,N_9573);
xor U12657 (N_12657,N_9381,N_11937);
and U12658 (N_12658,N_10166,N_9918);
nand U12659 (N_12659,N_9750,N_9721);
nand U12660 (N_12660,N_11849,N_10991);
or U12661 (N_12661,N_10442,N_10420);
nor U12662 (N_12662,N_9236,N_10474);
nand U12663 (N_12663,N_11039,N_10674);
nor U12664 (N_12664,N_11406,N_10219);
nand U12665 (N_12665,N_11511,N_10606);
and U12666 (N_12666,N_11271,N_11075);
nor U12667 (N_12667,N_9425,N_9885);
or U12668 (N_12668,N_11088,N_9578);
or U12669 (N_12669,N_9349,N_9716);
nor U12670 (N_12670,N_11220,N_10341);
nor U12671 (N_12671,N_9235,N_9925);
nand U12672 (N_12672,N_10385,N_10256);
and U12673 (N_12673,N_10455,N_9018);
nand U12674 (N_12674,N_9303,N_9832);
nand U12675 (N_12675,N_9883,N_11538);
and U12676 (N_12676,N_9266,N_9913);
nor U12677 (N_12677,N_10704,N_10163);
and U12678 (N_12678,N_9826,N_9755);
or U12679 (N_12679,N_9220,N_10695);
nor U12680 (N_12680,N_10673,N_11265);
and U12681 (N_12681,N_9243,N_9241);
and U12682 (N_12682,N_9352,N_10884);
and U12683 (N_12683,N_9818,N_11278);
nand U12684 (N_12684,N_10045,N_11357);
nor U12685 (N_12685,N_11647,N_11894);
and U12686 (N_12686,N_11903,N_11603);
and U12687 (N_12687,N_11917,N_11176);
or U12688 (N_12688,N_9717,N_9371);
or U12689 (N_12689,N_11954,N_11821);
and U12690 (N_12690,N_11237,N_11354);
or U12691 (N_12691,N_10689,N_10381);
or U12692 (N_12692,N_9184,N_11016);
nor U12693 (N_12693,N_9341,N_10644);
nor U12694 (N_12694,N_9308,N_9316);
and U12695 (N_12695,N_10056,N_10272);
xnor U12696 (N_12696,N_9705,N_9312);
nor U12697 (N_12697,N_10440,N_10094);
nor U12698 (N_12698,N_10599,N_9887);
or U12699 (N_12699,N_9673,N_11710);
or U12700 (N_12700,N_9164,N_9932);
and U12701 (N_12701,N_9355,N_9711);
nor U12702 (N_12702,N_11946,N_11139);
or U12703 (N_12703,N_10372,N_10808);
xnor U12704 (N_12704,N_11352,N_10595);
nor U12705 (N_12705,N_11662,N_11941);
nand U12706 (N_12706,N_11783,N_11440);
nand U12707 (N_12707,N_9121,N_10480);
and U12708 (N_12708,N_11678,N_11519);
nand U12709 (N_12709,N_9758,N_9554);
nor U12710 (N_12710,N_10542,N_9841);
xor U12711 (N_12711,N_9070,N_9796);
and U12712 (N_12712,N_9339,N_9757);
nor U12713 (N_12713,N_10511,N_11158);
and U12714 (N_12714,N_11744,N_10414);
nand U12715 (N_12715,N_9162,N_10882);
nand U12716 (N_12716,N_11679,N_11570);
nand U12717 (N_12717,N_9524,N_10544);
and U12718 (N_12718,N_10429,N_10006);
nor U12719 (N_12719,N_10826,N_10646);
nor U12720 (N_12720,N_9728,N_11404);
nand U12721 (N_12721,N_11631,N_11110);
nor U12722 (N_12722,N_10881,N_10368);
nand U12723 (N_12723,N_11367,N_11427);
nand U12724 (N_12724,N_10318,N_9326);
or U12725 (N_12725,N_11456,N_10469);
nand U12726 (N_12726,N_9156,N_11428);
nand U12727 (N_12727,N_11377,N_10863);
and U12728 (N_12728,N_10336,N_9869);
or U12729 (N_12729,N_9040,N_9701);
nand U12730 (N_12730,N_11563,N_9955);
nand U12731 (N_12731,N_10965,N_9998);
nand U12732 (N_12732,N_11153,N_9979);
or U12733 (N_12733,N_10654,N_9441);
nor U12734 (N_12734,N_11411,N_9817);
nand U12735 (N_12735,N_11667,N_10284);
nor U12736 (N_12736,N_9199,N_11080);
nand U12737 (N_12737,N_11596,N_9655);
and U12738 (N_12738,N_11027,N_11090);
xor U12739 (N_12739,N_11921,N_10686);
and U12740 (N_12740,N_10020,N_11435);
and U12741 (N_12741,N_11728,N_9277);
nand U12742 (N_12742,N_11072,N_11986);
and U12743 (N_12743,N_10459,N_9456);
nor U12744 (N_12744,N_11079,N_10165);
or U12745 (N_12745,N_9570,N_11227);
nand U12746 (N_12746,N_9969,N_10984);
or U12747 (N_12747,N_10002,N_11375);
and U12748 (N_12748,N_11147,N_10158);
and U12749 (N_12749,N_11668,N_9011);
or U12750 (N_12750,N_11503,N_9548);
nand U12751 (N_12751,N_10378,N_9240);
nor U12752 (N_12752,N_11281,N_9895);
and U12753 (N_12753,N_9891,N_9966);
or U12754 (N_12754,N_10433,N_11762);
nor U12755 (N_12755,N_10750,N_10278);
or U12756 (N_12756,N_11613,N_10356);
nand U12757 (N_12757,N_9902,N_11989);
and U12758 (N_12758,N_9299,N_11192);
nor U12759 (N_12759,N_10394,N_11127);
nor U12760 (N_12760,N_9939,N_10658);
nor U12761 (N_12761,N_10880,N_10717);
nor U12762 (N_12762,N_9180,N_10107);
nor U12763 (N_12763,N_10856,N_10978);
and U12764 (N_12764,N_11507,N_9195);
nand U12765 (N_12765,N_11012,N_10454);
and U12766 (N_12766,N_9436,N_11312);
or U12767 (N_12767,N_10294,N_9253);
nor U12768 (N_12768,N_9488,N_10719);
nor U12769 (N_12769,N_11288,N_9596);
nor U12770 (N_12770,N_10746,N_9847);
and U12771 (N_12771,N_10605,N_10263);
or U12772 (N_12772,N_10872,N_9109);
and U12773 (N_12773,N_11788,N_10949);
or U12774 (N_12774,N_9252,N_11199);
or U12775 (N_12775,N_10273,N_10151);
nand U12776 (N_12776,N_9604,N_11589);
or U12777 (N_12777,N_10172,N_9566);
and U12778 (N_12778,N_11370,N_10837);
and U12779 (N_12779,N_11988,N_10813);
and U12780 (N_12780,N_11180,N_11009);
and U12781 (N_12781,N_9963,N_10569);
or U12782 (N_12782,N_9638,N_11498);
and U12783 (N_12783,N_9498,N_9792);
nor U12784 (N_12784,N_11731,N_10781);
or U12785 (N_12785,N_9740,N_9143);
or U12786 (N_12786,N_9012,N_9679);
or U12787 (N_12787,N_11725,N_11300);
nor U12788 (N_12788,N_10116,N_11626);
or U12789 (N_12789,N_10085,N_11387);
or U12790 (N_12790,N_11928,N_11802);
nand U12791 (N_12791,N_9480,N_11515);
nand U12792 (N_12792,N_10291,N_9111);
nand U12793 (N_12793,N_11405,N_9977);
nor U12794 (N_12794,N_10950,N_11178);
and U12795 (N_12795,N_10657,N_10357);
nor U12796 (N_12796,N_11799,N_11259);
and U12797 (N_12797,N_10174,N_10242);
or U12798 (N_12798,N_9683,N_11721);
and U12799 (N_12799,N_10528,N_9894);
nor U12800 (N_12800,N_10444,N_10258);
nor U12801 (N_12801,N_10449,N_9748);
and U12802 (N_12802,N_10426,N_11780);
nor U12803 (N_12803,N_9497,N_11038);
or U12804 (N_12804,N_11331,N_11757);
nor U12805 (N_12805,N_9157,N_10299);
nand U12806 (N_12806,N_9225,N_11204);
nor U12807 (N_12807,N_9462,N_10691);
nand U12808 (N_12808,N_10396,N_10588);
nand U12809 (N_12809,N_9066,N_9761);
nor U12810 (N_12810,N_9810,N_11010);
or U12811 (N_12811,N_9057,N_11659);
nor U12812 (N_12812,N_9045,N_11773);
and U12813 (N_12813,N_11221,N_10545);
nor U12814 (N_12814,N_9039,N_10280);
or U12815 (N_12815,N_9602,N_10916);
or U12816 (N_12816,N_11733,N_10620);
nand U12817 (N_12817,N_9772,N_11429);
nand U12818 (N_12818,N_9187,N_10928);
nor U12819 (N_12819,N_11995,N_9437);
xnor U12820 (N_12820,N_9137,N_10524);
nor U12821 (N_12821,N_11804,N_11882);
and U12822 (N_12822,N_11712,N_9537);
or U12823 (N_12823,N_11461,N_10328);
nand U12824 (N_12824,N_9342,N_11485);
nor U12825 (N_12825,N_11095,N_11264);
nor U12826 (N_12826,N_11876,N_11856);
nand U12827 (N_12827,N_10296,N_9853);
nand U12828 (N_12828,N_10062,N_10457);
nor U12829 (N_12829,N_11409,N_10993);
and U12830 (N_12830,N_11976,N_9949);
and U12831 (N_12831,N_11314,N_10804);
and U12832 (N_12832,N_10775,N_10404);
and U12833 (N_12833,N_9793,N_10492);
nor U12834 (N_12834,N_11458,N_9864);
and U12835 (N_12835,N_9603,N_10682);
nand U12836 (N_12836,N_9633,N_9975);
and U12837 (N_12837,N_9546,N_11071);
and U12838 (N_12838,N_9706,N_11864);
nand U12839 (N_12839,N_9665,N_9205);
or U12840 (N_12840,N_10536,N_11776);
and U12841 (N_12841,N_10021,N_11309);
or U12842 (N_12842,N_9123,N_11363);
or U12843 (N_12843,N_11735,N_9680);
and U12844 (N_12844,N_10812,N_11482);
and U12845 (N_12845,N_10795,N_9641);
xnor U12846 (N_12846,N_11767,N_9560);
nand U12847 (N_12847,N_11291,N_9934);
and U12848 (N_12848,N_10637,N_10758);
nand U12849 (N_12849,N_9134,N_9659);
nand U12850 (N_12850,N_10762,N_9522);
nand U12851 (N_12851,N_10879,N_11225);
or U12852 (N_12852,N_10944,N_11398);
or U12853 (N_12853,N_11649,N_9653);
or U12854 (N_12854,N_9036,N_10203);
or U12855 (N_12855,N_9048,N_11673);
nand U12856 (N_12856,N_10053,N_11051);
nand U12857 (N_12857,N_9185,N_10705);
nand U12858 (N_12858,N_9431,N_11992);
nand U12859 (N_12859,N_11738,N_10430);
and U12860 (N_12860,N_11984,N_9196);
nor U12861 (N_12861,N_9209,N_9978);
and U12862 (N_12862,N_11417,N_10903);
nand U12863 (N_12863,N_10286,N_9795);
xor U12864 (N_12864,N_11359,N_9620);
or U12865 (N_12865,N_10358,N_10399);
nand U12866 (N_12866,N_11830,N_11308);
or U12867 (N_12867,N_10018,N_11923);
and U12868 (N_12868,N_11810,N_10154);
nand U12869 (N_12869,N_11286,N_10885);
and U12870 (N_12870,N_10828,N_9556);
nor U12871 (N_12871,N_9929,N_9950);
or U12872 (N_12872,N_9139,N_9424);
nor U12873 (N_12873,N_11320,N_10917);
nand U12874 (N_12874,N_10841,N_10927);
and U12875 (N_12875,N_11642,N_10519);
or U12876 (N_12876,N_9446,N_9595);
nor U12877 (N_12877,N_11316,N_9858);
or U12878 (N_12878,N_9927,N_9336);
or U12879 (N_12879,N_11270,N_11143);
nor U12880 (N_12880,N_9780,N_10685);
nor U12881 (N_12881,N_10529,N_11000);
and U12882 (N_12882,N_10901,N_9053);
nor U12883 (N_12883,N_9129,N_10102);
and U12884 (N_12884,N_10223,N_11284);
nand U12885 (N_12885,N_10677,N_10130);
or U12886 (N_12886,N_10495,N_9245);
nand U12887 (N_12887,N_9612,N_11183);
xnor U12888 (N_12888,N_9574,N_11193);
nand U12889 (N_12889,N_11217,N_11325);
nand U12890 (N_12890,N_10553,N_10926);
or U12891 (N_12891,N_10200,N_9008);
nand U12892 (N_12892,N_10967,N_11879);
or U12893 (N_12893,N_10445,N_11173);
or U12894 (N_12894,N_11643,N_10032);
and U12895 (N_12895,N_11552,N_10684);
nand U12896 (N_12896,N_11890,N_9459);
xnor U12897 (N_12897,N_9901,N_10059);
or U12898 (N_12898,N_9540,N_11247);
nor U12899 (N_12899,N_9021,N_11137);
nand U12900 (N_12900,N_11872,N_11536);
nor U12901 (N_12901,N_11472,N_11249);
nand U12902 (N_12902,N_10054,N_9551);
nor U12903 (N_12903,N_10339,N_11055);
or U12904 (N_12904,N_9080,N_11329);
nor U12905 (N_12905,N_11546,N_10168);
nor U12906 (N_12906,N_11770,N_11368);
nor U12907 (N_12907,N_9824,N_9943);
nand U12908 (N_12908,N_11058,N_9508);
nor U12909 (N_12909,N_11548,N_10930);
and U12910 (N_12910,N_10355,N_10471);
and U12911 (N_12911,N_11734,N_11803);
or U12912 (N_12912,N_10552,N_10895);
or U12913 (N_12913,N_11533,N_10912);
or U12914 (N_12914,N_9948,N_11298);
and U12915 (N_12915,N_9358,N_11243);
nor U12916 (N_12916,N_10313,N_11228);
and U12917 (N_12917,N_11869,N_11822);
nand U12918 (N_12918,N_9553,N_11232);
nand U12919 (N_12919,N_11163,N_9935);
and U12920 (N_12920,N_9666,N_11908);
or U12921 (N_12921,N_11036,N_9490);
nor U12922 (N_12922,N_11462,N_9112);
and U12923 (N_12923,N_9591,N_11301);
and U12924 (N_12924,N_10373,N_9896);
nand U12925 (N_12925,N_11393,N_9634);
nor U12926 (N_12926,N_10435,N_9110);
and U12927 (N_12927,N_10943,N_9348);
or U12928 (N_12928,N_10848,N_9857);
nand U12929 (N_12929,N_10001,N_11823);
nor U12930 (N_12930,N_10574,N_11537);
or U12931 (N_12931,N_11418,N_9083);
or U12932 (N_12932,N_11384,N_9811);
nor U12933 (N_12933,N_9501,N_10887);
nand U12934 (N_12934,N_10811,N_9676);
or U12935 (N_12935,N_11060,N_10181);
nand U12936 (N_12936,N_9898,N_9624);
nand U12937 (N_12937,N_11818,N_10460);
nand U12938 (N_12938,N_9393,N_10346);
nand U12939 (N_12939,N_9068,N_10493);
nand U12940 (N_12940,N_11559,N_10041);
nor U12941 (N_12941,N_11333,N_10938);
nand U12942 (N_12942,N_11664,N_9443);
or U12943 (N_12943,N_11275,N_10619);
and U12944 (N_12944,N_10543,N_9844);
nand U12945 (N_12945,N_10333,N_11414);
and U12946 (N_12946,N_9742,N_9870);
and U12947 (N_12947,N_9069,N_9800);
or U12948 (N_12948,N_10411,N_9464);
and U12949 (N_12949,N_10115,N_9532);
nor U12950 (N_12950,N_9610,N_10289);
and U12951 (N_12951,N_9838,N_9888);
nand U12952 (N_12952,N_9874,N_11115);
or U12953 (N_12953,N_11814,N_11895);
and U12954 (N_12954,N_11007,N_11064);
or U12955 (N_12955,N_9746,N_10196);
and U12956 (N_12956,N_10427,N_11444);
and U12957 (N_12957,N_11234,N_9166);
or U12958 (N_12958,N_9921,N_10729);
nand U12959 (N_12959,N_9822,N_11140);
and U12960 (N_12960,N_9569,N_11502);
or U12961 (N_12961,N_9762,N_11128);
and U12962 (N_12962,N_9465,N_11974);
nor U12963 (N_12963,N_9685,N_9345);
and U12964 (N_12964,N_9848,N_11065);
or U12965 (N_12965,N_11938,N_9073);
nor U12966 (N_12966,N_10632,N_10209);
nor U12967 (N_12967,N_10990,N_10303);
nand U12968 (N_12968,N_10679,N_10547);
or U12969 (N_12969,N_10057,N_10866);
or U12970 (N_12970,N_10266,N_11682);
and U12971 (N_12971,N_10484,N_9594);
nor U12972 (N_12972,N_11050,N_10514);
nor U12973 (N_12973,N_11499,N_11531);
nand U12974 (N_12974,N_11654,N_9178);
nand U12975 (N_12975,N_11703,N_11453);
and U12976 (N_12976,N_11490,N_9605);
nor U12977 (N_12977,N_11210,N_10447);
or U12978 (N_12978,N_11534,N_10106);
and U12979 (N_12979,N_11891,N_10298);
nor U12980 (N_12980,N_10241,N_11342);
nand U12981 (N_12981,N_10915,N_9670);
nor U12982 (N_12982,N_11119,N_10998);
nand U12983 (N_12983,N_11187,N_10779);
or U12984 (N_12984,N_11304,N_9165);
nand U12985 (N_12985,N_10824,N_9539);
nor U12986 (N_12986,N_10300,N_11229);
and U12987 (N_12987,N_9320,N_10787);
xor U12988 (N_12988,N_9262,N_10243);
and U12989 (N_12989,N_9037,N_10932);
or U12990 (N_12990,N_11282,N_10468);
nand U12991 (N_12991,N_10822,N_10551);
nor U12992 (N_12992,N_9014,N_10623);
or U12993 (N_12993,N_10815,N_11723);
or U12994 (N_12994,N_11772,N_11714);
and U12995 (N_12995,N_9704,N_10642);
or U12996 (N_12996,N_9078,N_10807);
and U12997 (N_12997,N_10858,N_10417);
nand U12998 (N_12998,N_9865,N_10254);
or U12999 (N_12999,N_10264,N_9773);
nand U13000 (N_13000,N_11420,N_11581);
nor U13001 (N_13001,N_11394,N_10190);
and U13002 (N_13002,N_11996,N_9799);
or U13003 (N_13003,N_10548,N_11877);
nand U13004 (N_13004,N_10617,N_9212);
and U13005 (N_13005,N_9942,N_9899);
nand U13006 (N_13006,N_11962,N_11853);
and U13007 (N_13007,N_11455,N_9071);
and U13008 (N_13008,N_10082,N_11262);
or U13009 (N_13009,N_10065,N_9599);
or U13010 (N_13010,N_10537,N_10122);
nand U13011 (N_13011,N_11525,N_11008);
nand U13012 (N_13012,N_9244,N_11980);
nand U13013 (N_13013,N_11141,N_10192);
and U13014 (N_13014,N_9421,N_11637);
nand U13015 (N_13015,N_9242,N_11540);
or U13016 (N_13016,N_11910,N_11748);
and U13017 (N_13017,N_11560,N_9327);
and U13018 (N_13018,N_9956,N_10026);
nor U13019 (N_13019,N_10017,N_9643);
nor U13020 (N_13020,N_10527,N_11048);
nor U13021 (N_13021,N_9854,N_10862);
and U13022 (N_13022,N_11318,N_11707);
nand U13023 (N_13023,N_10478,N_9147);
or U13024 (N_13024,N_10049,N_11019);
and U13025 (N_13025,N_10409,N_9333);
and U13026 (N_13026,N_9103,N_10964);
and U13027 (N_13027,N_10419,N_10276);
nand U13028 (N_13028,N_9510,N_9751);
nand U13029 (N_13029,N_9678,N_10819);
and U13030 (N_13030,N_10745,N_10314);
or U13031 (N_13031,N_10479,N_9226);
or U13032 (N_13032,N_10941,N_11774);
and U13033 (N_13033,N_10111,N_9359);
nor U13034 (N_13034,N_11566,N_9607);
nand U13035 (N_13035,N_9476,N_9689);
nor U13036 (N_13036,N_9953,N_9588);
nor U13037 (N_13037,N_10184,N_10046);
nand U13038 (N_13038,N_9304,N_10585);
and U13039 (N_13039,N_10834,N_11208);
nand U13040 (N_13040,N_10994,N_10175);
and U13041 (N_13041,N_9030,N_11189);
nand U13042 (N_13042,N_10135,N_9829);
nor U13043 (N_13043,N_9382,N_11074);
nand U13044 (N_13044,N_10786,N_9323);
or U13045 (N_13045,N_10676,N_11975);
or U13046 (N_13046,N_11274,N_10839);
and U13047 (N_13047,N_11948,N_10650);
or U13048 (N_13048,N_10798,N_9331);
or U13049 (N_13049,N_9770,N_9938);
and U13050 (N_13050,N_11296,N_11437);
or U13051 (N_13051,N_9700,N_11395);
nor U13052 (N_13052,N_9002,N_10749);
nor U13053 (N_13053,N_10251,N_10105);
and U13054 (N_13054,N_10390,N_10156);
or U13055 (N_13055,N_9347,N_9411);
nor U13056 (N_13056,N_10968,N_10715);
nor U13057 (N_13057,N_11979,N_10801);
and U13058 (N_13058,N_10330,N_10931);
nand U13059 (N_13059,N_11669,N_9256);
or U13060 (N_13060,N_10925,N_10269);
nor U13061 (N_13061,N_11236,N_9725);
or U13062 (N_13062,N_9986,N_10835);
nand U13063 (N_13063,N_11886,N_11939);
nand U13064 (N_13064,N_10075,N_9791);
xnor U13065 (N_13065,N_10012,N_10353);
nor U13066 (N_13066,N_11883,N_10029);
and U13067 (N_13067,N_9090,N_9450);
nor U13068 (N_13068,N_9876,N_9850);
nand U13069 (N_13069,N_10954,N_9962);
nand U13070 (N_13070,N_11765,N_11982);
nand U13071 (N_13071,N_9660,N_10150);
nand U13072 (N_13072,N_10891,N_9248);
and U13073 (N_13073,N_9936,N_10239);
nand U13074 (N_13074,N_9572,N_9138);
nor U13075 (N_13075,N_9454,N_10428);
or U13076 (N_13076,N_11392,N_11759);
nand U13077 (N_13077,N_9834,N_11901);
or U13078 (N_13078,N_10782,N_11149);
nand U13079 (N_13079,N_10515,N_11920);
nor U13080 (N_13080,N_10138,N_11235);
nor U13081 (N_13081,N_10756,N_10573);
or U13082 (N_13082,N_11013,N_9378);
and U13083 (N_13083,N_11126,N_10951);
or U13084 (N_13084,N_9403,N_11658);
and U13085 (N_13085,N_11932,N_9163);
nand U13086 (N_13086,N_9875,N_11862);
and U13087 (N_13087,N_11684,N_10665);
nand U13088 (N_13088,N_11689,N_9946);
nor U13089 (N_13089,N_11621,N_11063);
or U13090 (N_13090,N_11857,N_11542);
and U13091 (N_13091,N_9084,N_9449);
nor U13092 (N_13092,N_9699,N_11575);
nand U13093 (N_13093,N_11383,N_9846);
and U13094 (N_13094,N_11102,N_9724);
or U13095 (N_13095,N_11219,N_10058);
nand U13096 (N_13096,N_11963,N_11610);
and U13097 (N_13097,N_9995,N_11031);
and U13098 (N_13098,N_11332,N_11133);
nor U13099 (N_13099,N_11619,N_11484);
or U13100 (N_13100,N_11069,N_11959);
nand U13101 (N_13101,N_9125,N_9567);
nand U13102 (N_13102,N_11695,N_11640);
nand U13103 (N_13103,N_11256,N_11054);
nor U13104 (N_13104,N_11037,N_9994);
or U13105 (N_13105,N_10395,N_9075);
nor U13106 (N_13106,N_9190,N_10582);
nor U13107 (N_13107,N_9695,N_9951);
or U13108 (N_13108,N_9677,N_11053);
nand U13109 (N_13109,N_10301,N_10177);
or U13110 (N_13110,N_10508,N_10055);
and U13111 (N_13111,N_9769,N_11906);
or U13112 (N_13112,N_9774,N_9192);
or U13113 (N_13113,N_10688,N_11720);
nor U13114 (N_13114,N_9406,N_10448);
and U13115 (N_13115,N_10849,N_11805);
nand U13116 (N_13116,N_11162,N_10696);
or U13117 (N_13117,N_10713,N_11463);
or U13118 (N_13118,N_9232,N_11808);
nor U13119 (N_13119,N_9739,N_10332);
nor U13120 (N_13120,N_10234,N_9500);
nor U13121 (N_13121,N_11209,N_10760);
nor U13122 (N_13122,N_10918,N_11827);
and U13123 (N_13123,N_10942,N_11197);
nand U13124 (N_13124,N_9214,N_9094);
or U13125 (N_13125,N_10109,N_11706);
and U13126 (N_13126,N_9813,N_9733);
and U13127 (N_13127,N_9777,N_10902);
and U13128 (N_13128,N_9767,N_9910);
nand U13129 (N_13129,N_11618,N_9863);
or U13130 (N_13130,N_9642,N_10739);
or U13131 (N_13131,N_9439,N_10476);
nand U13132 (N_13132,N_11675,N_10022);
nand U13133 (N_13133,N_11687,N_10100);
or U13134 (N_13134,N_11557,N_10066);
nor U13135 (N_13135,N_10982,N_10503);
or U13136 (N_13136,N_10997,N_11452);
xnor U13137 (N_13137,N_10981,N_10443);
and U13138 (N_13138,N_9221,N_11196);
or U13139 (N_13139,N_10199,N_10132);
nand U13140 (N_13140,N_10622,N_9229);
nand U13141 (N_13141,N_9945,N_10236);
nor U13142 (N_13142,N_10274,N_10322);
and U13143 (N_13143,N_9468,N_11705);
and U13144 (N_13144,N_9552,N_11396);
nor U13145 (N_13145,N_11847,N_10089);
and U13146 (N_13146,N_10797,N_11572);
nand U13147 (N_13147,N_9035,N_10732);
nor U13148 (N_13148,N_9072,N_9674);
nand U13149 (N_13149,N_9429,N_11833);
and U13150 (N_13150,N_11913,N_9593);
nor U13151 (N_13151,N_10773,N_9720);
nand U13152 (N_13152,N_11685,N_10201);
and U13153 (N_13153,N_10146,N_9009);
nor U13154 (N_13154,N_9270,N_10173);
or U13155 (N_13155,N_10904,N_11322);
and U13156 (N_13156,N_9590,N_11002);
nor U13157 (N_13157,N_10465,N_11665);
and U13158 (N_13158,N_11763,N_10275);
and U13159 (N_13159,N_10093,N_9204);
nor U13160 (N_13160,N_9197,N_11446);
nor U13161 (N_13161,N_10402,N_11169);
and U13162 (N_13162,N_11319,N_10050);
or U13163 (N_13163,N_11439,N_11513);
nand U13164 (N_13164,N_9200,N_10669);
nor U13165 (N_13165,N_10262,N_10466);
nand U13166 (N_13166,N_9309,N_10643);
nor U13167 (N_13167,N_10434,N_9237);
nand U13168 (N_13168,N_9202,N_10040);
or U13169 (N_13169,N_10489,N_9941);
nand U13170 (N_13170,N_9261,N_11970);
and U13171 (N_13171,N_11837,N_10929);
and U13172 (N_13172,N_10609,N_9471);
nor U13173 (N_13173,N_10271,N_11999);
nor U13174 (N_13174,N_9389,N_9467);
nand U13175 (N_13175,N_11754,N_9362);
nor U13176 (N_13176,N_11134,N_10693);
nand U13177 (N_13177,N_11121,N_9354);
nor U13178 (N_13178,N_9809,N_9144);
nand U13179 (N_13179,N_10905,N_9872);
nand U13180 (N_13180,N_11242,N_10233);
nand U13181 (N_13181,N_10257,N_9198);
nor U13182 (N_13182,N_10405,N_9801);
nand U13183 (N_13183,N_9344,N_9259);
and U13184 (N_13184,N_9363,N_9374);
nor U13185 (N_13185,N_10329,N_10894);
nor U13186 (N_13186,N_11076,N_11489);
nor U13187 (N_13187,N_9172,N_9606);
nand U13188 (N_13188,N_11245,N_10876);
or U13189 (N_13189,N_9608,N_11491);
nand U13190 (N_13190,N_11279,N_9417);
and U13191 (N_13191,N_11014,N_10720);
xor U13192 (N_13192,N_11470,N_11340);
and U13193 (N_13193,N_9868,N_9768);
and U13194 (N_13194,N_10557,N_10424);
or U13195 (N_13195,N_10683,N_10418);
nand U13196 (N_13196,N_9158,N_9940);
xor U13197 (N_13197,N_11971,N_10576);
nor U13198 (N_13198,N_11070,N_9723);
or U13199 (N_13199,N_10244,N_9527);
or U13200 (N_13200,N_11812,N_9889);
or U13201 (N_13201,N_11778,N_9609);
nor U13202 (N_13202,N_10124,N_9734);
or U13203 (N_13203,N_10700,N_11690);
nor U13204 (N_13204,N_10833,N_11006);
or U13205 (N_13205,N_10464,N_10483);
nand U13206 (N_13206,N_11213,N_9671);
or U13207 (N_13207,N_10896,N_10439);
or U13208 (N_13208,N_9991,N_11924);
nor U13209 (N_13209,N_10800,N_11032);
nor U13210 (N_13210,N_11508,N_9458);
nor U13211 (N_13211,N_11608,N_10345);
or U13212 (N_13212,N_9043,N_11597);
nor U13213 (N_13213,N_9055,N_9096);
nand U13214 (N_13214,N_11501,N_9804);
or U13215 (N_13215,N_10316,N_10253);
nor U13216 (N_13216,N_9079,N_9741);
or U13217 (N_13217,N_10310,N_11600);
nand U13218 (N_13218,N_9519,N_11949);
xor U13219 (N_13219,N_11323,N_10525);
and U13220 (N_13220,N_11336,N_10507);
or U13221 (N_13221,N_11961,N_11993);
or U13222 (N_13222,N_10754,N_11114);
nand U13223 (N_13223,N_11464,N_10627);
nand U13224 (N_13224,N_9249,N_11292);
nand U13225 (N_13225,N_10593,N_9856);
and U13226 (N_13226,N_9338,N_9561);
nor U13227 (N_13227,N_11373,N_11516);
and U13228 (N_13228,N_9544,N_9900);
or U13229 (N_13229,N_11495,N_11925);
nand U13230 (N_13230,N_10067,N_10488);
or U13231 (N_13231,N_9217,N_11729);
nor U13232 (N_13232,N_10743,N_10616);
nand U13233 (N_13233,N_9086,N_11973);
nor U13234 (N_13234,N_11825,N_9408);
nand U13235 (N_13235,N_9516,N_10702);
and U13236 (N_13236,N_9547,N_9191);
nor U13237 (N_13237,N_9905,N_11442);
or U13238 (N_13238,N_9930,N_9124);
nor U13239 (N_13239,N_9208,N_9118);
and U13240 (N_13240,N_9218,N_10799);
and U13241 (N_13241,N_11260,N_9536);
and U13242 (N_13242,N_9142,N_10996);
nand U13243 (N_13243,N_11085,N_10957);
nand U13244 (N_13244,N_9149,N_9576);
and U13245 (N_13245,N_11430,N_11520);
nor U13246 (N_13246,N_11907,N_11184);
or U13247 (N_13247,N_9400,N_10681);
or U13248 (N_13248,N_10351,N_11719);
and U13249 (N_13249,N_10568,N_10796);
and U13250 (N_13250,N_11784,N_9580);
nor U13251 (N_13251,N_9926,N_10838);
and U13252 (N_13252,N_9332,N_10139);
nor U13253 (N_13253,N_11717,N_9193);
xor U13254 (N_13254,N_10567,N_11506);
nor U13255 (N_13255,N_9474,N_11942);
nor U13256 (N_13256,N_9970,N_11480);
nand U13257 (N_13257,N_11181,N_11627);
nand U13258 (N_13258,N_9778,N_9747);
and U13259 (N_13259,N_11130,N_11755);
and U13260 (N_13260,N_9160,N_10647);
and U13261 (N_13261,N_10556,N_11111);
or U13262 (N_13262,N_11978,N_9828);
and U13263 (N_13263,N_11066,N_11633);
nor U13264 (N_13264,N_10377,N_9231);
or U13265 (N_13265,N_10999,N_11887);
nor U13266 (N_13266,N_9438,N_10716);
nand U13267 (N_13267,N_9958,N_9015);
and U13268 (N_13268,N_10416,N_10245);
and U13269 (N_13269,N_9781,N_9365);
and U13270 (N_13270,N_11816,N_11361);
nor U13271 (N_13271,N_11541,N_11611);
nor U13272 (N_13272,N_9814,N_9821);
xor U13273 (N_13273,N_9102,N_10157);
or U13274 (N_13274,N_9321,N_9499);
nor U13275 (N_13275,N_10810,N_10728);
nand U13276 (N_13276,N_9511,N_11650);
or U13277 (N_13277,N_11241,N_10383);
nor U13278 (N_13278,N_9340,N_10759);
nor U13279 (N_13279,N_9044,N_11796);
and U13280 (N_13280,N_9223,N_9422);
and U13281 (N_13281,N_11752,N_9293);
or U13282 (N_13282,N_9067,N_9337);
nand U13283 (N_13283,N_10972,N_11004);
nor U13284 (N_13284,N_11615,N_9413);
nor U13285 (N_13285,N_10911,N_9100);
and U13286 (N_13286,N_10247,N_11025);
nor U13287 (N_13287,N_9155,N_10871);
or U13288 (N_13288,N_11091,N_10718);
nand U13289 (N_13289,N_9385,N_11374);
and U13290 (N_13290,N_11990,N_9227);
or U13291 (N_13291,N_10127,N_11644);
or U13292 (N_13292,N_10189,N_11625);
nor U13293 (N_13293,N_10517,N_10600);
nor U13294 (N_13294,N_9960,N_11376);
nor U13295 (N_13295,N_10847,N_11434);
nand U13296 (N_13296,N_9179,N_9402);
and U13297 (N_13297,N_10793,N_9194);
or U13298 (N_13298,N_11884,N_11958);
or U13299 (N_13299,N_9104,N_11258);
and U13300 (N_13300,N_9419,N_10806);
nor U13301 (N_13301,N_9426,N_10141);
and U13302 (N_13302,N_11526,N_9965);
nor U13303 (N_13303,N_10744,N_11175);
and U13304 (N_13304,N_11756,N_10230);
nor U13305 (N_13305,N_9065,N_11362);
and U13306 (N_13306,N_10520,N_10226);
or U13307 (N_13307,N_10752,N_9852);
and U13308 (N_13308,N_9807,N_9589);
nor U13309 (N_13309,N_11593,N_11693);
or U13310 (N_13310,N_9651,N_10875);
or U13311 (N_13311,N_11441,N_11107);
nor U13312 (N_13312,N_9988,N_11957);
or U13313 (N_13313,N_9658,N_11033);
or U13314 (N_13314,N_10376,N_11202);
and U13315 (N_13315,N_9046,N_11846);
nand U13316 (N_13316,N_11100,N_10306);
nor U13317 (N_13317,N_11736,N_11067);
and U13318 (N_13318,N_10618,N_11737);
or U13319 (N_13319,N_10893,N_10707);
or U13320 (N_13320,N_10117,N_10755);
and U13321 (N_13321,N_11135,N_11155);
and U13322 (N_13322,N_10534,N_11481);
nand U13323 (N_13323,N_11775,N_9823);
nor U13324 (N_13324,N_11806,N_9616);
nor U13325 (N_13325,N_11142,N_10104);
nand U13326 (N_13326,N_9618,N_10919);
or U13327 (N_13327,N_9301,N_11922);
and U13328 (N_13328,N_11677,N_11306);
and U13329 (N_13329,N_9054,N_10216);
nor U13330 (N_13330,N_11132,N_9518);
nor U13331 (N_13331,N_10521,N_9867);
and U13332 (N_13332,N_9586,N_10936);
nor U13333 (N_13333,N_9108,N_11045);
nor U13334 (N_13334,N_9825,N_11987);
nand U13335 (N_13335,N_9654,N_9692);
nand U13336 (N_13336,N_9006,N_9420);
nor U13337 (N_13337,N_9877,N_9115);
nor U13338 (N_13338,N_10741,N_10304);
or U13339 (N_13339,N_9367,N_10709);
nand U13340 (N_13340,N_9714,N_10182);
and U13341 (N_13341,N_11851,N_10295);
or U13342 (N_13342,N_10973,N_9409);
and U13343 (N_13343,N_11093,N_11170);
nor U13344 (N_13344,N_11584,N_9280);
nor U13345 (N_13345,N_10044,N_11438);
nand U13346 (N_13346,N_9528,N_10555);
and U13347 (N_13347,N_9615,N_10252);
nor U13348 (N_13348,N_9923,N_9289);
or U13349 (N_13349,N_10340,N_11410);
nand U13350 (N_13350,N_10211,N_10077);
nand U13351 (N_13351,N_10570,N_11413);
and U13352 (N_13352,N_9058,N_9906);
nand U13353 (N_13353,N_9771,N_10160);
and U13354 (N_13354,N_9427,N_9029);
or U13355 (N_13355,N_9502,N_9300);
and U13356 (N_13356,N_9911,N_11934);
nand U13357 (N_13357,N_11104,N_10842);
or U13358 (N_13358,N_10579,N_10814);
nor U13359 (N_13359,N_11898,N_9062);
nor U13360 (N_13360,N_9980,N_10790);
nor U13361 (N_13361,N_9691,N_10362);
nor U13362 (N_13362,N_10889,N_10210);
nand U13363 (N_13363,N_11313,N_9335);
or U13364 (N_13364,N_9313,N_9581);
nor U13365 (N_13365,N_11843,N_11764);
nor U13366 (N_13366,N_11753,N_10485);
and U13367 (N_13367,N_11861,N_9013);
nand U13368 (N_13368,N_10217,N_9492);
and U13369 (N_13369,N_10397,N_9463);
nand U13370 (N_13370,N_9276,N_10137);
nand U13371 (N_13371,N_10692,N_9983);
nand U13372 (N_13372,N_10401,N_10038);
nand U13373 (N_13373,N_11021,N_10119);
and U13374 (N_13374,N_9275,N_9627);
or U13375 (N_13375,N_9656,N_10751);
and U13376 (N_13376,N_9990,N_10614);
nand U13377 (N_13377,N_9565,N_10596);
or U13378 (N_13378,N_9370,N_11630);
and U13379 (N_13379,N_9207,N_10039);
and U13380 (N_13380,N_11473,N_11509);
nand U13381 (N_13381,N_10415,N_9496);
and U13382 (N_13382,N_9587,N_10821);
nand U13383 (N_13383,N_10027,N_10113);
nor U13384 (N_13384,N_10873,N_9288);
or U13385 (N_13385,N_9434,N_11981);
or U13386 (N_13386,N_10352,N_9285);
nor U13387 (N_13387,N_9788,N_10554);
or U13388 (N_13388,N_11539,N_11327);
or U13389 (N_13389,N_11792,N_11726);
nor U13390 (N_13390,N_10319,N_11653);
nor U13391 (N_13391,N_11854,N_11866);
or U13392 (N_13392,N_9186,N_11015);
nand U13393 (N_13393,N_11510,N_9401);
or U13394 (N_13394,N_9206,N_10735);
or U13395 (N_13395,N_9835,N_11124);
nand U13396 (N_13396,N_11500,N_9647);
or U13397 (N_13397,N_10711,N_9797);
and U13398 (N_13398,N_9533,N_11972);
or U13399 (N_13399,N_9188,N_9357);
nand U13400 (N_13400,N_10204,N_10853);
nor U13401 (N_13401,N_11297,N_9379);
nand U13402 (N_13402,N_10101,N_10194);
or U13403 (N_13403,N_9640,N_10670);
nand U13404 (N_13404,N_11638,N_10581);
nor U13405 (N_13405,N_10088,N_11571);
nor U13406 (N_13406,N_9350,N_11023);
nand U13407 (N_13407,N_9106,N_10178);
and U13408 (N_13408,N_9177,N_11769);
nand U13409 (N_13409,N_9579,N_10205);
nand U13410 (N_13410,N_10722,N_9893);
nor U13411 (N_13411,N_10898,N_11302);
or U13412 (N_13412,N_10277,N_11998);
and U13413 (N_13413,N_9050,N_11828);
nand U13414 (N_13414,N_11651,N_11268);
nor U13415 (N_13415,N_11969,N_9549);
nand U13416 (N_13416,N_9152,N_9059);
nor U13417 (N_13417,N_11579,N_10634);
or U13418 (N_13418,N_9644,N_9974);
or U13419 (N_13419,N_9314,N_11188);
or U13420 (N_13420,N_11811,N_9712);
nor U13421 (N_13421,N_9415,N_11082);
and U13422 (N_13422,N_9688,N_11768);
or U13423 (N_13423,N_10577,N_11561);
nand U13424 (N_13424,N_9455,N_10610);
and U13425 (N_13425,N_10016,N_11403);
and U13426 (N_13426,N_10477,N_10661);
or U13427 (N_13427,N_11867,N_11195);
or U13428 (N_13428,N_11250,N_9130);
and U13429 (N_13429,N_10687,N_10892);
or U13430 (N_13430,N_11801,N_10438);
and U13431 (N_13431,N_11061,N_10238);
and U13432 (N_13432,N_9052,N_9996);
nor U13433 (N_13433,N_11105,N_10152);
nor U13434 (N_13434,N_9866,N_9107);
and U13435 (N_13435,N_11443,N_11824);
or U13436 (N_13436,N_10030,N_10656);
or U13437 (N_13437,N_11555,N_11953);
and U13438 (N_13438,N_11785,N_11599);
nor U13439 (N_13439,N_10603,N_10028);
and U13440 (N_13440,N_10777,N_9154);
and U13441 (N_13441,N_10979,N_10946);
or U13442 (N_13442,N_9296,N_10363);
nand U13443 (N_13443,N_9028,N_11936);
or U13444 (N_13444,N_11203,N_9713);
nand U13445 (N_13445,N_9099,N_11912);
and U13446 (N_13446,N_10869,N_10778);
nand U13447 (N_13447,N_9764,N_11011);
or U13448 (N_13448,N_10025,N_10851);
or U13449 (N_13449,N_10292,N_9626);
nor U13450 (N_13450,N_10512,N_10910);
and U13451 (N_13451,N_10382,N_9798);
or U13452 (N_13452,N_11238,N_10193);
and U13453 (N_13453,N_10666,N_10159);
nor U13454 (N_13454,N_9815,N_9119);
and U13455 (N_13455,N_9120,N_10498);
and U13456 (N_13456,N_9042,N_11790);
or U13457 (N_13457,N_10974,N_11096);
and U13458 (N_13458,N_11348,N_11834);
nand U13459 (N_13459,N_10232,N_11798);
nor U13460 (N_13460,N_11200,N_11391);
or U13461 (N_13461,N_9736,N_9555);
nor U13462 (N_13462,N_10413,N_11062);
nor U13463 (N_13463,N_11791,N_10939);
or U13464 (N_13464,N_11580,N_9076);
nand U13465 (N_13465,N_11601,N_11781);
nand U13466 (N_13466,N_9448,N_9693);
nor U13467 (N_13467,N_11732,N_11751);
nor U13468 (N_13468,N_10265,N_10832);
or U13469 (N_13469,N_10770,N_10831);
and U13470 (N_13470,N_10437,N_10823);
nor U13471 (N_13471,N_11094,N_11412);
or U13472 (N_13472,N_9737,N_11761);
or U13473 (N_13473,N_9360,N_11929);
nand U13474 (N_13474,N_10197,N_10597);
nor U13475 (N_13475,N_10208,N_9805);
nand U13476 (N_13476,N_9395,N_10302);
nor U13477 (N_13477,N_9435,N_11777);
nand U13478 (N_13478,N_11117,N_10690);
or U13479 (N_13479,N_9176,N_9754);
xnor U13480 (N_13480,N_11739,N_10250);
nor U13481 (N_13481,N_9526,N_10672);
or U13482 (N_13482,N_10652,N_11671);
or U13483 (N_13483,N_11449,N_11101);
or U13484 (N_13484,N_11813,N_9812);
and U13485 (N_13485,N_10830,N_9600);
or U13486 (N_13486,N_11587,N_10921);
nand U13487 (N_13487,N_10436,N_10768);
xor U13488 (N_13488,N_11700,N_9477);
nor U13489 (N_13489,N_9286,N_10956);
nand U13490 (N_13490,N_10103,N_10297);
or U13491 (N_13491,N_9882,N_9684);
or U13492 (N_13492,N_11350,N_11881);
nand U13493 (N_13493,N_9993,N_9392);
or U13494 (N_13494,N_10817,N_9334);
and U13495 (N_13495,N_11224,N_11844);
or U13496 (N_13496,N_9375,N_10734);
and U13497 (N_13497,N_10123,N_10598);
nand U13498 (N_13498,N_11871,N_10861);
and U13499 (N_13499,N_10338,N_10850);
or U13500 (N_13500,N_11028,N_9130);
nor U13501 (N_13501,N_11300,N_9376);
and U13502 (N_13502,N_11756,N_10521);
nand U13503 (N_13503,N_11439,N_11777);
nor U13504 (N_13504,N_10467,N_10885);
nor U13505 (N_13505,N_11447,N_11963);
and U13506 (N_13506,N_9525,N_10863);
nand U13507 (N_13507,N_11089,N_11049);
or U13508 (N_13508,N_11398,N_9965);
nand U13509 (N_13509,N_10091,N_10548);
nor U13510 (N_13510,N_9633,N_11858);
or U13511 (N_13511,N_9676,N_9661);
and U13512 (N_13512,N_9828,N_9021);
nor U13513 (N_13513,N_9521,N_9183);
nor U13514 (N_13514,N_9906,N_9494);
or U13515 (N_13515,N_11261,N_11927);
or U13516 (N_13516,N_11294,N_9889);
and U13517 (N_13517,N_9996,N_10681);
nor U13518 (N_13518,N_10098,N_11692);
and U13519 (N_13519,N_10639,N_11737);
and U13520 (N_13520,N_9222,N_11073);
or U13521 (N_13521,N_11964,N_9123);
nor U13522 (N_13522,N_10140,N_11497);
nand U13523 (N_13523,N_10185,N_9210);
nand U13524 (N_13524,N_11919,N_10534);
nor U13525 (N_13525,N_10187,N_9187);
or U13526 (N_13526,N_10549,N_10895);
nand U13527 (N_13527,N_10204,N_11878);
and U13528 (N_13528,N_10572,N_11980);
nor U13529 (N_13529,N_11353,N_9339);
or U13530 (N_13530,N_10793,N_11995);
or U13531 (N_13531,N_9434,N_11483);
nor U13532 (N_13532,N_10929,N_9751);
or U13533 (N_13533,N_10044,N_9376);
nand U13534 (N_13534,N_9475,N_9181);
nor U13535 (N_13535,N_10306,N_11525);
nand U13536 (N_13536,N_9823,N_9950);
nand U13537 (N_13537,N_9651,N_9364);
or U13538 (N_13538,N_9966,N_9898);
and U13539 (N_13539,N_9688,N_10276);
or U13540 (N_13540,N_10893,N_11164);
nor U13541 (N_13541,N_9522,N_9446);
nor U13542 (N_13542,N_10205,N_11748);
or U13543 (N_13543,N_11837,N_10786);
and U13544 (N_13544,N_9489,N_11079);
or U13545 (N_13545,N_9940,N_10560);
nand U13546 (N_13546,N_9332,N_11502);
nand U13547 (N_13547,N_11062,N_9399);
nor U13548 (N_13548,N_10925,N_11901);
or U13549 (N_13549,N_10050,N_9354);
nor U13550 (N_13550,N_10842,N_9847);
and U13551 (N_13551,N_11617,N_11881);
nand U13552 (N_13552,N_9964,N_9493);
or U13553 (N_13553,N_11035,N_11870);
nand U13554 (N_13554,N_9656,N_10486);
nor U13555 (N_13555,N_11994,N_11578);
and U13556 (N_13556,N_9016,N_9270);
and U13557 (N_13557,N_11910,N_9513);
nor U13558 (N_13558,N_9228,N_9488);
and U13559 (N_13559,N_9139,N_11479);
nor U13560 (N_13560,N_9426,N_9494);
and U13561 (N_13561,N_10715,N_11861);
and U13562 (N_13562,N_10117,N_10052);
or U13563 (N_13563,N_9584,N_10838);
nand U13564 (N_13564,N_11416,N_11576);
nor U13565 (N_13565,N_9862,N_10258);
nand U13566 (N_13566,N_9593,N_10539);
nand U13567 (N_13567,N_11872,N_11736);
or U13568 (N_13568,N_9183,N_10693);
nor U13569 (N_13569,N_11753,N_11213);
nand U13570 (N_13570,N_10941,N_11866);
nor U13571 (N_13571,N_9953,N_10289);
nand U13572 (N_13572,N_10799,N_11625);
or U13573 (N_13573,N_11600,N_11555);
and U13574 (N_13574,N_11589,N_10376);
and U13575 (N_13575,N_10017,N_9985);
and U13576 (N_13576,N_9832,N_9392);
or U13577 (N_13577,N_10462,N_9482);
or U13578 (N_13578,N_10074,N_11273);
and U13579 (N_13579,N_9795,N_9183);
and U13580 (N_13580,N_10655,N_11647);
or U13581 (N_13581,N_9627,N_9775);
and U13582 (N_13582,N_10724,N_10944);
nor U13583 (N_13583,N_9707,N_9371);
nand U13584 (N_13584,N_11620,N_10128);
and U13585 (N_13585,N_10333,N_9763);
and U13586 (N_13586,N_9645,N_9318);
and U13587 (N_13587,N_10180,N_11305);
and U13588 (N_13588,N_10570,N_10535);
or U13589 (N_13589,N_9631,N_9024);
nor U13590 (N_13590,N_10768,N_11078);
nor U13591 (N_13591,N_11486,N_9804);
nand U13592 (N_13592,N_10554,N_11429);
and U13593 (N_13593,N_9547,N_9439);
nor U13594 (N_13594,N_11162,N_11927);
nor U13595 (N_13595,N_10147,N_11349);
and U13596 (N_13596,N_10578,N_11368);
nor U13597 (N_13597,N_9029,N_9369);
and U13598 (N_13598,N_9641,N_11576);
and U13599 (N_13599,N_11692,N_10648);
xor U13600 (N_13600,N_10014,N_9153);
nand U13601 (N_13601,N_11611,N_11369);
nor U13602 (N_13602,N_11178,N_10035);
and U13603 (N_13603,N_11613,N_11516);
nor U13604 (N_13604,N_10833,N_11894);
and U13605 (N_13605,N_11708,N_10664);
or U13606 (N_13606,N_11979,N_10087);
nor U13607 (N_13607,N_9929,N_11145);
or U13608 (N_13608,N_10795,N_10986);
and U13609 (N_13609,N_11264,N_11754);
nor U13610 (N_13610,N_10438,N_9937);
or U13611 (N_13611,N_9101,N_11920);
and U13612 (N_13612,N_11611,N_9575);
and U13613 (N_13613,N_10534,N_9822);
and U13614 (N_13614,N_9005,N_9568);
nor U13615 (N_13615,N_11358,N_11929);
nor U13616 (N_13616,N_9025,N_10951);
or U13617 (N_13617,N_9518,N_10184);
nand U13618 (N_13618,N_11142,N_9274);
and U13619 (N_13619,N_9787,N_9777);
and U13620 (N_13620,N_10247,N_9020);
nor U13621 (N_13621,N_9690,N_11874);
and U13622 (N_13622,N_11150,N_10870);
nor U13623 (N_13623,N_11904,N_11786);
nand U13624 (N_13624,N_11654,N_9729);
nand U13625 (N_13625,N_10520,N_11754);
and U13626 (N_13626,N_10483,N_11119);
and U13627 (N_13627,N_11048,N_10880);
or U13628 (N_13628,N_10516,N_9174);
or U13629 (N_13629,N_10853,N_10966);
and U13630 (N_13630,N_9091,N_10597);
nor U13631 (N_13631,N_9304,N_9110);
and U13632 (N_13632,N_9459,N_11932);
and U13633 (N_13633,N_9581,N_9102);
nand U13634 (N_13634,N_11087,N_11198);
and U13635 (N_13635,N_10521,N_10240);
nand U13636 (N_13636,N_10589,N_11882);
or U13637 (N_13637,N_11958,N_11052);
and U13638 (N_13638,N_9970,N_9433);
or U13639 (N_13639,N_11529,N_11019);
nand U13640 (N_13640,N_10423,N_11051);
or U13641 (N_13641,N_11563,N_9021);
or U13642 (N_13642,N_9252,N_11236);
or U13643 (N_13643,N_9062,N_11837);
and U13644 (N_13644,N_11215,N_9803);
nand U13645 (N_13645,N_11610,N_11511);
nand U13646 (N_13646,N_9222,N_10941);
and U13647 (N_13647,N_11211,N_9067);
or U13648 (N_13648,N_10600,N_9574);
and U13649 (N_13649,N_9643,N_9593);
nor U13650 (N_13650,N_9545,N_9243);
nor U13651 (N_13651,N_11786,N_11157);
or U13652 (N_13652,N_10806,N_9020);
nor U13653 (N_13653,N_9208,N_10361);
and U13654 (N_13654,N_9705,N_10202);
nand U13655 (N_13655,N_9499,N_9596);
nand U13656 (N_13656,N_9471,N_11895);
or U13657 (N_13657,N_10521,N_11493);
or U13658 (N_13658,N_10274,N_9526);
nand U13659 (N_13659,N_10049,N_11887);
nand U13660 (N_13660,N_9154,N_10977);
nand U13661 (N_13661,N_10000,N_9019);
and U13662 (N_13662,N_11650,N_9399);
nor U13663 (N_13663,N_11165,N_9631);
and U13664 (N_13664,N_10724,N_9540);
or U13665 (N_13665,N_9021,N_10341);
nand U13666 (N_13666,N_9410,N_11831);
and U13667 (N_13667,N_10370,N_10344);
and U13668 (N_13668,N_10222,N_9795);
or U13669 (N_13669,N_10349,N_11400);
or U13670 (N_13670,N_9276,N_10109);
nor U13671 (N_13671,N_9217,N_11601);
nand U13672 (N_13672,N_11179,N_9736);
or U13673 (N_13673,N_9125,N_10861);
and U13674 (N_13674,N_10064,N_10833);
nor U13675 (N_13675,N_9779,N_10583);
nand U13676 (N_13676,N_9720,N_11301);
nor U13677 (N_13677,N_10996,N_11341);
or U13678 (N_13678,N_9773,N_10515);
nand U13679 (N_13679,N_11112,N_10360);
nand U13680 (N_13680,N_11209,N_10735);
or U13681 (N_13681,N_9505,N_9551);
nor U13682 (N_13682,N_9166,N_9654);
nand U13683 (N_13683,N_9800,N_11630);
nor U13684 (N_13684,N_9892,N_10521);
nor U13685 (N_13685,N_11206,N_10435);
nand U13686 (N_13686,N_9583,N_9681);
and U13687 (N_13687,N_10824,N_9824);
and U13688 (N_13688,N_10268,N_9520);
nand U13689 (N_13689,N_10066,N_10969);
nand U13690 (N_13690,N_9987,N_9467);
or U13691 (N_13691,N_10752,N_9146);
nor U13692 (N_13692,N_9335,N_9418);
nor U13693 (N_13693,N_9639,N_10824);
or U13694 (N_13694,N_10667,N_9608);
nand U13695 (N_13695,N_11446,N_9763);
and U13696 (N_13696,N_9089,N_10535);
and U13697 (N_13697,N_9086,N_9353);
or U13698 (N_13698,N_9245,N_11416);
nor U13699 (N_13699,N_10512,N_11075);
or U13700 (N_13700,N_10048,N_9937);
nor U13701 (N_13701,N_9281,N_9041);
nor U13702 (N_13702,N_10815,N_10973);
nor U13703 (N_13703,N_11391,N_11430);
and U13704 (N_13704,N_11976,N_11536);
or U13705 (N_13705,N_9927,N_11542);
nor U13706 (N_13706,N_9162,N_11359);
nor U13707 (N_13707,N_9436,N_10313);
nor U13708 (N_13708,N_9189,N_10286);
or U13709 (N_13709,N_9697,N_10376);
or U13710 (N_13710,N_9404,N_10991);
or U13711 (N_13711,N_9889,N_9817);
xnor U13712 (N_13712,N_11206,N_11759);
nor U13713 (N_13713,N_11787,N_9077);
and U13714 (N_13714,N_11757,N_9631);
nor U13715 (N_13715,N_9378,N_10706);
and U13716 (N_13716,N_10666,N_9056);
nor U13717 (N_13717,N_11921,N_10488);
nor U13718 (N_13718,N_9808,N_9748);
nor U13719 (N_13719,N_10617,N_9572);
and U13720 (N_13720,N_9730,N_9595);
nand U13721 (N_13721,N_10934,N_9968);
nand U13722 (N_13722,N_11003,N_10065);
or U13723 (N_13723,N_9918,N_9270);
nand U13724 (N_13724,N_10687,N_9190);
nor U13725 (N_13725,N_10601,N_11624);
or U13726 (N_13726,N_10929,N_10687);
and U13727 (N_13727,N_11213,N_10855);
nand U13728 (N_13728,N_10159,N_11859);
and U13729 (N_13729,N_11954,N_10244);
nor U13730 (N_13730,N_9564,N_11489);
and U13731 (N_13731,N_10876,N_9180);
and U13732 (N_13732,N_11686,N_11832);
nor U13733 (N_13733,N_11599,N_10058);
or U13734 (N_13734,N_9559,N_9594);
and U13735 (N_13735,N_11262,N_9651);
nor U13736 (N_13736,N_9882,N_10264);
nor U13737 (N_13737,N_10026,N_10765);
nor U13738 (N_13738,N_9471,N_9468);
and U13739 (N_13739,N_11981,N_10119);
and U13740 (N_13740,N_9949,N_11149);
nand U13741 (N_13741,N_9619,N_11282);
nand U13742 (N_13742,N_9505,N_9167);
and U13743 (N_13743,N_11526,N_10509);
or U13744 (N_13744,N_9996,N_10389);
nand U13745 (N_13745,N_9634,N_11037);
or U13746 (N_13746,N_9882,N_11188);
nand U13747 (N_13747,N_11671,N_11509);
or U13748 (N_13748,N_9891,N_11657);
nand U13749 (N_13749,N_10427,N_11425);
nand U13750 (N_13750,N_10671,N_10689);
or U13751 (N_13751,N_9388,N_10871);
and U13752 (N_13752,N_9863,N_9181);
nor U13753 (N_13753,N_9381,N_9451);
nor U13754 (N_13754,N_9325,N_9021);
nand U13755 (N_13755,N_9662,N_9440);
nor U13756 (N_13756,N_10750,N_9919);
or U13757 (N_13757,N_11223,N_11629);
nand U13758 (N_13758,N_9872,N_9343);
nand U13759 (N_13759,N_9753,N_10352);
and U13760 (N_13760,N_9004,N_11311);
nor U13761 (N_13761,N_9549,N_10457);
nand U13762 (N_13762,N_10384,N_10606);
nand U13763 (N_13763,N_10415,N_11206);
or U13764 (N_13764,N_10694,N_9843);
and U13765 (N_13765,N_9237,N_10069);
nor U13766 (N_13766,N_11016,N_9414);
nand U13767 (N_13767,N_9413,N_11199);
nand U13768 (N_13768,N_10258,N_11537);
nor U13769 (N_13769,N_9010,N_10789);
and U13770 (N_13770,N_10308,N_11843);
nand U13771 (N_13771,N_9615,N_9278);
nor U13772 (N_13772,N_10073,N_10102);
or U13773 (N_13773,N_10877,N_11975);
and U13774 (N_13774,N_9323,N_11711);
nor U13775 (N_13775,N_9538,N_9448);
nand U13776 (N_13776,N_9817,N_10473);
nand U13777 (N_13777,N_11285,N_9727);
and U13778 (N_13778,N_9810,N_10139);
or U13779 (N_13779,N_9899,N_11128);
or U13780 (N_13780,N_10652,N_11723);
nor U13781 (N_13781,N_11491,N_11777);
nor U13782 (N_13782,N_10287,N_10357);
xor U13783 (N_13783,N_11049,N_11693);
or U13784 (N_13784,N_9991,N_9518);
nor U13785 (N_13785,N_11764,N_10854);
nand U13786 (N_13786,N_9470,N_10545);
nor U13787 (N_13787,N_9252,N_9304);
nor U13788 (N_13788,N_10052,N_10042);
and U13789 (N_13789,N_10905,N_11819);
nor U13790 (N_13790,N_10453,N_10011);
nand U13791 (N_13791,N_10060,N_9499);
nor U13792 (N_13792,N_9382,N_10205);
and U13793 (N_13793,N_10613,N_10985);
nand U13794 (N_13794,N_11222,N_9982);
and U13795 (N_13795,N_11936,N_10223);
and U13796 (N_13796,N_9103,N_10986);
or U13797 (N_13797,N_10440,N_9015);
nand U13798 (N_13798,N_11499,N_9060);
and U13799 (N_13799,N_10161,N_10677);
nand U13800 (N_13800,N_11253,N_10955);
and U13801 (N_13801,N_11342,N_10312);
and U13802 (N_13802,N_9570,N_10825);
nand U13803 (N_13803,N_9173,N_11461);
and U13804 (N_13804,N_10387,N_10411);
and U13805 (N_13805,N_9522,N_11889);
nand U13806 (N_13806,N_10685,N_11126);
or U13807 (N_13807,N_11366,N_10111);
nand U13808 (N_13808,N_10675,N_10935);
and U13809 (N_13809,N_9107,N_11337);
nor U13810 (N_13810,N_9331,N_11623);
nor U13811 (N_13811,N_11080,N_10423);
nand U13812 (N_13812,N_9323,N_10887);
and U13813 (N_13813,N_10268,N_11287);
nor U13814 (N_13814,N_11592,N_11571);
or U13815 (N_13815,N_11905,N_11870);
nand U13816 (N_13816,N_11836,N_10358);
nor U13817 (N_13817,N_10074,N_11927);
nand U13818 (N_13818,N_11960,N_11986);
nand U13819 (N_13819,N_11808,N_9143);
or U13820 (N_13820,N_10736,N_11246);
nand U13821 (N_13821,N_11934,N_10413);
nor U13822 (N_13822,N_10003,N_11795);
nor U13823 (N_13823,N_11941,N_10507);
nor U13824 (N_13824,N_11553,N_10168);
and U13825 (N_13825,N_10330,N_11700);
or U13826 (N_13826,N_9609,N_10997);
nand U13827 (N_13827,N_10682,N_11205);
and U13828 (N_13828,N_9635,N_9731);
and U13829 (N_13829,N_10900,N_10070);
and U13830 (N_13830,N_10998,N_11855);
nor U13831 (N_13831,N_11090,N_9093);
nor U13832 (N_13832,N_9821,N_10428);
or U13833 (N_13833,N_11046,N_10548);
nor U13834 (N_13834,N_9777,N_11080);
nand U13835 (N_13835,N_11448,N_9549);
or U13836 (N_13836,N_10912,N_11472);
nor U13837 (N_13837,N_9747,N_11708);
nand U13838 (N_13838,N_11368,N_11545);
nand U13839 (N_13839,N_9109,N_10514);
and U13840 (N_13840,N_10251,N_9550);
nand U13841 (N_13841,N_10151,N_9724);
nand U13842 (N_13842,N_11733,N_10914);
nor U13843 (N_13843,N_11218,N_10894);
nor U13844 (N_13844,N_10534,N_9786);
and U13845 (N_13845,N_10437,N_9209);
nor U13846 (N_13846,N_9710,N_10459);
nand U13847 (N_13847,N_11609,N_11641);
nor U13848 (N_13848,N_10936,N_11846);
and U13849 (N_13849,N_11081,N_10273);
nand U13850 (N_13850,N_10381,N_10652);
or U13851 (N_13851,N_11969,N_9566);
nor U13852 (N_13852,N_9314,N_11050);
and U13853 (N_13853,N_11967,N_11766);
nor U13854 (N_13854,N_10898,N_9414);
nor U13855 (N_13855,N_9329,N_11824);
nand U13856 (N_13856,N_9245,N_9939);
or U13857 (N_13857,N_9335,N_9206);
nand U13858 (N_13858,N_11969,N_9564);
nand U13859 (N_13859,N_9655,N_10055);
and U13860 (N_13860,N_9002,N_9483);
nand U13861 (N_13861,N_11013,N_11175);
and U13862 (N_13862,N_9596,N_9794);
or U13863 (N_13863,N_10331,N_10604);
nand U13864 (N_13864,N_10501,N_10156);
or U13865 (N_13865,N_9553,N_11883);
nand U13866 (N_13866,N_9453,N_10751);
nor U13867 (N_13867,N_9825,N_10518);
nand U13868 (N_13868,N_11736,N_10802);
or U13869 (N_13869,N_11056,N_11063);
nand U13870 (N_13870,N_10560,N_10590);
or U13871 (N_13871,N_10674,N_11386);
nor U13872 (N_13872,N_10863,N_10511);
and U13873 (N_13873,N_9181,N_10937);
or U13874 (N_13874,N_11851,N_11540);
nor U13875 (N_13875,N_10563,N_10756);
or U13876 (N_13876,N_9032,N_10396);
nand U13877 (N_13877,N_11053,N_10869);
nand U13878 (N_13878,N_9869,N_9993);
nand U13879 (N_13879,N_10722,N_10670);
or U13880 (N_13880,N_9770,N_11407);
or U13881 (N_13881,N_11267,N_11804);
nor U13882 (N_13882,N_11707,N_11948);
or U13883 (N_13883,N_10321,N_10198);
nand U13884 (N_13884,N_11399,N_11172);
nand U13885 (N_13885,N_11054,N_11656);
or U13886 (N_13886,N_10632,N_9384);
nand U13887 (N_13887,N_10757,N_11490);
nand U13888 (N_13888,N_10558,N_9031);
or U13889 (N_13889,N_9270,N_9176);
or U13890 (N_13890,N_10590,N_10889);
nand U13891 (N_13891,N_11153,N_9207);
or U13892 (N_13892,N_11018,N_11570);
nor U13893 (N_13893,N_10424,N_10833);
nand U13894 (N_13894,N_9535,N_9193);
and U13895 (N_13895,N_9864,N_11167);
nand U13896 (N_13896,N_11282,N_10929);
nor U13897 (N_13897,N_10146,N_9176);
and U13898 (N_13898,N_10622,N_10749);
nor U13899 (N_13899,N_11488,N_11953);
or U13900 (N_13900,N_10220,N_9960);
and U13901 (N_13901,N_9045,N_9201);
and U13902 (N_13902,N_10629,N_10419);
and U13903 (N_13903,N_9098,N_10657);
or U13904 (N_13904,N_11627,N_9339);
nand U13905 (N_13905,N_11191,N_9703);
nand U13906 (N_13906,N_10610,N_9264);
nand U13907 (N_13907,N_10338,N_10255);
or U13908 (N_13908,N_10123,N_11432);
and U13909 (N_13909,N_11195,N_9820);
xor U13910 (N_13910,N_10521,N_10681);
nand U13911 (N_13911,N_9466,N_9884);
nand U13912 (N_13912,N_10628,N_11232);
nor U13913 (N_13913,N_10088,N_9136);
nand U13914 (N_13914,N_11603,N_10985);
nor U13915 (N_13915,N_10372,N_11374);
nand U13916 (N_13916,N_9024,N_11742);
and U13917 (N_13917,N_9481,N_11432);
nor U13918 (N_13918,N_10789,N_9265);
nor U13919 (N_13919,N_10405,N_10143);
or U13920 (N_13920,N_10538,N_10018);
or U13921 (N_13921,N_11752,N_9947);
nand U13922 (N_13922,N_11755,N_10482);
or U13923 (N_13923,N_11467,N_10166);
nand U13924 (N_13924,N_11412,N_9557);
and U13925 (N_13925,N_11101,N_9562);
nor U13926 (N_13926,N_10199,N_9679);
or U13927 (N_13927,N_9888,N_10825);
nand U13928 (N_13928,N_10046,N_11186);
and U13929 (N_13929,N_9483,N_11835);
or U13930 (N_13930,N_9417,N_10722);
nand U13931 (N_13931,N_11904,N_10091);
nor U13932 (N_13932,N_11696,N_10290);
nor U13933 (N_13933,N_9627,N_10772);
or U13934 (N_13934,N_11780,N_11610);
nand U13935 (N_13935,N_9955,N_10753);
and U13936 (N_13936,N_11764,N_10598);
nor U13937 (N_13937,N_11049,N_9208);
nor U13938 (N_13938,N_9515,N_11282);
and U13939 (N_13939,N_10148,N_11993);
and U13940 (N_13940,N_9330,N_11392);
nand U13941 (N_13941,N_10091,N_10060);
nand U13942 (N_13942,N_11870,N_11632);
or U13943 (N_13943,N_11654,N_10109);
nor U13944 (N_13944,N_9060,N_10082);
nor U13945 (N_13945,N_10367,N_11357);
or U13946 (N_13946,N_11435,N_11702);
and U13947 (N_13947,N_11366,N_11946);
nor U13948 (N_13948,N_9994,N_11605);
and U13949 (N_13949,N_9271,N_11843);
or U13950 (N_13950,N_11166,N_10898);
xor U13951 (N_13951,N_10344,N_9863);
or U13952 (N_13952,N_9558,N_9598);
or U13953 (N_13953,N_11179,N_9554);
nand U13954 (N_13954,N_9305,N_11060);
nand U13955 (N_13955,N_9576,N_11391);
nor U13956 (N_13956,N_11960,N_9500);
or U13957 (N_13957,N_10403,N_10361);
or U13958 (N_13958,N_10408,N_9948);
xor U13959 (N_13959,N_10315,N_10279);
and U13960 (N_13960,N_11679,N_10794);
and U13961 (N_13961,N_9257,N_9185);
nor U13962 (N_13962,N_11487,N_11638);
nand U13963 (N_13963,N_10588,N_10447);
nor U13964 (N_13964,N_9844,N_10568);
nor U13965 (N_13965,N_11108,N_11537);
and U13966 (N_13966,N_10799,N_10092);
nand U13967 (N_13967,N_9092,N_11095);
nand U13968 (N_13968,N_11918,N_10516);
nand U13969 (N_13969,N_9540,N_10229);
nand U13970 (N_13970,N_9076,N_9309);
nor U13971 (N_13971,N_9700,N_10754);
nand U13972 (N_13972,N_10337,N_11411);
nor U13973 (N_13973,N_9304,N_10329);
and U13974 (N_13974,N_11375,N_11556);
and U13975 (N_13975,N_11604,N_10609);
nand U13976 (N_13976,N_9486,N_11909);
and U13977 (N_13977,N_9029,N_10750);
xnor U13978 (N_13978,N_10163,N_9857);
and U13979 (N_13979,N_11856,N_9264);
or U13980 (N_13980,N_9507,N_10478);
or U13981 (N_13981,N_10975,N_9042);
or U13982 (N_13982,N_10446,N_9516);
nor U13983 (N_13983,N_9472,N_9028);
or U13984 (N_13984,N_9657,N_11070);
nand U13985 (N_13985,N_9078,N_10822);
nor U13986 (N_13986,N_11220,N_10965);
and U13987 (N_13987,N_10871,N_10150);
or U13988 (N_13988,N_11872,N_9650);
nor U13989 (N_13989,N_10741,N_9832);
nand U13990 (N_13990,N_9462,N_10326);
nor U13991 (N_13991,N_10037,N_9903);
and U13992 (N_13992,N_10721,N_11149);
nor U13993 (N_13993,N_9239,N_9947);
or U13994 (N_13994,N_9856,N_10242);
or U13995 (N_13995,N_10850,N_11128);
nand U13996 (N_13996,N_10359,N_11515);
and U13997 (N_13997,N_9833,N_10008);
nand U13998 (N_13998,N_11502,N_11172);
and U13999 (N_13999,N_11725,N_11907);
and U14000 (N_14000,N_9596,N_9273);
nor U14001 (N_14001,N_10918,N_10014);
or U14002 (N_14002,N_11333,N_10106);
nor U14003 (N_14003,N_10544,N_11334);
and U14004 (N_14004,N_10937,N_10354);
or U14005 (N_14005,N_9280,N_11451);
and U14006 (N_14006,N_9933,N_9642);
and U14007 (N_14007,N_9563,N_10844);
nor U14008 (N_14008,N_9878,N_9684);
or U14009 (N_14009,N_11853,N_11642);
or U14010 (N_14010,N_10144,N_9258);
and U14011 (N_14011,N_11020,N_9276);
nand U14012 (N_14012,N_9457,N_10025);
or U14013 (N_14013,N_9608,N_10315);
xnor U14014 (N_14014,N_9221,N_11582);
or U14015 (N_14015,N_9926,N_9226);
nor U14016 (N_14016,N_10555,N_10208);
and U14017 (N_14017,N_9825,N_9635);
or U14018 (N_14018,N_11373,N_9811);
or U14019 (N_14019,N_10564,N_9476);
nand U14020 (N_14020,N_9729,N_11741);
or U14021 (N_14021,N_10886,N_11044);
or U14022 (N_14022,N_10276,N_9635);
nand U14023 (N_14023,N_10599,N_11935);
or U14024 (N_14024,N_9276,N_9404);
nand U14025 (N_14025,N_10969,N_10177);
nor U14026 (N_14026,N_10929,N_9094);
nand U14027 (N_14027,N_11359,N_9799);
nor U14028 (N_14028,N_9301,N_9994);
or U14029 (N_14029,N_11755,N_9446);
nand U14030 (N_14030,N_9398,N_10850);
or U14031 (N_14031,N_10466,N_10913);
nor U14032 (N_14032,N_10372,N_9233);
or U14033 (N_14033,N_11605,N_10261);
and U14034 (N_14034,N_9548,N_9581);
nor U14035 (N_14035,N_10965,N_9428);
and U14036 (N_14036,N_9681,N_9252);
and U14037 (N_14037,N_11221,N_10062);
nor U14038 (N_14038,N_11056,N_9852);
and U14039 (N_14039,N_11758,N_9095);
nand U14040 (N_14040,N_9381,N_9700);
nor U14041 (N_14041,N_10552,N_10596);
nor U14042 (N_14042,N_9094,N_9921);
nor U14043 (N_14043,N_10192,N_11015);
nor U14044 (N_14044,N_11148,N_10723);
and U14045 (N_14045,N_9689,N_9290);
nand U14046 (N_14046,N_10332,N_11881);
nor U14047 (N_14047,N_10259,N_11825);
or U14048 (N_14048,N_10983,N_9463);
nor U14049 (N_14049,N_11044,N_10688);
and U14050 (N_14050,N_9749,N_10322);
and U14051 (N_14051,N_10129,N_10219);
nand U14052 (N_14052,N_9261,N_10196);
nand U14053 (N_14053,N_11884,N_9648);
nand U14054 (N_14054,N_11637,N_10202);
nand U14055 (N_14055,N_9857,N_9620);
or U14056 (N_14056,N_10031,N_11740);
and U14057 (N_14057,N_11819,N_11740);
or U14058 (N_14058,N_9712,N_10651);
nor U14059 (N_14059,N_11598,N_10600);
nand U14060 (N_14060,N_11001,N_9205);
nand U14061 (N_14061,N_11128,N_9303);
or U14062 (N_14062,N_9194,N_10424);
nand U14063 (N_14063,N_11956,N_9675);
nor U14064 (N_14064,N_10797,N_10064);
and U14065 (N_14065,N_9081,N_10184);
nor U14066 (N_14066,N_9264,N_9869);
nor U14067 (N_14067,N_10767,N_9578);
nor U14068 (N_14068,N_9028,N_9279);
nand U14069 (N_14069,N_10125,N_11177);
nand U14070 (N_14070,N_10652,N_11349);
or U14071 (N_14071,N_9925,N_9283);
nor U14072 (N_14072,N_10878,N_11755);
nor U14073 (N_14073,N_10002,N_11100);
and U14074 (N_14074,N_9477,N_11889);
nand U14075 (N_14075,N_10813,N_11287);
nor U14076 (N_14076,N_10833,N_10380);
nand U14077 (N_14077,N_9495,N_9804);
or U14078 (N_14078,N_11633,N_10501);
nand U14079 (N_14079,N_9391,N_10370);
and U14080 (N_14080,N_9843,N_10311);
nor U14081 (N_14081,N_11357,N_9771);
nor U14082 (N_14082,N_10966,N_9329);
nand U14083 (N_14083,N_9843,N_9375);
and U14084 (N_14084,N_9615,N_9329);
and U14085 (N_14085,N_9417,N_9853);
or U14086 (N_14086,N_9451,N_11563);
and U14087 (N_14087,N_11312,N_9201);
and U14088 (N_14088,N_10259,N_9216);
nand U14089 (N_14089,N_11541,N_10291);
and U14090 (N_14090,N_10157,N_11384);
nand U14091 (N_14091,N_11103,N_10677);
and U14092 (N_14092,N_11366,N_9923);
or U14093 (N_14093,N_9923,N_11418);
nand U14094 (N_14094,N_9534,N_9999);
and U14095 (N_14095,N_10871,N_11865);
nor U14096 (N_14096,N_9871,N_9451);
nor U14097 (N_14097,N_10749,N_9062);
nor U14098 (N_14098,N_11316,N_9554);
and U14099 (N_14099,N_10384,N_11342);
nor U14100 (N_14100,N_11810,N_9835);
nor U14101 (N_14101,N_9521,N_10039);
nand U14102 (N_14102,N_11987,N_10565);
nor U14103 (N_14103,N_11364,N_11656);
and U14104 (N_14104,N_9411,N_11405);
or U14105 (N_14105,N_9797,N_9377);
and U14106 (N_14106,N_11753,N_10469);
and U14107 (N_14107,N_11386,N_9435);
or U14108 (N_14108,N_11908,N_10183);
nand U14109 (N_14109,N_11313,N_9436);
or U14110 (N_14110,N_9310,N_11615);
nand U14111 (N_14111,N_10584,N_10728);
nand U14112 (N_14112,N_11452,N_9227);
nor U14113 (N_14113,N_10457,N_10590);
and U14114 (N_14114,N_10921,N_9618);
nand U14115 (N_14115,N_9531,N_9864);
nand U14116 (N_14116,N_11777,N_11246);
nor U14117 (N_14117,N_11714,N_11817);
or U14118 (N_14118,N_9736,N_11525);
nor U14119 (N_14119,N_9230,N_9970);
nor U14120 (N_14120,N_9534,N_9936);
nand U14121 (N_14121,N_9914,N_11825);
and U14122 (N_14122,N_10515,N_11506);
and U14123 (N_14123,N_10912,N_9330);
and U14124 (N_14124,N_9986,N_11253);
nand U14125 (N_14125,N_10504,N_10239);
or U14126 (N_14126,N_11767,N_10040);
or U14127 (N_14127,N_10914,N_11203);
and U14128 (N_14128,N_11875,N_9130);
and U14129 (N_14129,N_9605,N_10974);
or U14130 (N_14130,N_11059,N_9966);
or U14131 (N_14131,N_9983,N_10681);
or U14132 (N_14132,N_10241,N_9886);
nand U14133 (N_14133,N_11485,N_11909);
or U14134 (N_14134,N_9114,N_9044);
and U14135 (N_14135,N_9964,N_11235);
or U14136 (N_14136,N_9405,N_11692);
or U14137 (N_14137,N_9164,N_10194);
or U14138 (N_14138,N_9425,N_11875);
or U14139 (N_14139,N_10819,N_9374);
nor U14140 (N_14140,N_11048,N_10554);
nand U14141 (N_14141,N_10596,N_10819);
nand U14142 (N_14142,N_9865,N_11754);
or U14143 (N_14143,N_11852,N_10823);
nor U14144 (N_14144,N_11475,N_10108);
nor U14145 (N_14145,N_9937,N_9773);
nand U14146 (N_14146,N_10627,N_10861);
nor U14147 (N_14147,N_9693,N_10600);
nand U14148 (N_14148,N_9584,N_10778);
nor U14149 (N_14149,N_10820,N_11261);
nand U14150 (N_14150,N_11170,N_9144);
nor U14151 (N_14151,N_11104,N_10983);
nand U14152 (N_14152,N_10148,N_11554);
nand U14153 (N_14153,N_11889,N_10034);
and U14154 (N_14154,N_11534,N_11284);
nand U14155 (N_14155,N_11060,N_11388);
or U14156 (N_14156,N_9646,N_10862);
and U14157 (N_14157,N_10477,N_11680);
and U14158 (N_14158,N_9801,N_11126);
and U14159 (N_14159,N_9590,N_9910);
nand U14160 (N_14160,N_11313,N_10435);
and U14161 (N_14161,N_11775,N_9686);
nor U14162 (N_14162,N_9373,N_10427);
and U14163 (N_14163,N_10654,N_10922);
nor U14164 (N_14164,N_10447,N_11668);
and U14165 (N_14165,N_9688,N_9695);
nor U14166 (N_14166,N_9602,N_11505);
or U14167 (N_14167,N_10908,N_9050);
nor U14168 (N_14168,N_10745,N_11653);
nand U14169 (N_14169,N_9820,N_11708);
nand U14170 (N_14170,N_10262,N_11765);
and U14171 (N_14171,N_9172,N_9906);
nor U14172 (N_14172,N_11009,N_10059);
nor U14173 (N_14173,N_11597,N_11769);
and U14174 (N_14174,N_10869,N_11610);
nand U14175 (N_14175,N_9546,N_11517);
nand U14176 (N_14176,N_11108,N_11279);
nand U14177 (N_14177,N_11208,N_11773);
nor U14178 (N_14178,N_9683,N_10848);
nand U14179 (N_14179,N_9042,N_9678);
and U14180 (N_14180,N_9415,N_9853);
and U14181 (N_14181,N_9009,N_10616);
nor U14182 (N_14182,N_10274,N_10451);
nor U14183 (N_14183,N_10773,N_11570);
nand U14184 (N_14184,N_11531,N_9956);
nor U14185 (N_14185,N_9327,N_9701);
or U14186 (N_14186,N_9170,N_10065);
or U14187 (N_14187,N_10350,N_11045);
nor U14188 (N_14188,N_9437,N_10632);
nand U14189 (N_14189,N_10645,N_10606);
or U14190 (N_14190,N_10159,N_10315);
nand U14191 (N_14191,N_9481,N_9058);
or U14192 (N_14192,N_9039,N_9834);
or U14193 (N_14193,N_10597,N_9964);
and U14194 (N_14194,N_10924,N_10801);
and U14195 (N_14195,N_11821,N_10064);
or U14196 (N_14196,N_11707,N_9670);
nor U14197 (N_14197,N_9305,N_10917);
nor U14198 (N_14198,N_9626,N_11784);
nand U14199 (N_14199,N_10073,N_10025);
nand U14200 (N_14200,N_10704,N_9597);
and U14201 (N_14201,N_9535,N_9378);
nand U14202 (N_14202,N_10862,N_10150);
and U14203 (N_14203,N_11904,N_11142);
nand U14204 (N_14204,N_9312,N_11327);
nand U14205 (N_14205,N_10142,N_10388);
and U14206 (N_14206,N_11811,N_11796);
and U14207 (N_14207,N_11561,N_9891);
nor U14208 (N_14208,N_11489,N_11135);
nor U14209 (N_14209,N_10128,N_9818);
nand U14210 (N_14210,N_9843,N_9778);
and U14211 (N_14211,N_10640,N_10057);
and U14212 (N_14212,N_9872,N_10915);
and U14213 (N_14213,N_9938,N_11553);
and U14214 (N_14214,N_10872,N_11921);
and U14215 (N_14215,N_9285,N_11441);
and U14216 (N_14216,N_9421,N_11228);
nand U14217 (N_14217,N_11410,N_11582);
and U14218 (N_14218,N_11934,N_9857);
nand U14219 (N_14219,N_9990,N_10466);
or U14220 (N_14220,N_11789,N_10420);
nand U14221 (N_14221,N_11692,N_10142);
or U14222 (N_14222,N_9499,N_10466);
and U14223 (N_14223,N_10383,N_10858);
and U14224 (N_14224,N_9201,N_9346);
nand U14225 (N_14225,N_10953,N_11213);
and U14226 (N_14226,N_9959,N_9729);
and U14227 (N_14227,N_9561,N_11912);
nor U14228 (N_14228,N_10673,N_11651);
nor U14229 (N_14229,N_9095,N_9832);
and U14230 (N_14230,N_11237,N_11145);
or U14231 (N_14231,N_11131,N_11251);
and U14232 (N_14232,N_10677,N_11916);
nor U14233 (N_14233,N_9791,N_10664);
nor U14234 (N_14234,N_10467,N_9640);
nand U14235 (N_14235,N_11758,N_9539);
or U14236 (N_14236,N_10865,N_9404);
and U14237 (N_14237,N_9517,N_11665);
and U14238 (N_14238,N_9208,N_10457);
and U14239 (N_14239,N_11377,N_11404);
nor U14240 (N_14240,N_11490,N_10930);
or U14241 (N_14241,N_9564,N_10647);
nand U14242 (N_14242,N_11761,N_10696);
or U14243 (N_14243,N_11688,N_11078);
nor U14244 (N_14244,N_10976,N_10187);
nand U14245 (N_14245,N_10399,N_11157);
nand U14246 (N_14246,N_9458,N_10556);
nand U14247 (N_14247,N_11378,N_9277);
and U14248 (N_14248,N_10659,N_11665);
and U14249 (N_14249,N_10718,N_9323);
nand U14250 (N_14250,N_9052,N_11461);
nand U14251 (N_14251,N_9874,N_10006);
nand U14252 (N_14252,N_10461,N_10492);
nand U14253 (N_14253,N_11816,N_11178);
nand U14254 (N_14254,N_11840,N_10904);
nor U14255 (N_14255,N_9068,N_11077);
or U14256 (N_14256,N_9707,N_11427);
nor U14257 (N_14257,N_10498,N_11227);
and U14258 (N_14258,N_11661,N_10402);
nor U14259 (N_14259,N_10716,N_9113);
and U14260 (N_14260,N_10718,N_10493);
nor U14261 (N_14261,N_10431,N_11354);
nor U14262 (N_14262,N_10998,N_9326);
nor U14263 (N_14263,N_9658,N_9719);
nand U14264 (N_14264,N_9737,N_10980);
nand U14265 (N_14265,N_10116,N_11110);
nor U14266 (N_14266,N_9375,N_11054);
nand U14267 (N_14267,N_10480,N_9252);
nor U14268 (N_14268,N_11030,N_10832);
or U14269 (N_14269,N_11805,N_11097);
nand U14270 (N_14270,N_9112,N_9860);
nor U14271 (N_14271,N_9658,N_9173);
and U14272 (N_14272,N_10806,N_9316);
and U14273 (N_14273,N_9795,N_11901);
nor U14274 (N_14274,N_10098,N_10897);
nand U14275 (N_14275,N_10645,N_10852);
or U14276 (N_14276,N_11658,N_11891);
nand U14277 (N_14277,N_10747,N_10422);
and U14278 (N_14278,N_11251,N_11151);
and U14279 (N_14279,N_11433,N_9533);
nor U14280 (N_14280,N_10703,N_11229);
or U14281 (N_14281,N_10530,N_11316);
and U14282 (N_14282,N_9818,N_10440);
nand U14283 (N_14283,N_11810,N_10214);
or U14284 (N_14284,N_10515,N_10930);
and U14285 (N_14285,N_10171,N_9654);
nand U14286 (N_14286,N_11202,N_11440);
or U14287 (N_14287,N_11134,N_10395);
and U14288 (N_14288,N_9912,N_9498);
nand U14289 (N_14289,N_10750,N_9787);
or U14290 (N_14290,N_11089,N_11728);
and U14291 (N_14291,N_10790,N_11404);
or U14292 (N_14292,N_11169,N_9881);
or U14293 (N_14293,N_9899,N_9529);
and U14294 (N_14294,N_9618,N_10329);
or U14295 (N_14295,N_11274,N_10550);
nor U14296 (N_14296,N_9908,N_9794);
nand U14297 (N_14297,N_10204,N_10991);
nand U14298 (N_14298,N_11221,N_10224);
nand U14299 (N_14299,N_10310,N_11238);
nor U14300 (N_14300,N_9027,N_10109);
nand U14301 (N_14301,N_11969,N_10987);
and U14302 (N_14302,N_10511,N_10311);
or U14303 (N_14303,N_11905,N_9502);
or U14304 (N_14304,N_10768,N_11412);
nand U14305 (N_14305,N_9515,N_10091);
or U14306 (N_14306,N_11154,N_9351);
xnor U14307 (N_14307,N_10010,N_10496);
or U14308 (N_14308,N_10351,N_11268);
and U14309 (N_14309,N_10111,N_10315);
nand U14310 (N_14310,N_9837,N_10324);
xnor U14311 (N_14311,N_10530,N_11903);
nor U14312 (N_14312,N_9569,N_9771);
nand U14313 (N_14313,N_11997,N_11304);
nor U14314 (N_14314,N_10608,N_11446);
nand U14315 (N_14315,N_11932,N_11600);
or U14316 (N_14316,N_9108,N_11203);
nor U14317 (N_14317,N_10683,N_10247);
and U14318 (N_14318,N_10916,N_10210);
nor U14319 (N_14319,N_10692,N_10133);
and U14320 (N_14320,N_9760,N_9958);
or U14321 (N_14321,N_11264,N_10352);
nor U14322 (N_14322,N_9338,N_11304);
or U14323 (N_14323,N_11086,N_11778);
nor U14324 (N_14324,N_10463,N_11750);
and U14325 (N_14325,N_9341,N_11724);
nand U14326 (N_14326,N_9902,N_10705);
and U14327 (N_14327,N_11316,N_10312);
nand U14328 (N_14328,N_9910,N_9480);
nand U14329 (N_14329,N_11748,N_11804);
nor U14330 (N_14330,N_9164,N_11803);
and U14331 (N_14331,N_11829,N_9596);
or U14332 (N_14332,N_9583,N_10919);
nor U14333 (N_14333,N_10488,N_9991);
nor U14334 (N_14334,N_10304,N_11796);
and U14335 (N_14335,N_11813,N_10199);
or U14336 (N_14336,N_10262,N_9474);
nor U14337 (N_14337,N_11105,N_11087);
and U14338 (N_14338,N_9255,N_11399);
or U14339 (N_14339,N_10655,N_10283);
and U14340 (N_14340,N_9699,N_10488);
nor U14341 (N_14341,N_11433,N_9429);
nor U14342 (N_14342,N_11783,N_10106);
nand U14343 (N_14343,N_9267,N_9528);
nand U14344 (N_14344,N_10142,N_10364);
nor U14345 (N_14345,N_9045,N_11551);
nor U14346 (N_14346,N_10545,N_11255);
or U14347 (N_14347,N_9805,N_10481);
nor U14348 (N_14348,N_9106,N_9856);
and U14349 (N_14349,N_10924,N_11647);
or U14350 (N_14350,N_10980,N_9992);
and U14351 (N_14351,N_9976,N_9777);
or U14352 (N_14352,N_10399,N_9718);
and U14353 (N_14353,N_9957,N_11363);
or U14354 (N_14354,N_9220,N_10572);
and U14355 (N_14355,N_11931,N_11076);
nand U14356 (N_14356,N_9049,N_9415);
and U14357 (N_14357,N_11258,N_9450);
nand U14358 (N_14358,N_9721,N_11090);
and U14359 (N_14359,N_10478,N_10472);
nor U14360 (N_14360,N_11573,N_10981);
nor U14361 (N_14361,N_9157,N_9887);
nand U14362 (N_14362,N_10593,N_10533);
nor U14363 (N_14363,N_11765,N_9781);
nor U14364 (N_14364,N_11632,N_9160);
nor U14365 (N_14365,N_11906,N_11343);
or U14366 (N_14366,N_11994,N_11434);
and U14367 (N_14367,N_9874,N_9124);
nor U14368 (N_14368,N_10884,N_11045);
or U14369 (N_14369,N_9591,N_9213);
nor U14370 (N_14370,N_11872,N_9822);
nand U14371 (N_14371,N_11737,N_11905);
nand U14372 (N_14372,N_10394,N_9991);
or U14373 (N_14373,N_11809,N_11271);
nor U14374 (N_14374,N_11788,N_11745);
or U14375 (N_14375,N_10179,N_10970);
or U14376 (N_14376,N_11944,N_11765);
or U14377 (N_14377,N_9259,N_10290);
nand U14378 (N_14378,N_11460,N_9905);
or U14379 (N_14379,N_9845,N_9624);
and U14380 (N_14380,N_10154,N_11204);
and U14381 (N_14381,N_10332,N_10859);
or U14382 (N_14382,N_10832,N_11373);
and U14383 (N_14383,N_9752,N_9441);
nor U14384 (N_14384,N_11878,N_11457);
and U14385 (N_14385,N_10594,N_9598);
xnor U14386 (N_14386,N_11895,N_9028);
nor U14387 (N_14387,N_11520,N_10884);
nand U14388 (N_14388,N_9160,N_10595);
nand U14389 (N_14389,N_11303,N_11388);
nor U14390 (N_14390,N_10560,N_9871);
or U14391 (N_14391,N_10200,N_9215);
nor U14392 (N_14392,N_10558,N_9821);
and U14393 (N_14393,N_10538,N_11550);
nor U14394 (N_14394,N_10580,N_11364);
and U14395 (N_14395,N_11871,N_11923);
nor U14396 (N_14396,N_10190,N_9728);
nor U14397 (N_14397,N_11484,N_11637);
nor U14398 (N_14398,N_9114,N_10203);
and U14399 (N_14399,N_11851,N_10188);
or U14400 (N_14400,N_10554,N_10515);
and U14401 (N_14401,N_10145,N_10823);
nand U14402 (N_14402,N_9710,N_9119);
nor U14403 (N_14403,N_11168,N_10727);
or U14404 (N_14404,N_11290,N_11502);
and U14405 (N_14405,N_9425,N_10125);
nor U14406 (N_14406,N_10287,N_11313);
and U14407 (N_14407,N_9590,N_10239);
and U14408 (N_14408,N_10638,N_9038);
and U14409 (N_14409,N_9196,N_9878);
nor U14410 (N_14410,N_9374,N_9659);
nand U14411 (N_14411,N_9858,N_11594);
nor U14412 (N_14412,N_11607,N_10178);
nor U14413 (N_14413,N_9664,N_10547);
and U14414 (N_14414,N_10965,N_10655);
xor U14415 (N_14415,N_10047,N_10451);
and U14416 (N_14416,N_11217,N_11113);
and U14417 (N_14417,N_9424,N_9123);
nand U14418 (N_14418,N_11230,N_11809);
nor U14419 (N_14419,N_11661,N_9477);
and U14420 (N_14420,N_9505,N_9843);
nor U14421 (N_14421,N_11661,N_10723);
nor U14422 (N_14422,N_10684,N_11228);
or U14423 (N_14423,N_10339,N_11691);
nor U14424 (N_14424,N_9769,N_9400);
nand U14425 (N_14425,N_11299,N_11187);
or U14426 (N_14426,N_11950,N_11186);
and U14427 (N_14427,N_9794,N_10878);
xnor U14428 (N_14428,N_10183,N_11983);
and U14429 (N_14429,N_9183,N_11190);
or U14430 (N_14430,N_9624,N_9047);
nor U14431 (N_14431,N_10341,N_11360);
and U14432 (N_14432,N_11617,N_11715);
and U14433 (N_14433,N_11133,N_10772);
or U14434 (N_14434,N_10807,N_10813);
nor U14435 (N_14435,N_9273,N_9288);
nor U14436 (N_14436,N_10980,N_10476);
nand U14437 (N_14437,N_11068,N_10640);
and U14438 (N_14438,N_11220,N_9679);
or U14439 (N_14439,N_9977,N_10813);
and U14440 (N_14440,N_11443,N_9359);
nand U14441 (N_14441,N_10074,N_10462);
and U14442 (N_14442,N_9356,N_11231);
or U14443 (N_14443,N_10600,N_11838);
and U14444 (N_14444,N_10139,N_11109);
or U14445 (N_14445,N_10818,N_9163);
nor U14446 (N_14446,N_11773,N_10063);
and U14447 (N_14447,N_11633,N_9294);
and U14448 (N_14448,N_11252,N_10369);
and U14449 (N_14449,N_9248,N_9444);
and U14450 (N_14450,N_11304,N_10713);
or U14451 (N_14451,N_9381,N_10236);
nor U14452 (N_14452,N_10465,N_11614);
or U14453 (N_14453,N_10553,N_9922);
nor U14454 (N_14454,N_9684,N_9191);
nand U14455 (N_14455,N_10662,N_9854);
nor U14456 (N_14456,N_10312,N_9594);
or U14457 (N_14457,N_11325,N_10403);
and U14458 (N_14458,N_11468,N_11969);
nor U14459 (N_14459,N_11299,N_9125);
nand U14460 (N_14460,N_9363,N_10132);
nand U14461 (N_14461,N_11060,N_10251);
nand U14462 (N_14462,N_9167,N_10292);
and U14463 (N_14463,N_9177,N_11980);
and U14464 (N_14464,N_10397,N_10782);
or U14465 (N_14465,N_9848,N_10656);
nand U14466 (N_14466,N_11582,N_9176);
and U14467 (N_14467,N_11923,N_9082);
nand U14468 (N_14468,N_9178,N_11248);
xor U14469 (N_14469,N_11850,N_10083);
nor U14470 (N_14470,N_9881,N_10554);
nand U14471 (N_14471,N_10975,N_11474);
nand U14472 (N_14472,N_10677,N_11043);
nor U14473 (N_14473,N_10922,N_10338);
nor U14474 (N_14474,N_11659,N_9976);
and U14475 (N_14475,N_10428,N_10714);
or U14476 (N_14476,N_11605,N_10792);
and U14477 (N_14477,N_9799,N_9634);
and U14478 (N_14478,N_11786,N_11855);
and U14479 (N_14479,N_10429,N_9609);
or U14480 (N_14480,N_10668,N_9825);
nor U14481 (N_14481,N_9126,N_10310);
nor U14482 (N_14482,N_9696,N_10061);
nor U14483 (N_14483,N_11205,N_10628);
and U14484 (N_14484,N_10805,N_11806);
and U14485 (N_14485,N_11815,N_9841);
nor U14486 (N_14486,N_10359,N_9144);
and U14487 (N_14487,N_10683,N_11341);
nand U14488 (N_14488,N_9697,N_10842);
or U14489 (N_14489,N_9793,N_9239);
and U14490 (N_14490,N_9156,N_11524);
or U14491 (N_14491,N_9094,N_11431);
or U14492 (N_14492,N_10176,N_10127);
nand U14493 (N_14493,N_11535,N_9313);
or U14494 (N_14494,N_10126,N_10708);
nand U14495 (N_14495,N_9669,N_11762);
or U14496 (N_14496,N_10971,N_9269);
and U14497 (N_14497,N_10405,N_10584);
and U14498 (N_14498,N_9810,N_11220);
nor U14499 (N_14499,N_9698,N_9730);
nor U14500 (N_14500,N_9469,N_10007);
or U14501 (N_14501,N_9284,N_11110);
nor U14502 (N_14502,N_9285,N_11985);
and U14503 (N_14503,N_9897,N_11573);
and U14504 (N_14504,N_10404,N_11065);
or U14505 (N_14505,N_10206,N_10578);
nand U14506 (N_14506,N_11859,N_11259);
or U14507 (N_14507,N_11733,N_9540);
and U14508 (N_14508,N_11731,N_10122);
xor U14509 (N_14509,N_11679,N_11063);
nor U14510 (N_14510,N_10435,N_11590);
nor U14511 (N_14511,N_9508,N_11907);
nand U14512 (N_14512,N_9143,N_11026);
nand U14513 (N_14513,N_10170,N_11898);
or U14514 (N_14514,N_9557,N_11888);
nand U14515 (N_14515,N_10684,N_9008);
or U14516 (N_14516,N_9484,N_10851);
and U14517 (N_14517,N_11401,N_11754);
or U14518 (N_14518,N_10520,N_10688);
or U14519 (N_14519,N_10181,N_11553);
and U14520 (N_14520,N_10048,N_9677);
nand U14521 (N_14521,N_9843,N_10087);
nand U14522 (N_14522,N_11306,N_9729);
or U14523 (N_14523,N_10032,N_11327);
and U14524 (N_14524,N_9191,N_10798);
or U14525 (N_14525,N_9507,N_9762);
or U14526 (N_14526,N_9708,N_9431);
or U14527 (N_14527,N_9674,N_9482);
nor U14528 (N_14528,N_9708,N_11245);
nand U14529 (N_14529,N_9680,N_9784);
and U14530 (N_14530,N_11640,N_11133);
nand U14531 (N_14531,N_11931,N_10549);
and U14532 (N_14532,N_10970,N_9508);
or U14533 (N_14533,N_9347,N_11372);
nand U14534 (N_14534,N_11092,N_9223);
or U14535 (N_14535,N_9976,N_9216);
or U14536 (N_14536,N_9749,N_9048);
and U14537 (N_14537,N_11326,N_9617);
or U14538 (N_14538,N_9702,N_10336);
and U14539 (N_14539,N_11702,N_9617);
nand U14540 (N_14540,N_10732,N_9012);
xnor U14541 (N_14541,N_9602,N_11122);
or U14542 (N_14542,N_9033,N_10313);
nand U14543 (N_14543,N_11406,N_11336);
or U14544 (N_14544,N_9965,N_11125);
or U14545 (N_14545,N_9432,N_11286);
nor U14546 (N_14546,N_10687,N_9030);
and U14547 (N_14547,N_9088,N_9790);
nand U14548 (N_14548,N_9791,N_10556);
and U14549 (N_14549,N_11027,N_11792);
nor U14550 (N_14550,N_9902,N_10132);
nor U14551 (N_14551,N_9988,N_10308);
nor U14552 (N_14552,N_9536,N_9173);
nand U14553 (N_14553,N_10237,N_10142);
or U14554 (N_14554,N_9080,N_11370);
and U14555 (N_14555,N_9265,N_9670);
and U14556 (N_14556,N_9271,N_11355);
or U14557 (N_14557,N_10130,N_9577);
and U14558 (N_14558,N_10937,N_10393);
nand U14559 (N_14559,N_9118,N_11699);
and U14560 (N_14560,N_11051,N_11206);
nand U14561 (N_14561,N_11055,N_11901);
nand U14562 (N_14562,N_9994,N_11786);
and U14563 (N_14563,N_11371,N_11743);
nand U14564 (N_14564,N_10023,N_11468);
nor U14565 (N_14565,N_9215,N_10428);
and U14566 (N_14566,N_11125,N_11056);
and U14567 (N_14567,N_9424,N_10711);
nand U14568 (N_14568,N_10264,N_10853);
and U14569 (N_14569,N_10339,N_11819);
nor U14570 (N_14570,N_10977,N_10519);
and U14571 (N_14571,N_10090,N_9905);
nand U14572 (N_14572,N_11562,N_11116);
and U14573 (N_14573,N_10906,N_9641);
nand U14574 (N_14574,N_9469,N_11148);
and U14575 (N_14575,N_10523,N_11143);
or U14576 (N_14576,N_11506,N_10409);
and U14577 (N_14577,N_10545,N_11245);
nor U14578 (N_14578,N_10762,N_10780);
nand U14579 (N_14579,N_11432,N_11250);
or U14580 (N_14580,N_11607,N_10508);
or U14581 (N_14581,N_9976,N_11658);
or U14582 (N_14582,N_10746,N_9880);
and U14583 (N_14583,N_11679,N_11850);
and U14584 (N_14584,N_9065,N_10019);
nor U14585 (N_14585,N_10587,N_11675);
nor U14586 (N_14586,N_10877,N_9344);
or U14587 (N_14587,N_11848,N_9369);
nor U14588 (N_14588,N_11409,N_11049);
or U14589 (N_14589,N_11444,N_9987);
or U14590 (N_14590,N_11693,N_11295);
and U14591 (N_14591,N_11480,N_9267);
nor U14592 (N_14592,N_11769,N_9750);
nor U14593 (N_14593,N_9266,N_10010);
nor U14594 (N_14594,N_11074,N_9696);
and U14595 (N_14595,N_9989,N_11776);
or U14596 (N_14596,N_11495,N_9062);
nor U14597 (N_14597,N_9994,N_10210);
or U14598 (N_14598,N_9933,N_11081);
and U14599 (N_14599,N_11226,N_9326);
and U14600 (N_14600,N_9509,N_10385);
or U14601 (N_14601,N_10031,N_11607);
nor U14602 (N_14602,N_9766,N_10861);
or U14603 (N_14603,N_9128,N_10001);
or U14604 (N_14604,N_9872,N_10168);
or U14605 (N_14605,N_10547,N_11288);
or U14606 (N_14606,N_11561,N_11218);
nor U14607 (N_14607,N_10504,N_11105);
or U14608 (N_14608,N_10439,N_11125);
nor U14609 (N_14609,N_10853,N_9486);
nand U14610 (N_14610,N_9671,N_11757);
nand U14611 (N_14611,N_9092,N_9206);
nand U14612 (N_14612,N_9460,N_11105);
or U14613 (N_14613,N_10970,N_10945);
nand U14614 (N_14614,N_9030,N_9273);
nand U14615 (N_14615,N_10697,N_10971);
nor U14616 (N_14616,N_11497,N_9199);
or U14617 (N_14617,N_10760,N_9295);
and U14618 (N_14618,N_9195,N_10550);
and U14619 (N_14619,N_11737,N_9324);
and U14620 (N_14620,N_11583,N_11249);
and U14621 (N_14621,N_9765,N_11333);
and U14622 (N_14622,N_11295,N_10438);
nand U14623 (N_14623,N_11424,N_9138);
nor U14624 (N_14624,N_9681,N_9708);
or U14625 (N_14625,N_11560,N_9408);
or U14626 (N_14626,N_9412,N_11625);
nor U14627 (N_14627,N_10272,N_11368);
or U14628 (N_14628,N_11234,N_10873);
and U14629 (N_14629,N_11648,N_11544);
nand U14630 (N_14630,N_10184,N_10300);
nor U14631 (N_14631,N_11314,N_10583);
nor U14632 (N_14632,N_10349,N_11141);
nand U14633 (N_14633,N_9326,N_10211);
nand U14634 (N_14634,N_10754,N_11027);
and U14635 (N_14635,N_11599,N_9499);
or U14636 (N_14636,N_9315,N_10468);
or U14637 (N_14637,N_10143,N_11021);
or U14638 (N_14638,N_11925,N_9575);
nor U14639 (N_14639,N_11035,N_10854);
nor U14640 (N_14640,N_10433,N_11215);
nand U14641 (N_14641,N_10809,N_10222);
nand U14642 (N_14642,N_9662,N_11559);
nand U14643 (N_14643,N_11900,N_9288);
or U14644 (N_14644,N_11518,N_9174);
or U14645 (N_14645,N_10765,N_9251);
or U14646 (N_14646,N_11942,N_10542);
nor U14647 (N_14647,N_10467,N_9745);
nand U14648 (N_14648,N_10560,N_10669);
nor U14649 (N_14649,N_11772,N_11738);
nor U14650 (N_14650,N_10421,N_11671);
and U14651 (N_14651,N_10516,N_11204);
or U14652 (N_14652,N_11841,N_9304);
nand U14653 (N_14653,N_11037,N_10174);
and U14654 (N_14654,N_11973,N_10611);
nand U14655 (N_14655,N_11955,N_11361);
or U14656 (N_14656,N_10112,N_9440);
and U14657 (N_14657,N_10486,N_9144);
nor U14658 (N_14658,N_9026,N_10148);
nand U14659 (N_14659,N_9699,N_11208);
nand U14660 (N_14660,N_10735,N_11139);
and U14661 (N_14661,N_10775,N_9996);
or U14662 (N_14662,N_11299,N_10211);
nand U14663 (N_14663,N_9880,N_10339);
nand U14664 (N_14664,N_10506,N_10192);
nand U14665 (N_14665,N_11356,N_9240);
or U14666 (N_14666,N_9759,N_11640);
nand U14667 (N_14667,N_9710,N_9232);
or U14668 (N_14668,N_10981,N_11865);
or U14669 (N_14669,N_9318,N_11048);
or U14670 (N_14670,N_9602,N_10895);
nand U14671 (N_14671,N_10995,N_11866);
or U14672 (N_14672,N_9898,N_10157);
nand U14673 (N_14673,N_10761,N_11680);
nor U14674 (N_14674,N_11975,N_9635);
or U14675 (N_14675,N_10396,N_9192);
and U14676 (N_14676,N_9689,N_10443);
or U14677 (N_14677,N_11159,N_9872);
nor U14678 (N_14678,N_9005,N_9148);
nor U14679 (N_14679,N_10720,N_10281);
or U14680 (N_14680,N_9913,N_10558);
or U14681 (N_14681,N_11220,N_9615);
and U14682 (N_14682,N_10079,N_11867);
nand U14683 (N_14683,N_11945,N_9800);
or U14684 (N_14684,N_9033,N_9590);
or U14685 (N_14685,N_11794,N_10057);
nor U14686 (N_14686,N_11886,N_10072);
and U14687 (N_14687,N_9910,N_10790);
nand U14688 (N_14688,N_11173,N_11244);
nor U14689 (N_14689,N_9821,N_10653);
nor U14690 (N_14690,N_9647,N_11094);
nand U14691 (N_14691,N_11807,N_9834);
nand U14692 (N_14692,N_11202,N_11717);
nand U14693 (N_14693,N_10914,N_9616);
nand U14694 (N_14694,N_10066,N_11269);
nor U14695 (N_14695,N_9846,N_11370);
or U14696 (N_14696,N_9929,N_9115);
nand U14697 (N_14697,N_10707,N_10500);
and U14698 (N_14698,N_9805,N_10732);
nor U14699 (N_14699,N_10266,N_10350);
nor U14700 (N_14700,N_10197,N_9665);
or U14701 (N_14701,N_9014,N_9199);
nor U14702 (N_14702,N_9095,N_11281);
nand U14703 (N_14703,N_11057,N_9560);
xor U14704 (N_14704,N_9248,N_10693);
nand U14705 (N_14705,N_11139,N_11161);
nand U14706 (N_14706,N_10069,N_10840);
and U14707 (N_14707,N_9441,N_9612);
and U14708 (N_14708,N_10232,N_11118);
and U14709 (N_14709,N_11424,N_9516);
nand U14710 (N_14710,N_9171,N_9521);
or U14711 (N_14711,N_10508,N_10295);
nor U14712 (N_14712,N_11830,N_11199);
or U14713 (N_14713,N_10739,N_9568);
nor U14714 (N_14714,N_10923,N_10525);
or U14715 (N_14715,N_10678,N_9507);
nand U14716 (N_14716,N_11360,N_9823);
or U14717 (N_14717,N_10905,N_9301);
nand U14718 (N_14718,N_10270,N_10612);
nand U14719 (N_14719,N_9626,N_11862);
nand U14720 (N_14720,N_10481,N_9678);
nand U14721 (N_14721,N_11850,N_10609);
and U14722 (N_14722,N_11730,N_10699);
and U14723 (N_14723,N_10406,N_9342);
nand U14724 (N_14724,N_9107,N_11387);
nand U14725 (N_14725,N_11256,N_10771);
nand U14726 (N_14726,N_11477,N_10308);
nand U14727 (N_14727,N_10608,N_10102);
nor U14728 (N_14728,N_11475,N_11260);
nor U14729 (N_14729,N_9149,N_9798);
or U14730 (N_14730,N_9734,N_9843);
and U14731 (N_14731,N_11254,N_9697);
or U14732 (N_14732,N_10599,N_10530);
nand U14733 (N_14733,N_11655,N_10598);
nor U14734 (N_14734,N_10882,N_9738);
nand U14735 (N_14735,N_10874,N_10148);
and U14736 (N_14736,N_9242,N_9390);
and U14737 (N_14737,N_9313,N_11624);
nand U14738 (N_14738,N_11453,N_11775);
and U14739 (N_14739,N_9165,N_9669);
and U14740 (N_14740,N_11414,N_10338);
nand U14741 (N_14741,N_10520,N_10742);
or U14742 (N_14742,N_11845,N_11916);
nand U14743 (N_14743,N_10898,N_9104);
or U14744 (N_14744,N_10498,N_10607);
nand U14745 (N_14745,N_10361,N_11652);
nand U14746 (N_14746,N_11702,N_10550);
and U14747 (N_14747,N_10211,N_9794);
or U14748 (N_14748,N_10946,N_11731);
nand U14749 (N_14749,N_10967,N_10250);
and U14750 (N_14750,N_9068,N_9232);
nor U14751 (N_14751,N_11891,N_11913);
or U14752 (N_14752,N_11974,N_11925);
and U14753 (N_14753,N_11459,N_10395);
and U14754 (N_14754,N_11610,N_11573);
and U14755 (N_14755,N_10970,N_9576);
and U14756 (N_14756,N_11259,N_11595);
nand U14757 (N_14757,N_9980,N_9567);
and U14758 (N_14758,N_11647,N_10478);
nor U14759 (N_14759,N_10984,N_9240);
nor U14760 (N_14760,N_11962,N_9530);
nand U14761 (N_14761,N_10873,N_11831);
and U14762 (N_14762,N_9674,N_10989);
or U14763 (N_14763,N_9821,N_11608);
and U14764 (N_14764,N_10899,N_9877);
nand U14765 (N_14765,N_11628,N_9827);
nand U14766 (N_14766,N_11824,N_10367);
nand U14767 (N_14767,N_11583,N_11513);
nand U14768 (N_14768,N_11345,N_11024);
and U14769 (N_14769,N_11818,N_9974);
and U14770 (N_14770,N_10502,N_9840);
and U14771 (N_14771,N_11801,N_10698);
xnor U14772 (N_14772,N_11264,N_10626);
or U14773 (N_14773,N_9755,N_11267);
or U14774 (N_14774,N_10702,N_9794);
and U14775 (N_14775,N_11313,N_10795);
and U14776 (N_14776,N_10016,N_9903);
nand U14777 (N_14777,N_11041,N_10190);
and U14778 (N_14778,N_10198,N_9858);
and U14779 (N_14779,N_10472,N_11751);
nor U14780 (N_14780,N_10520,N_10177);
and U14781 (N_14781,N_10546,N_10977);
and U14782 (N_14782,N_10128,N_11805);
or U14783 (N_14783,N_11235,N_9385);
nand U14784 (N_14784,N_10577,N_11493);
or U14785 (N_14785,N_11395,N_9469);
nand U14786 (N_14786,N_9107,N_10499);
and U14787 (N_14787,N_11616,N_11182);
and U14788 (N_14788,N_10116,N_10377);
or U14789 (N_14789,N_10784,N_10048);
or U14790 (N_14790,N_9142,N_10312);
and U14791 (N_14791,N_9262,N_9300);
or U14792 (N_14792,N_9371,N_11470);
nor U14793 (N_14793,N_10889,N_10926);
and U14794 (N_14794,N_10455,N_11906);
nor U14795 (N_14795,N_10222,N_10455);
or U14796 (N_14796,N_11716,N_10750);
or U14797 (N_14797,N_9660,N_9114);
and U14798 (N_14798,N_9212,N_10057);
and U14799 (N_14799,N_9377,N_10695);
and U14800 (N_14800,N_9162,N_11709);
and U14801 (N_14801,N_10723,N_11408);
and U14802 (N_14802,N_9476,N_9057);
nand U14803 (N_14803,N_10939,N_11269);
or U14804 (N_14804,N_11077,N_9513);
nor U14805 (N_14805,N_9257,N_11980);
nand U14806 (N_14806,N_11905,N_11795);
xnor U14807 (N_14807,N_11682,N_11952);
or U14808 (N_14808,N_9475,N_11951);
nor U14809 (N_14809,N_11764,N_11290);
and U14810 (N_14810,N_9931,N_10922);
nand U14811 (N_14811,N_11678,N_10133);
and U14812 (N_14812,N_10815,N_11806);
nand U14813 (N_14813,N_9345,N_11489);
and U14814 (N_14814,N_10256,N_10441);
nand U14815 (N_14815,N_9170,N_11836);
or U14816 (N_14816,N_11272,N_11712);
nand U14817 (N_14817,N_9897,N_9071);
nand U14818 (N_14818,N_11635,N_11479);
xnor U14819 (N_14819,N_9701,N_10653);
and U14820 (N_14820,N_9924,N_10292);
nand U14821 (N_14821,N_11509,N_10519);
nor U14822 (N_14822,N_9804,N_11722);
nand U14823 (N_14823,N_9314,N_9082);
nor U14824 (N_14824,N_10564,N_9809);
nor U14825 (N_14825,N_10225,N_9069);
or U14826 (N_14826,N_11141,N_10674);
nand U14827 (N_14827,N_11266,N_9525);
or U14828 (N_14828,N_10669,N_9258);
nor U14829 (N_14829,N_11037,N_10806);
nor U14830 (N_14830,N_11125,N_11153);
nand U14831 (N_14831,N_10559,N_10766);
or U14832 (N_14832,N_10836,N_9334);
or U14833 (N_14833,N_11855,N_11823);
nor U14834 (N_14834,N_11936,N_9653);
nand U14835 (N_14835,N_10046,N_9159);
and U14836 (N_14836,N_9773,N_10083);
and U14837 (N_14837,N_11980,N_9092);
nor U14838 (N_14838,N_10388,N_11694);
nor U14839 (N_14839,N_11343,N_9389);
nor U14840 (N_14840,N_11661,N_10262);
or U14841 (N_14841,N_9025,N_11345);
nor U14842 (N_14842,N_9924,N_9930);
or U14843 (N_14843,N_10042,N_10343);
nand U14844 (N_14844,N_10315,N_10189);
or U14845 (N_14845,N_11893,N_11330);
or U14846 (N_14846,N_10571,N_9761);
nand U14847 (N_14847,N_11938,N_10859);
or U14848 (N_14848,N_11672,N_11149);
and U14849 (N_14849,N_9080,N_9537);
nor U14850 (N_14850,N_9007,N_10104);
nand U14851 (N_14851,N_11990,N_9746);
or U14852 (N_14852,N_9341,N_10610);
or U14853 (N_14853,N_9134,N_10614);
nand U14854 (N_14854,N_11181,N_10928);
nand U14855 (N_14855,N_10357,N_10648);
nand U14856 (N_14856,N_9164,N_10034);
or U14857 (N_14857,N_11802,N_10925);
nor U14858 (N_14858,N_11187,N_10962);
nand U14859 (N_14859,N_9515,N_10831);
nor U14860 (N_14860,N_9207,N_9539);
nand U14861 (N_14861,N_11702,N_10176);
nand U14862 (N_14862,N_9260,N_10792);
and U14863 (N_14863,N_10207,N_11050);
and U14864 (N_14864,N_11035,N_10811);
nand U14865 (N_14865,N_11715,N_11725);
and U14866 (N_14866,N_10620,N_10035);
nor U14867 (N_14867,N_11992,N_9688);
or U14868 (N_14868,N_9238,N_9794);
or U14869 (N_14869,N_10456,N_9803);
and U14870 (N_14870,N_10247,N_10625);
nor U14871 (N_14871,N_10944,N_11061);
nor U14872 (N_14872,N_9945,N_11373);
nor U14873 (N_14873,N_9106,N_10267);
or U14874 (N_14874,N_9291,N_9808);
nand U14875 (N_14875,N_11950,N_10684);
nand U14876 (N_14876,N_10968,N_10713);
nor U14877 (N_14877,N_10738,N_10628);
and U14878 (N_14878,N_10671,N_9200);
or U14879 (N_14879,N_9307,N_9821);
nand U14880 (N_14880,N_11631,N_10551);
nand U14881 (N_14881,N_11426,N_11381);
or U14882 (N_14882,N_9460,N_11973);
nand U14883 (N_14883,N_11336,N_11732);
or U14884 (N_14884,N_10156,N_11734);
nor U14885 (N_14885,N_11539,N_9846);
and U14886 (N_14886,N_10904,N_10017);
and U14887 (N_14887,N_11500,N_9810);
and U14888 (N_14888,N_9563,N_10383);
nor U14889 (N_14889,N_9752,N_9881);
and U14890 (N_14890,N_9484,N_9010);
and U14891 (N_14891,N_10937,N_11175);
and U14892 (N_14892,N_10923,N_9125);
or U14893 (N_14893,N_11279,N_9872);
xor U14894 (N_14894,N_9589,N_10290);
nor U14895 (N_14895,N_10130,N_10161);
and U14896 (N_14896,N_10659,N_11963);
and U14897 (N_14897,N_11171,N_9568);
or U14898 (N_14898,N_11668,N_10772);
nor U14899 (N_14899,N_11770,N_11815);
and U14900 (N_14900,N_9662,N_11154);
or U14901 (N_14901,N_11797,N_9844);
and U14902 (N_14902,N_9550,N_11589);
nand U14903 (N_14903,N_11930,N_9282);
nor U14904 (N_14904,N_10981,N_9059);
and U14905 (N_14905,N_9913,N_11576);
nor U14906 (N_14906,N_11554,N_10857);
and U14907 (N_14907,N_10261,N_10269);
or U14908 (N_14908,N_11317,N_9428);
and U14909 (N_14909,N_9539,N_11035);
and U14910 (N_14910,N_11581,N_9831);
and U14911 (N_14911,N_9298,N_10421);
or U14912 (N_14912,N_11342,N_10753);
nand U14913 (N_14913,N_10394,N_10270);
nand U14914 (N_14914,N_9721,N_9788);
or U14915 (N_14915,N_9076,N_10694);
or U14916 (N_14916,N_10238,N_9004);
nor U14917 (N_14917,N_9668,N_11669);
and U14918 (N_14918,N_10793,N_9733);
and U14919 (N_14919,N_9742,N_10145);
nor U14920 (N_14920,N_11513,N_11527);
and U14921 (N_14921,N_9074,N_9985);
nor U14922 (N_14922,N_10193,N_11941);
nand U14923 (N_14923,N_11263,N_11087);
or U14924 (N_14924,N_10366,N_11419);
and U14925 (N_14925,N_9526,N_10267);
and U14926 (N_14926,N_9835,N_10020);
or U14927 (N_14927,N_9103,N_11955);
and U14928 (N_14928,N_10566,N_9128);
nor U14929 (N_14929,N_9292,N_10098);
nand U14930 (N_14930,N_10346,N_9224);
nand U14931 (N_14931,N_11645,N_9399);
and U14932 (N_14932,N_10552,N_11657);
nand U14933 (N_14933,N_10886,N_10084);
nand U14934 (N_14934,N_9071,N_9888);
nor U14935 (N_14935,N_9455,N_9591);
nand U14936 (N_14936,N_10020,N_11847);
nor U14937 (N_14937,N_10779,N_9639);
nor U14938 (N_14938,N_10520,N_11472);
or U14939 (N_14939,N_9173,N_10458);
nor U14940 (N_14940,N_10034,N_9630);
nor U14941 (N_14941,N_11190,N_9722);
nand U14942 (N_14942,N_10142,N_9528);
and U14943 (N_14943,N_9522,N_11040);
nor U14944 (N_14944,N_10676,N_10681);
nand U14945 (N_14945,N_11557,N_10634);
and U14946 (N_14946,N_10783,N_10560);
nand U14947 (N_14947,N_9869,N_11297);
nand U14948 (N_14948,N_9626,N_11370);
nand U14949 (N_14949,N_10187,N_9468);
and U14950 (N_14950,N_10728,N_10151);
nor U14951 (N_14951,N_11134,N_11010);
or U14952 (N_14952,N_11102,N_10017);
or U14953 (N_14953,N_11205,N_10404);
nor U14954 (N_14954,N_11436,N_10809);
or U14955 (N_14955,N_11420,N_10963);
or U14956 (N_14956,N_11149,N_10980);
nor U14957 (N_14957,N_9252,N_10302);
or U14958 (N_14958,N_9411,N_10422);
nand U14959 (N_14959,N_11411,N_11918);
nor U14960 (N_14960,N_10197,N_9202);
or U14961 (N_14961,N_9889,N_11584);
and U14962 (N_14962,N_11253,N_10142);
nor U14963 (N_14963,N_10903,N_10607);
nor U14964 (N_14964,N_11971,N_9889);
nand U14965 (N_14965,N_10585,N_9603);
and U14966 (N_14966,N_11220,N_11042);
nand U14967 (N_14967,N_9515,N_11761);
nor U14968 (N_14968,N_10672,N_11592);
nor U14969 (N_14969,N_11348,N_11757);
nor U14970 (N_14970,N_11781,N_11186);
and U14971 (N_14971,N_11498,N_9377);
or U14972 (N_14972,N_9993,N_9825);
nand U14973 (N_14973,N_9590,N_9128);
nand U14974 (N_14974,N_9672,N_10264);
or U14975 (N_14975,N_9650,N_10363);
nor U14976 (N_14976,N_10758,N_11424);
nor U14977 (N_14977,N_9367,N_9703);
or U14978 (N_14978,N_9918,N_9466);
and U14979 (N_14979,N_10443,N_9001);
nor U14980 (N_14980,N_11098,N_11024);
or U14981 (N_14981,N_10707,N_11194);
and U14982 (N_14982,N_11531,N_10057);
nor U14983 (N_14983,N_9156,N_9847);
nand U14984 (N_14984,N_9528,N_9935);
and U14985 (N_14985,N_10355,N_10832);
or U14986 (N_14986,N_10374,N_10999);
nand U14987 (N_14987,N_11149,N_9997);
nor U14988 (N_14988,N_9107,N_10839);
or U14989 (N_14989,N_10719,N_11316);
nand U14990 (N_14990,N_9337,N_10345);
nand U14991 (N_14991,N_9930,N_11963);
or U14992 (N_14992,N_9704,N_11967);
nand U14993 (N_14993,N_10458,N_9459);
or U14994 (N_14994,N_10771,N_11964);
nor U14995 (N_14995,N_10157,N_11449);
nor U14996 (N_14996,N_9181,N_10443);
or U14997 (N_14997,N_10853,N_11902);
and U14998 (N_14998,N_10594,N_9066);
and U14999 (N_14999,N_11579,N_10741);
and UO_0 (O_0,N_12683,N_12553);
nand UO_1 (O_1,N_13536,N_13130);
or UO_2 (O_2,N_12637,N_14259);
and UO_3 (O_3,N_12982,N_13301);
or UO_4 (O_4,N_14565,N_14919);
nor UO_5 (O_5,N_12459,N_12908);
nand UO_6 (O_6,N_13261,N_14521);
or UO_7 (O_7,N_13495,N_12787);
and UO_8 (O_8,N_13725,N_12007);
and UO_9 (O_9,N_12162,N_13432);
and UO_10 (O_10,N_12545,N_12979);
or UO_11 (O_11,N_12548,N_12572);
and UO_12 (O_12,N_14747,N_13383);
or UO_13 (O_13,N_12618,N_14878);
and UO_14 (O_14,N_12074,N_12730);
and UO_15 (O_15,N_13463,N_14978);
and UO_16 (O_16,N_13135,N_14831);
or UO_17 (O_17,N_14769,N_12053);
nand UO_18 (O_18,N_12764,N_13291);
nand UO_19 (O_19,N_14455,N_14116);
and UO_20 (O_20,N_14395,N_13281);
nor UO_21 (O_21,N_14266,N_13413);
nor UO_22 (O_22,N_14039,N_13029);
or UO_23 (O_23,N_12639,N_12839);
or UO_24 (O_24,N_12851,N_14588);
nor UO_25 (O_25,N_14037,N_12172);
or UO_26 (O_26,N_14572,N_14056);
nand UO_27 (O_27,N_14518,N_12139);
nor UO_28 (O_28,N_13238,N_13232);
or UO_29 (O_29,N_14091,N_13353);
or UO_30 (O_30,N_14360,N_14048);
and UO_31 (O_31,N_14967,N_13020);
nor UO_32 (O_32,N_12344,N_13717);
or UO_33 (O_33,N_14494,N_12242);
and UO_34 (O_34,N_12924,N_14851);
and UO_35 (O_35,N_12781,N_13943);
and UO_36 (O_36,N_12030,N_14064);
or UO_37 (O_37,N_14102,N_14576);
nand UO_38 (O_38,N_13501,N_12083);
and UO_39 (O_39,N_12786,N_14748);
and UO_40 (O_40,N_13877,N_13103);
and UO_41 (O_41,N_14844,N_12697);
or UO_42 (O_42,N_12339,N_13551);
nor UO_43 (O_43,N_12492,N_14160);
xnor UO_44 (O_44,N_12080,N_12811);
nand UO_45 (O_45,N_14819,N_13438);
or UO_46 (O_46,N_14589,N_13409);
or UO_47 (O_47,N_14886,N_13191);
and UO_48 (O_48,N_13671,N_13168);
and UO_49 (O_49,N_14935,N_12992);
and UO_50 (O_50,N_13543,N_13740);
nand UO_51 (O_51,N_13530,N_12834);
or UO_52 (O_52,N_13042,N_13842);
nor UO_53 (O_53,N_12830,N_12850);
nor UO_54 (O_54,N_14881,N_12766);
nand UO_55 (O_55,N_13480,N_13726);
nor UO_56 (O_56,N_12441,N_13751);
or UO_57 (O_57,N_13123,N_13069);
nor UO_58 (O_58,N_12825,N_13639);
nand UO_59 (O_59,N_13695,N_13876);
nor UO_60 (O_60,N_13679,N_12563);
or UO_61 (O_61,N_12779,N_12909);
and UO_62 (O_62,N_12867,N_12058);
and UO_63 (O_63,N_14045,N_14568);
xnor UO_64 (O_64,N_14816,N_12327);
and UO_65 (O_65,N_13444,N_14439);
or UO_66 (O_66,N_12422,N_14793);
nor UO_67 (O_67,N_14168,N_12624);
and UO_68 (O_68,N_13562,N_14250);
nor UO_69 (O_69,N_14574,N_12930);
or UO_70 (O_70,N_14185,N_13979);
or UO_71 (O_71,N_14535,N_13882);
and UO_72 (O_72,N_13361,N_13402);
nand UO_73 (O_73,N_13164,N_14800);
nor UO_74 (O_74,N_14854,N_12842);
nor UO_75 (O_75,N_14614,N_13110);
nor UO_76 (O_76,N_13371,N_13455);
or UO_77 (O_77,N_13124,N_14128);
nand UO_78 (O_78,N_13412,N_13381);
or UO_79 (O_79,N_12958,N_14660);
nor UO_80 (O_80,N_13484,N_12535);
and UO_81 (O_81,N_14483,N_14941);
and UO_82 (O_82,N_12975,N_12325);
or UO_83 (O_83,N_14170,N_12345);
and UO_84 (O_84,N_12282,N_12064);
nor UO_85 (O_85,N_13280,N_14108);
and UO_86 (O_86,N_12050,N_12686);
or UO_87 (O_87,N_12440,N_12451);
and UO_88 (O_88,N_12854,N_13584);
or UO_89 (O_89,N_13023,N_12102);
nor UO_90 (O_90,N_12833,N_13903);
nor UO_91 (O_91,N_14791,N_13490);
and UO_92 (O_92,N_14221,N_13324);
or UO_93 (O_93,N_12216,N_13532);
nand UO_94 (O_94,N_12933,N_14384);
and UO_95 (O_95,N_14964,N_13149);
nand UO_96 (O_96,N_13346,N_12285);
and UO_97 (O_97,N_13479,N_12439);
nor UO_98 (O_98,N_13190,N_13460);
and UO_99 (O_99,N_14686,N_13223);
or UO_100 (O_100,N_13090,N_14396);
and UO_101 (O_101,N_13678,N_14488);
and UO_102 (O_102,N_12034,N_12749);
xnor UO_103 (O_103,N_12201,N_13183);
nand UO_104 (O_104,N_14921,N_12466);
nor UO_105 (O_105,N_13665,N_13384);
nor UO_106 (O_106,N_13696,N_14290);
and UO_107 (O_107,N_13061,N_12799);
and UO_108 (O_108,N_13772,N_14449);
or UO_109 (O_109,N_12628,N_14173);
nand UO_110 (O_110,N_12679,N_13812);
nand UO_111 (O_111,N_12197,N_14106);
and UO_112 (O_112,N_14874,N_12525);
and UO_113 (O_113,N_14968,N_14047);
and UO_114 (O_114,N_14436,N_13959);
or UO_115 (O_115,N_14234,N_13635);
and UO_116 (O_116,N_14666,N_14688);
nand UO_117 (O_117,N_12420,N_12801);
or UO_118 (O_118,N_13956,N_13286);
nand UO_119 (O_119,N_12045,N_14226);
or UO_120 (O_120,N_12130,N_13390);
or UO_121 (O_121,N_12554,N_13252);
nor UO_122 (O_122,N_13598,N_13411);
nand UO_123 (O_123,N_14678,N_12215);
and UO_124 (O_124,N_14241,N_12230);
nor UO_125 (O_125,N_12990,N_12136);
and UO_126 (O_126,N_13711,N_12086);
or UO_127 (O_127,N_13937,N_12263);
or UO_128 (O_128,N_12612,N_13940);
and UO_129 (O_129,N_12134,N_14993);
nand UO_130 (O_130,N_14710,N_14562);
nand UO_131 (O_131,N_13850,N_13887);
and UO_132 (O_132,N_14302,N_12415);
or UO_133 (O_133,N_14619,N_13827);
and UO_134 (O_134,N_14719,N_14304);
or UO_135 (O_135,N_14520,N_13486);
nor UO_136 (O_136,N_13985,N_13995);
nand UO_137 (O_137,N_14277,N_13156);
nor UO_138 (O_138,N_13008,N_12988);
or UO_139 (O_139,N_14780,N_13583);
and UO_140 (O_140,N_14732,N_14848);
nor UO_141 (O_141,N_13356,N_13893);
and UO_142 (O_142,N_13556,N_12667);
or UO_143 (O_143,N_14708,N_14069);
nand UO_144 (O_144,N_14997,N_13651);
or UO_145 (O_145,N_12425,N_14492);
and UO_146 (O_146,N_14669,N_14319);
or UO_147 (O_147,N_14852,N_14639);
or UO_148 (O_148,N_12721,N_14388);
nor UO_149 (O_149,N_12722,N_12835);
nand UO_150 (O_150,N_13227,N_14104);
nor UO_151 (O_151,N_12755,N_12497);
nor UO_152 (O_152,N_14672,N_13716);
or UO_153 (O_153,N_12557,N_13749);
or UO_154 (O_154,N_14510,N_12129);
and UO_155 (O_155,N_13660,N_12896);
xnor UO_156 (O_156,N_13563,N_14677);
nor UO_157 (O_157,N_14784,N_14552);
and UO_158 (O_158,N_14165,N_14201);
nor UO_159 (O_159,N_13265,N_12915);
or UO_160 (O_160,N_14254,N_14391);
nand UO_161 (O_161,N_12538,N_12537);
nor UO_162 (O_162,N_12812,N_14286);
and UO_163 (O_163,N_14136,N_14551);
or UO_164 (O_164,N_12310,N_14306);
or UO_165 (O_165,N_12181,N_14785);
and UO_166 (O_166,N_13987,N_13976);
nor UO_167 (O_167,N_13552,N_13923);
or UO_168 (O_168,N_12632,N_14138);
nand UO_169 (O_169,N_12360,N_13761);
or UO_170 (O_170,N_12144,N_13092);
nand UO_171 (O_171,N_14316,N_12886);
nand UO_172 (O_172,N_13694,N_13058);
nor UO_173 (O_173,N_13091,N_12752);
and UO_174 (O_174,N_14973,N_12790);
nand UO_175 (O_175,N_12324,N_12318);
or UO_176 (O_176,N_12665,N_13690);
and UO_177 (O_177,N_13147,N_14346);
and UO_178 (O_178,N_12206,N_13133);
nand UO_179 (O_179,N_13429,N_14216);
or UO_180 (O_180,N_14801,N_13874);
nand UO_181 (O_181,N_13853,N_13992);
and UO_182 (O_182,N_13632,N_12288);
and UO_183 (O_183,N_14808,N_12974);
and UO_184 (O_184,N_14654,N_14125);
and UO_185 (O_185,N_12925,N_13759);
or UO_186 (O_186,N_12556,N_14726);
nor UO_187 (O_187,N_13382,N_12753);
or UO_188 (O_188,N_14385,N_12294);
and UO_189 (O_189,N_14390,N_12750);
nor UO_190 (O_190,N_12902,N_14853);
and UO_191 (O_191,N_12953,N_12555);
nor UO_192 (O_192,N_14541,N_14132);
or UO_193 (O_193,N_12617,N_14904);
and UO_194 (O_194,N_13854,N_13684);
and UO_195 (O_195,N_14673,N_14189);
nand UO_196 (O_196,N_12037,N_14841);
nor UO_197 (O_197,N_14053,N_13752);
nor UO_198 (O_198,N_13952,N_13268);
nor UO_199 (O_199,N_12253,N_13861);
nor UO_200 (O_200,N_13006,N_12533);
and UO_201 (O_201,N_12245,N_12499);
nand UO_202 (O_202,N_12368,N_14087);
nor UO_203 (O_203,N_12237,N_14190);
or UO_204 (O_204,N_12448,N_14187);
or UO_205 (O_205,N_13834,N_14075);
or UO_206 (O_206,N_14466,N_12770);
nand UO_207 (O_207,N_12212,N_14570);
or UO_208 (O_208,N_13811,N_12540);
and UO_209 (O_209,N_12587,N_12341);
or UO_210 (O_210,N_14662,N_13662);
or UO_211 (O_211,N_13450,N_14479);
nor UO_212 (O_212,N_13293,N_13314);
and UO_213 (O_213,N_13546,N_13847);
or UO_214 (O_214,N_12493,N_13054);
nand UO_215 (O_215,N_12380,N_14295);
nor UO_216 (O_216,N_12771,N_13278);
and UO_217 (O_217,N_13554,N_14827);
nand UO_218 (O_218,N_14725,N_13735);
or UO_219 (O_219,N_13487,N_13819);
nor UO_220 (O_220,N_13106,N_14507);
and UO_221 (O_221,N_13626,N_14776);
and UO_222 (O_222,N_13407,N_14786);
nor UO_223 (O_223,N_12168,N_13604);
or UO_224 (O_224,N_12932,N_12071);
nand UO_225 (O_225,N_13951,N_12396);
and UO_226 (O_226,N_13055,N_12106);
or UO_227 (O_227,N_12916,N_14749);
nand UO_228 (O_228,N_12987,N_14199);
or UO_229 (O_229,N_12240,N_14743);
nand UO_230 (O_230,N_14958,N_12120);
and UO_231 (O_231,N_13277,N_12137);
and UO_232 (O_232,N_14322,N_14006);
and UO_233 (O_233,N_12250,N_13445);
and UO_234 (O_234,N_13814,N_12507);
nand UO_235 (O_235,N_14086,N_14717);
and UO_236 (O_236,N_12797,N_12276);
nor UO_237 (O_237,N_13362,N_13722);
nand UO_238 (O_238,N_12414,N_14214);
nand UO_239 (O_239,N_14381,N_14327);
or UO_240 (O_240,N_13978,N_14947);
nand UO_241 (O_241,N_13083,N_13049);
and UO_242 (O_242,N_14358,N_12211);
nor UO_243 (O_243,N_12574,N_14705);
and UO_244 (O_244,N_14498,N_13755);
and UO_245 (O_245,N_14171,N_12528);
and UO_246 (O_246,N_13786,N_13097);
nand UO_247 (O_247,N_14410,N_13521);
nor UO_248 (O_248,N_12482,N_13003);
nor UO_249 (O_249,N_14680,N_13677);
nor UO_250 (O_250,N_14580,N_12534);
nand UO_251 (O_251,N_12596,N_12798);
or UO_252 (O_252,N_13715,N_13573);
or UO_253 (O_253,N_14446,N_14134);
nor UO_254 (O_254,N_13137,N_12523);
or UO_255 (O_255,N_13829,N_14735);
and UO_256 (O_256,N_13802,N_12911);
nand UO_257 (O_257,N_14975,N_13576);
nor UO_258 (O_258,N_13166,N_14882);
or UO_259 (O_259,N_13197,N_14228);
nand UO_260 (O_260,N_12702,N_13421);
and UO_261 (O_261,N_14901,N_13560);
nor UO_262 (O_262,N_13306,N_14811);
nand UO_263 (O_263,N_14247,N_13060);
or UO_264 (O_264,N_12619,N_14714);
and UO_265 (O_265,N_13880,N_13770);
and UO_266 (O_266,N_14105,N_14865);
or UO_267 (O_267,N_14100,N_13084);
and UO_268 (O_268,N_13121,N_12849);
nand UO_269 (O_269,N_14411,N_13505);
or UO_270 (O_270,N_14746,N_13958);
and UO_271 (O_271,N_12822,N_12061);
nor UO_272 (O_272,N_14500,N_14657);
nand UO_273 (O_273,N_12783,N_12235);
and UO_274 (O_274,N_14573,N_12984);
or UO_275 (O_275,N_14712,N_12936);
or UO_276 (O_276,N_13212,N_13736);
or UO_277 (O_277,N_14179,N_14379);
or UO_278 (O_278,N_14276,N_13840);
and UO_279 (O_279,N_13035,N_12186);
nand UO_280 (O_280,N_13763,N_12377);
nand UO_281 (O_281,N_14202,N_14974);
nor UO_282 (O_282,N_14354,N_12550);
nor UO_283 (O_283,N_13417,N_14505);
nand UO_284 (O_284,N_13435,N_14015);
nand UO_285 (O_285,N_12163,N_13247);
nor UO_286 (O_286,N_12154,N_14465);
and UO_287 (O_287,N_13406,N_14602);
nand UO_288 (O_288,N_12336,N_14691);
or UO_289 (O_289,N_13119,N_14945);
nand UO_290 (O_290,N_14009,N_13270);
and UO_291 (O_291,N_14055,N_14699);
and UO_292 (O_292,N_14151,N_12855);
nor UO_293 (O_293,N_14166,N_12692);
nor UO_294 (O_294,N_13920,N_12320);
and UO_295 (O_295,N_12452,N_12880);
and UO_296 (O_296,N_12435,N_13145);
nand UO_297 (O_297,N_14547,N_14989);
or UO_298 (O_298,N_12899,N_13585);
nand UO_299 (O_299,N_14509,N_13437);
nand UO_300 (O_300,N_13509,N_14493);
nand UO_301 (O_301,N_14907,N_14491);
nand UO_302 (O_302,N_13013,N_12551);
and UO_303 (O_303,N_13670,N_14647);
or UO_304 (O_304,N_14137,N_12765);
nor UO_305 (O_305,N_14689,N_14652);
nor UO_306 (O_306,N_12814,N_13482);
or UO_307 (O_307,N_12273,N_14164);
nand UO_308 (O_308,N_12893,N_14453);
and UO_309 (O_309,N_14835,N_12028);
and UO_310 (O_310,N_13698,N_14549);
nand UO_311 (O_311,N_13875,N_12810);
and UO_312 (O_312,N_12238,N_12881);
or UO_313 (O_313,N_13713,N_12733);
and UO_314 (O_314,N_14133,N_14774);
nor UO_315 (O_315,N_14583,N_13625);
or UO_316 (O_316,N_12701,N_13969);
and UO_317 (O_317,N_13082,N_14367);
nand UO_318 (O_318,N_12606,N_12910);
and UO_319 (O_319,N_14879,N_13424);
nand UO_320 (O_320,N_14406,N_14750);
nor UO_321 (O_321,N_13204,N_12657);
and UO_322 (O_322,N_12141,N_14068);
nand UO_323 (O_323,N_14093,N_12438);
and UO_324 (O_324,N_14739,N_13640);
and UO_325 (O_325,N_14523,N_13897);
or UO_326 (O_326,N_14681,N_14764);
nor UO_327 (O_327,N_13174,N_12705);
and UO_328 (O_328,N_12200,N_14584);
nand UO_329 (O_329,N_14107,N_14145);
nor UO_330 (O_330,N_14153,N_12542);
nand UO_331 (O_331,N_14722,N_14161);
nor UO_332 (O_332,N_13768,N_12152);
nor UO_333 (O_333,N_13224,N_12042);
nor UO_334 (O_334,N_14707,N_12605);
and UO_335 (O_335,N_12309,N_12195);
nor UO_336 (O_336,N_12623,N_14273);
or UO_337 (O_337,N_14352,N_13701);
or UO_338 (O_338,N_12408,N_14423);
or UO_339 (O_339,N_12473,N_14641);
and UO_340 (O_340,N_13890,N_12708);
or UO_341 (O_341,N_12860,N_14034);
nor UO_342 (O_342,N_13271,N_12664);
nand UO_343 (O_343,N_14545,N_13544);
nor UO_344 (O_344,N_12960,N_13313);
nand UO_345 (O_345,N_13955,N_14289);
and UO_346 (O_346,N_13970,N_13099);
and UO_347 (O_347,N_13275,N_13192);
nor UO_348 (O_348,N_14083,N_13433);
or UO_349 (O_349,N_14099,N_13799);
and UO_350 (O_350,N_14649,N_13400);
nand UO_351 (O_351,N_12391,N_12434);
and UO_352 (O_352,N_12189,N_13366);
and UO_353 (O_353,N_14752,N_14976);
nor UO_354 (O_354,N_13915,N_14771);
nor UO_355 (O_355,N_14617,N_13865);
or UO_356 (O_356,N_14790,N_14194);
nor UO_357 (O_357,N_14251,N_14581);
nor UO_358 (O_358,N_12374,N_12808);
and UO_359 (O_359,N_14338,N_12496);
nand UO_360 (O_360,N_12455,N_12944);
nand UO_361 (O_361,N_12820,N_13900);
and UO_362 (O_362,N_14868,N_14903);
nor UO_363 (O_363,N_12476,N_12026);
xor UO_364 (O_364,N_13687,N_13986);
and UO_365 (O_365,N_13493,N_14309);
nand UO_366 (O_366,N_13352,N_13373);
nor UO_367 (O_367,N_12062,N_12871);
and UO_368 (O_368,N_12922,N_13938);
nor UO_369 (O_369,N_13385,N_12760);
or UO_370 (O_370,N_12888,N_13650);
nand UO_371 (O_371,N_14524,N_13253);
nor UO_372 (O_372,N_13578,N_14114);
nand UO_373 (O_373,N_13870,N_12486);
nor UO_374 (O_374,N_12449,N_13685);
nand UO_375 (O_375,N_13916,N_12337);
nor UO_376 (O_376,N_12609,N_14996);
nor UO_377 (O_377,N_14939,N_13977);
or UO_378 (O_378,N_12373,N_14644);
and UO_379 (O_379,N_13838,N_14920);
or UO_380 (O_380,N_12196,N_13471);
or UO_381 (O_381,N_12367,N_12681);
or UO_382 (O_382,N_12308,N_12502);
and UO_383 (O_383,N_12052,N_12983);
nor UO_384 (O_384,N_14307,N_13781);
nor UO_385 (O_385,N_13194,N_14761);
or UO_386 (O_386,N_13264,N_13776);
and UO_387 (O_387,N_14017,N_12478);
nand UO_388 (O_388,N_13209,N_14877);
nand UO_389 (O_389,N_13791,N_12358);
nor UO_390 (O_390,N_14632,N_13141);
and UO_391 (O_391,N_14329,N_12109);
and UO_392 (O_392,N_13185,N_13872);
and UO_393 (O_393,N_13581,N_12720);
nand UO_394 (O_394,N_12277,N_13279);
or UO_395 (O_395,N_12468,N_13451);
or UO_396 (O_396,N_13007,N_12219);
and UO_397 (O_397,N_13410,N_14427);
or UO_398 (O_398,N_12445,N_13300);
nand UO_399 (O_399,N_12539,N_13467);
nand UO_400 (O_400,N_12464,N_14067);
or UO_401 (O_401,N_14540,N_13052);
nand UO_402 (O_402,N_14667,N_14721);
or UO_403 (O_403,N_12387,N_12359);
nor UO_404 (O_404,N_14817,N_13704);
nor UO_405 (O_405,N_13188,N_12937);
or UO_406 (O_406,N_14536,N_14078);
nor UO_407 (O_407,N_12182,N_12920);
or UO_408 (O_408,N_12316,N_14651);
nor UO_409 (O_409,N_14419,N_12218);
or UO_410 (O_410,N_14548,N_13912);
nor UO_411 (O_411,N_12031,N_12393);
and UO_412 (O_412,N_13967,N_12104);
nor UO_413 (O_413,N_14859,N_13608);
nand UO_414 (O_414,N_12207,N_12500);
nor UO_415 (O_415,N_12430,N_13873);
nand UO_416 (O_416,N_13334,N_13964);
nand UO_417 (O_417,N_12389,N_12291);
nand UO_418 (O_418,N_12398,N_13004);
nand UO_419 (O_419,N_12576,N_13729);
nand UO_420 (O_420,N_12194,N_14624);
nor UO_421 (O_421,N_13215,N_13442);
nor UO_422 (O_422,N_12520,N_14040);
nor UO_423 (O_423,N_12188,N_12929);
nand UO_424 (O_424,N_14842,N_14713);
or UO_425 (O_425,N_13966,N_12517);
or UO_426 (O_426,N_13221,N_14495);
and UO_427 (O_427,N_13071,N_14336);
nor UO_428 (O_428,N_14715,N_12123);
nand UO_429 (O_429,N_13528,N_13021);
nand UO_430 (O_430,N_13456,N_13533);
nand UO_431 (O_431,N_14060,N_14755);
and UO_432 (O_432,N_14013,N_13350);
nand UO_433 (O_433,N_14288,N_12895);
nor UO_434 (O_434,N_13102,N_12780);
nand UO_435 (O_435,N_12068,N_14422);
nand UO_436 (O_436,N_14528,N_13804);
and UO_437 (O_437,N_12119,N_12223);
nor UO_438 (O_438,N_12952,N_13093);
or UO_439 (O_439,N_13683,N_14534);
or UO_440 (O_440,N_12856,N_13100);
nor UO_441 (O_441,N_14267,N_13053);
nand UO_442 (O_442,N_13594,N_13045);
nand UO_443 (O_443,N_13512,N_13918);
and UO_444 (O_444,N_12180,N_12234);
and UO_445 (O_445,N_12647,N_12460);
and UO_446 (O_446,N_13165,N_12643);
and UO_447 (O_447,N_13862,N_13138);
or UO_448 (O_448,N_14071,N_12529);
xor UO_449 (O_449,N_14058,N_13550);
nor UO_450 (O_450,N_13750,N_14292);
nor UO_451 (O_451,N_13094,N_14402);
nand UO_452 (O_452,N_14450,N_13559);
nand UO_453 (O_453,N_12997,N_12055);
or UO_454 (O_454,N_13311,N_13038);
or UO_455 (O_455,N_14249,N_12477);
and UO_456 (O_456,N_13089,N_14608);
nand UO_457 (O_457,N_13997,N_13901);
and UO_458 (O_458,N_14012,N_12541);
nor UO_459 (O_459,N_12513,N_14861);
nand UO_460 (O_460,N_13282,N_14730);
or UO_461 (O_461,N_12480,N_12652);
nand UO_462 (O_462,N_12133,N_13234);
nor UO_463 (O_463,N_12066,N_14377);
and UO_464 (O_464,N_13499,N_13290);
nand UO_465 (O_465,N_12405,N_14413);
nand UO_466 (O_466,N_12254,N_12942);
or UO_467 (O_467,N_14910,N_12763);
and UO_468 (O_468,N_13675,N_13262);
nand UO_469 (O_469,N_13700,N_13333);
or UO_470 (O_470,N_12257,N_12883);
nor UO_471 (O_471,N_14020,N_13283);
or UO_472 (O_472,N_14183,N_13960);
and UO_473 (O_473,N_12735,N_14312);
or UO_474 (O_474,N_12791,N_14155);
nand UO_475 (O_475,N_13513,N_13886);
and UO_476 (O_476,N_14701,N_13464);
or UO_477 (O_477,N_12424,N_14629);
or UO_478 (O_478,N_12272,N_13538);
or UO_479 (O_479,N_12311,N_14582);
and UO_480 (O_480,N_12584,N_13498);
nand UO_481 (O_481,N_14962,N_14598);
nor UO_482 (O_482,N_12018,N_13201);
nand UO_483 (O_483,N_13179,N_14026);
or UO_484 (O_484,N_14872,N_12560);
nand UO_485 (O_485,N_14777,N_14731);
nand UO_486 (O_486,N_13048,N_13496);
nand UO_487 (O_487,N_14981,N_14330);
or UO_488 (O_488,N_14522,N_14404);
nor UO_489 (O_489,N_13941,N_13375);
and UO_490 (O_490,N_13401,N_12829);
or UO_491 (O_491,N_12543,N_14397);
or UO_492 (O_492,N_13558,N_14796);
or UO_493 (O_493,N_13758,N_13965);
nor UO_494 (O_494,N_13974,N_13624);
nand UO_495 (O_495,N_14952,N_13387);
or UO_496 (O_496,N_12383,N_12229);
and UO_497 (O_497,N_12178,N_14866);
nand UO_498 (O_498,N_12734,N_12577);
and UO_499 (O_499,N_12140,N_12857);
nand UO_500 (O_500,N_14511,N_14938);
nand UO_501 (O_501,N_13611,N_13601);
nor UO_502 (O_502,N_14979,N_14825);
nor UO_503 (O_503,N_14613,N_12699);
and UO_504 (O_504,N_13936,N_12522);
or UO_505 (O_505,N_14196,N_13393);
nor UO_506 (O_506,N_12912,N_12029);
nor UO_507 (O_507,N_13222,N_12578);
or UO_508 (O_508,N_14248,N_12192);
nand UO_509 (O_509,N_14659,N_13643);
or UO_510 (O_510,N_13591,N_12190);
or UO_511 (O_511,N_12661,N_14059);
or UO_512 (O_512,N_12267,N_13125);
and UO_513 (O_513,N_14625,N_13753);
nand UO_514 (O_514,N_13186,N_12084);
nor UO_515 (O_515,N_13888,N_14113);
and UO_516 (O_516,N_12845,N_14265);
nand UO_517 (O_517,N_14308,N_14516);
or UO_518 (O_518,N_14029,N_13351);
or UO_519 (O_519,N_14437,N_14019);
and UO_520 (O_520,N_14257,N_13285);
or UO_521 (O_521,N_13065,N_13173);
and UO_522 (O_522,N_12570,N_14127);
and UO_523 (O_523,N_12530,N_14252);
nand UO_524 (O_524,N_14923,N_13681);
nor UO_525 (O_525,N_13619,N_14043);
nand UO_526 (O_526,N_13502,N_14418);
nor UO_527 (O_527,N_14604,N_13308);
nor UO_528 (O_528,N_12268,N_13294);
nor UO_529 (O_529,N_14256,N_13792);
or UO_530 (O_530,N_13878,N_12082);
or UO_531 (O_531,N_12846,N_12917);
or UO_532 (O_532,N_13636,N_12595);
nand UO_533 (O_533,N_13266,N_14334);
or UO_534 (O_534,N_14564,N_14766);
nand UO_535 (O_535,N_14481,N_13833);
nand UO_536 (O_536,N_13746,N_13195);
nand UO_537 (O_537,N_14373,N_12298);
nand UO_538 (O_538,N_14463,N_12159);
nand UO_539 (O_539,N_14955,N_12299);
or UO_540 (O_540,N_12091,N_13259);
nand UO_541 (O_541,N_13358,N_13810);
nand UO_542 (O_542,N_14569,N_14931);
nor UO_543 (O_543,N_14467,N_13386);
nand UO_544 (O_544,N_13789,N_12655);
or UO_545 (O_545,N_14880,N_12634);
nand UO_546 (O_546,N_13949,N_13068);
or UO_547 (O_547,N_13218,N_12488);
nor UO_548 (O_548,N_12103,N_14805);
nor UO_549 (O_549,N_14345,N_13365);
nor UO_550 (O_550,N_12041,N_12409);
nor UO_551 (O_551,N_12264,N_13516);
and UO_552 (O_552,N_12934,N_14943);
nand UO_553 (O_553,N_12868,N_12989);
nor UO_554 (O_554,N_13254,N_13771);
and UO_555 (O_555,N_13708,N_14407);
or UO_556 (O_556,N_12003,N_12390);
and UO_557 (O_557,N_12889,N_12817);
and UO_558 (O_558,N_14870,N_13564);
nor UO_559 (O_559,N_13140,N_14553);
and UO_560 (O_560,N_12890,N_12012);
nor UO_561 (O_561,N_13523,N_13835);
and UO_562 (O_562,N_13322,N_14698);
nand UO_563 (O_563,N_13040,N_14706);
nor UO_564 (O_564,N_14095,N_12711);
nand UO_565 (O_565,N_12155,N_13710);
and UO_566 (O_566,N_13744,N_13086);
nor UO_567 (O_567,N_14143,N_14366);
nor UO_568 (O_568,N_12796,N_13593);
or UO_569 (O_569,N_14300,N_12458);
nand UO_570 (O_570,N_14860,N_12950);
and UO_571 (O_571,N_14115,N_13911);
nor UO_572 (O_572,N_13263,N_12411);
or UO_573 (O_573,N_13963,N_14834);
nor UO_574 (O_574,N_14728,N_13064);
nor UO_575 (O_575,N_13132,N_13009);
nand UO_576 (O_576,N_14471,N_14224);
and UO_577 (O_577,N_12597,N_12354);
or UO_578 (O_578,N_14150,N_13288);
and UO_579 (O_579,N_13659,N_14839);
nand UO_580 (O_580,N_13800,N_12069);
and UO_581 (O_581,N_12521,N_12590);
and UO_582 (O_582,N_14030,N_14084);
or UO_583 (O_583,N_14081,N_14661);
nand UO_584 (O_584,N_12504,N_12032);
nand UO_585 (O_585,N_14092,N_13778);
and UO_586 (O_586,N_12005,N_12802);
and UO_587 (O_587,N_12739,N_14229);
nor UO_588 (O_588,N_12056,N_12125);
and UO_589 (O_589,N_14464,N_13397);
or UO_590 (O_590,N_13907,N_12748);
or UO_591 (O_591,N_13414,N_12020);
nor UO_592 (O_592,N_13515,N_12147);
or UO_593 (O_593,N_14124,N_13524);
nor UO_594 (O_594,N_12094,N_13545);
or UO_595 (O_595,N_13014,N_12173);
nand UO_596 (O_596,N_13742,N_14895);
and UO_597 (O_597,N_14995,N_13806);
nor UO_598 (O_598,N_14959,N_14736);
or UO_599 (O_599,N_14648,N_12099);
nor UO_600 (O_600,N_14566,N_12295);
nor UO_601 (O_601,N_12397,N_14264);
nand UO_602 (O_602,N_12048,N_13830);
or UO_603 (O_603,N_12232,N_14533);
or UO_604 (O_604,N_14441,N_12290);
nor UO_605 (O_605,N_14798,N_13507);
and UO_606 (O_606,N_13196,N_13289);
or UO_607 (O_607,N_14814,N_13000);
or UO_608 (O_608,N_14121,N_13112);
nor UO_609 (O_609,N_14775,N_12809);
or UO_610 (O_610,N_12171,N_14129);
nor UO_611 (O_611,N_12687,N_12593);
nand UO_612 (O_612,N_13914,N_13844);
nor UO_613 (O_613,N_12292,N_13453);
and UO_614 (O_614,N_12759,N_14956);
nand UO_615 (O_615,N_12406,N_14826);
and UO_616 (O_616,N_14237,N_14222);
nor UO_617 (O_617,N_12970,N_14531);
xor UO_618 (O_618,N_14514,N_14460);
or UO_619 (O_619,N_14754,N_14260);
nand UO_620 (O_620,N_14044,N_12227);
nor UO_621 (O_621,N_13628,N_14832);
nand UO_622 (O_622,N_13026,N_13320);
nand UO_623 (O_623,N_12421,N_12343);
nand UO_624 (O_624,N_13982,N_14633);
and UO_625 (O_625,N_14656,N_12670);
or UO_626 (O_626,N_13692,N_13826);
and UO_627 (O_627,N_14760,N_14900);
or UO_628 (O_628,N_12305,N_13404);
nand UO_629 (O_629,N_13469,N_13056);
or UO_630 (O_630,N_14906,N_13323);
and UO_631 (O_631,N_13648,N_13723);
nand UO_632 (O_632,N_13883,N_12913);
or UO_633 (O_633,N_12379,N_13654);
or UO_634 (O_634,N_13175,N_14812);
and UO_635 (O_635,N_13927,N_14139);
nand UO_636 (O_636,N_12688,N_13709);
nor UO_637 (O_637,N_12089,N_12033);
nand UO_638 (O_638,N_12142,N_14175);
nor UO_639 (O_639,N_12816,N_12220);
nand UO_640 (O_640,N_13131,N_14451);
and UO_641 (O_641,N_13503,N_12284);
nand UO_642 (O_642,N_14543,N_14085);
or UO_643 (O_643,N_13730,N_12717);
nand UO_644 (O_644,N_14490,N_12959);
nor UO_645 (O_645,N_14035,N_12401);
nor UO_646 (O_646,N_12536,N_13531);
and UO_647 (O_647,N_14837,N_13318);
nor UO_648 (O_648,N_12625,N_13793);
nand UO_649 (O_649,N_13572,N_13919);
nand UO_650 (O_650,N_14429,N_13483);
nand UO_651 (O_651,N_12407,N_13561);
or UO_652 (O_652,N_13714,N_12662);
and UO_653 (O_653,N_14847,N_14169);
nand UO_654 (O_654,N_12145,N_13721);
and UO_655 (O_655,N_12704,N_13425);
and UO_656 (O_656,N_12185,N_12261);
nor UO_657 (O_657,N_13330,N_14922);
and UO_658 (O_658,N_13154,N_13299);
and UO_659 (O_659,N_12579,N_14664);
or UO_660 (O_660,N_13539,N_14884);
nor UO_661 (O_661,N_13863,N_12600);
nor UO_662 (O_662,N_13249,N_14405);
nand UO_663 (O_663,N_14002,N_13688);
nand UO_664 (O_664,N_14753,N_12673);
or UO_665 (O_665,N_12741,N_13120);
nand UO_666 (O_666,N_14342,N_13213);
nor UO_667 (O_667,N_14845,N_14041);
nand UO_668 (O_668,N_14970,N_14212);
nor UO_669 (O_669,N_14687,N_14403);
and UO_670 (O_670,N_14890,N_12977);
or UO_671 (O_671,N_13163,N_12350);
or UO_672 (O_672,N_14615,N_14733);
nor UO_673 (O_673,N_12636,N_14949);
or UO_674 (O_674,N_12143,N_12225);
nand UO_675 (O_675,N_14486,N_12111);
nor UO_676 (O_676,N_14089,N_14577);
nor UO_677 (O_677,N_13649,N_13780);
nor UO_678 (O_678,N_12392,N_13085);
or UO_679 (O_679,N_13151,N_12241);
nand UO_680 (O_680,N_13537,N_14090);
and UO_681 (O_681,N_14944,N_12231);
and UO_682 (O_682,N_12450,N_13569);
nand UO_683 (O_683,N_12386,N_14770);
nand UO_684 (O_684,N_14571,N_13764);
nand UO_685 (O_685,N_12426,N_12465);
and UO_686 (O_686,N_14062,N_13022);
nor UO_687 (O_687,N_14783,N_14645);
nand UO_688 (O_688,N_13818,N_13975);
nor UO_689 (O_689,N_13743,N_13128);
nor UO_690 (O_690,N_14223,N_13187);
nand UO_691 (O_691,N_13566,N_12093);
and UO_692 (O_692,N_12718,N_12805);
nand UO_693 (O_693,N_14435,N_14293);
and UO_694 (O_694,N_13950,N_12645);
nand UO_695 (O_695,N_14781,N_14530);
nand UO_696 (O_696,N_12827,N_12736);
nand UO_697 (O_697,N_13015,N_13345);
or UO_698 (O_698,N_12601,N_12063);
or UO_699 (O_699,N_13517,N_13615);
or UO_700 (O_700,N_13160,N_12124);
nand UO_701 (O_701,N_12611,N_14028);
nor UO_702 (O_702,N_13666,N_12745);
nor UO_703 (O_703,N_13557,N_12901);
and UO_704 (O_704,N_13592,N_13329);
nor UO_705 (O_705,N_12585,N_14263);
or UO_706 (O_706,N_12485,N_13305);
nand UO_707 (O_707,N_12249,N_13565);
nor UO_708 (O_708,N_12985,N_14317);
nor UO_709 (O_709,N_14156,N_14557);
nor UO_710 (O_710,N_12274,N_12402);
or UO_711 (O_711,N_12728,N_14579);
or UO_712 (O_712,N_14003,N_12598);
and UO_713 (O_713,N_14515,N_12244);
nand UO_714 (O_714,N_14809,N_13292);
nor UO_715 (O_715,N_14176,N_14112);
nor UO_716 (O_716,N_13555,N_13599);
nor UO_717 (O_717,N_12519,N_13932);
nor UO_718 (O_718,N_12353,N_14912);
and UO_719 (O_719,N_12051,N_13113);
and UO_720 (O_720,N_13645,N_14502);
nand UO_721 (O_721,N_14799,N_12203);
xor UO_722 (O_722,N_14454,N_12331);
or UO_723 (O_723,N_13219,N_13142);
and UO_724 (O_724,N_13674,N_12561);
nor UO_725 (O_725,N_12454,N_14188);
and UO_726 (O_726,N_13779,N_12546);
or UO_727 (O_727,N_13150,N_12602);
or UO_728 (O_728,N_13474,N_14443);
nor UO_729 (O_729,N_12304,N_14262);
or UO_730 (O_730,N_13757,N_14773);
or UO_731 (O_731,N_14258,N_12967);
or UO_732 (O_732,N_13989,N_14314);
or UO_733 (O_733,N_14430,N_14897);
nand UO_734 (O_734,N_14909,N_12644);
and UO_735 (O_735,N_14496,N_13734);
nor UO_736 (O_736,N_12986,N_14742);
nand UO_737 (O_737,N_13889,N_12199);
nand UO_738 (O_738,N_14274,N_14409);
nor UO_739 (O_739,N_13379,N_13646);
nand UO_740 (O_740,N_14593,N_13618);
or UO_741 (O_741,N_14272,N_12947);
and UO_742 (O_742,N_13245,N_12092);
nand UO_743 (O_743,N_14616,N_13707);
nand UO_744 (O_744,N_14740,N_12236);
or UO_745 (O_745,N_14014,N_13848);
nor UO_746 (O_746,N_14054,N_14695);
or UO_747 (O_747,N_12991,N_13198);
xnor UO_748 (O_748,N_13816,N_14804);
nand UO_749 (O_749,N_12118,N_12315);
and UO_750 (O_750,N_12626,N_14361);
nor UO_751 (O_751,N_12737,N_13111);
or UO_752 (O_752,N_12117,N_14525);
nand UO_753 (O_753,N_13237,N_14117);
or UO_754 (O_754,N_12076,N_12583);
and UO_755 (O_755,N_14122,N_12491);
xor UO_756 (O_756,N_14324,N_13851);
xor UO_757 (O_757,N_12754,N_13845);
nand UO_758 (O_758,N_12075,N_12691);
nand UO_759 (O_759,N_14599,N_12296);
or UO_760 (O_760,N_14782,N_13458);
or UO_761 (O_761,N_12676,N_13570);
nand UO_762 (O_762,N_13884,N_14597);
nor UO_763 (O_763,N_12135,N_13449);
and UO_764 (O_764,N_13446,N_13813);
and UO_765 (O_765,N_13269,N_12900);
and UO_766 (O_766,N_13993,N_14933);
or UO_767 (O_767,N_13041,N_12689);
nand UO_768 (O_768,N_12222,N_12187);
nand UO_769 (O_769,N_13481,N_13858);
nor UO_770 (O_770,N_14332,N_14126);
nor UO_771 (O_771,N_13657,N_12874);
or UO_772 (O_772,N_14807,N_12882);
or UO_773 (O_773,N_13439,N_12160);
and UO_774 (O_774,N_14738,N_13988);
and UO_775 (O_775,N_13307,N_14445);
nor UO_776 (O_776,N_12349,N_13428);
and UO_777 (O_777,N_14779,N_12714);
nor UO_778 (O_778,N_12758,N_13339);
and UO_779 (O_779,N_14503,N_14810);
and UO_780 (O_780,N_12418,N_12726);
nor UO_781 (O_781,N_14323,N_12177);
or UO_782 (O_782,N_14198,N_13898);
nor UO_783 (O_783,N_12047,N_14693);
or UO_784 (O_784,N_13535,N_13705);
nor UO_785 (O_785,N_13617,N_14946);
and UO_786 (O_786,N_12621,N_12044);
or UO_787 (O_787,N_14298,N_13766);
or UO_788 (O_788,N_13177,N_13321);
nor UO_789 (O_789,N_12126,N_12941);
nand UO_790 (O_790,N_14983,N_12259);
nand UO_791 (O_791,N_14350,N_12604);
and UO_792 (O_792,N_12338,N_12594);
or UO_793 (O_793,N_14745,N_14928);
nor UO_794 (O_794,N_12462,N_13902);
or UO_795 (O_795,N_14073,N_14356);
nor UO_796 (O_796,N_13343,N_12127);
nand UO_797 (O_797,N_12040,N_13036);
nor UO_798 (O_798,N_13357,N_14301);
nor UO_799 (O_799,N_13945,N_12956);
or UO_800 (O_800,N_14927,N_14937);
or UO_801 (O_801,N_13595,N_13210);
and UO_802 (O_802,N_12972,N_12633);
and UO_803 (O_803,N_13368,N_12246);
nand UO_804 (O_804,N_13108,N_14794);
or UO_805 (O_805,N_12019,N_12384);
nor UO_806 (O_806,N_13167,N_13367);
or UO_807 (O_807,N_13331,N_12364);
nor UO_808 (O_808,N_13568,N_13669);
nand UO_809 (O_809,N_12614,N_14246);
or UO_810 (O_810,N_12024,N_14193);
nor UO_811 (O_811,N_14815,N_14763);
and UO_812 (O_812,N_12951,N_14458);
or UO_813 (O_813,N_13680,N_12794);
nor UO_814 (O_814,N_13586,N_14977);
or UO_815 (O_815,N_12965,N_12248);
and UO_816 (O_816,N_14024,N_14372);
and UO_817 (O_817,N_14050,N_14011);
or UO_818 (O_818,N_12116,N_13691);
nor UO_819 (O_819,N_13609,N_12509);
or UO_820 (O_820,N_13105,N_13376);
or UO_821 (O_821,N_12432,N_14607);
nor UO_822 (O_822,N_13774,N_12558);
or UO_823 (O_823,N_14555,N_12629);
or UO_824 (O_824,N_12531,N_14461);
nand UO_825 (O_825,N_12954,N_14538);
nand UO_826 (O_826,N_14271,N_12375);
and UO_827 (O_827,N_14061,N_13984);
and UO_828 (O_828,N_14374,N_12372);
or UO_829 (O_829,N_14595,N_12586);
or UO_830 (O_830,N_12348,N_13998);
nand UO_831 (O_831,N_13074,N_12690);
nor UO_832 (O_832,N_12164,N_14357);
nor UO_833 (O_833,N_13697,N_13741);
or UO_834 (O_834,N_12490,N_13948);
or UO_835 (O_835,N_13739,N_12654);
nand UO_836 (O_836,N_13231,N_12156);
or UO_837 (O_837,N_14217,N_13824);
nor UO_838 (O_838,N_14820,N_12326);
and UO_839 (O_839,N_14382,N_13857);
nand UO_840 (O_840,N_13762,N_13822);
or UO_841 (O_841,N_12088,N_14398);
or UO_842 (O_842,N_13616,N_13341);
nand UO_843 (O_843,N_13540,N_12463);
and UO_844 (O_844,N_12903,N_14972);
or UO_845 (O_845,N_12487,N_13240);
nand UO_846 (O_846,N_14177,N_12723);
and UO_847 (O_847,N_14141,N_13821);
or UO_848 (O_848,N_12228,N_12884);
nor UO_849 (O_849,N_13718,N_14741);
nor UO_850 (O_850,N_13756,N_14376);
nor UO_851 (O_851,N_14351,N_13335);
and UO_852 (O_852,N_12751,N_13392);
nor UO_853 (O_853,N_14802,N_13328);
and UO_854 (O_854,N_14038,N_13939);
or UO_855 (O_855,N_12575,N_13109);
xor UO_856 (O_856,N_13754,N_12844);
or UO_857 (O_857,N_13096,N_13596);
and UO_858 (O_858,N_13947,N_14149);
or UO_859 (O_859,N_13719,N_14718);
or UO_860 (O_860,N_12729,N_14025);
nor UO_861 (O_861,N_13302,N_14867);
xor UO_862 (O_862,N_13017,N_13807);
nand UO_863 (O_863,N_12824,N_14925);
nand UO_864 (O_864,N_12381,N_14873);
nor UO_865 (O_865,N_14836,N_14005);
or UO_866 (O_866,N_14915,N_12351);
or UO_867 (O_867,N_13760,N_13922);
nor UO_868 (O_868,N_13623,N_12891);
nor UO_869 (O_869,N_12658,N_13737);
or UO_870 (O_870,N_12121,N_13803);
and UO_871 (O_871,N_14077,N_13801);
or UO_872 (O_872,N_14414,N_13607);
nand UO_873 (O_873,N_14362,N_14813);
nor UO_874 (O_874,N_14833,N_14954);
or UO_875 (O_875,N_13909,N_14830);
nand UO_876 (O_876,N_14797,N_14079);
or UO_877 (O_877,N_13024,N_12501);
nor UO_878 (O_878,N_13363,N_12376);
nor UO_879 (O_879,N_12732,N_13787);
or UO_880 (O_880,N_14225,N_14665);
or UO_881 (O_881,N_14154,N_12897);
nand UO_882 (O_882,N_13001,N_14474);
nor UO_883 (O_883,N_12792,N_12789);
and UO_884 (O_884,N_13610,N_13693);
nor UO_885 (O_885,N_12877,N_12429);
and UO_886 (O_886,N_12447,N_12352);
nand UO_887 (O_887,N_12795,N_12262);
nor UO_888 (O_888,N_13485,N_14365);
nand UO_889 (O_889,N_13633,N_12793);
and UO_890 (O_890,N_14072,N_12511);
nor UO_891 (O_891,N_13019,N_12183);
or UO_892 (O_892,N_12108,N_12524);
nand UO_893 (O_893,N_14986,N_14328);
nand UO_894 (O_894,N_14990,N_12512);
nand UO_895 (O_895,N_14905,N_13208);
and UO_896 (O_896,N_14008,N_14601);
nor UO_897 (O_897,N_12289,N_13310);
nor UO_898 (O_898,N_12684,N_14759);
or UO_899 (O_899,N_13189,N_14144);
nor UO_900 (O_900,N_12057,N_14758);
nand UO_901 (O_901,N_13929,N_13388);
nand UO_902 (O_902,N_14452,N_14157);
nand UO_903 (O_903,N_12090,N_13733);
or UO_904 (O_904,N_12762,N_13885);
or UO_905 (O_905,N_12322,N_14275);
and UO_906 (O_906,N_14299,N_14709);
nor UO_907 (O_907,N_14152,N_14296);
nor UO_908 (O_908,N_13046,N_13202);
nor UO_909 (O_909,N_14610,N_12323);
nand UO_910 (O_910,N_12224,N_14051);
nor UO_911 (O_911,N_13891,N_12015);
or UO_912 (O_912,N_14027,N_12544);
nor UO_913 (O_913,N_13904,N_12371);
or UO_914 (O_914,N_13867,N_14683);
or UO_915 (O_915,N_14966,N_14723);
or UO_916 (O_916,N_13391,N_13258);
and UO_917 (O_917,N_12838,N_14778);
or UO_918 (O_918,N_14109,N_12731);
or UO_919 (O_919,N_13457,N_12907);
nand UO_920 (O_920,N_12526,N_14855);
nand UO_921 (O_921,N_13452,N_13241);
and UO_922 (O_922,N_12054,N_14103);
or UO_923 (O_923,N_12873,N_14389);
or UO_924 (O_924,N_14261,N_12035);
nor UO_925 (O_925,N_12128,N_12649);
or UO_926 (O_926,N_14756,N_14146);
and UO_927 (O_927,N_13246,N_14394);
or UO_928 (O_928,N_12841,N_12875);
nand UO_929 (O_929,N_13364,N_14070);
nor UO_930 (O_930,N_12498,N_13928);
or UO_931 (O_931,N_12869,N_12962);
and UO_932 (O_932,N_14432,N_12060);
nand UO_933 (O_933,N_12945,N_14478);
nor UO_934 (O_934,N_13567,N_14982);
and UO_935 (O_935,N_14612,N_12918);
nor UO_936 (O_936,N_12079,N_14280);
nor UO_937 (O_937,N_13798,N_13423);
or UO_938 (O_938,N_13476,N_12388);
and UO_939 (O_939,N_13274,N_14364);
or UO_940 (O_940,N_13703,N_14448);
nor UO_941 (O_941,N_12776,N_12709);
or UO_942 (O_942,N_13589,N_13002);
nand UO_943 (O_943,N_12923,N_14605);
or UO_944 (O_944,N_12948,N_13999);
or UO_945 (O_945,N_12417,N_13547);
nor UO_946 (O_946,N_12333,N_13720);
nand UO_947 (O_947,N_14896,N_13372);
and UO_948 (O_948,N_13686,N_14120);
and UO_949 (O_949,N_13860,N_14462);
and UO_950 (O_950,N_12313,N_13217);
nor UO_951 (O_951,N_12804,N_14517);
or UO_952 (O_952,N_12279,N_12680);
nor UO_953 (O_953,N_14147,N_13063);
or UO_954 (O_954,N_12803,N_12217);
nor UO_955 (O_955,N_13647,N_14621);
nand UO_956 (O_956,N_12994,N_12674);
nor UO_957 (O_957,N_13441,N_14018);
or UO_958 (O_958,N_13534,N_14702);
nand UO_959 (O_959,N_13018,N_13706);
or UO_960 (O_960,N_13634,N_14850);
nor UO_961 (O_961,N_13422,N_12049);
nand UO_962 (O_962,N_12395,N_14849);
nand UO_963 (O_963,N_12562,N_14159);
xnor UO_964 (O_964,N_12659,N_14131);
or UO_965 (O_965,N_14278,N_14233);
or UO_966 (O_966,N_14347,N_12788);
nand UO_967 (O_967,N_12165,N_12870);
nor UO_968 (O_968,N_14951,N_12413);
and UO_969 (O_969,N_12608,N_12184);
nand UO_970 (O_970,N_12693,N_12098);
nand UO_971 (O_971,N_12046,N_13689);
and UO_972 (O_972,N_14856,N_13582);
nand UO_973 (O_973,N_12115,N_14846);
and UO_974 (O_974,N_12510,N_13051);
or UO_975 (O_975,N_13152,N_13931);
nand UO_976 (O_976,N_14684,N_14191);
nor UO_977 (O_977,N_14269,N_12025);
and UO_978 (O_978,N_14716,N_14646);
nor UO_979 (O_979,N_14679,N_13101);
or UO_980 (O_980,N_14477,N_12747);
nand UO_981 (O_981,N_13360,N_12677);
nor UO_982 (O_982,N_13699,N_12355);
nor UO_983 (O_983,N_12996,N_14331);
and UO_984 (O_984,N_14963,N_13529);
nand UO_985 (O_985,N_13553,N_13243);
and UO_986 (O_986,N_13066,N_14917);
and UO_987 (O_987,N_14609,N_14400);
nor UO_988 (O_988,N_12226,N_14140);
or UO_989 (O_989,N_12342,N_12131);
nor UO_990 (O_990,N_14529,N_13426);
nor UO_991 (O_991,N_13434,N_14101);
and UO_992 (O_992,N_12744,N_14297);
nand UO_993 (O_993,N_13228,N_13378);
nor UO_994 (O_994,N_12081,N_14627);
and UO_995 (O_995,N_13248,N_13580);
nand UO_996 (O_996,N_12568,N_12706);
nor UO_997 (O_997,N_12549,N_12004);
nor UO_998 (O_998,N_14343,N_13472);
or UO_999 (O_999,N_14424,N_12821);
and UO_1000 (O_1000,N_12831,N_12955);
and UO_1001 (O_1001,N_12998,N_12861);
and UO_1002 (O_1002,N_14828,N_13415);
or UO_1003 (O_1003,N_12635,N_12642);
and UO_1004 (O_1004,N_14703,N_14353);
and UO_1005 (O_1005,N_12999,N_12939);
nand UO_1006 (O_1006,N_14994,N_14349);
or UO_1007 (O_1007,N_14532,N_13355);
and UO_1008 (O_1008,N_14482,N_13348);
and UO_1009 (O_1009,N_12506,N_12696);
and UO_1010 (O_1010,N_12743,N_14918);
nand UO_1011 (O_1011,N_12150,N_14519);
nand UO_1012 (O_1012,N_12146,N_13788);
nor UO_1013 (O_1013,N_14578,N_12565);
or UO_1014 (O_1014,N_14426,N_12627);
or UO_1015 (O_1015,N_14370,N_14438);
and UO_1016 (O_1016,N_12016,N_14697);
nand UO_1017 (O_1017,N_13416,N_14871);
nand UO_1018 (O_1018,N_12700,N_14757);
nand UO_1019 (O_1019,N_14235,N_12014);
or UO_1020 (O_1020,N_13340,N_13921);
and UO_1021 (O_1021,N_13954,N_13957);
or UO_1022 (O_1022,N_13655,N_14858);
and UO_1023 (O_1023,N_12270,N_12157);
nor UO_1024 (O_1024,N_14806,N_14724);
nor UO_1025 (O_1025,N_12410,N_12966);
nand UO_1026 (O_1026,N_14603,N_12457);
and UO_1027 (O_1027,N_14333,N_13574);
and UO_1028 (O_1028,N_12210,N_14930);
nor UO_1029 (O_1029,N_12369,N_14207);
nor UO_1030 (O_1030,N_13775,N_12515);
and UO_1031 (O_1031,N_14670,N_12481);
nor UO_1032 (O_1032,N_14023,N_12707);
nand UO_1033 (O_1033,N_12169,N_14110);
nor UO_1034 (O_1034,N_12980,N_13296);
nand UO_1035 (O_1035,N_14685,N_13374);
or UO_1036 (O_1036,N_12768,N_13603);
xnor UO_1037 (O_1037,N_12101,N_14232);
and UO_1038 (O_1038,N_13169,N_13661);
nor UO_1039 (O_1039,N_12547,N_13078);
nand UO_1040 (O_1040,N_13895,N_13155);
nor UO_1041 (O_1041,N_12437,N_13866);
nor UO_1042 (O_1042,N_12784,N_13587);
nor UO_1043 (O_1043,N_14310,N_13317);
and UO_1044 (O_1044,N_13408,N_13354);
and UO_1045 (O_1045,N_13178,N_13032);
nand UO_1046 (O_1046,N_12483,N_13664);
nor UO_1047 (O_1047,N_13251,N_12971);
and UO_1048 (O_1048,N_12404,N_13295);
nand UO_1049 (O_1049,N_13114,N_13027);
or UO_1050 (O_1050,N_14355,N_13039);
nand UO_1051 (O_1051,N_14255,N_13081);
and UO_1052 (O_1052,N_13403,N_13841);
and UO_1053 (O_1053,N_14399,N_12252);
nand UO_1054 (O_1054,N_13738,N_13656);
or UO_1055 (O_1055,N_13962,N_12303);
nand UO_1056 (O_1056,N_13732,N_12399);
nor UO_1057 (O_1057,N_13702,N_12885);
or UO_1058 (O_1058,N_14655,N_13727);
or UO_1059 (O_1059,N_14097,N_12769);
xor UO_1060 (O_1060,N_13466,N_14527);
nor UO_1061 (O_1061,N_13012,N_14640);
nand UO_1062 (O_1062,N_14442,N_13526);
and UO_1063 (O_1063,N_14957,N_13033);
and UO_1064 (O_1064,N_14556,N_14969);
and UO_1065 (O_1065,N_12712,N_14219);
nand UO_1066 (O_1066,N_12470,N_13783);
or UO_1067 (O_1067,N_13855,N_14668);
nor UO_1068 (O_1068,N_12761,N_13588);
or UO_1069 (O_1069,N_12973,N_12321);
nor UO_1070 (O_1070,N_13492,N_14751);
nand UO_1071 (O_1071,N_12400,N_14618);
and UO_1072 (O_1072,N_14052,N_14638);
nand UO_1073 (O_1073,N_14066,N_14984);
and UO_1074 (O_1074,N_12110,N_13627);
nor UO_1075 (O_1075,N_12356,N_14063);
nor UO_1076 (O_1076,N_13079,N_12085);
nand UO_1077 (O_1077,N_13930,N_13005);
and UO_1078 (O_1078,N_13207,N_12330);
nor UO_1079 (O_1079,N_13454,N_12107);
and UO_1080 (O_1080,N_14487,N_12011);
and UO_1081 (O_1081,N_13548,N_12738);
or UO_1082 (O_1082,N_14208,N_14539);
nand UO_1083 (O_1083,N_14885,N_13117);
or UO_1084 (O_1084,N_14393,N_12158);
or UO_1085 (O_1085,N_12319,N_12715);
nand UO_1086 (O_1086,N_12806,N_12022);
nor UO_1087 (O_1087,N_13220,N_12832);
and UO_1088 (O_1088,N_12963,N_14704);
and UO_1089 (O_1089,N_14899,N_12166);
and UO_1090 (O_1090,N_12474,N_13206);
nor UO_1091 (O_1091,N_14282,N_12767);
and UO_1092 (O_1092,N_13606,N_14472);
nor UO_1093 (O_1093,N_14369,N_13242);
or UO_1094 (O_1094,N_13653,N_12823);
or UO_1095 (O_1095,N_12281,N_12021);
nor UO_1096 (O_1096,N_12265,N_12059);
and UO_1097 (O_1097,N_12710,N_14182);
nor UO_1098 (O_1098,N_13157,N_13057);
and UO_1099 (O_1099,N_12191,N_13642);
nand UO_1100 (O_1100,N_13211,N_12328);
or UO_1101 (O_1101,N_13255,N_12995);
or UO_1102 (O_1102,N_14682,N_13579);
or UO_1103 (O_1103,N_14891,N_14767);
xor UO_1104 (O_1104,N_13159,N_12964);
and UO_1105 (O_1105,N_12122,N_13337);
nor UO_1106 (O_1106,N_13846,N_12444);
nor UO_1107 (O_1107,N_14094,N_14315);
nand UO_1108 (O_1108,N_13809,N_13832);
nor UO_1109 (O_1109,N_12862,N_12818);
nor UO_1110 (O_1110,N_14606,N_12622);
nand UO_1111 (O_1111,N_14428,N_12170);
and UO_1112 (O_1112,N_13652,N_12837);
or UO_1113 (O_1113,N_12719,N_12105);
nor UO_1114 (O_1114,N_12275,N_13828);
or UO_1115 (O_1115,N_13134,N_14239);
nor UO_1116 (O_1116,N_14894,N_14953);
or UO_1117 (O_1117,N_13462,N_13638);
or UO_1118 (O_1118,N_12589,N_14634);
and UO_1119 (O_1119,N_12208,N_12566);
and UO_1120 (O_1120,N_13620,N_12179);
nand UO_1121 (O_1121,N_13427,N_13777);
or UO_1122 (O_1122,N_12419,N_13637);
and UO_1123 (O_1123,N_14242,N_13864);
nor UO_1124 (O_1124,N_12247,N_13990);
nor UO_1125 (O_1125,N_12603,N_12138);
or UO_1126 (O_1126,N_13199,N_14971);
nand UO_1127 (O_1127,N_13470,N_12876);
nor UO_1128 (O_1128,N_13067,N_14001);
and UO_1129 (O_1129,N_13129,N_12630);
or UO_1130 (O_1130,N_13273,N_12456);
and UO_1131 (O_1131,N_14663,N_13075);
or UO_1132 (O_1132,N_13748,N_14010);
nand UO_1133 (O_1133,N_12039,N_12638);
and UO_1134 (O_1134,N_13506,N_12898);
nor UO_1135 (O_1135,N_12112,N_14215);
and UO_1136 (O_1136,N_13953,N_14696);
nor UO_1137 (O_1137,N_13181,N_12001);
and UO_1138 (O_1138,N_12981,N_14934);
nand UO_1139 (O_1139,N_14484,N_12573);
nand UO_1140 (O_1140,N_14932,N_13500);
or UO_1141 (O_1141,N_13913,N_14631);
and UO_1142 (O_1142,N_14111,N_13602);
nand UO_1143 (O_1143,N_14325,N_13973);
nand UO_1144 (O_1144,N_14768,N_12017);
nor UO_1145 (O_1145,N_13316,N_12592);
nor UO_1146 (O_1146,N_12620,N_12826);
and UO_1147 (O_1147,N_12070,N_14862);
or UO_1148 (O_1148,N_14636,N_14209);
or UO_1149 (O_1149,N_12251,N_12892);
nand UO_1150 (O_1150,N_12233,N_12256);
nor UO_1151 (O_1151,N_13298,N_13944);
or UO_1152 (O_1152,N_12660,N_14238);
and UO_1153 (O_1153,N_13575,N_14711);
or UO_1154 (O_1154,N_13059,N_14447);
nor UO_1155 (O_1155,N_12385,N_12489);
nor UO_1156 (O_1156,N_14795,N_12935);
nand UO_1157 (O_1157,N_13050,N_14016);
nor UO_1158 (O_1158,N_13996,N_12943);
and UO_1159 (O_1159,N_14594,N_13510);
and UO_1160 (O_1160,N_13267,N_13784);
nand UO_1161 (O_1161,N_13136,N_14049);
or UO_1162 (O_1162,N_13257,N_12302);
or UO_1163 (O_1163,N_14468,N_13522);
or UO_1164 (O_1164,N_14180,N_13235);
nand UO_1165 (O_1165,N_13153,N_13148);
or UO_1166 (O_1166,N_14065,N_13095);
nand UO_1167 (O_1167,N_14908,N_12209);
nand UO_1168 (O_1168,N_13881,N_14596);
and UO_1169 (O_1169,N_14172,N_13796);
and UO_1170 (O_1170,N_12149,N_13831);
nand UO_1171 (O_1171,N_13016,N_13892);
nor UO_1172 (O_1172,N_13176,N_12174);
nand UO_1173 (O_1173,N_12097,N_12518);
nand UO_1174 (O_1174,N_13491,N_13030);
nor UO_1175 (O_1175,N_13073,N_14135);
or UO_1176 (O_1176,N_14042,N_14339);
nor UO_1177 (O_1177,N_14546,N_13605);
nand UO_1178 (O_1178,N_14178,N_14998);
nand UO_1179 (O_1179,N_13144,N_14501);
nand UO_1180 (O_1180,N_13342,N_13398);
nand UO_1181 (O_1181,N_13072,N_13180);
and UO_1182 (O_1182,N_13667,N_14181);
or UO_1183 (O_1183,N_13284,N_14818);
or UO_1184 (O_1184,N_14980,N_14913);
nand UO_1185 (O_1185,N_12361,N_12433);
and UO_1186 (O_1186,N_14916,N_13629);
nor UO_1187 (O_1187,N_13028,N_14658);
nand UO_1188 (O_1188,N_12938,N_12859);
and UO_1189 (O_1189,N_14281,N_13459);
or UO_1190 (O_1190,N_13519,N_13338);
nand UO_1191 (O_1191,N_12394,N_14340);
nand UO_1192 (O_1192,N_13226,N_14893);
or UO_1193 (O_1193,N_12293,N_12334);
or UO_1194 (O_1194,N_12239,N_14470);
nand UO_1195 (O_1195,N_13239,N_14637);
nor UO_1196 (O_1196,N_14245,N_14526);
nand UO_1197 (O_1197,N_13782,N_14268);
nand UO_1198 (O_1198,N_12694,N_13044);
or UO_1199 (O_1199,N_13448,N_13933);
nand UO_1200 (O_1200,N_13107,N_13571);
or UO_1201 (O_1201,N_13676,N_14270);
nor UO_1202 (O_1202,N_13380,N_12591);
nand UO_1203 (O_1203,N_14046,N_13614);
or UO_1204 (O_1204,N_13597,N_12672);
or UO_1205 (O_1205,N_14744,N_14765);
nand UO_1206 (O_1206,N_13127,N_14204);
nand UO_1207 (O_1207,N_12286,N_14720);
and UO_1208 (O_1208,N_12650,N_14499);
or UO_1209 (O_1209,N_13961,N_14218);
or UO_1210 (O_1210,N_12993,N_13968);
and UO_1211 (O_1211,N_13418,N_14420);
or UO_1212 (O_1212,N_13088,N_12716);
nand UO_1213 (O_1213,N_13326,N_12815);
or UO_1214 (O_1214,N_13600,N_14401);
and UO_1215 (O_1215,N_13272,N_12847);
and UO_1216 (O_1216,N_13905,N_12742);
and UO_1217 (O_1217,N_12280,N_14821);
nor UO_1218 (O_1218,N_14864,N_12271);
nand UO_1219 (O_1219,N_13116,N_12836);
and UO_1220 (O_1220,N_14590,N_14371);
nand UO_1221 (O_1221,N_13820,N_12894);
or UO_1222 (O_1222,N_13672,N_12297);
and UO_1223 (O_1223,N_12887,N_14902);
nand UO_1224 (O_1224,N_13146,N_13203);
or UO_1225 (O_1225,N_13477,N_13256);
and UO_1226 (O_1226,N_13443,N_13118);
and UO_1227 (O_1227,N_14287,N_14082);
nor UO_1228 (O_1228,N_13825,N_12863);
or UO_1229 (O_1229,N_13162,N_14174);
nor UO_1230 (O_1230,N_13244,N_13010);
or UO_1231 (O_1231,N_12472,N_14244);
nand UO_1232 (O_1232,N_12724,N_13332);
nor UO_1233 (O_1233,N_14650,N_12243);
or UO_1234 (O_1234,N_13934,N_13972);
or UO_1235 (O_1235,N_13430,N_13325);
nand UO_1236 (O_1236,N_14203,N_12027);
and UO_1237 (O_1237,N_13795,N_12800);
nand UO_1238 (O_1238,N_14635,N_12904);
or UO_1239 (O_1239,N_12484,N_12631);
or UO_1240 (O_1240,N_14291,N_14033);
or UO_1241 (O_1241,N_12378,N_13171);
nor UO_1242 (O_1242,N_12968,N_12114);
or UO_1243 (O_1243,N_14575,N_12006);
nor UO_1244 (O_1244,N_13465,N_13658);
or UO_1245 (O_1245,N_14007,N_13869);
nor UO_1246 (O_1246,N_13527,N_14829);
or UO_1247 (O_1247,N_13815,N_12193);
and UO_1248 (O_1248,N_13590,N_13473);
and UO_1249 (O_1249,N_14476,N_14320);
or UO_1250 (O_1250,N_13405,N_12668);
nor UO_1251 (O_1251,N_12616,N_12100);
and UO_1252 (O_1252,N_12685,N_14611);
or UO_1253 (O_1253,N_14911,N_14227);
and UO_1254 (O_1254,N_13336,N_13946);
nor UO_1255 (O_1255,N_12819,N_14200);
or UO_1256 (O_1256,N_14375,N_13104);
or UO_1257 (O_1257,N_14205,N_14585);
and UO_1258 (O_1258,N_13076,N_12852);
or UO_1259 (O_1259,N_12740,N_13899);
or UO_1260 (O_1260,N_14559,N_13794);
nor UO_1261 (O_1261,N_12151,N_14321);
or UO_1262 (O_1262,N_13843,N_12362);
and UO_1263 (O_1263,N_12940,N_12043);
or UO_1264 (O_1264,N_14508,N_14337);
nand UO_1265 (O_1265,N_12926,N_13668);
or UO_1266 (O_1266,N_13233,N_14700);
or UO_1267 (O_1267,N_14857,N_13525);
nand UO_1268 (O_1268,N_12340,N_14987);
or UO_1269 (O_1269,N_13785,N_13917);
nor UO_1270 (O_1270,N_13037,N_12278);
and UO_1271 (O_1271,N_12077,N_12365);
nor UO_1272 (O_1272,N_14387,N_13497);
nor UO_1273 (O_1273,N_12905,N_13817);
nor UO_1274 (O_1274,N_12775,N_14475);
xor UO_1275 (O_1275,N_12588,N_14434);
or UO_1276 (O_1276,N_12782,N_14253);
nor UO_1277 (O_1277,N_12671,N_13852);
or UO_1278 (O_1278,N_12370,N_14341);
nand UO_1279 (O_1279,N_12161,N_12571);
and UO_1280 (O_1280,N_12919,N_12840);
or UO_1281 (O_1281,N_14560,N_13980);
or UO_1282 (O_1282,N_14497,N_14675);
and UO_1283 (O_1283,N_12865,N_13942);
or UO_1284 (O_1284,N_14031,N_13062);
nor UO_1285 (O_1285,N_12906,N_14561);
or UO_1286 (O_1286,N_12653,N_12008);
nor UO_1287 (O_1287,N_13926,N_14000);
nor UO_1288 (O_1288,N_12363,N_12403);
or UO_1289 (O_1289,N_12221,N_12848);
nand UO_1290 (O_1290,N_13447,N_12656);
and UO_1291 (O_1291,N_13216,N_14392);
nor UO_1292 (O_1292,N_12461,N_13431);
nor UO_1293 (O_1293,N_12153,N_13994);
nor UO_1294 (O_1294,N_13143,N_13773);
nand UO_1295 (O_1295,N_13745,N_12828);
or UO_1296 (O_1296,N_14822,N_13369);
nand UO_1297 (O_1297,N_14425,N_14789);
nor UO_1298 (O_1298,N_12306,N_12269);
or UO_1299 (O_1299,N_13260,N_12931);
and UO_1300 (O_1300,N_13115,N_12300);
and UO_1301 (O_1301,N_13440,N_13839);
and UO_1302 (O_1302,N_14294,N_12009);
nor UO_1303 (O_1303,N_14620,N_12777);
or UO_1304 (O_1304,N_12641,N_12346);
and UO_1305 (O_1305,N_12527,N_14444);
nand UO_1306 (O_1306,N_13225,N_14192);
nor UO_1307 (O_1307,N_12678,N_12167);
nor UO_1308 (O_1308,N_13488,N_13359);
or UO_1309 (O_1309,N_12813,N_13797);
or UO_1310 (O_1310,N_12148,N_14383);
or UO_1311 (O_1311,N_13621,N_14243);
or UO_1312 (O_1312,N_12772,N_13031);
nor UO_1313 (O_1313,N_14433,N_12335);
and UO_1314 (O_1314,N_13856,N_12213);
and UO_1315 (O_1315,N_13230,N_14313);
and UO_1316 (O_1316,N_12773,N_12072);
nor UO_1317 (O_1317,N_12357,N_13494);
nand UO_1318 (O_1318,N_13478,N_14513);
and UO_1319 (O_1319,N_14863,N_12471);
and UO_1320 (O_1320,N_13475,N_13805);
and UO_1321 (O_1321,N_12552,N_14843);
or UO_1322 (O_1322,N_12613,N_12382);
nand UO_1323 (O_1323,N_13312,N_14211);
nor UO_1324 (O_1324,N_14080,N_12427);
nand UO_1325 (O_1325,N_14914,N_12095);
and UO_1326 (O_1326,N_12301,N_12469);
nor UO_1327 (O_1327,N_14788,N_13389);
or UO_1328 (O_1328,N_13287,N_14032);
nand UO_1329 (O_1329,N_14148,N_14772);
nand UO_1330 (O_1330,N_12914,N_14305);
nor UO_1331 (O_1331,N_13047,N_13158);
and UO_1332 (O_1332,N_12412,N_12976);
or UO_1333 (O_1333,N_13910,N_14875);
and UO_1334 (O_1334,N_14459,N_14158);
and UO_1335 (O_1335,N_12307,N_12416);
and UO_1336 (O_1336,N_12969,N_12675);
and UO_1337 (O_1337,N_14380,N_14960);
or UO_1338 (O_1338,N_14130,N_12516);
or UO_1339 (O_1339,N_12648,N_12610);
nor UO_1340 (O_1340,N_12067,N_14421);
or UO_1341 (O_1341,N_12957,N_14961);
and UO_1342 (O_1342,N_13396,N_14892);
or UO_1343 (O_1343,N_14363,N_13663);
nand UO_1344 (O_1344,N_14803,N_14888);
or UO_1345 (O_1345,N_14195,N_13631);
and UO_1346 (O_1346,N_12495,N_13613);
nor UO_1347 (O_1347,N_14600,N_12646);
or UO_1348 (O_1348,N_13468,N_14303);
nand UO_1349 (O_1349,N_13122,N_14279);
nand UO_1350 (O_1350,N_12669,N_14163);
or UO_1351 (O_1351,N_13077,N_12946);
nor UO_1352 (O_1352,N_14197,N_13161);
nand UO_1353 (O_1353,N_14622,N_12508);
or UO_1354 (O_1354,N_13236,N_14628);
or UO_1355 (O_1355,N_12255,N_14762);
and UO_1356 (O_1356,N_14642,N_13747);
and UO_1357 (O_1357,N_13011,N_12807);
nor UO_1358 (O_1358,N_12564,N_12214);
nor UO_1359 (O_1359,N_12698,N_14985);
nor UO_1360 (O_1360,N_14119,N_13377);
nor UO_1361 (O_1361,N_13344,N_13983);
and UO_1362 (O_1362,N_12036,N_13200);
nand UO_1363 (O_1363,N_14480,N_14824);
nor UO_1364 (O_1364,N_12332,N_14592);
and UO_1365 (O_1365,N_14924,N_14694);
nand UO_1366 (O_1366,N_12503,N_12774);
or UO_1367 (O_1367,N_12569,N_12921);
nand UO_1368 (O_1368,N_14335,N_14240);
or UO_1369 (O_1369,N_14318,N_14623);
and UO_1370 (O_1370,N_13349,N_13399);
nand UO_1371 (O_1371,N_14230,N_12202);
nand UO_1372 (O_1372,N_13879,N_13139);
nor UO_1373 (O_1373,N_12928,N_12260);
and UO_1374 (O_1374,N_12580,N_12961);
nor UO_1375 (O_1375,N_12615,N_14118);
nor UO_1376 (O_1376,N_13622,N_14123);
and UO_1377 (O_1377,N_12785,N_14558);
or UO_1378 (O_1378,N_13250,N_12283);
and UO_1379 (O_1379,N_14926,N_13808);
or UO_1380 (O_1380,N_14940,N_12453);
nor UO_1381 (O_1381,N_13327,N_12423);
nor UO_1382 (O_1382,N_14213,N_13518);
nor UO_1383 (O_1383,N_13304,N_12927);
nand UO_1384 (O_1384,N_12757,N_13394);
nor UO_1385 (O_1385,N_12002,N_14690);
and UO_1386 (O_1386,N_14162,N_13908);
and UO_1387 (O_1387,N_14542,N_12431);
or UO_1388 (O_1388,N_12023,N_12666);
or UO_1389 (O_1389,N_13170,N_14186);
or UO_1390 (O_1390,N_14378,N_12176);
and UO_1391 (O_1391,N_12599,N_13924);
and UO_1392 (O_1392,N_12607,N_14876);
or UO_1393 (O_1393,N_14022,N_14988);
nand UO_1394 (O_1394,N_13682,N_13214);
and UO_1395 (O_1395,N_13043,N_12853);
or UO_1396 (O_1396,N_13673,N_12663);
nand UO_1397 (O_1397,N_12559,N_12087);
and UO_1398 (O_1398,N_13728,N_12582);
nand UO_1399 (O_1399,N_14869,N_13868);
and UO_1400 (O_1400,N_13508,N_14456);
and UO_1401 (O_1401,N_14210,N_14283);
and UO_1402 (O_1402,N_12778,N_13871);
or UO_1403 (O_1403,N_12843,N_14563);
nor UO_1404 (O_1404,N_12532,N_14004);
or UO_1405 (O_1405,N_12073,N_12013);
or UO_1406 (O_1406,N_14936,N_13172);
nand UO_1407 (O_1407,N_13612,N_14485);
and UO_1408 (O_1408,N_12366,N_12266);
nand UO_1409 (O_1409,N_13935,N_13511);
or UO_1410 (O_1410,N_13896,N_14236);
nor UO_1411 (O_1411,N_14889,N_14473);
or UO_1412 (O_1412,N_13849,N_13823);
nor UO_1413 (O_1413,N_12467,N_14883);
nand UO_1414 (O_1414,N_12312,N_14088);
nand UO_1415 (O_1415,N_13767,N_14206);
or UO_1416 (O_1416,N_14469,N_13182);
and UO_1417 (O_1417,N_12581,N_12258);
or UO_1418 (O_1418,N_14440,N_12198);
nand UO_1419 (O_1419,N_13461,N_12866);
or UO_1420 (O_1420,N_14412,N_14929);
nor UO_1421 (O_1421,N_14096,N_14348);
nand UO_1422 (O_1422,N_12428,N_12651);
and UO_1423 (O_1423,N_12727,N_14167);
nand UO_1424 (O_1424,N_12065,N_12442);
nand UO_1425 (O_1425,N_13436,N_14737);
or UO_1426 (O_1426,N_13370,N_13087);
or UO_1427 (O_1427,N_14098,N_12703);
or UO_1428 (O_1428,N_14792,N_14630);
nand UO_1429 (O_1429,N_13098,N_13541);
xor UO_1430 (O_1430,N_13276,N_14416);
nand UO_1431 (O_1431,N_13205,N_13347);
nor UO_1432 (O_1432,N_12746,N_14550);
or UO_1433 (O_1433,N_12978,N_12205);
or UO_1434 (O_1434,N_12872,N_13303);
nor UO_1435 (O_1435,N_13126,N_12475);
and UO_1436 (O_1436,N_13319,N_13765);
nor UO_1437 (O_1437,N_13080,N_14992);
nor UO_1438 (O_1438,N_12446,N_13790);
nor UO_1439 (O_1439,N_13859,N_13981);
nand UO_1440 (O_1440,N_14965,N_14076);
or UO_1441 (O_1441,N_14727,N_14457);
and UO_1442 (O_1442,N_12443,N_12078);
or UO_1443 (O_1443,N_14408,N_12682);
nor UO_1444 (O_1444,N_12314,N_14021);
and UO_1445 (O_1445,N_12713,N_14386);
nor UO_1446 (O_1446,N_14626,N_14823);
nor UO_1447 (O_1447,N_12879,N_13419);
nor UO_1448 (O_1448,N_14036,N_14999);
nand UO_1449 (O_1449,N_13025,N_14676);
and UO_1450 (O_1450,N_12505,N_13630);
or UO_1451 (O_1451,N_12878,N_13309);
or UO_1452 (O_1452,N_14729,N_12204);
nand UO_1453 (O_1453,N_14991,N_12038);
nor UO_1454 (O_1454,N_14587,N_13034);
nand UO_1455 (O_1455,N_13641,N_12567);
nand UO_1456 (O_1456,N_12113,N_14506);
nand UO_1457 (O_1457,N_12756,N_14948);
nand UO_1458 (O_1458,N_14417,N_13712);
and UO_1459 (O_1459,N_13549,N_13577);
nand UO_1460 (O_1460,N_14142,N_13184);
nand UO_1461 (O_1461,N_14311,N_14567);
nand UO_1462 (O_1462,N_14942,N_12514);
nand UO_1463 (O_1463,N_13836,N_13971);
nand UO_1464 (O_1464,N_14898,N_14489);
or UO_1465 (O_1465,N_13297,N_12494);
xnor UO_1466 (O_1466,N_14950,N_14285);
nand UO_1467 (O_1467,N_14671,N_13520);
nand UO_1468 (O_1468,N_13315,N_12640);
nor UO_1469 (O_1469,N_14368,N_13395);
or UO_1470 (O_1470,N_13769,N_14359);
and UO_1471 (O_1471,N_12329,N_13193);
nand UO_1472 (O_1472,N_14057,N_12317);
and UO_1473 (O_1473,N_13514,N_14220);
and UO_1474 (O_1474,N_13420,N_14838);
nor UO_1475 (O_1475,N_12436,N_13070);
nor UO_1476 (O_1476,N_14512,N_14231);
or UO_1477 (O_1477,N_13925,N_13837);
nand UO_1478 (O_1478,N_14734,N_13991);
and UO_1479 (O_1479,N_12287,N_14586);
and UO_1480 (O_1480,N_12479,N_13542);
nand UO_1481 (O_1481,N_14554,N_13489);
or UO_1482 (O_1482,N_14840,N_13894);
nor UO_1483 (O_1483,N_14504,N_12010);
nor UO_1484 (O_1484,N_13644,N_14643);
nand UO_1485 (O_1485,N_14787,N_14537);
nor UO_1486 (O_1486,N_14284,N_14674);
nand UO_1487 (O_1487,N_14415,N_14074);
or UO_1488 (O_1488,N_14326,N_14591);
and UO_1489 (O_1489,N_12175,N_12096);
nand UO_1490 (O_1490,N_14653,N_14692);
nand UO_1491 (O_1491,N_14544,N_12695);
nor UO_1492 (O_1492,N_14184,N_12949);
nor UO_1493 (O_1493,N_13906,N_13731);
nand UO_1494 (O_1494,N_12858,N_12132);
nand UO_1495 (O_1495,N_13724,N_14887);
nor UO_1496 (O_1496,N_12000,N_12864);
nand UO_1497 (O_1497,N_13229,N_12725);
and UO_1498 (O_1498,N_12347,N_14344);
or UO_1499 (O_1499,N_13504,N_14431);
and UO_1500 (O_1500,N_12884,N_13203);
nor UO_1501 (O_1501,N_14612,N_13467);
or UO_1502 (O_1502,N_14213,N_14858);
nor UO_1503 (O_1503,N_12710,N_14871);
nor UO_1504 (O_1504,N_13442,N_12461);
or UO_1505 (O_1505,N_12160,N_13388);
or UO_1506 (O_1506,N_12020,N_13123);
nor UO_1507 (O_1507,N_12318,N_13988);
nand UO_1508 (O_1508,N_12066,N_12143);
nand UO_1509 (O_1509,N_14553,N_13899);
nor UO_1510 (O_1510,N_12503,N_14332);
nor UO_1511 (O_1511,N_12139,N_13859);
nor UO_1512 (O_1512,N_12624,N_14928);
and UO_1513 (O_1513,N_14782,N_12597);
nor UO_1514 (O_1514,N_14376,N_13772);
xor UO_1515 (O_1515,N_14351,N_13453);
nand UO_1516 (O_1516,N_14032,N_14616);
and UO_1517 (O_1517,N_12263,N_14017);
or UO_1518 (O_1518,N_12783,N_13586);
or UO_1519 (O_1519,N_12807,N_12046);
nand UO_1520 (O_1520,N_12017,N_12753);
nand UO_1521 (O_1521,N_14978,N_13683);
or UO_1522 (O_1522,N_14990,N_12355);
nand UO_1523 (O_1523,N_13507,N_12425);
nand UO_1524 (O_1524,N_14480,N_13412);
or UO_1525 (O_1525,N_13119,N_13921);
nor UO_1526 (O_1526,N_12178,N_13031);
or UO_1527 (O_1527,N_14354,N_14523);
or UO_1528 (O_1528,N_13280,N_12733);
nor UO_1529 (O_1529,N_14766,N_12226);
and UO_1530 (O_1530,N_12309,N_14616);
or UO_1531 (O_1531,N_12046,N_14185);
nor UO_1532 (O_1532,N_13186,N_14756);
nor UO_1533 (O_1533,N_12006,N_12902);
and UO_1534 (O_1534,N_12500,N_14605);
nand UO_1535 (O_1535,N_12395,N_13012);
and UO_1536 (O_1536,N_12032,N_14564);
or UO_1537 (O_1537,N_14554,N_12074);
or UO_1538 (O_1538,N_14876,N_12960);
nand UO_1539 (O_1539,N_13038,N_13101);
or UO_1540 (O_1540,N_13917,N_13787);
nand UO_1541 (O_1541,N_12808,N_12893);
and UO_1542 (O_1542,N_14427,N_12929);
and UO_1543 (O_1543,N_13951,N_14855);
or UO_1544 (O_1544,N_14169,N_13904);
xnor UO_1545 (O_1545,N_12493,N_13038);
or UO_1546 (O_1546,N_12537,N_12206);
and UO_1547 (O_1547,N_12054,N_12951);
or UO_1548 (O_1548,N_13183,N_13128);
and UO_1549 (O_1549,N_13993,N_12824);
nand UO_1550 (O_1550,N_13038,N_14711);
nand UO_1551 (O_1551,N_14888,N_14554);
or UO_1552 (O_1552,N_13557,N_12069);
or UO_1553 (O_1553,N_14372,N_13439);
nor UO_1554 (O_1554,N_13819,N_13958);
or UO_1555 (O_1555,N_13949,N_14590);
nor UO_1556 (O_1556,N_12821,N_14747);
or UO_1557 (O_1557,N_14729,N_12334);
or UO_1558 (O_1558,N_12321,N_14213);
or UO_1559 (O_1559,N_13827,N_12564);
nand UO_1560 (O_1560,N_12382,N_13239);
and UO_1561 (O_1561,N_14504,N_12316);
or UO_1562 (O_1562,N_13041,N_13396);
nand UO_1563 (O_1563,N_14531,N_14390);
and UO_1564 (O_1564,N_12670,N_13123);
and UO_1565 (O_1565,N_12899,N_13493);
nand UO_1566 (O_1566,N_13315,N_14582);
nand UO_1567 (O_1567,N_12734,N_13292);
nor UO_1568 (O_1568,N_12089,N_12235);
nor UO_1569 (O_1569,N_13208,N_12946);
and UO_1570 (O_1570,N_12617,N_13477);
nor UO_1571 (O_1571,N_12201,N_13768);
and UO_1572 (O_1572,N_12896,N_13848);
xnor UO_1573 (O_1573,N_14260,N_14767);
and UO_1574 (O_1574,N_12335,N_13749);
nor UO_1575 (O_1575,N_12310,N_12911);
nor UO_1576 (O_1576,N_12243,N_14291);
nor UO_1577 (O_1577,N_12324,N_14944);
or UO_1578 (O_1578,N_13194,N_14581);
nor UO_1579 (O_1579,N_12028,N_14681);
or UO_1580 (O_1580,N_14912,N_14579);
and UO_1581 (O_1581,N_12210,N_12466);
and UO_1582 (O_1582,N_13724,N_12556);
nor UO_1583 (O_1583,N_12403,N_13924);
or UO_1584 (O_1584,N_14196,N_12250);
nand UO_1585 (O_1585,N_13724,N_12079);
and UO_1586 (O_1586,N_13935,N_13221);
or UO_1587 (O_1587,N_12839,N_14593);
and UO_1588 (O_1588,N_14681,N_12624);
nand UO_1589 (O_1589,N_13470,N_12540);
nand UO_1590 (O_1590,N_12385,N_14126);
nand UO_1591 (O_1591,N_13642,N_12916);
nand UO_1592 (O_1592,N_12757,N_13386);
and UO_1593 (O_1593,N_12405,N_13841);
and UO_1594 (O_1594,N_12411,N_14346);
nand UO_1595 (O_1595,N_14569,N_14241);
xor UO_1596 (O_1596,N_13904,N_13712);
and UO_1597 (O_1597,N_12243,N_14086);
or UO_1598 (O_1598,N_13285,N_14519);
nand UO_1599 (O_1599,N_13284,N_14837);
nor UO_1600 (O_1600,N_12376,N_12285);
or UO_1601 (O_1601,N_12391,N_13105);
and UO_1602 (O_1602,N_12545,N_14828);
nand UO_1603 (O_1603,N_13474,N_13149);
nand UO_1604 (O_1604,N_12715,N_14729);
or UO_1605 (O_1605,N_14562,N_13733);
xnor UO_1606 (O_1606,N_12776,N_13721);
and UO_1607 (O_1607,N_14756,N_14261);
or UO_1608 (O_1608,N_12536,N_14449);
nand UO_1609 (O_1609,N_14662,N_14916);
and UO_1610 (O_1610,N_12377,N_14464);
and UO_1611 (O_1611,N_12648,N_14926);
nand UO_1612 (O_1612,N_13194,N_13956);
or UO_1613 (O_1613,N_13426,N_12705);
and UO_1614 (O_1614,N_14646,N_14117);
and UO_1615 (O_1615,N_13019,N_12596);
nor UO_1616 (O_1616,N_14979,N_13901);
nand UO_1617 (O_1617,N_14469,N_14977);
and UO_1618 (O_1618,N_13687,N_14530);
nor UO_1619 (O_1619,N_14580,N_12225);
and UO_1620 (O_1620,N_14298,N_12700);
and UO_1621 (O_1621,N_14965,N_14344);
nand UO_1622 (O_1622,N_14038,N_13597);
nand UO_1623 (O_1623,N_13696,N_12118);
nor UO_1624 (O_1624,N_13517,N_13893);
and UO_1625 (O_1625,N_12273,N_13527);
xor UO_1626 (O_1626,N_12937,N_13317);
nand UO_1627 (O_1627,N_12119,N_13070);
or UO_1628 (O_1628,N_13702,N_13404);
or UO_1629 (O_1629,N_14619,N_14590);
or UO_1630 (O_1630,N_13058,N_14868);
nand UO_1631 (O_1631,N_14674,N_14389);
or UO_1632 (O_1632,N_12586,N_14115);
and UO_1633 (O_1633,N_12620,N_14118);
nor UO_1634 (O_1634,N_13491,N_14132);
nand UO_1635 (O_1635,N_14199,N_13235);
or UO_1636 (O_1636,N_13023,N_12390);
nand UO_1637 (O_1637,N_12725,N_12292);
nor UO_1638 (O_1638,N_12689,N_13403);
nor UO_1639 (O_1639,N_14787,N_12528);
nor UO_1640 (O_1640,N_12937,N_14250);
nand UO_1641 (O_1641,N_14081,N_12011);
and UO_1642 (O_1642,N_12248,N_12960);
nor UO_1643 (O_1643,N_14366,N_12150);
nor UO_1644 (O_1644,N_13678,N_12956);
or UO_1645 (O_1645,N_12715,N_14232);
and UO_1646 (O_1646,N_13743,N_14150);
and UO_1647 (O_1647,N_12026,N_13732);
or UO_1648 (O_1648,N_13988,N_14463);
nor UO_1649 (O_1649,N_13166,N_13341);
or UO_1650 (O_1650,N_14381,N_12972);
or UO_1651 (O_1651,N_12459,N_13374);
nand UO_1652 (O_1652,N_13324,N_13409);
and UO_1653 (O_1653,N_13218,N_13403);
and UO_1654 (O_1654,N_12902,N_13471);
and UO_1655 (O_1655,N_14244,N_12166);
nor UO_1656 (O_1656,N_13967,N_14544);
and UO_1657 (O_1657,N_13465,N_13823);
or UO_1658 (O_1658,N_12464,N_14462);
or UO_1659 (O_1659,N_12772,N_12304);
or UO_1660 (O_1660,N_13423,N_14808);
nand UO_1661 (O_1661,N_12770,N_13116);
and UO_1662 (O_1662,N_12201,N_13815);
nand UO_1663 (O_1663,N_13860,N_13341);
nand UO_1664 (O_1664,N_14449,N_12116);
or UO_1665 (O_1665,N_12893,N_14164);
nor UO_1666 (O_1666,N_14603,N_13804);
nor UO_1667 (O_1667,N_12937,N_12179);
and UO_1668 (O_1668,N_12864,N_13574);
nand UO_1669 (O_1669,N_13485,N_14204);
or UO_1670 (O_1670,N_13429,N_14817);
or UO_1671 (O_1671,N_12173,N_14804);
or UO_1672 (O_1672,N_13887,N_12222);
and UO_1673 (O_1673,N_12470,N_13418);
nor UO_1674 (O_1674,N_14269,N_14716);
nor UO_1675 (O_1675,N_12819,N_12962);
or UO_1676 (O_1676,N_14010,N_14486);
nor UO_1677 (O_1677,N_13921,N_12665);
nor UO_1678 (O_1678,N_12719,N_14934);
nand UO_1679 (O_1679,N_12360,N_13916);
nor UO_1680 (O_1680,N_13675,N_12803);
nand UO_1681 (O_1681,N_13681,N_14374);
and UO_1682 (O_1682,N_14383,N_12703);
and UO_1683 (O_1683,N_12588,N_14683);
or UO_1684 (O_1684,N_12661,N_12946);
or UO_1685 (O_1685,N_13890,N_14635);
and UO_1686 (O_1686,N_12329,N_12357);
nand UO_1687 (O_1687,N_12213,N_13476);
nor UO_1688 (O_1688,N_14164,N_12697);
and UO_1689 (O_1689,N_13509,N_14648);
or UO_1690 (O_1690,N_13777,N_14891);
nand UO_1691 (O_1691,N_13006,N_12915);
nor UO_1692 (O_1692,N_12278,N_12639);
nor UO_1693 (O_1693,N_13537,N_14046);
nor UO_1694 (O_1694,N_14884,N_14644);
and UO_1695 (O_1695,N_13268,N_12541);
nor UO_1696 (O_1696,N_13508,N_14919);
and UO_1697 (O_1697,N_12907,N_14837);
nor UO_1698 (O_1698,N_12327,N_12430);
and UO_1699 (O_1699,N_12257,N_14005);
nor UO_1700 (O_1700,N_13744,N_14140);
and UO_1701 (O_1701,N_12415,N_13982);
or UO_1702 (O_1702,N_13187,N_14651);
xor UO_1703 (O_1703,N_12116,N_13228);
nor UO_1704 (O_1704,N_14647,N_12728);
nand UO_1705 (O_1705,N_13951,N_13713);
and UO_1706 (O_1706,N_12494,N_12529);
or UO_1707 (O_1707,N_14131,N_12781);
nand UO_1708 (O_1708,N_14526,N_13340);
nor UO_1709 (O_1709,N_12579,N_13653);
and UO_1710 (O_1710,N_14604,N_14594);
nor UO_1711 (O_1711,N_13535,N_14404);
nand UO_1712 (O_1712,N_14708,N_13869);
or UO_1713 (O_1713,N_12120,N_13156);
nand UO_1714 (O_1714,N_14395,N_13684);
and UO_1715 (O_1715,N_14928,N_13206);
nand UO_1716 (O_1716,N_13018,N_12187);
nand UO_1717 (O_1717,N_12346,N_12926);
or UO_1718 (O_1718,N_13980,N_12477);
nand UO_1719 (O_1719,N_14808,N_13120);
and UO_1720 (O_1720,N_14878,N_12404);
nand UO_1721 (O_1721,N_14319,N_14441);
nor UO_1722 (O_1722,N_14247,N_12218);
nor UO_1723 (O_1723,N_12053,N_12064);
or UO_1724 (O_1724,N_14001,N_12012);
nor UO_1725 (O_1725,N_13046,N_12799);
nand UO_1726 (O_1726,N_13390,N_13431);
and UO_1727 (O_1727,N_13721,N_13317);
nand UO_1728 (O_1728,N_14645,N_14832);
or UO_1729 (O_1729,N_13847,N_14696);
or UO_1730 (O_1730,N_14842,N_12860);
or UO_1731 (O_1731,N_13753,N_13571);
nor UO_1732 (O_1732,N_12547,N_14391);
nor UO_1733 (O_1733,N_12463,N_14812);
or UO_1734 (O_1734,N_12162,N_12825);
and UO_1735 (O_1735,N_13732,N_12927);
or UO_1736 (O_1736,N_14242,N_12283);
or UO_1737 (O_1737,N_12498,N_14052);
and UO_1738 (O_1738,N_13379,N_14684);
or UO_1739 (O_1739,N_14872,N_14325);
or UO_1740 (O_1740,N_14748,N_14915);
nor UO_1741 (O_1741,N_12920,N_13545);
nand UO_1742 (O_1742,N_14021,N_12094);
nor UO_1743 (O_1743,N_13892,N_13242);
or UO_1744 (O_1744,N_14148,N_14951);
nor UO_1745 (O_1745,N_13979,N_13252);
or UO_1746 (O_1746,N_12174,N_14172);
and UO_1747 (O_1747,N_13628,N_12321);
nand UO_1748 (O_1748,N_12531,N_12949);
xnor UO_1749 (O_1749,N_14012,N_14011);
nor UO_1750 (O_1750,N_13951,N_13461);
nand UO_1751 (O_1751,N_12201,N_12167);
or UO_1752 (O_1752,N_12315,N_14682);
nor UO_1753 (O_1753,N_13189,N_14790);
and UO_1754 (O_1754,N_12213,N_14488);
or UO_1755 (O_1755,N_13922,N_14614);
and UO_1756 (O_1756,N_13916,N_12479);
nor UO_1757 (O_1757,N_12296,N_13617);
nand UO_1758 (O_1758,N_13242,N_12387);
and UO_1759 (O_1759,N_13841,N_12756);
nand UO_1760 (O_1760,N_12102,N_14452);
and UO_1761 (O_1761,N_13293,N_14420);
nor UO_1762 (O_1762,N_13041,N_12611);
or UO_1763 (O_1763,N_13488,N_14758);
and UO_1764 (O_1764,N_12818,N_13372);
and UO_1765 (O_1765,N_13447,N_12820);
and UO_1766 (O_1766,N_13637,N_12921);
nand UO_1767 (O_1767,N_12661,N_12789);
or UO_1768 (O_1768,N_14497,N_12802);
nor UO_1769 (O_1769,N_13689,N_13714);
nand UO_1770 (O_1770,N_13650,N_14230);
nand UO_1771 (O_1771,N_14823,N_12399);
nand UO_1772 (O_1772,N_12957,N_14695);
and UO_1773 (O_1773,N_12012,N_13320);
nor UO_1774 (O_1774,N_12254,N_13195);
and UO_1775 (O_1775,N_12620,N_13369);
or UO_1776 (O_1776,N_13739,N_12769);
and UO_1777 (O_1777,N_13795,N_13501);
nand UO_1778 (O_1778,N_13765,N_14923);
or UO_1779 (O_1779,N_14504,N_13452);
or UO_1780 (O_1780,N_14656,N_14276);
nor UO_1781 (O_1781,N_14309,N_14421);
and UO_1782 (O_1782,N_12684,N_14100);
nor UO_1783 (O_1783,N_13527,N_12564);
nand UO_1784 (O_1784,N_13023,N_12789);
nand UO_1785 (O_1785,N_12625,N_13044);
or UO_1786 (O_1786,N_14709,N_13816);
and UO_1787 (O_1787,N_12376,N_12950);
nor UO_1788 (O_1788,N_14528,N_13815);
nor UO_1789 (O_1789,N_14054,N_14066);
nand UO_1790 (O_1790,N_14442,N_13580);
or UO_1791 (O_1791,N_14511,N_13110);
and UO_1792 (O_1792,N_13641,N_14374);
nor UO_1793 (O_1793,N_14960,N_13059);
nand UO_1794 (O_1794,N_13935,N_14761);
and UO_1795 (O_1795,N_12275,N_13227);
nor UO_1796 (O_1796,N_13764,N_13873);
nand UO_1797 (O_1797,N_12019,N_14767);
nand UO_1798 (O_1798,N_14576,N_14541);
nor UO_1799 (O_1799,N_14516,N_12508);
and UO_1800 (O_1800,N_13293,N_13395);
nor UO_1801 (O_1801,N_14121,N_14106);
or UO_1802 (O_1802,N_12456,N_13361);
or UO_1803 (O_1803,N_14645,N_12167);
nand UO_1804 (O_1804,N_13978,N_13699);
and UO_1805 (O_1805,N_12758,N_12183);
or UO_1806 (O_1806,N_13737,N_14506);
nand UO_1807 (O_1807,N_14242,N_13534);
and UO_1808 (O_1808,N_12182,N_14261);
xnor UO_1809 (O_1809,N_14828,N_12981);
nor UO_1810 (O_1810,N_13397,N_12612);
nand UO_1811 (O_1811,N_12573,N_13274);
and UO_1812 (O_1812,N_12387,N_13290);
or UO_1813 (O_1813,N_13930,N_13185);
or UO_1814 (O_1814,N_12032,N_13262);
or UO_1815 (O_1815,N_12591,N_12388);
nor UO_1816 (O_1816,N_12435,N_12198);
nor UO_1817 (O_1817,N_13010,N_13174);
nor UO_1818 (O_1818,N_14506,N_12680);
nor UO_1819 (O_1819,N_13827,N_14765);
nand UO_1820 (O_1820,N_13518,N_14446);
or UO_1821 (O_1821,N_14749,N_12336);
nand UO_1822 (O_1822,N_14605,N_13406);
or UO_1823 (O_1823,N_12878,N_13654);
nor UO_1824 (O_1824,N_12918,N_14346);
nand UO_1825 (O_1825,N_13081,N_14488);
nand UO_1826 (O_1826,N_14962,N_13859);
and UO_1827 (O_1827,N_12471,N_14350);
and UO_1828 (O_1828,N_12705,N_12084);
and UO_1829 (O_1829,N_13542,N_14202);
or UO_1830 (O_1830,N_12344,N_13333);
nand UO_1831 (O_1831,N_14459,N_14299);
or UO_1832 (O_1832,N_12433,N_12268);
nand UO_1833 (O_1833,N_12944,N_12762);
nor UO_1834 (O_1834,N_14721,N_14164);
and UO_1835 (O_1835,N_12364,N_14853);
and UO_1836 (O_1836,N_13694,N_12597);
and UO_1837 (O_1837,N_13781,N_13085);
or UO_1838 (O_1838,N_12297,N_13627);
or UO_1839 (O_1839,N_12958,N_13031);
and UO_1840 (O_1840,N_14213,N_12593);
and UO_1841 (O_1841,N_12521,N_14978);
and UO_1842 (O_1842,N_13694,N_13880);
or UO_1843 (O_1843,N_14117,N_12914);
or UO_1844 (O_1844,N_13949,N_14168);
nand UO_1845 (O_1845,N_13170,N_12867);
or UO_1846 (O_1846,N_14934,N_14298);
and UO_1847 (O_1847,N_14877,N_12640);
nor UO_1848 (O_1848,N_12483,N_13242);
or UO_1849 (O_1849,N_14984,N_13075);
or UO_1850 (O_1850,N_13341,N_12232);
nand UO_1851 (O_1851,N_13116,N_13224);
nor UO_1852 (O_1852,N_14463,N_12365);
or UO_1853 (O_1853,N_13087,N_12950);
nand UO_1854 (O_1854,N_14496,N_14626);
nand UO_1855 (O_1855,N_14114,N_13302);
nor UO_1856 (O_1856,N_14569,N_13917);
nor UO_1857 (O_1857,N_14634,N_14994);
or UO_1858 (O_1858,N_14827,N_14503);
or UO_1859 (O_1859,N_12073,N_13940);
nor UO_1860 (O_1860,N_12334,N_13085);
and UO_1861 (O_1861,N_13013,N_12065);
nor UO_1862 (O_1862,N_13866,N_12473);
or UO_1863 (O_1863,N_12279,N_13827);
or UO_1864 (O_1864,N_14500,N_14775);
or UO_1865 (O_1865,N_12078,N_13930);
nor UO_1866 (O_1866,N_12794,N_12774);
and UO_1867 (O_1867,N_12582,N_12066);
and UO_1868 (O_1868,N_14547,N_12252);
nor UO_1869 (O_1869,N_13464,N_14473);
nand UO_1870 (O_1870,N_13880,N_13401);
and UO_1871 (O_1871,N_14538,N_12253);
and UO_1872 (O_1872,N_12008,N_12236);
nor UO_1873 (O_1873,N_12814,N_12322);
nand UO_1874 (O_1874,N_12123,N_14026);
nor UO_1875 (O_1875,N_13325,N_14430);
nand UO_1876 (O_1876,N_13135,N_14778);
nor UO_1877 (O_1877,N_12701,N_13999);
nand UO_1878 (O_1878,N_14703,N_14532);
or UO_1879 (O_1879,N_14291,N_13529);
and UO_1880 (O_1880,N_13370,N_13243);
nand UO_1881 (O_1881,N_13961,N_14195);
and UO_1882 (O_1882,N_12264,N_12468);
nor UO_1883 (O_1883,N_13039,N_13085);
and UO_1884 (O_1884,N_13629,N_13073);
and UO_1885 (O_1885,N_14085,N_13950);
and UO_1886 (O_1886,N_14303,N_14677);
or UO_1887 (O_1887,N_14652,N_13532);
and UO_1888 (O_1888,N_13941,N_13688);
nor UO_1889 (O_1889,N_13034,N_14229);
or UO_1890 (O_1890,N_12264,N_12938);
and UO_1891 (O_1891,N_14378,N_12960);
xnor UO_1892 (O_1892,N_13504,N_12487);
and UO_1893 (O_1893,N_12817,N_13325);
nor UO_1894 (O_1894,N_12220,N_14397);
nand UO_1895 (O_1895,N_12482,N_12934);
or UO_1896 (O_1896,N_12576,N_14717);
nor UO_1897 (O_1897,N_14793,N_13547);
or UO_1898 (O_1898,N_12604,N_14296);
nor UO_1899 (O_1899,N_12087,N_13585);
nand UO_1900 (O_1900,N_12147,N_13790);
and UO_1901 (O_1901,N_13733,N_12107);
nand UO_1902 (O_1902,N_14850,N_14120);
and UO_1903 (O_1903,N_13019,N_14538);
or UO_1904 (O_1904,N_13175,N_13011);
nand UO_1905 (O_1905,N_13381,N_12463);
nand UO_1906 (O_1906,N_13847,N_14528);
or UO_1907 (O_1907,N_12263,N_13232);
nor UO_1908 (O_1908,N_14921,N_13524);
or UO_1909 (O_1909,N_13949,N_12109);
nor UO_1910 (O_1910,N_13026,N_13801);
and UO_1911 (O_1911,N_13046,N_14623);
nor UO_1912 (O_1912,N_13171,N_12464);
or UO_1913 (O_1913,N_13057,N_14969);
nor UO_1914 (O_1914,N_13896,N_12871);
nand UO_1915 (O_1915,N_12977,N_13076);
and UO_1916 (O_1916,N_12390,N_14946);
and UO_1917 (O_1917,N_13504,N_13935);
and UO_1918 (O_1918,N_13667,N_13217);
nor UO_1919 (O_1919,N_12937,N_12820);
nor UO_1920 (O_1920,N_14922,N_13145);
nand UO_1921 (O_1921,N_14614,N_12358);
nor UO_1922 (O_1922,N_13137,N_13677);
xnor UO_1923 (O_1923,N_13488,N_12180);
and UO_1924 (O_1924,N_12021,N_14658);
and UO_1925 (O_1925,N_14925,N_13728);
or UO_1926 (O_1926,N_12900,N_14146);
nand UO_1927 (O_1927,N_14576,N_14922);
nand UO_1928 (O_1928,N_14648,N_13498);
nor UO_1929 (O_1929,N_13369,N_13694);
nor UO_1930 (O_1930,N_14778,N_14979);
or UO_1931 (O_1931,N_12892,N_12055);
nor UO_1932 (O_1932,N_12614,N_12499);
and UO_1933 (O_1933,N_12392,N_12025);
nor UO_1934 (O_1934,N_12180,N_14989);
nor UO_1935 (O_1935,N_14378,N_14658);
nor UO_1936 (O_1936,N_12803,N_13673);
and UO_1937 (O_1937,N_12945,N_12889);
nor UO_1938 (O_1938,N_14310,N_14561);
or UO_1939 (O_1939,N_13165,N_12402);
or UO_1940 (O_1940,N_12911,N_14599);
or UO_1941 (O_1941,N_13644,N_13953);
or UO_1942 (O_1942,N_12693,N_12836);
nand UO_1943 (O_1943,N_13634,N_13873);
or UO_1944 (O_1944,N_13191,N_12563);
and UO_1945 (O_1945,N_12341,N_13082);
and UO_1946 (O_1946,N_14213,N_13623);
and UO_1947 (O_1947,N_12762,N_13004);
and UO_1948 (O_1948,N_14257,N_12283);
or UO_1949 (O_1949,N_12583,N_13885);
and UO_1950 (O_1950,N_12772,N_14002);
nor UO_1951 (O_1951,N_12700,N_13039);
or UO_1952 (O_1952,N_12324,N_12001);
nor UO_1953 (O_1953,N_12684,N_12286);
nand UO_1954 (O_1954,N_13121,N_14462);
or UO_1955 (O_1955,N_12739,N_14212);
and UO_1956 (O_1956,N_13131,N_12389);
nor UO_1957 (O_1957,N_13726,N_13350);
or UO_1958 (O_1958,N_13199,N_13107);
nor UO_1959 (O_1959,N_12587,N_13342);
or UO_1960 (O_1960,N_13962,N_13785);
and UO_1961 (O_1961,N_12494,N_14734);
or UO_1962 (O_1962,N_12417,N_14826);
nor UO_1963 (O_1963,N_14422,N_14775);
nand UO_1964 (O_1964,N_13095,N_14440);
nor UO_1965 (O_1965,N_13556,N_12562);
nor UO_1966 (O_1966,N_13303,N_14267);
and UO_1967 (O_1967,N_14735,N_12995);
nor UO_1968 (O_1968,N_13206,N_14932);
or UO_1969 (O_1969,N_12341,N_12344);
and UO_1970 (O_1970,N_14761,N_13202);
nor UO_1971 (O_1971,N_12350,N_14031);
or UO_1972 (O_1972,N_12125,N_14801);
nand UO_1973 (O_1973,N_12001,N_13559);
nand UO_1974 (O_1974,N_13212,N_13302);
or UO_1975 (O_1975,N_12895,N_12151);
or UO_1976 (O_1976,N_14054,N_13077);
and UO_1977 (O_1977,N_13693,N_12647);
nor UO_1978 (O_1978,N_14075,N_12719);
xor UO_1979 (O_1979,N_12765,N_14382);
nor UO_1980 (O_1980,N_14542,N_14451);
nor UO_1981 (O_1981,N_14768,N_13535);
nor UO_1982 (O_1982,N_12138,N_12491);
nor UO_1983 (O_1983,N_12653,N_12460);
nand UO_1984 (O_1984,N_13482,N_14993);
nor UO_1985 (O_1985,N_12505,N_12398);
nand UO_1986 (O_1986,N_12708,N_14359);
nor UO_1987 (O_1987,N_13827,N_12534);
nor UO_1988 (O_1988,N_12290,N_13515);
nor UO_1989 (O_1989,N_14165,N_13708);
and UO_1990 (O_1990,N_13995,N_13243);
nor UO_1991 (O_1991,N_14747,N_12103);
and UO_1992 (O_1992,N_14890,N_14061);
nor UO_1993 (O_1993,N_13042,N_12215);
nor UO_1994 (O_1994,N_13849,N_14597);
nor UO_1995 (O_1995,N_14988,N_13082);
nor UO_1996 (O_1996,N_14809,N_14195);
nand UO_1997 (O_1997,N_14798,N_12727);
nor UO_1998 (O_1998,N_12717,N_13393);
nor UO_1999 (O_1999,N_13685,N_12355);
endmodule