module basic_1000_10000_1500_50_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_86,In_438);
and U1 (N_1,In_39,In_185);
or U2 (N_2,In_357,In_969);
nand U3 (N_3,In_790,In_267);
nand U4 (N_4,In_749,In_446);
nand U5 (N_5,In_872,In_799);
nand U6 (N_6,In_36,In_552);
nand U7 (N_7,In_4,In_873);
nand U8 (N_8,In_6,In_852);
or U9 (N_9,In_380,In_459);
xnor U10 (N_10,In_254,In_468);
nand U11 (N_11,In_609,In_440);
nor U12 (N_12,In_278,In_309);
nor U13 (N_13,In_783,In_867);
nor U14 (N_14,In_302,In_500);
nand U15 (N_15,In_788,In_526);
nor U16 (N_16,In_818,In_83);
and U17 (N_17,In_522,In_305);
nand U18 (N_18,In_976,In_660);
and U19 (N_19,In_212,In_166);
or U20 (N_20,In_71,In_194);
nor U21 (N_21,In_327,In_745);
and U22 (N_22,In_883,In_579);
nor U23 (N_23,In_82,In_805);
nand U24 (N_24,In_504,In_283);
nor U25 (N_25,In_957,In_333);
or U26 (N_26,In_493,In_454);
nor U27 (N_27,In_699,In_251);
or U28 (N_28,In_938,In_501);
nand U29 (N_29,In_926,In_404);
or U30 (N_30,In_59,In_203);
and U31 (N_31,In_310,In_847);
nor U32 (N_32,In_763,In_915);
and U33 (N_33,In_591,In_663);
and U34 (N_34,In_94,In_625);
nor U35 (N_35,In_292,In_256);
nand U36 (N_36,In_375,In_131);
nor U37 (N_37,In_686,In_61);
nand U38 (N_38,In_328,In_144);
and U39 (N_39,In_447,In_416);
and U40 (N_40,In_18,In_627);
nor U41 (N_41,In_920,In_40);
and U42 (N_42,In_979,In_257);
and U43 (N_43,In_260,In_177);
nor U44 (N_44,In_693,In_518);
and U45 (N_45,In_602,In_608);
nor U46 (N_46,In_628,In_372);
nand U47 (N_47,In_713,In_760);
nand U48 (N_48,In_258,In_350);
or U49 (N_49,In_48,In_918);
or U50 (N_50,In_529,In_678);
nor U51 (N_51,In_630,In_572);
nor U52 (N_52,In_953,In_961);
xnor U53 (N_53,In_596,In_561);
and U54 (N_54,In_263,In_234);
nand U55 (N_55,In_820,In_181);
or U56 (N_56,In_174,In_288);
and U57 (N_57,In_385,In_394);
or U58 (N_58,In_189,In_368);
and U59 (N_59,In_742,In_943);
nand U60 (N_60,In_248,In_449);
nor U61 (N_61,In_925,In_472);
and U62 (N_62,In_183,In_530);
xnor U63 (N_63,In_574,In_272);
nand U64 (N_64,In_941,In_800);
nor U65 (N_65,In_866,In_746);
or U66 (N_66,In_549,In_452);
or U67 (N_67,In_296,In_707);
nand U68 (N_68,In_448,In_268);
and U69 (N_69,In_455,In_589);
nor U70 (N_70,In_25,In_668);
and U71 (N_71,In_963,In_215);
nand U72 (N_72,In_999,In_240);
xor U73 (N_73,In_17,In_191);
nand U74 (N_74,In_116,In_422);
xnor U75 (N_75,In_261,In_541);
nor U76 (N_76,In_726,In_559);
nor U77 (N_77,In_13,In_532);
nor U78 (N_78,In_67,In_954);
nand U79 (N_79,In_8,In_885);
or U80 (N_80,In_58,In_893);
or U81 (N_81,In_667,In_271);
or U82 (N_82,In_496,In_764);
nand U83 (N_83,In_233,In_970);
or U84 (N_84,In_169,In_806);
nor U85 (N_85,In_875,In_362);
or U86 (N_86,In_619,In_64);
or U87 (N_87,In_655,In_562);
nand U88 (N_88,In_47,In_733);
nor U89 (N_89,In_694,In_192);
nor U90 (N_90,In_980,In_340);
nor U91 (N_91,In_535,In_218);
nor U92 (N_92,In_499,In_924);
nor U93 (N_93,In_457,In_408);
nand U94 (N_94,In_626,In_117);
or U95 (N_95,In_402,In_836);
nand U96 (N_96,In_276,In_364);
or U97 (N_97,In_179,In_456);
or U98 (N_98,In_382,In_275);
and U99 (N_99,In_978,In_365);
nor U100 (N_100,In_149,In_486);
or U101 (N_101,In_928,In_343);
or U102 (N_102,In_986,In_141);
nor U103 (N_103,In_615,In_994);
and U104 (N_104,In_880,In_75);
or U105 (N_105,In_570,In_88);
nor U106 (N_106,In_546,In_286);
nor U107 (N_107,In_871,In_613);
nand U108 (N_108,In_462,In_844);
nor U109 (N_109,In_821,In_200);
and U110 (N_110,In_564,In_510);
or U111 (N_111,In_768,In_264);
and U112 (N_112,In_139,In_284);
or U113 (N_113,In_709,In_172);
and U114 (N_114,In_441,In_491);
or U115 (N_115,In_654,In_160);
nor U116 (N_116,In_736,In_273);
and U117 (N_117,In_933,In_837);
nor U118 (N_118,In_600,In_962);
and U119 (N_119,In_931,In_330);
nor U120 (N_120,In_831,In_474);
or U121 (N_121,In_984,In_940);
and U122 (N_122,In_803,In_358);
or U123 (N_123,In_665,In_405);
nor U124 (N_124,In_796,In_823);
and U125 (N_125,In_658,In_731);
and U126 (N_126,In_503,In_539);
nor U127 (N_127,In_817,In_31);
nor U128 (N_128,In_639,In_460);
or U129 (N_129,In_996,In_725);
nor U130 (N_130,In_566,In_188);
nor U131 (N_131,In_308,In_41);
or U132 (N_132,In_27,In_555);
nor U133 (N_133,In_96,In_680);
nor U134 (N_134,In_683,In_700);
nor U135 (N_135,In_519,In_133);
or U136 (N_136,In_765,In_85);
or U137 (N_137,In_479,In_87);
or U138 (N_138,In_193,In_390);
and U139 (N_139,In_672,In_576);
and U140 (N_140,In_524,In_319);
nand U141 (N_141,In_826,In_793);
and U142 (N_142,In_214,In_485);
nand U143 (N_143,In_345,In_137);
or U144 (N_144,In_10,In_974);
nor U145 (N_145,In_12,In_740);
nor U146 (N_146,In_685,In_662);
nand U147 (N_147,In_274,In_293);
or U148 (N_148,In_482,In_331);
nand U149 (N_149,In_761,In_159);
xor U150 (N_150,In_673,In_597);
and U151 (N_151,In_550,In_766);
nand U152 (N_152,In_142,In_516);
nand U153 (N_153,In_987,In_723);
and U154 (N_154,In_509,In_495);
xor U155 (N_155,In_311,In_32);
nand U156 (N_156,In_0,In_729);
nor U157 (N_157,In_966,In_81);
and U158 (N_158,In_130,In_593);
xnor U159 (N_159,In_949,In_666);
nand U160 (N_160,In_923,In_582);
nand U161 (N_161,In_538,In_900);
nand U162 (N_162,In_476,In_477);
and U163 (N_163,In_605,In_815);
nor U164 (N_164,In_860,In_548);
nor U165 (N_165,In_718,In_414);
and U166 (N_166,In_363,In_878);
xor U167 (N_167,In_512,In_968);
nand U168 (N_168,In_982,In_488);
nor U169 (N_169,In_786,In_209);
nor U170 (N_170,In_415,In_389);
and U171 (N_171,In_62,In_124);
nand U172 (N_172,In_315,In_198);
nand U173 (N_173,In_249,In_134);
nor U174 (N_174,In_377,In_676);
nor U175 (N_175,In_927,In_601);
nor U176 (N_176,In_703,In_262);
nor U177 (N_177,In_802,In_287);
nor U178 (N_178,In_877,In_281);
and U179 (N_179,In_858,In_577);
nand U180 (N_180,In_688,In_103);
and U181 (N_181,In_184,In_584);
nor U182 (N_182,In_235,In_53);
and U183 (N_183,In_640,In_199);
nand U184 (N_184,In_341,In_644);
nor U185 (N_185,In_16,In_161);
nor U186 (N_186,In_279,In_669);
and U187 (N_187,In_956,In_621);
xor U188 (N_188,In_451,In_480);
and U189 (N_189,In_536,In_913);
nand U190 (N_190,In_643,In_635);
nand U191 (N_191,In_527,In_945);
nor U192 (N_192,In_517,In_386);
and U193 (N_193,In_917,In_939);
nand U194 (N_194,In_899,In_722);
nand U195 (N_195,In_612,In_430);
or U196 (N_196,In_881,In_219);
or U197 (N_197,In_239,In_861);
nor U198 (N_198,In_972,In_370);
and U199 (N_199,In_56,In_417);
and U200 (N_200,In_471,In_180);
and U201 (N_201,In_306,In_946);
and U202 (N_202,In_3,In_421);
nor U203 (N_203,N_196,In_997);
nand U204 (N_204,In_171,In_674);
or U205 (N_205,In_778,N_26);
nor U206 (N_206,In_383,In_458);
or U207 (N_207,In_929,N_111);
and U208 (N_208,In_808,In_592);
nor U209 (N_209,In_779,N_191);
nand U210 (N_210,In_294,In_428);
nand U211 (N_211,In_716,In_696);
nand U212 (N_212,In_907,In_981);
and U213 (N_213,In_51,In_659);
or U214 (N_214,In_897,N_173);
nand U215 (N_215,In_326,N_199);
nand U216 (N_216,In_352,In_28);
nand U217 (N_217,In_342,In_178);
nand U218 (N_218,In_425,In_588);
nand U219 (N_219,In_348,In_2);
nor U220 (N_220,N_39,In_114);
nand U221 (N_221,N_12,In_698);
and U222 (N_222,In_490,N_163);
or U223 (N_223,In_366,N_113);
nand U224 (N_224,In_487,In_226);
nor U225 (N_225,N_161,In_231);
or U226 (N_226,N_192,In_632);
nor U227 (N_227,In_842,In_955);
nand U228 (N_228,In_834,In_759);
nand U229 (N_229,In_886,In_657);
nor U230 (N_230,In_195,N_62);
and U231 (N_231,In_229,In_176);
and U232 (N_232,In_754,N_7);
nand U233 (N_233,In_201,In_104);
or U234 (N_234,In_896,N_190);
and U235 (N_235,In_747,In_413);
nand U236 (N_236,N_162,In_599);
and U237 (N_237,In_113,In_398);
nand U238 (N_238,In_905,In_967);
and U239 (N_239,N_168,In_156);
nand U240 (N_240,N_45,In_316);
or U241 (N_241,In_167,N_20);
and U242 (N_242,In_537,In_473);
nand U243 (N_243,In_424,In_521);
nand U244 (N_244,In_610,In_638);
nor U245 (N_245,In_429,N_129);
nand U246 (N_246,In_323,In_687);
nor U247 (N_247,In_126,In_433);
nor U248 (N_248,In_182,N_60);
nor U249 (N_249,In_838,In_965);
and U250 (N_250,In_656,In_937);
and U251 (N_251,In_387,N_132);
and U252 (N_252,N_151,N_147);
nand U253 (N_253,In_888,In_265);
nor U254 (N_254,In_206,N_165);
or U255 (N_255,In_848,In_393);
nor U256 (N_256,N_138,In_775);
xnor U257 (N_257,In_849,In_771);
and U258 (N_258,In_461,In_162);
and U259 (N_259,N_194,In_355);
or U260 (N_260,N_87,In_551);
nand U261 (N_261,In_186,In_606);
or U262 (N_262,In_136,In_406);
nand U263 (N_263,In_435,In_734);
and U264 (N_264,N_180,N_121);
nand U265 (N_265,N_46,In_300);
and U266 (N_266,N_94,In_902);
or U267 (N_267,In_641,N_169);
nor U268 (N_268,In_128,In_297);
and U269 (N_269,In_313,In_908);
nand U270 (N_270,N_116,In_367);
or U271 (N_271,N_40,In_135);
nand U272 (N_272,In_857,In_906);
or U273 (N_273,N_179,In_89);
nand U274 (N_274,N_198,N_125);
nand U275 (N_275,In_557,In_418);
nand U276 (N_276,N_117,In_998);
and U277 (N_277,In_715,In_228);
nor U278 (N_278,In_629,In_360);
and U279 (N_279,In_840,In_34);
nor U280 (N_280,N_32,In_507);
nor U281 (N_281,N_41,In_554);
and U282 (N_282,N_50,In_318);
nor U283 (N_283,In_569,In_735);
or U284 (N_284,In_420,In_324);
nand U285 (N_285,N_184,N_103);
or U286 (N_286,In_502,In_453);
and U287 (N_287,N_85,In_371);
nand U288 (N_288,N_59,N_64);
nor U289 (N_289,In_769,In_814);
or U290 (N_290,In_391,In_781);
nand U291 (N_291,In_72,In_197);
nand U292 (N_292,N_38,In_622);
nand U293 (N_293,In_110,In_791);
and U294 (N_294,In_339,N_183);
or U295 (N_295,In_708,In_813);
and U296 (N_296,In_618,In_870);
nand U297 (N_297,In_993,In_758);
and U298 (N_298,In_533,In_646);
or U299 (N_299,In_792,In_243);
and U300 (N_300,In_798,In_334);
or U301 (N_301,N_110,In_173);
nand U302 (N_302,In_210,In_738);
nand U303 (N_303,In_361,In_780);
nand U304 (N_304,In_498,N_78);
or U305 (N_305,N_95,In_120);
or U306 (N_306,In_587,N_126);
or U307 (N_307,In_839,N_11);
nor U308 (N_308,N_72,In_384);
or U309 (N_309,N_80,In_648);
nor U310 (N_310,In_301,N_67);
and U311 (N_311,In_822,In_964);
and U312 (N_312,In_270,In_767);
and U313 (N_313,In_168,In_583);
nand U314 (N_314,N_93,In_743);
nand U315 (N_315,N_176,In_804);
and U316 (N_316,N_79,In_221);
xnor U317 (N_317,In_95,In_105);
or U318 (N_318,In_912,In_921);
nand U319 (N_319,In_565,N_100);
xor U320 (N_320,In_483,In_481);
nand U321 (N_321,In_388,In_238);
or U322 (N_322,In_190,In_155);
nand U323 (N_323,N_155,In_187);
nand U324 (N_324,N_58,N_63);
xnor U325 (N_325,In_236,In_789);
or U326 (N_326,In_304,In_637);
and U327 (N_327,In_374,N_29);
and U328 (N_328,In_801,In_427);
and U329 (N_329,In_730,In_732);
nand U330 (N_330,In_397,N_120);
nand U331 (N_331,In_671,N_3);
or U332 (N_332,N_28,In_409);
or U333 (N_333,N_92,In_494);
or U334 (N_334,N_193,N_101);
and U335 (N_335,In_910,In_381);
nand U336 (N_336,N_18,In_623);
and U337 (N_337,N_136,In_157);
nor U338 (N_338,In_977,In_354);
nand U339 (N_339,N_88,In_7);
and U340 (N_340,In_988,N_71);
nand U341 (N_341,N_91,In_400);
or U342 (N_342,N_104,N_144);
nor U343 (N_343,In_146,In_148);
nand U344 (N_344,In_266,In_60);
nand U345 (N_345,In_332,In_846);
and U346 (N_346,N_152,In_299);
or U347 (N_347,In_211,In_691);
or U348 (N_348,N_84,In_598);
or U349 (N_349,In_603,In_695);
or U350 (N_350,N_119,N_86);
and U351 (N_351,In_369,In_80);
nor U352 (N_352,In_50,In_111);
and U353 (N_353,N_35,N_97);
nand U354 (N_354,In_807,N_0);
nor U355 (N_355,N_81,In_207);
and U356 (N_356,In_336,In_633);
or U357 (N_357,In_720,N_51);
or U358 (N_358,In_985,In_531);
nor U359 (N_359,N_31,In_947);
nand U360 (N_360,In_351,In_403);
nor U361 (N_361,In_558,In_9);
nor U362 (N_362,N_124,In_344);
xnor U363 (N_363,N_102,In_614);
nand U364 (N_364,In_690,In_950);
and U365 (N_365,In_337,In_904);
and U366 (N_366,In_320,N_53);
xor U367 (N_367,In_478,In_109);
nor U368 (N_368,In_845,In_661);
and U369 (N_369,In_125,N_6);
nor U370 (N_370,In_353,In_919);
and U371 (N_371,In_54,In_70);
nand U372 (N_372,In_119,In_100);
nand U373 (N_373,In_784,N_21);
xor U374 (N_374,In_329,N_73);
and U375 (N_375,In_68,N_107);
and U376 (N_376,In_827,In_443);
nor U377 (N_377,In_898,In_84);
nand U378 (N_378,N_10,In_43);
nor U379 (N_379,In_255,In_205);
and U380 (N_380,In_35,In_291);
and U381 (N_381,N_105,In_810);
nor U382 (N_382,In_702,In_63);
or U383 (N_383,In_108,In_140);
nor U384 (N_384,In_824,In_399);
nor U385 (N_385,N_114,In_830);
nor U386 (N_386,N_23,In_739);
nand U387 (N_387,In_123,In_122);
and U388 (N_388,In_5,In_98);
or U389 (N_389,In_379,In_289);
or U390 (N_390,In_77,In_989);
nor U391 (N_391,N_130,In_651);
nand U392 (N_392,In_508,In_412);
nor U393 (N_393,N_82,In_762);
nor U394 (N_394,In_511,In_202);
nor U395 (N_395,In_321,In_90);
and U396 (N_396,In_138,In_282);
nand U397 (N_397,In_213,In_505);
or U398 (N_398,In_556,In_465);
and U399 (N_399,In_607,In_692);
or U400 (N_400,In_143,N_318);
nand U401 (N_401,In_542,N_240);
and U402 (N_402,N_330,In_909);
nand U403 (N_403,In_751,In_719);
or U404 (N_404,N_57,N_374);
nor U405 (N_405,In_401,In_737);
or U406 (N_406,N_47,N_296);
nor U407 (N_407,N_314,In_890);
or U408 (N_408,In_816,N_244);
and U409 (N_409,In_595,N_291);
nor U410 (N_410,In_647,N_380);
nor U411 (N_411,N_44,N_289);
nand U412 (N_412,In_952,In_423);
nand U413 (N_413,In_664,In_545);
nand U414 (N_414,In_170,In_445);
or U415 (N_415,In_129,N_260);
and U416 (N_416,N_137,N_281);
nor U417 (N_417,In_825,N_167);
and U418 (N_418,In_497,In_835);
nand U419 (N_419,In_853,In_29);
or U420 (N_420,In_217,N_310);
and U421 (N_421,N_372,N_204);
nand U422 (N_422,In_594,In_704);
nand U423 (N_423,In_145,In_863);
or U424 (N_424,N_282,N_75);
nand U425 (N_425,N_337,N_272);
or U426 (N_426,In_944,In_1);
nor U427 (N_427,In_204,In_753);
nand U428 (N_428,N_207,In_489);
nand U429 (N_429,In_948,In_426);
or U430 (N_430,In_24,In_891);
and U431 (N_431,In_241,In_752);
nor U432 (N_432,In_958,N_370);
or U433 (N_433,N_224,N_321);
nand U434 (N_434,In_20,N_389);
and U435 (N_435,N_279,In_514);
and U436 (N_436,N_384,N_166);
and U437 (N_437,N_213,In_466);
or U438 (N_438,In_101,N_182);
or U439 (N_439,In_121,In_396);
nor U440 (N_440,N_232,N_208);
or U441 (N_441,N_24,In_611);
and U442 (N_442,In_620,In_991);
and U443 (N_443,N_329,N_70);
nand U444 (N_444,In_714,N_333);
and U445 (N_445,In_484,N_301);
and U446 (N_446,N_302,In_652);
or U447 (N_447,N_241,N_344);
nand U448 (N_448,N_178,In_76);
and U449 (N_449,N_36,N_42);
or U450 (N_450,In_227,N_33);
or U451 (N_451,N_254,In_645);
or U452 (N_452,In_112,N_292);
or U453 (N_453,In_677,N_186);
or U454 (N_454,In_617,N_66);
nand U455 (N_455,N_331,In_795);
nor U456 (N_456,In_33,In_894);
nor U457 (N_457,In_44,N_259);
nand U458 (N_458,In_165,In_728);
nor U459 (N_459,In_772,N_256);
and U460 (N_460,N_228,N_61);
and U461 (N_461,N_357,In_223);
and U462 (N_462,In_220,N_139);
or U463 (N_463,In_450,In_568);
nor U464 (N_464,N_251,N_397);
and U465 (N_465,In_540,In_819);
and U466 (N_466,In_757,N_262);
or U467 (N_467,N_171,N_170);
nor U468 (N_468,In_851,N_383);
and U469 (N_469,In_701,N_188);
and U470 (N_470,N_149,In_935);
and U471 (N_471,N_358,In_573);
or U472 (N_472,N_369,In_411);
nor U473 (N_473,In_895,In_46);
nand U474 (N_474,In_553,In_520);
xor U475 (N_475,In_843,N_392);
nand U476 (N_476,In_932,N_158);
nor U477 (N_477,In_49,In_392);
xnor U478 (N_478,In_469,N_209);
nand U479 (N_479,N_246,N_303);
and U480 (N_480,N_157,In_250);
nand U481 (N_481,N_252,N_148);
nor U482 (N_482,N_231,In_679);
nor U483 (N_483,In_253,N_49);
and U484 (N_484,N_211,In_829);
and U485 (N_485,N_112,N_395);
nor U486 (N_486,In_436,N_141);
xnor U487 (N_487,In_575,N_320);
nor U488 (N_488,In_544,N_68);
and U489 (N_489,N_17,In_439);
or U490 (N_490,In_727,In_528);
or U491 (N_491,N_172,N_309);
nand U492 (N_492,In_653,N_356);
or U493 (N_493,N_365,N_277);
and U494 (N_494,In_356,N_307);
and U495 (N_495,N_269,N_378);
nor U496 (N_496,N_229,In_298);
nand U497 (N_497,N_215,N_69);
and U498 (N_498,N_388,In_208);
or U499 (N_499,N_298,N_249);
nor U500 (N_500,In_684,N_350);
nor U501 (N_501,In_616,N_263);
or U502 (N_502,N_293,In_252);
nand U503 (N_503,N_223,In_395);
and U504 (N_504,In_99,N_236);
nand U505 (N_505,N_177,N_323);
nor U506 (N_506,N_122,In_314);
and U507 (N_507,N_327,N_218);
or U508 (N_508,In_785,N_96);
and U509 (N_509,N_237,N_349);
nor U510 (N_510,N_54,N_390);
and U511 (N_511,N_250,N_345);
nand U512 (N_512,N_385,N_242);
and U513 (N_513,N_195,In_78);
and U514 (N_514,N_160,In_335);
and U515 (N_515,N_83,In_523);
and U516 (N_516,In_776,In_65);
and U517 (N_517,N_13,N_219);
and U518 (N_518,N_290,N_352);
nor U519 (N_519,N_266,In_869);
or U520 (N_520,N_43,N_368);
nand U521 (N_521,In_936,N_348);
or U522 (N_522,N_367,In_922);
or U523 (N_523,N_156,N_164);
nor U524 (N_524,N_273,In_710);
nand U525 (N_525,N_9,N_37);
nor U526 (N_526,In_724,N_214);
nand U527 (N_527,In_280,N_27);
and U528 (N_528,In_52,In_164);
nor U529 (N_529,In_960,N_150);
and U530 (N_530,In_876,N_297);
nand U531 (N_531,In_879,In_543);
or U532 (N_532,N_271,In_850);
or U533 (N_533,N_265,In_983);
nand U534 (N_534,In_325,N_366);
nand U535 (N_535,In_990,N_77);
nor U536 (N_536,In_624,N_371);
or U537 (N_537,N_339,N_258);
and U538 (N_538,In_432,In_246);
or U539 (N_539,In_642,N_145);
nor U540 (N_540,In_995,In_444);
nand U541 (N_541,N_135,N_375);
and U542 (N_542,N_308,N_230);
and U543 (N_543,In_222,In_91);
nor U544 (N_544,N_131,In_604);
nand U545 (N_545,In_74,N_295);
nor U546 (N_546,N_133,N_270);
or U547 (N_547,N_288,N_159);
or U548 (N_548,In_756,In_230);
nor U549 (N_549,N_285,N_346);
nor U550 (N_550,In_748,N_226);
nand U551 (N_551,In_911,In_901);
or U552 (N_552,N_15,In_682);
and U553 (N_553,N_200,In_11);
and U554 (N_554,In_492,N_322);
or U555 (N_555,N_74,In_578);
or U556 (N_556,In_285,In_410);
nor U557 (N_557,In_127,N_278);
nor U558 (N_558,In_23,In_721);
nand U559 (N_559,In_307,N_394);
nor U560 (N_560,N_235,N_393);
and U561 (N_561,N_360,N_123);
or U562 (N_562,N_274,N_227);
or U563 (N_563,In_705,N_233);
or U564 (N_564,N_185,In_244);
or U565 (N_565,N_353,N_239);
nand U566 (N_566,In_914,In_649);
and U567 (N_567,In_464,In_349);
nor U568 (N_568,In_650,In_470);
nand U569 (N_569,In_862,N_342);
or U570 (N_570,N_108,In_959);
nor U571 (N_571,N_324,In_66);
or U572 (N_572,In_269,In_153);
nor U573 (N_573,N_206,In_290);
nand U574 (N_574,In_118,N_217);
or U575 (N_575,In_437,In_163);
nand U576 (N_576,N_118,N_355);
or U577 (N_577,In_744,In_859);
or U578 (N_578,In_152,N_205);
or U579 (N_579,N_134,N_127);
nor U580 (N_580,N_338,N_341);
or U581 (N_581,In_689,In_868);
or U582 (N_582,In_216,In_874);
xor U583 (N_583,N_247,In_15);
or U584 (N_584,In_277,In_547);
and U585 (N_585,N_248,N_89);
nand U586 (N_586,In_841,N_283);
xnor U587 (N_587,In_634,In_232);
nor U588 (N_588,N_76,N_311);
nor U589 (N_589,N_335,N_14);
or U590 (N_590,N_30,N_99);
or U591 (N_591,In_22,In_590);
or U592 (N_592,In_563,In_196);
and U593 (N_593,In_675,N_312);
nor U594 (N_594,N_398,N_1);
xnor U595 (N_595,N_65,In_475);
or U596 (N_596,In_378,In_338);
nor U597 (N_597,In_797,In_463);
or U598 (N_598,N_326,In_741);
nor U599 (N_599,In_513,In_856);
nand U600 (N_600,N_583,N_513);
nand U601 (N_601,In_865,N_313);
nor U602 (N_602,N_452,N_336);
nand U603 (N_603,N_565,N_462);
nand U604 (N_604,In_750,N_430);
or U605 (N_605,In_107,N_434);
nor U606 (N_606,N_568,N_377);
and U607 (N_607,N_594,N_586);
or U608 (N_608,N_572,N_280);
nand U609 (N_609,N_484,N_496);
or U610 (N_610,In_887,N_421);
and U611 (N_611,N_559,N_573);
or U612 (N_612,N_284,N_493);
or U613 (N_613,N_234,N_448);
or U614 (N_614,N_401,In_102);
and U615 (N_615,N_590,In_832);
nor U616 (N_616,N_347,N_479);
or U617 (N_617,N_512,In_567);
or U618 (N_618,N_517,N_332);
nand U619 (N_619,N_560,N_90);
nor U620 (N_620,N_48,N_592);
and U621 (N_621,N_245,N_576);
nand U622 (N_622,N_525,N_596);
xor U623 (N_623,N_376,N_548);
nor U624 (N_624,In_30,In_434);
nand U625 (N_625,N_522,N_457);
and U626 (N_626,N_521,N_482);
nor U627 (N_627,N_449,N_403);
and U628 (N_628,In_515,N_411);
nor U629 (N_629,N_467,In_864);
or U630 (N_630,N_515,In_55);
and U631 (N_631,N_540,N_593);
nand U632 (N_632,In_942,N_472);
nor U633 (N_633,N_547,In_79);
or U634 (N_634,N_423,N_386);
nand U635 (N_635,In_934,In_42);
xnor U636 (N_636,N_537,N_581);
nor U637 (N_637,In_525,N_514);
or U638 (N_638,In_782,N_534);
and U639 (N_639,N_541,N_599);
xor U640 (N_640,In_631,In_322);
nor U641 (N_641,N_299,N_429);
or U642 (N_642,In_903,In_154);
nor U643 (N_643,In_971,N_408);
or U644 (N_644,N_334,N_294);
nor U645 (N_645,N_98,N_264);
and U646 (N_646,In_115,N_220);
or U647 (N_647,N_536,In_106);
nor U648 (N_648,N_415,N_529);
nor U649 (N_649,N_439,N_465);
or U650 (N_650,N_340,N_585);
or U651 (N_651,N_556,In_697);
or U652 (N_652,N_563,In_975);
or U653 (N_653,In_37,In_19);
and U654 (N_654,N_531,N_470);
nand U655 (N_655,N_526,In_882);
and U656 (N_656,In_317,N_533);
or U657 (N_657,N_474,N_570);
and U658 (N_658,N_319,N_407);
or U659 (N_659,N_528,N_399);
or U660 (N_660,N_406,N_437);
or U661 (N_661,In_833,N_580);
and U662 (N_662,N_417,N_428);
nor U663 (N_663,In_951,N_498);
or U664 (N_664,N_443,In_773);
nand U665 (N_665,N_499,N_516);
and U666 (N_666,N_431,N_197);
and U667 (N_667,N_450,In_930);
or U668 (N_668,N_400,N_454);
nand U669 (N_669,N_497,N_210);
nor U670 (N_670,N_480,N_509);
nand U671 (N_671,N_487,N_490);
nand U672 (N_672,In_373,N_115);
and U673 (N_673,N_523,N_276);
nor U674 (N_674,In_69,In_92);
or U675 (N_675,N_142,N_469);
and U676 (N_676,N_511,In_347);
or U677 (N_677,N_589,In_787);
or U678 (N_678,N_410,N_549);
nor U679 (N_679,In_811,N_52);
nand U680 (N_680,N_558,In_534);
or U681 (N_681,N_304,N_238);
nor U682 (N_682,N_212,In_770);
and U683 (N_683,N_477,In_506);
or U684 (N_684,In_467,N_577);
xnor U685 (N_685,N_508,N_574);
nand U686 (N_686,In_774,N_422);
nand U687 (N_687,N_552,In_97);
or U688 (N_688,In_889,N_456);
nor U689 (N_689,In_892,N_519);
or U690 (N_690,N_561,N_261);
nor U691 (N_691,N_535,N_253);
xor U692 (N_692,N_564,N_409);
nand U693 (N_693,N_544,N_488);
nor U694 (N_694,N_181,N_328);
nand U695 (N_695,N_475,N_257);
and U696 (N_696,N_494,N_567);
nand U697 (N_697,N_557,In_706);
and U698 (N_698,In_73,N_451);
nor U699 (N_699,N_575,N_8);
nor U700 (N_700,N_507,In_636);
nor U701 (N_701,N_550,N_34);
and U702 (N_702,In_854,In_755);
nand U703 (N_703,N_305,N_351);
nand U704 (N_704,N_379,N_187);
or U705 (N_705,N_538,N_146);
nand U706 (N_706,N_591,N_267);
and U707 (N_707,N_363,N_587);
nand U708 (N_708,N_584,N_143);
or U709 (N_709,N_413,In_794);
or U710 (N_710,N_438,N_588);
nor U711 (N_711,N_566,N_554);
or U712 (N_712,N_343,N_202);
or U713 (N_713,In_711,N_446);
nand U714 (N_714,N_325,N_444);
or U715 (N_715,In_670,N_471);
and U716 (N_716,N_414,N_359);
or U717 (N_717,N_455,In_247);
or U718 (N_718,N_396,N_530);
and U719 (N_719,N_2,N_569);
nor U720 (N_720,N_203,N_504);
or U721 (N_721,In_21,N_579);
and U722 (N_722,In_150,N_476);
or U723 (N_723,N_286,N_491);
nor U724 (N_724,N_453,In_681);
nand U725 (N_725,In_580,N_432);
or U726 (N_726,In_359,In_442);
or U727 (N_727,N_578,In_571);
and U728 (N_728,N_364,N_300);
nand U729 (N_729,In_346,N_425);
nand U730 (N_730,N_464,N_402);
and U731 (N_731,N_354,In_586);
nand U732 (N_732,N_543,N_315);
and U733 (N_733,In_712,N_532);
or U734 (N_734,N_221,N_502);
nand U735 (N_735,N_109,In_158);
and U736 (N_736,N_436,N_468);
or U737 (N_737,In_147,N_404);
and U738 (N_738,N_25,In_26);
nor U739 (N_739,In_14,N_466);
nor U740 (N_740,N_460,N_416);
nor U741 (N_741,N_553,N_222);
nor U742 (N_742,N_268,N_419);
nand U743 (N_743,N_539,In_884);
nor U744 (N_744,N_140,N_216);
nor U745 (N_745,N_495,In_777);
nand U746 (N_746,N_418,N_442);
nor U747 (N_747,N_22,In_242);
nand U748 (N_748,N_16,N_500);
or U749 (N_749,In_245,N_412);
and U750 (N_750,N_154,In_973);
or U751 (N_751,N_381,In_585);
nand U752 (N_752,N_463,N_546);
or U753 (N_753,N_373,N_551);
or U754 (N_754,In_45,N_597);
nor U755 (N_755,N_459,N_518);
and U756 (N_756,In_407,N_433);
or U757 (N_757,In_812,N_524);
nand U758 (N_758,N_458,N_362);
nor U759 (N_759,N_255,In_237);
and U760 (N_760,N_361,N_56);
nor U761 (N_761,N_201,In_224);
and U762 (N_762,N_153,In_431);
nand U763 (N_763,N_542,N_175);
nor U764 (N_764,N_5,N_445);
and U765 (N_765,N_501,N_440);
and U766 (N_766,N_391,N_317);
and U767 (N_767,N_225,In_303);
nor U768 (N_768,In_809,N_287);
and U769 (N_769,In_295,N_55);
and U770 (N_770,N_555,In_38);
nand U771 (N_771,N_486,In_855);
or U772 (N_772,N_243,N_427);
nor U773 (N_773,In_828,In_132);
nand U774 (N_774,N_441,N_189);
nand U775 (N_775,In_175,In_419);
and U776 (N_776,In_717,In_916);
nor U777 (N_777,N_582,N_420);
nand U778 (N_778,N_426,N_562);
nor U779 (N_779,In_581,N_106);
xnor U780 (N_780,In_992,N_503);
or U781 (N_781,N_492,N_520);
xnor U782 (N_782,N_316,N_481);
nand U783 (N_783,In_312,N_485);
nor U784 (N_784,N_478,In_376);
and U785 (N_785,N_473,N_275);
and U786 (N_786,N_4,N_510);
nand U787 (N_787,N_435,N_424);
nand U788 (N_788,N_571,N_306);
and U789 (N_789,N_387,N_595);
nor U790 (N_790,In_151,N_489);
nand U791 (N_791,N_405,N_174);
or U792 (N_792,N_527,N_19);
nor U793 (N_793,N_382,N_505);
or U794 (N_794,In_57,N_545);
xnor U795 (N_795,N_447,N_506);
nor U796 (N_796,In_560,In_259);
or U797 (N_797,In_225,N_598);
nand U798 (N_798,N_128,In_93);
nand U799 (N_799,N_461,N_483);
or U800 (N_800,N_761,N_702);
and U801 (N_801,N_627,N_687);
nor U802 (N_802,N_725,N_683);
nand U803 (N_803,N_607,N_736);
nor U804 (N_804,N_769,N_614);
nor U805 (N_805,N_692,N_704);
nor U806 (N_806,N_643,N_654);
and U807 (N_807,N_726,N_611);
nand U808 (N_808,N_652,N_685);
nor U809 (N_809,N_723,N_688);
nor U810 (N_810,N_783,N_637);
nor U811 (N_811,N_764,N_749);
nand U812 (N_812,N_710,N_631);
nor U813 (N_813,N_779,N_613);
nand U814 (N_814,N_600,N_663);
or U815 (N_815,N_644,N_707);
or U816 (N_816,N_632,N_698);
xor U817 (N_817,N_778,N_605);
and U818 (N_818,N_601,N_750);
nand U819 (N_819,N_691,N_695);
and U820 (N_820,N_732,N_799);
nor U821 (N_821,N_686,N_630);
nor U822 (N_822,N_676,N_672);
nor U823 (N_823,N_673,N_603);
nand U824 (N_824,N_773,N_677);
or U825 (N_825,N_713,N_689);
nor U826 (N_826,N_634,N_739);
or U827 (N_827,N_609,N_712);
and U828 (N_828,N_645,N_638);
nor U829 (N_829,N_765,N_651);
xor U830 (N_830,N_690,N_618);
or U831 (N_831,N_744,N_795);
or U832 (N_832,N_746,N_727);
and U833 (N_833,N_711,N_655);
nand U834 (N_834,N_653,N_706);
and U835 (N_835,N_745,N_766);
or U836 (N_836,N_657,N_714);
nor U837 (N_837,N_756,N_753);
or U838 (N_838,N_741,N_784);
or U839 (N_839,N_716,N_771);
and U840 (N_840,N_738,N_785);
nor U841 (N_841,N_602,N_625);
nand U842 (N_842,N_719,N_722);
or U843 (N_843,N_610,N_742);
nor U844 (N_844,N_735,N_708);
or U845 (N_845,N_640,N_668);
or U846 (N_846,N_791,N_701);
nor U847 (N_847,N_734,N_684);
nor U848 (N_848,N_786,N_767);
nor U849 (N_849,N_670,N_642);
and U850 (N_850,N_620,N_661);
or U851 (N_851,N_737,N_626);
or U852 (N_852,N_649,N_754);
and U853 (N_853,N_720,N_665);
xor U854 (N_854,N_615,N_669);
nand U855 (N_855,N_647,N_790);
nor U856 (N_856,N_758,N_721);
nand U857 (N_857,N_787,N_656);
and U858 (N_858,N_703,N_633);
nor U859 (N_859,N_780,N_662);
and U860 (N_860,N_717,N_659);
nor U861 (N_861,N_635,N_660);
and U862 (N_862,N_666,N_798);
or U863 (N_863,N_733,N_793);
nor U864 (N_864,N_789,N_728);
xnor U865 (N_865,N_748,N_752);
or U866 (N_866,N_762,N_782);
and U867 (N_867,N_792,N_650);
nand U868 (N_868,N_681,N_697);
nand U869 (N_869,N_641,N_622);
nand U870 (N_870,N_604,N_619);
and U871 (N_871,N_608,N_678);
or U872 (N_872,N_731,N_740);
or U873 (N_873,N_664,N_743);
and U874 (N_874,N_694,N_730);
nor U875 (N_875,N_776,N_755);
and U876 (N_876,N_636,N_612);
nand U877 (N_877,N_777,N_718);
and U878 (N_878,N_770,N_705);
and U879 (N_879,N_680,N_629);
or U880 (N_880,N_699,N_763);
nor U881 (N_881,N_675,N_772);
nor U882 (N_882,N_606,N_724);
nor U883 (N_883,N_768,N_646);
xnor U884 (N_884,N_729,N_682);
or U885 (N_885,N_747,N_693);
nor U886 (N_886,N_796,N_667);
and U887 (N_887,N_775,N_628);
or U888 (N_888,N_679,N_624);
nand U889 (N_889,N_757,N_639);
or U890 (N_890,N_751,N_760);
nor U891 (N_891,N_648,N_621);
or U892 (N_892,N_715,N_709);
nor U893 (N_893,N_700,N_759);
xnor U894 (N_894,N_671,N_617);
and U895 (N_895,N_623,N_696);
and U896 (N_896,N_616,N_774);
nor U897 (N_897,N_794,N_658);
and U898 (N_898,N_797,N_788);
xnor U899 (N_899,N_674,N_781);
nand U900 (N_900,N_700,N_673);
nor U901 (N_901,N_686,N_711);
nand U902 (N_902,N_670,N_652);
nor U903 (N_903,N_772,N_771);
xnor U904 (N_904,N_711,N_799);
and U905 (N_905,N_661,N_617);
nand U906 (N_906,N_646,N_728);
nand U907 (N_907,N_628,N_679);
nor U908 (N_908,N_601,N_620);
nor U909 (N_909,N_613,N_624);
nand U910 (N_910,N_751,N_793);
or U911 (N_911,N_667,N_785);
and U912 (N_912,N_614,N_741);
and U913 (N_913,N_725,N_721);
nor U914 (N_914,N_648,N_742);
and U915 (N_915,N_782,N_620);
nand U916 (N_916,N_643,N_661);
nand U917 (N_917,N_761,N_676);
nand U918 (N_918,N_612,N_772);
and U919 (N_919,N_768,N_686);
and U920 (N_920,N_727,N_748);
nor U921 (N_921,N_781,N_616);
and U922 (N_922,N_609,N_645);
or U923 (N_923,N_601,N_682);
nand U924 (N_924,N_680,N_619);
nand U925 (N_925,N_732,N_717);
nor U926 (N_926,N_636,N_666);
and U927 (N_927,N_714,N_696);
nand U928 (N_928,N_715,N_732);
nor U929 (N_929,N_778,N_686);
and U930 (N_930,N_698,N_610);
xnor U931 (N_931,N_699,N_713);
nand U932 (N_932,N_719,N_791);
xnor U933 (N_933,N_709,N_674);
and U934 (N_934,N_640,N_693);
nand U935 (N_935,N_620,N_656);
nor U936 (N_936,N_745,N_710);
and U937 (N_937,N_686,N_667);
nand U938 (N_938,N_721,N_618);
nand U939 (N_939,N_727,N_749);
or U940 (N_940,N_745,N_773);
and U941 (N_941,N_738,N_659);
nand U942 (N_942,N_670,N_768);
and U943 (N_943,N_774,N_692);
nor U944 (N_944,N_613,N_607);
and U945 (N_945,N_603,N_759);
or U946 (N_946,N_680,N_794);
nor U947 (N_947,N_765,N_610);
nand U948 (N_948,N_786,N_732);
or U949 (N_949,N_623,N_766);
and U950 (N_950,N_605,N_767);
or U951 (N_951,N_663,N_788);
or U952 (N_952,N_771,N_697);
nand U953 (N_953,N_730,N_734);
or U954 (N_954,N_744,N_663);
nor U955 (N_955,N_762,N_676);
xor U956 (N_956,N_733,N_720);
and U957 (N_957,N_713,N_690);
nand U958 (N_958,N_718,N_655);
nor U959 (N_959,N_712,N_628);
and U960 (N_960,N_793,N_766);
or U961 (N_961,N_778,N_770);
or U962 (N_962,N_759,N_722);
nand U963 (N_963,N_683,N_729);
nor U964 (N_964,N_640,N_665);
and U965 (N_965,N_700,N_778);
nor U966 (N_966,N_695,N_757);
nor U967 (N_967,N_740,N_783);
nor U968 (N_968,N_624,N_716);
nand U969 (N_969,N_770,N_654);
or U970 (N_970,N_746,N_768);
nand U971 (N_971,N_694,N_717);
nand U972 (N_972,N_722,N_665);
or U973 (N_973,N_777,N_784);
nand U974 (N_974,N_727,N_620);
or U975 (N_975,N_752,N_783);
or U976 (N_976,N_600,N_634);
or U977 (N_977,N_795,N_626);
nand U978 (N_978,N_700,N_620);
xnor U979 (N_979,N_766,N_724);
or U980 (N_980,N_673,N_727);
nand U981 (N_981,N_685,N_610);
nand U982 (N_982,N_673,N_729);
and U983 (N_983,N_680,N_678);
nand U984 (N_984,N_785,N_646);
nand U985 (N_985,N_707,N_709);
and U986 (N_986,N_768,N_699);
nand U987 (N_987,N_711,N_759);
and U988 (N_988,N_672,N_765);
and U989 (N_989,N_619,N_665);
or U990 (N_990,N_761,N_626);
nand U991 (N_991,N_748,N_703);
and U992 (N_992,N_601,N_676);
or U993 (N_993,N_741,N_607);
nand U994 (N_994,N_742,N_624);
and U995 (N_995,N_697,N_650);
nor U996 (N_996,N_680,N_719);
nor U997 (N_997,N_621,N_773);
and U998 (N_998,N_739,N_669);
nor U999 (N_999,N_669,N_797);
and U1000 (N_1000,N_941,N_867);
nor U1001 (N_1001,N_895,N_850);
or U1002 (N_1002,N_959,N_969);
or U1003 (N_1003,N_978,N_990);
nor U1004 (N_1004,N_858,N_911);
and U1005 (N_1005,N_920,N_957);
nor U1006 (N_1006,N_890,N_902);
and U1007 (N_1007,N_862,N_965);
nor U1008 (N_1008,N_861,N_886);
and U1009 (N_1009,N_879,N_853);
nand U1010 (N_1010,N_881,N_851);
and U1011 (N_1011,N_952,N_975);
nand U1012 (N_1012,N_817,N_918);
or U1013 (N_1013,N_982,N_874);
and U1014 (N_1014,N_909,N_905);
xor U1015 (N_1015,N_926,N_958);
or U1016 (N_1016,N_806,N_816);
nand U1017 (N_1017,N_838,N_908);
nand U1018 (N_1018,N_876,N_972);
nand U1019 (N_1019,N_812,N_821);
nor U1020 (N_1020,N_855,N_822);
nor U1021 (N_1021,N_996,N_930);
nand U1022 (N_1022,N_814,N_983);
or U1023 (N_1023,N_848,N_942);
nand U1024 (N_1024,N_877,N_882);
and U1025 (N_1025,N_875,N_927);
and U1026 (N_1026,N_832,N_960);
xnor U1027 (N_1027,N_809,N_894);
xnor U1028 (N_1028,N_906,N_924);
nor U1029 (N_1029,N_815,N_897);
nor U1030 (N_1030,N_863,N_804);
nand U1031 (N_1031,N_981,N_846);
nand U1032 (N_1032,N_864,N_899);
or U1033 (N_1033,N_950,N_992);
nand U1034 (N_1034,N_998,N_868);
and U1035 (N_1035,N_961,N_834);
nand U1036 (N_1036,N_811,N_878);
nand U1037 (N_1037,N_896,N_953);
or U1038 (N_1038,N_844,N_968);
and U1039 (N_1039,N_948,N_856);
or U1040 (N_1040,N_800,N_839);
or U1041 (N_1041,N_980,N_921);
nand U1042 (N_1042,N_873,N_925);
nand U1043 (N_1043,N_987,N_944);
nor U1044 (N_1044,N_813,N_802);
and U1045 (N_1045,N_956,N_966);
and U1046 (N_1046,N_826,N_912);
nand U1047 (N_1047,N_887,N_993);
or U1048 (N_1048,N_847,N_820);
nand U1049 (N_1049,N_986,N_995);
and U1050 (N_1050,N_999,N_989);
nor U1051 (N_1051,N_932,N_922);
xnor U1052 (N_1052,N_801,N_964);
and U1053 (N_1053,N_955,N_841);
xnor U1054 (N_1054,N_833,N_971);
nand U1055 (N_1055,N_883,N_892);
nor U1056 (N_1056,N_829,N_880);
and U1057 (N_1057,N_974,N_991);
nor U1058 (N_1058,N_836,N_940);
and U1059 (N_1059,N_891,N_939);
or U1060 (N_1060,N_962,N_977);
and U1061 (N_1061,N_818,N_949);
and U1062 (N_1062,N_866,N_963);
nand U1063 (N_1063,N_951,N_945);
or U1064 (N_1064,N_916,N_943);
nor U1065 (N_1065,N_828,N_973);
and U1066 (N_1066,N_985,N_935);
or U1067 (N_1067,N_937,N_825);
and U1068 (N_1068,N_888,N_917);
or U1069 (N_1069,N_857,N_859);
or U1070 (N_1070,N_840,N_913);
or U1071 (N_1071,N_854,N_903);
and U1072 (N_1072,N_823,N_946);
and U1073 (N_1073,N_967,N_872);
nor U1074 (N_1074,N_810,N_984);
nand U1075 (N_1075,N_900,N_947);
nand U1076 (N_1076,N_842,N_919);
or U1077 (N_1077,N_914,N_871);
xor U1078 (N_1078,N_928,N_931);
nor U1079 (N_1079,N_893,N_852);
nor U1080 (N_1080,N_845,N_805);
nand U1081 (N_1081,N_819,N_827);
nor U1082 (N_1082,N_830,N_869);
and U1083 (N_1083,N_865,N_835);
nor U1084 (N_1084,N_933,N_929);
nand U1085 (N_1085,N_889,N_988);
and U1086 (N_1086,N_970,N_849);
nand U1087 (N_1087,N_954,N_831);
nor U1088 (N_1088,N_807,N_910);
nor U1089 (N_1089,N_923,N_904);
xnor U1090 (N_1090,N_901,N_808);
or U1091 (N_1091,N_997,N_885);
or U1092 (N_1092,N_803,N_994);
xnor U1093 (N_1093,N_898,N_934);
nand U1094 (N_1094,N_976,N_824);
or U1095 (N_1095,N_837,N_938);
or U1096 (N_1096,N_915,N_860);
nor U1097 (N_1097,N_870,N_843);
nand U1098 (N_1098,N_884,N_907);
nand U1099 (N_1099,N_979,N_936);
nor U1100 (N_1100,N_949,N_992);
and U1101 (N_1101,N_846,N_906);
nor U1102 (N_1102,N_800,N_874);
nor U1103 (N_1103,N_898,N_997);
nand U1104 (N_1104,N_877,N_893);
nor U1105 (N_1105,N_996,N_850);
nor U1106 (N_1106,N_906,N_881);
nand U1107 (N_1107,N_821,N_978);
and U1108 (N_1108,N_838,N_889);
or U1109 (N_1109,N_841,N_974);
or U1110 (N_1110,N_962,N_828);
nand U1111 (N_1111,N_919,N_967);
or U1112 (N_1112,N_947,N_811);
nor U1113 (N_1113,N_881,N_829);
and U1114 (N_1114,N_875,N_931);
and U1115 (N_1115,N_904,N_912);
and U1116 (N_1116,N_853,N_982);
and U1117 (N_1117,N_983,N_913);
nor U1118 (N_1118,N_868,N_937);
or U1119 (N_1119,N_947,N_834);
nor U1120 (N_1120,N_947,N_868);
or U1121 (N_1121,N_864,N_830);
nor U1122 (N_1122,N_835,N_855);
and U1123 (N_1123,N_927,N_902);
or U1124 (N_1124,N_800,N_892);
nor U1125 (N_1125,N_915,N_872);
nand U1126 (N_1126,N_942,N_813);
or U1127 (N_1127,N_992,N_813);
nand U1128 (N_1128,N_979,N_805);
and U1129 (N_1129,N_975,N_962);
nand U1130 (N_1130,N_924,N_883);
nand U1131 (N_1131,N_808,N_821);
or U1132 (N_1132,N_831,N_957);
nor U1133 (N_1133,N_858,N_826);
and U1134 (N_1134,N_822,N_946);
xnor U1135 (N_1135,N_946,N_988);
nand U1136 (N_1136,N_993,N_918);
nor U1137 (N_1137,N_874,N_904);
or U1138 (N_1138,N_847,N_904);
and U1139 (N_1139,N_952,N_803);
nor U1140 (N_1140,N_841,N_884);
and U1141 (N_1141,N_964,N_979);
nor U1142 (N_1142,N_873,N_805);
nand U1143 (N_1143,N_836,N_863);
nor U1144 (N_1144,N_961,N_995);
nor U1145 (N_1145,N_808,N_957);
nand U1146 (N_1146,N_965,N_883);
nand U1147 (N_1147,N_901,N_846);
and U1148 (N_1148,N_959,N_945);
or U1149 (N_1149,N_849,N_851);
nor U1150 (N_1150,N_868,N_933);
nor U1151 (N_1151,N_850,N_891);
nor U1152 (N_1152,N_900,N_876);
nor U1153 (N_1153,N_892,N_841);
and U1154 (N_1154,N_926,N_950);
or U1155 (N_1155,N_953,N_993);
and U1156 (N_1156,N_984,N_815);
nor U1157 (N_1157,N_846,N_873);
and U1158 (N_1158,N_926,N_949);
or U1159 (N_1159,N_894,N_832);
or U1160 (N_1160,N_894,N_959);
and U1161 (N_1161,N_954,N_805);
and U1162 (N_1162,N_864,N_850);
or U1163 (N_1163,N_883,N_893);
nor U1164 (N_1164,N_846,N_988);
nor U1165 (N_1165,N_933,N_974);
nor U1166 (N_1166,N_833,N_947);
and U1167 (N_1167,N_801,N_955);
and U1168 (N_1168,N_995,N_923);
or U1169 (N_1169,N_840,N_876);
nor U1170 (N_1170,N_957,N_924);
nand U1171 (N_1171,N_860,N_828);
nor U1172 (N_1172,N_971,N_964);
and U1173 (N_1173,N_900,N_930);
nand U1174 (N_1174,N_811,N_834);
nor U1175 (N_1175,N_822,N_902);
nor U1176 (N_1176,N_945,N_985);
nand U1177 (N_1177,N_921,N_961);
nor U1178 (N_1178,N_872,N_863);
nand U1179 (N_1179,N_823,N_949);
and U1180 (N_1180,N_982,N_850);
and U1181 (N_1181,N_862,N_847);
or U1182 (N_1182,N_893,N_966);
nor U1183 (N_1183,N_800,N_847);
nand U1184 (N_1184,N_877,N_924);
or U1185 (N_1185,N_831,N_981);
nand U1186 (N_1186,N_940,N_956);
and U1187 (N_1187,N_975,N_954);
nand U1188 (N_1188,N_975,N_821);
nand U1189 (N_1189,N_823,N_869);
or U1190 (N_1190,N_956,N_845);
nor U1191 (N_1191,N_880,N_916);
nor U1192 (N_1192,N_828,N_997);
and U1193 (N_1193,N_868,N_972);
nand U1194 (N_1194,N_947,N_872);
and U1195 (N_1195,N_802,N_818);
and U1196 (N_1196,N_887,N_999);
and U1197 (N_1197,N_898,N_888);
nor U1198 (N_1198,N_935,N_806);
nor U1199 (N_1199,N_974,N_948);
nand U1200 (N_1200,N_1027,N_1036);
nor U1201 (N_1201,N_1149,N_1007);
nor U1202 (N_1202,N_1015,N_1024);
or U1203 (N_1203,N_1099,N_1054);
nor U1204 (N_1204,N_1004,N_1079);
nor U1205 (N_1205,N_1044,N_1063);
or U1206 (N_1206,N_1093,N_1077);
and U1207 (N_1207,N_1033,N_1194);
nor U1208 (N_1208,N_1069,N_1083);
or U1209 (N_1209,N_1096,N_1135);
or U1210 (N_1210,N_1049,N_1037);
or U1211 (N_1211,N_1086,N_1022);
or U1212 (N_1212,N_1104,N_1160);
and U1213 (N_1213,N_1188,N_1140);
or U1214 (N_1214,N_1006,N_1182);
nand U1215 (N_1215,N_1047,N_1155);
or U1216 (N_1216,N_1040,N_1073);
nand U1217 (N_1217,N_1020,N_1081);
or U1218 (N_1218,N_1090,N_1060);
or U1219 (N_1219,N_1137,N_1108);
nand U1220 (N_1220,N_1016,N_1088);
and U1221 (N_1221,N_1032,N_1176);
nor U1222 (N_1222,N_1118,N_1117);
and U1223 (N_1223,N_1144,N_1112);
nand U1224 (N_1224,N_1165,N_1065);
nand U1225 (N_1225,N_1008,N_1166);
or U1226 (N_1226,N_1197,N_1168);
and U1227 (N_1227,N_1130,N_1121);
nor U1228 (N_1228,N_1053,N_1179);
nand U1229 (N_1229,N_1046,N_1116);
and U1230 (N_1230,N_1074,N_1119);
and U1231 (N_1231,N_1031,N_1000);
or U1232 (N_1232,N_1056,N_1156);
xnor U1233 (N_1233,N_1068,N_1059);
nor U1234 (N_1234,N_1126,N_1014);
nor U1235 (N_1235,N_1186,N_1002);
nand U1236 (N_1236,N_1064,N_1180);
and U1237 (N_1237,N_1185,N_1174);
nand U1238 (N_1238,N_1178,N_1043);
xnor U1239 (N_1239,N_1010,N_1092);
or U1240 (N_1240,N_1061,N_1013);
nor U1241 (N_1241,N_1017,N_1019);
nor U1242 (N_1242,N_1038,N_1162);
xnor U1243 (N_1243,N_1091,N_1183);
and U1244 (N_1244,N_1184,N_1175);
or U1245 (N_1245,N_1058,N_1035);
nor U1246 (N_1246,N_1158,N_1152);
nand U1247 (N_1247,N_1127,N_1018);
or U1248 (N_1248,N_1164,N_1173);
and U1249 (N_1249,N_1029,N_1101);
nand U1250 (N_1250,N_1028,N_1089);
or U1251 (N_1251,N_1169,N_1134);
nor U1252 (N_1252,N_1129,N_1196);
or U1253 (N_1253,N_1005,N_1094);
or U1254 (N_1254,N_1138,N_1041);
nand U1255 (N_1255,N_1153,N_1095);
and U1256 (N_1256,N_1071,N_1170);
nand U1257 (N_1257,N_1132,N_1021);
or U1258 (N_1258,N_1111,N_1026);
xnor U1259 (N_1259,N_1193,N_1115);
or U1260 (N_1260,N_1191,N_1039);
or U1261 (N_1261,N_1114,N_1051);
or U1262 (N_1262,N_1192,N_1190);
xor U1263 (N_1263,N_1082,N_1098);
or U1264 (N_1264,N_1177,N_1009);
or U1265 (N_1265,N_1151,N_1199);
and U1266 (N_1266,N_1122,N_1030);
and U1267 (N_1267,N_1034,N_1084);
nor U1268 (N_1268,N_1163,N_1001);
nor U1269 (N_1269,N_1146,N_1011);
and U1270 (N_1270,N_1105,N_1085);
or U1271 (N_1271,N_1110,N_1159);
or U1272 (N_1272,N_1150,N_1147);
nor U1273 (N_1273,N_1025,N_1131);
nand U1274 (N_1274,N_1045,N_1070);
nor U1275 (N_1275,N_1120,N_1198);
nand U1276 (N_1276,N_1042,N_1050);
nand U1277 (N_1277,N_1076,N_1055);
nor U1278 (N_1278,N_1113,N_1154);
and U1279 (N_1279,N_1125,N_1145);
nor U1280 (N_1280,N_1133,N_1078);
and U1281 (N_1281,N_1181,N_1057);
or U1282 (N_1282,N_1103,N_1167);
nand U1283 (N_1283,N_1066,N_1171);
and U1284 (N_1284,N_1143,N_1172);
xnor U1285 (N_1285,N_1012,N_1067);
nor U1286 (N_1286,N_1023,N_1195);
and U1287 (N_1287,N_1080,N_1062);
nand U1288 (N_1288,N_1141,N_1139);
and U1289 (N_1289,N_1187,N_1189);
and U1290 (N_1290,N_1052,N_1109);
xor U1291 (N_1291,N_1148,N_1087);
or U1292 (N_1292,N_1100,N_1123);
and U1293 (N_1293,N_1124,N_1048);
nand U1294 (N_1294,N_1072,N_1142);
and U1295 (N_1295,N_1128,N_1003);
nand U1296 (N_1296,N_1157,N_1075);
nor U1297 (N_1297,N_1107,N_1136);
nor U1298 (N_1298,N_1102,N_1106);
nand U1299 (N_1299,N_1161,N_1097);
and U1300 (N_1300,N_1070,N_1121);
and U1301 (N_1301,N_1070,N_1095);
and U1302 (N_1302,N_1083,N_1054);
or U1303 (N_1303,N_1018,N_1095);
nand U1304 (N_1304,N_1068,N_1161);
and U1305 (N_1305,N_1125,N_1134);
and U1306 (N_1306,N_1057,N_1193);
nand U1307 (N_1307,N_1057,N_1011);
nor U1308 (N_1308,N_1168,N_1029);
nand U1309 (N_1309,N_1145,N_1031);
or U1310 (N_1310,N_1051,N_1108);
and U1311 (N_1311,N_1187,N_1154);
and U1312 (N_1312,N_1102,N_1180);
or U1313 (N_1313,N_1157,N_1084);
nand U1314 (N_1314,N_1051,N_1073);
and U1315 (N_1315,N_1111,N_1144);
nor U1316 (N_1316,N_1181,N_1097);
or U1317 (N_1317,N_1152,N_1008);
nand U1318 (N_1318,N_1078,N_1057);
or U1319 (N_1319,N_1084,N_1038);
nand U1320 (N_1320,N_1107,N_1074);
and U1321 (N_1321,N_1122,N_1057);
nor U1322 (N_1322,N_1026,N_1179);
or U1323 (N_1323,N_1069,N_1053);
or U1324 (N_1324,N_1081,N_1038);
or U1325 (N_1325,N_1119,N_1071);
or U1326 (N_1326,N_1143,N_1030);
nor U1327 (N_1327,N_1157,N_1022);
or U1328 (N_1328,N_1154,N_1057);
or U1329 (N_1329,N_1075,N_1114);
and U1330 (N_1330,N_1195,N_1096);
and U1331 (N_1331,N_1036,N_1183);
nor U1332 (N_1332,N_1167,N_1075);
nor U1333 (N_1333,N_1007,N_1062);
or U1334 (N_1334,N_1101,N_1122);
and U1335 (N_1335,N_1024,N_1180);
nand U1336 (N_1336,N_1052,N_1120);
or U1337 (N_1337,N_1114,N_1191);
xor U1338 (N_1338,N_1019,N_1132);
nand U1339 (N_1339,N_1080,N_1185);
nor U1340 (N_1340,N_1179,N_1105);
or U1341 (N_1341,N_1136,N_1040);
nand U1342 (N_1342,N_1120,N_1193);
nand U1343 (N_1343,N_1129,N_1070);
nor U1344 (N_1344,N_1125,N_1168);
or U1345 (N_1345,N_1077,N_1005);
nor U1346 (N_1346,N_1168,N_1127);
or U1347 (N_1347,N_1017,N_1117);
nor U1348 (N_1348,N_1039,N_1169);
nor U1349 (N_1349,N_1140,N_1042);
or U1350 (N_1350,N_1018,N_1040);
nor U1351 (N_1351,N_1157,N_1138);
and U1352 (N_1352,N_1172,N_1023);
nand U1353 (N_1353,N_1103,N_1011);
nor U1354 (N_1354,N_1160,N_1074);
or U1355 (N_1355,N_1047,N_1028);
nand U1356 (N_1356,N_1147,N_1112);
or U1357 (N_1357,N_1046,N_1013);
and U1358 (N_1358,N_1077,N_1197);
nand U1359 (N_1359,N_1043,N_1087);
nand U1360 (N_1360,N_1129,N_1180);
nand U1361 (N_1361,N_1178,N_1172);
or U1362 (N_1362,N_1041,N_1157);
and U1363 (N_1363,N_1128,N_1151);
or U1364 (N_1364,N_1125,N_1141);
nand U1365 (N_1365,N_1092,N_1193);
or U1366 (N_1366,N_1142,N_1158);
nor U1367 (N_1367,N_1083,N_1096);
and U1368 (N_1368,N_1178,N_1008);
and U1369 (N_1369,N_1160,N_1154);
and U1370 (N_1370,N_1052,N_1074);
and U1371 (N_1371,N_1107,N_1187);
and U1372 (N_1372,N_1033,N_1118);
nor U1373 (N_1373,N_1004,N_1111);
nand U1374 (N_1374,N_1140,N_1088);
nand U1375 (N_1375,N_1183,N_1142);
nand U1376 (N_1376,N_1193,N_1104);
nand U1377 (N_1377,N_1161,N_1114);
or U1378 (N_1378,N_1199,N_1008);
or U1379 (N_1379,N_1077,N_1182);
nand U1380 (N_1380,N_1031,N_1106);
and U1381 (N_1381,N_1130,N_1166);
or U1382 (N_1382,N_1055,N_1113);
nor U1383 (N_1383,N_1082,N_1109);
or U1384 (N_1384,N_1118,N_1031);
nor U1385 (N_1385,N_1129,N_1095);
nand U1386 (N_1386,N_1076,N_1179);
nor U1387 (N_1387,N_1074,N_1076);
or U1388 (N_1388,N_1030,N_1048);
nand U1389 (N_1389,N_1015,N_1198);
or U1390 (N_1390,N_1198,N_1139);
and U1391 (N_1391,N_1154,N_1198);
nor U1392 (N_1392,N_1107,N_1071);
nor U1393 (N_1393,N_1075,N_1015);
and U1394 (N_1394,N_1198,N_1025);
nor U1395 (N_1395,N_1090,N_1193);
nand U1396 (N_1396,N_1053,N_1079);
and U1397 (N_1397,N_1028,N_1138);
or U1398 (N_1398,N_1026,N_1070);
nor U1399 (N_1399,N_1006,N_1168);
nor U1400 (N_1400,N_1253,N_1203);
nor U1401 (N_1401,N_1282,N_1367);
or U1402 (N_1402,N_1278,N_1284);
nand U1403 (N_1403,N_1246,N_1239);
or U1404 (N_1404,N_1262,N_1204);
nor U1405 (N_1405,N_1382,N_1306);
nand U1406 (N_1406,N_1290,N_1329);
or U1407 (N_1407,N_1370,N_1383);
or U1408 (N_1408,N_1327,N_1345);
xor U1409 (N_1409,N_1321,N_1254);
and U1410 (N_1410,N_1311,N_1332);
nand U1411 (N_1411,N_1341,N_1315);
and U1412 (N_1412,N_1309,N_1368);
nand U1413 (N_1413,N_1335,N_1344);
nand U1414 (N_1414,N_1399,N_1364);
nor U1415 (N_1415,N_1219,N_1376);
nor U1416 (N_1416,N_1355,N_1291);
nor U1417 (N_1417,N_1387,N_1287);
nor U1418 (N_1418,N_1374,N_1285);
and U1419 (N_1419,N_1277,N_1273);
or U1420 (N_1420,N_1233,N_1221);
or U1421 (N_1421,N_1371,N_1396);
and U1422 (N_1422,N_1214,N_1394);
nand U1423 (N_1423,N_1350,N_1234);
or U1424 (N_1424,N_1385,N_1244);
nor U1425 (N_1425,N_1328,N_1207);
nor U1426 (N_1426,N_1237,N_1236);
nor U1427 (N_1427,N_1378,N_1210);
or U1428 (N_1428,N_1353,N_1257);
nand U1429 (N_1429,N_1208,N_1326);
or U1430 (N_1430,N_1361,N_1238);
and U1431 (N_1431,N_1227,N_1302);
or U1432 (N_1432,N_1331,N_1389);
nand U1433 (N_1433,N_1354,N_1220);
or U1434 (N_1434,N_1242,N_1314);
or U1435 (N_1435,N_1252,N_1232);
nor U1436 (N_1436,N_1395,N_1325);
or U1437 (N_1437,N_1338,N_1248);
or U1438 (N_1438,N_1391,N_1323);
nor U1439 (N_1439,N_1366,N_1264);
or U1440 (N_1440,N_1322,N_1348);
or U1441 (N_1441,N_1343,N_1258);
or U1442 (N_1442,N_1243,N_1272);
nor U1443 (N_1443,N_1360,N_1263);
xor U1444 (N_1444,N_1283,N_1268);
nand U1445 (N_1445,N_1212,N_1205);
and U1446 (N_1446,N_1265,N_1267);
nand U1447 (N_1447,N_1280,N_1351);
nand U1448 (N_1448,N_1392,N_1365);
xnor U1449 (N_1449,N_1393,N_1359);
and U1450 (N_1450,N_1336,N_1206);
nand U1451 (N_1451,N_1226,N_1320);
and U1452 (N_1452,N_1307,N_1379);
or U1453 (N_1453,N_1358,N_1384);
nor U1454 (N_1454,N_1362,N_1346);
nand U1455 (N_1455,N_1276,N_1299);
or U1456 (N_1456,N_1223,N_1398);
xnor U1457 (N_1457,N_1303,N_1304);
nor U1458 (N_1458,N_1289,N_1241);
nand U1459 (N_1459,N_1380,N_1308);
and U1460 (N_1460,N_1247,N_1286);
or U1461 (N_1461,N_1349,N_1255);
nand U1462 (N_1462,N_1261,N_1375);
nor U1463 (N_1463,N_1270,N_1347);
or U1464 (N_1464,N_1240,N_1319);
nor U1465 (N_1465,N_1386,N_1269);
nor U1466 (N_1466,N_1259,N_1313);
nand U1467 (N_1467,N_1224,N_1275);
nand U1468 (N_1468,N_1305,N_1213);
xnor U1469 (N_1469,N_1266,N_1300);
nor U1470 (N_1470,N_1388,N_1377);
nor U1471 (N_1471,N_1217,N_1340);
or U1472 (N_1472,N_1324,N_1256);
nor U1473 (N_1473,N_1294,N_1373);
or U1474 (N_1474,N_1352,N_1317);
or U1475 (N_1475,N_1249,N_1229);
or U1476 (N_1476,N_1369,N_1333);
and U1477 (N_1477,N_1200,N_1231);
nand U1478 (N_1478,N_1372,N_1312);
and U1479 (N_1479,N_1260,N_1281);
nand U1480 (N_1480,N_1250,N_1209);
nand U1481 (N_1481,N_1296,N_1216);
nand U1482 (N_1482,N_1228,N_1235);
or U1483 (N_1483,N_1222,N_1288);
or U1484 (N_1484,N_1339,N_1301);
nor U1485 (N_1485,N_1357,N_1202);
nand U1486 (N_1486,N_1356,N_1211);
nor U1487 (N_1487,N_1293,N_1245);
nor U1488 (N_1488,N_1337,N_1215);
nor U1489 (N_1489,N_1251,N_1295);
and U1490 (N_1490,N_1274,N_1230);
or U1491 (N_1491,N_1342,N_1297);
nor U1492 (N_1492,N_1397,N_1279);
nand U1493 (N_1493,N_1316,N_1330);
and U1494 (N_1494,N_1201,N_1292);
nor U1495 (N_1495,N_1334,N_1310);
or U1496 (N_1496,N_1225,N_1271);
or U1497 (N_1497,N_1363,N_1390);
nand U1498 (N_1498,N_1318,N_1298);
nor U1499 (N_1499,N_1218,N_1381);
and U1500 (N_1500,N_1338,N_1219);
and U1501 (N_1501,N_1396,N_1356);
and U1502 (N_1502,N_1268,N_1351);
or U1503 (N_1503,N_1379,N_1237);
nor U1504 (N_1504,N_1330,N_1355);
nor U1505 (N_1505,N_1233,N_1379);
or U1506 (N_1506,N_1265,N_1241);
or U1507 (N_1507,N_1283,N_1289);
xor U1508 (N_1508,N_1366,N_1234);
and U1509 (N_1509,N_1228,N_1251);
or U1510 (N_1510,N_1281,N_1276);
xnor U1511 (N_1511,N_1360,N_1298);
and U1512 (N_1512,N_1393,N_1263);
nand U1513 (N_1513,N_1326,N_1330);
nand U1514 (N_1514,N_1372,N_1343);
and U1515 (N_1515,N_1385,N_1390);
and U1516 (N_1516,N_1278,N_1360);
nor U1517 (N_1517,N_1314,N_1215);
and U1518 (N_1518,N_1328,N_1336);
and U1519 (N_1519,N_1238,N_1210);
or U1520 (N_1520,N_1229,N_1320);
nor U1521 (N_1521,N_1394,N_1370);
nor U1522 (N_1522,N_1321,N_1275);
or U1523 (N_1523,N_1297,N_1223);
or U1524 (N_1524,N_1337,N_1209);
nand U1525 (N_1525,N_1283,N_1292);
xor U1526 (N_1526,N_1224,N_1238);
and U1527 (N_1527,N_1249,N_1226);
or U1528 (N_1528,N_1321,N_1258);
nand U1529 (N_1529,N_1227,N_1317);
and U1530 (N_1530,N_1221,N_1247);
nand U1531 (N_1531,N_1379,N_1212);
and U1532 (N_1532,N_1295,N_1321);
nor U1533 (N_1533,N_1320,N_1231);
and U1534 (N_1534,N_1256,N_1343);
or U1535 (N_1535,N_1288,N_1363);
and U1536 (N_1536,N_1282,N_1301);
or U1537 (N_1537,N_1335,N_1362);
or U1538 (N_1538,N_1298,N_1306);
nor U1539 (N_1539,N_1303,N_1206);
nand U1540 (N_1540,N_1383,N_1363);
and U1541 (N_1541,N_1211,N_1207);
nand U1542 (N_1542,N_1212,N_1342);
or U1543 (N_1543,N_1368,N_1380);
or U1544 (N_1544,N_1397,N_1212);
and U1545 (N_1545,N_1224,N_1241);
nor U1546 (N_1546,N_1269,N_1316);
or U1547 (N_1547,N_1210,N_1259);
or U1548 (N_1548,N_1330,N_1204);
nor U1549 (N_1549,N_1236,N_1311);
nor U1550 (N_1550,N_1226,N_1391);
nor U1551 (N_1551,N_1327,N_1265);
or U1552 (N_1552,N_1312,N_1351);
nand U1553 (N_1553,N_1328,N_1259);
nor U1554 (N_1554,N_1351,N_1230);
or U1555 (N_1555,N_1339,N_1308);
nand U1556 (N_1556,N_1369,N_1277);
or U1557 (N_1557,N_1206,N_1370);
and U1558 (N_1558,N_1233,N_1282);
nor U1559 (N_1559,N_1349,N_1251);
nor U1560 (N_1560,N_1320,N_1344);
nand U1561 (N_1561,N_1305,N_1363);
nor U1562 (N_1562,N_1324,N_1340);
nand U1563 (N_1563,N_1325,N_1373);
nor U1564 (N_1564,N_1363,N_1273);
nand U1565 (N_1565,N_1215,N_1370);
nor U1566 (N_1566,N_1338,N_1281);
and U1567 (N_1567,N_1385,N_1320);
nand U1568 (N_1568,N_1208,N_1217);
nand U1569 (N_1569,N_1267,N_1275);
nand U1570 (N_1570,N_1242,N_1367);
and U1571 (N_1571,N_1213,N_1233);
or U1572 (N_1572,N_1309,N_1282);
and U1573 (N_1573,N_1223,N_1218);
and U1574 (N_1574,N_1208,N_1256);
nand U1575 (N_1575,N_1295,N_1316);
nor U1576 (N_1576,N_1225,N_1279);
nor U1577 (N_1577,N_1219,N_1252);
and U1578 (N_1578,N_1366,N_1392);
or U1579 (N_1579,N_1337,N_1380);
or U1580 (N_1580,N_1344,N_1346);
nand U1581 (N_1581,N_1258,N_1297);
and U1582 (N_1582,N_1233,N_1353);
nor U1583 (N_1583,N_1354,N_1254);
or U1584 (N_1584,N_1241,N_1232);
and U1585 (N_1585,N_1318,N_1202);
nor U1586 (N_1586,N_1354,N_1304);
nand U1587 (N_1587,N_1238,N_1229);
and U1588 (N_1588,N_1350,N_1397);
and U1589 (N_1589,N_1344,N_1216);
nor U1590 (N_1590,N_1278,N_1293);
or U1591 (N_1591,N_1241,N_1207);
nand U1592 (N_1592,N_1296,N_1300);
nand U1593 (N_1593,N_1311,N_1389);
and U1594 (N_1594,N_1364,N_1219);
or U1595 (N_1595,N_1279,N_1286);
or U1596 (N_1596,N_1300,N_1356);
nand U1597 (N_1597,N_1342,N_1210);
nor U1598 (N_1598,N_1232,N_1203);
or U1599 (N_1599,N_1261,N_1212);
nor U1600 (N_1600,N_1459,N_1508);
or U1601 (N_1601,N_1443,N_1503);
and U1602 (N_1602,N_1436,N_1540);
or U1603 (N_1603,N_1546,N_1406);
nor U1604 (N_1604,N_1589,N_1556);
nor U1605 (N_1605,N_1599,N_1451);
nand U1606 (N_1606,N_1563,N_1438);
or U1607 (N_1607,N_1554,N_1410);
nor U1608 (N_1608,N_1463,N_1550);
nor U1609 (N_1609,N_1448,N_1577);
or U1610 (N_1610,N_1455,N_1560);
nand U1611 (N_1611,N_1505,N_1502);
nand U1612 (N_1612,N_1529,N_1452);
nor U1613 (N_1613,N_1524,N_1461);
nor U1614 (N_1614,N_1402,N_1581);
xnor U1615 (N_1615,N_1594,N_1500);
and U1616 (N_1616,N_1439,N_1471);
xor U1617 (N_1617,N_1535,N_1539);
xnor U1618 (N_1618,N_1458,N_1591);
xnor U1619 (N_1619,N_1430,N_1510);
or U1620 (N_1620,N_1479,N_1475);
or U1621 (N_1621,N_1498,N_1568);
or U1622 (N_1622,N_1584,N_1570);
or U1623 (N_1623,N_1553,N_1483);
nand U1624 (N_1624,N_1499,N_1480);
or U1625 (N_1625,N_1476,N_1428);
nor U1626 (N_1626,N_1543,N_1544);
nand U1627 (N_1627,N_1495,N_1561);
or U1628 (N_1628,N_1464,N_1460);
nor U1629 (N_1629,N_1533,N_1442);
nand U1630 (N_1630,N_1401,N_1441);
nand U1631 (N_1631,N_1413,N_1579);
nor U1632 (N_1632,N_1588,N_1587);
nor U1633 (N_1633,N_1528,N_1586);
or U1634 (N_1634,N_1456,N_1467);
nor U1635 (N_1635,N_1478,N_1582);
nor U1636 (N_1636,N_1477,N_1523);
nand U1637 (N_1637,N_1411,N_1538);
or U1638 (N_1638,N_1468,N_1519);
nor U1639 (N_1639,N_1501,N_1592);
nor U1640 (N_1640,N_1527,N_1565);
nand U1641 (N_1641,N_1403,N_1444);
or U1642 (N_1642,N_1525,N_1492);
nand U1643 (N_1643,N_1494,N_1427);
and U1644 (N_1644,N_1432,N_1558);
or U1645 (N_1645,N_1429,N_1437);
and U1646 (N_1646,N_1440,N_1484);
nor U1647 (N_1647,N_1555,N_1578);
nand U1648 (N_1648,N_1512,N_1418);
or U1649 (N_1649,N_1474,N_1504);
xor U1650 (N_1650,N_1521,N_1470);
nand U1651 (N_1651,N_1590,N_1489);
or U1652 (N_1652,N_1445,N_1572);
or U1653 (N_1653,N_1423,N_1407);
nor U1654 (N_1654,N_1419,N_1569);
or U1655 (N_1655,N_1531,N_1447);
nand U1656 (N_1656,N_1454,N_1559);
nor U1657 (N_1657,N_1416,N_1564);
nor U1658 (N_1658,N_1575,N_1493);
and U1659 (N_1659,N_1549,N_1420);
or U1660 (N_1660,N_1583,N_1542);
nand U1661 (N_1661,N_1551,N_1469);
and U1662 (N_1662,N_1409,N_1536);
or U1663 (N_1663,N_1598,N_1424);
or U1664 (N_1664,N_1482,N_1450);
or U1665 (N_1665,N_1574,N_1415);
xnor U1666 (N_1666,N_1537,N_1518);
and U1667 (N_1667,N_1408,N_1473);
nor U1668 (N_1668,N_1431,N_1490);
nor U1669 (N_1669,N_1435,N_1485);
or U1670 (N_1670,N_1541,N_1496);
or U1671 (N_1671,N_1453,N_1412);
nand U1672 (N_1672,N_1400,N_1421);
nand U1673 (N_1673,N_1488,N_1547);
nand U1674 (N_1674,N_1457,N_1449);
nand U1675 (N_1675,N_1595,N_1593);
and U1676 (N_1676,N_1511,N_1426);
or U1677 (N_1677,N_1520,N_1433);
or U1678 (N_1678,N_1517,N_1405);
and U1679 (N_1679,N_1497,N_1404);
nor U1680 (N_1680,N_1466,N_1585);
nor U1681 (N_1681,N_1491,N_1557);
and U1682 (N_1682,N_1526,N_1516);
and U1683 (N_1683,N_1566,N_1514);
and U1684 (N_1684,N_1486,N_1472);
or U1685 (N_1685,N_1462,N_1532);
or U1686 (N_1686,N_1446,N_1425);
nand U1687 (N_1687,N_1548,N_1481);
nand U1688 (N_1688,N_1597,N_1562);
and U1689 (N_1689,N_1515,N_1571);
or U1690 (N_1690,N_1580,N_1552);
and U1691 (N_1691,N_1465,N_1506);
and U1692 (N_1692,N_1434,N_1545);
or U1693 (N_1693,N_1596,N_1513);
or U1694 (N_1694,N_1567,N_1417);
nand U1695 (N_1695,N_1534,N_1487);
nor U1696 (N_1696,N_1530,N_1573);
or U1697 (N_1697,N_1509,N_1576);
or U1698 (N_1698,N_1422,N_1507);
nand U1699 (N_1699,N_1414,N_1522);
nand U1700 (N_1700,N_1533,N_1496);
or U1701 (N_1701,N_1549,N_1589);
nand U1702 (N_1702,N_1550,N_1599);
and U1703 (N_1703,N_1516,N_1428);
or U1704 (N_1704,N_1585,N_1411);
nand U1705 (N_1705,N_1523,N_1495);
nor U1706 (N_1706,N_1468,N_1490);
nand U1707 (N_1707,N_1511,N_1410);
or U1708 (N_1708,N_1521,N_1595);
xor U1709 (N_1709,N_1460,N_1403);
nor U1710 (N_1710,N_1498,N_1567);
nor U1711 (N_1711,N_1477,N_1469);
nor U1712 (N_1712,N_1566,N_1598);
and U1713 (N_1713,N_1550,N_1509);
nand U1714 (N_1714,N_1544,N_1405);
nor U1715 (N_1715,N_1506,N_1417);
nor U1716 (N_1716,N_1581,N_1476);
or U1717 (N_1717,N_1446,N_1535);
and U1718 (N_1718,N_1557,N_1514);
nand U1719 (N_1719,N_1558,N_1472);
nand U1720 (N_1720,N_1439,N_1553);
nor U1721 (N_1721,N_1430,N_1442);
nand U1722 (N_1722,N_1540,N_1456);
nor U1723 (N_1723,N_1508,N_1463);
nor U1724 (N_1724,N_1557,N_1533);
nor U1725 (N_1725,N_1545,N_1515);
nand U1726 (N_1726,N_1552,N_1517);
nor U1727 (N_1727,N_1466,N_1481);
or U1728 (N_1728,N_1570,N_1460);
or U1729 (N_1729,N_1486,N_1564);
nor U1730 (N_1730,N_1534,N_1510);
and U1731 (N_1731,N_1467,N_1461);
nand U1732 (N_1732,N_1586,N_1508);
or U1733 (N_1733,N_1491,N_1514);
nor U1734 (N_1734,N_1423,N_1442);
xnor U1735 (N_1735,N_1451,N_1435);
and U1736 (N_1736,N_1562,N_1435);
nor U1737 (N_1737,N_1578,N_1562);
nor U1738 (N_1738,N_1482,N_1484);
or U1739 (N_1739,N_1565,N_1532);
nand U1740 (N_1740,N_1515,N_1510);
and U1741 (N_1741,N_1462,N_1505);
or U1742 (N_1742,N_1494,N_1469);
and U1743 (N_1743,N_1500,N_1526);
and U1744 (N_1744,N_1469,N_1552);
nand U1745 (N_1745,N_1574,N_1559);
or U1746 (N_1746,N_1548,N_1562);
nor U1747 (N_1747,N_1562,N_1424);
nor U1748 (N_1748,N_1585,N_1417);
or U1749 (N_1749,N_1429,N_1512);
nor U1750 (N_1750,N_1436,N_1542);
or U1751 (N_1751,N_1438,N_1428);
and U1752 (N_1752,N_1475,N_1423);
and U1753 (N_1753,N_1517,N_1473);
or U1754 (N_1754,N_1545,N_1497);
or U1755 (N_1755,N_1485,N_1505);
and U1756 (N_1756,N_1488,N_1492);
nor U1757 (N_1757,N_1434,N_1438);
xor U1758 (N_1758,N_1517,N_1564);
nand U1759 (N_1759,N_1540,N_1548);
nor U1760 (N_1760,N_1509,N_1496);
or U1761 (N_1761,N_1545,N_1574);
nor U1762 (N_1762,N_1581,N_1555);
or U1763 (N_1763,N_1509,N_1412);
nor U1764 (N_1764,N_1472,N_1550);
nand U1765 (N_1765,N_1514,N_1532);
or U1766 (N_1766,N_1474,N_1400);
or U1767 (N_1767,N_1539,N_1599);
nor U1768 (N_1768,N_1433,N_1540);
and U1769 (N_1769,N_1411,N_1508);
nand U1770 (N_1770,N_1510,N_1475);
nand U1771 (N_1771,N_1561,N_1569);
nor U1772 (N_1772,N_1401,N_1407);
nand U1773 (N_1773,N_1439,N_1432);
or U1774 (N_1774,N_1495,N_1423);
nand U1775 (N_1775,N_1528,N_1512);
nor U1776 (N_1776,N_1540,N_1459);
nand U1777 (N_1777,N_1446,N_1471);
or U1778 (N_1778,N_1478,N_1408);
and U1779 (N_1779,N_1507,N_1593);
and U1780 (N_1780,N_1516,N_1512);
nor U1781 (N_1781,N_1447,N_1479);
and U1782 (N_1782,N_1453,N_1574);
nor U1783 (N_1783,N_1456,N_1517);
nor U1784 (N_1784,N_1500,N_1519);
and U1785 (N_1785,N_1468,N_1561);
nor U1786 (N_1786,N_1539,N_1417);
and U1787 (N_1787,N_1437,N_1464);
and U1788 (N_1788,N_1472,N_1434);
nor U1789 (N_1789,N_1421,N_1437);
nand U1790 (N_1790,N_1409,N_1589);
nand U1791 (N_1791,N_1468,N_1474);
and U1792 (N_1792,N_1405,N_1469);
and U1793 (N_1793,N_1443,N_1546);
and U1794 (N_1794,N_1590,N_1434);
nand U1795 (N_1795,N_1527,N_1425);
nand U1796 (N_1796,N_1472,N_1516);
or U1797 (N_1797,N_1552,N_1546);
nor U1798 (N_1798,N_1462,N_1507);
and U1799 (N_1799,N_1434,N_1513);
xor U1800 (N_1800,N_1769,N_1714);
nor U1801 (N_1801,N_1705,N_1768);
nand U1802 (N_1802,N_1749,N_1686);
and U1803 (N_1803,N_1736,N_1763);
or U1804 (N_1804,N_1703,N_1678);
nand U1805 (N_1805,N_1708,N_1781);
and U1806 (N_1806,N_1764,N_1724);
or U1807 (N_1807,N_1786,N_1795);
nand U1808 (N_1808,N_1718,N_1777);
nand U1809 (N_1809,N_1791,N_1788);
or U1810 (N_1810,N_1771,N_1612);
or U1811 (N_1811,N_1731,N_1711);
and U1812 (N_1812,N_1739,N_1726);
nand U1813 (N_1813,N_1691,N_1631);
nor U1814 (N_1814,N_1706,N_1615);
nand U1815 (N_1815,N_1798,N_1765);
or U1816 (N_1816,N_1735,N_1600);
and U1817 (N_1817,N_1619,N_1784);
nor U1818 (N_1818,N_1681,N_1758);
nand U1819 (N_1819,N_1650,N_1617);
nand U1820 (N_1820,N_1740,N_1693);
or U1821 (N_1821,N_1719,N_1672);
nand U1822 (N_1822,N_1609,N_1661);
or U1823 (N_1823,N_1762,N_1653);
and U1824 (N_1824,N_1674,N_1683);
nor U1825 (N_1825,N_1737,N_1639);
nand U1826 (N_1826,N_1642,N_1715);
nor U1827 (N_1827,N_1746,N_1742);
nor U1828 (N_1828,N_1638,N_1685);
nor U1829 (N_1829,N_1659,N_1687);
nor U1830 (N_1830,N_1689,N_1603);
or U1831 (N_1831,N_1780,N_1644);
nand U1832 (N_1832,N_1745,N_1695);
nand U1833 (N_1833,N_1774,N_1665);
nor U1834 (N_1834,N_1618,N_1649);
xnor U1835 (N_1835,N_1709,N_1744);
or U1836 (N_1836,N_1645,N_1799);
nand U1837 (N_1837,N_1680,N_1608);
nand U1838 (N_1838,N_1782,N_1716);
nand U1839 (N_1839,N_1792,N_1675);
nor U1840 (N_1840,N_1663,N_1722);
nor U1841 (N_1841,N_1669,N_1775);
nand U1842 (N_1842,N_1628,N_1641);
nand U1843 (N_1843,N_1699,N_1629);
or U1844 (N_1844,N_1658,N_1622);
nor U1845 (N_1845,N_1757,N_1747);
nor U1846 (N_1846,N_1729,N_1767);
nand U1847 (N_1847,N_1738,N_1700);
nand U1848 (N_1848,N_1643,N_1698);
nand U1849 (N_1849,N_1741,N_1694);
nor U1850 (N_1850,N_1621,N_1696);
and U1851 (N_1851,N_1704,N_1730);
nand U1852 (N_1852,N_1654,N_1766);
xnor U1853 (N_1853,N_1790,N_1620);
nand U1854 (N_1854,N_1721,N_1601);
or U1855 (N_1855,N_1688,N_1614);
nor U1856 (N_1856,N_1734,N_1793);
and U1857 (N_1857,N_1727,N_1712);
and U1858 (N_1858,N_1717,N_1677);
nor U1859 (N_1859,N_1713,N_1673);
and U1860 (N_1860,N_1660,N_1637);
or U1861 (N_1861,N_1760,N_1627);
or U1862 (N_1862,N_1682,N_1640);
nand U1863 (N_1863,N_1783,N_1647);
or U1864 (N_1864,N_1668,N_1676);
nor U1865 (N_1865,N_1606,N_1657);
or U1866 (N_1866,N_1759,N_1728);
nor U1867 (N_1867,N_1701,N_1623);
nor U1868 (N_1868,N_1761,N_1797);
nand U1869 (N_1869,N_1607,N_1754);
nor U1870 (N_1870,N_1725,N_1692);
nor U1871 (N_1871,N_1616,N_1646);
and U1872 (N_1872,N_1733,N_1662);
or U1873 (N_1873,N_1656,N_1755);
nor U1874 (N_1874,N_1748,N_1671);
and U1875 (N_1875,N_1732,N_1789);
or U1876 (N_1876,N_1778,N_1787);
and U1877 (N_1877,N_1720,N_1604);
nor U1878 (N_1878,N_1632,N_1707);
nand U1879 (N_1879,N_1690,N_1785);
nand U1880 (N_1880,N_1756,N_1684);
nand U1881 (N_1881,N_1651,N_1794);
or U1882 (N_1882,N_1613,N_1776);
nand U1883 (N_1883,N_1723,N_1648);
nand U1884 (N_1884,N_1670,N_1602);
nand U1885 (N_1885,N_1633,N_1655);
and U1886 (N_1886,N_1753,N_1605);
and U1887 (N_1887,N_1664,N_1702);
nor U1888 (N_1888,N_1679,N_1630);
nor U1889 (N_1889,N_1611,N_1624);
nor U1890 (N_1890,N_1751,N_1750);
nand U1891 (N_1891,N_1652,N_1635);
and U1892 (N_1892,N_1636,N_1743);
nor U1893 (N_1893,N_1610,N_1710);
nand U1894 (N_1894,N_1773,N_1634);
xor U1895 (N_1895,N_1667,N_1772);
and U1896 (N_1896,N_1626,N_1666);
and U1897 (N_1897,N_1625,N_1779);
and U1898 (N_1898,N_1796,N_1770);
nor U1899 (N_1899,N_1752,N_1697);
nand U1900 (N_1900,N_1669,N_1768);
nor U1901 (N_1901,N_1750,N_1766);
and U1902 (N_1902,N_1603,N_1768);
or U1903 (N_1903,N_1603,N_1691);
or U1904 (N_1904,N_1733,N_1706);
nor U1905 (N_1905,N_1774,N_1731);
nand U1906 (N_1906,N_1666,N_1667);
and U1907 (N_1907,N_1709,N_1702);
or U1908 (N_1908,N_1648,N_1655);
nor U1909 (N_1909,N_1757,N_1611);
nand U1910 (N_1910,N_1724,N_1653);
nand U1911 (N_1911,N_1784,N_1637);
nor U1912 (N_1912,N_1606,N_1626);
and U1913 (N_1913,N_1709,N_1730);
or U1914 (N_1914,N_1760,N_1664);
and U1915 (N_1915,N_1621,N_1743);
or U1916 (N_1916,N_1660,N_1601);
nand U1917 (N_1917,N_1634,N_1682);
or U1918 (N_1918,N_1748,N_1613);
or U1919 (N_1919,N_1791,N_1639);
or U1920 (N_1920,N_1746,N_1684);
or U1921 (N_1921,N_1700,N_1733);
and U1922 (N_1922,N_1744,N_1662);
nor U1923 (N_1923,N_1726,N_1725);
or U1924 (N_1924,N_1746,N_1744);
and U1925 (N_1925,N_1686,N_1600);
nor U1926 (N_1926,N_1717,N_1751);
nor U1927 (N_1927,N_1622,N_1718);
nor U1928 (N_1928,N_1743,N_1706);
and U1929 (N_1929,N_1766,N_1623);
nand U1930 (N_1930,N_1775,N_1634);
or U1931 (N_1931,N_1682,N_1623);
or U1932 (N_1932,N_1667,N_1790);
nand U1933 (N_1933,N_1742,N_1786);
nand U1934 (N_1934,N_1783,N_1657);
nor U1935 (N_1935,N_1667,N_1600);
nor U1936 (N_1936,N_1604,N_1697);
and U1937 (N_1937,N_1676,N_1642);
or U1938 (N_1938,N_1683,N_1654);
nor U1939 (N_1939,N_1638,N_1634);
xnor U1940 (N_1940,N_1618,N_1784);
nor U1941 (N_1941,N_1739,N_1612);
nor U1942 (N_1942,N_1668,N_1612);
nor U1943 (N_1943,N_1728,N_1736);
nor U1944 (N_1944,N_1745,N_1746);
or U1945 (N_1945,N_1694,N_1691);
or U1946 (N_1946,N_1753,N_1736);
or U1947 (N_1947,N_1761,N_1697);
nand U1948 (N_1948,N_1706,N_1670);
and U1949 (N_1949,N_1628,N_1656);
nor U1950 (N_1950,N_1655,N_1611);
xnor U1951 (N_1951,N_1741,N_1664);
nand U1952 (N_1952,N_1781,N_1771);
nand U1953 (N_1953,N_1643,N_1624);
nand U1954 (N_1954,N_1712,N_1753);
xnor U1955 (N_1955,N_1650,N_1712);
nor U1956 (N_1956,N_1651,N_1731);
nand U1957 (N_1957,N_1722,N_1653);
and U1958 (N_1958,N_1661,N_1614);
and U1959 (N_1959,N_1785,N_1744);
or U1960 (N_1960,N_1650,N_1610);
nor U1961 (N_1961,N_1734,N_1757);
or U1962 (N_1962,N_1618,N_1635);
nand U1963 (N_1963,N_1683,N_1691);
or U1964 (N_1964,N_1697,N_1731);
and U1965 (N_1965,N_1686,N_1695);
and U1966 (N_1966,N_1790,N_1650);
or U1967 (N_1967,N_1671,N_1750);
and U1968 (N_1968,N_1772,N_1745);
or U1969 (N_1969,N_1664,N_1609);
nor U1970 (N_1970,N_1661,N_1786);
or U1971 (N_1971,N_1779,N_1703);
or U1972 (N_1972,N_1796,N_1634);
and U1973 (N_1973,N_1600,N_1700);
or U1974 (N_1974,N_1661,N_1748);
and U1975 (N_1975,N_1699,N_1618);
or U1976 (N_1976,N_1722,N_1750);
or U1977 (N_1977,N_1753,N_1622);
and U1978 (N_1978,N_1765,N_1687);
nand U1979 (N_1979,N_1730,N_1620);
nor U1980 (N_1980,N_1652,N_1657);
xnor U1981 (N_1981,N_1619,N_1608);
and U1982 (N_1982,N_1696,N_1702);
and U1983 (N_1983,N_1682,N_1658);
or U1984 (N_1984,N_1629,N_1744);
and U1985 (N_1985,N_1603,N_1631);
xnor U1986 (N_1986,N_1775,N_1744);
xor U1987 (N_1987,N_1732,N_1614);
nor U1988 (N_1988,N_1610,N_1718);
or U1989 (N_1989,N_1765,N_1776);
and U1990 (N_1990,N_1617,N_1701);
or U1991 (N_1991,N_1698,N_1610);
or U1992 (N_1992,N_1707,N_1636);
nand U1993 (N_1993,N_1755,N_1744);
and U1994 (N_1994,N_1790,N_1797);
or U1995 (N_1995,N_1770,N_1624);
nand U1996 (N_1996,N_1705,N_1674);
nor U1997 (N_1997,N_1794,N_1655);
nor U1998 (N_1998,N_1676,N_1775);
nor U1999 (N_1999,N_1601,N_1754);
and U2000 (N_2000,N_1908,N_1885);
nor U2001 (N_2001,N_1985,N_1835);
nor U2002 (N_2002,N_1860,N_1935);
or U2003 (N_2003,N_1897,N_1868);
nand U2004 (N_2004,N_1877,N_1929);
nor U2005 (N_2005,N_1883,N_1841);
and U2006 (N_2006,N_1804,N_1831);
nor U2007 (N_2007,N_1816,N_1991);
and U2008 (N_2008,N_1887,N_1822);
nor U2009 (N_2009,N_1959,N_1881);
nor U2010 (N_2010,N_1968,N_1924);
nand U2011 (N_2011,N_1847,N_1920);
xor U2012 (N_2012,N_1916,N_1905);
nor U2013 (N_2013,N_1919,N_1862);
and U2014 (N_2014,N_1928,N_1801);
and U2015 (N_2015,N_1806,N_1923);
and U2016 (N_2016,N_1839,N_1848);
or U2017 (N_2017,N_1938,N_1954);
or U2018 (N_2018,N_1828,N_1833);
xor U2019 (N_2019,N_1844,N_1875);
and U2020 (N_2020,N_1953,N_1840);
or U2021 (N_2021,N_1931,N_1970);
and U2022 (N_2022,N_1886,N_1879);
nand U2023 (N_2023,N_1937,N_1936);
and U2024 (N_2024,N_1819,N_1882);
nor U2025 (N_2025,N_1942,N_1854);
nand U2026 (N_2026,N_1825,N_1855);
and U2027 (N_2027,N_1974,N_1966);
or U2028 (N_2028,N_1986,N_1981);
nor U2029 (N_2029,N_1832,N_1914);
or U2030 (N_2030,N_1809,N_1960);
nor U2031 (N_2031,N_1805,N_1863);
nor U2032 (N_2032,N_1814,N_1909);
nand U2033 (N_2033,N_1904,N_1918);
or U2034 (N_2034,N_1964,N_1846);
nor U2035 (N_2035,N_1823,N_1997);
and U2036 (N_2036,N_1927,N_1910);
or U2037 (N_2037,N_1926,N_1913);
nor U2038 (N_2038,N_1827,N_1945);
or U2039 (N_2039,N_1977,N_1951);
nor U2040 (N_2040,N_1849,N_1955);
nand U2041 (N_2041,N_1911,N_1851);
and U2042 (N_2042,N_1917,N_1890);
and U2043 (N_2043,N_1808,N_1907);
xnor U2044 (N_2044,N_1817,N_1915);
nor U2045 (N_2045,N_1989,N_1821);
and U2046 (N_2046,N_1940,N_1880);
and U2047 (N_2047,N_1973,N_1999);
nand U2048 (N_2048,N_1826,N_1894);
nand U2049 (N_2049,N_1956,N_1812);
nand U2050 (N_2050,N_1998,N_1990);
nor U2051 (N_2051,N_1933,N_1962);
xor U2052 (N_2052,N_1869,N_1952);
nor U2053 (N_2053,N_1946,N_1872);
or U2054 (N_2054,N_1906,N_1899);
nand U2055 (N_2055,N_1864,N_1934);
nor U2056 (N_2056,N_1963,N_1810);
nor U2057 (N_2057,N_1961,N_1878);
or U2058 (N_2058,N_1856,N_1902);
and U2059 (N_2059,N_1836,N_1976);
or U2060 (N_2060,N_1884,N_1893);
or U2061 (N_2061,N_1993,N_1967);
nand U2062 (N_2062,N_1866,N_1818);
xor U2063 (N_2063,N_1957,N_1925);
or U2064 (N_2064,N_1852,N_1859);
nand U2065 (N_2065,N_1895,N_1921);
xnor U2066 (N_2066,N_1858,N_1912);
nor U2067 (N_2067,N_1861,N_1969);
nor U2068 (N_2068,N_1820,N_1871);
or U2069 (N_2069,N_1950,N_1994);
nand U2070 (N_2070,N_1975,N_1829);
and U2071 (N_2071,N_1978,N_1896);
and U2072 (N_2072,N_1947,N_1892);
or U2073 (N_2073,N_1803,N_1811);
nor U2074 (N_2074,N_1802,N_1965);
and U2075 (N_2075,N_1807,N_1932);
nand U2076 (N_2076,N_1980,N_1992);
or U2077 (N_2077,N_1988,N_1984);
xor U2078 (N_2078,N_1888,N_1867);
or U2079 (N_2079,N_1948,N_1837);
and U2080 (N_2080,N_1996,N_1853);
nand U2081 (N_2081,N_1901,N_1944);
and U2082 (N_2082,N_1949,N_1900);
nor U2083 (N_2083,N_1995,N_1845);
or U2084 (N_2084,N_1939,N_1815);
nand U2085 (N_2085,N_1983,N_1873);
or U2086 (N_2086,N_1838,N_1874);
nand U2087 (N_2087,N_1987,N_1850);
nand U2088 (N_2088,N_1982,N_1834);
or U2089 (N_2089,N_1898,N_1903);
nand U2090 (N_2090,N_1958,N_1870);
or U2091 (N_2091,N_1843,N_1800);
or U2092 (N_2092,N_1979,N_1876);
and U2093 (N_2093,N_1971,N_1830);
nand U2094 (N_2094,N_1813,N_1842);
and U2095 (N_2095,N_1943,N_1972);
nor U2096 (N_2096,N_1889,N_1824);
or U2097 (N_2097,N_1857,N_1891);
nand U2098 (N_2098,N_1941,N_1922);
nor U2099 (N_2099,N_1865,N_1930);
nand U2100 (N_2100,N_1912,N_1991);
and U2101 (N_2101,N_1998,N_1866);
and U2102 (N_2102,N_1801,N_1885);
and U2103 (N_2103,N_1834,N_1844);
or U2104 (N_2104,N_1822,N_1970);
nand U2105 (N_2105,N_1801,N_1927);
and U2106 (N_2106,N_1815,N_1965);
nor U2107 (N_2107,N_1936,N_1912);
or U2108 (N_2108,N_1945,N_1835);
nor U2109 (N_2109,N_1927,N_1898);
nor U2110 (N_2110,N_1891,N_1864);
or U2111 (N_2111,N_1978,N_1909);
or U2112 (N_2112,N_1824,N_1864);
nand U2113 (N_2113,N_1944,N_1899);
nor U2114 (N_2114,N_1841,N_1834);
nand U2115 (N_2115,N_1900,N_1956);
nor U2116 (N_2116,N_1841,N_1809);
nand U2117 (N_2117,N_1820,N_1869);
nor U2118 (N_2118,N_1920,N_1923);
or U2119 (N_2119,N_1933,N_1993);
or U2120 (N_2120,N_1923,N_1897);
nor U2121 (N_2121,N_1961,N_1824);
nor U2122 (N_2122,N_1858,N_1877);
and U2123 (N_2123,N_1879,N_1896);
or U2124 (N_2124,N_1862,N_1908);
or U2125 (N_2125,N_1872,N_1925);
and U2126 (N_2126,N_1906,N_1863);
xnor U2127 (N_2127,N_1956,N_1966);
nand U2128 (N_2128,N_1881,N_1969);
xor U2129 (N_2129,N_1858,N_1866);
nor U2130 (N_2130,N_1827,N_1856);
or U2131 (N_2131,N_1823,N_1870);
and U2132 (N_2132,N_1829,N_1934);
or U2133 (N_2133,N_1877,N_1882);
and U2134 (N_2134,N_1824,N_1999);
nor U2135 (N_2135,N_1808,N_1855);
and U2136 (N_2136,N_1960,N_1936);
nor U2137 (N_2137,N_1837,N_1936);
or U2138 (N_2138,N_1881,N_1817);
or U2139 (N_2139,N_1889,N_1875);
nor U2140 (N_2140,N_1973,N_1997);
nand U2141 (N_2141,N_1931,N_1966);
xnor U2142 (N_2142,N_1916,N_1980);
or U2143 (N_2143,N_1961,N_1956);
nand U2144 (N_2144,N_1838,N_1945);
nand U2145 (N_2145,N_1830,N_1839);
nand U2146 (N_2146,N_1817,N_1888);
or U2147 (N_2147,N_1835,N_1829);
and U2148 (N_2148,N_1961,N_1963);
xor U2149 (N_2149,N_1881,N_1821);
or U2150 (N_2150,N_1868,N_1984);
or U2151 (N_2151,N_1814,N_1869);
and U2152 (N_2152,N_1946,N_1949);
nand U2153 (N_2153,N_1812,N_1819);
xor U2154 (N_2154,N_1933,N_1845);
nor U2155 (N_2155,N_1946,N_1846);
nor U2156 (N_2156,N_1927,N_1949);
or U2157 (N_2157,N_1981,N_1815);
xnor U2158 (N_2158,N_1844,N_1917);
nor U2159 (N_2159,N_1989,N_1949);
and U2160 (N_2160,N_1973,N_1863);
or U2161 (N_2161,N_1894,N_1845);
nand U2162 (N_2162,N_1883,N_1877);
or U2163 (N_2163,N_1864,N_1990);
nor U2164 (N_2164,N_1804,N_1850);
and U2165 (N_2165,N_1999,N_1893);
nand U2166 (N_2166,N_1996,N_1891);
or U2167 (N_2167,N_1911,N_1857);
or U2168 (N_2168,N_1987,N_1991);
nor U2169 (N_2169,N_1846,N_1954);
nand U2170 (N_2170,N_1966,N_1998);
nand U2171 (N_2171,N_1970,N_1932);
nor U2172 (N_2172,N_1965,N_1893);
or U2173 (N_2173,N_1860,N_1996);
and U2174 (N_2174,N_1927,N_1941);
or U2175 (N_2175,N_1909,N_1900);
and U2176 (N_2176,N_1912,N_1930);
or U2177 (N_2177,N_1810,N_1900);
or U2178 (N_2178,N_1998,N_1979);
nor U2179 (N_2179,N_1805,N_1862);
nor U2180 (N_2180,N_1866,N_1909);
nand U2181 (N_2181,N_1953,N_1942);
nor U2182 (N_2182,N_1831,N_1866);
nor U2183 (N_2183,N_1948,N_1942);
nor U2184 (N_2184,N_1855,N_1957);
nor U2185 (N_2185,N_1876,N_1836);
nor U2186 (N_2186,N_1882,N_1876);
and U2187 (N_2187,N_1911,N_1871);
or U2188 (N_2188,N_1832,N_1996);
nor U2189 (N_2189,N_1835,N_1915);
nand U2190 (N_2190,N_1816,N_1949);
and U2191 (N_2191,N_1945,N_1930);
or U2192 (N_2192,N_1950,N_1924);
and U2193 (N_2193,N_1949,N_1837);
and U2194 (N_2194,N_1898,N_1816);
nand U2195 (N_2195,N_1892,N_1835);
or U2196 (N_2196,N_1875,N_1964);
nand U2197 (N_2197,N_1947,N_1977);
or U2198 (N_2198,N_1857,N_1876);
or U2199 (N_2199,N_1837,N_1855);
or U2200 (N_2200,N_2136,N_2122);
nand U2201 (N_2201,N_2114,N_2007);
or U2202 (N_2202,N_2177,N_2124);
and U2203 (N_2203,N_2085,N_2148);
or U2204 (N_2204,N_2029,N_2131);
and U2205 (N_2205,N_2077,N_2076);
and U2206 (N_2206,N_2127,N_2082);
nand U2207 (N_2207,N_2067,N_2183);
nand U2208 (N_2208,N_2010,N_2176);
and U2209 (N_2209,N_2078,N_2035);
nand U2210 (N_2210,N_2090,N_2143);
or U2211 (N_2211,N_2141,N_2045);
and U2212 (N_2212,N_2180,N_2062);
or U2213 (N_2213,N_2072,N_2015);
or U2214 (N_2214,N_2043,N_2137);
nand U2215 (N_2215,N_2102,N_2151);
and U2216 (N_2216,N_2094,N_2088);
or U2217 (N_2217,N_2188,N_2116);
nor U2218 (N_2218,N_2018,N_2026);
or U2219 (N_2219,N_2028,N_2179);
nand U2220 (N_2220,N_2139,N_2111);
nor U2221 (N_2221,N_2110,N_2003);
nand U2222 (N_2222,N_2173,N_2187);
nor U2223 (N_2223,N_2021,N_2162);
or U2224 (N_2224,N_2195,N_2009);
xor U2225 (N_2225,N_2032,N_2115);
nor U2226 (N_2226,N_2123,N_2100);
or U2227 (N_2227,N_2112,N_2095);
nor U2228 (N_2228,N_2099,N_2184);
or U2229 (N_2229,N_2103,N_2134);
and U2230 (N_2230,N_2121,N_2074);
or U2231 (N_2231,N_2070,N_2169);
nand U2232 (N_2232,N_2055,N_2025);
or U2233 (N_2233,N_2101,N_2089);
nand U2234 (N_2234,N_2069,N_2059);
or U2235 (N_2235,N_2036,N_2181);
xnor U2236 (N_2236,N_2050,N_2000);
nand U2237 (N_2237,N_2109,N_2024);
xnor U2238 (N_2238,N_2152,N_2163);
nor U2239 (N_2239,N_2149,N_2033);
nand U2240 (N_2240,N_2040,N_2133);
xnor U2241 (N_2241,N_2166,N_2061);
nand U2242 (N_2242,N_2150,N_2093);
and U2243 (N_2243,N_2087,N_2005);
nand U2244 (N_2244,N_2135,N_2119);
nor U2245 (N_2245,N_2189,N_2198);
or U2246 (N_2246,N_2190,N_2052);
and U2247 (N_2247,N_2017,N_2084);
or U2248 (N_2248,N_2038,N_2118);
and U2249 (N_2249,N_2171,N_2182);
or U2250 (N_2250,N_2022,N_2104);
or U2251 (N_2251,N_2091,N_2004);
xnor U2252 (N_2252,N_2154,N_2108);
nand U2253 (N_2253,N_2128,N_2063);
nor U2254 (N_2254,N_2081,N_2153);
nor U2255 (N_2255,N_2051,N_2146);
nand U2256 (N_2256,N_2107,N_2020);
and U2257 (N_2257,N_2164,N_2129);
nand U2258 (N_2258,N_2039,N_2083);
xnor U2259 (N_2259,N_2175,N_2161);
nor U2260 (N_2260,N_2193,N_2044);
nand U2261 (N_2261,N_2034,N_2086);
nor U2262 (N_2262,N_2002,N_2012);
nor U2263 (N_2263,N_2054,N_2056);
and U2264 (N_2264,N_2001,N_2068);
or U2265 (N_2265,N_2156,N_2157);
and U2266 (N_2266,N_2008,N_2160);
nand U2267 (N_2267,N_2159,N_2142);
xor U2268 (N_2268,N_2178,N_2046);
nor U2269 (N_2269,N_2075,N_2126);
nand U2270 (N_2270,N_2138,N_2064);
or U2271 (N_2271,N_2019,N_2196);
or U2272 (N_2272,N_2047,N_2106);
and U2273 (N_2273,N_2092,N_2174);
nor U2274 (N_2274,N_2132,N_2120);
or U2275 (N_2275,N_2192,N_2096);
or U2276 (N_2276,N_2042,N_2144);
or U2277 (N_2277,N_2105,N_2117);
nor U2278 (N_2278,N_2170,N_2145);
xnor U2279 (N_2279,N_2155,N_2186);
and U2280 (N_2280,N_2066,N_2071);
nand U2281 (N_2281,N_2016,N_2060);
nand U2282 (N_2282,N_2073,N_2079);
nand U2283 (N_2283,N_2053,N_2065);
nand U2284 (N_2284,N_2197,N_2027);
nand U2285 (N_2285,N_2006,N_2037);
nand U2286 (N_2286,N_2147,N_2191);
nand U2287 (N_2287,N_2113,N_2057);
nand U2288 (N_2288,N_2194,N_2023);
nand U2289 (N_2289,N_2049,N_2058);
nand U2290 (N_2290,N_2158,N_2172);
and U2291 (N_2291,N_2011,N_2031);
nand U2292 (N_2292,N_2098,N_2185);
nor U2293 (N_2293,N_2048,N_2030);
or U2294 (N_2294,N_2014,N_2080);
and U2295 (N_2295,N_2013,N_2167);
and U2296 (N_2296,N_2130,N_2165);
or U2297 (N_2297,N_2199,N_2097);
and U2298 (N_2298,N_2125,N_2140);
xor U2299 (N_2299,N_2168,N_2041);
and U2300 (N_2300,N_2010,N_2110);
or U2301 (N_2301,N_2142,N_2178);
and U2302 (N_2302,N_2133,N_2122);
and U2303 (N_2303,N_2120,N_2017);
nand U2304 (N_2304,N_2040,N_2080);
and U2305 (N_2305,N_2133,N_2018);
or U2306 (N_2306,N_2163,N_2096);
nor U2307 (N_2307,N_2114,N_2125);
nor U2308 (N_2308,N_2188,N_2158);
and U2309 (N_2309,N_2183,N_2097);
nand U2310 (N_2310,N_2194,N_2106);
nor U2311 (N_2311,N_2023,N_2022);
nand U2312 (N_2312,N_2043,N_2037);
nor U2313 (N_2313,N_2161,N_2037);
nand U2314 (N_2314,N_2106,N_2195);
nand U2315 (N_2315,N_2060,N_2022);
nand U2316 (N_2316,N_2188,N_2011);
or U2317 (N_2317,N_2179,N_2039);
or U2318 (N_2318,N_2141,N_2162);
xor U2319 (N_2319,N_2156,N_2119);
nor U2320 (N_2320,N_2167,N_2053);
or U2321 (N_2321,N_2173,N_2165);
or U2322 (N_2322,N_2057,N_2089);
or U2323 (N_2323,N_2030,N_2036);
or U2324 (N_2324,N_2199,N_2150);
nor U2325 (N_2325,N_2029,N_2056);
and U2326 (N_2326,N_2009,N_2149);
or U2327 (N_2327,N_2100,N_2047);
nor U2328 (N_2328,N_2027,N_2075);
nor U2329 (N_2329,N_2153,N_2113);
nand U2330 (N_2330,N_2038,N_2162);
and U2331 (N_2331,N_2103,N_2100);
or U2332 (N_2332,N_2123,N_2182);
or U2333 (N_2333,N_2103,N_2163);
nor U2334 (N_2334,N_2146,N_2079);
nand U2335 (N_2335,N_2078,N_2126);
nor U2336 (N_2336,N_2072,N_2120);
nand U2337 (N_2337,N_2009,N_2079);
and U2338 (N_2338,N_2154,N_2130);
nand U2339 (N_2339,N_2132,N_2022);
nor U2340 (N_2340,N_2166,N_2025);
nand U2341 (N_2341,N_2151,N_2010);
nand U2342 (N_2342,N_2078,N_2015);
nand U2343 (N_2343,N_2002,N_2138);
and U2344 (N_2344,N_2046,N_2101);
nand U2345 (N_2345,N_2084,N_2011);
nand U2346 (N_2346,N_2195,N_2180);
and U2347 (N_2347,N_2097,N_2188);
nor U2348 (N_2348,N_2078,N_2181);
nand U2349 (N_2349,N_2117,N_2145);
or U2350 (N_2350,N_2068,N_2088);
nor U2351 (N_2351,N_2055,N_2049);
and U2352 (N_2352,N_2004,N_2139);
or U2353 (N_2353,N_2065,N_2176);
or U2354 (N_2354,N_2014,N_2143);
xnor U2355 (N_2355,N_2148,N_2068);
nor U2356 (N_2356,N_2179,N_2162);
nand U2357 (N_2357,N_2033,N_2098);
nor U2358 (N_2358,N_2131,N_2026);
nor U2359 (N_2359,N_2031,N_2104);
nand U2360 (N_2360,N_2109,N_2160);
or U2361 (N_2361,N_2159,N_2102);
or U2362 (N_2362,N_2121,N_2019);
or U2363 (N_2363,N_2004,N_2178);
and U2364 (N_2364,N_2179,N_2176);
or U2365 (N_2365,N_2091,N_2120);
or U2366 (N_2366,N_2159,N_2153);
or U2367 (N_2367,N_2024,N_2051);
or U2368 (N_2368,N_2014,N_2065);
nor U2369 (N_2369,N_2045,N_2175);
nand U2370 (N_2370,N_2009,N_2139);
nand U2371 (N_2371,N_2162,N_2005);
nand U2372 (N_2372,N_2190,N_2145);
or U2373 (N_2373,N_2113,N_2074);
nor U2374 (N_2374,N_2058,N_2165);
or U2375 (N_2375,N_2115,N_2127);
nand U2376 (N_2376,N_2170,N_2009);
nand U2377 (N_2377,N_2053,N_2024);
nand U2378 (N_2378,N_2159,N_2107);
or U2379 (N_2379,N_2161,N_2060);
and U2380 (N_2380,N_2110,N_2184);
or U2381 (N_2381,N_2013,N_2082);
or U2382 (N_2382,N_2161,N_2008);
nand U2383 (N_2383,N_2053,N_2140);
nor U2384 (N_2384,N_2045,N_2104);
nor U2385 (N_2385,N_2035,N_2104);
and U2386 (N_2386,N_2186,N_2030);
and U2387 (N_2387,N_2161,N_2134);
nand U2388 (N_2388,N_2058,N_2019);
and U2389 (N_2389,N_2182,N_2073);
nor U2390 (N_2390,N_2188,N_2062);
xnor U2391 (N_2391,N_2016,N_2123);
nor U2392 (N_2392,N_2103,N_2044);
and U2393 (N_2393,N_2019,N_2079);
nand U2394 (N_2394,N_2026,N_2140);
or U2395 (N_2395,N_2056,N_2116);
nor U2396 (N_2396,N_2044,N_2146);
nand U2397 (N_2397,N_2024,N_2157);
and U2398 (N_2398,N_2134,N_2085);
or U2399 (N_2399,N_2184,N_2008);
nor U2400 (N_2400,N_2361,N_2294);
or U2401 (N_2401,N_2399,N_2218);
nand U2402 (N_2402,N_2339,N_2392);
and U2403 (N_2403,N_2315,N_2211);
nor U2404 (N_2404,N_2202,N_2396);
nor U2405 (N_2405,N_2223,N_2235);
nand U2406 (N_2406,N_2351,N_2205);
nor U2407 (N_2407,N_2216,N_2219);
nor U2408 (N_2408,N_2367,N_2230);
nand U2409 (N_2409,N_2299,N_2380);
nand U2410 (N_2410,N_2206,N_2311);
nor U2411 (N_2411,N_2328,N_2213);
or U2412 (N_2412,N_2336,N_2329);
nor U2413 (N_2413,N_2395,N_2314);
and U2414 (N_2414,N_2278,N_2261);
and U2415 (N_2415,N_2243,N_2266);
or U2416 (N_2416,N_2276,N_2309);
nor U2417 (N_2417,N_2267,N_2300);
or U2418 (N_2418,N_2391,N_2238);
nand U2419 (N_2419,N_2225,N_2305);
nor U2420 (N_2420,N_2227,N_2322);
and U2421 (N_2421,N_2386,N_2360);
or U2422 (N_2422,N_2249,N_2247);
and U2423 (N_2423,N_2272,N_2203);
and U2424 (N_2424,N_2286,N_2368);
nor U2425 (N_2425,N_2217,N_2275);
or U2426 (N_2426,N_2332,N_2274);
and U2427 (N_2427,N_2372,N_2341);
nor U2428 (N_2428,N_2295,N_2264);
xnor U2429 (N_2429,N_2240,N_2383);
or U2430 (N_2430,N_2317,N_2224);
or U2431 (N_2431,N_2262,N_2338);
xor U2432 (N_2432,N_2226,N_2304);
and U2433 (N_2433,N_2285,N_2237);
and U2434 (N_2434,N_2355,N_2302);
nand U2435 (N_2435,N_2365,N_2371);
or U2436 (N_2436,N_2231,N_2385);
nand U2437 (N_2437,N_2320,N_2318);
or U2438 (N_2438,N_2335,N_2331);
or U2439 (N_2439,N_2236,N_2250);
and U2440 (N_2440,N_2324,N_2333);
or U2441 (N_2441,N_2384,N_2390);
nand U2442 (N_2442,N_2345,N_2233);
nor U2443 (N_2443,N_2290,N_2270);
or U2444 (N_2444,N_2228,N_2291);
or U2445 (N_2445,N_2271,N_2248);
nand U2446 (N_2446,N_2357,N_2352);
and U2447 (N_2447,N_2340,N_2347);
or U2448 (N_2448,N_2200,N_2337);
nor U2449 (N_2449,N_2389,N_2349);
nand U2450 (N_2450,N_2292,N_2222);
nor U2451 (N_2451,N_2239,N_2207);
and U2452 (N_2452,N_2310,N_2381);
and U2453 (N_2453,N_2374,N_2287);
nor U2454 (N_2454,N_2398,N_2387);
xor U2455 (N_2455,N_2353,N_2356);
or U2456 (N_2456,N_2229,N_2369);
nand U2457 (N_2457,N_2246,N_2253);
or U2458 (N_2458,N_2346,N_2343);
nand U2459 (N_2459,N_2354,N_2215);
and U2460 (N_2460,N_2394,N_2279);
or U2461 (N_2461,N_2312,N_2313);
nand U2462 (N_2462,N_2366,N_2297);
nor U2463 (N_2463,N_2280,N_2208);
and U2464 (N_2464,N_2263,N_2373);
and U2465 (N_2465,N_2393,N_2260);
or U2466 (N_2466,N_2362,N_2220);
nand U2467 (N_2467,N_2283,N_2289);
nor U2468 (N_2468,N_2214,N_2342);
and U2469 (N_2469,N_2378,N_2388);
nand U2470 (N_2470,N_2375,N_2259);
nand U2471 (N_2471,N_2258,N_2308);
nor U2472 (N_2472,N_2363,N_2370);
or U2473 (N_2473,N_2284,N_2209);
nand U2474 (N_2474,N_2204,N_2334);
nand U2475 (N_2475,N_2293,N_2254);
and U2476 (N_2476,N_2282,N_2256);
nand U2477 (N_2477,N_2325,N_2301);
and U2478 (N_2478,N_2382,N_2298);
and U2479 (N_2479,N_2210,N_2281);
nand U2480 (N_2480,N_2201,N_2234);
nor U2481 (N_2481,N_2358,N_2221);
nor U2482 (N_2482,N_2316,N_2364);
nor U2483 (N_2483,N_2327,N_2348);
or U2484 (N_2484,N_2376,N_2251);
or U2485 (N_2485,N_2307,N_2244);
nand U2486 (N_2486,N_2321,N_2212);
or U2487 (N_2487,N_2330,N_2326);
or U2488 (N_2488,N_2377,N_2245);
nand U2489 (N_2489,N_2252,N_2397);
or U2490 (N_2490,N_2257,N_2268);
nand U2491 (N_2491,N_2277,N_2306);
nor U2492 (N_2492,N_2319,N_2379);
nor U2493 (N_2493,N_2273,N_2265);
or U2494 (N_2494,N_2232,N_2255);
and U2495 (N_2495,N_2323,N_2303);
xor U2496 (N_2496,N_2344,N_2242);
nor U2497 (N_2497,N_2241,N_2296);
or U2498 (N_2498,N_2359,N_2288);
nand U2499 (N_2499,N_2350,N_2269);
nor U2500 (N_2500,N_2261,N_2237);
or U2501 (N_2501,N_2329,N_2252);
nand U2502 (N_2502,N_2360,N_2319);
or U2503 (N_2503,N_2335,N_2301);
and U2504 (N_2504,N_2242,N_2224);
nand U2505 (N_2505,N_2303,N_2207);
or U2506 (N_2506,N_2250,N_2300);
nor U2507 (N_2507,N_2255,N_2216);
nor U2508 (N_2508,N_2337,N_2227);
nor U2509 (N_2509,N_2343,N_2316);
and U2510 (N_2510,N_2220,N_2207);
nand U2511 (N_2511,N_2310,N_2208);
nor U2512 (N_2512,N_2361,N_2288);
and U2513 (N_2513,N_2393,N_2325);
and U2514 (N_2514,N_2328,N_2337);
nor U2515 (N_2515,N_2275,N_2263);
and U2516 (N_2516,N_2325,N_2239);
nor U2517 (N_2517,N_2245,N_2279);
or U2518 (N_2518,N_2321,N_2313);
or U2519 (N_2519,N_2271,N_2283);
nand U2520 (N_2520,N_2310,N_2231);
nor U2521 (N_2521,N_2294,N_2373);
nand U2522 (N_2522,N_2236,N_2364);
nor U2523 (N_2523,N_2299,N_2210);
and U2524 (N_2524,N_2341,N_2367);
nor U2525 (N_2525,N_2296,N_2382);
and U2526 (N_2526,N_2304,N_2294);
nand U2527 (N_2527,N_2253,N_2273);
or U2528 (N_2528,N_2382,N_2240);
or U2529 (N_2529,N_2254,N_2355);
or U2530 (N_2530,N_2285,N_2306);
and U2531 (N_2531,N_2287,N_2248);
and U2532 (N_2532,N_2246,N_2267);
or U2533 (N_2533,N_2200,N_2246);
and U2534 (N_2534,N_2387,N_2306);
nor U2535 (N_2535,N_2200,N_2208);
nand U2536 (N_2536,N_2279,N_2365);
and U2537 (N_2537,N_2364,N_2361);
or U2538 (N_2538,N_2314,N_2217);
nor U2539 (N_2539,N_2390,N_2362);
nor U2540 (N_2540,N_2259,N_2357);
nand U2541 (N_2541,N_2306,N_2223);
nand U2542 (N_2542,N_2361,N_2296);
nor U2543 (N_2543,N_2227,N_2399);
or U2544 (N_2544,N_2348,N_2363);
nor U2545 (N_2545,N_2351,N_2227);
nor U2546 (N_2546,N_2337,N_2313);
or U2547 (N_2547,N_2237,N_2367);
nor U2548 (N_2548,N_2370,N_2338);
and U2549 (N_2549,N_2390,N_2200);
or U2550 (N_2550,N_2360,N_2371);
or U2551 (N_2551,N_2298,N_2229);
nor U2552 (N_2552,N_2290,N_2235);
nand U2553 (N_2553,N_2350,N_2346);
nand U2554 (N_2554,N_2335,N_2278);
nand U2555 (N_2555,N_2238,N_2389);
nor U2556 (N_2556,N_2204,N_2393);
nand U2557 (N_2557,N_2255,N_2200);
and U2558 (N_2558,N_2223,N_2340);
xor U2559 (N_2559,N_2248,N_2346);
nor U2560 (N_2560,N_2321,N_2370);
nand U2561 (N_2561,N_2237,N_2210);
or U2562 (N_2562,N_2256,N_2377);
and U2563 (N_2563,N_2279,N_2324);
and U2564 (N_2564,N_2321,N_2211);
nand U2565 (N_2565,N_2291,N_2297);
or U2566 (N_2566,N_2348,N_2300);
or U2567 (N_2567,N_2316,N_2314);
or U2568 (N_2568,N_2289,N_2354);
and U2569 (N_2569,N_2322,N_2312);
and U2570 (N_2570,N_2392,N_2298);
nand U2571 (N_2571,N_2366,N_2395);
nand U2572 (N_2572,N_2207,N_2328);
and U2573 (N_2573,N_2204,N_2200);
nor U2574 (N_2574,N_2243,N_2350);
nand U2575 (N_2575,N_2296,N_2385);
nor U2576 (N_2576,N_2351,N_2320);
nor U2577 (N_2577,N_2213,N_2224);
and U2578 (N_2578,N_2273,N_2319);
nand U2579 (N_2579,N_2285,N_2371);
or U2580 (N_2580,N_2251,N_2266);
nand U2581 (N_2581,N_2321,N_2233);
and U2582 (N_2582,N_2284,N_2227);
nor U2583 (N_2583,N_2293,N_2222);
nor U2584 (N_2584,N_2383,N_2210);
or U2585 (N_2585,N_2391,N_2388);
nand U2586 (N_2586,N_2384,N_2304);
or U2587 (N_2587,N_2351,N_2387);
nor U2588 (N_2588,N_2295,N_2293);
nand U2589 (N_2589,N_2373,N_2332);
nor U2590 (N_2590,N_2230,N_2348);
and U2591 (N_2591,N_2311,N_2369);
nor U2592 (N_2592,N_2226,N_2376);
or U2593 (N_2593,N_2296,N_2391);
nor U2594 (N_2594,N_2324,N_2222);
nor U2595 (N_2595,N_2228,N_2231);
and U2596 (N_2596,N_2206,N_2308);
or U2597 (N_2597,N_2388,N_2384);
nand U2598 (N_2598,N_2224,N_2311);
nand U2599 (N_2599,N_2214,N_2210);
and U2600 (N_2600,N_2512,N_2508);
or U2601 (N_2601,N_2555,N_2583);
and U2602 (N_2602,N_2463,N_2485);
and U2603 (N_2603,N_2588,N_2577);
or U2604 (N_2604,N_2525,N_2514);
nand U2605 (N_2605,N_2529,N_2576);
or U2606 (N_2606,N_2516,N_2416);
and U2607 (N_2607,N_2584,N_2560);
nand U2608 (N_2608,N_2455,N_2476);
or U2609 (N_2609,N_2412,N_2450);
nor U2610 (N_2610,N_2597,N_2535);
or U2611 (N_2611,N_2470,N_2498);
nand U2612 (N_2612,N_2472,N_2441);
nand U2613 (N_2613,N_2545,N_2487);
or U2614 (N_2614,N_2561,N_2547);
nand U2615 (N_2615,N_2581,N_2549);
and U2616 (N_2616,N_2411,N_2464);
nand U2617 (N_2617,N_2518,N_2417);
nand U2618 (N_2618,N_2539,N_2474);
nand U2619 (N_2619,N_2400,N_2510);
nand U2620 (N_2620,N_2590,N_2460);
and U2621 (N_2621,N_2552,N_2537);
nand U2622 (N_2622,N_2505,N_2488);
nand U2623 (N_2623,N_2509,N_2420);
nor U2624 (N_2624,N_2407,N_2458);
and U2625 (N_2625,N_2502,N_2503);
xor U2626 (N_2626,N_2595,N_2515);
nand U2627 (N_2627,N_2406,N_2469);
and U2628 (N_2628,N_2478,N_2570);
nand U2629 (N_2629,N_2456,N_2447);
nor U2630 (N_2630,N_2489,N_2538);
and U2631 (N_2631,N_2586,N_2497);
nor U2632 (N_2632,N_2452,N_2499);
nor U2633 (N_2633,N_2580,N_2421);
nor U2634 (N_2634,N_2507,N_2449);
or U2635 (N_2635,N_2462,N_2433);
nor U2636 (N_2636,N_2536,N_2480);
and U2637 (N_2637,N_2427,N_2454);
nand U2638 (N_2638,N_2435,N_2568);
xor U2639 (N_2639,N_2453,N_2541);
and U2640 (N_2640,N_2591,N_2496);
or U2641 (N_2641,N_2443,N_2429);
nand U2642 (N_2642,N_2511,N_2596);
nand U2643 (N_2643,N_2431,N_2520);
or U2644 (N_2644,N_2504,N_2532);
nor U2645 (N_2645,N_2594,N_2461);
or U2646 (N_2646,N_2418,N_2425);
and U2647 (N_2647,N_2519,N_2424);
or U2648 (N_2648,N_2436,N_2543);
nand U2649 (N_2649,N_2553,N_2523);
or U2650 (N_2650,N_2402,N_2530);
or U2651 (N_2651,N_2559,N_2565);
nand U2652 (N_2652,N_2527,N_2528);
nor U2653 (N_2653,N_2569,N_2526);
nor U2654 (N_2654,N_2459,N_2524);
nor U2655 (N_2655,N_2494,N_2414);
and U2656 (N_2656,N_2546,N_2408);
nand U2657 (N_2657,N_2554,N_2432);
and U2658 (N_2658,N_2467,N_2423);
nor U2659 (N_2659,N_2403,N_2599);
and U2660 (N_2660,N_2548,N_2567);
nand U2661 (N_2661,N_2562,N_2540);
and U2662 (N_2662,N_2491,N_2517);
nor U2663 (N_2663,N_2405,N_2468);
nor U2664 (N_2664,N_2434,N_2493);
and U2665 (N_2665,N_2558,N_2426);
or U2666 (N_2666,N_2448,N_2531);
or U2667 (N_2667,N_2593,N_2575);
and U2668 (N_2668,N_2582,N_2563);
or U2669 (N_2669,N_2483,N_2544);
and U2670 (N_2670,N_2589,N_2404);
and U2671 (N_2671,N_2430,N_2444);
or U2672 (N_2672,N_2446,N_2445);
nand U2673 (N_2673,N_2439,N_2579);
nor U2674 (N_2674,N_2564,N_2466);
or U2675 (N_2675,N_2592,N_2501);
or U2676 (N_2676,N_2513,N_2542);
and U2677 (N_2677,N_2486,N_2521);
or U2678 (N_2678,N_2587,N_2410);
or U2679 (N_2679,N_2522,N_2438);
nor U2680 (N_2680,N_2475,N_2556);
nand U2681 (N_2681,N_2419,N_2415);
nand U2682 (N_2682,N_2571,N_2534);
or U2683 (N_2683,N_2551,N_2465);
and U2684 (N_2684,N_2574,N_2506);
or U2685 (N_2685,N_2492,N_2413);
or U2686 (N_2686,N_2495,N_2500);
nor U2687 (N_2687,N_2440,N_2481);
nor U2688 (N_2688,N_2557,N_2457);
and U2689 (N_2689,N_2484,N_2598);
or U2690 (N_2690,N_2451,N_2490);
nor U2691 (N_2691,N_2479,N_2477);
and U2692 (N_2692,N_2578,N_2428);
nor U2693 (N_2693,N_2482,N_2401);
and U2694 (N_2694,N_2422,N_2473);
nor U2695 (N_2695,N_2471,N_2550);
nor U2696 (N_2696,N_2437,N_2572);
and U2697 (N_2697,N_2442,N_2585);
nand U2698 (N_2698,N_2533,N_2573);
and U2699 (N_2699,N_2409,N_2566);
xor U2700 (N_2700,N_2578,N_2478);
xor U2701 (N_2701,N_2571,N_2417);
and U2702 (N_2702,N_2455,N_2529);
or U2703 (N_2703,N_2549,N_2535);
nor U2704 (N_2704,N_2484,N_2510);
nor U2705 (N_2705,N_2577,N_2570);
and U2706 (N_2706,N_2507,N_2536);
nor U2707 (N_2707,N_2538,N_2404);
xor U2708 (N_2708,N_2544,N_2563);
nor U2709 (N_2709,N_2428,N_2527);
nor U2710 (N_2710,N_2548,N_2429);
and U2711 (N_2711,N_2585,N_2471);
nor U2712 (N_2712,N_2447,N_2406);
nor U2713 (N_2713,N_2582,N_2543);
nor U2714 (N_2714,N_2423,N_2492);
nand U2715 (N_2715,N_2557,N_2406);
nand U2716 (N_2716,N_2516,N_2492);
nor U2717 (N_2717,N_2569,N_2567);
nand U2718 (N_2718,N_2478,N_2401);
nor U2719 (N_2719,N_2596,N_2422);
and U2720 (N_2720,N_2413,N_2474);
or U2721 (N_2721,N_2444,N_2405);
or U2722 (N_2722,N_2441,N_2575);
nor U2723 (N_2723,N_2440,N_2482);
nor U2724 (N_2724,N_2551,N_2579);
nor U2725 (N_2725,N_2503,N_2407);
nor U2726 (N_2726,N_2590,N_2501);
or U2727 (N_2727,N_2424,N_2501);
and U2728 (N_2728,N_2433,N_2510);
nand U2729 (N_2729,N_2476,N_2555);
or U2730 (N_2730,N_2552,N_2439);
nor U2731 (N_2731,N_2505,N_2519);
or U2732 (N_2732,N_2478,N_2511);
or U2733 (N_2733,N_2400,N_2548);
xnor U2734 (N_2734,N_2513,N_2547);
nor U2735 (N_2735,N_2419,N_2475);
nand U2736 (N_2736,N_2472,N_2560);
and U2737 (N_2737,N_2598,N_2417);
nor U2738 (N_2738,N_2526,N_2589);
nor U2739 (N_2739,N_2506,N_2572);
nor U2740 (N_2740,N_2582,N_2533);
and U2741 (N_2741,N_2440,N_2500);
and U2742 (N_2742,N_2486,N_2411);
nand U2743 (N_2743,N_2425,N_2494);
nand U2744 (N_2744,N_2452,N_2496);
nor U2745 (N_2745,N_2407,N_2463);
nor U2746 (N_2746,N_2559,N_2582);
nand U2747 (N_2747,N_2479,N_2570);
and U2748 (N_2748,N_2511,N_2421);
xor U2749 (N_2749,N_2421,N_2457);
nor U2750 (N_2750,N_2599,N_2587);
or U2751 (N_2751,N_2512,N_2472);
and U2752 (N_2752,N_2424,N_2550);
and U2753 (N_2753,N_2488,N_2582);
and U2754 (N_2754,N_2571,N_2598);
and U2755 (N_2755,N_2452,N_2461);
or U2756 (N_2756,N_2513,N_2543);
nor U2757 (N_2757,N_2458,N_2493);
nand U2758 (N_2758,N_2419,N_2567);
or U2759 (N_2759,N_2595,N_2423);
nand U2760 (N_2760,N_2435,N_2467);
or U2761 (N_2761,N_2467,N_2580);
nand U2762 (N_2762,N_2522,N_2542);
or U2763 (N_2763,N_2478,N_2543);
nor U2764 (N_2764,N_2579,N_2476);
nor U2765 (N_2765,N_2545,N_2536);
and U2766 (N_2766,N_2429,N_2578);
nor U2767 (N_2767,N_2540,N_2535);
and U2768 (N_2768,N_2490,N_2532);
nand U2769 (N_2769,N_2419,N_2527);
nand U2770 (N_2770,N_2445,N_2569);
nor U2771 (N_2771,N_2494,N_2462);
and U2772 (N_2772,N_2462,N_2454);
nand U2773 (N_2773,N_2499,N_2545);
and U2774 (N_2774,N_2500,N_2485);
nand U2775 (N_2775,N_2543,N_2406);
nor U2776 (N_2776,N_2584,N_2578);
and U2777 (N_2777,N_2566,N_2511);
or U2778 (N_2778,N_2439,N_2461);
and U2779 (N_2779,N_2541,N_2404);
or U2780 (N_2780,N_2414,N_2418);
and U2781 (N_2781,N_2449,N_2593);
or U2782 (N_2782,N_2523,N_2552);
and U2783 (N_2783,N_2482,N_2592);
and U2784 (N_2784,N_2434,N_2460);
nor U2785 (N_2785,N_2582,N_2517);
nor U2786 (N_2786,N_2404,N_2458);
nor U2787 (N_2787,N_2436,N_2459);
and U2788 (N_2788,N_2403,N_2503);
or U2789 (N_2789,N_2586,N_2517);
and U2790 (N_2790,N_2436,N_2537);
and U2791 (N_2791,N_2576,N_2469);
nand U2792 (N_2792,N_2407,N_2564);
or U2793 (N_2793,N_2514,N_2531);
and U2794 (N_2794,N_2541,N_2579);
nor U2795 (N_2795,N_2472,N_2506);
nor U2796 (N_2796,N_2440,N_2531);
nor U2797 (N_2797,N_2499,N_2408);
nor U2798 (N_2798,N_2450,N_2481);
and U2799 (N_2799,N_2425,N_2471);
nor U2800 (N_2800,N_2650,N_2631);
nor U2801 (N_2801,N_2678,N_2779);
nor U2802 (N_2802,N_2743,N_2619);
nand U2803 (N_2803,N_2679,N_2682);
or U2804 (N_2804,N_2791,N_2642);
nor U2805 (N_2805,N_2633,N_2794);
nand U2806 (N_2806,N_2721,N_2783);
and U2807 (N_2807,N_2748,N_2752);
or U2808 (N_2808,N_2742,N_2618);
or U2809 (N_2809,N_2747,N_2627);
and U2810 (N_2810,N_2683,N_2640);
and U2811 (N_2811,N_2692,N_2646);
nor U2812 (N_2812,N_2621,N_2775);
and U2813 (N_2813,N_2770,N_2781);
and U2814 (N_2814,N_2704,N_2762);
nand U2815 (N_2815,N_2637,N_2700);
nor U2816 (N_2816,N_2788,N_2703);
or U2817 (N_2817,N_2699,N_2668);
nand U2818 (N_2818,N_2665,N_2720);
nand U2819 (N_2819,N_2758,N_2790);
and U2820 (N_2820,N_2728,N_2709);
and U2821 (N_2821,N_2629,N_2702);
or U2822 (N_2822,N_2691,N_2714);
nor U2823 (N_2823,N_2707,N_2745);
nand U2824 (N_2824,N_2751,N_2687);
and U2825 (N_2825,N_2765,N_2705);
nand U2826 (N_2826,N_2656,N_2738);
or U2827 (N_2827,N_2663,N_2706);
nor U2828 (N_2828,N_2772,N_2757);
nand U2829 (N_2829,N_2648,N_2754);
nor U2830 (N_2830,N_2773,N_2649);
or U2831 (N_2831,N_2603,N_2763);
or U2832 (N_2832,N_2639,N_2712);
or U2833 (N_2833,N_2761,N_2744);
or U2834 (N_2834,N_2673,N_2734);
nor U2835 (N_2835,N_2667,N_2630);
nor U2836 (N_2836,N_2787,N_2643);
or U2837 (N_2837,N_2750,N_2601);
and U2838 (N_2838,N_2749,N_2614);
or U2839 (N_2839,N_2661,N_2680);
nand U2840 (N_2840,N_2769,N_2622);
or U2841 (N_2841,N_2670,N_2776);
and U2842 (N_2842,N_2708,N_2777);
or U2843 (N_2843,N_2654,N_2644);
nand U2844 (N_2844,N_2625,N_2792);
nor U2845 (N_2845,N_2632,N_2789);
or U2846 (N_2846,N_2722,N_2652);
nand U2847 (N_2847,N_2647,N_2624);
or U2848 (N_2848,N_2684,N_2732);
nand U2849 (N_2849,N_2780,N_2676);
nor U2850 (N_2850,N_2784,N_2753);
nand U2851 (N_2851,N_2701,N_2604);
nand U2852 (N_2852,N_2795,N_2739);
nand U2853 (N_2853,N_2685,N_2612);
and U2854 (N_2854,N_2608,N_2730);
and U2855 (N_2855,N_2797,N_2737);
nor U2856 (N_2856,N_2716,N_2609);
and U2857 (N_2857,N_2710,N_2713);
nand U2858 (N_2858,N_2616,N_2759);
and U2859 (N_2859,N_2767,N_2740);
or U2860 (N_2860,N_2696,N_2600);
xor U2861 (N_2861,N_2617,N_2666);
and U2862 (N_2862,N_2690,N_2686);
nor U2863 (N_2863,N_2755,N_2674);
nand U2864 (N_2864,N_2669,N_2694);
or U2865 (N_2865,N_2636,N_2764);
or U2866 (N_2866,N_2611,N_2785);
nand U2867 (N_2867,N_2613,N_2727);
and U2868 (N_2868,N_2606,N_2653);
and U2869 (N_2869,N_2651,N_2723);
and U2870 (N_2870,N_2726,N_2638);
nor U2871 (N_2871,N_2655,N_2681);
or U2872 (N_2872,N_2766,N_2731);
and U2873 (N_2873,N_2698,N_2733);
or U2874 (N_2874,N_2658,N_2715);
nand U2875 (N_2875,N_2689,N_2641);
nand U2876 (N_2876,N_2634,N_2695);
xor U2877 (N_2877,N_2623,N_2756);
or U2878 (N_2878,N_2693,N_2672);
nor U2879 (N_2879,N_2717,N_2736);
or U2880 (N_2880,N_2782,N_2760);
and U2881 (N_2881,N_2796,N_2798);
nand U2882 (N_2882,N_2718,N_2688);
or U2883 (N_2883,N_2697,N_2793);
nor U2884 (N_2884,N_2778,N_2677);
nor U2885 (N_2885,N_2607,N_2799);
nand U2886 (N_2886,N_2741,N_2729);
or U2887 (N_2887,N_2605,N_2771);
nor U2888 (N_2888,N_2774,N_2635);
nor U2889 (N_2889,N_2711,N_2746);
nor U2890 (N_2890,N_2735,N_2719);
and U2891 (N_2891,N_2657,N_2664);
or U2892 (N_2892,N_2724,N_2660);
or U2893 (N_2893,N_2626,N_2662);
and U2894 (N_2894,N_2725,N_2610);
and U2895 (N_2895,N_2615,N_2620);
nor U2896 (N_2896,N_2628,N_2768);
and U2897 (N_2897,N_2602,N_2671);
and U2898 (N_2898,N_2786,N_2675);
nand U2899 (N_2899,N_2659,N_2645);
and U2900 (N_2900,N_2649,N_2719);
nand U2901 (N_2901,N_2735,N_2681);
nor U2902 (N_2902,N_2672,N_2783);
nand U2903 (N_2903,N_2759,N_2742);
or U2904 (N_2904,N_2641,N_2758);
nand U2905 (N_2905,N_2617,N_2758);
or U2906 (N_2906,N_2744,N_2680);
or U2907 (N_2907,N_2783,N_2683);
and U2908 (N_2908,N_2618,N_2782);
nor U2909 (N_2909,N_2735,N_2778);
or U2910 (N_2910,N_2627,N_2722);
or U2911 (N_2911,N_2680,N_2759);
and U2912 (N_2912,N_2621,N_2750);
and U2913 (N_2913,N_2676,N_2786);
nor U2914 (N_2914,N_2691,N_2692);
nor U2915 (N_2915,N_2674,N_2732);
nand U2916 (N_2916,N_2781,N_2723);
nor U2917 (N_2917,N_2642,N_2738);
nand U2918 (N_2918,N_2756,N_2669);
nor U2919 (N_2919,N_2611,N_2693);
and U2920 (N_2920,N_2673,N_2726);
and U2921 (N_2921,N_2652,N_2614);
or U2922 (N_2922,N_2641,N_2667);
or U2923 (N_2923,N_2790,N_2792);
nor U2924 (N_2924,N_2639,N_2606);
or U2925 (N_2925,N_2630,N_2631);
nand U2926 (N_2926,N_2692,N_2700);
and U2927 (N_2927,N_2764,N_2791);
and U2928 (N_2928,N_2718,N_2771);
nor U2929 (N_2929,N_2707,N_2753);
or U2930 (N_2930,N_2607,N_2645);
and U2931 (N_2931,N_2752,N_2668);
and U2932 (N_2932,N_2775,N_2776);
or U2933 (N_2933,N_2627,N_2719);
nor U2934 (N_2934,N_2651,N_2702);
and U2935 (N_2935,N_2717,N_2600);
and U2936 (N_2936,N_2603,N_2680);
and U2937 (N_2937,N_2688,N_2672);
or U2938 (N_2938,N_2652,N_2762);
xnor U2939 (N_2939,N_2643,N_2650);
and U2940 (N_2940,N_2738,N_2773);
nand U2941 (N_2941,N_2623,N_2734);
nand U2942 (N_2942,N_2780,N_2670);
nor U2943 (N_2943,N_2738,N_2763);
nand U2944 (N_2944,N_2756,N_2695);
or U2945 (N_2945,N_2696,N_2770);
nand U2946 (N_2946,N_2774,N_2742);
nand U2947 (N_2947,N_2796,N_2605);
or U2948 (N_2948,N_2780,N_2631);
and U2949 (N_2949,N_2610,N_2649);
or U2950 (N_2950,N_2674,N_2643);
or U2951 (N_2951,N_2700,N_2705);
and U2952 (N_2952,N_2737,N_2642);
and U2953 (N_2953,N_2606,N_2709);
nor U2954 (N_2954,N_2656,N_2743);
and U2955 (N_2955,N_2630,N_2654);
nand U2956 (N_2956,N_2699,N_2631);
or U2957 (N_2957,N_2734,N_2681);
nor U2958 (N_2958,N_2781,N_2776);
nor U2959 (N_2959,N_2767,N_2783);
nor U2960 (N_2960,N_2606,N_2782);
and U2961 (N_2961,N_2686,N_2679);
or U2962 (N_2962,N_2717,N_2700);
xor U2963 (N_2963,N_2700,N_2606);
nor U2964 (N_2964,N_2760,N_2608);
nand U2965 (N_2965,N_2707,N_2717);
nor U2966 (N_2966,N_2644,N_2735);
and U2967 (N_2967,N_2682,N_2730);
and U2968 (N_2968,N_2721,N_2789);
or U2969 (N_2969,N_2798,N_2669);
nor U2970 (N_2970,N_2777,N_2766);
or U2971 (N_2971,N_2604,N_2615);
nand U2972 (N_2972,N_2625,N_2676);
or U2973 (N_2973,N_2662,N_2671);
and U2974 (N_2974,N_2663,N_2700);
nor U2975 (N_2975,N_2642,N_2778);
and U2976 (N_2976,N_2771,N_2686);
and U2977 (N_2977,N_2793,N_2681);
or U2978 (N_2978,N_2697,N_2778);
or U2979 (N_2979,N_2743,N_2730);
nand U2980 (N_2980,N_2741,N_2620);
nand U2981 (N_2981,N_2669,N_2771);
nand U2982 (N_2982,N_2730,N_2648);
and U2983 (N_2983,N_2600,N_2611);
or U2984 (N_2984,N_2705,N_2734);
and U2985 (N_2985,N_2621,N_2716);
or U2986 (N_2986,N_2666,N_2766);
or U2987 (N_2987,N_2714,N_2784);
nand U2988 (N_2988,N_2669,N_2687);
nand U2989 (N_2989,N_2655,N_2746);
or U2990 (N_2990,N_2779,N_2676);
and U2991 (N_2991,N_2729,N_2726);
nand U2992 (N_2992,N_2668,N_2783);
nor U2993 (N_2993,N_2614,N_2689);
and U2994 (N_2994,N_2726,N_2767);
xnor U2995 (N_2995,N_2642,N_2707);
or U2996 (N_2996,N_2626,N_2636);
or U2997 (N_2997,N_2640,N_2773);
nor U2998 (N_2998,N_2743,N_2708);
and U2999 (N_2999,N_2606,N_2707);
xor U3000 (N_3000,N_2932,N_2884);
and U3001 (N_3001,N_2915,N_2944);
or U3002 (N_3002,N_2807,N_2968);
or U3003 (N_3003,N_2847,N_2939);
nor U3004 (N_3004,N_2816,N_2806);
nor U3005 (N_3005,N_2888,N_2920);
nand U3006 (N_3006,N_2892,N_2859);
nor U3007 (N_3007,N_2981,N_2809);
nor U3008 (N_3008,N_2900,N_2867);
nand U3009 (N_3009,N_2837,N_2829);
nand U3010 (N_3010,N_2972,N_2985);
nor U3011 (N_3011,N_2827,N_2865);
and U3012 (N_3012,N_2952,N_2903);
nand U3013 (N_3013,N_2820,N_2836);
or U3014 (N_3014,N_2853,N_2995);
or U3015 (N_3015,N_2879,N_2845);
nand U3016 (N_3016,N_2934,N_2860);
nand U3017 (N_3017,N_2902,N_2899);
and U3018 (N_3018,N_2964,N_2931);
and U3019 (N_3019,N_2916,N_2921);
nand U3020 (N_3020,N_2800,N_2925);
or U3021 (N_3021,N_2864,N_2855);
and U3022 (N_3022,N_2835,N_2804);
nor U3023 (N_3023,N_2866,N_2911);
or U3024 (N_3024,N_2828,N_2815);
nor U3025 (N_3025,N_2950,N_2844);
nand U3026 (N_3026,N_2974,N_2830);
xnor U3027 (N_3027,N_2848,N_2989);
nor U3028 (N_3028,N_2923,N_2913);
nand U3029 (N_3029,N_2808,N_2843);
and U3030 (N_3030,N_2849,N_2928);
nor U3031 (N_3031,N_2881,N_2918);
and U3032 (N_3032,N_2980,N_2992);
or U3033 (N_3033,N_2929,N_2873);
or U3034 (N_3034,N_2998,N_2948);
or U3035 (N_3035,N_2838,N_2875);
nand U3036 (N_3036,N_2890,N_2810);
or U3037 (N_3037,N_2924,N_2825);
or U3038 (N_3038,N_2870,N_2941);
nor U3039 (N_3039,N_2993,N_2821);
and U3040 (N_3040,N_2880,N_2930);
nor U3041 (N_3041,N_2937,N_2908);
nor U3042 (N_3042,N_2882,N_2973);
xnor U3043 (N_3043,N_2904,N_2817);
and U3044 (N_3044,N_2874,N_2907);
nand U3045 (N_3045,N_2818,N_2851);
and U3046 (N_3046,N_2905,N_2834);
or U3047 (N_3047,N_2858,N_2802);
or U3048 (N_3048,N_2803,N_2951);
nand U3049 (N_3049,N_2922,N_2927);
nand U3050 (N_3050,N_2906,N_2954);
nand U3051 (N_3051,N_2994,N_2958);
or U3052 (N_3052,N_2957,N_2979);
nor U3053 (N_3053,N_2893,N_2971);
or U3054 (N_3054,N_2987,N_2955);
and U3055 (N_3055,N_2811,N_2831);
and U3056 (N_3056,N_2943,N_2850);
and U3057 (N_3057,N_2871,N_2886);
or U3058 (N_3058,N_2878,N_2986);
nand U3059 (N_3059,N_2909,N_2805);
or U3060 (N_3060,N_2997,N_2938);
nor U3061 (N_3061,N_2833,N_2897);
nand U3062 (N_3062,N_2822,N_2854);
and U3063 (N_3063,N_2935,N_2977);
nand U3064 (N_3064,N_2856,N_2953);
or U3065 (N_3065,N_2872,N_2945);
nand U3066 (N_3066,N_2967,N_2883);
nor U3067 (N_3067,N_2990,N_2869);
nand U3068 (N_3068,N_2975,N_2960);
nor U3069 (N_3069,N_2970,N_2801);
nor U3070 (N_3070,N_2868,N_2912);
nand U3071 (N_3071,N_2963,N_2910);
or U3072 (N_3072,N_2996,N_2876);
nand U3073 (N_3073,N_2946,N_2942);
and U3074 (N_3074,N_2984,N_2824);
or U3075 (N_3075,N_2949,N_2826);
and U3076 (N_3076,N_2917,N_2956);
and U3077 (N_3077,N_2933,N_2962);
or U3078 (N_3078,N_2926,N_2991);
or U3079 (N_3079,N_2919,N_2842);
or U3080 (N_3080,N_2840,N_2969);
and U3081 (N_3081,N_2863,N_2812);
or U3082 (N_3082,N_2940,N_2936);
nand U3083 (N_3083,N_2982,N_2961);
nor U3084 (N_3084,N_2894,N_2999);
and U3085 (N_3085,N_2959,N_2813);
nand U3086 (N_3086,N_2901,N_2841);
or U3087 (N_3087,N_2947,N_2814);
nor U3088 (N_3088,N_2898,N_2839);
nor U3089 (N_3089,N_2852,N_2891);
or U3090 (N_3090,N_2857,N_2978);
nand U3091 (N_3091,N_2846,N_2877);
xnor U3092 (N_3092,N_2983,N_2823);
nand U3093 (N_3093,N_2988,N_2914);
nor U3094 (N_3094,N_2861,N_2976);
nand U3095 (N_3095,N_2832,N_2885);
and U3096 (N_3096,N_2895,N_2966);
nand U3097 (N_3097,N_2889,N_2896);
or U3098 (N_3098,N_2819,N_2862);
nor U3099 (N_3099,N_2965,N_2887);
nor U3100 (N_3100,N_2905,N_2826);
nand U3101 (N_3101,N_2978,N_2877);
nor U3102 (N_3102,N_2817,N_2894);
or U3103 (N_3103,N_2966,N_2885);
nor U3104 (N_3104,N_2994,N_2877);
nor U3105 (N_3105,N_2829,N_2828);
and U3106 (N_3106,N_2958,N_2944);
and U3107 (N_3107,N_2938,N_2840);
or U3108 (N_3108,N_2824,N_2812);
or U3109 (N_3109,N_2994,N_2853);
or U3110 (N_3110,N_2879,N_2886);
nand U3111 (N_3111,N_2960,N_2976);
and U3112 (N_3112,N_2893,N_2922);
and U3113 (N_3113,N_2933,N_2813);
nand U3114 (N_3114,N_2970,N_2919);
nor U3115 (N_3115,N_2858,N_2981);
and U3116 (N_3116,N_2860,N_2835);
and U3117 (N_3117,N_2939,N_2857);
nor U3118 (N_3118,N_2945,N_2995);
or U3119 (N_3119,N_2983,N_2819);
nor U3120 (N_3120,N_2951,N_2967);
nand U3121 (N_3121,N_2869,N_2993);
nor U3122 (N_3122,N_2875,N_2885);
nor U3123 (N_3123,N_2816,N_2955);
nor U3124 (N_3124,N_2971,N_2911);
nand U3125 (N_3125,N_2910,N_2891);
nor U3126 (N_3126,N_2803,N_2813);
and U3127 (N_3127,N_2906,N_2926);
or U3128 (N_3128,N_2832,N_2953);
nand U3129 (N_3129,N_2966,N_2801);
nand U3130 (N_3130,N_2854,N_2887);
nor U3131 (N_3131,N_2977,N_2804);
nor U3132 (N_3132,N_2819,N_2969);
nand U3133 (N_3133,N_2943,N_2895);
nor U3134 (N_3134,N_2852,N_2902);
nand U3135 (N_3135,N_2813,N_2925);
nand U3136 (N_3136,N_2841,N_2892);
nand U3137 (N_3137,N_2872,N_2979);
nand U3138 (N_3138,N_2833,N_2822);
and U3139 (N_3139,N_2994,N_2930);
nand U3140 (N_3140,N_2937,N_2999);
nand U3141 (N_3141,N_2922,N_2992);
nand U3142 (N_3142,N_2884,N_2885);
nor U3143 (N_3143,N_2843,N_2936);
or U3144 (N_3144,N_2898,N_2949);
nand U3145 (N_3145,N_2873,N_2820);
nand U3146 (N_3146,N_2952,N_2885);
nand U3147 (N_3147,N_2997,N_2817);
nand U3148 (N_3148,N_2833,N_2886);
nor U3149 (N_3149,N_2973,N_2827);
or U3150 (N_3150,N_2945,N_2814);
xnor U3151 (N_3151,N_2832,N_2874);
or U3152 (N_3152,N_2923,N_2802);
nand U3153 (N_3153,N_2931,N_2988);
and U3154 (N_3154,N_2953,N_2829);
nor U3155 (N_3155,N_2988,N_2871);
nand U3156 (N_3156,N_2908,N_2942);
and U3157 (N_3157,N_2961,N_2905);
nand U3158 (N_3158,N_2925,N_2978);
nand U3159 (N_3159,N_2808,N_2961);
nand U3160 (N_3160,N_2855,N_2950);
nand U3161 (N_3161,N_2886,N_2812);
or U3162 (N_3162,N_2977,N_2885);
nor U3163 (N_3163,N_2901,N_2879);
or U3164 (N_3164,N_2802,N_2972);
nand U3165 (N_3165,N_2864,N_2867);
nand U3166 (N_3166,N_2834,N_2822);
or U3167 (N_3167,N_2835,N_2874);
or U3168 (N_3168,N_2801,N_2883);
nor U3169 (N_3169,N_2861,N_2808);
nor U3170 (N_3170,N_2895,N_2886);
nand U3171 (N_3171,N_2902,N_2989);
and U3172 (N_3172,N_2859,N_2801);
nand U3173 (N_3173,N_2836,N_2807);
or U3174 (N_3174,N_2964,N_2822);
nor U3175 (N_3175,N_2824,N_2801);
nor U3176 (N_3176,N_2807,N_2863);
xnor U3177 (N_3177,N_2828,N_2825);
or U3178 (N_3178,N_2937,N_2912);
nor U3179 (N_3179,N_2920,N_2840);
and U3180 (N_3180,N_2984,N_2906);
or U3181 (N_3181,N_2910,N_2892);
or U3182 (N_3182,N_2827,N_2848);
nand U3183 (N_3183,N_2886,N_2965);
nor U3184 (N_3184,N_2924,N_2976);
and U3185 (N_3185,N_2829,N_2806);
or U3186 (N_3186,N_2966,N_2841);
nor U3187 (N_3187,N_2899,N_2981);
nand U3188 (N_3188,N_2980,N_2939);
or U3189 (N_3189,N_2922,N_2907);
and U3190 (N_3190,N_2902,N_2813);
nand U3191 (N_3191,N_2840,N_2949);
nand U3192 (N_3192,N_2870,N_2806);
or U3193 (N_3193,N_2997,N_2876);
and U3194 (N_3194,N_2956,N_2918);
or U3195 (N_3195,N_2916,N_2855);
or U3196 (N_3196,N_2895,N_2923);
nand U3197 (N_3197,N_2967,N_2970);
or U3198 (N_3198,N_2828,N_2850);
or U3199 (N_3199,N_2840,N_2828);
nor U3200 (N_3200,N_3073,N_3138);
nand U3201 (N_3201,N_3025,N_3186);
nor U3202 (N_3202,N_3074,N_3049);
and U3203 (N_3203,N_3008,N_3188);
nor U3204 (N_3204,N_3195,N_3164);
or U3205 (N_3205,N_3129,N_3178);
nand U3206 (N_3206,N_3004,N_3193);
and U3207 (N_3207,N_3168,N_3132);
or U3208 (N_3208,N_3190,N_3034);
nand U3209 (N_3209,N_3179,N_3023);
nand U3210 (N_3210,N_3029,N_3010);
and U3211 (N_3211,N_3069,N_3050);
nor U3212 (N_3212,N_3169,N_3128);
nor U3213 (N_3213,N_3007,N_3058);
nand U3214 (N_3214,N_3119,N_3006);
and U3215 (N_3215,N_3002,N_3101);
nor U3216 (N_3216,N_3198,N_3114);
and U3217 (N_3217,N_3012,N_3059);
or U3218 (N_3218,N_3135,N_3160);
or U3219 (N_3219,N_3127,N_3071);
nand U3220 (N_3220,N_3107,N_3123);
or U3221 (N_3221,N_3094,N_3156);
nor U3222 (N_3222,N_3053,N_3180);
or U3223 (N_3223,N_3040,N_3104);
or U3224 (N_3224,N_3052,N_3078);
nor U3225 (N_3225,N_3185,N_3153);
nor U3226 (N_3226,N_3175,N_3191);
and U3227 (N_3227,N_3054,N_3147);
and U3228 (N_3228,N_3083,N_3192);
nand U3229 (N_3229,N_3019,N_3072);
nor U3230 (N_3230,N_3044,N_3144);
and U3231 (N_3231,N_3009,N_3171);
nand U3232 (N_3232,N_3056,N_3199);
or U3233 (N_3233,N_3027,N_3082);
and U3234 (N_3234,N_3124,N_3063);
nor U3235 (N_3235,N_3174,N_3099);
or U3236 (N_3236,N_3084,N_3194);
and U3237 (N_3237,N_3172,N_3041);
nand U3238 (N_3238,N_3045,N_3140);
and U3239 (N_3239,N_3105,N_3079);
nand U3240 (N_3240,N_3157,N_3116);
nor U3241 (N_3241,N_3035,N_3061);
nor U3242 (N_3242,N_3043,N_3089);
nand U3243 (N_3243,N_3076,N_3005);
nor U3244 (N_3244,N_3154,N_3096);
or U3245 (N_3245,N_3048,N_3130);
nand U3246 (N_3246,N_3015,N_3032);
xor U3247 (N_3247,N_3093,N_3000);
nor U3248 (N_3248,N_3021,N_3117);
nand U3249 (N_3249,N_3057,N_3031);
and U3250 (N_3250,N_3095,N_3163);
or U3251 (N_3251,N_3003,N_3033);
nor U3252 (N_3252,N_3197,N_3017);
or U3253 (N_3253,N_3039,N_3110);
or U3254 (N_3254,N_3088,N_3139);
nor U3255 (N_3255,N_3155,N_3108);
nand U3256 (N_3256,N_3065,N_3067);
xnor U3257 (N_3257,N_3134,N_3036);
nand U3258 (N_3258,N_3196,N_3150);
nand U3259 (N_3259,N_3176,N_3136);
and U3260 (N_3260,N_3022,N_3149);
or U3261 (N_3261,N_3014,N_3001);
nand U3262 (N_3262,N_3080,N_3087);
nor U3263 (N_3263,N_3024,N_3030);
or U3264 (N_3264,N_3097,N_3189);
nand U3265 (N_3265,N_3181,N_3055);
nor U3266 (N_3266,N_3018,N_3103);
nand U3267 (N_3267,N_3081,N_3133);
nand U3268 (N_3268,N_3098,N_3091);
nor U3269 (N_3269,N_3020,N_3026);
nor U3270 (N_3270,N_3062,N_3166);
or U3271 (N_3271,N_3120,N_3085);
nand U3272 (N_3272,N_3141,N_3060);
xor U3273 (N_3273,N_3028,N_3106);
or U3274 (N_3274,N_3038,N_3162);
nand U3275 (N_3275,N_3143,N_3077);
nand U3276 (N_3276,N_3145,N_3161);
nand U3277 (N_3277,N_3075,N_3126);
nand U3278 (N_3278,N_3151,N_3064);
nand U3279 (N_3279,N_3152,N_3148);
or U3280 (N_3280,N_3170,N_3070);
or U3281 (N_3281,N_3165,N_3125);
or U3282 (N_3282,N_3158,N_3068);
or U3283 (N_3283,N_3173,N_3090);
nand U3284 (N_3284,N_3066,N_3146);
nand U3285 (N_3285,N_3086,N_3118);
and U3286 (N_3286,N_3142,N_3037);
or U3287 (N_3287,N_3159,N_3112);
nor U3288 (N_3288,N_3182,N_3137);
nand U3289 (N_3289,N_3115,N_3121);
or U3290 (N_3290,N_3187,N_3016);
and U3291 (N_3291,N_3047,N_3100);
nand U3292 (N_3292,N_3131,N_3122);
nor U3293 (N_3293,N_3102,N_3184);
or U3294 (N_3294,N_3183,N_3092);
nor U3295 (N_3295,N_3177,N_3113);
and U3296 (N_3296,N_3042,N_3109);
and U3297 (N_3297,N_3011,N_3046);
nand U3298 (N_3298,N_3167,N_3013);
nor U3299 (N_3299,N_3111,N_3051);
nor U3300 (N_3300,N_3003,N_3009);
nor U3301 (N_3301,N_3188,N_3002);
or U3302 (N_3302,N_3012,N_3017);
nor U3303 (N_3303,N_3162,N_3052);
nand U3304 (N_3304,N_3005,N_3159);
nor U3305 (N_3305,N_3151,N_3026);
nor U3306 (N_3306,N_3196,N_3039);
or U3307 (N_3307,N_3121,N_3036);
nand U3308 (N_3308,N_3025,N_3093);
nor U3309 (N_3309,N_3136,N_3148);
and U3310 (N_3310,N_3139,N_3194);
and U3311 (N_3311,N_3067,N_3186);
nor U3312 (N_3312,N_3036,N_3168);
xor U3313 (N_3313,N_3027,N_3179);
nand U3314 (N_3314,N_3089,N_3148);
nand U3315 (N_3315,N_3176,N_3161);
nor U3316 (N_3316,N_3031,N_3006);
and U3317 (N_3317,N_3074,N_3107);
and U3318 (N_3318,N_3146,N_3137);
nand U3319 (N_3319,N_3167,N_3131);
nand U3320 (N_3320,N_3076,N_3157);
or U3321 (N_3321,N_3172,N_3158);
or U3322 (N_3322,N_3009,N_3032);
nor U3323 (N_3323,N_3135,N_3174);
and U3324 (N_3324,N_3129,N_3197);
or U3325 (N_3325,N_3015,N_3029);
or U3326 (N_3326,N_3097,N_3000);
or U3327 (N_3327,N_3140,N_3092);
or U3328 (N_3328,N_3133,N_3068);
nand U3329 (N_3329,N_3143,N_3092);
xnor U3330 (N_3330,N_3153,N_3194);
or U3331 (N_3331,N_3087,N_3075);
or U3332 (N_3332,N_3021,N_3087);
nor U3333 (N_3333,N_3135,N_3129);
and U3334 (N_3334,N_3175,N_3021);
nor U3335 (N_3335,N_3102,N_3034);
nand U3336 (N_3336,N_3105,N_3183);
or U3337 (N_3337,N_3029,N_3067);
or U3338 (N_3338,N_3185,N_3089);
nor U3339 (N_3339,N_3146,N_3197);
nor U3340 (N_3340,N_3112,N_3158);
nor U3341 (N_3341,N_3118,N_3114);
or U3342 (N_3342,N_3038,N_3176);
nor U3343 (N_3343,N_3075,N_3169);
or U3344 (N_3344,N_3132,N_3024);
nand U3345 (N_3345,N_3188,N_3122);
nor U3346 (N_3346,N_3082,N_3073);
and U3347 (N_3347,N_3131,N_3100);
or U3348 (N_3348,N_3171,N_3031);
xor U3349 (N_3349,N_3176,N_3107);
or U3350 (N_3350,N_3159,N_3182);
and U3351 (N_3351,N_3144,N_3025);
nand U3352 (N_3352,N_3010,N_3018);
nor U3353 (N_3353,N_3064,N_3007);
or U3354 (N_3354,N_3084,N_3167);
nand U3355 (N_3355,N_3139,N_3125);
nor U3356 (N_3356,N_3090,N_3040);
or U3357 (N_3357,N_3034,N_3189);
and U3358 (N_3358,N_3096,N_3152);
and U3359 (N_3359,N_3116,N_3161);
or U3360 (N_3360,N_3052,N_3088);
or U3361 (N_3361,N_3062,N_3093);
or U3362 (N_3362,N_3186,N_3166);
and U3363 (N_3363,N_3074,N_3192);
nor U3364 (N_3364,N_3011,N_3018);
nor U3365 (N_3365,N_3148,N_3004);
and U3366 (N_3366,N_3150,N_3159);
and U3367 (N_3367,N_3135,N_3057);
and U3368 (N_3368,N_3094,N_3124);
and U3369 (N_3369,N_3090,N_3023);
or U3370 (N_3370,N_3127,N_3157);
or U3371 (N_3371,N_3141,N_3154);
or U3372 (N_3372,N_3150,N_3084);
nor U3373 (N_3373,N_3123,N_3194);
nand U3374 (N_3374,N_3175,N_3129);
nor U3375 (N_3375,N_3086,N_3180);
and U3376 (N_3376,N_3145,N_3019);
xnor U3377 (N_3377,N_3093,N_3075);
nor U3378 (N_3378,N_3010,N_3013);
or U3379 (N_3379,N_3003,N_3049);
and U3380 (N_3380,N_3090,N_3059);
and U3381 (N_3381,N_3049,N_3154);
or U3382 (N_3382,N_3066,N_3004);
nand U3383 (N_3383,N_3194,N_3176);
nand U3384 (N_3384,N_3004,N_3168);
and U3385 (N_3385,N_3133,N_3042);
or U3386 (N_3386,N_3150,N_3112);
nor U3387 (N_3387,N_3079,N_3002);
or U3388 (N_3388,N_3012,N_3123);
or U3389 (N_3389,N_3104,N_3087);
nor U3390 (N_3390,N_3043,N_3133);
nor U3391 (N_3391,N_3068,N_3161);
nor U3392 (N_3392,N_3034,N_3139);
nand U3393 (N_3393,N_3087,N_3041);
and U3394 (N_3394,N_3064,N_3036);
or U3395 (N_3395,N_3103,N_3056);
nand U3396 (N_3396,N_3141,N_3019);
and U3397 (N_3397,N_3033,N_3022);
xor U3398 (N_3398,N_3072,N_3023);
nand U3399 (N_3399,N_3017,N_3087);
nor U3400 (N_3400,N_3363,N_3288);
nor U3401 (N_3401,N_3371,N_3311);
and U3402 (N_3402,N_3294,N_3259);
and U3403 (N_3403,N_3337,N_3367);
or U3404 (N_3404,N_3340,N_3204);
nand U3405 (N_3405,N_3347,N_3332);
or U3406 (N_3406,N_3290,N_3201);
nand U3407 (N_3407,N_3235,N_3368);
nand U3408 (N_3408,N_3260,N_3310);
or U3409 (N_3409,N_3345,N_3309);
and U3410 (N_3410,N_3273,N_3252);
or U3411 (N_3411,N_3227,N_3276);
nor U3412 (N_3412,N_3391,N_3268);
nor U3413 (N_3413,N_3356,N_3314);
or U3414 (N_3414,N_3326,N_3302);
nand U3415 (N_3415,N_3343,N_3240);
nor U3416 (N_3416,N_3202,N_3389);
nand U3417 (N_3417,N_3321,N_3362);
or U3418 (N_3418,N_3366,N_3306);
nand U3419 (N_3419,N_3346,N_3331);
or U3420 (N_3420,N_3258,N_3219);
or U3421 (N_3421,N_3298,N_3315);
nand U3422 (N_3422,N_3358,N_3220);
xor U3423 (N_3423,N_3323,N_3297);
or U3424 (N_3424,N_3262,N_3365);
nor U3425 (N_3425,N_3399,N_3300);
nor U3426 (N_3426,N_3206,N_3388);
nor U3427 (N_3427,N_3247,N_3378);
nand U3428 (N_3428,N_3211,N_3242);
nor U3429 (N_3429,N_3316,N_3210);
or U3430 (N_3430,N_3243,N_3231);
nand U3431 (N_3431,N_3244,N_3233);
and U3432 (N_3432,N_3359,N_3364);
and U3433 (N_3433,N_3215,N_3327);
nand U3434 (N_3434,N_3301,N_3248);
or U3435 (N_3435,N_3349,N_3223);
nor U3436 (N_3436,N_3336,N_3353);
nor U3437 (N_3437,N_3373,N_3269);
nand U3438 (N_3438,N_3267,N_3305);
nand U3439 (N_3439,N_3376,N_3312);
nor U3440 (N_3440,N_3387,N_3313);
and U3441 (N_3441,N_3357,N_3380);
nand U3442 (N_3442,N_3350,N_3338);
nor U3443 (N_3443,N_3341,N_3304);
nand U3444 (N_3444,N_3342,N_3249);
and U3445 (N_3445,N_3214,N_3246);
nand U3446 (N_3446,N_3395,N_3281);
nor U3447 (N_3447,N_3284,N_3217);
and U3448 (N_3448,N_3381,N_3320);
nand U3449 (N_3449,N_3209,N_3299);
or U3450 (N_3450,N_3228,N_3216);
or U3451 (N_3451,N_3295,N_3285);
nand U3452 (N_3452,N_3329,N_3339);
nor U3453 (N_3453,N_3351,N_3270);
or U3454 (N_3454,N_3344,N_3212);
nor U3455 (N_3455,N_3397,N_3287);
nor U3456 (N_3456,N_3334,N_3232);
or U3457 (N_3457,N_3279,N_3335);
nor U3458 (N_3458,N_3251,N_3348);
or U3459 (N_3459,N_3322,N_3318);
xor U3460 (N_3460,N_3245,N_3272);
xor U3461 (N_3461,N_3250,N_3317);
nand U3462 (N_3462,N_3255,N_3271);
nor U3463 (N_3463,N_3325,N_3375);
nand U3464 (N_3464,N_3328,N_3278);
or U3465 (N_3465,N_3225,N_3222);
nor U3466 (N_3466,N_3283,N_3239);
nand U3467 (N_3467,N_3370,N_3354);
nor U3468 (N_3468,N_3324,N_3352);
and U3469 (N_3469,N_3254,N_3307);
nor U3470 (N_3470,N_3208,N_3280);
and U3471 (N_3471,N_3286,N_3275);
and U3472 (N_3472,N_3390,N_3277);
nand U3473 (N_3473,N_3253,N_3385);
nor U3474 (N_3474,N_3213,N_3374);
nand U3475 (N_3475,N_3221,N_3382);
nor U3476 (N_3476,N_3257,N_3224);
nand U3477 (N_3477,N_3355,N_3282);
or U3478 (N_3478,N_3308,N_3393);
nor U3479 (N_3479,N_3296,N_3203);
and U3480 (N_3480,N_3234,N_3265);
nor U3481 (N_3481,N_3372,N_3200);
nor U3482 (N_3482,N_3377,N_3333);
nor U3483 (N_3483,N_3379,N_3266);
or U3484 (N_3484,N_3207,N_3291);
or U3485 (N_3485,N_3237,N_3261);
and U3486 (N_3486,N_3386,N_3274);
nand U3487 (N_3487,N_3292,N_3319);
nand U3488 (N_3488,N_3238,N_3236);
and U3489 (N_3489,N_3230,N_3289);
and U3490 (N_3490,N_3384,N_3229);
and U3491 (N_3491,N_3293,N_3361);
xor U3492 (N_3492,N_3330,N_3241);
nand U3493 (N_3493,N_3264,N_3360);
or U3494 (N_3494,N_3398,N_3263);
or U3495 (N_3495,N_3396,N_3218);
nor U3496 (N_3496,N_3369,N_3392);
nand U3497 (N_3497,N_3256,N_3205);
or U3498 (N_3498,N_3303,N_3383);
nor U3499 (N_3499,N_3226,N_3394);
or U3500 (N_3500,N_3225,N_3300);
nand U3501 (N_3501,N_3323,N_3200);
xnor U3502 (N_3502,N_3359,N_3288);
or U3503 (N_3503,N_3330,N_3263);
nand U3504 (N_3504,N_3323,N_3221);
nor U3505 (N_3505,N_3225,N_3211);
or U3506 (N_3506,N_3332,N_3217);
or U3507 (N_3507,N_3365,N_3225);
nand U3508 (N_3508,N_3353,N_3378);
or U3509 (N_3509,N_3272,N_3213);
or U3510 (N_3510,N_3228,N_3201);
nor U3511 (N_3511,N_3311,N_3258);
nand U3512 (N_3512,N_3237,N_3254);
nand U3513 (N_3513,N_3366,N_3229);
or U3514 (N_3514,N_3397,N_3238);
nor U3515 (N_3515,N_3335,N_3282);
and U3516 (N_3516,N_3265,N_3352);
nor U3517 (N_3517,N_3272,N_3294);
or U3518 (N_3518,N_3394,N_3255);
nand U3519 (N_3519,N_3257,N_3200);
and U3520 (N_3520,N_3220,N_3371);
nand U3521 (N_3521,N_3221,N_3347);
nand U3522 (N_3522,N_3308,N_3389);
and U3523 (N_3523,N_3252,N_3340);
and U3524 (N_3524,N_3363,N_3221);
nor U3525 (N_3525,N_3305,N_3333);
and U3526 (N_3526,N_3239,N_3204);
nor U3527 (N_3527,N_3282,N_3306);
nor U3528 (N_3528,N_3201,N_3226);
nand U3529 (N_3529,N_3314,N_3341);
nand U3530 (N_3530,N_3234,N_3299);
and U3531 (N_3531,N_3343,N_3261);
and U3532 (N_3532,N_3399,N_3309);
and U3533 (N_3533,N_3381,N_3263);
or U3534 (N_3534,N_3327,N_3286);
and U3535 (N_3535,N_3314,N_3359);
nand U3536 (N_3536,N_3335,N_3315);
and U3537 (N_3537,N_3300,N_3363);
nor U3538 (N_3538,N_3282,N_3349);
nand U3539 (N_3539,N_3287,N_3382);
or U3540 (N_3540,N_3268,N_3265);
and U3541 (N_3541,N_3249,N_3377);
or U3542 (N_3542,N_3224,N_3370);
and U3543 (N_3543,N_3271,N_3222);
or U3544 (N_3544,N_3208,N_3322);
and U3545 (N_3545,N_3219,N_3372);
or U3546 (N_3546,N_3218,N_3342);
and U3547 (N_3547,N_3249,N_3270);
or U3548 (N_3548,N_3232,N_3285);
nand U3549 (N_3549,N_3386,N_3282);
nor U3550 (N_3550,N_3233,N_3293);
nor U3551 (N_3551,N_3253,N_3240);
or U3552 (N_3552,N_3240,N_3260);
and U3553 (N_3553,N_3229,N_3236);
or U3554 (N_3554,N_3226,N_3211);
and U3555 (N_3555,N_3346,N_3271);
and U3556 (N_3556,N_3381,N_3275);
nand U3557 (N_3557,N_3313,N_3304);
and U3558 (N_3558,N_3325,N_3296);
and U3559 (N_3559,N_3273,N_3383);
nor U3560 (N_3560,N_3298,N_3364);
nor U3561 (N_3561,N_3316,N_3319);
nor U3562 (N_3562,N_3328,N_3256);
xor U3563 (N_3563,N_3386,N_3296);
nand U3564 (N_3564,N_3306,N_3319);
nand U3565 (N_3565,N_3374,N_3372);
or U3566 (N_3566,N_3326,N_3328);
nand U3567 (N_3567,N_3217,N_3307);
nor U3568 (N_3568,N_3268,N_3240);
and U3569 (N_3569,N_3334,N_3386);
nand U3570 (N_3570,N_3360,N_3285);
nand U3571 (N_3571,N_3381,N_3329);
and U3572 (N_3572,N_3324,N_3330);
and U3573 (N_3573,N_3312,N_3330);
or U3574 (N_3574,N_3372,N_3261);
nor U3575 (N_3575,N_3346,N_3294);
or U3576 (N_3576,N_3207,N_3341);
nor U3577 (N_3577,N_3309,N_3248);
or U3578 (N_3578,N_3264,N_3242);
nor U3579 (N_3579,N_3290,N_3212);
nand U3580 (N_3580,N_3371,N_3378);
and U3581 (N_3581,N_3397,N_3361);
and U3582 (N_3582,N_3204,N_3359);
nor U3583 (N_3583,N_3291,N_3322);
or U3584 (N_3584,N_3231,N_3399);
and U3585 (N_3585,N_3264,N_3385);
and U3586 (N_3586,N_3379,N_3381);
nand U3587 (N_3587,N_3294,N_3205);
and U3588 (N_3588,N_3383,N_3379);
nor U3589 (N_3589,N_3334,N_3303);
or U3590 (N_3590,N_3354,N_3230);
nand U3591 (N_3591,N_3326,N_3307);
nand U3592 (N_3592,N_3367,N_3319);
or U3593 (N_3593,N_3208,N_3254);
and U3594 (N_3594,N_3255,N_3233);
nand U3595 (N_3595,N_3322,N_3298);
nor U3596 (N_3596,N_3201,N_3296);
and U3597 (N_3597,N_3372,N_3379);
nand U3598 (N_3598,N_3266,N_3372);
or U3599 (N_3599,N_3317,N_3307);
nand U3600 (N_3600,N_3466,N_3573);
nand U3601 (N_3601,N_3443,N_3403);
nand U3602 (N_3602,N_3490,N_3464);
or U3603 (N_3603,N_3459,N_3432);
and U3604 (N_3604,N_3502,N_3436);
nand U3605 (N_3605,N_3518,N_3472);
and U3606 (N_3606,N_3590,N_3587);
and U3607 (N_3607,N_3450,N_3461);
and U3608 (N_3608,N_3441,N_3408);
nand U3609 (N_3609,N_3440,N_3560);
nor U3610 (N_3610,N_3534,N_3539);
nor U3611 (N_3611,N_3444,N_3582);
and U3612 (N_3612,N_3484,N_3498);
nor U3613 (N_3613,N_3427,N_3561);
or U3614 (N_3614,N_3467,N_3419);
nand U3615 (N_3615,N_3423,N_3562);
and U3616 (N_3616,N_3533,N_3412);
nand U3617 (N_3617,N_3433,N_3566);
or U3618 (N_3618,N_3445,N_3485);
nor U3619 (N_3619,N_3448,N_3487);
nand U3620 (N_3620,N_3543,N_3532);
and U3621 (N_3621,N_3486,N_3557);
and U3622 (N_3622,N_3411,N_3535);
nor U3623 (N_3623,N_3591,N_3507);
nor U3624 (N_3624,N_3586,N_3559);
nor U3625 (N_3625,N_3402,N_3439);
or U3626 (N_3626,N_3584,N_3568);
or U3627 (N_3627,N_3465,N_3596);
and U3628 (N_3628,N_3552,N_3531);
nor U3629 (N_3629,N_3434,N_3455);
and U3630 (N_3630,N_3580,N_3567);
or U3631 (N_3631,N_3544,N_3488);
nor U3632 (N_3632,N_3469,N_3482);
and U3633 (N_3633,N_3574,N_3504);
and U3634 (N_3634,N_3447,N_3516);
nor U3635 (N_3635,N_3569,N_3506);
nor U3636 (N_3636,N_3478,N_3548);
and U3637 (N_3637,N_3442,N_3483);
nor U3638 (N_3638,N_3514,N_3409);
nand U3639 (N_3639,N_3546,N_3416);
nand U3640 (N_3640,N_3576,N_3500);
and U3641 (N_3641,N_3431,N_3474);
nand U3642 (N_3642,N_3457,N_3446);
nor U3643 (N_3643,N_3594,N_3541);
nand U3644 (N_3644,N_3425,N_3463);
nand U3645 (N_3645,N_3523,N_3493);
nor U3646 (N_3646,N_3526,N_3537);
or U3647 (N_3647,N_3542,N_3400);
and U3648 (N_3648,N_3565,N_3499);
nor U3649 (N_3649,N_3522,N_3401);
nor U3650 (N_3650,N_3492,N_3438);
xor U3651 (N_3651,N_3406,N_3420);
nand U3652 (N_3652,N_3512,N_3525);
nand U3653 (N_3653,N_3451,N_3413);
and U3654 (N_3654,N_3527,N_3536);
nand U3655 (N_3655,N_3480,N_3583);
and U3656 (N_3656,N_3599,N_3538);
nor U3657 (N_3657,N_3564,N_3579);
or U3658 (N_3658,N_3481,N_3404);
and U3659 (N_3659,N_3460,N_3515);
and U3660 (N_3660,N_3456,N_3475);
nand U3661 (N_3661,N_3571,N_3572);
nand U3662 (N_3662,N_3593,N_3553);
or U3663 (N_3663,N_3528,N_3556);
or U3664 (N_3664,N_3417,N_3428);
or U3665 (N_3665,N_3554,N_3421);
nor U3666 (N_3666,N_3578,N_3414);
nor U3667 (N_3667,N_3549,N_3517);
or U3668 (N_3668,N_3415,N_3510);
nand U3669 (N_3669,N_3477,N_3430);
or U3670 (N_3670,N_3422,N_3470);
or U3671 (N_3671,N_3407,N_3476);
xnor U3672 (N_3672,N_3563,N_3452);
and U3673 (N_3673,N_3503,N_3429);
and U3674 (N_3674,N_3405,N_3454);
and U3675 (N_3675,N_3530,N_3589);
and U3676 (N_3676,N_3437,N_3435);
nand U3677 (N_3677,N_3551,N_3426);
nand U3678 (N_3678,N_3509,N_3462);
or U3679 (N_3679,N_3555,N_3592);
nor U3680 (N_3680,N_3453,N_3575);
nand U3681 (N_3681,N_3496,N_3540);
or U3682 (N_3682,N_3570,N_3519);
or U3683 (N_3683,N_3558,N_3550);
or U3684 (N_3684,N_3491,N_3468);
nor U3685 (N_3685,N_3513,N_3505);
nand U3686 (N_3686,N_3424,N_3501);
or U3687 (N_3687,N_3529,N_3458);
nand U3688 (N_3688,N_3479,N_3577);
or U3689 (N_3689,N_3495,N_3597);
and U3690 (N_3690,N_3521,N_3494);
nor U3691 (N_3691,N_3581,N_3511);
and U3692 (N_3692,N_3508,N_3520);
and U3693 (N_3693,N_3595,N_3588);
nor U3694 (N_3694,N_3418,N_3497);
and U3695 (N_3695,N_3524,N_3545);
nor U3696 (N_3696,N_3598,N_3473);
or U3697 (N_3697,N_3471,N_3449);
nand U3698 (N_3698,N_3547,N_3585);
and U3699 (N_3699,N_3410,N_3489);
and U3700 (N_3700,N_3565,N_3521);
and U3701 (N_3701,N_3566,N_3589);
nor U3702 (N_3702,N_3416,N_3570);
or U3703 (N_3703,N_3457,N_3479);
and U3704 (N_3704,N_3542,N_3591);
and U3705 (N_3705,N_3421,N_3401);
and U3706 (N_3706,N_3581,N_3538);
and U3707 (N_3707,N_3534,N_3439);
nand U3708 (N_3708,N_3475,N_3444);
nand U3709 (N_3709,N_3537,N_3543);
and U3710 (N_3710,N_3489,N_3464);
nand U3711 (N_3711,N_3480,N_3407);
or U3712 (N_3712,N_3466,N_3440);
or U3713 (N_3713,N_3520,N_3567);
nor U3714 (N_3714,N_3588,N_3518);
nor U3715 (N_3715,N_3536,N_3508);
nand U3716 (N_3716,N_3446,N_3518);
nor U3717 (N_3717,N_3502,N_3551);
nor U3718 (N_3718,N_3487,N_3471);
or U3719 (N_3719,N_3465,N_3458);
or U3720 (N_3720,N_3428,N_3544);
nor U3721 (N_3721,N_3522,N_3564);
nand U3722 (N_3722,N_3437,N_3428);
or U3723 (N_3723,N_3582,N_3500);
nor U3724 (N_3724,N_3471,N_3575);
or U3725 (N_3725,N_3430,N_3517);
and U3726 (N_3726,N_3484,N_3521);
or U3727 (N_3727,N_3540,N_3421);
xnor U3728 (N_3728,N_3522,N_3484);
or U3729 (N_3729,N_3582,N_3537);
nor U3730 (N_3730,N_3462,N_3517);
or U3731 (N_3731,N_3452,N_3559);
or U3732 (N_3732,N_3537,N_3585);
and U3733 (N_3733,N_3595,N_3477);
and U3734 (N_3734,N_3575,N_3526);
and U3735 (N_3735,N_3408,N_3529);
and U3736 (N_3736,N_3551,N_3444);
or U3737 (N_3737,N_3584,N_3535);
or U3738 (N_3738,N_3432,N_3537);
or U3739 (N_3739,N_3412,N_3577);
and U3740 (N_3740,N_3421,N_3587);
nor U3741 (N_3741,N_3457,N_3535);
nor U3742 (N_3742,N_3447,N_3473);
nand U3743 (N_3743,N_3536,N_3529);
nor U3744 (N_3744,N_3585,N_3517);
nand U3745 (N_3745,N_3586,N_3577);
and U3746 (N_3746,N_3518,N_3476);
and U3747 (N_3747,N_3548,N_3450);
and U3748 (N_3748,N_3414,N_3594);
xor U3749 (N_3749,N_3411,N_3454);
or U3750 (N_3750,N_3557,N_3583);
and U3751 (N_3751,N_3497,N_3529);
and U3752 (N_3752,N_3418,N_3531);
nor U3753 (N_3753,N_3553,N_3444);
nand U3754 (N_3754,N_3524,N_3581);
or U3755 (N_3755,N_3596,N_3400);
nand U3756 (N_3756,N_3534,N_3596);
nand U3757 (N_3757,N_3515,N_3468);
nor U3758 (N_3758,N_3427,N_3506);
or U3759 (N_3759,N_3537,N_3542);
and U3760 (N_3760,N_3433,N_3510);
nand U3761 (N_3761,N_3442,N_3511);
nor U3762 (N_3762,N_3462,N_3482);
or U3763 (N_3763,N_3505,N_3558);
nand U3764 (N_3764,N_3545,N_3488);
nand U3765 (N_3765,N_3447,N_3579);
or U3766 (N_3766,N_3420,N_3533);
nor U3767 (N_3767,N_3589,N_3410);
nand U3768 (N_3768,N_3531,N_3550);
or U3769 (N_3769,N_3455,N_3467);
nor U3770 (N_3770,N_3554,N_3437);
nand U3771 (N_3771,N_3572,N_3563);
and U3772 (N_3772,N_3419,N_3499);
or U3773 (N_3773,N_3474,N_3575);
or U3774 (N_3774,N_3553,N_3485);
and U3775 (N_3775,N_3411,N_3459);
or U3776 (N_3776,N_3521,N_3441);
or U3777 (N_3777,N_3585,N_3576);
nor U3778 (N_3778,N_3426,N_3491);
and U3779 (N_3779,N_3513,N_3582);
nor U3780 (N_3780,N_3597,N_3541);
or U3781 (N_3781,N_3588,N_3543);
xnor U3782 (N_3782,N_3456,N_3413);
and U3783 (N_3783,N_3492,N_3567);
nor U3784 (N_3784,N_3408,N_3492);
nor U3785 (N_3785,N_3454,N_3472);
and U3786 (N_3786,N_3527,N_3552);
nor U3787 (N_3787,N_3470,N_3531);
or U3788 (N_3788,N_3407,N_3433);
nor U3789 (N_3789,N_3528,N_3427);
nand U3790 (N_3790,N_3516,N_3428);
nor U3791 (N_3791,N_3498,N_3577);
and U3792 (N_3792,N_3495,N_3498);
nor U3793 (N_3793,N_3489,N_3496);
nand U3794 (N_3794,N_3472,N_3453);
and U3795 (N_3795,N_3429,N_3448);
and U3796 (N_3796,N_3422,N_3428);
nand U3797 (N_3797,N_3595,N_3513);
and U3798 (N_3798,N_3431,N_3435);
nand U3799 (N_3799,N_3438,N_3553);
and U3800 (N_3800,N_3745,N_3682);
xor U3801 (N_3801,N_3740,N_3760);
and U3802 (N_3802,N_3652,N_3757);
nor U3803 (N_3803,N_3704,N_3731);
or U3804 (N_3804,N_3642,N_3724);
nor U3805 (N_3805,N_3636,N_3791);
nand U3806 (N_3806,N_3606,N_3735);
nor U3807 (N_3807,N_3696,N_3793);
and U3808 (N_3808,N_3644,N_3756);
or U3809 (N_3809,N_3738,N_3621);
nor U3810 (N_3810,N_3774,N_3714);
nand U3811 (N_3811,N_3732,N_3773);
nor U3812 (N_3812,N_3695,N_3656);
nor U3813 (N_3813,N_3789,N_3675);
nand U3814 (N_3814,N_3726,N_3790);
nand U3815 (N_3815,N_3612,N_3669);
or U3816 (N_3816,N_3658,N_3622);
nor U3817 (N_3817,N_3602,N_3619);
and U3818 (N_3818,N_3637,N_3722);
or U3819 (N_3819,N_3625,N_3672);
or U3820 (N_3820,N_3787,N_3650);
nand U3821 (N_3821,N_3721,N_3635);
or U3822 (N_3822,N_3616,N_3706);
nand U3823 (N_3823,N_3786,N_3799);
and U3824 (N_3824,N_3605,N_3788);
nand U3825 (N_3825,N_3729,N_3678);
or U3826 (N_3826,N_3780,N_3700);
nand U3827 (N_3827,N_3633,N_3727);
or U3828 (N_3828,N_3664,N_3628);
nand U3829 (N_3829,N_3614,N_3660);
or U3830 (N_3830,N_3734,N_3776);
nor U3831 (N_3831,N_3792,N_3610);
nor U3832 (N_3832,N_3781,N_3620);
nand U3833 (N_3833,N_3618,N_3691);
and U3834 (N_3834,N_3778,N_3643);
or U3835 (N_3835,N_3654,N_3779);
nor U3836 (N_3836,N_3683,N_3744);
nor U3837 (N_3837,N_3715,N_3647);
and U3838 (N_3838,N_3608,N_3689);
nor U3839 (N_3839,N_3684,N_3638);
nor U3840 (N_3840,N_3690,N_3677);
nor U3841 (N_3841,N_3733,N_3626);
and U3842 (N_3842,N_3708,N_3679);
and U3843 (N_3843,N_3659,N_3766);
and U3844 (N_3844,N_3746,N_3667);
nor U3845 (N_3845,N_3748,N_3767);
nand U3846 (N_3846,N_3701,N_3728);
xnor U3847 (N_3847,N_3685,N_3604);
nand U3848 (N_3848,N_3603,N_3761);
and U3849 (N_3849,N_3775,N_3751);
and U3850 (N_3850,N_3752,N_3661);
nor U3851 (N_3851,N_3777,N_3743);
xnor U3852 (N_3852,N_3765,N_3764);
nand U3853 (N_3853,N_3617,N_3710);
nand U3854 (N_3854,N_3693,N_3623);
nor U3855 (N_3855,N_3783,N_3662);
nand U3856 (N_3856,N_3649,N_3739);
and U3857 (N_3857,N_3611,N_3671);
or U3858 (N_3858,N_3698,N_3736);
nand U3859 (N_3859,N_3725,N_3657);
nor U3860 (N_3860,N_3795,N_3640);
nand U3861 (N_3861,N_3754,N_3601);
nand U3862 (N_3862,N_3785,N_3607);
nor U3863 (N_3863,N_3742,N_3755);
or U3864 (N_3864,N_3703,N_3627);
and U3865 (N_3865,N_3707,N_3613);
nor U3866 (N_3866,N_3651,N_3702);
nor U3867 (N_3867,N_3782,N_3758);
nand U3868 (N_3868,N_3609,N_3753);
nor U3869 (N_3869,N_3673,N_3784);
xor U3870 (N_3870,N_3768,N_3674);
nand U3871 (N_3871,N_3713,N_3716);
nand U3872 (N_3872,N_3630,N_3641);
nand U3873 (N_3873,N_3747,N_3771);
nor U3874 (N_3874,N_3711,N_3718);
or U3875 (N_3875,N_3705,N_3680);
or U3876 (N_3876,N_3759,N_3634);
nor U3877 (N_3877,N_3645,N_3670);
nand U3878 (N_3878,N_3750,N_3600);
or U3879 (N_3879,N_3639,N_3772);
or U3880 (N_3880,N_3688,N_3697);
nor U3881 (N_3881,N_3712,N_3709);
nor U3882 (N_3882,N_3749,N_3723);
nand U3883 (N_3883,N_3692,N_3632);
nand U3884 (N_3884,N_3687,N_3763);
xor U3885 (N_3885,N_3686,N_3653);
and U3886 (N_3886,N_3631,N_3741);
and U3887 (N_3887,N_3796,N_3681);
or U3888 (N_3888,N_3648,N_3769);
nor U3889 (N_3889,N_3615,N_3624);
xnor U3890 (N_3890,N_3699,N_3737);
and U3891 (N_3891,N_3762,N_3794);
or U3892 (N_3892,N_3798,N_3719);
nor U3893 (N_3893,N_3770,N_3676);
nand U3894 (N_3894,N_3730,N_3668);
nor U3895 (N_3895,N_3655,N_3720);
and U3896 (N_3896,N_3629,N_3666);
nor U3897 (N_3897,N_3646,N_3797);
and U3898 (N_3898,N_3717,N_3694);
nand U3899 (N_3899,N_3663,N_3665);
or U3900 (N_3900,N_3611,N_3772);
nand U3901 (N_3901,N_3793,N_3736);
and U3902 (N_3902,N_3698,N_3727);
or U3903 (N_3903,N_3778,N_3674);
nand U3904 (N_3904,N_3750,N_3728);
nor U3905 (N_3905,N_3619,N_3642);
and U3906 (N_3906,N_3628,N_3739);
nand U3907 (N_3907,N_3709,N_3746);
nand U3908 (N_3908,N_3764,N_3741);
or U3909 (N_3909,N_3657,N_3681);
and U3910 (N_3910,N_3714,N_3735);
nand U3911 (N_3911,N_3759,N_3753);
and U3912 (N_3912,N_3737,N_3608);
or U3913 (N_3913,N_3762,N_3738);
or U3914 (N_3914,N_3696,N_3644);
xor U3915 (N_3915,N_3621,N_3733);
nor U3916 (N_3916,N_3786,N_3782);
nand U3917 (N_3917,N_3709,N_3725);
or U3918 (N_3918,N_3773,N_3796);
nor U3919 (N_3919,N_3614,N_3639);
nand U3920 (N_3920,N_3694,N_3646);
or U3921 (N_3921,N_3689,N_3616);
and U3922 (N_3922,N_3734,N_3659);
and U3923 (N_3923,N_3783,N_3796);
and U3924 (N_3924,N_3626,N_3797);
nor U3925 (N_3925,N_3690,N_3715);
and U3926 (N_3926,N_3702,N_3645);
and U3927 (N_3927,N_3630,N_3778);
nand U3928 (N_3928,N_3738,N_3633);
nor U3929 (N_3929,N_3712,N_3667);
nor U3930 (N_3930,N_3657,N_3757);
nand U3931 (N_3931,N_3724,N_3671);
and U3932 (N_3932,N_3698,N_3787);
and U3933 (N_3933,N_3729,N_3612);
and U3934 (N_3934,N_3617,N_3752);
or U3935 (N_3935,N_3603,N_3635);
or U3936 (N_3936,N_3639,N_3703);
nor U3937 (N_3937,N_3711,N_3726);
nor U3938 (N_3938,N_3620,N_3727);
xor U3939 (N_3939,N_3606,N_3749);
or U3940 (N_3940,N_3629,N_3779);
nand U3941 (N_3941,N_3791,N_3633);
xor U3942 (N_3942,N_3797,N_3609);
nor U3943 (N_3943,N_3791,N_3759);
nand U3944 (N_3944,N_3668,N_3714);
nor U3945 (N_3945,N_3708,N_3750);
and U3946 (N_3946,N_3782,N_3777);
nand U3947 (N_3947,N_3783,N_3750);
or U3948 (N_3948,N_3680,N_3778);
nand U3949 (N_3949,N_3707,N_3752);
and U3950 (N_3950,N_3614,N_3616);
and U3951 (N_3951,N_3761,N_3765);
nand U3952 (N_3952,N_3793,N_3795);
and U3953 (N_3953,N_3605,N_3648);
xor U3954 (N_3954,N_3770,N_3639);
or U3955 (N_3955,N_3666,N_3692);
nor U3956 (N_3956,N_3645,N_3772);
or U3957 (N_3957,N_3737,N_3739);
or U3958 (N_3958,N_3735,N_3622);
and U3959 (N_3959,N_3640,N_3735);
nor U3960 (N_3960,N_3684,N_3650);
nor U3961 (N_3961,N_3787,N_3703);
nor U3962 (N_3962,N_3674,N_3770);
or U3963 (N_3963,N_3624,N_3742);
nand U3964 (N_3964,N_3713,N_3664);
or U3965 (N_3965,N_3683,N_3643);
xor U3966 (N_3966,N_3724,N_3631);
and U3967 (N_3967,N_3702,N_3606);
nor U3968 (N_3968,N_3707,N_3690);
nand U3969 (N_3969,N_3745,N_3714);
nand U3970 (N_3970,N_3634,N_3663);
nand U3971 (N_3971,N_3600,N_3604);
and U3972 (N_3972,N_3745,N_3628);
nor U3973 (N_3973,N_3670,N_3625);
and U3974 (N_3974,N_3620,N_3634);
and U3975 (N_3975,N_3749,N_3733);
nand U3976 (N_3976,N_3733,N_3771);
and U3977 (N_3977,N_3702,N_3692);
and U3978 (N_3978,N_3639,N_3673);
and U3979 (N_3979,N_3709,N_3710);
nor U3980 (N_3980,N_3782,N_3719);
or U3981 (N_3981,N_3694,N_3743);
or U3982 (N_3982,N_3718,N_3688);
nor U3983 (N_3983,N_3693,N_3741);
nand U3984 (N_3984,N_3688,N_3652);
nor U3985 (N_3985,N_3666,N_3764);
nand U3986 (N_3986,N_3616,N_3733);
nand U3987 (N_3987,N_3706,N_3653);
nor U3988 (N_3988,N_3704,N_3623);
and U3989 (N_3989,N_3628,N_3635);
or U3990 (N_3990,N_3688,N_3682);
and U3991 (N_3991,N_3705,N_3752);
or U3992 (N_3992,N_3624,N_3678);
or U3993 (N_3993,N_3794,N_3752);
and U3994 (N_3994,N_3686,N_3789);
or U3995 (N_3995,N_3619,N_3775);
nor U3996 (N_3996,N_3653,N_3737);
or U3997 (N_3997,N_3764,N_3646);
nand U3998 (N_3998,N_3677,N_3691);
or U3999 (N_3999,N_3689,N_3736);
and U4000 (N_4000,N_3940,N_3826);
or U4001 (N_4001,N_3889,N_3811);
nor U4002 (N_4002,N_3829,N_3843);
nand U4003 (N_4003,N_3855,N_3924);
or U4004 (N_4004,N_3925,N_3866);
nor U4005 (N_4005,N_3819,N_3905);
nand U4006 (N_4006,N_3931,N_3974);
or U4007 (N_4007,N_3941,N_3833);
or U4008 (N_4008,N_3993,N_3888);
and U4009 (N_4009,N_3876,N_3805);
or U4010 (N_4010,N_3995,N_3842);
and U4011 (N_4011,N_3887,N_3918);
or U4012 (N_4012,N_3987,N_3903);
and U4013 (N_4013,N_3927,N_3992);
or U4014 (N_4014,N_3875,N_3822);
nand U4015 (N_4015,N_3912,N_3898);
or U4016 (N_4016,N_3914,N_3864);
nor U4017 (N_4017,N_3951,N_3823);
nor U4018 (N_4018,N_3943,N_3944);
and U4019 (N_4019,N_3856,N_3921);
nand U4020 (N_4020,N_3910,N_3849);
or U4021 (N_4021,N_3945,N_3970);
nand U4022 (N_4022,N_3880,N_3817);
nor U4023 (N_4023,N_3844,N_3813);
nor U4024 (N_4024,N_3956,N_3892);
nor U4025 (N_4025,N_3872,N_3854);
nand U4026 (N_4026,N_3942,N_3932);
nor U4027 (N_4027,N_3969,N_3908);
and U4028 (N_4028,N_3965,N_3865);
nor U4029 (N_4029,N_3859,N_3824);
and U4030 (N_4030,N_3895,N_3950);
nor U4031 (N_4031,N_3988,N_3953);
or U4032 (N_4032,N_3860,N_3897);
nand U4033 (N_4033,N_3922,N_3919);
nand U4034 (N_4034,N_3847,N_3907);
nand U4035 (N_4035,N_3996,N_3963);
or U4036 (N_4036,N_3935,N_3947);
and U4037 (N_4037,N_3915,N_3899);
and U4038 (N_4038,N_3853,N_3836);
xnor U4039 (N_4039,N_3870,N_3939);
xnor U4040 (N_4040,N_3948,N_3830);
nand U4041 (N_4041,N_3896,N_3851);
or U4042 (N_4042,N_3858,N_3985);
nand U4043 (N_4043,N_3968,N_3983);
and U4044 (N_4044,N_3928,N_3874);
or U4045 (N_4045,N_3909,N_3937);
nor U4046 (N_4046,N_3920,N_3952);
nor U4047 (N_4047,N_3804,N_3801);
or U4048 (N_4048,N_3820,N_3906);
xnor U4049 (N_4049,N_3877,N_3846);
or U4050 (N_4050,N_3902,N_3807);
nand U4051 (N_4051,N_3867,N_3900);
nor U4052 (N_4052,N_3984,N_3971);
nand U4053 (N_4053,N_3871,N_3998);
nand U4054 (N_4054,N_3954,N_3913);
nor U4055 (N_4055,N_3882,N_3839);
nor U4056 (N_4056,N_3989,N_3962);
nor U4057 (N_4057,N_3868,N_3977);
nor U4058 (N_4058,N_3972,N_3917);
nor U4059 (N_4059,N_3904,N_3981);
nand U4060 (N_4060,N_3982,N_3929);
or U4061 (N_4061,N_3828,N_3891);
and U4062 (N_4062,N_3934,N_3840);
and U4063 (N_4063,N_3806,N_3815);
or U4064 (N_4064,N_3926,N_3886);
nand U4065 (N_4065,N_3994,N_3957);
or U4066 (N_4066,N_3831,N_3814);
or U4067 (N_4067,N_3808,N_3979);
nand U4068 (N_4068,N_3838,N_3938);
and U4069 (N_4069,N_3997,N_3841);
nor U4070 (N_4070,N_3894,N_3873);
nor U4071 (N_4071,N_3818,N_3936);
or U4072 (N_4072,N_3863,N_3810);
nand U4073 (N_4073,N_3857,N_3881);
nand U4074 (N_4074,N_3973,N_3800);
nor U4075 (N_4075,N_3893,N_3827);
nand U4076 (N_4076,N_3834,N_3835);
xnor U4077 (N_4077,N_3802,N_3869);
nor U4078 (N_4078,N_3809,N_3991);
and U4079 (N_4079,N_3883,N_3911);
nor U4080 (N_4080,N_3878,N_3879);
and U4081 (N_4081,N_3933,N_3852);
and U4082 (N_4082,N_3850,N_3976);
or U4083 (N_4083,N_3848,N_3955);
or U4084 (N_4084,N_3990,N_3890);
nand U4085 (N_4085,N_3978,N_3986);
or U4086 (N_4086,N_3949,N_3967);
or U4087 (N_4087,N_3980,N_3958);
and U4088 (N_4088,N_3825,N_3930);
and U4089 (N_4089,N_3960,N_3862);
and U4090 (N_4090,N_3946,N_3999);
nor U4091 (N_4091,N_3975,N_3845);
and U4092 (N_4092,N_3832,N_3837);
and U4093 (N_4093,N_3812,N_3959);
nor U4094 (N_4094,N_3861,N_3803);
nor U4095 (N_4095,N_3816,N_3961);
nor U4096 (N_4096,N_3901,N_3964);
nand U4097 (N_4097,N_3923,N_3966);
nand U4098 (N_4098,N_3885,N_3821);
nand U4099 (N_4099,N_3884,N_3916);
and U4100 (N_4100,N_3975,N_3952);
nor U4101 (N_4101,N_3855,N_3948);
nor U4102 (N_4102,N_3991,N_3837);
and U4103 (N_4103,N_3973,N_3902);
xor U4104 (N_4104,N_3931,N_3926);
nand U4105 (N_4105,N_3921,N_3909);
and U4106 (N_4106,N_3832,N_3863);
nor U4107 (N_4107,N_3971,N_3844);
nand U4108 (N_4108,N_3897,N_3979);
and U4109 (N_4109,N_3982,N_3864);
and U4110 (N_4110,N_3841,N_3821);
and U4111 (N_4111,N_3865,N_3832);
and U4112 (N_4112,N_3800,N_3886);
xor U4113 (N_4113,N_3968,N_3970);
or U4114 (N_4114,N_3980,N_3925);
xor U4115 (N_4115,N_3961,N_3943);
nor U4116 (N_4116,N_3988,N_3840);
nand U4117 (N_4117,N_3902,N_3903);
or U4118 (N_4118,N_3911,N_3810);
nand U4119 (N_4119,N_3888,N_3933);
nand U4120 (N_4120,N_3953,N_3945);
nor U4121 (N_4121,N_3805,N_3949);
nand U4122 (N_4122,N_3981,N_3954);
or U4123 (N_4123,N_3972,N_3855);
nand U4124 (N_4124,N_3991,N_3956);
or U4125 (N_4125,N_3979,N_3815);
nor U4126 (N_4126,N_3995,N_3860);
or U4127 (N_4127,N_3957,N_3818);
nor U4128 (N_4128,N_3851,N_3978);
nor U4129 (N_4129,N_3880,N_3928);
nor U4130 (N_4130,N_3927,N_3924);
and U4131 (N_4131,N_3945,N_3983);
or U4132 (N_4132,N_3853,N_3882);
and U4133 (N_4133,N_3963,N_3910);
nor U4134 (N_4134,N_3855,N_3863);
nor U4135 (N_4135,N_3991,N_3817);
nor U4136 (N_4136,N_3986,N_3871);
nor U4137 (N_4137,N_3989,N_3815);
nand U4138 (N_4138,N_3813,N_3819);
nor U4139 (N_4139,N_3839,N_3909);
nor U4140 (N_4140,N_3902,N_3974);
or U4141 (N_4141,N_3929,N_3843);
nand U4142 (N_4142,N_3852,N_3859);
or U4143 (N_4143,N_3837,N_3927);
nor U4144 (N_4144,N_3815,N_3960);
or U4145 (N_4145,N_3857,N_3912);
nand U4146 (N_4146,N_3896,N_3903);
nand U4147 (N_4147,N_3949,N_3828);
or U4148 (N_4148,N_3924,N_3823);
or U4149 (N_4149,N_3852,N_3977);
or U4150 (N_4150,N_3943,N_3903);
nor U4151 (N_4151,N_3982,N_3893);
nor U4152 (N_4152,N_3971,N_3998);
and U4153 (N_4153,N_3921,N_3811);
nand U4154 (N_4154,N_3828,N_3941);
nor U4155 (N_4155,N_3973,N_3896);
or U4156 (N_4156,N_3982,N_3855);
and U4157 (N_4157,N_3869,N_3811);
or U4158 (N_4158,N_3960,N_3851);
and U4159 (N_4159,N_3898,N_3925);
and U4160 (N_4160,N_3854,N_3879);
nand U4161 (N_4161,N_3999,N_3945);
or U4162 (N_4162,N_3889,N_3925);
or U4163 (N_4163,N_3829,N_3961);
or U4164 (N_4164,N_3973,N_3832);
nor U4165 (N_4165,N_3884,N_3922);
or U4166 (N_4166,N_3897,N_3971);
and U4167 (N_4167,N_3848,N_3853);
or U4168 (N_4168,N_3984,N_3860);
or U4169 (N_4169,N_3824,N_3928);
and U4170 (N_4170,N_3931,N_3849);
and U4171 (N_4171,N_3947,N_3999);
nor U4172 (N_4172,N_3926,N_3957);
nand U4173 (N_4173,N_3860,N_3867);
nand U4174 (N_4174,N_3987,N_3931);
nand U4175 (N_4175,N_3821,N_3819);
or U4176 (N_4176,N_3822,N_3907);
nor U4177 (N_4177,N_3846,N_3816);
or U4178 (N_4178,N_3896,N_3858);
and U4179 (N_4179,N_3875,N_3886);
and U4180 (N_4180,N_3875,N_3873);
and U4181 (N_4181,N_3948,N_3936);
and U4182 (N_4182,N_3951,N_3936);
and U4183 (N_4183,N_3839,N_3997);
nand U4184 (N_4184,N_3803,N_3996);
or U4185 (N_4185,N_3995,N_3887);
or U4186 (N_4186,N_3993,N_3937);
nand U4187 (N_4187,N_3846,N_3989);
or U4188 (N_4188,N_3881,N_3811);
nor U4189 (N_4189,N_3969,N_3982);
nor U4190 (N_4190,N_3898,N_3989);
nand U4191 (N_4191,N_3866,N_3800);
xor U4192 (N_4192,N_3881,N_3934);
and U4193 (N_4193,N_3803,N_3995);
xor U4194 (N_4194,N_3917,N_3907);
nand U4195 (N_4195,N_3814,N_3966);
or U4196 (N_4196,N_3832,N_3921);
nand U4197 (N_4197,N_3926,N_3941);
and U4198 (N_4198,N_3923,N_3917);
and U4199 (N_4199,N_3955,N_3842);
nor U4200 (N_4200,N_4071,N_4129);
nand U4201 (N_4201,N_4111,N_4118);
or U4202 (N_4202,N_4063,N_4130);
nor U4203 (N_4203,N_4089,N_4030);
nor U4204 (N_4204,N_4079,N_4047);
or U4205 (N_4205,N_4038,N_4134);
or U4206 (N_4206,N_4198,N_4023);
nand U4207 (N_4207,N_4153,N_4195);
nor U4208 (N_4208,N_4192,N_4150);
or U4209 (N_4209,N_4191,N_4138);
nand U4210 (N_4210,N_4035,N_4090);
or U4211 (N_4211,N_4028,N_4143);
nor U4212 (N_4212,N_4097,N_4092);
and U4213 (N_4213,N_4070,N_4175);
and U4214 (N_4214,N_4137,N_4127);
or U4215 (N_4215,N_4147,N_4187);
and U4216 (N_4216,N_4006,N_4178);
nor U4217 (N_4217,N_4121,N_4069);
nand U4218 (N_4218,N_4057,N_4123);
and U4219 (N_4219,N_4048,N_4081);
nand U4220 (N_4220,N_4019,N_4180);
or U4221 (N_4221,N_4155,N_4052);
nand U4222 (N_4222,N_4073,N_4076);
nand U4223 (N_4223,N_4128,N_4003);
nand U4224 (N_4224,N_4193,N_4190);
nand U4225 (N_4225,N_4002,N_4160);
and U4226 (N_4226,N_4102,N_4167);
nor U4227 (N_4227,N_4042,N_4086);
and U4228 (N_4228,N_4098,N_4120);
or U4229 (N_4229,N_4074,N_4106);
nand U4230 (N_4230,N_4169,N_4091);
or U4231 (N_4231,N_4114,N_4037);
and U4232 (N_4232,N_4109,N_4001);
nor U4233 (N_4233,N_4016,N_4154);
and U4234 (N_4234,N_4075,N_4027);
nand U4235 (N_4235,N_4033,N_4012);
nor U4236 (N_4236,N_4105,N_4124);
nand U4237 (N_4237,N_4148,N_4055);
nor U4238 (N_4238,N_4100,N_4049);
nand U4239 (N_4239,N_4108,N_4131);
nor U4240 (N_4240,N_4110,N_4010);
nand U4241 (N_4241,N_4043,N_4197);
and U4242 (N_4242,N_4007,N_4067);
nor U4243 (N_4243,N_4009,N_4044);
and U4244 (N_4244,N_4025,N_4041);
and U4245 (N_4245,N_4166,N_4117);
or U4246 (N_4246,N_4181,N_4112);
nand U4247 (N_4247,N_4161,N_4036);
nor U4248 (N_4248,N_4056,N_4176);
nand U4249 (N_4249,N_4095,N_4194);
nand U4250 (N_4250,N_4078,N_4144);
nand U4251 (N_4251,N_4093,N_4189);
xor U4252 (N_4252,N_4011,N_4045);
xor U4253 (N_4253,N_4141,N_4151);
nor U4254 (N_4254,N_4096,N_4013);
nor U4255 (N_4255,N_4179,N_4116);
or U4256 (N_4256,N_4185,N_4061);
nand U4257 (N_4257,N_4024,N_4159);
and U4258 (N_4258,N_4029,N_4196);
and U4259 (N_4259,N_4083,N_4170);
nand U4260 (N_4260,N_4177,N_4026);
nor U4261 (N_4261,N_4119,N_4152);
and U4262 (N_4262,N_4162,N_4107);
nand U4263 (N_4263,N_4164,N_4064);
nor U4264 (N_4264,N_4077,N_4031);
nor U4265 (N_4265,N_4183,N_4080);
or U4266 (N_4266,N_4173,N_4103);
xnor U4267 (N_4267,N_4054,N_4018);
nor U4268 (N_4268,N_4115,N_4085);
nand U4269 (N_4269,N_4140,N_4017);
xnor U4270 (N_4270,N_4146,N_4072);
and U4271 (N_4271,N_4199,N_4058);
and U4272 (N_4272,N_4039,N_4099);
or U4273 (N_4273,N_4186,N_4015);
or U4274 (N_4274,N_4184,N_4132);
nand U4275 (N_4275,N_4032,N_4004);
nand U4276 (N_4276,N_4021,N_4142);
nand U4277 (N_4277,N_4157,N_4022);
or U4278 (N_4278,N_4084,N_4158);
and U4279 (N_4279,N_4122,N_4133);
or U4280 (N_4280,N_4014,N_4126);
nor U4281 (N_4281,N_4062,N_4165);
nor U4282 (N_4282,N_4051,N_4034);
nor U4283 (N_4283,N_4008,N_4046);
or U4284 (N_4284,N_4101,N_4068);
xor U4285 (N_4285,N_4135,N_4059);
and U4286 (N_4286,N_4053,N_4145);
nand U4287 (N_4287,N_4113,N_4087);
and U4288 (N_4288,N_4000,N_4139);
or U4289 (N_4289,N_4104,N_4188);
and U4290 (N_4290,N_4082,N_4149);
or U4291 (N_4291,N_4040,N_4182);
and U4292 (N_4292,N_4172,N_4136);
nand U4293 (N_4293,N_4163,N_4088);
nor U4294 (N_4294,N_4168,N_4174);
and U4295 (N_4295,N_4171,N_4094);
or U4296 (N_4296,N_4060,N_4066);
and U4297 (N_4297,N_4020,N_4125);
nand U4298 (N_4298,N_4156,N_4050);
and U4299 (N_4299,N_4065,N_4005);
or U4300 (N_4300,N_4068,N_4088);
or U4301 (N_4301,N_4041,N_4177);
and U4302 (N_4302,N_4145,N_4080);
or U4303 (N_4303,N_4007,N_4010);
nand U4304 (N_4304,N_4121,N_4118);
and U4305 (N_4305,N_4071,N_4139);
nand U4306 (N_4306,N_4093,N_4104);
or U4307 (N_4307,N_4041,N_4119);
and U4308 (N_4308,N_4156,N_4018);
or U4309 (N_4309,N_4146,N_4170);
or U4310 (N_4310,N_4000,N_4071);
nor U4311 (N_4311,N_4166,N_4136);
nor U4312 (N_4312,N_4138,N_4061);
nor U4313 (N_4313,N_4073,N_4100);
and U4314 (N_4314,N_4053,N_4065);
and U4315 (N_4315,N_4110,N_4106);
xnor U4316 (N_4316,N_4179,N_4160);
nor U4317 (N_4317,N_4105,N_4195);
nor U4318 (N_4318,N_4076,N_4161);
nor U4319 (N_4319,N_4192,N_4084);
and U4320 (N_4320,N_4042,N_4149);
or U4321 (N_4321,N_4007,N_4197);
nor U4322 (N_4322,N_4056,N_4025);
nor U4323 (N_4323,N_4068,N_4057);
or U4324 (N_4324,N_4113,N_4099);
or U4325 (N_4325,N_4106,N_4012);
nand U4326 (N_4326,N_4004,N_4044);
nor U4327 (N_4327,N_4151,N_4008);
nor U4328 (N_4328,N_4154,N_4194);
nor U4329 (N_4329,N_4042,N_4060);
xnor U4330 (N_4330,N_4106,N_4100);
nand U4331 (N_4331,N_4067,N_4073);
nor U4332 (N_4332,N_4052,N_4028);
nor U4333 (N_4333,N_4045,N_4065);
and U4334 (N_4334,N_4003,N_4111);
nand U4335 (N_4335,N_4098,N_4012);
nor U4336 (N_4336,N_4054,N_4021);
or U4337 (N_4337,N_4138,N_4116);
nand U4338 (N_4338,N_4019,N_4062);
nor U4339 (N_4339,N_4160,N_4198);
or U4340 (N_4340,N_4053,N_4019);
or U4341 (N_4341,N_4055,N_4194);
or U4342 (N_4342,N_4151,N_4059);
nor U4343 (N_4343,N_4115,N_4190);
nor U4344 (N_4344,N_4045,N_4184);
nand U4345 (N_4345,N_4144,N_4009);
and U4346 (N_4346,N_4001,N_4159);
nor U4347 (N_4347,N_4054,N_4092);
nand U4348 (N_4348,N_4144,N_4179);
nand U4349 (N_4349,N_4122,N_4168);
or U4350 (N_4350,N_4123,N_4146);
or U4351 (N_4351,N_4017,N_4003);
or U4352 (N_4352,N_4141,N_4131);
nor U4353 (N_4353,N_4161,N_4176);
or U4354 (N_4354,N_4145,N_4092);
nor U4355 (N_4355,N_4014,N_4008);
and U4356 (N_4356,N_4177,N_4133);
and U4357 (N_4357,N_4125,N_4120);
nand U4358 (N_4358,N_4180,N_4058);
nand U4359 (N_4359,N_4146,N_4055);
nand U4360 (N_4360,N_4169,N_4038);
nand U4361 (N_4361,N_4148,N_4105);
and U4362 (N_4362,N_4139,N_4028);
and U4363 (N_4363,N_4000,N_4181);
nand U4364 (N_4364,N_4099,N_4035);
nand U4365 (N_4365,N_4190,N_4078);
or U4366 (N_4366,N_4197,N_4115);
xnor U4367 (N_4367,N_4059,N_4183);
nor U4368 (N_4368,N_4175,N_4099);
nand U4369 (N_4369,N_4113,N_4126);
and U4370 (N_4370,N_4044,N_4020);
nor U4371 (N_4371,N_4099,N_4146);
nand U4372 (N_4372,N_4140,N_4170);
nor U4373 (N_4373,N_4146,N_4063);
and U4374 (N_4374,N_4140,N_4156);
and U4375 (N_4375,N_4077,N_4185);
xor U4376 (N_4376,N_4158,N_4017);
or U4377 (N_4377,N_4085,N_4187);
or U4378 (N_4378,N_4177,N_4008);
or U4379 (N_4379,N_4103,N_4048);
nand U4380 (N_4380,N_4170,N_4073);
and U4381 (N_4381,N_4189,N_4080);
nor U4382 (N_4382,N_4120,N_4131);
or U4383 (N_4383,N_4123,N_4154);
or U4384 (N_4384,N_4130,N_4099);
nor U4385 (N_4385,N_4046,N_4082);
or U4386 (N_4386,N_4199,N_4143);
or U4387 (N_4387,N_4105,N_4035);
and U4388 (N_4388,N_4036,N_4014);
nand U4389 (N_4389,N_4045,N_4198);
or U4390 (N_4390,N_4044,N_4158);
and U4391 (N_4391,N_4179,N_4159);
or U4392 (N_4392,N_4076,N_4196);
nor U4393 (N_4393,N_4175,N_4075);
nor U4394 (N_4394,N_4104,N_4028);
nand U4395 (N_4395,N_4074,N_4116);
or U4396 (N_4396,N_4190,N_4004);
nor U4397 (N_4397,N_4029,N_4096);
nand U4398 (N_4398,N_4078,N_4044);
nand U4399 (N_4399,N_4093,N_4162);
nand U4400 (N_4400,N_4378,N_4227);
and U4401 (N_4401,N_4360,N_4332);
and U4402 (N_4402,N_4330,N_4287);
or U4403 (N_4403,N_4363,N_4214);
or U4404 (N_4404,N_4293,N_4318);
and U4405 (N_4405,N_4376,N_4337);
xor U4406 (N_4406,N_4362,N_4246);
or U4407 (N_4407,N_4372,N_4326);
and U4408 (N_4408,N_4264,N_4260);
and U4409 (N_4409,N_4284,N_4240);
nand U4410 (N_4410,N_4224,N_4300);
and U4411 (N_4411,N_4285,N_4253);
and U4412 (N_4412,N_4309,N_4218);
nand U4413 (N_4413,N_4223,N_4368);
and U4414 (N_4414,N_4395,N_4250);
and U4415 (N_4415,N_4234,N_4207);
or U4416 (N_4416,N_4328,N_4365);
and U4417 (N_4417,N_4296,N_4236);
and U4418 (N_4418,N_4259,N_4382);
and U4419 (N_4419,N_4277,N_4267);
and U4420 (N_4420,N_4205,N_4222);
or U4421 (N_4421,N_4203,N_4262);
or U4422 (N_4422,N_4320,N_4212);
nand U4423 (N_4423,N_4298,N_4294);
nand U4424 (N_4424,N_4334,N_4299);
nor U4425 (N_4425,N_4393,N_4225);
nor U4426 (N_4426,N_4273,N_4398);
xor U4427 (N_4427,N_4341,N_4353);
or U4428 (N_4428,N_4208,N_4317);
or U4429 (N_4429,N_4321,N_4306);
nor U4430 (N_4430,N_4319,N_4391);
nor U4431 (N_4431,N_4270,N_4333);
or U4432 (N_4432,N_4279,N_4385);
nand U4433 (N_4433,N_4244,N_4297);
nand U4434 (N_4434,N_4338,N_4359);
nor U4435 (N_4435,N_4219,N_4308);
nor U4436 (N_4436,N_4350,N_4217);
nor U4437 (N_4437,N_4375,N_4263);
xor U4438 (N_4438,N_4245,N_4381);
nand U4439 (N_4439,N_4291,N_4276);
or U4440 (N_4440,N_4388,N_4315);
nor U4441 (N_4441,N_4280,N_4386);
or U4442 (N_4442,N_4367,N_4323);
or U4443 (N_4443,N_4229,N_4283);
and U4444 (N_4444,N_4202,N_4380);
nand U4445 (N_4445,N_4210,N_4241);
nor U4446 (N_4446,N_4220,N_4397);
and U4447 (N_4447,N_4226,N_4364);
nor U4448 (N_4448,N_4331,N_4288);
nand U4449 (N_4449,N_4206,N_4373);
nor U4450 (N_4450,N_4383,N_4374);
nor U4451 (N_4451,N_4344,N_4261);
nand U4452 (N_4452,N_4265,N_4235);
or U4453 (N_4453,N_4242,N_4336);
nor U4454 (N_4454,N_4237,N_4357);
nor U4455 (N_4455,N_4390,N_4272);
and U4456 (N_4456,N_4213,N_4351);
and U4457 (N_4457,N_4313,N_4312);
nor U4458 (N_4458,N_4399,N_4215);
or U4459 (N_4459,N_4369,N_4271);
nand U4460 (N_4460,N_4329,N_4371);
and U4461 (N_4461,N_4352,N_4275);
and U4462 (N_4462,N_4282,N_4304);
and U4463 (N_4463,N_4396,N_4233);
or U4464 (N_4464,N_4258,N_4325);
or U4465 (N_4465,N_4370,N_4266);
nand U4466 (N_4466,N_4340,N_4286);
or U4467 (N_4467,N_4204,N_4232);
and U4468 (N_4468,N_4200,N_4354);
nand U4469 (N_4469,N_4379,N_4384);
nand U4470 (N_4470,N_4252,N_4268);
and U4471 (N_4471,N_4349,N_4255);
or U4472 (N_4472,N_4389,N_4238);
nor U4473 (N_4473,N_4366,N_4256);
nand U4474 (N_4474,N_4301,N_4355);
or U4475 (N_4475,N_4348,N_4231);
and U4476 (N_4476,N_4269,N_4251);
nand U4477 (N_4477,N_4247,N_4322);
nand U4478 (N_4478,N_4307,N_4316);
or U4479 (N_4479,N_4394,N_4311);
nand U4480 (N_4480,N_4239,N_4305);
xor U4481 (N_4481,N_4335,N_4295);
nor U4482 (N_4482,N_4361,N_4281);
and U4483 (N_4483,N_4302,N_4201);
nand U4484 (N_4484,N_4377,N_4358);
and U4485 (N_4485,N_4254,N_4257);
and U4486 (N_4486,N_4278,N_4327);
nor U4487 (N_4487,N_4324,N_4387);
nand U4488 (N_4488,N_4345,N_4230);
nor U4489 (N_4489,N_4228,N_4346);
and U4490 (N_4490,N_4347,N_4243);
and U4491 (N_4491,N_4310,N_4248);
and U4492 (N_4492,N_4290,N_4249);
nand U4493 (N_4493,N_4274,N_4342);
or U4494 (N_4494,N_4211,N_4303);
and U4495 (N_4495,N_4392,N_4216);
nand U4496 (N_4496,N_4292,N_4289);
or U4497 (N_4497,N_4356,N_4221);
or U4498 (N_4498,N_4339,N_4314);
or U4499 (N_4499,N_4209,N_4343);
nand U4500 (N_4500,N_4269,N_4304);
or U4501 (N_4501,N_4264,N_4223);
and U4502 (N_4502,N_4355,N_4366);
and U4503 (N_4503,N_4270,N_4339);
nor U4504 (N_4504,N_4399,N_4344);
and U4505 (N_4505,N_4288,N_4214);
and U4506 (N_4506,N_4267,N_4305);
or U4507 (N_4507,N_4210,N_4345);
or U4508 (N_4508,N_4289,N_4379);
and U4509 (N_4509,N_4273,N_4207);
and U4510 (N_4510,N_4336,N_4214);
nand U4511 (N_4511,N_4336,N_4253);
nand U4512 (N_4512,N_4240,N_4294);
nand U4513 (N_4513,N_4383,N_4275);
or U4514 (N_4514,N_4296,N_4394);
nand U4515 (N_4515,N_4290,N_4235);
or U4516 (N_4516,N_4203,N_4253);
nor U4517 (N_4517,N_4292,N_4359);
nor U4518 (N_4518,N_4312,N_4347);
xnor U4519 (N_4519,N_4230,N_4210);
nor U4520 (N_4520,N_4301,N_4365);
and U4521 (N_4521,N_4242,N_4250);
or U4522 (N_4522,N_4351,N_4241);
and U4523 (N_4523,N_4378,N_4237);
nor U4524 (N_4524,N_4344,N_4379);
and U4525 (N_4525,N_4284,N_4324);
and U4526 (N_4526,N_4270,N_4264);
nand U4527 (N_4527,N_4388,N_4345);
nor U4528 (N_4528,N_4334,N_4306);
or U4529 (N_4529,N_4375,N_4311);
nor U4530 (N_4530,N_4348,N_4219);
or U4531 (N_4531,N_4393,N_4313);
nand U4532 (N_4532,N_4306,N_4235);
or U4533 (N_4533,N_4388,N_4372);
and U4534 (N_4534,N_4299,N_4360);
xnor U4535 (N_4535,N_4237,N_4232);
or U4536 (N_4536,N_4282,N_4265);
nand U4537 (N_4537,N_4359,N_4243);
nor U4538 (N_4538,N_4342,N_4335);
or U4539 (N_4539,N_4333,N_4328);
or U4540 (N_4540,N_4275,N_4316);
and U4541 (N_4541,N_4385,N_4368);
or U4542 (N_4542,N_4362,N_4378);
nor U4543 (N_4543,N_4330,N_4373);
and U4544 (N_4544,N_4304,N_4362);
and U4545 (N_4545,N_4251,N_4210);
nor U4546 (N_4546,N_4336,N_4284);
or U4547 (N_4547,N_4328,N_4258);
and U4548 (N_4548,N_4287,N_4323);
nand U4549 (N_4549,N_4260,N_4334);
nand U4550 (N_4550,N_4320,N_4367);
nor U4551 (N_4551,N_4274,N_4356);
and U4552 (N_4552,N_4385,N_4200);
or U4553 (N_4553,N_4224,N_4327);
and U4554 (N_4554,N_4326,N_4201);
and U4555 (N_4555,N_4242,N_4218);
xnor U4556 (N_4556,N_4225,N_4295);
xnor U4557 (N_4557,N_4399,N_4338);
nor U4558 (N_4558,N_4236,N_4285);
nor U4559 (N_4559,N_4229,N_4212);
nor U4560 (N_4560,N_4241,N_4237);
or U4561 (N_4561,N_4327,N_4256);
and U4562 (N_4562,N_4242,N_4370);
and U4563 (N_4563,N_4397,N_4296);
and U4564 (N_4564,N_4313,N_4203);
and U4565 (N_4565,N_4223,N_4280);
nor U4566 (N_4566,N_4370,N_4372);
or U4567 (N_4567,N_4369,N_4381);
and U4568 (N_4568,N_4272,N_4393);
xor U4569 (N_4569,N_4238,N_4286);
nor U4570 (N_4570,N_4329,N_4246);
and U4571 (N_4571,N_4303,N_4314);
and U4572 (N_4572,N_4340,N_4225);
nor U4573 (N_4573,N_4326,N_4324);
nor U4574 (N_4574,N_4378,N_4348);
nor U4575 (N_4575,N_4207,N_4390);
and U4576 (N_4576,N_4380,N_4216);
nor U4577 (N_4577,N_4272,N_4327);
nor U4578 (N_4578,N_4319,N_4258);
nor U4579 (N_4579,N_4305,N_4339);
and U4580 (N_4580,N_4318,N_4303);
or U4581 (N_4581,N_4383,N_4203);
nor U4582 (N_4582,N_4267,N_4249);
or U4583 (N_4583,N_4296,N_4305);
and U4584 (N_4584,N_4326,N_4395);
nand U4585 (N_4585,N_4349,N_4280);
nor U4586 (N_4586,N_4337,N_4351);
nand U4587 (N_4587,N_4299,N_4394);
nor U4588 (N_4588,N_4299,N_4263);
or U4589 (N_4589,N_4378,N_4295);
nor U4590 (N_4590,N_4240,N_4351);
or U4591 (N_4591,N_4269,N_4279);
nor U4592 (N_4592,N_4376,N_4331);
nand U4593 (N_4593,N_4202,N_4266);
nor U4594 (N_4594,N_4287,N_4344);
xnor U4595 (N_4595,N_4355,N_4377);
nor U4596 (N_4596,N_4397,N_4265);
nor U4597 (N_4597,N_4241,N_4305);
nor U4598 (N_4598,N_4287,N_4364);
nor U4599 (N_4599,N_4256,N_4374);
and U4600 (N_4600,N_4402,N_4400);
nor U4601 (N_4601,N_4493,N_4463);
nand U4602 (N_4602,N_4404,N_4513);
nand U4603 (N_4603,N_4491,N_4512);
and U4604 (N_4604,N_4505,N_4470);
nor U4605 (N_4605,N_4432,N_4587);
nand U4606 (N_4606,N_4436,N_4516);
or U4607 (N_4607,N_4537,N_4549);
and U4608 (N_4608,N_4517,N_4554);
nor U4609 (N_4609,N_4419,N_4582);
or U4610 (N_4610,N_4462,N_4452);
or U4611 (N_4611,N_4577,N_4571);
nor U4612 (N_4612,N_4599,N_4465);
and U4613 (N_4613,N_4448,N_4523);
nor U4614 (N_4614,N_4471,N_4563);
and U4615 (N_4615,N_4475,N_4578);
or U4616 (N_4616,N_4502,N_4559);
and U4617 (N_4617,N_4459,N_4514);
and U4618 (N_4618,N_4440,N_4418);
or U4619 (N_4619,N_4497,N_4449);
and U4620 (N_4620,N_4406,N_4480);
nor U4621 (N_4621,N_4543,N_4446);
nand U4622 (N_4622,N_4501,N_4489);
nand U4623 (N_4623,N_4434,N_4539);
and U4624 (N_4624,N_4466,N_4585);
nor U4625 (N_4625,N_4534,N_4529);
nand U4626 (N_4626,N_4427,N_4525);
and U4627 (N_4627,N_4518,N_4458);
nor U4628 (N_4628,N_4415,N_4438);
or U4629 (N_4629,N_4424,N_4533);
and U4630 (N_4630,N_4545,N_4423);
and U4631 (N_4631,N_4408,N_4414);
nand U4632 (N_4632,N_4498,N_4556);
and U4633 (N_4633,N_4528,N_4433);
xor U4634 (N_4634,N_4588,N_4495);
and U4635 (N_4635,N_4494,N_4457);
nand U4636 (N_4636,N_4576,N_4580);
and U4637 (N_4637,N_4439,N_4488);
nand U4638 (N_4638,N_4544,N_4420);
nand U4639 (N_4639,N_4492,N_4565);
and U4640 (N_4640,N_4429,N_4486);
and U4641 (N_4641,N_4481,N_4431);
nor U4642 (N_4642,N_4574,N_4410);
nand U4643 (N_4643,N_4567,N_4451);
or U4644 (N_4644,N_4583,N_4435);
and U4645 (N_4645,N_4536,N_4592);
and U4646 (N_4646,N_4569,N_4511);
nand U4647 (N_4647,N_4417,N_4409);
nor U4648 (N_4648,N_4590,N_4566);
nand U4649 (N_4649,N_4535,N_4530);
or U4650 (N_4650,N_4548,N_4468);
and U4651 (N_4651,N_4560,N_4485);
and U4652 (N_4652,N_4586,N_4526);
or U4653 (N_4653,N_4447,N_4561);
or U4654 (N_4654,N_4461,N_4455);
and U4655 (N_4655,N_4496,N_4469);
nand U4656 (N_4656,N_4507,N_4521);
nor U4657 (N_4657,N_4482,N_4542);
or U4658 (N_4658,N_4437,N_4428);
or U4659 (N_4659,N_4568,N_4581);
nand U4660 (N_4660,N_4456,N_4503);
and U4661 (N_4661,N_4441,N_4520);
and U4662 (N_4662,N_4477,N_4522);
or U4663 (N_4663,N_4527,N_4555);
and U4664 (N_4664,N_4474,N_4584);
and U4665 (N_4665,N_4524,N_4553);
or U4666 (N_4666,N_4572,N_4579);
or U4667 (N_4667,N_4500,N_4573);
or U4668 (N_4668,N_4467,N_4484);
or U4669 (N_4669,N_4506,N_4464);
nand U4670 (N_4670,N_4479,N_4401);
or U4671 (N_4671,N_4531,N_4490);
and U4672 (N_4672,N_4421,N_4564);
and U4673 (N_4673,N_4422,N_4453);
and U4674 (N_4674,N_4546,N_4416);
or U4675 (N_4675,N_4595,N_4413);
nor U4676 (N_4676,N_4472,N_4443);
or U4677 (N_4677,N_4541,N_4483);
or U4678 (N_4678,N_4454,N_4450);
or U4679 (N_4679,N_4596,N_4473);
nand U4680 (N_4680,N_4547,N_4550);
or U4681 (N_4681,N_4412,N_4460);
or U4682 (N_4682,N_4407,N_4598);
and U4683 (N_4683,N_4504,N_4403);
nor U4684 (N_4684,N_4442,N_4570);
nor U4685 (N_4685,N_4510,N_4426);
nand U4686 (N_4686,N_4487,N_4476);
and U4687 (N_4687,N_4478,N_4508);
nor U4688 (N_4688,N_4597,N_4551);
nand U4689 (N_4689,N_4430,N_4515);
and U4690 (N_4690,N_4532,N_4562);
and U4691 (N_4691,N_4538,N_4557);
nand U4692 (N_4692,N_4499,N_4519);
nand U4693 (N_4693,N_4445,N_4575);
nor U4694 (N_4694,N_4509,N_4591);
nor U4695 (N_4695,N_4593,N_4425);
and U4696 (N_4696,N_4405,N_4589);
nor U4697 (N_4697,N_4594,N_4444);
or U4698 (N_4698,N_4552,N_4558);
and U4699 (N_4699,N_4540,N_4411);
nand U4700 (N_4700,N_4446,N_4535);
nor U4701 (N_4701,N_4592,N_4598);
or U4702 (N_4702,N_4431,N_4573);
nor U4703 (N_4703,N_4528,N_4472);
nand U4704 (N_4704,N_4499,N_4501);
nand U4705 (N_4705,N_4566,N_4470);
or U4706 (N_4706,N_4563,N_4441);
and U4707 (N_4707,N_4430,N_4414);
and U4708 (N_4708,N_4481,N_4526);
or U4709 (N_4709,N_4588,N_4485);
or U4710 (N_4710,N_4502,N_4458);
nand U4711 (N_4711,N_4417,N_4547);
nand U4712 (N_4712,N_4527,N_4519);
nor U4713 (N_4713,N_4552,N_4519);
nor U4714 (N_4714,N_4441,N_4506);
nand U4715 (N_4715,N_4504,N_4498);
nand U4716 (N_4716,N_4487,N_4488);
nand U4717 (N_4717,N_4473,N_4489);
or U4718 (N_4718,N_4536,N_4514);
nand U4719 (N_4719,N_4436,N_4550);
or U4720 (N_4720,N_4444,N_4423);
and U4721 (N_4721,N_4410,N_4559);
nand U4722 (N_4722,N_4533,N_4431);
nand U4723 (N_4723,N_4564,N_4581);
nor U4724 (N_4724,N_4424,N_4503);
or U4725 (N_4725,N_4594,N_4551);
or U4726 (N_4726,N_4435,N_4596);
and U4727 (N_4727,N_4404,N_4556);
and U4728 (N_4728,N_4444,N_4506);
nor U4729 (N_4729,N_4475,N_4415);
and U4730 (N_4730,N_4447,N_4529);
or U4731 (N_4731,N_4569,N_4514);
nand U4732 (N_4732,N_4587,N_4500);
nand U4733 (N_4733,N_4491,N_4511);
and U4734 (N_4734,N_4512,N_4585);
or U4735 (N_4735,N_4527,N_4461);
or U4736 (N_4736,N_4455,N_4578);
nand U4737 (N_4737,N_4573,N_4583);
nor U4738 (N_4738,N_4544,N_4490);
nand U4739 (N_4739,N_4533,N_4593);
and U4740 (N_4740,N_4589,N_4599);
nand U4741 (N_4741,N_4511,N_4545);
and U4742 (N_4742,N_4556,N_4551);
and U4743 (N_4743,N_4598,N_4416);
and U4744 (N_4744,N_4425,N_4478);
nand U4745 (N_4745,N_4496,N_4486);
nor U4746 (N_4746,N_4439,N_4524);
nand U4747 (N_4747,N_4400,N_4511);
or U4748 (N_4748,N_4425,N_4421);
or U4749 (N_4749,N_4544,N_4448);
or U4750 (N_4750,N_4488,N_4442);
and U4751 (N_4751,N_4506,N_4453);
or U4752 (N_4752,N_4561,N_4415);
nand U4753 (N_4753,N_4474,N_4433);
or U4754 (N_4754,N_4486,N_4487);
nor U4755 (N_4755,N_4574,N_4502);
and U4756 (N_4756,N_4405,N_4552);
nand U4757 (N_4757,N_4512,N_4575);
nor U4758 (N_4758,N_4420,N_4414);
xor U4759 (N_4759,N_4427,N_4559);
nand U4760 (N_4760,N_4503,N_4546);
or U4761 (N_4761,N_4433,N_4440);
and U4762 (N_4762,N_4568,N_4526);
and U4763 (N_4763,N_4467,N_4495);
and U4764 (N_4764,N_4569,N_4506);
nand U4765 (N_4765,N_4511,N_4563);
or U4766 (N_4766,N_4493,N_4429);
or U4767 (N_4767,N_4519,N_4560);
nor U4768 (N_4768,N_4425,N_4576);
xnor U4769 (N_4769,N_4526,N_4508);
nand U4770 (N_4770,N_4456,N_4530);
and U4771 (N_4771,N_4425,N_4442);
nor U4772 (N_4772,N_4593,N_4423);
nand U4773 (N_4773,N_4561,N_4414);
nor U4774 (N_4774,N_4413,N_4401);
or U4775 (N_4775,N_4567,N_4461);
nand U4776 (N_4776,N_4435,N_4592);
or U4777 (N_4777,N_4555,N_4409);
nand U4778 (N_4778,N_4454,N_4430);
nor U4779 (N_4779,N_4505,N_4543);
and U4780 (N_4780,N_4588,N_4451);
and U4781 (N_4781,N_4426,N_4415);
and U4782 (N_4782,N_4471,N_4413);
and U4783 (N_4783,N_4578,N_4562);
nor U4784 (N_4784,N_4591,N_4527);
nor U4785 (N_4785,N_4439,N_4519);
nand U4786 (N_4786,N_4551,N_4434);
xor U4787 (N_4787,N_4443,N_4580);
and U4788 (N_4788,N_4589,N_4539);
and U4789 (N_4789,N_4435,N_4526);
nor U4790 (N_4790,N_4531,N_4450);
nand U4791 (N_4791,N_4472,N_4440);
nor U4792 (N_4792,N_4549,N_4573);
or U4793 (N_4793,N_4543,N_4564);
nand U4794 (N_4794,N_4441,N_4587);
or U4795 (N_4795,N_4577,N_4472);
or U4796 (N_4796,N_4592,N_4422);
nor U4797 (N_4797,N_4581,N_4588);
or U4798 (N_4798,N_4552,N_4463);
nor U4799 (N_4799,N_4580,N_4571);
nand U4800 (N_4800,N_4620,N_4775);
or U4801 (N_4801,N_4708,N_4641);
nand U4802 (N_4802,N_4698,N_4729);
and U4803 (N_4803,N_4759,N_4762);
nand U4804 (N_4804,N_4716,N_4676);
nor U4805 (N_4805,N_4747,N_4619);
or U4806 (N_4806,N_4640,N_4794);
or U4807 (N_4807,N_4621,N_4723);
or U4808 (N_4808,N_4616,N_4774);
or U4809 (N_4809,N_4637,N_4769);
and U4810 (N_4810,N_4609,N_4665);
or U4811 (N_4811,N_4684,N_4766);
and U4812 (N_4812,N_4755,N_4672);
nand U4813 (N_4813,N_4670,N_4720);
or U4814 (N_4814,N_4781,N_4688);
or U4815 (N_4815,N_4668,N_4791);
and U4816 (N_4816,N_4651,N_4711);
nand U4817 (N_4817,N_4683,N_4702);
nor U4818 (N_4818,N_4602,N_4777);
and U4819 (N_4819,N_4606,N_4601);
nor U4820 (N_4820,N_4732,N_4611);
or U4821 (N_4821,N_4780,N_4615);
and U4822 (N_4822,N_4704,N_4669);
and U4823 (N_4823,N_4790,N_4715);
and U4824 (N_4824,N_4658,N_4632);
xnor U4825 (N_4825,N_4737,N_4771);
or U4826 (N_4826,N_4625,N_4663);
nand U4827 (N_4827,N_4795,N_4779);
and U4828 (N_4828,N_4763,N_4649);
nor U4829 (N_4829,N_4754,N_4783);
nor U4830 (N_4830,N_4660,N_4736);
nand U4831 (N_4831,N_4657,N_4682);
or U4832 (N_4832,N_4655,N_4607);
and U4833 (N_4833,N_4675,N_4624);
nor U4834 (N_4834,N_4696,N_4734);
nor U4835 (N_4835,N_4667,N_4659);
or U4836 (N_4836,N_4642,N_4765);
or U4837 (N_4837,N_4604,N_4745);
nand U4838 (N_4838,N_4697,N_4728);
or U4839 (N_4839,N_4768,N_4610);
and U4840 (N_4840,N_4756,N_4695);
nand U4841 (N_4841,N_4646,N_4612);
nand U4842 (N_4842,N_4626,N_4798);
nand U4843 (N_4843,N_4636,N_4664);
nor U4844 (N_4844,N_4710,N_4635);
nor U4845 (N_4845,N_4752,N_4654);
nor U4846 (N_4846,N_4713,N_4787);
and U4847 (N_4847,N_4694,N_4679);
nand U4848 (N_4848,N_4693,N_4797);
and U4849 (N_4849,N_4746,N_4700);
and U4850 (N_4850,N_4760,N_4623);
nand U4851 (N_4851,N_4703,N_4674);
nand U4852 (N_4852,N_4753,N_4719);
nor U4853 (N_4853,N_4796,N_4742);
nand U4854 (N_4854,N_4714,N_4722);
and U4855 (N_4855,N_4792,N_4613);
or U4856 (N_4856,N_4717,N_4749);
nor U4857 (N_4857,N_4788,N_4744);
or U4858 (N_4858,N_4724,N_4718);
and U4859 (N_4859,N_4699,N_4608);
nand U4860 (N_4860,N_4761,N_4644);
and U4861 (N_4861,N_4605,N_4782);
and U4862 (N_4862,N_4627,N_4633);
xnor U4863 (N_4863,N_4776,N_4631);
or U4864 (N_4864,N_4691,N_4689);
and U4865 (N_4865,N_4630,N_4673);
or U4866 (N_4866,N_4600,N_4740);
or U4867 (N_4867,N_4645,N_4687);
nor U4868 (N_4868,N_4733,N_4735);
or U4869 (N_4869,N_4638,N_4634);
nor U4870 (N_4870,N_4773,N_4731);
nor U4871 (N_4871,N_4793,N_4758);
xnor U4872 (N_4872,N_4772,N_4789);
or U4873 (N_4873,N_4725,N_4639);
nand U4874 (N_4874,N_4730,N_4629);
nor U4875 (N_4875,N_4757,N_4690);
or U4876 (N_4876,N_4726,N_4706);
or U4877 (N_4877,N_4786,N_4677);
nor U4878 (N_4878,N_4721,N_4705);
nand U4879 (N_4879,N_4686,N_4750);
or U4880 (N_4880,N_4628,N_4785);
and U4881 (N_4881,N_4709,N_4656);
and U4882 (N_4882,N_4618,N_4603);
and U4883 (N_4883,N_4681,N_4770);
and U4884 (N_4884,N_4678,N_4751);
and U4885 (N_4885,N_4764,N_4767);
nor U4886 (N_4886,N_4666,N_4648);
nor U4887 (N_4887,N_4653,N_4741);
nor U4888 (N_4888,N_4701,N_4739);
nor U4889 (N_4889,N_4685,N_4614);
or U4890 (N_4890,N_4799,N_4662);
or U4891 (N_4891,N_4661,N_4748);
and U4892 (N_4892,N_4692,N_4622);
nand U4893 (N_4893,N_4650,N_4671);
nor U4894 (N_4894,N_4652,N_4778);
nor U4895 (N_4895,N_4784,N_4647);
nand U4896 (N_4896,N_4738,N_4617);
nor U4897 (N_4897,N_4707,N_4727);
or U4898 (N_4898,N_4680,N_4743);
nor U4899 (N_4899,N_4712,N_4643);
nand U4900 (N_4900,N_4712,N_4785);
nand U4901 (N_4901,N_4734,N_4720);
nand U4902 (N_4902,N_4636,N_4637);
and U4903 (N_4903,N_4717,N_4647);
or U4904 (N_4904,N_4680,N_4705);
nor U4905 (N_4905,N_4779,N_4747);
nor U4906 (N_4906,N_4627,N_4720);
and U4907 (N_4907,N_4666,N_4698);
nor U4908 (N_4908,N_4798,N_4649);
xor U4909 (N_4909,N_4727,N_4611);
nor U4910 (N_4910,N_4672,N_4702);
or U4911 (N_4911,N_4658,N_4795);
and U4912 (N_4912,N_4791,N_4736);
nor U4913 (N_4913,N_4728,N_4735);
nand U4914 (N_4914,N_4722,N_4655);
nor U4915 (N_4915,N_4751,N_4736);
and U4916 (N_4916,N_4672,N_4798);
or U4917 (N_4917,N_4743,N_4616);
or U4918 (N_4918,N_4660,N_4798);
nor U4919 (N_4919,N_4673,N_4623);
nor U4920 (N_4920,N_4718,N_4747);
nand U4921 (N_4921,N_4611,N_4740);
nor U4922 (N_4922,N_4674,N_4777);
nor U4923 (N_4923,N_4605,N_4768);
nand U4924 (N_4924,N_4629,N_4699);
nand U4925 (N_4925,N_4628,N_4764);
nand U4926 (N_4926,N_4607,N_4721);
nand U4927 (N_4927,N_4655,N_4637);
and U4928 (N_4928,N_4669,N_4628);
and U4929 (N_4929,N_4683,N_4666);
nor U4930 (N_4930,N_4675,N_4681);
or U4931 (N_4931,N_4768,N_4744);
and U4932 (N_4932,N_4637,N_4700);
nor U4933 (N_4933,N_4642,N_4721);
nor U4934 (N_4934,N_4620,N_4603);
nand U4935 (N_4935,N_4676,N_4645);
nand U4936 (N_4936,N_4713,N_4760);
nand U4937 (N_4937,N_4762,N_4678);
nand U4938 (N_4938,N_4741,N_4730);
nand U4939 (N_4939,N_4724,N_4752);
or U4940 (N_4940,N_4683,N_4721);
or U4941 (N_4941,N_4728,N_4719);
nand U4942 (N_4942,N_4602,N_4717);
and U4943 (N_4943,N_4792,N_4662);
or U4944 (N_4944,N_4687,N_4719);
or U4945 (N_4945,N_4677,N_4643);
nand U4946 (N_4946,N_4736,N_4716);
or U4947 (N_4947,N_4723,N_4730);
or U4948 (N_4948,N_4794,N_4753);
nor U4949 (N_4949,N_4782,N_4710);
or U4950 (N_4950,N_4777,N_4756);
or U4951 (N_4951,N_4753,N_4774);
or U4952 (N_4952,N_4605,N_4794);
or U4953 (N_4953,N_4756,N_4758);
nor U4954 (N_4954,N_4623,N_4713);
nand U4955 (N_4955,N_4774,N_4724);
nor U4956 (N_4956,N_4700,N_4620);
or U4957 (N_4957,N_4728,N_4790);
and U4958 (N_4958,N_4613,N_4609);
and U4959 (N_4959,N_4765,N_4684);
xor U4960 (N_4960,N_4770,N_4682);
or U4961 (N_4961,N_4712,N_4792);
or U4962 (N_4962,N_4625,N_4767);
or U4963 (N_4963,N_4792,N_4683);
xor U4964 (N_4964,N_4626,N_4728);
or U4965 (N_4965,N_4662,N_4766);
nand U4966 (N_4966,N_4791,N_4684);
nor U4967 (N_4967,N_4762,N_4715);
nand U4968 (N_4968,N_4797,N_4777);
or U4969 (N_4969,N_4704,N_4686);
nand U4970 (N_4970,N_4733,N_4771);
nor U4971 (N_4971,N_4678,N_4698);
or U4972 (N_4972,N_4777,N_4682);
or U4973 (N_4973,N_4723,N_4764);
and U4974 (N_4974,N_4786,N_4788);
or U4975 (N_4975,N_4655,N_4715);
and U4976 (N_4976,N_4741,N_4689);
nand U4977 (N_4977,N_4787,N_4629);
or U4978 (N_4978,N_4779,N_4797);
nand U4979 (N_4979,N_4610,N_4736);
and U4980 (N_4980,N_4631,N_4735);
nor U4981 (N_4981,N_4700,N_4683);
nand U4982 (N_4982,N_4728,N_4723);
nor U4983 (N_4983,N_4717,N_4707);
nand U4984 (N_4984,N_4675,N_4767);
or U4985 (N_4985,N_4792,N_4720);
or U4986 (N_4986,N_4608,N_4636);
nor U4987 (N_4987,N_4798,N_4684);
and U4988 (N_4988,N_4778,N_4721);
and U4989 (N_4989,N_4670,N_4792);
nor U4990 (N_4990,N_4723,N_4666);
nand U4991 (N_4991,N_4776,N_4689);
and U4992 (N_4992,N_4754,N_4732);
nor U4993 (N_4993,N_4738,N_4616);
nor U4994 (N_4994,N_4700,N_4655);
or U4995 (N_4995,N_4778,N_4693);
or U4996 (N_4996,N_4717,N_4688);
or U4997 (N_4997,N_4742,N_4730);
and U4998 (N_4998,N_4771,N_4642);
or U4999 (N_4999,N_4706,N_4656);
nand U5000 (N_5000,N_4869,N_4862);
nand U5001 (N_5001,N_4943,N_4931);
xnor U5002 (N_5002,N_4861,N_4957);
nand U5003 (N_5003,N_4928,N_4836);
nand U5004 (N_5004,N_4956,N_4823);
nor U5005 (N_5005,N_4840,N_4803);
nand U5006 (N_5006,N_4872,N_4999);
nor U5007 (N_5007,N_4968,N_4980);
nand U5008 (N_5008,N_4981,N_4835);
xor U5009 (N_5009,N_4936,N_4822);
nor U5010 (N_5010,N_4874,N_4886);
nand U5011 (N_5011,N_4992,N_4850);
nand U5012 (N_5012,N_4844,N_4989);
nand U5013 (N_5013,N_4892,N_4826);
nor U5014 (N_5014,N_4800,N_4962);
nand U5015 (N_5015,N_4967,N_4893);
and U5016 (N_5016,N_4847,N_4876);
nor U5017 (N_5017,N_4903,N_4960);
and U5018 (N_5018,N_4924,N_4839);
nand U5019 (N_5019,N_4873,N_4906);
and U5020 (N_5020,N_4841,N_4814);
and U5021 (N_5021,N_4813,N_4922);
nand U5022 (N_5022,N_4934,N_4938);
nor U5023 (N_5023,N_4908,N_4883);
or U5024 (N_5024,N_4902,N_4988);
nand U5025 (N_5025,N_4818,N_4849);
nor U5026 (N_5026,N_4946,N_4911);
nor U5027 (N_5027,N_4901,N_4949);
or U5028 (N_5028,N_4819,N_4935);
and U5029 (N_5029,N_4890,N_4939);
or U5030 (N_5030,N_4945,N_4804);
nand U5031 (N_5031,N_4976,N_4858);
nand U5032 (N_5032,N_4987,N_4973);
or U5033 (N_5033,N_4947,N_4966);
nand U5034 (N_5034,N_4891,N_4910);
or U5035 (N_5035,N_4909,N_4871);
xor U5036 (N_5036,N_4926,N_4831);
nor U5037 (N_5037,N_4843,N_4953);
nand U5038 (N_5038,N_4888,N_4896);
or U5039 (N_5039,N_4940,N_4856);
nor U5040 (N_5040,N_4870,N_4829);
and U5041 (N_5041,N_4952,N_4864);
or U5042 (N_5042,N_4972,N_4961);
and U5043 (N_5043,N_4985,N_4964);
nand U5044 (N_5044,N_4994,N_4827);
and U5045 (N_5045,N_4885,N_4820);
nor U5046 (N_5046,N_4955,N_4833);
nand U5047 (N_5047,N_4837,N_4997);
and U5048 (N_5048,N_4852,N_4937);
or U5049 (N_5049,N_4895,N_4817);
and U5050 (N_5050,N_4950,N_4904);
nand U5051 (N_5051,N_4915,N_4854);
nor U5052 (N_5052,N_4907,N_4979);
and U5053 (N_5053,N_4948,N_4986);
and U5054 (N_5054,N_4842,N_4851);
nand U5055 (N_5055,N_4916,N_4942);
nor U5056 (N_5056,N_4917,N_4824);
and U5057 (N_5057,N_4923,N_4808);
and U5058 (N_5058,N_4900,N_4912);
or U5059 (N_5059,N_4930,N_4878);
nand U5060 (N_5060,N_4815,N_4963);
and U5061 (N_5061,N_4845,N_4919);
nand U5062 (N_5062,N_4801,N_4880);
or U5063 (N_5063,N_4970,N_4991);
xor U5064 (N_5064,N_4834,N_4863);
nor U5065 (N_5065,N_4913,N_4898);
and U5066 (N_5066,N_4995,N_4887);
nor U5067 (N_5067,N_4899,N_4846);
nor U5068 (N_5068,N_4965,N_4905);
nand U5069 (N_5069,N_4832,N_4889);
nor U5070 (N_5070,N_4812,N_4802);
and U5071 (N_5071,N_4810,N_4866);
nand U5072 (N_5072,N_4925,N_4816);
nor U5073 (N_5073,N_4867,N_4879);
nand U5074 (N_5074,N_4877,N_4932);
nor U5075 (N_5075,N_4933,N_4811);
nand U5076 (N_5076,N_4807,N_4881);
or U5077 (N_5077,N_4865,N_4982);
or U5078 (N_5078,N_4984,N_4920);
nand U5079 (N_5079,N_4859,N_4921);
or U5080 (N_5080,N_4828,N_4914);
and U5081 (N_5081,N_4830,N_4805);
xnor U5082 (N_5082,N_4868,N_4977);
nor U5083 (N_5083,N_4848,N_4806);
nand U5084 (N_5084,N_4929,N_4951);
nand U5085 (N_5085,N_4860,N_4959);
nor U5086 (N_5086,N_4884,N_4927);
or U5087 (N_5087,N_4918,N_4954);
or U5088 (N_5088,N_4882,N_4983);
nand U5089 (N_5089,N_4958,N_4974);
nand U5090 (N_5090,N_4998,N_4894);
or U5091 (N_5091,N_4825,N_4993);
nor U5092 (N_5092,N_4975,N_4838);
and U5093 (N_5093,N_4855,N_4821);
nor U5094 (N_5094,N_4944,N_4996);
or U5095 (N_5095,N_4941,N_4990);
nand U5096 (N_5096,N_4875,N_4857);
or U5097 (N_5097,N_4853,N_4809);
or U5098 (N_5098,N_4969,N_4897);
or U5099 (N_5099,N_4978,N_4971);
or U5100 (N_5100,N_4877,N_4960);
nand U5101 (N_5101,N_4897,N_4826);
nor U5102 (N_5102,N_4840,N_4957);
nand U5103 (N_5103,N_4868,N_4938);
and U5104 (N_5104,N_4979,N_4818);
nor U5105 (N_5105,N_4802,N_4835);
or U5106 (N_5106,N_4855,N_4922);
nor U5107 (N_5107,N_4935,N_4938);
or U5108 (N_5108,N_4994,N_4967);
nor U5109 (N_5109,N_4961,N_4850);
xor U5110 (N_5110,N_4843,N_4848);
nor U5111 (N_5111,N_4971,N_4910);
nor U5112 (N_5112,N_4926,N_4917);
or U5113 (N_5113,N_4973,N_4818);
nand U5114 (N_5114,N_4966,N_4995);
nor U5115 (N_5115,N_4989,N_4849);
and U5116 (N_5116,N_4956,N_4986);
or U5117 (N_5117,N_4913,N_4970);
or U5118 (N_5118,N_4931,N_4848);
and U5119 (N_5119,N_4935,N_4942);
xnor U5120 (N_5120,N_4866,N_4890);
or U5121 (N_5121,N_4905,N_4923);
nor U5122 (N_5122,N_4885,N_4845);
nand U5123 (N_5123,N_4926,N_4852);
nand U5124 (N_5124,N_4828,N_4845);
and U5125 (N_5125,N_4948,N_4969);
and U5126 (N_5126,N_4828,N_4818);
nand U5127 (N_5127,N_4809,N_4879);
and U5128 (N_5128,N_4913,N_4955);
nand U5129 (N_5129,N_4998,N_4810);
nor U5130 (N_5130,N_4851,N_4947);
nand U5131 (N_5131,N_4953,N_4976);
nor U5132 (N_5132,N_4947,N_4883);
nand U5133 (N_5133,N_4839,N_4826);
nand U5134 (N_5134,N_4872,N_4916);
and U5135 (N_5135,N_4991,N_4833);
and U5136 (N_5136,N_4855,N_4904);
or U5137 (N_5137,N_4918,N_4906);
or U5138 (N_5138,N_4941,N_4927);
nand U5139 (N_5139,N_4975,N_4929);
or U5140 (N_5140,N_4994,N_4909);
nand U5141 (N_5141,N_4845,N_4869);
or U5142 (N_5142,N_4944,N_4818);
nor U5143 (N_5143,N_4957,N_4863);
nor U5144 (N_5144,N_4852,N_4882);
xor U5145 (N_5145,N_4926,N_4964);
or U5146 (N_5146,N_4960,N_4926);
nand U5147 (N_5147,N_4985,N_4912);
nand U5148 (N_5148,N_4860,N_4884);
or U5149 (N_5149,N_4899,N_4971);
nand U5150 (N_5150,N_4912,N_4939);
and U5151 (N_5151,N_4911,N_4988);
and U5152 (N_5152,N_4892,N_4801);
nor U5153 (N_5153,N_4940,N_4986);
or U5154 (N_5154,N_4831,N_4955);
nand U5155 (N_5155,N_4806,N_4861);
xor U5156 (N_5156,N_4882,N_4884);
nor U5157 (N_5157,N_4807,N_4874);
nand U5158 (N_5158,N_4879,N_4949);
and U5159 (N_5159,N_4804,N_4843);
nand U5160 (N_5160,N_4992,N_4942);
nand U5161 (N_5161,N_4813,N_4803);
nand U5162 (N_5162,N_4968,N_4864);
or U5163 (N_5163,N_4899,N_4974);
and U5164 (N_5164,N_4939,N_4843);
nand U5165 (N_5165,N_4812,N_4846);
or U5166 (N_5166,N_4973,N_4962);
and U5167 (N_5167,N_4891,N_4949);
and U5168 (N_5168,N_4852,N_4821);
or U5169 (N_5169,N_4941,N_4805);
or U5170 (N_5170,N_4906,N_4907);
nand U5171 (N_5171,N_4890,N_4857);
or U5172 (N_5172,N_4834,N_4991);
or U5173 (N_5173,N_4881,N_4966);
nand U5174 (N_5174,N_4879,N_4853);
xnor U5175 (N_5175,N_4976,N_4979);
xnor U5176 (N_5176,N_4979,N_4986);
or U5177 (N_5177,N_4816,N_4943);
and U5178 (N_5178,N_4915,N_4816);
and U5179 (N_5179,N_4934,N_4806);
xor U5180 (N_5180,N_4952,N_4924);
or U5181 (N_5181,N_4876,N_4934);
and U5182 (N_5182,N_4886,N_4983);
and U5183 (N_5183,N_4803,N_4839);
nand U5184 (N_5184,N_4805,N_4837);
and U5185 (N_5185,N_4969,N_4901);
nand U5186 (N_5186,N_4910,N_4816);
and U5187 (N_5187,N_4841,N_4929);
nor U5188 (N_5188,N_4801,N_4804);
nor U5189 (N_5189,N_4889,N_4923);
or U5190 (N_5190,N_4980,N_4828);
and U5191 (N_5191,N_4981,N_4993);
nor U5192 (N_5192,N_4988,N_4925);
and U5193 (N_5193,N_4852,N_4940);
nand U5194 (N_5194,N_4944,N_4960);
or U5195 (N_5195,N_4871,N_4908);
nand U5196 (N_5196,N_4944,N_4901);
nand U5197 (N_5197,N_4998,N_4956);
nor U5198 (N_5198,N_4959,N_4807);
or U5199 (N_5199,N_4856,N_4835);
and U5200 (N_5200,N_5147,N_5144);
or U5201 (N_5201,N_5045,N_5158);
or U5202 (N_5202,N_5106,N_5102);
and U5203 (N_5203,N_5098,N_5035);
xnor U5204 (N_5204,N_5041,N_5151);
nand U5205 (N_5205,N_5128,N_5038);
nor U5206 (N_5206,N_5112,N_5056);
or U5207 (N_5207,N_5066,N_5085);
or U5208 (N_5208,N_5131,N_5141);
nand U5209 (N_5209,N_5100,N_5118);
or U5210 (N_5210,N_5074,N_5119);
or U5211 (N_5211,N_5108,N_5148);
or U5212 (N_5212,N_5026,N_5116);
nand U5213 (N_5213,N_5165,N_5010);
nor U5214 (N_5214,N_5019,N_5022);
and U5215 (N_5215,N_5189,N_5024);
nand U5216 (N_5216,N_5187,N_5132);
or U5217 (N_5217,N_5073,N_5050);
and U5218 (N_5218,N_5068,N_5043);
and U5219 (N_5219,N_5160,N_5006);
and U5220 (N_5220,N_5140,N_5058);
nand U5221 (N_5221,N_5153,N_5152);
or U5222 (N_5222,N_5081,N_5000);
and U5223 (N_5223,N_5007,N_5062);
and U5224 (N_5224,N_5099,N_5166);
and U5225 (N_5225,N_5054,N_5084);
nand U5226 (N_5226,N_5157,N_5192);
nand U5227 (N_5227,N_5018,N_5125);
or U5228 (N_5228,N_5037,N_5191);
or U5229 (N_5229,N_5103,N_5134);
nor U5230 (N_5230,N_5036,N_5053);
nand U5231 (N_5231,N_5154,N_5076);
and U5232 (N_5232,N_5156,N_5096);
xnor U5233 (N_5233,N_5002,N_5030);
nand U5234 (N_5234,N_5190,N_5193);
and U5235 (N_5235,N_5114,N_5090);
nor U5236 (N_5236,N_5111,N_5137);
or U5237 (N_5237,N_5175,N_5162);
nor U5238 (N_5238,N_5104,N_5195);
or U5239 (N_5239,N_5001,N_5070);
or U5240 (N_5240,N_5163,N_5133);
or U5241 (N_5241,N_5060,N_5149);
or U5242 (N_5242,N_5199,N_5013);
nand U5243 (N_5243,N_5105,N_5124);
and U5244 (N_5244,N_5186,N_5020);
nand U5245 (N_5245,N_5123,N_5177);
and U5246 (N_5246,N_5179,N_5176);
nor U5247 (N_5247,N_5184,N_5004);
nor U5248 (N_5248,N_5122,N_5092);
nand U5249 (N_5249,N_5078,N_5172);
nand U5250 (N_5250,N_5129,N_5047);
and U5251 (N_5251,N_5097,N_5029);
nand U5252 (N_5252,N_5017,N_5057);
and U5253 (N_5253,N_5159,N_5015);
or U5254 (N_5254,N_5178,N_5196);
or U5255 (N_5255,N_5059,N_5126);
and U5256 (N_5256,N_5061,N_5009);
or U5257 (N_5257,N_5113,N_5127);
xnor U5258 (N_5258,N_5197,N_5171);
and U5259 (N_5259,N_5049,N_5091);
nor U5260 (N_5260,N_5136,N_5048);
or U5261 (N_5261,N_5033,N_5005);
and U5262 (N_5262,N_5130,N_5032);
and U5263 (N_5263,N_5142,N_5077);
and U5264 (N_5264,N_5089,N_5031);
and U5265 (N_5265,N_5063,N_5003);
nor U5266 (N_5266,N_5071,N_5121);
nand U5267 (N_5267,N_5095,N_5042);
nor U5268 (N_5268,N_5083,N_5094);
nor U5269 (N_5269,N_5052,N_5025);
nor U5270 (N_5270,N_5067,N_5167);
nand U5271 (N_5271,N_5107,N_5109);
and U5272 (N_5272,N_5117,N_5170);
nand U5273 (N_5273,N_5155,N_5046);
nand U5274 (N_5274,N_5194,N_5027);
nand U5275 (N_5275,N_5145,N_5012);
nand U5276 (N_5276,N_5168,N_5034);
nor U5277 (N_5277,N_5138,N_5023);
or U5278 (N_5278,N_5088,N_5008);
and U5279 (N_5279,N_5174,N_5082);
or U5280 (N_5280,N_5169,N_5075);
or U5281 (N_5281,N_5173,N_5120);
nand U5282 (N_5282,N_5101,N_5146);
nand U5283 (N_5283,N_5021,N_5011);
or U5284 (N_5284,N_5115,N_5080);
nor U5285 (N_5285,N_5072,N_5143);
nand U5286 (N_5286,N_5093,N_5016);
or U5287 (N_5287,N_5028,N_5069);
nand U5288 (N_5288,N_5039,N_5181);
nand U5289 (N_5289,N_5086,N_5188);
xor U5290 (N_5290,N_5183,N_5185);
nor U5291 (N_5291,N_5161,N_5180);
or U5292 (N_5292,N_5079,N_5065);
and U5293 (N_5293,N_5164,N_5110);
or U5294 (N_5294,N_5014,N_5087);
or U5295 (N_5295,N_5064,N_5135);
nor U5296 (N_5296,N_5139,N_5150);
nor U5297 (N_5297,N_5040,N_5198);
or U5298 (N_5298,N_5182,N_5051);
nor U5299 (N_5299,N_5055,N_5044);
and U5300 (N_5300,N_5180,N_5162);
nand U5301 (N_5301,N_5142,N_5167);
or U5302 (N_5302,N_5101,N_5087);
or U5303 (N_5303,N_5152,N_5007);
nand U5304 (N_5304,N_5184,N_5089);
nor U5305 (N_5305,N_5134,N_5078);
nand U5306 (N_5306,N_5039,N_5189);
nand U5307 (N_5307,N_5081,N_5023);
or U5308 (N_5308,N_5116,N_5175);
nor U5309 (N_5309,N_5033,N_5138);
and U5310 (N_5310,N_5128,N_5187);
and U5311 (N_5311,N_5018,N_5100);
and U5312 (N_5312,N_5042,N_5062);
and U5313 (N_5313,N_5181,N_5182);
and U5314 (N_5314,N_5139,N_5116);
and U5315 (N_5315,N_5010,N_5073);
nor U5316 (N_5316,N_5178,N_5199);
nand U5317 (N_5317,N_5164,N_5071);
and U5318 (N_5318,N_5082,N_5193);
nor U5319 (N_5319,N_5187,N_5102);
nor U5320 (N_5320,N_5173,N_5104);
xnor U5321 (N_5321,N_5085,N_5064);
and U5322 (N_5322,N_5125,N_5162);
and U5323 (N_5323,N_5132,N_5055);
nand U5324 (N_5324,N_5135,N_5027);
nor U5325 (N_5325,N_5041,N_5146);
xnor U5326 (N_5326,N_5085,N_5142);
and U5327 (N_5327,N_5060,N_5152);
nand U5328 (N_5328,N_5039,N_5043);
and U5329 (N_5329,N_5191,N_5134);
nor U5330 (N_5330,N_5097,N_5124);
nor U5331 (N_5331,N_5148,N_5160);
nor U5332 (N_5332,N_5034,N_5119);
or U5333 (N_5333,N_5122,N_5020);
and U5334 (N_5334,N_5083,N_5033);
nor U5335 (N_5335,N_5078,N_5024);
or U5336 (N_5336,N_5097,N_5066);
nand U5337 (N_5337,N_5075,N_5061);
and U5338 (N_5338,N_5028,N_5193);
nand U5339 (N_5339,N_5039,N_5025);
nand U5340 (N_5340,N_5056,N_5040);
nor U5341 (N_5341,N_5146,N_5107);
and U5342 (N_5342,N_5119,N_5101);
and U5343 (N_5343,N_5005,N_5060);
nor U5344 (N_5344,N_5000,N_5110);
or U5345 (N_5345,N_5179,N_5054);
nor U5346 (N_5346,N_5006,N_5143);
and U5347 (N_5347,N_5010,N_5016);
and U5348 (N_5348,N_5008,N_5104);
and U5349 (N_5349,N_5013,N_5152);
or U5350 (N_5350,N_5129,N_5162);
and U5351 (N_5351,N_5010,N_5088);
and U5352 (N_5352,N_5014,N_5192);
and U5353 (N_5353,N_5115,N_5146);
nand U5354 (N_5354,N_5032,N_5155);
and U5355 (N_5355,N_5198,N_5022);
nor U5356 (N_5356,N_5167,N_5191);
and U5357 (N_5357,N_5065,N_5125);
and U5358 (N_5358,N_5192,N_5103);
or U5359 (N_5359,N_5094,N_5117);
or U5360 (N_5360,N_5052,N_5142);
and U5361 (N_5361,N_5131,N_5080);
nand U5362 (N_5362,N_5132,N_5080);
xor U5363 (N_5363,N_5189,N_5022);
or U5364 (N_5364,N_5075,N_5006);
or U5365 (N_5365,N_5057,N_5099);
nor U5366 (N_5366,N_5091,N_5192);
or U5367 (N_5367,N_5020,N_5060);
or U5368 (N_5368,N_5069,N_5059);
nand U5369 (N_5369,N_5140,N_5177);
or U5370 (N_5370,N_5005,N_5042);
or U5371 (N_5371,N_5068,N_5102);
or U5372 (N_5372,N_5065,N_5083);
nand U5373 (N_5373,N_5074,N_5008);
or U5374 (N_5374,N_5197,N_5141);
and U5375 (N_5375,N_5003,N_5011);
nand U5376 (N_5376,N_5182,N_5070);
nand U5377 (N_5377,N_5020,N_5021);
and U5378 (N_5378,N_5008,N_5070);
nor U5379 (N_5379,N_5010,N_5151);
nand U5380 (N_5380,N_5158,N_5148);
xnor U5381 (N_5381,N_5098,N_5027);
nand U5382 (N_5382,N_5128,N_5057);
nand U5383 (N_5383,N_5068,N_5024);
or U5384 (N_5384,N_5039,N_5032);
nand U5385 (N_5385,N_5118,N_5187);
nor U5386 (N_5386,N_5133,N_5141);
nor U5387 (N_5387,N_5141,N_5184);
nand U5388 (N_5388,N_5096,N_5126);
or U5389 (N_5389,N_5178,N_5106);
nand U5390 (N_5390,N_5179,N_5178);
nor U5391 (N_5391,N_5035,N_5013);
nand U5392 (N_5392,N_5085,N_5138);
or U5393 (N_5393,N_5052,N_5042);
nor U5394 (N_5394,N_5136,N_5110);
nand U5395 (N_5395,N_5145,N_5048);
nand U5396 (N_5396,N_5186,N_5176);
nor U5397 (N_5397,N_5098,N_5090);
nand U5398 (N_5398,N_5169,N_5155);
nor U5399 (N_5399,N_5153,N_5146);
and U5400 (N_5400,N_5310,N_5300);
nand U5401 (N_5401,N_5276,N_5215);
nand U5402 (N_5402,N_5337,N_5328);
nor U5403 (N_5403,N_5244,N_5285);
and U5404 (N_5404,N_5303,N_5335);
nand U5405 (N_5405,N_5367,N_5237);
and U5406 (N_5406,N_5395,N_5216);
nand U5407 (N_5407,N_5295,N_5206);
and U5408 (N_5408,N_5281,N_5384);
nand U5409 (N_5409,N_5272,N_5380);
and U5410 (N_5410,N_5347,N_5266);
or U5411 (N_5411,N_5325,N_5357);
and U5412 (N_5412,N_5238,N_5280);
or U5413 (N_5413,N_5296,N_5340);
and U5414 (N_5414,N_5293,N_5366);
or U5415 (N_5415,N_5329,N_5223);
and U5416 (N_5416,N_5372,N_5332);
or U5417 (N_5417,N_5230,N_5373);
xnor U5418 (N_5418,N_5211,N_5381);
nand U5419 (N_5419,N_5256,N_5364);
and U5420 (N_5420,N_5336,N_5309);
nor U5421 (N_5421,N_5284,N_5341);
nor U5422 (N_5422,N_5360,N_5379);
and U5423 (N_5423,N_5301,N_5369);
or U5424 (N_5424,N_5339,N_5290);
or U5425 (N_5425,N_5353,N_5229);
nand U5426 (N_5426,N_5291,N_5231);
and U5427 (N_5427,N_5304,N_5343);
nor U5428 (N_5428,N_5277,N_5330);
nand U5429 (N_5429,N_5208,N_5393);
and U5430 (N_5430,N_5308,N_5365);
or U5431 (N_5431,N_5307,N_5242);
or U5432 (N_5432,N_5288,N_5265);
nand U5433 (N_5433,N_5349,N_5258);
nand U5434 (N_5434,N_5200,N_5394);
nor U5435 (N_5435,N_5204,N_5214);
and U5436 (N_5436,N_5371,N_5386);
nand U5437 (N_5437,N_5399,N_5270);
or U5438 (N_5438,N_5225,N_5207);
and U5439 (N_5439,N_5359,N_5220);
and U5440 (N_5440,N_5368,N_5283);
or U5441 (N_5441,N_5322,N_5338);
nor U5442 (N_5442,N_5385,N_5354);
nand U5443 (N_5443,N_5247,N_5370);
or U5444 (N_5444,N_5217,N_5389);
nand U5445 (N_5445,N_5375,N_5352);
and U5446 (N_5446,N_5203,N_5299);
and U5447 (N_5447,N_5344,N_5377);
or U5448 (N_5448,N_5234,N_5254);
or U5449 (N_5449,N_5317,N_5387);
nand U5450 (N_5450,N_5226,N_5252);
nor U5451 (N_5451,N_5239,N_5356);
nand U5452 (N_5452,N_5311,N_5326);
or U5453 (N_5453,N_5363,N_5355);
nand U5454 (N_5454,N_5397,N_5263);
nor U5455 (N_5455,N_5224,N_5221);
and U5456 (N_5456,N_5333,N_5320);
nand U5457 (N_5457,N_5294,N_5378);
or U5458 (N_5458,N_5228,N_5313);
nand U5459 (N_5459,N_5305,N_5271);
nor U5460 (N_5460,N_5323,N_5348);
or U5461 (N_5461,N_5334,N_5345);
and U5462 (N_5462,N_5398,N_5302);
and U5463 (N_5463,N_5262,N_5241);
or U5464 (N_5464,N_5315,N_5282);
or U5465 (N_5465,N_5261,N_5321);
nor U5466 (N_5466,N_5209,N_5318);
xor U5467 (N_5467,N_5362,N_5374);
and U5468 (N_5468,N_5286,N_5289);
nand U5469 (N_5469,N_5264,N_5253);
and U5470 (N_5470,N_5312,N_5213);
nor U5471 (N_5471,N_5350,N_5298);
or U5472 (N_5472,N_5331,N_5248);
and U5473 (N_5473,N_5383,N_5324);
nor U5474 (N_5474,N_5235,N_5269);
or U5475 (N_5475,N_5251,N_5245);
nand U5476 (N_5476,N_5314,N_5205);
and U5477 (N_5477,N_5240,N_5278);
and U5478 (N_5478,N_5358,N_5232);
nand U5479 (N_5479,N_5292,N_5361);
xnor U5480 (N_5480,N_5273,N_5279);
or U5481 (N_5481,N_5259,N_5257);
nor U5482 (N_5482,N_5319,N_5351);
nor U5483 (N_5483,N_5246,N_5227);
nor U5484 (N_5484,N_5202,N_5268);
and U5485 (N_5485,N_5316,N_5243);
or U5486 (N_5486,N_5342,N_5249);
nor U5487 (N_5487,N_5222,N_5233);
xor U5488 (N_5488,N_5274,N_5390);
nor U5489 (N_5489,N_5236,N_5297);
or U5490 (N_5490,N_5212,N_5388);
nor U5491 (N_5491,N_5327,N_5275);
nand U5492 (N_5492,N_5382,N_5346);
or U5493 (N_5493,N_5250,N_5391);
and U5494 (N_5494,N_5210,N_5392);
or U5495 (N_5495,N_5201,N_5260);
and U5496 (N_5496,N_5376,N_5306);
nor U5497 (N_5497,N_5219,N_5287);
and U5498 (N_5498,N_5396,N_5255);
nand U5499 (N_5499,N_5218,N_5267);
and U5500 (N_5500,N_5360,N_5341);
and U5501 (N_5501,N_5233,N_5296);
or U5502 (N_5502,N_5282,N_5335);
nand U5503 (N_5503,N_5213,N_5369);
or U5504 (N_5504,N_5274,N_5391);
and U5505 (N_5505,N_5352,N_5229);
or U5506 (N_5506,N_5221,N_5204);
and U5507 (N_5507,N_5356,N_5207);
nor U5508 (N_5508,N_5391,N_5253);
nor U5509 (N_5509,N_5207,N_5384);
or U5510 (N_5510,N_5340,N_5206);
or U5511 (N_5511,N_5240,N_5372);
nand U5512 (N_5512,N_5374,N_5257);
or U5513 (N_5513,N_5286,N_5355);
or U5514 (N_5514,N_5333,N_5356);
or U5515 (N_5515,N_5300,N_5313);
nand U5516 (N_5516,N_5337,N_5362);
or U5517 (N_5517,N_5305,N_5328);
or U5518 (N_5518,N_5380,N_5305);
or U5519 (N_5519,N_5296,N_5355);
and U5520 (N_5520,N_5315,N_5305);
or U5521 (N_5521,N_5357,N_5291);
nor U5522 (N_5522,N_5231,N_5263);
nor U5523 (N_5523,N_5271,N_5211);
and U5524 (N_5524,N_5352,N_5261);
or U5525 (N_5525,N_5285,N_5380);
nor U5526 (N_5526,N_5276,N_5236);
or U5527 (N_5527,N_5263,N_5277);
and U5528 (N_5528,N_5269,N_5274);
or U5529 (N_5529,N_5261,N_5385);
nor U5530 (N_5530,N_5354,N_5226);
nand U5531 (N_5531,N_5258,N_5290);
nand U5532 (N_5532,N_5374,N_5286);
nand U5533 (N_5533,N_5316,N_5268);
and U5534 (N_5534,N_5368,N_5345);
and U5535 (N_5535,N_5350,N_5385);
and U5536 (N_5536,N_5212,N_5234);
xnor U5537 (N_5537,N_5283,N_5323);
nor U5538 (N_5538,N_5206,N_5211);
nand U5539 (N_5539,N_5221,N_5395);
or U5540 (N_5540,N_5305,N_5253);
or U5541 (N_5541,N_5274,N_5348);
nand U5542 (N_5542,N_5284,N_5391);
and U5543 (N_5543,N_5280,N_5219);
nor U5544 (N_5544,N_5283,N_5397);
nand U5545 (N_5545,N_5316,N_5284);
and U5546 (N_5546,N_5261,N_5335);
nand U5547 (N_5547,N_5270,N_5201);
nand U5548 (N_5548,N_5315,N_5279);
nor U5549 (N_5549,N_5237,N_5329);
nor U5550 (N_5550,N_5335,N_5365);
and U5551 (N_5551,N_5250,N_5398);
or U5552 (N_5552,N_5344,N_5205);
nor U5553 (N_5553,N_5209,N_5381);
xnor U5554 (N_5554,N_5323,N_5389);
and U5555 (N_5555,N_5370,N_5267);
nand U5556 (N_5556,N_5346,N_5370);
and U5557 (N_5557,N_5352,N_5346);
nor U5558 (N_5558,N_5344,N_5206);
or U5559 (N_5559,N_5213,N_5204);
or U5560 (N_5560,N_5362,N_5270);
nor U5561 (N_5561,N_5274,N_5385);
nand U5562 (N_5562,N_5215,N_5336);
nand U5563 (N_5563,N_5381,N_5341);
nand U5564 (N_5564,N_5247,N_5228);
nor U5565 (N_5565,N_5272,N_5291);
nand U5566 (N_5566,N_5279,N_5359);
nor U5567 (N_5567,N_5325,N_5282);
or U5568 (N_5568,N_5376,N_5264);
and U5569 (N_5569,N_5240,N_5243);
nor U5570 (N_5570,N_5272,N_5221);
nor U5571 (N_5571,N_5223,N_5284);
and U5572 (N_5572,N_5318,N_5236);
or U5573 (N_5573,N_5278,N_5368);
nor U5574 (N_5574,N_5203,N_5346);
nor U5575 (N_5575,N_5305,N_5396);
nand U5576 (N_5576,N_5262,N_5215);
or U5577 (N_5577,N_5243,N_5378);
and U5578 (N_5578,N_5346,N_5301);
and U5579 (N_5579,N_5331,N_5301);
nand U5580 (N_5580,N_5275,N_5339);
or U5581 (N_5581,N_5340,N_5365);
nor U5582 (N_5582,N_5338,N_5346);
or U5583 (N_5583,N_5320,N_5326);
nor U5584 (N_5584,N_5207,N_5313);
or U5585 (N_5585,N_5330,N_5280);
and U5586 (N_5586,N_5207,N_5338);
or U5587 (N_5587,N_5282,N_5219);
nor U5588 (N_5588,N_5303,N_5383);
nand U5589 (N_5589,N_5295,N_5354);
and U5590 (N_5590,N_5297,N_5232);
xor U5591 (N_5591,N_5226,N_5294);
and U5592 (N_5592,N_5353,N_5250);
or U5593 (N_5593,N_5253,N_5205);
nor U5594 (N_5594,N_5354,N_5281);
nand U5595 (N_5595,N_5317,N_5303);
or U5596 (N_5596,N_5308,N_5318);
and U5597 (N_5597,N_5272,N_5294);
or U5598 (N_5598,N_5357,N_5220);
or U5599 (N_5599,N_5340,N_5273);
and U5600 (N_5600,N_5412,N_5583);
nand U5601 (N_5601,N_5507,N_5433);
nor U5602 (N_5602,N_5581,N_5545);
nand U5603 (N_5603,N_5520,N_5506);
or U5604 (N_5604,N_5510,N_5411);
and U5605 (N_5605,N_5477,N_5423);
nor U5606 (N_5606,N_5593,N_5453);
nand U5607 (N_5607,N_5525,N_5558);
or U5608 (N_5608,N_5511,N_5447);
or U5609 (N_5609,N_5562,N_5574);
and U5610 (N_5610,N_5535,N_5564);
nand U5611 (N_5611,N_5484,N_5554);
or U5612 (N_5612,N_5552,N_5408);
and U5613 (N_5613,N_5572,N_5424);
nand U5614 (N_5614,N_5565,N_5584);
nand U5615 (N_5615,N_5529,N_5464);
nand U5616 (N_5616,N_5560,N_5595);
nand U5617 (N_5617,N_5589,N_5566);
and U5618 (N_5618,N_5547,N_5480);
nor U5619 (N_5619,N_5542,N_5556);
nand U5620 (N_5620,N_5540,N_5435);
or U5621 (N_5621,N_5561,N_5452);
nor U5622 (N_5622,N_5430,N_5549);
and U5623 (N_5623,N_5505,N_5519);
nand U5624 (N_5624,N_5439,N_5587);
or U5625 (N_5625,N_5489,N_5596);
nand U5626 (N_5626,N_5557,N_5450);
and U5627 (N_5627,N_5448,N_5479);
or U5628 (N_5628,N_5509,N_5444);
nor U5629 (N_5629,N_5577,N_5481);
nor U5630 (N_5630,N_5537,N_5592);
nor U5631 (N_5631,N_5528,N_5418);
or U5632 (N_5632,N_5585,N_5404);
and U5633 (N_5633,N_5534,N_5555);
or U5634 (N_5634,N_5533,N_5413);
nor U5635 (N_5635,N_5573,N_5449);
nor U5636 (N_5636,N_5475,N_5499);
and U5637 (N_5637,N_5586,N_5512);
or U5638 (N_5638,N_5590,N_5419);
or U5639 (N_5639,N_5491,N_5454);
nor U5640 (N_5640,N_5594,N_5472);
nand U5641 (N_5641,N_5523,N_5410);
or U5642 (N_5642,N_5429,N_5548);
nand U5643 (N_5643,N_5403,N_5446);
nand U5644 (N_5644,N_5567,N_5437);
or U5645 (N_5645,N_5417,N_5569);
or U5646 (N_5646,N_5400,N_5456);
nor U5647 (N_5647,N_5597,N_5451);
and U5648 (N_5648,N_5527,N_5427);
nor U5649 (N_5649,N_5508,N_5498);
nand U5650 (N_5650,N_5471,N_5582);
and U5651 (N_5651,N_5482,N_5405);
nor U5652 (N_5652,N_5473,N_5468);
and U5653 (N_5653,N_5436,N_5467);
or U5654 (N_5654,N_5459,N_5531);
nor U5655 (N_5655,N_5493,N_5541);
or U5656 (N_5656,N_5538,N_5500);
nand U5657 (N_5657,N_5492,N_5463);
and U5658 (N_5658,N_5474,N_5470);
nand U5659 (N_5659,N_5536,N_5571);
nand U5660 (N_5660,N_5425,N_5422);
nand U5661 (N_5661,N_5461,N_5440);
nor U5662 (N_5662,N_5563,N_5460);
nor U5663 (N_5663,N_5504,N_5434);
and U5664 (N_5664,N_5465,N_5416);
nor U5665 (N_5665,N_5522,N_5515);
nor U5666 (N_5666,N_5490,N_5544);
or U5667 (N_5667,N_5438,N_5469);
nand U5668 (N_5668,N_5501,N_5513);
or U5669 (N_5669,N_5526,N_5441);
or U5670 (N_5670,N_5455,N_5550);
or U5671 (N_5671,N_5503,N_5495);
or U5672 (N_5672,N_5426,N_5406);
and U5673 (N_5673,N_5532,N_5524);
nand U5674 (N_5674,N_5517,N_5543);
nand U5675 (N_5675,N_5575,N_5466);
and U5676 (N_5676,N_5591,N_5485);
and U5677 (N_5677,N_5570,N_5559);
nor U5678 (N_5678,N_5445,N_5443);
xnor U5679 (N_5679,N_5431,N_5487);
or U5680 (N_5680,N_5402,N_5553);
nor U5681 (N_5681,N_5476,N_5432);
or U5682 (N_5682,N_5457,N_5580);
nor U5683 (N_5683,N_5420,N_5428);
nand U5684 (N_5684,N_5478,N_5598);
nand U5685 (N_5685,N_5539,N_5483);
or U5686 (N_5686,N_5462,N_5486);
nor U5687 (N_5687,N_5599,N_5421);
and U5688 (N_5688,N_5516,N_5514);
nand U5689 (N_5689,N_5414,N_5497);
and U5690 (N_5690,N_5568,N_5488);
nand U5691 (N_5691,N_5409,N_5494);
or U5692 (N_5692,N_5579,N_5415);
nand U5693 (N_5693,N_5442,N_5551);
nor U5694 (N_5694,N_5578,N_5518);
xor U5695 (N_5695,N_5458,N_5496);
nand U5696 (N_5696,N_5401,N_5521);
and U5697 (N_5697,N_5407,N_5588);
nor U5698 (N_5698,N_5502,N_5546);
nor U5699 (N_5699,N_5576,N_5530);
or U5700 (N_5700,N_5540,N_5593);
and U5701 (N_5701,N_5483,N_5455);
or U5702 (N_5702,N_5547,N_5548);
nor U5703 (N_5703,N_5566,N_5424);
nand U5704 (N_5704,N_5446,N_5503);
nor U5705 (N_5705,N_5511,N_5561);
nand U5706 (N_5706,N_5457,N_5436);
nor U5707 (N_5707,N_5459,N_5533);
nor U5708 (N_5708,N_5459,N_5568);
or U5709 (N_5709,N_5524,N_5442);
nand U5710 (N_5710,N_5551,N_5411);
nand U5711 (N_5711,N_5537,N_5476);
nand U5712 (N_5712,N_5405,N_5531);
or U5713 (N_5713,N_5421,N_5575);
nand U5714 (N_5714,N_5531,N_5518);
nand U5715 (N_5715,N_5467,N_5488);
and U5716 (N_5716,N_5433,N_5474);
nand U5717 (N_5717,N_5566,N_5439);
and U5718 (N_5718,N_5476,N_5492);
nor U5719 (N_5719,N_5480,N_5577);
nor U5720 (N_5720,N_5456,N_5485);
or U5721 (N_5721,N_5491,N_5463);
and U5722 (N_5722,N_5496,N_5549);
nand U5723 (N_5723,N_5508,N_5431);
or U5724 (N_5724,N_5442,N_5431);
nor U5725 (N_5725,N_5509,N_5513);
xor U5726 (N_5726,N_5520,N_5559);
or U5727 (N_5727,N_5541,N_5543);
xor U5728 (N_5728,N_5435,N_5507);
nand U5729 (N_5729,N_5472,N_5452);
nor U5730 (N_5730,N_5549,N_5484);
or U5731 (N_5731,N_5534,N_5596);
nand U5732 (N_5732,N_5479,N_5559);
nor U5733 (N_5733,N_5537,N_5591);
nor U5734 (N_5734,N_5465,N_5411);
nand U5735 (N_5735,N_5524,N_5506);
or U5736 (N_5736,N_5487,N_5581);
nand U5737 (N_5737,N_5593,N_5530);
nand U5738 (N_5738,N_5553,N_5549);
nor U5739 (N_5739,N_5566,N_5434);
nor U5740 (N_5740,N_5543,N_5524);
and U5741 (N_5741,N_5428,N_5589);
nor U5742 (N_5742,N_5422,N_5437);
and U5743 (N_5743,N_5404,N_5469);
xor U5744 (N_5744,N_5582,N_5514);
or U5745 (N_5745,N_5579,N_5542);
nor U5746 (N_5746,N_5465,N_5460);
nor U5747 (N_5747,N_5512,N_5418);
or U5748 (N_5748,N_5563,N_5447);
nand U5749 (N_5749,N_5528,N_5434);
or U5750 (N_5750,N_5489,N_5542);
or U5751 (N_5751,N_5489,N_5517);
xnor U5752 (N_5752,N_5429,N_5462);
and U5753 (N_5753,N_5405,N_5489);
nor U5754 (N_5754,N_5417,N_5592);
and U5755 (N_5755,N_5477,N_5536);
nand U5756 (N_5756,N_5544,N_5456);
or U5757 (N_5757,N_5446,N_5505);
nor U5758 (N_5758,N_5432,N_5588);
nor U5759 (N_5759,N_5401,N_5456);
nor U5760 (N_5760,N_5440,N_5578);
nand U5761 (N_5761,N_5487,N_5476);
nand U5762 (N_5762,N_5433,N_5552);
and U5763 (N_5763,N_5406,N_5413);
nor U5764 (N_5764,N_5423,N_5461);
nand U5765 (N_5765,N_5571,N_5477);
and U5766 (N_5766,N_5461,N_5596);
and U5767 (N_5767,N_5420,N_5507);
and U5768 (N_5768,N_5594,N_5476);
nor U5769 (N_5769,N_5522,N_5530);
nor U5770 (N_5770,N_5434,N_5512);
nor U5771 (N_5771,N_5453,N_5514);
and U5772 (N_5772,N_5562,N_5458);
and U5773 (N_5773,N_5489,N_5598);
and U5774 (N_5774,N_5422,N_5441);
and U5775 (N_5775,N_5580,N_5462);
nor U5776 (N_5776,N_5448,N_5532);
nand U5777 (N_5777,N_5402,N_5439);
xnor U5778 (N_5778,N_5512,N_5475);
and U5779 (N_5779,N_5558,N_5492);
nand U5780 (N_5780,N_5511,N_5421);
xnor U5781 (N_5781,N_5531,N_5578);
nor U5782 (N_5782,N_5568,N_5401);
and U5783 (N_5783,N_5576,N_5443);
and U5784 (N_5784,N_5432,N_5517);
and U5785 (N_5785,N_5433,N_5461);
or U5786 (N_5786,N_5441,N_5519);
and U5787 (N_5787,N_5408,N_5415);
nand U5788 (N_5788,N_5439,N_5517);
and U5789 (N_5789,N_5461,N_5404);
nand U5790 (N_5790,N_5561,N_5527);
xor U5791 (N_5791,N_5481,N_5568);
nor U5792 (N_5792,N_5566,N_5490);
or U5793 (N_5793,N_5462,N_5574);
nor U5794 (N_5794,N_5416,N_5404);
nor U5795 (N_5795,N_5497,N_5432);
or U5796 (N_5796,N_5516,N_5433);
nor U5797 (N_5797,N_5574,N_5420);
nor U5798 (N_5798,N_5430,N_5478);
xor U5799 (N_5799,N_5463,N_5560);
nor U5800 (N_5800,N_5688,N_5782);
and U5801 (N_5801,N_5638,N_5717);
and U5802 (N_5802,N_5628,N_5654);
nand U5803 (N_5803,N_5612,N_5622);
and U5804 (N_5804,N_5765,N_5726);
nand U5805 (N_5805,N_5798,N_5696);
xnor U5806 (N_5806,N_5625,N_5646);
nor U5807 (N_5807,N_5775,N_5602);
and U5808 (N_5808,N_5663,N_5670);
nor U5809 (N_5809,N_5751,N_5614);
or U5810 (N_5810,N_5732,N_5637);
and U5811 (N_5811,N_5675,N_5705);
nor U5812 (N_5812,N_5655,N_5746);
or U5813 (N_5813,N_5716,N_5710);
nor U5814 (N_5814,N_5785,N_5615);
and U5815 (N_5815,N_5649,N_5668);
or U5816 (N_5816,N_5647,N_5728);
nor U5817 (N_5817,N_5661,N_5767);
or U5818 (N_5818,N_5747,N_5677);
and U5819 (N_5819,N_5764,N_5773);
nor U5820 (N_5820,N_5621,N_5691);
nand U5821 (N_5821,N_5632,N_5666);
nor U5822 (N_5822,N_5617,N_5695);
nand U5823 (N_5823,N_5650,N_5757);
or U5824 (N_5824,N_5703,N_5680);
and U5825 (N_5825,N_5715,N_5772);
nand U5826 (N_5826,N_5748,N_5673);
or U5827 (N_5827,N_5712,N_5722);
and U5828 (N_5828,N_5708,N_5641);
or U5829 (N_5829,N_5687,N_5724);
nand U5830 (N_5830,N_5718,N_5657);
nand U5831 (N_5831,N_5627,N_5642);
nor U5832 (N_5832,N_5603,N_5733);
nand U5833 (N_5833,N_5743,N_5636);
and U5834 (N_5834,N_5684,N_5634);
nand U5835 (N_5835,N_5788,N_5692);
or U5836 (N_5836,N_5750,N_5660);
and U5837 (N_5837,N_5601,N_5643);
nor U5838 (N_5838,N_5653,N_5674);
xnor U5839 (N_5839,N_5709,N_5701);
nand U5840 (N_5840,N_5699,N_5608);
and U5841 (N_5841,N_5793,N_5790);
and U5842 (N_5842,N_5753,N_5781);
or U5843 (N_5843,N_5662,N_5763);
nor U5844 (N_5844,N_5734,N_5783);
nor U5845 (N_5845,N_5635,N_5706);
and U5846 (N_5846,N_5776,N_5707);
or U5847 (N_5847,N_5607,N_5784);
or U5848 (N_5848,N_5774,N_5623);
nand U5849 (N_5849,N_5780,N_5685);
or U5850 (N_5850,N_5762,N_5754);
nand U5851 (N_5851,N_5604,N_5629);
nand U5852 (N_5852,N_5698,N_5609);
and U5853 (N_5853,N_5624,N_5766);
or U5854 (N_5854,N_5620,N_5669);
and U5855 (N_5855,N_5752,N_5659);
nand U5856 (N_5856,N_5664,N_5606);
and U5857 (N_5857,N_5678,N_5679);
and U5858 (N_5858,N_5720,N_5714);
nand U5859 (N_5859,N_5742,N_5711);
nor U5860 (N_5860,N_5791,N_5789);
and U5861 (N_5861,N_5769,N_5713);
nor U5862 (N_5862,N_5690,N_5656);
and U5863 (N_5863,N_5741,N_5744);
and U5864 (N_5864,N_5723,N_5600);
nor U5865 (N_5865,N_5749,N_5619);
nand U5866 (N_5866,N_5768,N_5702);
nor U5867 (N_5867,N_5796,N_5787);
nand U5868 (N_5868,N_5770,N_5738);
and U5869 (N_5869,N_5755,N_5760);
nor U5870 (N_5870,N_5739,N_5777);
nor U5871 (N_5871,N_5651,N_5644);
nand U5872 (N_5872,N_5616,N_5693);
nand U5873 (N_5873,N_5737,N_5756);
nor U5874 (N_5874,N_5745,N_5731);
and U5875 (N_5875,N_5697,N_5648);
nand U5876 (N_5876,N_5671,N_5652);
and U5877 (N_5877,N_5792,N_5672);
nand U5878 (N_5878,N_5771,N_5719);
and U5879 (N_5879,N_5676,N_5639);
nor U5880 (N_5880,N_5740,N_5758);
and U5881 (N_5881,N_5729,N_5799);
nand U5882 (N_5882,N_5730,N_5658);
nor U5883 (N_5883,N_5794,N_5683);
nor U5884 (N_5884,N_5700,N_5682);
xor U5885 (N_5885,N_5633,N_5631);
nand U5886 (N_5886,N_5727,N_5665);
or U5887 (N_5887,N_5681,N_5626);
and U5888 (N_5888,N_5618,N_5761);
and U5889 (N_5889,N_5797,N_5640);
and U5890 (N_5890,N_5667,N_5611);
nand U5891 (N_5891,N_5689,N_5735);
and U5892 (N_5892,N_5704,N_5694);
nand U5893 (N_5893,N_5786,N_5795);
nand U5894 (N_5894,N_5613,N_5721);
nor U5895 (N_5895,N_5645,N_5759);
or U5896 (N_5896,N_5778,N_5630);
or U5897 (N_5897,N_5779,N_5736);
nor U5898 (N_5898,N_5686,N_5725);
or U5899 (N_5899,N_5605,N_5610);
nand U5900 (N_5900,N_5798,N_5698);
and U5901 (N_5901,N_5715,N_5769);
nand U5902 (N_5902,N_5632,N_5604);
and U5903 (N_5903,N_5604,N_5796);
and U5904 (N_5904,N_5727,N_5620);
nor U5905 (N_5905,N_5603,N_5625);
and U5906 (N_5906,N_5640,N_5796);
or U5907 (N_5907,N_5791,N_5652);
and U5908 (N_5908,N_5774,N_5663);
and U5909 (N_5909,N_5717,N_5675);
and U5910 (N_5910,N_5788,N_5689);
or U5911 (N_5911,N_5734,N_5702);
nor U5912 (N_5912,N_5629,N_5792);
or U5913 (N_5913,N_5666,N_5748);
or U5914 (N_5914,N_5786,N_5722);
or U5915 (N_5915,N_5643,N_5782);
and U5916 (N_5916,N_5684,N_5733);
nand U5917 (N_5917,N_5643,N_5739);
and U5918 (N_5918,N_5648,N_5619);
nand U5919 (N_5919,N_5686,N_5660);
nor U5920 (N_5920,N_5760,N_5771);
nand U5921 (N_5921,N_5781,N_5745);
xor U5922 (N_5922,N_5733,N_5676);
nand U5923 (N_5923,N_5689,N_5723);
and U5924 (N_5924,N_5666,N_5641);
nor U5925 (N_5925,N_5746,N_5620);
xor U5926 (N_5926,N_5729,N_5653);
and U5927 (N_5927,N_5620,N_5662);
nor U5928 (N_5928,N_5791,N_5736);
or U5929 (N_5929,N_5752,N_5638);
and U5930 (N_5930,N_5715,N_5675);
or U5931 (N_5931,N_5783,N_5634);
or U5932 (N_5932,N_5704,N_5678);
or U5933 (N_5933,N_5736,N_5623);
and U5934 (N_5934,N_5788,N_5718);
nor U5935 (N_5935,N_5724,N_5618);
nand U5936 (N_5936,N_5736,N_5690);
nor U5937 (N_5937,N_5624,N_5731);
or U5938 (N_5938,N_5701,N_5691);
nand U5939 (N_5939,N_5745,N_5637);
nand U5940 (N_5940,N_5609,N_5620);
or U5941 (N_5941,N_5607,N_5708);
and U5942 (N_5942,N_5731,N_5799);
nand U5943 (N_5943,N_5634,N_5747);
or U5944 (N_5944,N_5753,N_5718);
nand U5945 (N_5945,N_5770,N_5665);
or U5946 (N_5946,N_5701,N_5649);
or U5947 (N_5947,N_5766,N_5721);
nand U5948 (N_5948,N_5736,N_5748);
and U5949 (N_5949,N_5654,N_5756);
nand U5950 (N_5950,N_5630,N_5633);
nand U5951 (N_5951,N_5742,N_5764);
xor U5952 (N_5952,N_5764,N_5687);
nor U5953 (N_5953,N_5730,N_5677);
nor U5954 (N_5954,N_5632,N_5772);
nand U5955 (N_5955,N_5746,N_5777);
nand U5956 (N_5956,N_5653,N_5675);
or U5957 (N_5957,N_5784,N_5679);
or U5958 (N_5958,N_5776,N_5604);
and U5959 (N_5959,N_5748,N_5773);
nor U5960 (N_5960,N_5683,N_5754);
or U5961 (N_5961,N_5726,N_5794);
and U5962 (N_5962,N_5646,N_5651);
and U5963 (N_5963,N_5622,N_5661);
nor U5964 (N_5964,N_5771,N_5779);
nand U5965 (N_5965,N_5664,N_5608);
and U5966 (N_5966,N_5615,N_5610);
nor U5967 (N_5967,N_5661,N_5609);
or U5968 (N_5968,N_5779,N_5618);
nor U5969 (N_5969,N_5695,N_5609);
nand U5970 (N_5970,N_5727,N_5790);
and U5971 (N_5971,N_5798,N_5742);
or U5972 (N_5972,N_5602,N_5723);
and U5973 (N_5973,N_5761,N_5721);
nand U5974 (N_5974,N_5683,N_5712);
nor U5975 (N_5975,N_5652,N_5609);
and U5976 (N_5976,N_5727,N_5607);
nor U5977 (N_5977,N_5685,N_5644);
or U5978 (N_5978,N_5691,N_5770);
nor U5979 (N_5979,N_5762,N_5678);
or U5980 (N_5980,N_5732,N_5652);
or U5981 (N_5981,N_5754,N_5743);
and U5982 (N_5982,N_5644,N_5625);
nor U5983 (N_5983,N_5708,N_5692);
nand U5984 (N_5984,N_5608,N_5767);
nand U5985 (N_5985,N_5616,N_5740);
and U5986 (N_5986,N_5685,N_5763);
xor U5987 (N_5987,N_5714,N_5611);
nor U5988 (N_5988,N_5713,N_5771);
nand U5989 (N_5989,N_5675,N_5677);
or U5990 (N_5990,N_5600,N_5795);
or U5991 (N_5991,N_5695,N_5668);
and U5992 (N_5992,N_5793,N_5794);
nand U5993 (N_5993,N_5693,N_5791);
or U5994 (N_5994,N_5787,N_5778);
nand U5995 (N_5995,N_5675,N_5735);
nand U5996 (N_5996,N_5732,N_5759);
and U5997 (N_5997,N_5713,N_5668);
and U5998 (N_5998,N_5676,N_5654);
nor U5999 (N_5999,N_5729,N_5762);
nor U6000 (N_6000,N_5832,N_5840);
nand U6001 (N_6001,N_5970,N_5962);
and U6002 (N_6002,N_5874,N_5895);
nand U6003 (N_6003,N_5806,N_5825);
or U6004 (N_6004,N_5887,N_5995);
or U6005 (N_6005,N_5842,N_5977);
or U6006 (N_6006,N_5921,N_5916);
nand U6007 (N_6007,N_5903,N_5989);
nand U6008 (N_6008,N_5841,N_5915);
nand U6009 (N_6009,N_5848,N_5867);
and U6010 (N_6010,N_5890,N_5966);
and U6011 (N_6011,N_5967,N_5932);
nor U6012 (N_6012,N_5885,N_5873);
nor U6013 (N_6013,N_5991,N_5843);
nor U6014 (N_6014,N_5815,N_5870);
nor U6015 (N_6015,N_5868,N_5853);
nand U6016 (N_6016,N_5944,N_5951);
and U6017 (N_6017,N_5802,N_5892);
or U6018 (N_6018,N_5845,N_5830);
and U6019 (N_6019,N_5947,N_5985);
or U6020 (N_6020,N_5898,N_5902);
and U6021 (N_6021,N_5877,N_5955);
nand U6022 (N_6022,N_5931,N_5837);
nand U6023 (N_6023,N_5864,N_5942);
nand U6024 (N_6024,N_5922,N_5835);
and U6025 (N_6025,N_5984,N_5974);
and U6026 (N_6026,N_5987,N_5838);
nor U6027 (N_6027,N_5833,N_5846);
or U6028 (N_6028,N_5899,N_5928);
and U6029 (N_6029,N_5959,N_5847);
xnor U6030 (N_6030,N_5904,N_5956);
nor U6031 (N_6031,N_5935,N_5986);
and U6032 (N_6032,N_5816,N_5896);
or U6033 (N_6033,N_5945,N_5957);
and U6034 (N_6034,N_5858,N_5836);
nor U6035 (N_6035,N_5851,N_5905);
and U6036 (N_6036,N_5934,N_5844);
nor U6037 (N_6037,N_5924,N_5981);
nand U6038 (N_6038,N_5807,N_5879);
or U6039 (N_6039,N_5950,N_5997);
nor U6040 (N_6040,N_5855,N_5949);
or U6041 (N_6041,N_5961,N_5866);
or U6042 (N_6042,N_5882,N_5814);
nor U6043 (N_6043,N_5818,N_5834);
nor U6044 (N_6044,N_5828,N_5875);
or U6045 (N_6045,N_5865,N_5958);
and U6046 (N_6046,N_5952,N_5943);
nand U6047 (N_6047,N_5983,N_5960);
or U6048 (N_6048,N_5876,N_5859);
and U6049 (N_6049,N_5831,N_5948);
xor U6050 (N_6050,N_5999,N_5979);
and U6051 (N_6051,N_5886,N_5976);
or U6052 (N_6052,N_5897,N_5857);
nor U6053 (N_6053,N_5860,N_5996);
nand U6054 (N_6054,N_5972,N_5880);
nand U6055 (N_6055,N_5936,N_5888);
and U6056 (N_6056,N_5988,N_5881);
xnor U6057 (N_6057,N_5920,N_5964);
and U6058 (N_6058,N_5809,N_5893);
or U6059 (N_6059,N_5819,N_5990);
xnor U6060 (N_6060,N_5805,N_5965);
nor U6061 (N_6061,N_5939,N_5808);
or U6062 (N_6062,N_5852,N_5803);
or U6063 (N_6063,N_5827,N_5817);
nand U6064 (N_6064,N_5938,N_5813);
and U6065 (N_6065,N_5810,N_5884);
nor U6066 (N_6066,N_5980,N_5918);
nor U6067 (N_6067,N_5971,N_5993);
nor U6068 (N_6068,N_5953,N_5909);
nand U6069 (N_6069,N_5871,N_5878);
nor U6070 (N_6070,N_5969,N_5992);
and U6071 (N_6071,N_5925,N_5926);
nor U6072 (N_6072,N_5839,N_5849);
nor U6073 (N_6073,N_5973,N_5927);
and U6074 (N_6074,N_5941,N_5946);
nand U6075 (N_6075,N_5824,N_5923);
and U6076 (N_6076,N_5906,N_5863);
or U6077 (N_6077,N_5917,N_5912);
and U6078 (N_6078,N_5856,N_5968);
or U6079 (N_6079,N_5933,N_5911);
nor U6080 (N_6080,N_5889,N_5894);
or U6081 (N_6081,N_5929,N_5900);
nor U6082 (N_6082,N_5891,N_5801);
nand U6083 (N_6083,N_5908,N_5883);
nand U6084 (N_6084,N_5910,N_5998);
or U6085 (N_6085,N_5861,N_5850);
and U6086 (N_6086,N_5869,N_5978);
or U6087 (N_6087,N_5913,N_5982);
nand U6088 (N_6088,N_5930,N_5812);
and U6089 (N_6089,N_5901,N_5862);
nor U6090 (N_6090,N_5994,N_5975);
or U6091 (N_6091,N_5829,N_5811);
nor U6092 (N_6092,N_5800,N_5919);
and U6093 (N_6093,N_5872,N_5821);
and U6094 (N_6094,N_5940,N_5822);
xnor U6095 (N_6095,N_5914,N_5954);
and U6096 (N_6096,N_5854,N_5804);
nor U6097 (N_6097,N_5907,N_5963);
nand U6098 (N_6098,N_5937,N_5820);
nor U6099 (N_6099,N_5826,N_5823);
or U6100 (N_6100,N_5984,N_5875);
nor U6101 (N_6101,N_5959,N_5854);
and U6102 (N_6102,N_5970,N_5951);
nand U6103 (N_6103,N_5853,N_5971);
or U6104 (N_6104,N_5972,N_5840);
nand U6105 (N_6105,N_5869,N_5952);
or U6106 (N_6106,N_5879,N_5804);
nor U6107 (N_6107,N_5904,N_5932);
or U6108 (N_6108,N_5890,N_5879);
nand U6109 (N_6109,N_5867,N_5820);
and U6110 (N_6110,N_5933,N_5890);
nor U6111 (N_6111,N_5914,N_5919);
or U6112 (N_6112,N_5962,N_5994);
nor U6113 (N_6113,N_5950,N_5966);
or U6114 (N_6114,N_5891,N_5896);
nor U6115 (N_6115,N_5901,N_5971);
nand U6116 (N_6116,N_5801,N_5803);
and U6117 (N_6117,N_5974,N_5923);
nor U6118 (N_6118,N_5846,N_5939);
nand U6119 (N_6119,N_5971,N_5968);
and U6120 (N_6120,N_5974,N_5925);
nor U6121 (N_6121,N_5830,N_5860);
and U6122 (N_6122,N_5817,N_5936);
nand U6123 (N_6123,N_5839,N_5868);
or U6124 (N_6124,N_5822,N_5834);
nand U6125 (N_6125,N_5873,N_5818);
nor U6126 (N_6126,N_5941,N_5932);
xor U6127 (N_6127,N_5980,N_5981);
or U6128 (N_6128,N_5886,N_5968);
and U6129 (N_6129,N_5898,N_5862);
or U6130 (N_6130,N_5873,N_5970);
nor U6131 (N_6131,N_5959,N_5957);
nor U6132 (N_6132,N_5922,N_5942);
or U6133 (N_6133,N_5894,N_5954);
or U6134 (N_6134,N_5905,N_5857);
nor U6135 (N_6135,N_5808,N_5863);
and U6136 (N_6136,N_5959,N_5816);
nor U6137 (N_6137,N_5885,N_5895);
nand U6138 (N_6138,N_5904,N_5971);
or U6139 (N_6139,N_5980,N_5948);
and U6140 (N_6140,N_5880,N_5976);
nand U6141 (N_6141,N_5929,N_5974);
nor U6142 (N_6142,N_5841,N_5973);
nand U6143 (N_6143,N_5973,N_5899);
xor U6144 (N_6144,N_5969,N_5852);
nand U6145 (N_6145,N_5819,N_5891);
nor U6146 (N_6146,N_5886,N_5930);
or U6147 (N_6147,N_5970,N_5938);
and U6148 (N_6148,N_5888,N_5841);
or U6149 (N_6149,N_5978,N_5800);
nor U6150 (N_6150,N_5876,N_5861);
and U6151 (N_6151,N_5935,N_5921);
or U6152 (N_6152,N_5919,N_5939);
and U6153 (N_6153,N_5947,N_5917);
and U6154 (N_6154,N_5908,N_5877);
nor U6155 (N_6155,N_5938,N_5833);
or U6156 (N_6156,N_5843,N_5874);
nor U6157 (N_6157,N_5832,N_5904);
nand U6158 (N_6158,N_5990,N_5875);
and U6159 (N_6159,N_5925,N_5880);
or U6160 (N_6160,N_5933,N_5931);
and U6161 (N_6161,N_5815,N_5813);
or U6162 (N_6162,N_5836,N_5862);
and U6163 (N_6163,N_5896,N_5854);
and U6164 (N_6164,N_5969,N_5870);
nor U6165 (N_6165,N_5994,N_5845);
xor U6166 (N_6166,N_5876,N_5910);
and U6167 (N_6167,N_5998,N_5855);
nand U6168 (N_6168,N_5992,N_5931);
nor U6169 (N_6169,N_5901,N_5838);
nand U6170 (N_6170,N_5866,N_5896);
nor U6171 (N_6171,N_5953,N_5894);
and U6172 (N_6172,N_5829,N_5951);
nor U6173 (N_6173,N_5871,N_5940);
and U6174 (N_6174,N_5857,N_5941);
nand U6175 (N_6175,N_5915,N_5909);
or U6176 (N_6176,N_5953,N_5951);
or U6177 (N_6177,N_5935,N_5970);
nand U6178 (N_6178,N_5862,N_5824);
nand U6179 (N_6179,N_5869,N_5913);
xor U6180 (N_6180,N_5879,N_5982);
and U6181 (N_6181,N_5851,N_5915);
nand U6182 (N_6182,N_5913,N_5807);
nor U6183 (N_6183,N_5992,N_5807);
nand U6184 (N_6184,N_5860,N_5808);
and U6185 (N_6185,N_5953,N_5927);
or U6186 (N_6186,N_5873,N_5991);
and U6187 (N_6187,N_5994,N_5971);
nor U6188 (N_6188,N_5944,N_5830);
nor U6189 (N_6189,N_5956,N_5896);
and U6190 (N_6190,N_5947,N_5999);
and U6191 (N_6191,N_5905,N_5814);
and U6192 (N_6192,N_5872,N_5838);
nor U6193 (N_6193,N_5955,N_5951);
nor U6194 (N_6194,N_5868,N_5964);
nor U6195 (N_6195,N_5857,N_5917);
nand U6196 (N_6196,N_5862,N_5944);
or U6197 (N_6197,N_5937,N_5956);
or U6198 (N_6198,N_5951,N_5958);
nor U6199 (N_6199,N_5889,N_5971);
nor U6200 (N_6200,N_6001,N_6016);
nand U6201 (N_6201,N_6124,N_6179);
nor U6202 (N_6202,N_6052,N_6126);
or U6203 (N_6203,N_6091,N_6088);
or U6204 (N_6204,N_6133,N_6024);
and U6205 (N_6205,N_6144,N_6171);
nor U6206 (N_6206,N_6116,N_6027);
and U6207 (N_6207,N_6136,N_6031);
nand U6208 (N_6208,N_6077,N_6123);
and U6209 (N_6209,N_6109,N_6093);
nand U6210 (N_6210,N_6064,N_6142);
nor U6211 (N_6211,N_6197,N_6161);
and U6212 (N_6212,N_6021,N_6046);
nand U6213 (N_6213,N_6100,N_6134);
xor U6214 (N_6214,N_6048,N_6112);
and U6215 (N_6215,N_6043,N_6164);
nand U6216 (N_6216,N_6113,N_6135);
nand U6217 (N_6217,N_6045,N_6128);
and U6218 (N_6218,N_6009,N_6014);
or U6219 (N_6219,N_6106,N_6121);
and U6220 (N_6220,N_6033,N_6063);
nor U6221 (N_6221,N_6096,N_6075);
nand U6222 (N_6222,N_6102,N_6094);
nor U6223 (N_6223,N_6032,N_6087);
nand U6224 (N_6224,N_6019,N_6192);
nor U6225 (N_6225,N_6114,N_6074);
and U6226 (N_6226,N_6198,N_6049);
nand U6227 (N_6227,N_6071,N_6130);
and U6228 (N_6228,N_6017,N_6003);
nor U6229 (N_6229,N_6006,N_6040);
and U6230 (N_6230,N_6062,N_6129);
or U6231 (N_6231,N_6187,N_6067);
nor U6232 (N_6232,N_6007,N_6173);
nor U6233 (N_6233,N_6054,N_6150);
and U6234 (N_6234,N_6195,N_6018);
nor U6235 (N_6235,N_6181,N_6110);
or U6236 (N_6236,N_6176,N_6182);
nand U6237 (N_6237,N_6120,N_6042);
or U6238 (N_6238,N_6189,N_6131);
or U6239 (N_6239,N_6037,N_6188);
nand U6240 (N_6240,N_6023,N_6029);
nor U6241 (N_6241,N_6056,N_6084);
or U6242 (N_6242,N_6149,N_6175);
or U6243 (N_6243,N_6036,N_6039);
xnor U6244 (N_6244,N_6183,N_6082);
nor U6245 (N_6245,N_6068,N_6066);
nand U6246 (N_6246,N_6153,N_6119);
or U6247 (N_6247,N_6141,N_6107);
nand U6248 (N_6248,N_6165,N_6015);
or U6249 (N_6249,N_6061,N_6089);
or U6250 (N_6250,N_6000,N_6101);
nor U6251 (N_6251,N_6057,N_6050);
and U6252 (N_6252,N_6103,N_6085);
nand U6253 (N_6253,N_6163,N_6079);
nand U6254 (N_6254,N_6172,N_6041);
nor U6255 (N_6255,N_6156,N_6090);
or U6256 (N_6256,N_6080,N_6105);
nor U6257 (N_6257,N_6004,N_6022);
or U6258 (N_6258,N_6058,N_6122);
nor U6259 (N_6259,N_6073,N_6025);
and U6260 (N_6260,N_6132,N_6159);
nand U6261 (N_6261,N_6193,N_6104);
nor U6262 (N_6262,N_6035,N_6083);
nor U6263 (N_6263,N_6180,N_6047);
nand U6264 (N_6264,N_6154,N_6098);
or U6265 (N_6265,N_6166,N_6152);
or U6266 (N_6266,N_6169,N_6138);
nand U6267 (N_6267,N_6162,N_6034);
nor U6268 (N_6268,N_6012,N_6081);
nor U6269 (N_6269,N_6028,N_6196);
and U6270 (N_6270,N_6011,N_6118);
and U6271 (N_6271,N_6008,N_6139);
nor U6272 (N_6272,N_6117,N_6145);
or U6273 (N_6273,N_6070,N_6038);
nor U6274 (N_6274,N_6146,N_6055);
or U6275 (N_6275,N_6092,N_6095);
nor U6276 (N_6276,N_6026,N_6147);
nor U6277 (N_6277,N_6051,N_6137);
and U6278 (N_6278,N_6157,N_6072);
and U6279 (N_6279,N_6190,N_6151);
and U6280 (N_6280,N_6125,N_6191);
nand U6281 (N_6281,N_6097,N_6002);
and U6282 (N_6282,N_6010,N_6158);
or U6283 (N_6283,N_6167,N_6044);
and U6284 (N_6284,N_6155,N_6148);
nor U6285 (N_6285,N_6186,N_6199);
or U6286 (N_6286,N_6013,N_6086);
nor U6287 (N_6287,N_6170,N_6005);
and U6288 (N_6288,N_6078,N_6099);
and U6289 (N_6289,N_6127,N_6143);
and U6290 (N_6290,N_6184,N_6194);
and U6291 (N_6291,N_6053,N_6140);
nand U6292 (N_6292,N_6174,N_6115);
or U6293 (N_6293,N_6076,N_6160);
nand U6294 (N_6294,N_6069,N_6168);
or U6295 (N_6295,N_6059,N_6020);
nor U6296 (N_6296,N_6177,N_6108);
or U6297 (N_6297,N_6178,N_6185);
or U6298 (N_6298,N_6030,N_6060);
or U6299 (N_6299,N_6111,N_6065);
nand U6300 (N_6300,N_6058,N_6073);
and U6301 (N_6301,N_6191,N_6135);
nand U6302 (N_6302,N_6084,N_6088);
nand U6303 (N_6303,N_6160,N_6050);
nor U6304 (N_6304,N_6022,N_6185);
or U6305 (N_6305,N_6127,N_6110);
nand U6306 (N_6306,N_6006,N_6089);
nand U6307 (N_6307,N_6084,N_6150);
or U6308 (N_6308,N_6191,N_6042);
nor U6309 (N_6309,N_6016,N_6168);
and U6310 (N_6310,N_6136,N_6052);
nor U6311 (N_6311,N_6195,N_6181);
nor U6312 (N_6312,N_6055,N_6095);
nor U6313 (N_6313,N_6020,N_6084);
xnor U6314 (N_6314,N_6157,N_6087);
and U6315 (N_6315,N_6079,N_6090);
or U6316 (N_6316,N_6151,N_6034);
or U6317 (N_6317,N_6188,N_6121);
nor U6318 (N_6318,N_6175,N_6148);
or U6319 (N_6319,N_6098,N_6129);
or U6320 (N_6320,N_6118,N_6055);
nor U6321 (N_6321,N_6185,N_6091);
nand U6322 (N_6322,N_6061,N_6084);
nand U6323 (N_6323,N_6110,N_6000);
or U6324 (N_6324,N_6005,N_6138);
and U6325 (N_6325,N_6082,N_6012);
or U6326 (N_6326,N_6048,N_6142);
and U6327 (N_6327,N_6054,N_6013);
nor U6328 (N_6328,N_6010,N_6134);
and U6329 (N_6329,N_6049,N_6180);
and U6330 (N_6330,N_6172,N_6096);
xnor U6331 (N_6331,N_6048,N_6025);
and U6332 (N_6332,N_6110,N_6018);
xor U6333 (N_6333,N_6029,N_6063);
and U6334 (N_6334,N_6056,N_6107);
nand U6335 (N_6335,N_6160,N_6132);
nand U6336 (N_6336,N_6124,N_6015);
nor U6337 (N_6337,N_6083,N_6072);
nand U6338 (N_6338,N_6106,N_6147);
or U6339 (N_6339,N_6014,N_6006);
xor U6340 (N_6340,N_6194,N_6170);
nand U6341 (N_6341,N_6175,N_6106);
or U6342 (N_6342,N_6132,N_6038);
or U6343 (N_6343,N_6074,N_6031);
and U6344 (N_6344,N_6062,N_6159);
or U6345 (N_6345,N_6066,N_6029);
or U6346 (N_6346,N_6055,N_6187);
nand U6347 (N_6347,N_6045,N_6169);
nand U6348 (N_6348,N_6188,N_6080);
nor U6349 (N_6349,N_6152,N_6194);
nor U6350 (N_6350,N_6111,N_6076);
nor U6351 (N_6351,N_6187,N_6158);
and U6352 (N_6352,N_6118,N_6126);
and U6353 (N_6353,N_6122,N_6036);
and U6354 (N_6354,N_6171,N_6136);
and U6355 (N_6355,N_6107,N_6012);
nor U6356 (N_6356,N_6162,N_6176);
nor U6357 (N_6357,N_6103,N_6199);
or U6358 (N_6358,N_6182,N_6102);
nor U6359 (N_6359,N_6027,N_6052);
xor U6360 (N_6360,N_6108,N_6068);
or U6361 (N_6361,N_6113,N_6031);
nor U6362 (N_6362,N_6006,N_6047);
nor U6363 (N_6363,N_6134,N_6074);
or U6364 (N_6364,N_6058,N_6161);
nand U6365 (N_6365,N_6193,N_6041);
and U6366 (N_6366,N_6145,N_6128);
nand U6367 (N_6367,N_6015,N_6178);
nor U6368 (N_6368,N_6165,N_6138);
nand U6369 (N_6369,N_6199,N_6131);
and U6370 (N_6370,N_6082,N_6115);
or U6371 (N_6371,N_6170,N_6133);
or U6372 (N_6372,N_6167,N_6072);
or U6373 (N_6373,N_6049,N_6087);
nor U6374 (N_6374,N_6187,N_6175);
or U6375 (N_6375,N_6057,N_6074);
nor U6376 (N_6376,N_6157,N_6106);
and U6377 (N_6377,N_6087,N_6037);
nand U6378 (N_6378,N_6026,N_6040);
nor U6379 (N_6379,N_6119,N_6108);
nand U6380 (N_6380,N_6072,N_6123);
nand U6381 (N_6381,N_6045,N_6138);
and U6382 (N_6382,N_6166,N_6108);
and U6383 (N_6383,N_6138,N_6104);
and U6384 (N_6384,N_6026,N_6167);
xnor U6385 (N_6385,N_6033,N_6001);
nor U6386 (N_6386,N_6029,N_6007);
nand U6387 (N_6387,N_6182,N_6192);
nand U6388 (N_6388,N_6084,N_6157);
and U6389 (N_6389,N_6049,N_6189);
nor U6390 (N_6390,N_6167,N_6057);
or U6391 (N_6391,N_6149,N_6148);
nor U6392 (N_6392,N_6170,N_6125);
nor U6393 (N_6393,N_6179,N_6007);
and U6394 (N_6394,N_6139,N_6128);
nor U6395 (N_6395,N_6093,N_6007);
nor U6396 (N_6396,N_6185,N_6187);
or U6397 (N_6397,N_6194,N_6169);
and U6398 (N_6398,N_6165,N_6166);
and U6399 (N_6399,N_6099,N_6096);
nor U6400 (N_6400,N_6296,N_6310);
xnor U6401 (N_6401,N_6294,N_6297);
nand U6402 (N_6402,N_6312,N_6210);
nor U6403 (N_6403,N_6289,N_6309);
or U6404 (N_6404,N_6261,N_6337);
and U6405 (N_6405,N_6318,N_6230);
or U6406 (N_6406,N_6211,N_6320);
and U6407 (N_6407,N_6332,N_6399);
nand U6408 (N_6408,N_6398,N_6262);
or U6409 (N_6409,N_6253,N_6300);
nor U6410 (N_6410,N_6377,N_6287);
or U6411 (N_6411,N_6385,N_6393);
and U6412 (N_6412,N_6351,N_6246);
nand U6413 (N_6413,N_6223,N_6201);
and U6414 (N_6414,N_6389,N_6380);
nor U6415 (N_6415,N_6390,N_6254);
or U6416 (N_6416,N_6365,N_6267);
nand U6417 (N_6417,N_6364,N_6306);
or U6418 (N_6418,N_6238,N_6224);
and U6419 (N_6419,N_6383,N_6241);
nor U6420 (N_6420,N_6266,N_6301);
and U6421 (N_6421,N_6295,N_6208);
nor U6422 (N_6422,N_6329,N_6378);
or U6423 (N_6423,N_6379,N_6249);
nand U6424 (N_6424,N_6245,N_6353);
and U6425 (N_6425,N_6326,N_6299);
or U6426 (N_6426,N_6252,N_6273);
nor U6427 (N_6427,N_6319,N_6366);
nor U6428 (N_6428,N_6317,N_6363);
and U6429 (N_6429,N_6298,N_6316);
xnor U6430 (N_6430,N_6392,N_6214);
nand U6431 (N_6431,N_6235,N_6209);
and U6432 (N_6432,N_6282,N_6216);
and U6433 (N_6433,N_6331,N_6275);
or U6434 (N_6434,N_6362,N_6292);
or U6435 (N_6435,N_6341,N_6370);
or U6436 (N_6436,N_6369,N_6345);
nor U6437 (N_6437,N_6270,N_6397);
nand U6438 (N_6438,N_6325,N_6225);
and U6439 (N_6439,N_6330,N_6227);
nor U6440 (N_6440,N_6367,N_6202);
or U6441 (N_6441,N_6356,N_6229);
and U6442 (N_6442,N_6373,N_6286);
or U6443 (N_6443,N_6308,N_6217);
nand U6444 (N_6444,N_6347,N_6339);
and U6445 (N_6445,N_6268,N_6361);
nor U6446 (N_6446,N_6352,N_6234);
nand U6447 (N_6447,N_6260,N_6384);
or U6448 (N_6448,N_6307,N_6205);
and U6449 (N_6449,N_6204,N_6344);
nor U6450 (N_6450,N_6371,N_6396);
nand U6451 (N_6451,N_6338,N_6304);
and U6452 (N_6452,N_6281,N_6322);
or U6453 (N_6453,N_6265,N_6251);
xor U6454 (N_6454,N_6324,N_6239);
and U6455 (N_6455,N_6315,N_6313);
nand U6456 (N_6456,N_6323,N_6242);
nor U6457 (N_6457,N_6333,N_6382);
or U6458 (N_6458,N_6250,N_6368);
nor U6459 (N_6459,N_6231,N_6255);
and U6460 (N_6460,N_6271,N_6219);
nand U6461 (N_6461,N_6342,N_6256);
nand U6462 (N_6462,N_6206,N_6213);
nand U6463 (N_6463,N_6259,N_6293);
or U6464 (N_6464,N_6215,N_6305);
or U6465 (N_6465,N_6340,N_6276);
nand U6466 (N_6466,N_6355,N_6236);
nor U6467 (N_6467,N_6248,N_6376);
nor U6468 (N_6468,N_6334,N_6327);
or U6469 (N_6469,N_6228,N_6200);
nand U6470 (N_6470,N_6388,N_6328);
or U6471 (N_6471,N_6277,N_6391);
or U6472 (N_6472,N_6284,N_6358);
or U6473 (N_6473,N_6272,N_6274);
or U6474 (N_6474,N_6346,N_6243);
nand U6475 (N_6475,N_6220,N_6381);
or U6476 (N_6476,N_6386,N_6375);
and U6477 (N_6477,N_6343,N_6247);
or U6478 (N_6478,N_6240,N_6314);
and U6479 (N_6479,N_6218,N_6233);
nor U6480 (N_6480,N_6278,N_6232);
and U6481 (N_6481,N_6244,N_6237);
nand U6482 (N_6482,N_6264,N_6257);
and U6483 (N_6483,N_6203,N_6258);
nor U6484 (N_6484,N_6394,N_6279);
nand U6485 (N_6485,N_6349,N_6207);
nor U6486 (N_6486,N_6311,N_6336);
nand U6487 (N_6487,N_6222,N_6212);
nor U6488 (N_6488,N_6226,N_6285);
and U6489 (N_6489,N_6372,N_6302);
or U6490 (N_6490,N_6290,N_6283);
nor U6491 (N_6491,N_6335,N_6350);
or U6492 (N_6492,N_6303,N_6354);
xnor U6493 (N_6493,N_6360,N_6288);
and U6494 (N_6494,N_6263,N_6348);
nand U6495 (N_6495,N_6357,N_6387);
nand U6496 (N_6496,N_6280,N_6395);
or U6497 (N_6497,N_6221,N_6269);
or U6498 (N_6498,N_6321,N_6374);
and U6499 (N_6499,N_6359,N_6291);
and U6500 (N_6500,N_6361,N_6342);
nor U6501 (N_6501,N_6366,N_6298);
and U6502 (N_6502,N_6220,N_6339);
or U6503 (N_6503,N_6376,N_6226);
nand U6504 (N_6504,N_6282,N_6346);
or U6505 (N_6505,N_6273,N_6390);
nand U6506 (N_6506,N_6390,N_6335);
nor U6507 (N_6507,N_6257,N_6313);
and U6508 (N_6508,N_6283,N_6247);
and U6509 (N_6509,N_6264,N_6207);
or U6510 (N_6510,N_6348,N_6394);
nor U6511 (N_6511,N_6290,N_6214);
or U6512 (N_6512,N_6336,N_6215);
and U6513 (N_6513,N_6357,N_6350);
nand U6514 (N_6514,N_6335,N_6205);
nor U6515 (N_6515,N_6389,N_6272);
nand U6516 (N_6516,N_6248,N_6260);
nor U6517 (N_6517,N_6248,N_6308);
or U6518 (N_6518,N_6242,N_6387);
nand U6519 (N_6519,N_6298,N_6370);
and U6520 (N_6520,N_6353,N_6250);
nand U6521 (N_6521,N_6234,N_6210);
and U6522 (N_6522,N_6219,N_6233);
and U6523 (N_6523,N_6277,N_6398);
or U6524 (N_6524,N_6355,N_6222);
and U6525 (N_6525,N_6377,N_6262);
nor U6526 (N_6526,N_6319,N_6218);
nor U6527 (N_6527,N_6328,N_6282);
xor U6528 (N_6528,N_6387,N_6247);
nand U6529 (N_6529,N_6365,N_6362);
nor U6530 (N_6530,N_6359,N_6337);
and U6531 (N_6531,N_6369,N_6273);
nor U6532 (N_6532,N_6359,N_6299);
or U6533 (N_6533,N_6344,N_6319);
nand U6534 (N_6534,N_6298,N_6331);
nor U6535 (N_6535,N_6255,N_6357);
nand U6536 (N_6536,N_6343,N_6221);
nor U6537 (N_6537,N_6208,N_6213);
and U6538 (N_6538,N_6225,N_6322);
nand U6539 (N_6539,N_6285,N_6296);
nand U6540 (N_6540,N_6297,N_6338);
nor U6541 (N_6541,N_6230,N_6234);
nand U6542 (N_6542,N_6228,N_6256);
or U6543 (N_6543,N_6356,N_6305);
nor U6544 (N_6544,N_6316,N_6349);
and U6545 (N_6545,N_6348,N_6283);
nand U6546 (N_6546,N_6267,N_6399);
nand U6547 (N_6547,N_6215,N_6367);
and U6548 (N_6548,N_6386,N_6235);
nand U6549 (N_6549,N_6390,N_6271);
nor U6550 (N_6550,N_6301,N_6231);
nor U6551 (N_6551,N_6318,N_6396);
nand U6552 (N_6552,N_6382,N_6367);
or U6553 (N_6553,N_6378,N_6382);
nand U6554 (N_6554,N_6318,N_6312);
nor U6555 (N_6555,N_6371,N_6202);
or U6556 (N_6556,N_6255,N_6342);
nor U6557 (N_6557,N_6264,N_6334);
nand U6558 (N_6558,N_6245,N_6320);
nand U6559 (N_6559,N_6259,N_6372);
or U6560 (N_6560,N_6206,N_6220);
or U6561 (N_6561,N_6207,N_6259);
nor U6562 (N_6562,N_6208,N_6315);
and U6563 (N_6563,N_6365,N_6317);
nor U6564 (N_6564,N_6241,N_6294);
nor U6565 (N_6565,N_6215,N_6313);
xor U6566 (N_6566,N_6254,N_6305);
nand U6567 (N_6567,N_6286,N_6328);
nand U6568 (N_6568,N_6242,N_6248);
nand U6569 (N_6569,N_6232,N_6227);
nand U6570 (N_6570,N_6267,N_6206);
nor U6571 (N_6571,N_6218,N_6308);
nor U6572 (N_6572,N_6228,N_6378);
or U6573 (N_6573,N_6244,N_6352);
nand U6574 (N_6574,N_6395,N_6372);
nand U6575 (N_6575,N_6242,N_6328);
or U6576 (N_6576,N_6392,N_6241);
and U6577 (N_6577,N_6236,N_6365);
or U6578 (N_6578,N_6318,N_6334);
or U6579 (N_6579,N_6327,N_6204);
nor U6580 (N_6580,N_6207,N_6360);
or U6581 (N_6581,N_6338,N_6323);
and U6582 (N_6582,N_6389,N_6371);
nor U6583 (N_6583,N_6303,N_6310);
or U6584 (N_6584,N_6377,N_6382);
or U6585 (N_6585,N_6237,N_6247);
nor U6586 (N_6586,N_6242,N_6206);
nor U6587 (N_6587,N_6289,N_6319);
and U6588 (N_6588,N_6327,N_6396);
nand U6589 (N_6589,N_6230,N_6358);
or U6590 (N_6590,N_6239,N_6340);
or U6591 (N_6591,N_6206,N_6321);
or U6592 (N_6592,N_6389,N_6329);
nand U6593 (N_6593,N_6265,N_6327);
nand U6594 (N_6594,N_6249,N_6283);
or U6595 (N_6595,N_6285,N_6307);
xnor U6596 (N_6596,N_6242,N_6357);
nand U6597 (N_6597,N_6268,N_6390);
nor U6598 (N_6598,N_6320,N_6264);
nand U6599 (N_6599,N_6327,N_6222);
nor U6600 (N_6600,N_6426,N_6521);
nor U6601 (N_6601,N_6492,N_6496);
nor U6602 (N_6602,N_6558,N_6550);
or U6603 (N_6603,N_6402,N_6522);
or U6604 (N_6604,N_6452,N_6578);
or U6605 (N_6605,N_6527,N_6571);
nand U6606 (N_6606,N_6579,N_6546);
nand U6607 (N_6607,N_6548,N_6432);
and U6608 (N_6608,N_6598,N_6480);
or U6609 (N_6609,N_6505,N_6560);
or U6610 (N_6610,N_6435,N_6586);
nor U6611 (N_6611,N_6420,N_6563);
and U6612 (N_6612,N_6434,N_6436);
xor U6613 (N_6613,N_6516,N_6576);
nand U6614 (N_6614,N_6543,N_6449);
nor U6615 (N_6615,N_6499,N_6568);
and U6616 (N_6616,N_6493,N_6468);
xor U6617 (N_6617,N_6472,N_6534);
and U6618 (N_6618,N_6514,N_6556);
or U6619 (N_6619,N_6474,N_6554);
and U6620 (N_6620,N_6573,N_6559);
or U6621 (N_6621,N_6495,N_6528);
nand U6622 (N_6622,N_6484,N_6589);
and U6623 (N_6623,N_6450,N_6411);
nor U6624 (N_6624,N_6539,N_6460);
nor U6625 (N_6625,N_6570,N_6467);
or U6626 (N_6626,N_6588,N_6557);
or U6627 (N_6627,N_6425,N_6567);
and U6628 (N_6628,N_6476,N_6544);
and U6629 (N_6629,N_6575,N_6400);
nand U6630 (N_6630,N_6442,N_6502);
or U6631 (N_6631,N_6405,N_6465);
nand U6632 (N_6632,N_6423,N_6433);
nor U6633 (N_6633,N_6403,N_6424);
nor U6634 (N_6634,N_6591,N_6574);
nor U6635 (N_6635,N_6459,N_6566);
and U6636 (N_6636,N_6483,N_6469);
and U6637 (N_6637,N_6585,N_6594);
nor U6638 (N_6638,N_6438,N_6498);
nand U6639 (N_6639,N_6491,N_6583);
or U6640 (N_6640,N_6526,N_6512);
or U6641 (N_6641,N_6440,N_6551);
and U6642 (N_6642,N_6475,N_6487);
and U6643 (N_6643,N_6552,N_6580);
or U6644 (N_6644,N_6482,N_6596);
nor U6645 (N_6645,N_6533,N_6525);
nand U6646 (N_6646,N_6553,N_6451);
nor U6647 (N_6647,N_6429,N_6523);
or U6648 (N_6648,N_6538,N_6455);
nand U6649 (N_6649,N_6417,N_6503);
nand U6650 (N_6650,N_6584,N_6509);
and U6651 (N_6651,N_6457,N_6444);
xor U6652 (N_6652,N_6414,N_6581);
or U6653 (N_6653,N_6443,N_6413);
and U6654 (N_6654,N_6416,N_6464);
or U6655 (N_6655,N_6564,N_6510);
nor U6656 (N_6656,N_6478,N_6486);
or U6657 (N_6657,N_6448,N_6587);
nor U6658 (N_6658,N_6439,N_6595);
nand U6659 (N_6659,N_6406,N_6508);
nand U6660 (N_6660,N_6485,N_6407);
and U6661 (N_6661,N_6542,N_6463);
nor U6662 (N_6662,N_6410,N_6456);
nor U6663 (N_6663,N_6497,N_6428);
or U6664 (N_6664,N_6561,N_6519);
or U6665 (N_6665,N_6536,N_6592);
and U6666 (N_6666,N_6565,N_6488);
nand U6667 (N_6667,N_6430,N_6507);
nand U6668 (N_6668,N_6530,N_6513);
nand U6669 (N_6669,N_6415,N_6408);
and U6670 (N_6670,N_6494,N_6477);
or U6671 (N_6671,N_6453,N_6532);
nand U6672 (N_6672,N_6540,N_6471);
or U6673 (N_6673,N_6599,N_6412);
xnor U6674 (N_6674,N_6517,N_6582);
nand U6675 (N_6675,N_6419,N_6489);
and U6676 (N_6676,N_6404,N_6555);
nand U6677 (N_6677,N_6501,N_6431);
and U6678 (N_6678,N_6506,N_6545);
nor U6679 (N_6679,N_6421,N_6597);
nand U6680 (N_6680,N_6593,N_6473);
nor U6681 (N_6681,N_6445,N_6504);
and U6682 (N_6682,N_6535,N_6515);
nand U6683 (N_6683,N_6490,N_6470);
nor U6684 (N_6684,N_6458,N_6447);
and U6685 (N_6685,N_6549,N_6562);
and U6686 (N_6686,N_6524,N_6590);
and U6687 (N_6687,N_6437,N_6418);
and U6688 (N_6688,N_6441,N_6461);
or U6689 (N_6689,N_6541,N_6401);
or U6690 (N_6690,N_6518,N_6466);
and U6691 (N_6691,N_6547,N_6462);
or U6692 (N_6692,N_6537,N_6446);
or U6693 (N_6693,N_6511,N_6454);
or U6694 (N_6694,N_6422,N_6520);
or U6695 (N_6695,N_6569,N_6500);
or U6696 (N_6696,N_6481,N_6577);
nand U6697 (N_6697,N_6529,N_6427);
and U6698 (N_6698,N_6572,N_6409);
or U6699 (N_6699,N_6531,N_6479);
or U6700 (N_6700,N_6404,N_6577);
or U6701 (N_6701,N_6512,N_6470);
and U6702 (N_6702,N_6543,N_6434);
or U6703 (N_6703,N_6481,N_6579);
nor U6704 (N_6704,N_6546,N_6446);
nor U6705 (N_6705,N_6474,N_6518);
or U6706 (N_6706,N_6578,N_6457);
nand U6707 (N_6707,N_6527,N_6448);
and U6708 (N_6708,N_6485,N_6538);
nor U6709 (N_6709,N_6565,N_6490);
nand U6710 (N_6710,N_6417,N_6544);
nor U6711 (N_6711,N_6542,N_6404);
and U6712 (N_6712,N_6554,N_6432);
nand U6713 (N_6713,N_6543,N_6529);
nand U6714 (N_6714,N_6492,N_6591);
nand U6715 (N_6715,N_6442,N_6407);
or U6716 (N_6716,N_6482,N_6479);
nor U6717 (N_6717,N_6485,N_6563);
or U6718 (N_6718,N_6548,N_6525);
and U6719 (N_6719,N_6556,N_6407);
and U6720 (N_6720,N_6581,N_6456);
and U6721 (N_6721,N_6592,N_6576);
or U6722 (N_6722,N_6576,N_6430);
nor U6723 (N_6723,N_6520,N_6487);
nor U6724 (N_6724,N_6581,N_6593);
or U6725 (N_6725,N_6581,N_6513);
and U6726 (N_6726,N_6589,N_6451);
and U6727 (N_6727,N_6520,N_6564);
nor U6728 (N_6728,N_6531,N_6409);
or U6729 (N_6729,N_6589,N_6463);
and U6730 (N_6730,N_6421,N_6550);
nand U6731 (N_6731,N_6450,N_6553);
nand U6732 (N_6732,N_6596,N_6461);
and U6733 (N_6733,N_6440,N_6479);
or U6734 (N_6734,N_6465,N_6404);
nand U6735 (N_6735,N_6489,N_6425);
or U6736 (N_6736,N_6545,N_6548);
and U6737 (N_6737,N_6418,N_6511);
nor U6738 (N_6738,N_6502,N_6448);
or U6739 (N_6739,N_6591,N_6565);
nand U6740 (N_6740,N_6463,N_6592);
and U6741 (N_6741,N_6419,N_6596);
or U6742 (N_6742,N_6514,N_6518);
and U6743 (N_6743,N_6425,N_6599);
nor U6744 (N_6744,N_6409,N_6481);
nand U6745 (N_6745,N_6496,N_6512);
nand U6746 (N_6746,N_6598,N_6419);
or U6747 (N_6747,N_6499,N_6541);
or U6748 (N_6748,N_6501,N_6566);
and U6749 (N_6749,N_6435,N_6517);
or U6750 (N_6750,N_6458,N_6408);
or U6751 (N_6751,N_6444,N_6560);
or U6752 (N_6752,N_6588,N_6429);
nor U6753 (N_6753,N_6576,N_6535);
nor U6754 (N_6754,N_6477,N_6526);
nor U6755 (N_6755,N_6477,N_6530);
or U6756 (N_6756,N_6437,N_6527);
nor U6757 (N_6757,N_6526,N_6568);
and U6758 (N_6758,N_6421,N_6590);
and U6759 (N_6759,N_6451,N_6409);
nand U6760 (N_6760,N_6431,N_6404);
nor U6761 (N_6761,N_6471,N_6407);
nor U6762 (N_6762,N_6558,N_6581);
or U6763 (N_6763,N_6532,N_6490);
nor U6764 (N_6764,N_6563,N_6533);
or U6765 (N_6765,N_6531,N_6592);
nor U6766 (N_6766,N_6531,N_6590);
or U6767 (N_6767,N_6509,N_6537);
nor U6768 (N_6768,N_6487,N_6499);
and U6769 (N_6769,N_6596,N_6577);
nor U6770 (N_6770,N_6509,N_6494);
nor U6771 (N_6771,N_6512,N_6505);
or U6772 (N_6772,N_6413,N_6400);
nand U6773 (N_6773,N_6423,N_6560);
and U6774 (N_6774,N_6565,N_6439);
or U6775 (N_6775,N_6565,N_6433);
nor U6776 (N_6776,N_6410,N_6469);
nand U6777 (N_6777,N_6571,N_6591);
and U6778 (N_6778,N_6522,N_6592);
nand U6779 (N_6779,N_6531,N_6447);
and U6780 (N_6780,N_6589,N_6565);
and U6781 (N_6781,N_6411,N_6525);
and U6782 (N_6782,N_6539,N_6475);
nor U6783 (N_6783,N_6578,N_6479);
nand U6784 (N_6784,N_6580,N_6426);
nor U6785 (N_6785,N_6443,N_6455);
nor U6786 (N_6786,N_6584,N_6544);
or U6787 (N_6787,N_6481,N_6594);
or U6788 (N_6788,N_6595,N_6404);
nor U6789 (N_6789,N_6489,N_6511);
or U6790 (N_6790,N_6546,N_6492);
nor U6791 (N_6791,N_6557,N_6450);
and U6792 (N_6792,N_6502,N_6581);
and U6793 (N_6793,N_6409,N_6401);
and U6794 (N_6794,N_6546,N_6404);
nand U6795 (N_6795,N_6592,N_6406);
nor U6796 (N_6796,N_6568,N_6446);
or U6797 (N_6797,N_6509,N_6483);
and U6798 (N_6798,N_6447,N_6413);
or U6799 (N_6799,N_6461,N_6509);
or U6800 (N_6800,N_6732,N_6778);
nor U6801 (N_6801,N_6722,N_6715);
nor U6802 (N_6802,N_6701,N_6608);
nor U6803 (N_6803,N_6746,N_6748);
nand U6804 (N_6804,N_6643,N_6607);
or U6805 (N_6805,N_6777,N_6648);
xor U6806 (N_6806,N_6791,N_6736);
or U6807 (N_6807,N_6633,N_6689);
xnor U6808 (N_6808,N_6794,N_6642);
and U6809 (N_6809,N_6638,N_6729);
nor U6810 (N_6810,N_6668,N_6693);
nor U6811 (N_6811,N_6750,N_6757);
and U6812 (N_6812,N_6711,N_6710);
and U6813 (N_6813,N_6658,N_6627);
or U6814 (N_6814,N_6673,N_6762);
nand U6815 (N_6815,N_6790,N_6730);
or U6816 (N_6816,N_6703,N_6604);
nand U6817 (N_6817,N_6612,N_6725);
or U6818 (N_6818,N_6665,N_6626);
or U6819 (N_6819,N_6610,N_6797);
or U6820 (N_6820,N_6600,N_6744);
and U6821 (N_6821,N_6619,N_6760);
or U6822 (N_6822,N_6796,N_6766);
nor U6823 (N_6823,N_6664,N_6678);
or U6824 (N_6824,N_6763,N_6754);
nor U6825 (N_6825,N_6647,N_6646);
nor U6826 (N_6826,N_6683,N_6785);
and U6827 (N_6827,N_6764,N_6702);
nor U6828 (N_6828,N_6654,N_6759);
nand U6829 (N_6829,N_6623,N_6779);
nand U6830 (N_6830,N_6603,N_6685);
and U6831 (N_6831,N_6625,N_6798);
or U6832 (N_6832,N_6752,N_6696);
nand U6833 (N_6833,N_6650,N_6672);
and U6834 (N_6834,N_6629,N_6712);
and U6835 (N_6835,N_6720,N_6691);
or U6836 (N_6836,N_6774,N_6613);
or U6837 (N_6837,N_6709,N_6758);
or U6838 (N_6838,N_6700,N_6768);
nor U6839 (N_6839,N_6679,N_6721);
nor U6840 (N_6840,N_6639,N_6780);
or U6841 (N_6841,N_6783,N_6751);
or U6842 (N_6842,N_6765,N_6697);
or U6843 (N_6843,N_6649,N_6659);
and U6844 (N_6844,N_6753,N_6770);
nor U6845 (N_6845,N_6792,N_6793);
or U6846 (N_6846,N_6769,N_6747);
and U6847 (N_6847,N_6724,N_6788);
or U6848 (N_6848,N_6742,N_6628);
nand U6849 (N_6849,N_6740,N_6695);
or U6850 (N_6850,N_6781,N_6726);
nand U6851 (N_6851,N_6674,N_6728);
xor U6852 (N_6852,N_6745,N_6741);
xnor U6853 (N_6853,N_6630,N_6611);
and U6854 (N_6854,N_6690,N_6718);
and U6855 (N_6855,N_6615,N_6714);
and U6856 (N_6856,N_6743,N_6621);
and U6857 (N_6857,N_6707,N_6620);
nor U6858 (N_6858,N_6635,N_6622);
or U6859 (N_6859,N_6789,N_6708);
or U6860 (N_6860,N_6716,N_6776);
nor U6861 (N_6861,N_6755,N_6737);
and U6862 (N_6862,N_6680,N_6739);
or U6863 (N_6863,N_6636,N_6631);
and U6864 (N_6864,N_6699,N_6661);
or U6865 (N_6865,N_6634,N_6662);
and U6866 (N_6866,N_6681,N_6601);
or U6867 (N_6867,N_6795,N_6651);
nand U6868 (N_6868,N_6706,N_6655);
xnor U6869 (N_6869,N_6773,N_6660);
or U6870 (N_6870,N_6767,N_6645);
xnor U6871 (N_6871,N_6644,N_6675);
nor U6872 (N_6872,N_6713,N_6676);
and U6873 (N_6873,N_6670,N_6671);
nand U6874 (N_6874,N_6684,N_6775);
or U6875 (N_6875,N_6688,N_6749);
nand U6876 (N_6876,N_6632,N_6733);
nand U6877 (N_6877,N_6799,N_6605);
nand U6878 (N_6878,N_6669,N_6641);
and U6879 (N_6879,N_6652,N_6772);
nor U6880 (N_6880,N_6771,N_6687);
and U6881 (N_6881,N_6787,N_6738);
xor U6882 (N_6882,N_6698,N_6734);
or U6883 (N_6883,N_6602,N_6618);
nand U6884 (N_6884,N_6606,N_6653);
and U6885 (N_6885,N_6784,N_6666);
and U6886 (N_6886,N_6692,N_6616);
nor U6887 (N_6887,N_6682,N_6731);
and U6888 (N_6888,N_6723,N_6704);
and U6889 (N_6889,N_6735,N_6761);
and U6890 (N_6890,N_6640,N_6656);
and U6891 (N_6891,N_6782,N_6756);
or U6892 (N_6892,N_6694,N_6717);
xnor U6893 (N_6893,N_6614,N_6677);
nor U6894 (N_6894,N_6609,N_6686);
xnor U6895 (N_6895,N_6617,N_6786);
nor U6896 (N_6896,N_6667,N_6719);
nor U6897 (N_6897,N_6727,N_6705);
nand U6898 (N_6898,N_6637,N_6663);
and U6899 (N_6899,N_6657,N_6624);
or U6900 (N_6900,N_6738,N_6690);
nand U6901 (N_6901,N_6708,N_6688);
or U6902 (N_6902,N_6759,N_6718);
and U6903 (N_6903,N_6778,N_6683);
and U6904 (N_6904,N_6666,N_6704);
and U6905 (N_6905,N_6697,N_6687);
nor U6906 (N_6906,N_6748,N_6794);
and U6907 (N_6907,N_6753,N_6680);
nor U6908 (N_6908,N_6751,N_6726);
or U6909 (N_6909,N_6628,N_6763);
or U6910 (N_6910,N_6762,N_6613);
or U6911 (N_6911,N_6643,N_6743);
and U6912 (N_6912,N_6729,N_6797);
and U6913 (N_6913,N_6685,N_6691);
xnor U6914 (N_6914,N_6637,N_6696);
or U6915 (N_6915,N_6606,N_6761);
and U6916 (N_6916,N_6738,N_6759);
nand U6917 (N_6917,N_6645,N_6763);
nor U6918 (N_6918,N_6670,N_6730);
and U6919 (N_6919,N_6737,N_6663);
nand U6920 (N_6920,N_6651,N_6796);
and U6921 (N_6921,N_6682,N_6671);
and U6922 (N_6922,N_6766,N_6650);
nand U6923 (N_6923,N_6725,N_6667);
nor U6924 (N_6924,N_6638,N_6751);
nand U6925 (N_6925,N_6715,N_6619);
nor U6926 (N_6926,N_6673,N_6672);
or U6927 (N_6927,N_6753,N_6708);
or U6928 (N_6928,N_6795,N_6738);
and U6929 (N_6929,N_6798,N_6765);
nand U6930 (N_6930,N_6678,N_6681);
xor U6931 (N_6931,N_6797,N_6665);
nor U6932 (N_6932,N_6709,N_6644);
nor U6933 (N_6933,N_6760,N_6737);
or U6934 (N_6934,N_6670,N_6776);
nor U6935 (N_6935,N_6684,N_6620);
nand U6936 (N_6936,N_6635,N_6614);
and U6937 (N_6937,N_6644,N_6622);
nand U6938 (N_6938,N_6727,N_6691);
and U6939 (N_6939,N_6768,N_6772);
and U6940 (N_6940,N_6737,N_6784);
or U6941 (N_6941,N_6720,N_6779);
nor U6942 (N_6942,N_6794,N_6746);
and U6943 (N_6943,N_6738,N_6680);
and U6944 (N_6944,N_6794,N_6768);
and U6945 (N_6945,N_6642,N_6709);
and U6946 (N_6946,N_6706,N_6645);
and U6947 (N_6947,N_6662,N_6732);
and U6948 (N_6948,N_6714,N_6762);
nand U6949 (N_6949,N_6799,N_6747);
nor U6950 (N_6950,N_6794,N_6711);
and U6951 (N_6951,N_6603,N_6792);
nor U6952 (N_6952,N_6723,N_6646);
and U6953 (N_6953,N_6741,N_6608);
or U6954 (N_6954,N_6757,N_6706);
nand U6955 (N_6955,N_6730,N_6792);
nor U6956 (N_6956,N_6756,N_6649);
and U6957 (N_6957,N_6700,N_6612);
and U6958 (N_6958,N_6796,N_6627);
nand U6959 (N_6959,N_6716,N_6740);
or U6960 (N_6960,N_6729,N_6607);
nand U6961 (N_6961,N_6778,N_6613);
nand U6962 (N_6962,N_6636,N_6635);
and U6963 (N_6963,N_6674,N_6798);
nand U6964 (N_6964,N_6736,N_6641);
nor U6965 (N_6965,N_6799,N_6609);
nor U6966 (N_6966,N_6695,N_6630);
and U6967 (N_6967,N_6652,N_6663);
nor U6968 (N_6968,N_6727,N_6750);
nand U6969 (N_6969,N_6679,N_6740);
nor U6970 (N_6970,N_6714,N_6617);
and U6971 (N_6971,N_6702,N_6751);
or U6972 (N_6972,N_6648,N_6634);
nor U6973 (N_6973,N_6696,N_6615);
and U6974 (N_6974,N_6625,N_6709);
or U6975 (N_6975,N_6790,N_6784);
nand U6976 (N_6976,N_6747,N_6627);
nand U6977 (N_6977,N_6776,N_6799);
nor U6978 (N_6978,N_6789,N_6717);
and U6979 (N_6979,N_6662,N_6624);
and U6980 (N_6980,N_6642,N_6748);
and U6981 (N_6981,N_6618,N_6715);
nand U6982 (N_6982,N_6614,N_6784);
and U6983 (N_6983,N_6730,N_6706);
or U6984 (N_6984,N_6634,N_6600);
and U6985 (N_6985,N_6644,N_6751);
or U6986 (N_6986,N_6677,N_6675);
or U6987 (N_6987,N_6795,N_6697);
nor U6988 (N_6988,N_6698,N_6755);
nand U6989 (N_6989,N_6641,N_6771);
or U6990 (N_6990,N_6681,N_6690);
or U6991 (N_6991,N_6691,N_6629);
nor U6992 (N_6992,N_6682,N_6677);
nand U6993 (N_6993,N_6615,N_6787);
or U6994 (N_6994,N_6749,N_6721);
xor U6995 (N_6995,N_6673,N_6600);
and U6996 (N_6996,N_6697,N_6626);
or U6997 (N_6997,N_6641,N_6790);
nor U6998 (N_6998,N_6685,N_6736);
nor U6999 (N_6999,N_6758,N_6796);
nor U7000 (N_7000,N_6884,N_6994);
nand U7001 (N_7001,N_6982,N_6870);
nand U7002 (N_7002,N_6991,N_6907);
nor U7003 (N_7003,N_6826,N_6865);
nor U7004 (N_7004,N_6872,N_6952);
nor U7005 (N_7005,N_6959,N_6802);
or U7006 (N_7006,N_6891,N_6823);
nand U7007 (N_7007,N_6873,N_6833);
or U7008 (N_7008,N_6938,N_6875);
nor U7009 (N_7009,N_6964,N_6941);
nand U7010 (N_7010,N_6898,N_6830);
or U7011 (N_7011,N_6852,N_6888);
or U7012 (N_7012,N_6990,N_6837);
nor U7013 (N_7013,N_6935,N_6943);
nand U7014 (N_7014,N_6804,N_6809);
xor U7015 (N_7015,N_6945,N_6912);
nor U7016 (N_7016,N_6831,N_6933);
and U7017 (N_7017,N_6874,N_6810);
nor U7018 (N_7018,N_6866,N_6842);
nor U7019 (N_7019,N_6855,N_6817);
and U7020 (N_7020,N_6954,N_6993);
nand U7021 (N_7021,N_6909,N_6868);
xnor U7022 (N_7022,N_6905,N_6906);
nand U7023 (N_7023,N_6886,N_6829);
and U7024 (N_7024,N_6895,N_6820);
nand U7025 (N_7025,N_6960,N_6998);
nand U7026 (N_7026,N_6983,N_6913);
and U7027 (N_7027,N_6858,N_6996);
nand U7028 (N_7028,N_6966,N_6924);
and U7029 (N_7029,N_6890,N_6972);
and U7030 (N_7030,N_6897,N_6834);
and U7031 (N_7031,N_6963,N_6977);
and U7032 (N_7032,N_6989,N_6818);
or U7033 (N_7033,N_6976,N_6944);
nand U7034 (N_7034,N_6930,N_6808);
nor U7035 (N_7035,N_6979,N_6995);
or U7036 (N_7036,N_6928,N_6961);
nand U7037 (N_7037,N_6971,N_6997);
nor U7038 (N_7038,N_6860,N_6851);
nor U7039 (N_7039,N_6840,N_6848);
and U7040 (N_7040,N_6816,N_6919);
xor U7041 (N_7041,N_6850,N_6958);
and U7042 (N_7042,N_6942,N_6968);
nor U7043 (N_7043,N_6927,N_6992);
xor U7044 (N_7044,N_6864,N_6969);
nor U7045 (N_7045,N_6974,N_6843);
nor U7046 (N_7046,N_6880,N_6846);
and U7047 (N_7047,N_6955,N_6832);
nand U7048 (N_7048,N_6814,N_6970);
nor U7049 (N_7049,N_6853,N_6915);
nor U7050 (N_7050,N_6800,N_6908);
nand U7051 (N_7051,N_6867,N_6980);
and U7052 (N_7052,N_6937,N_6836);
nor U7053 (N_7053,N_6896,N_6967);
nor U7054 (N_7054,N_6981,N_6835);
or U7055 (N_7055,N_6861,N_6920);
nand U7056 (N_7056,N_6921,N_6871);
or U7057 (N_7057,N_6819,N_6940);
nand U7058 (N_7058,N_6910,N_6984);
nor U7059 (N_7059,N_6887,N_6929);
or U7060 (N_7060,N_6885,N_6988);
or U7061 (N_7061,N_6917,N_6881);
or U7062 (N_7062,N_6939,N_6923);
nor U7063 (N_7063,N_6893,N_6877);
nand U7064 (N_7064,N_6911,N_6918);
nand U7065 (N_7065,N_6805,N_6806);
nor U7066 (N_7066,N_6838,N_6953);
or U7067 (N_7067,N_6841,N_6932);
nand U7068 (N_7068,N_6985,N_6856);
nor U7069 (N_7069,N_6822,N_6812);
or U7070 (N_7070,N_6825,N_6878);
or U7071 (N_7071,N_6849,N_6889);
and U7072 (N_7072,N_6899,N_6987);
nor U7073 (N_7073,N_6902,N_6882);
nor U7074 (N_7074,N_6815,N_6916);
nor U7075 (N_7075,N_6859,N_6892);
nor U7076 (N_7076,N_6844,N_6801);
and U7077 (N_7077,N_6973,N_6862);
nor U7078 (N_7078,N_6965,N_6956);
or U7079 (N_7079,N_6962,N_6951);
and U7080 (N_7080,N_6946,N_6957);
nor U7081 (N_7081,N_6936,N_6869);
nand U7082 (N_7082,N_6978,N_6900);
nor U7083 (N_7083,N_6807,N_6845);
or U7084 (N_7084,N_6854,N_6925);
nand U7085 (N_7085,N_6821,N_6999);
and U7086 (N_7086,N_6883,N_6811);
nor U7087 (N_7087,N_6828,N_6894);
or U7088 (N_7088,N_6975,N_6824);
and U7089 (N_7089,N_6926,N_6847);
nor U7090 (N_7090,N_6931,N_6803);
or U7091 (N_7091,N_6949,N_6813);
and U7092 (N_7092,N_6922,N_6863);
nor U7093 (N_7093,N_6857,N_6986);
nand U7094 (N_7094,N_6827,N_6901);
nor U7095 (N_7095,N_6839,N_6934);
nand U7096 (N_7096,N_6879,N_6950);
nor U7097 (N_7097,N_6947,N_6904);
and U7098 (N_7098,N_6948,N_6876);
nand U7099 (N_7099,N_6903,N_6914);
nand U7100 (N_7100,N_6866,N_6917);
and U7101 (N_7101,N_6850,N_6982);
or U7102 (N_7102,N_6922,N_6951);
xnor U7103 (N_7103,N_6813,N_6969);
or U7104 (N_7104,N_6992,N_6852);
or U7105 (N_7105,N_6813,N_6927);
nand U7106 (N_7106,N_6864,N_6982);
nor U7107 (N_7107,N_6932,N_6858);
nor U7108 (N_7108,N_6844,N_6921);
and U7109 (N_7109,N_6815,N_6810);
and U7110 (N_7110,N_6993,N_6887);
and U7111 (N_7111,N_6918,N_6821);
or U7112 (N_7112,N_6842,N_6966);
and U7113 (N_7113,N_6930,N_6836);
and U7114 (N_7114,N_6875,N_6922);
and U7115 (N_7115,N_6900,N_6912);
or U7116 (N_7116,N_6880,N_6834);
and U7117 (N_7117,N_6914,N_6848);
xor U7118 (N_7118,N_6971,N_6890);
and U7119 (N_7119,N_6845,N_6852);
or U7120 (N_7120,N_6983,N_6903);
and U7121 (N_7121,N_6950,N_6909);
or U7122 (N_7122,N_6876,N_6871);
or U7123 (N_7123,N_6931,N_6893);
nor U7124 (N_7124,N_6957,N_6840);
and U7125 (N_7125,N_6960,N_6945);
or U7126 (N_7126,N_6823,N_6870);
and U7127 (N_7127,N_6826,N_6972);
or U7128 (N_7128,N_6884,N_6974);
and U7129 (N_7129,N_6886,N_6812);
and U7130 (N_7130,N_6843,N_6980);
nand U7131 (N_7131,N_6951,N_6865);
nand U7132 (N_7132,N_6878,N_6812);
nor U7133 (N_7133,N_6854,N_6810);
nand U7134 (N_7134,N_6945,N_6894);
nand U7135 (N_7135,N_6846,N_6830);
and U7136 (N_7136,N_6948,N_6968);
or U7137 (N_7137,N_6827,N_6807);
nand U7138 (N_7138,N_6946,N_6813);
and U7139 (N_7139,N_6823,N_6845);
or U7140 (N_7140,N_6996,N_6862);
and U7141 (N_7141,N_6981,N_6852);
nor U7142 (N_7142,N_6855,N_6882);
nand U7143 (N_7143,N_6947,N_6873);
nand U7144 (N_7144,N_6889,N_6958);
nand U7145 (N_7145,N_6935,N_6829);
nor U7146 (N_7146,N_6862,N_6848);
nor U7147 (N_7147,N_6851,N_6957);
nor U7148 (N_7148,N_6875,N_6941);
nand U7149 (N_7149,N_6869,N_6868);
and U7150 (N_7150,N_6851,N_6984);
and U7151 (N_7151,N_6810,N_6975);
nand U7152 (N_7152,N_6983,N_6855);
nor U7153 (N_7153,N_6865,N_6971);
nor U7154 (N_7154,N_6922,N_6952);
nor U7155 (N_7155,N_6999,N_6857);
and U7156 (N_7156,N_6957,N_6806);
nor U7157 (N_7157,N_6800,N_6933);
nor U7158 (N_7158,N_6882,N_6910);
and U7159 (N_7159,N_6803,N_6893);
or U7160 (N_7160,N_6987,N_6813);
and U7161 (N_7161,N_6899,N_6989);
nor U7162 (N_7162,N_6994,N_6829);
nor U7163 (N_7163,N_6846,N_6822);
or U7164 (N_7164,N_6888,N_6971);
or U7165 (N_7165,N_6975,N_6985);
or U7166 (N_7166,N_6919,N_6923);
nand U7167 (N_7167,N_6810,N_6951);
nand U7168 (N_7168,N_6835,N_6806);
or U7169 (N_7169,N_6952,N_6951);
or U7170 (N_7170,N_6875,N_6807);
nor U7171 (N_7171,N_6972,N_6840);
nand U7172 (N_7172,N_6954,N_6955);
and U7173 (N_7173,N_6814,N_6903);
and U7174 (N_7174,N_6965,N_6842);
or U7175 (N_7175,N_6898,N_6952);
and U7176 (N_7176,N_6846,N_6983);
and U7177 (N_7177,N_6868,N_6945);
nand U7178 (N_7178,N_6966,N_6974);
nand U7179 (N_7179,N_6838,N_6897);
nand U7180 (N_7180,N_6994,N_6844);
nor U7181 (N_7181,N_6882,N_6913);
nand U7182 (N_7182,N_6897,N_6825);
nand U7183 (N_7183,N_6989,N_6878);
or U7184 (N_7184,N_6906,N_6847);
nor U7185 (N_7185,N_6960,N_6901);
and U7186 (N_7186,N_6913,N_6806);
or U7187 (N_7187,N_6915,N_6983);
nor U7188 (N_7188,N_6836,N_6837);
or U7189 (N_7189,N_6931,N_6937);
nand U7190 (N_7190,N_6906,N_6833);
and U7191 (N_7191,N_6924,N_6984);
nor U7192 (N_7192,N_6893,N_6853);
nand U7193 (N_7193,N_6923,N_6955);
nor U7194 (N_7194,N_6894,N_6801);
and U7195 (N_7195,N_6862,N_6956);
and U7196 (N_7196,N_6916,N_6816);
and U7197 (N_7197,N_6938,N_6929);
nand U7198 (N_7198,N_6947,N_6908);
and U7199 (N_7199,N_6840,N_6930);
and U7200 (N_7200,N_7181,N_7169);
nand U7201 (N_7201,N_7178,N_7044);
and U7202 (N_7202,N_7147,N_7173);
and U7203 (N_7203,N_7096,N_7174);
and U7204 (N_7204,N_7047,N_7001);
nor U7205 (N_7205,N_7087,N_7120);
nand U7206 (N_7206,N_7146,N_7075);
or U7207 (N_7207,N_7003,N_7086);
nand U7208 (N_7208,N_7078,N_7062);
or U7209 (N_7209,N_7068,N_7106);
nand U7210 (N_7210,N_7130,N_7186);
nand U7211 (N_7211,N_7183,N_7193);
xnor U7212 (N_7212,N_7065,N_7032);
and U7213 (N_7213,N_7150,N_7105);
and U7214 (N_7214,N_7163,N_7012);
nand U7215 (N_7215,N_7117,N_7058);
nand U7216 (N_7216,N_7164,N_7172);
or U7217 (N_7217,N_7092,N_7110);
nor U7218 (N_7218,N_7119,N_7094);
and U7219 (N_7219,N_7069,N_7165);
nor U7220 (N_7220,N_7064,N_7074);
nand U7221 (N_7221,N_7160,N_7030);
and U7222 (N_7222,N_7148,N_7052);
nor U7223 (N_7223,N_7066,N_7070);
nor U7224 (N_7224,N_7152,N_7157);
and U7225 (N_7225,N_7054,N_7133);
and U7226 (N_7226,N_7084,N_7031);
and U7227 (N_7227,N_7112,N_7190);
xor U7228 (N_7228,N_7161,N_7077);
nor U7229 (N_7229,N_7091,N_7144);
nor U7230 (N_7230,N_7038,N_7145);
nor U7231 (N_7231,N_7015,N_7033);
and U7232 (N_7232,N_7184,N_7081);
and U7233 (N_7233,N_7080,N_7121);
nand U7234 (N_7234,N_7140,N_7175);
nor U7235 (N_7235,N_7107,N_7170);
and U7236 (N_7236,N_7019,N_7051);
and U7237 (N_7237,N_7135,N_7138);
nand U7238 (N_7238,N_7125,N_7109);
nand U7239 (N_7239,N_7000,N_7071);
nor U7240 (N_7240,N_7176,N_7100);
or U7241 (N_7241,N_7020,N_7002);
nand U7242 (N_7242,N_7131,N_7059);
nor U7243 (N_7243,N_7085,N_7057);
xor U7244 (N_7244,N_7056,N_7010);
nor U7245 (N_7245,N_7192,N_7142);
nor U7246 (N_7246,N_7113,N_7154);
nor U7247 (N_7247,N_7045,N_7014);
nand U7248 (N_7248,N_7123,N_7180);
nor U7249 (N_7249,N_7053,N_7095);
nor U7250 (N_7250,N_7049,N_7028);
or U7251 (N_7251,N_7179,N_7016);
and U7252 (N_7252,N_7060,N_7067);
nor U7253 (N_7253,N_7034,N_7006);
and U7254 (N_7254,N_7041,N_7166);
or U7255 (N_7255,N_7168,N_7025);
nand U7256 (N_7256,N_7017,N_7026);
and U7257 (N_7257,N_7188,N_7022);
nand U7258 (N_7258,N_7196,N_7156);
or U7259 (N_7259,N_7050,N_7004);
or U7260 (N_7260,N_7073,N_7018);
nand U7261 (N_7261,N_7013,N_7029);
and U7262 (N_7262,N_7055,N_7090);
or U7263 (N_7263,N_7037,N_7141);
and U7264 (N_7264,N_7143,N_7108);
nand U7265 (N_7265,N_7027,N_7035);
nand U7266 (N_7266,N_7111,N_7177);
nor U7267 (N_7267,N_7153,N_7083);
nor U7268 (N_7268,N_7102,N_7007);
nand U7269 (N_7269,N_7089,N_7199);
and U7270 (N_7270,N_7097,N_7115);
or U7271 (N_7271,N_7195,N_7005);
nand U7272 (N_7272,N_7009,N_7039);
nor U7273 (N_7273,N_7101,N_7122);
and U7274 (N_7274,N_7023,N_7036);
nor U7275 (N_7275,N_7103,N_7191);
nand U7276 (N_7276,N_7116,N_7139);
nor U7277 (N_7277,N_7132,N_7061);
and U7278 (N_7278,N_7118,N_7126);
or U7279 (N_7279,N_7046,N_7158);
or U7280 (N_7280,N_7048,N_7197);
nand U7281 (N_7281,N_7008,N_7082);
or U7282 (N_7282,N_7024,N_7137);
nand U7283 (N_7283,N_7128,N_7043);
nand U7284 (N_7284,N_7155,N_7098);
xor U7285 (N_7285,N_7189,N_7040);
nand U7286 (N_7286,N_7021,N_7079);
and U7287 (N_7287,N_7042,N_7104);
or U7288 (N_7288,N_7063,N_7129);
or U7289 (N_7289,N_7159,N_7167);
xnor U7290 (N_7290,N_7093,N_7194);
or U7291 (N_7291,N_7011,N_7162);
or U7292 (N_7292,N_7187,N_7099);
nor U7293 (N_7293,N_7124,N_7182);
nand U7294 (N_7294,N_7171,N_7072);
and U7295 (N_7295,N_7134,N_7198);
nor U7296 (N_7296,N_7114,N_7127);
and U7297 (N_7297,N_7185,N_7076);
nand U7298 (N_7298,N_7088,N_7136);
or U7299 (N_7299,N_7151,N_7149);
nor U7300 (N_7300,N_7078,N_7181);
nor U7301 (N_7301,N_7136,N_7182);
nand U7302 (N_7302,N_7020,N_7070);
nand U7303 (N_7303,N_7174,N_7184);
or U7304 (N_7304,N_7179,N_7192);
nor U7305 (N_7305,N_7114,N_7047);
nor U7306 (N_7306,N_7110,N_7160);
and U7307 (N_7307,N_7080,N_7144);
or U7308 (N_7308,N_7000,N_7156);
or U7309 (N_7309,N_7173,N_7162);
nor U7310 (N_7310,N_7109,N_7051);
or U7311 (N_7311,N_7174,N_7084);
or U7312 (N_7312,N_7064,N_7194);
or U7313 (N_7313,N_7130,N_7007);
nand U7314 (N_7314,N_7164,N_7008);
nand U7315 (N_7315,N_7165,N_7018);
or U7316 (N_7316,N_7055,N_7007);
nor U7317 (N_7317,N_7103,N_7163);
and U7318 (N_7318,N_7141,N_7026);
or U7319 (N_7319,N_7019,N_7121);
and U7320 (N_7320,N_7125,N_7088);
nand U7321 (N_7321,N_7135,N_7146);
nand U7322 (N_7322,N_7127,N_7052);
nor U7323 (N_7323,N_7158,N_7165);
nor U7324 (N_7324,N_7193,N_7014);
xnor U7325 (N_7325,N_7028,N_7149);
nand U7326 (N_7326,N_7154,N_7139);
or U7327 (N_7327,N_7180,N_7079);
nand U7328 (N_7328,N_7059,N_7051);
and U7329 (N_7329,N_7044,N_7168);
nand U7330 (N_7330,N_7102,N_7155);
nand U7331 (N_7331,N_7032,N_7160);
nand U7332 (N_7332,N_7112,N_7159);
nand U7333 (N_7333,N_7185,N_7050);
nor U7334 (N_7334,N_7125,N_7142);
or U7335 (N_7335,N_7077,N_7192);
or U7336 (N_7336,N_7068,N_7082);
nor U7337 (N_7337,N_7095,N_7115);
nand U7338 (N_7338,N_7101,N_7012);
nand U7339 (N_7339,N_7197,N_7020);
nand U7340 (N_7340,N_7075,N_7076);
and U7341 (N_7341,N_7006,N_7153);
nor U7342 (N_7342,N_7055,N_7185);
or U7343 (N_7343,N_7197,N_7122);
or U7344 (N_7344,N_7007,N_7042);
nand U7345 (N_7345,N_7190,N_7136);
nor U7346 (N_7346,N_7135,N_7002);
and U7347 (N_7347,N_7134,N_7185);
nand U7348 (N_7348,N_7004,N_7117);
and U7349 (N_7349,N_7049,N_7179);
nand U7350 (N_7350,N_7047,N_7136);
nand U7351 (N_7351,N_7110,N_7050);
and U7352 (N_7352,N_7107,N_7025);
and U7353 (N_7353,N_7096,N_7147);
or U7354 (N_7354,N_7138,N_7151);
nand U7355 (N_7355,N_7026,N_7156);
or U7356 (N_7356,N_7044,N_7004);
or U7357 (N_7357,N_7078,N_7027);
and U7358 (N_7358,N_7181,N_7005);
nor U7359 (N_7359,N_7160,N_7059);
nor U7360 (N_7360,N_7154,N_7199);
or U7361 (N_7361,N_7149,N_7180);
nand U7362 (N_7362,N_7065,N_7198);
nor U7363 (N_7363,N_7141,N_7032);
nor U7364 (N_7364,N_7142,N_7066);
nand U7365 (N_7365,N_7134,N_7094);
and U7366 (N_7366,N_7109,N_7150);
nor U7367 (N_7367,N_7197,N_7109);
and U7368 (N_7368,N_7042,N_7044);
or U7369 (N_7369,N_7041,N_7035);
nor U7370 (N_7370,N_7159,N_7186);
nor U7371 (N_7371,N_7042,N_7165);
or U7372 (N_7372,N_7105,N_7165);
or U7373 (N_7373,N_7004,N_7055);
or U7374 (N_7374,N_7016,N_7157);
nand U7375 (N_7375,N_7130,N_7082);
nand U7376 (N_7376,N_7057,N_7051);
nand U7377 (N_7377,N_7063,N_7185);
or U7378 (N_7378,N_7104,N_7073);
nor U7379 (N_7379,N_7150,N_7164);
or U7380 (N_7380,N_7064,N_7163);
nand U7381 (N_7381,N_7117,N_7166);
nand U7382 (N_7382,N_7094,N_7159);
and U7383 (N_7383,N_7000,N_7031);
nor U7384 (N_7384,N_7159,N_7176);
nand U7385 (N_7385,N_7054,N_7135);
and U7386 (N_7386,N_7051,N_7143);
and U7387 (N_7387,N_7193,N_7166);
or U7388 (N_7388,N_7174,N_7142);
nor U7389 (N_7389,N_7027,N_7104);
or U7390 (N_7390,N_7089,N_7111);
nand U7391 (N_7391,N_7179,N_7184);
nand U7392 (N_7392,N_7077,N_7102);
nor U7393 (N_7393,N_7064,N_7155);
nand U7394 (N_7394,N_7194,N_7107);
xor U7395 (N_7395,N_7102,N_7054);
and U7396 (N_7396,N_7101,N_7092);
and U7397 (N_7397,N_7100,N_7022);
and U7398 (N_7398,N_7156,N_7011);
and U7399 (N_7399,N_7192,N_7128);
and U7400 (N_7400,N_7303,N_7378);
and U7401 (N_7401,N_7293,N_7371);
nor U7402 (N_7402,N_7324,N_7284);
or U7403 (N_7403,N_7304,N_7297);
and U7404 (N_7404,N_7323,N_7399);
and U7405 (N_7405,N_7238,N_7215);
and U7406 (N_7406,N_7310,N_7338);
nor U7407 (N_7407,N_7203,N_7241);
nor U7408 (N_7408,N_7397,N_7329);
or U7409 (N_7409,N_7246,N_7318);
nand U7410 (N_7410,N_7382,N_7229);
nor U7411 (N_7411,N_7283,N_7377);
nor U7412 (N_7412,N_7279,N_7392);
nand U7413 (N_7413,N_7332,N_7317);
or U7414 (N_7414,N_7295,N_7352);
or U7415 (N_7415,N_7253,N_7263);
nor U7416 (N_7416,N_7398,N_7250);
nand U7417 (N_7417,N_7313,N_7341);
or U7418 (N_7418,N_7208,N_7372);
or U7419 (N_7419,N_7335,N_7376);
or U7420 (N_7420,N_7389,N_7243);
nand U7421 (N_7421,N_7218,N_7268);
nand U7422 (N_7422,N_7307,N_7254);
and U7423 (N_7423,N_7278,N_7275);
or U7424 (N_7424,N_7365,N_7237);
nor U7425 (N_7425,N_7211,N_7395);
or U7426 (N_7426,N_7367,N_7343);
nor U7427 (N_7427,N_7230,N_7280);
nand U7428 (N_7428,N_7384,N_7281);
xor U7429 (N_7429,N_7345,N_7291);
nor U7430 (N_7430,N_7287,N_7260);
and U7431 (N_7431,N_7388,N_7233);
nor U7432 (N_7432,N_7272,N_7370);
nor U7433 (N_7433,N_7270,N_7213);
nand U7434 (N_7434,N_7257,N_7259);
and U7435 (N_7435,N_7312,N_7315);
or U7436 (N_7436,N_7207,N_7245);
nand U7437 (N_7437,N_7276,N_7346);
and U7438 (N_7438,N_7311,N_7214);
and U7439 (N_7439,N_7348,N_7242);
and U7440 (N_7440,N_7220,N_7361);
and U7441 (N_7441,N_7256,N_7383);
nand U7442 (N_7442,N_7262,N_7201);
nand U7443 (N_7443,N_7342,N_7349);
or U7444 (N_7444,N_7255,N_7248);
nand U7445 (N_7445,N_7296,N_7277);
xor U7446 (N_7446,N_7269,N_7351);
nand U7447 (N_7447,N_7337,N_7327);
or U7448 (N_7448,N_7290,N_7212);
nor U7449 (N_7449,N_7266,N_7223);
or U7450 (N_7450,N_7299,N_7357);
or U7451 (N_7451,N_7339,N_7350);
or U7452 (N_7452,N_7267,N_7288);
and U7453 (N_7453,N_7217,N_7302);
nand U7454 (N_7454,N_7334,N_7273);
or U7455 (N_7455,N_7228,N_7387);
xor U7456 (N_7456,N_7309,N_7355);
or U7457 (N_7457,N_7251,N_7204);
or U7458 (N_7458,N_7219,N_7359);
nand U7459 (N_7459,N_7285,N_7271);
and U7460 (N_7460,N_7247,N_7385);
nor U7461 (N_7461,N_7325,N_7320);
xor U7462 (N_7462,N_7354,N_7356);
and U7463 (N_7463,N_7210,N_7374);
and U7464 (N_7464,N_7234,N_7227);
or U7465 (N_7465,N_7373,N_7347);
nor U7466 (N_7466,N_7336,N_7200);
nand U7467 (N_7467,N_7236,N_7202);
or U7468 (N_7468,N_7344,N_7235);
nor U7469 (N_7469,N_7221,N_7239);
nor U7470 (N_7470,N_7396,N_7340);
nand U7471 (N_7471,N_7333,N_7319);
and U7472 (N_7472,N_7375,N_7390);
or U7473 (N_7473,N_7393,N_7326);
xor U7474 (N_7474,N_7362,N_7353);
nand U7475 (N_7475,N_7289,N_7294);
nand U7476 (N_7476,N_7301,N_7394);
or U7477 (N_7477,N_7331,N_7322);
and U7478 (N_7478,N_7380,N_7358);
nor U7479 (N_7479,N_7232,N_7381);
nand U7480 (N_7480,N_7205,N_7265);
or U7481 (N_7481,N_7391,N_7206);
nand U7482 (N_7482,N_7363,N_7298);
nand U7483 (N_7483,N_7282,N_7274);
nor U7484 (N_7484,N_7386,N_7328);
nand U7485 (N_7485,N_7226,N_7368);
nand U7486 (N_7486,N_7369,N_7321);
nand U7487 (N_7487,N_7225,N_7300);
nor U7488 (N_7488,N_7264,N_7216);
nand U7489 (N_7489,N_7249,N_7252);
or U7490 (N_7490,N_7244,N_7316);
nand U7491 (N_7491,N_7224,N_7308);
nor U7492 (N_7492,N_7261,N_7286);
xnor U7493 (N_7493,N_7305,N_7330);
nor U7494 (N_7494,N_7292,N_7231);
or U7495 (N_7495,N_7360,N_7222);
or U7496 (N_7496,N_7364,N_7314);
or U7497 (N_7497,N_7240,N_7366);
xnor U7498 (N_7498,N_7306,N_7258);
nor U7499 (N_7499,N_7379,N_7209);
or U7500 (N_7500,N_7314,N_7333);
nand U7501 (N_7501,N_7385,N_7290);
or U7502 (N_7502,N_7228,N_7243);
nand U7503 (N_7503,N_7302,N_7312);
and U7504 (N_7504,N_7349,N_7296);
and U7505 (N_7505,N_7300,N_7204);
or U7506 (N_7506,N_7209,N_7280);
and U7507 (N_7507,N_7399,N_7386);
and U7508 (N_7508,N_7326,N_7385);
nor U7509 (N_7509,N_7214,N_7284);
and U7510 (N_7510,N_7338,N_7337);
or U7511 (N_7511,N_7289,N_7211);
or U7512 (N_7512,N_7202,N_7229);
and U7513 (N_7513,N_7203,N_7334);
nor U7514 (N_7514,N_7211,N_7213);
or U7515 (N_7515,N_7254,N_7368);
nand U7516 (N_7516,N_7383,N_7354);
nand U7517 (N_7517,N_7381,N_7314);
and U7518 (N_7518,N_7201,N_7346);
nor U7519 (N_7519,N_7306,N_7374);
xor U7520 (N_7520,N_7201,N_7314);
xor U7521 (N_7521,N_7344,N_7368);
nor U7522 (N_7522,N_7270,N_7303);
and U7523 (N_7523,N_7329,N_7267);
nand U7524 (N_7524,N_7327,N_7365);
nand U7525 (N_7525,N_7314,N_7338);
xor U7526 (N_7526,N_7234,N_7200);
and U7527 (N_7527,N_7215,N_7369);
and U7528 (N_7528,N_7221,N_7312);
and U7529 (N_7529,N_7240,N_7244);
nand U7530 (N_7530,N_7246,N_7370);
nand U7531 (N_7531,N_7344,N_7290);
nor U7532 (N_7532,N_7309,N_7315);
nor U7533 (N_7533,N_7284,N_7388);
and U7534 (N_7534,N_7382,N_7247);
and U7535 (N_7535,N_7325,N_7362);
nor U7536 (N_7536,N_7217,N_7228);
nor U7537 (N_7537,N_7222,N_7215);
nor U7538 (N_7538,N_7208,N_7289);
or U7539 (N_7539,N_7352,N_7211);
and U7540 (N_7540,N_7344,N_7289);
xor U7541 (N_7541,N_7354,N_7254);
nor U7542 (N_7542,N_7330,N_7364);
or U7543 (N_7543,N_7392,N_7255);
nand U7544 (N_7544,N_7281,N_7201);
nand U7545 (N_7545,N_7360,N_7395);
or U7546 (N_7546,N_7217,N_7316);
nand U7547 (N_7547,N_7353,N_7381);
or U7548 (N_7548,N_7260,N_7240);
or U7549 (N_7549,N_7282,N_7205);
or U7550 (N_7550,N_7276,N_7291);
nand U7551 (N_7551,N_7299,N_7324);
nand U7552 (N_7552,N_7390,N_7343);
nor U7553 (N_7553,N_7221,N_7331);
or U7554 (N_7554,N_7270,N_7391);
and U7555 (N_7555,N_7375,N_7383);
nand U7556 (N_7556,N_7360,N_7275);
nor U7557 (N_7557,N_7227,N_7207);
nand U7558 (N_7558,N_7374,N_7230);
or U7559 (N_7559,N_7257,N_7206);
nand U7560 (N_7560,N_7236,N_7263);
or U7561 (N_7561,N_7226,N_7327);
or U7562 (N_7562,N_7245,N_7292);
nand U7563 (N_7563,N_7391,N_7267);
nor U7564 (N_7564,N_7207,N_7308);
and U7565 (N_7565,N_7346,N_7367);
xor U7566 (N_7566,N_7330,N_7362);
and U7567 (N_7567,N_7265,N_7251);
nor U7568 (N_7568,N_7292,N_7398);
nor U7569 (N_7569,N_7266,N_7271);
or U7570 (N_7570,N_7334,N_7291);
and U7571 (N_7571,N_7326,N_7266);
nand U7572 (N_7572,N_7333,N_7372);
and U7573 (N_7573,N_7395,N_7303);
or U7574 (N_7574,N_7341,N_7271);
nor U7575 (N_7575,N_7368,N_7277);
nor U7576 (N_7576,N_7310,N_7347);
nor U7577 (N_7577,N_7264,N_7302);
nand U7578 (N_7578,N_7212,N_7364);
and U7579 (N_7579,N_7331,N_7378);
nand U7580 (N_7580,N_7346,N_7249);
nor U7581 (N_7581,N_7308,N_7251);
nor U7582 (N_7582,N_7345,N_7256);
nand U7583 (N_7583,N_7359,N_7222);
and U7584 (N_7584,N_7220,N_7385);
or U7585 (N_7585,N_7218,N_7276);
nor U7586 (N_7586,N_7297,N_7224);
and U7587 (N_7587,N_7306,N_7369);
nor U7588 (N_7588,N_7293,N_7258);
nand U7589 (N_7589,N_7288,N_7343);
and U7590 (N_7590,N_7250,N_7335);
and U7591 (N_7591,N_7376,N_7316);
or U7592 (N_7592,N_7307,N_7323);
nand U7593 (N_7593,N_7244,N_7379);
and U7594 (N_7594,N_7323,N_7372);
nor U7595 (N_7595,N_7203,N_7386);
and U7596 (N_7596,N_7233,N_7277);
nor U7597 (N_7597,N_7327,N_7293);
nor U7598 (N_7598,N_7260,N_7272);
nor U7599 (N_7599,N_7227,N_7322);
nor U7600 (N_7600,N_7570,N_7595);
nor U7601 (N_7601,N_7492,N_7454);
nor U7602 (N_7602,N_7512,N_7448);
or U7603 (N_7603,N_7515,N_7554);
nand U7604 (N_7604,N_7551,N_7547);
or U7605 (N_7605,N_7510,N_7536);
or U7606 (N_7606,N_7452,N_7412);
nor U7607 (N_7607,N_7479,N_7577);
or U7608 (N_7608,N_7499,N_7453);
or U7609 (N_7609,N_7578,N_7470);
or U7610 (N_7610,N_7420,N_7565);
xnor U7611 (N_7611,N_7500,N_7569);
or U7612 (N_7612,N_7415,N_7407);
nor U7613 (N_7613,N_7509,N_7550);
or U7614 (N_7614,N_7481,N_7418);
or U7615 (N_7615,N_7523,N_7444);
nand U7616 (N_7616,N_7588,N_7506);
xor U7617 (N_7617,N_7482,N_7438);
and U7618 (N_7618,N_7439,N_7540);
nor U7619 (N_7619,N_7513,N_7432);
or U7620 (N_7620,N_7502,N_7450);
or U7621 (N_7621,N_7404,N_7562);
nand U7622 (N_7622,N_7596,N_7576);
xor U7623 (N_7623,N_7514,N_7528);
or U7624 (N_7624,N_7477,N_7590);
and U7625 (N_7625,N_7429,N_7445);
nor U7626 (N_7626,N_7497,N_7451);
nor U7627 (N_7627,N_7521,N_7517);
or U7628 (N_7628,N_7440,N_7427);
or U7629 (N_7629,N_7449,N_7443);
and U7630 (N_7630,N_7431,N_7469);
and U7631 (N_7631,N_7423,N_7435);
nor U7632 (N_7632,N_7486,N_7543);
nand U7633 (N_7633,N_7422,N_7561);
nand U7634 (N_7634,N_7413,N_7507);
nor U7635 (N_7635,N_7518,N_7498);
and U7636 (N_7636,N_7574,N_7476);
and U7637 (N_7637,N_7530,N_7546);
or U7638 (N_7638,N_7433,N_7579);
or U7639 (N_7639,N_7471,N_7573);
nor U7640 (N_7640,N_7527,N_7472);
and U7641 (N_7641,N_7417,N_7409);
and U7642 (N_7642,N_7566,N_7549);
and U7643 (N_7643,N_7511,N_7463);
nor U7644 (N_7644,N_7456,N_7411);
or U7645 (N_7645,N_7465,N_7437);
and U7646 (N_7646,N_7504,N_7589);
nor U7647 (N_7647,N_7494,N_7458);
nand U7648 (N_7648,N_7559,N_7406);
and U7649 (N_7649,N_7583,N_7582);
and U7650 (N_7650,N_7410,N_7503);
nand U7651 (N_7651,N_7544,N_7442);
or U7652 (N_7652,N_7400,N_7403);
or U7653 (N_7653,N_7493,N_7421);
and U7654 (N_7654,N_7446,N_7560);
nand U7655 (N_7655,N_7462,N_7484);
nand U7656 (N_7656,N_7466,N_7485);
or U7657 (N_7657,N_7594,N_7541);
and U7658 (N_7658,N_7581,N_7496);
nor U7659 (N_7659,N_7414,N_7531);
nor U7660 (N_7660,N_7534,N_7402);
or U7661 (N_7661,N_7478,N_7473);
or U7662 (N_7662,N_7533,N_7508);
and U7663 (N_7663,N_7556,N_7436);
nor U7664 (N_7664,N_7592,N_7572);
or U7665 (N_7665,N_7424,N_7571);
nand U7666 (N_7666,N_7416,N_7524);
and U7667 (N_7667,N_7520,N_7430);
or U7668 (N_7668,N_7419,N_7401);
nand U7669 (N_7669,N_7584,N_7428);
and U7670 (N_7670,N_7405,N_7487);
nor U7671 (N_7671,N_7459,N_7548);
and U7672 (N_7672,N_7563,N_7558);
nand U7673 (N_7673,N_7447,N_7529);
nand U7674 (N_7674,N_7585,N_7467);
nor U7675 (N_7675,N_7455,N_7593);
nor U7676 (N_7676,N_7542,N_7599);
and U7677 (N_7677,N_7538,N_7460);
and U7678 (N_7678,N_7580,N_7525);
or U7679 (N_7679,N_7537,N_7490);
nand U7680 (N_7680,N_7426,N_7434);
or U7681 (N_7681,N_7553,N_7597);
nor U7682 (N_7682,N_7575,N_7522);
nor U7683 (N_7683,N_7591,N_7489);
and U7684 (N_7684,N_7480,N_7408);
nand U7685 (N_7685,N_7568,N_7468);
nand U7686 (N_7686,N_7526,N_7491);
nor U7687 (N_7687,N_7557,N_7516);
nand U7688 (N_7688,N_7535,N_7495);
or U7689 (N_7689,N_7461,N_7483);
xor U7690 (N_7690,N_7598,N_7505);
and U7691 (N_7691,N_7564,N_7425);
and U7692 (N_7692,N_7501,N_7457);
and U7693 (N_7693,N_7475,N_7587);
or U7694 (N_7694,N_7539,N_7474);
and U7695 (N_7695,N_7586,N_7545);
nor U7696 (N_7696,N_7519,N_7488);
nor U7697 (N_7697,N_7555,N_7552);
nor U7698 (N_7698,N_7567,N_7441);
and U7699 (N_7699,N_7532,N_7464);
or U7700 (N_7700,N_7513,N_7536);
and U7701 (N_7701,N_7599,N_7459);
or U7702 (N_7702,N_7446,N_7569);
nor U7703 (N_7703,N_7591,N_7494);
nor U7704 (N_7704,N_7457,N_7517);
nor U7705 (N_7705,N_7584,N_7426);
nand U7706 (N_7706,N_7569,N_7586);
nand U7707 (N_7707,N_7424,N_7435);
nand U7708 (N_7708,N_7400,N_7558);
nand U7709 (N_7709,N_7404,N_7470);
nor U7710 (N_7710,N_7498,N_7401);
nand U7711 (N_7711,N_7567,N_7495);
and U7712 (N_7712,N_7560,N_7536);
nor U7713 (N_7713,N_7464,N_7423);
nor U7714 (N_7714,N_7463,N_7458);
or U7715 (N_7715,N_7589,N_7573);
or U7716 (N_7716,N_7550,N_7491);
nand U7717 (N_7717,N_7402,N_7462);
nand U7718 (N_7718,N_7459,N_7483);
or U7719 (N_7719,N_7488,N_7523);
nor U7720 (N_7720,N_7599,N_7556);
and U7721 (N_7721,N_7429,N_7479);
or U7722 (N_7722,N_7429,N_7502);
xor U7723 (N_7723,N_7501,N_7432);
and U7724 (N_7724,N_7451,N_7437);
and U7725 (N_7725,N_7431,N_7592);
and U7726 (N_7726,N_7564,N_7491);
and U7727 (N_7727,N_7469,N_7430);
and U7728 (N_7728,N_7587,N_7403);
nand U7729 (N_7729,N_7402,N_7490);
and U7730 (N_7730,N_7491,N_7486);
nand U7731 (N_7731,N_7449,N_7512);
nand U7732 (N_7732,N_7509,N_7549);
nor U7733 (N_7733,N_7509,N_7558);
or U7734 (N_7734,N_7409,N_7584);
nor U7735 (N_7735,N_7577,N_7542);
or U7736 (N_7736,N_7429,N_7576);
nand U7737 (N_7737,N_7451,N_7426);
nor U7738 (N_7738,N_7548,N_7476);
or U7739 (N_7739,N_7538,N_7433);
or U7740 (N_7740,N_7576,N_7588);
or U7741 (N_7741,N_7592,N_7470);
nand U7742 (N_7742,N_7466,N_7488);
and U7743 (N_7743,N_7531,N_7488);
nor U7744 (N_7744,N_7494,N_7483);
nand U7745 (N_7745,N_7509,N_7463);
nand U7746 (N_7746,N_7599,N_7555);
and U7747 (N_7747,N_7598,N_7499);
nor U7748 (N_7748,N_7521,N_7571);
or U7749 (N_7749,N_7436,N_7586);
or U7750 (N_7750,N_7412,N_7544);
nand U7751 (N_7751,N_7470,N_7556);
or U7752 (N_7752,N_7423,N_7574);
or U7753 (N_7753,N_7452,N_7471);
and U7754 (N_7754,N_7509,N_7581);
nor U7755 (N_7755,N_7573,N_7401);
or U7756 (N_7756,N_7545,N_7588);
or U7757 (N_7757,N_7461,N_7428);
and U7758 (N_7758,N_7526,N_7463);
nand U7759 (N_7759,N_7431,N_7413);
or U7760 (N_7760,N_7560,N_7591);
nor U7761 (N_7761,N_7412,N_7551);
nand U7762 (N_7762,N_7496,N_7507);
xor U7763 (N_7763,N_7442,N_7471);
nor U7764 (N_7764,N_7443,N_7592);
nor U7765 (N_7765,N_7594,N_7505);
nor U7766 (N_7766,N_7546,N_7446);
or U7767 (N_7767,N_7505,N_7514);
nor U7768 (N_7768,N_7466,N_7400);
nand U7769 (N_7769,N_7523,N_7565);
nand U7770 (N_7770,N_7555,N_7545);
nand U7771 (N_7771,N_7583,N_7576);
nor U7772 (N_7772,N_7533,N_7427);
or U7773 (N_7773,N_7519,N_7414);
or U7774 (N_7774,N_7470,N_7437);
and U7775 (N_7775,N_7539,N_7491);
nand U7776 (N_7776,N_7558,N_7507);
nor U7777 (N_7777,N_7506,N_7516);
or U7778 (N_7778,N_7563,N_7473);
nor U7779 (N_7779,N_7535,N_7419);
nor U7780 (N_7780,N_7501,N_7472);
and U7781 (N_7781,N_7559,N_7442);
nor U7782 (N_7782,N_7473,N_7524);
nor U7783 (N_7783,N_7544,N_7491);
or U7784 (N_7784,N_7556,N_7481);
and U7785 (N_7785,N_7559,N_7494);
nor U7786 (N_7786,N_7407,N_7401);
nand U7787 (N_7787,N_7405,N_7457);
nand U7788 (N_7788,N_7416,N_7572);
and U7789 (N_7789,N_7563,N_7529);
and U7790 (N_7790,N_7425,N_7545);
and U7791 (N_7791,N_7564,N_7495);
nand U7792 (N_7792,N_7486,N_7535);
or U7793 (N_7793,N_7508,N_7418);
or U7794 (N_7794,N_7436,N_7482);
and U7795 (N_7795,N_7496,N_7526);
nor U7796 (N_7796,N_7526,N_7445);
nor U7797 (N_7797,N_7453,N_7580);
nand U7798 (N_7798,N_7465,N_7459);
or U7799 (N_7799,N_7576,N_7407);
and U7800 (N_7800,N_7648,N_7730);
or U7801 (N_7801,N_7635,N_7766);
nor U7802 (N_7802,N_7614,N_7627);
or U7803 (N_7803,N_7675,N_7640);
nand U7804 (N_7804,N_7787,N_7637);
nor U7805 (N_7805,N_7795,N_7779);
xor U7806 (N_7806,N_7645,N_7747);
nand U7807 (N_7807,N_7647,N_7789);
nor U7808 (N_7808,N_7683,N_7642);
nor U7809 (N_7809,N_7735,N_7678);
or U7810 (N_7810,N_7691,N_7703);
nand U7811 (N_7811,N_7781,N_7764);
and U7812 (N_7812,N_7743,N_7639);
or U7813 (N_7813,N_7757,N_7667);
and U7814 (N_7814,N_7721,N_7776);
or U7815 (N_7815,N_7649,N_7794);
nor U7816 (N_7816,N_7708,N_7613);
and U7817 (N_7817,N_7632,N_7710);
and U7818 (N_7818,N_7713,N_7609);
or U7819 (N_7819,N_7755,N_7748);
nand U7820 (N_7820,N_7686,N_7744);
xnor U7821 (N_7821,N_7726,N_7716);
nand U7822 (N_7822,N_7671,N_7601);
nor U7823 (N_7823,N_7669,N_7623);
or U7824 (N_7824,N_7604,N_7692);
or U7825 (N_7825,N_7799,N_7754);
and U7826 (N_7826,N_7783,N_7780);
and U7827 (N_7827,N_7651,N_7670);
nand U7828 (N_7828,N_7600,N_7786);
nor U7829 (N_7829,N_7631,N_7778);
nand U7830 (N_7830,N_7619,N_7700);
nand U7831 (N_7831,N_7681,N_7694);
nand U7832 (N_7832,N_7750,N_7602);
or U7833 (N_7833,N_7676,N_7665);
nor U7834 (N_7834,N_7773,N_7620);
nand U7835 (N_7835,N_7608,N_7607);
xnor U7836 (N_7836,N_7654,N_7634);
and U7837 (N_7837,N_7693,N_7785);
xor U7838 (N_7838,N_7762,N_7734);
and U7839 (N_7839,N_7680,N_7701);
and U7840 (N_7840,N_7659,N_7624);
nor U7841 (N_7841,N_7740,N_7769);
nor U7842 (N_7842,N_7771,N_7630);
and U7843 (N_7843,N_7768,N_7626);
and U7844 (N_7844,N_7695,N_7749);
nand U7845 (N_7845,N_7760,N_7663);
or U7846 (N_7846,N_7666,N_7603);
nor U7847 (N_7847,N_7690,N_7796);
and U7848 (N_7848,N_7798,N_7706);
nor U7849 (N_7849,N_7605,N_7793);
nor U7850 (N_7850,N_7739,N_7775);
nand U7851 (N_7851,N_7628,N_7724);
nor U7852 (N_7852,N_7633,N_7790);
nand U7853 (N_7853,N_7759,N_7688);
and U7854 (N_7854,N_7705,N_7758);
nor U7855 (N_7855,N_7714,N_7711);
and U7856 (N_7856,N_7615,N_7732);
nand U7857 (N_7857,N_7772,N_7636);
nor U7858 (N_7858,N_7718,N_7660);
or U7859 (N_7859,N_7712,N_7767);
xnor U7860 (N_7860,N_7717,N_7606);
or U7861 (N_7861,N_7737,N_7731);
nand U7862 (N_7862,N_7753,N_7657);
nand U7863 (N_7863,N_7622,N_7650);
nor U7864 (N_7864,N_7728,N_7738);
nand U7865 (N_7865,N_7644,N_7611);
nor U7866 (N_7866,N_7733,N_7797);
and U7867 (N_7867,N_7697,N_7662);
or U7868 (N_7868,N_7610,N_7707);
nand U7869 (N_7869,N_7655,N_7638);
or U7870 (N_7870,N_7621,N_7677);
nor U7871 (N_7871,N_7653,N_7745);
or U7872 (N_7872,N_7646,N_7661);
nand U7873 (N_7873,N_7777,N_7702);
xor U7874 (N_7874,N_7682,N_7679);
nor U7875 (N_7875,N_7656,N_7641);
nor U7876 (N_7876,N_7756,N_7696);
or U7877 (N_7877,N_7723,N_7765);
nand U7878 (N_7878,N_7782,N_7770);
and U7879 (N_7879,N_7684,N_7652);
nand U7880 (N_7880,N_7725,N_7719);
nand U7881 (N_7881,N_7784,N_7698);
nor U7882 (N_7882,N_7672,N_7612);
and U7883 (N_7883,N_7741,N_7746);
nand U7884 (N_7884,N_7727,N_7715);
or U7885 (N_7885,N_7673,N_7788);
and U7886 (N_7886,N_7616,N_7689);
nor U7887 (N_7887,N_7704,N_7742);
nand U7888 (N_7888,N_7664,N_7774);
and U7889 (N_7889,N_7763,N_7729);
and U7890 (N_7890,N_7617,N_7668);
nor U7891 (N_7891,N_7722,N_7658);
nor U7892 (N_7892,N_7699,N_7752);
and U7893 (N_7893,N_7736,N_7685);
or U7894 (N_7894,N_7761,N_7791);
or U7895 (N_7895,N_7618,N_7709);
nand U7896 (N_7896,N_7687,N_7643);
nand U7897 (N_7897,N_7625,N_7751);
and U7898 (N_7898,N_7720,N_7792);
and U7899 (N_7899,N_7674,N_7629);
and U7900 (N_7900,N_7618,N_7607);
nor U7901 (N_7901,N_7745,N_7713);
nand U7902 (N_7902,N_7760,N_7603);
nor U7903 (N_7903,N_7754,N_7679);
nand U7904 (N_7904,N_7613,N_7634);
and U7905 (N_7905,N_7691,N_7667);
nor U7906 (N_7906,N_7738,N_7699);
and U7907 (N_7907,N_7669,N_7718);
xnor U7908 (N_7908,N_7631,N_7623);
nand U7909 (N_7909,N_7604,N_7729);
and U7910 (N_7910,N_7676,N_7732);
nor U7911 (N_7911,N_7678,N_7746);
nand U7912 (N_7912,N_7620,N_7642);
or U7913 (N_7913,N_7643,N_7774);
nor U7914 (N_7914,N_7732,N_7670);
or U7915 (N_7915,N_7786,N_7753);
and U7916 (N_7916,N_7690,N_7636);
or U7917 (N_7917,N_7771,N_7729);
xor U7918 (N_7918,N_7614,N_7659);
xnor U7919 (N_7919,N_7694,N_7638);
or U7920 (N_7920,N_7780,N_7763);
nand U7921 (N_7921,N_7645,N_7789);
nor U7922 (N_7922,N_7649,N_7778);
nor U7923 (N_7923,N_7711,N_7682);
or U7924 (N_7924,N_7715,N_7747);
nor U7925 (N_7925,N_7640,N_7798);
nor U7926 (N_7926,N_7629,N_7787);
nor U7927 (N_7927,N_7791,N_7783);
nand U7928 (N_7928,N_7703,N_7613);
xor U7929 (N_7929,N_7794,N_7603);
and U7930 (N_7930,N_7764,N_7701);
nor U7931 (N_7931,N_7612,N_7790);
nor U7932 (N_7932,N_7796,N_7775);
or U7933 (N_7933,N_7656,N_7738);
nor U7934 (N_7934,N_7742,N_7692);
and U7935 (N_7935,N_7635,N_7746);
or U7936 (N_7936,N_7751,N_7766);
or U7937 (N_7937,N_7685,N_7695);
nand U7938 (N_7938,N_7682,N_7735);
nor U7939 (N_7939,N_7606,N_7652);
and U7940 (N_7940,N_7679,N_7768);
and U7941 (N_7941,N_7694,N_7724);
nand U7942 (N_7942,N_7703,N_7709);
nor U7943 (N_7943,N_7714,N_7700);
nand U7944 (N_7944,N_7787,N_7662);
nor U7945 (N_7945,N_7674,N_7718);
nand U7946 (N_7946,N_7632,N_7638);
or U7947 (N_7947,N_7614,N_7678);
or U7948 (N_7948,N_7674,N_7643);
nor U7949 (N_7949,N_7651,N_7729);
and U7950 (N_7950,N_7677,N_7799);
nor U7951 (N_7951,N_7603,N_7693);
nand U7952 (N_7952,N_7635,N_7609);
nor U7953 (N_7953,N_7664,N_7705);
and U7954 (N_7954,N_7751,N_7614);
and U7955 (N_7955,N_7606,N_7690);
nand U7956 (N_7956,N_7757,N_7765);
nand U7957 (N_7957,N_7783,N_7683);
or U7958 (N_7958,N_7648,N_7794);
or U7959 (N_7959,N_7606,N_7642);
or U7960 (N_7960,N_7681,N_7778);
nand U7961 (N_7961,N_7726,N_7621);
nor U7962 (N_7962,N_7793,N_7663);
nand U7963 (N_7963,N_7660,N_7629);
and U7964 (N_7964,N_7725,N_7644);
nand U7965 (N_7965,N_7653,N_7693);
nor U7966 (N_7966,N_7670,N_7758);
nand U7967 (N_7967,N_7753,N_7648);
or U7968 (N_7968,N_7647,N_7661);
nor U7969 (N_7969,N_7722,N_7628);
or U7970 (N_7970,N_7746,N_7674);
nor U7971 (N_7971,N_7763,N_7743);
nand U7972 (N_7972,N_7633,N_7748);
xnor U7973 (N_7973,N_7726,N_7677);
nor U7974 (N_7974,N_7781,N_7633);
and U7975 (N_7975,N_7756,N_7607);
and U7976 (N_7976,N_7719,N_7783);
and U7977 (N_7977,N_7603,N_7673);
and U7978 (N_7978,N_7623,N_7656);
or U7979 (N_7979,N_7794,N_7778);
nand U7980 (N_7980,N_7687,N_7742);
or U7981 (N_7981,N_7763,N_7792);
and U7982 (N_7982,N_7641,N_7638);
and U7983 (N_7983,N_7757,N_7619);
and U7984 (N_7984,N_7667,N_7604);
nand U7985 (N_7985,N_7701,N_7676);
nand U7986 (N_7986,N_7746,N_7602);
nand U7987 (N_7987,N_7772,N_7758);
and U7988 (N_7988,N_7663,N_7670);
nand U7989 (N_7989,N_7609,N_7610);
or U7990 (N_7990,N_7776,N_7630);
and U7991 (N_7991,N_7657,N_7767);
nor U7992 (N_7992,N_7755,N_7762);
and U7993 (N_7993,N_7776,N_7766);
or U7994 (N_7994,N_7614,N_7782);
nand U7995 (N_7995,N_7675,N_7653);
nor U7996 (N_7996,N_7693,N_7688);
nor U7997 (N_7997,N_7683,N_7787);
nand U7998 (N_7998,N_7637,N_7648);
nor U7999 (N_7999,N_7739,N_7601);
xor U8000 (N_8000,N_7872,N_7902);
and U8001 (N_8001,N_7854,N_7873);
and U8002 (N_8002,N_7940,N_7827);
nor U8003 (N_8003,N_7859,N_7843);
and U8004 (N_8004,N_7971,N_7945);
xor U8005 (N_8005,N_7907,N_7861);
nor U8006 (N_8006,N_7863,N_7958);
nand U8007 (N_8007,N_7977,N_7949);
nor U8008 (N_8008,N_7813,N_7838);
or U8009 (N_8009,N_7850,N_7981);
nor U8010 (N_8010,N_7928,N_7944);
nand U8011 (N_8011,N_7806,N_7908);
nor U8012 (N_8012,N_7932,N_7978);
or U8013 (N_8013,N_7925,N_7966);
or U8014 (N_8014,N_7990,N_7921);
and U8015 (N_8015,N_7953,N_7807);
and U8016 (N_8016,N_7996,N_7820);
nor U8017 (N_8017,N_7951,N_7826);
nand U8018 (N_8018,N_7892,N_7871);
or U8019 (N_8019,N_7832,N_7917);
or U8020 (N_8020,N_7800,N_7961);
and U8021 (N_8021,N_7954,N_7965);
nand U8022 (N_8022,N_7963,N_7867);
and U8023 (N_8023,N_7803,N_7969);
and U8024 (N_8024,N_7909,N_7984);
or U8025 (N_8025,N_7979,N_7903);
nand U8026 (N_8026,N_7877,N_7889);
nand U8027 (N_8027,N_7960,N_7988);
nor U8028 (N_8028,N_7912,N_7851);
and U8029 (N_8029,N_7989,N_7881);
nand U8030 (N_8030,N_7972,N_7992);
nor U8031 (N_8031,N_7930,N_7878);
xnor U8032 (N_8032,N_7923,N_7842);
or U8033 (N_8033,N_7950,N_7997);
or U8034 (N_8034,N_7916,N_7823);
and U8035 (N_8035,N_7991,N_7887);
and U8036 (N_8036,N_7973,N_7905);
nand U8037 (N_8037,N_7847,N_7821);
or U8038 (N_8038,N_7924,N_7883);
nor U8039 (N_8039,N_7955,N_7938);
nand U8040 (N_8040,N_7957,N_7809);
and U8041 (N_8041,N_7824,N_7865);
and U8042 (N_8042,N_7937,N_7880);
or U8043 (N_8043,N_7913,N_7819);
nor U8044 (N_8044,N_7844,N_7980);
nor U8045 (N_8045,N_7837,N_7993);
and U8046 (N_8046,N_7956,N_7841);
nor U8047 (N_8047,N_7920,N_7895);
or U8048 (N_8048,N_7967,N_7968);
or U8049 (N_8049,N_7939,N_7933);
or U8050 (N_8050,N_7910,N_7868);
or U8051 (N_8051,N_7896,N_7846);
and U8052 (N_8052,N_7879,N_7936);
and U8053 (N_8053,N_7869,N_7948);
nor U8054 (N_8054,N_7946,N_7845);
and U8055 (N_8055,N_7810,N_7964);
and U8056 (N_8056,N_7974,N_7983);
nand U8057 (N_8057,N_7822,N_7839);
or U8058 (N_8058,N_7911,N_7994);
xnor U8059 (N_8059,N_7982,N_7906);
nor U8060 (N_8060,N_7855,N_7853);
nor U8061 (N_8061,N_7901,N_7828);
and U8062 (N_8062,N_7849,N_7833);
or U8063 (N_8063,N_7995,N_7898);
nor U8064 (N_8064,N_7888,N_7857);
nor U8065 (N_8065,N_7840,N_7970);
and U8066 (N_8066,N_7935,N_7922);
nor U8067 (N_8067,N_7904,N_7914);
or U8068 (N_8068,N_7897,N_7947);
nand U8069 (N_8069,N_7926,N_7862);
or U8070 (N_8070,N_7830,N_7858);
nand U8071 (N_8071,N_7801,N_7866);
and U8072 (N_8072,N_7811,N_7816);
and U8073 (N_8073,N_7804,N_7985);
and U8074 (N_8074,N_7856,N_7805);
nor U8075 (N_8075,N_7942,N_7831);
nand U8076 (N_8076,N_7874,N_7986);
nand U8077 (N_8077,N_7919,N_7900);
or U8078 (N_8078,N_7812,N_7952);
and U8079 (N_8079,N_7802,N_7894);
and U8080 (N_8080,N_7918,N_7891);
and U8081 (N_8081,N_7829,N_7836);
and U8082 (N_8082,N_7975,N_7817);
or U8083 (N_8083,N_7870,N_7834);
nor U8084 (N_8084,N_7962,N_7876);
or U8085 (N_8085,N_7941,N_7808);
and U8086 (N_8086,N_7860,N_7884);
or U8087 (N_8087,N_7852,N_7848);
nand U8088 (N_8088,N_7931,N_7893);
nor U8089 (N_8089,N_7929,N_7899);
and U8090 (N_8090,N_7825,N_7814);
nor U8091 (N_8091,N_7998,N_7864);
nor U8092 (N_8092,N_7886,N_7943);
nor U8093 (N_8093,N_7999,N_7875);
nand U8094 (N_8094,N_7959,N_7885);
xor U8095 (N_8095,N_7927,N_7815);
and U8096 (N_8096,N_7915,N_7818);
nor U8097 (N_8097,N_7835,N_7934);
nor U8098 (N_8098,N_7987,N_7976);
or U8099 (N_8099,N_7890,N_7882);
nor U8100 (N_8100,N_7910,N_7960);
nand U8101 (N_8101,N_7995,N_7965);
or U8102 (N_8102,N_7903,N_7852);
nand U8103 (N_8103,N_7976,N_7916);
and U8104 (N_8104,N_7989,N_7890);
or U8105 (N_8105,N_7807,N_7907);
or U8106 (N_8106,N_7825,N_7812);
nor U8107 (N_8107,N_7946,N_7971);
nand U8108 (N_8108,N_7852,N_7800);
and U8109 (N_8109,N_7832,N_7983);
and U8110 (N_8110,N_7947,N_7987);
or U8111 (N_8111,N_7843,N_7874);
nor U8112 (N_8112,N_7822,N_7819);
or U8113 (N_8113,N_7960,N_7974);
and U8114 (N_8114,N_7931,N_7899);
nand U8115 (N_8115,N_7821,N_7842);
nand U8116 (N_8116,N_7961,N_7952);
nor U8117 (N_8117,N_7999,N_7990);
or U8118 (N_8118,N_7933,N_7936);
nor U8119 (N_8119,N_7881,N_7938);
nor U8120 (N_8120,N_7859,N_7980);
and U8121 (N_8121,N_7967,N_7949);
and U8122 (N_8122,N_7861,N_7828);
and U8123 (N_8123,N_7967,N_7940);
and U8124 (N_8124,N_7935,N_7920);
and U8125 (N_8125,N_7805,N_7967);
nor U8126 (N_8126,N_7944,N_7846);
or U8127 (N_8127,N_7954,N_7875);
and U8128 (N_8128,N_7858,N_7809);
nand U8129 (N_8129,N_7877,N_7923);
nor U8130 (N_8130,N_7892,N_7982);
or U8131 (N_8131,N_7954,N_7932);
or U8132 (N_8132,N_7850,N_7847);
nand U8133 (N_8133,N_7955,N_7924);
and U8134 (N_8134,N_7899,N_7809);
nor U8135 (N_8135,N_7961,N_7921);
or U8136 (N_8136,N_7946,N_7872);
nor U8137 (N_8137,N_7830,N_7816);
and U8138 (N_8138,N_7801,N_7904);
or U8139 (N_8139,N_7936,N_7973);
or U8140 (N_8140,N_7973,N_7883);
nor U8141 (N_8141,N_7808,N_7835);
and U8142 (N_8142,N_7906,N_7888);
nor U8143 (N_8143,N_7871,N_7810);
nand U8144 (N_8144,N_7986,N_7865);
xnor U8145 (N_8145,N_7854,N_7996);
nand U8146 (N_8146,N_7858,N_7925);
nand U8147 (N_8147,N_7830,N_7941);
and U8148 (N_8148,N_7922,N_7814);
nand U8149 (N_8149,N_7919,N_7852);
nor U8150 (N_8150,N_7804,N_7945);
xnor U8151 (N_8151,N_7959,N_7998);
nand U8152 (N_8152,N_7857,N_7903);
nand U8153 (N_8153,N_7961,N_7844);
and U8154 (N_8154,N_7806,N_7832);
nand U8155 (N_8155,N_7862,N_7861);
nand U8156 (N_8156,N_7817,N_7853);
or U8157 (N_8157,N_7992,N_7814);
nand U8158 (N_8158,N_7939,N_7873);
and U8159 (N_8159,N_7906,N_7823);
nand U8160 (N_8160,N_7995,N_7820);
nor U8161 (N_8161,N_7867,N_7992);
nor U8162 (N_8162,N_7834,N_7809);
or U8163 (N_8163,N_7967,N_7900);
and U8164 (N_8164,N_7828,N_7940);
and U8165 (N_8165,N_7827,N_7802);
and U8166 (N_8166,N_7826,N_7960);
or U8167 (N_8167,N_7984,N_7940);
or U8168 (N_8168,N_7921,N_7967);
xor U8169 (N_8169,N_7850,N_7862);
or U8170 (N_8170,N_7956,N_7856);
nand U8171 (N_8171,N_7980,N_7983);
nand U8172 (N_8172,N_7896,N_7959);
nand U8173 (N_8173,N_7931,N_7848);
xor U8174 (N_8174,N_7984,N_7943);
or U8175 (N_8175,N_7901,N_7948);
or U8176 (N_8176,N_7986,N_7825);
or U8177 (N_8177,N_7927,N_7892);
and U8178 (N_8178,N_7840,N_7801);
nand U8179 (N_8179,N_7979,N_7976);
nand U8180 (N_8180,N_7827,N_7844);
nor U8181 (N_8181,N_7837,N_7958);
nor U8182 (N_8182,N_7887,N_7908);
or U8183 (N_8183,N_7903,N_7901);
or U8184 (N_8184,N_7894,N_7989);
or U8185 (N_8185,N_7892,N_7948);
or U8186 (N_8186,N_7975,N_7859);
and U8187 (N_8187,N_7908,N_7998);
nor U8188 (N_8188,N_7811,N_7876);
and U8189 (N_8189,N_7807,N_7965);
nor U8190 (N_8190,N_7858,N_7907);
nor U8191 (N_8191,N_7841,N_7819);
and U8192 (N_8192,N_7802,N_7935);
and U8193 (N_8193,N_7870,N_7800);
nand U8194 (N_8194,N_7867,N_7864);
and U8195 (N_8195,N_7945,N_7923);
nand U8196 (N_8196,N_7975,N_7965);
nor U8197 (N_8197,N_7927,N_7884);
nor U8198 (N_8198,N_7950,N_7827);
nand U8199 (N_8199,N_7976,N_7820);
or U8200 (N_8200,N_8158,N_8098);
nand U8201 (N_8201,N_8119,N_8066);
and U8202 (N_8202,N_8029,N_8062);
nor U8203 (N_8203,N_8072,N_8190);
xor U8204 (N_8204,N_8179,N_8199);
nor U8205 (N_8205,N_8183,N_8165);
xnor U8206 (N_8206,N_8016,N_8111);
or U8207 (N_8207,N_8030,N_8055);
nor U8208 (N_8208,N_8083,N_8163);
nand U8209 (N_8209,N_8189,N_8151);
nor U8210 (N_8210,N_8156,N_8187);
nand U8211 (N_8211,N_8037,N_8079);
or U8212 (N_8212,N_8057,N_8000);
and U8213 (N_8213,N_8121,N_8112);
nor U8214 (N_8214,N_8070,N_8047);
nor U8215 (N_8215,N_8039,N_8193);
and U8216 (N_8216,N_8097,N_8052);
nor U8217 (N_8217,N_8049,N_8050);
and U8218 (N_8218,N_8136,N_8195);
nand U8219 (N_8219,N_8006,N_8056);
xnor U8220 (N_8220,N_8027,N_8007);
nand U8221 (N_8221,N_8107,N_8146);
nand U8222 (N_8222,N_8142,N_8101);
and U8223 (N_8223,N_8108,N_8078);
nand U8224 (N_8224,N_8105,N_8024);
nor U8225 (N_8225,N_8026,N_8003);
nand U8226 (N_8226,N_8014,N_8133);
or U8227 (N_8227,N_8095,N_8035);
nand U8228 (N_8228,N_8086,N_8106);
nand U8229 (N_8229,N_8167,N_8162);
and U8230 (N_8230,N_8140,N_8011);
nor U8231 (N_8231,N_8132,N_8071);
nand U8232 (N_8232,N_8082,N_8090);
and U8233 (N_8233,N_8170,N_8012);
nor U8234 (N_8234,N_8021,N_8164);
xnor U8235 (N_8235,N_8064,N_8159);
nand U8236 (N_8236,N_8010,N_8061);
or U8237 (N_8237,N_8185,N_8131);
nor U8238 (N_8238,N_8194,N_8143);
or U8239 (N_8239,N_8096,N_8155);
or U8240 (N_8240,N_8019,N_8102);
or U8241 (N_8241,N_8113,N_8045);
or U8242 (N_8242,N_8174,N_8104);
nor U8243 (N_8243,N_8139,N_8171);
nor U8244 (N_8244,N_8188,N_8022);
nand U8245 (N_8245,N_8196,N_8161);
nor U8246 (N_8246,N_8128,N_8089);
nor U8247 (N_8247,N_8100,N_8028);
and U8248 (N_8248,N_8127,N_8123);
nor U8249 (N_8249,N_8120,N_8150);
or U8250 (N_8250,N_8130,N_8075);
and U8251 (N_8251,N_8059,N_8002);
and U8252 (N_8252,N_8129,N_8152);
nand U8253 (N_8253,N_8177,N_8192);
or U8254 (N_8254,N_8091,N_8160);
nor U8255 (N_8255,N_8042,N_8141);
and U8256 (N_8256,N_8099,N_8168);
nor U8257 (N_8257,N_8001,N_8068);
or U8258 (N_8258,N_8043,N_8038);
nand U8259 (N_8259,N_8060,N_8125);
nor U8260 (N_8260,N_8145,N_8053);
and U8261 (N_8261,N_8094,N_8109);
nand U8262 (N_8262,N_8184,N_8093);
or U8263 (N_8263,N_8173,N_8025);
or U8264 (N_8264,N_8138,N_8054);
nand U8265 (N_8265,N_8137,N_8069);
or U8266 (N_8266,N_8110,N_8081);
nand U8267 (N_8267,N_8077,N_8046);
or U8268 (N_8268,N_8122,N_8087);
nand U8269 (N_8269,N_8124,N_8153);
or U8270 (N_8270,N_8033,N_8048);
nor U8271 (N_8271,N_8017,N_8197);
nand U8272 (N_8272,N_8041,N_8181);
and U8273 (N_8273,N_8015,N_8009);
and U8274 (N_8274,N_8013,N_8115);
nor U8275 (N_8275,N_8116,N_8076);
nand U8276 (N_8276,N_8080,N_8065);
or U8277 (N_8277,N_8023,N_8018);
nor U8278 (N_8278,N_8117,N_8126);
and U8279 (N_8279,N_8074,N_8147);
and U8280 (N_8280,N_8044,N_8198);
nand U8281 (N_8281,N_8180,N_8051);
nand U8282 (N_8282,N_8135,N_8118);
nand U8283 (N_8283,N_8114,N_8172);
and U8284 (N_8284,N_8008,N_8166);
and U8285 (N_8285,N_8182,N_8134);
nand U8286 (N_8286,N_8088,N_8175);
and U8287 (N_8287,N_8032,N_8157);
or U8288 (N_8288,N_8005,N_8063);
or U8289 (N_8289,N_8031,N_8186);
or U8290 (N_8290,N_8178,N_8169);
nor U8291 (N_8291,N_8034,N_8084);
nor U8292 (N_8292,N_8176,N_8149);
nand U8293 (N_8293,N_8040,N_8092);
nand U8294 (N_8294,N_8191,N_8073);
xnor U8295 (N_8295,N_8144,N_8058);
or U8296 (N_8296,N_8085,N_8036);
xnor U8297 (N_8297,N_8020,N_8148);
nand U8298 (N_8298,N_8067,N_8004);
and U8299 (N_8299,N_8154,N_8103);
nand U8300 (N_8300,N_8172,N_8115);
nor U8301 (N_8301,N_8145,N_8013);
or U8302 (N_8302,N_8037,N_8031);
and U8303 (N_8303,N_8128,N_8018);
and U8304 (N_8304,N_8132,N_8172);
and U8305 (N_8305,N_8195,N_8058);
nand U8306 (N_8306,N_8155,N_8049);
or U8307 (N_8307,N_8044,N_8131);
and U8308 (N_8308,N_8148,N_8184);
nand U8309 (N_8309,N_8073,N_8027);
xor U8310 (N_8310,N_8162,N_8135);
nand U8311 (N_8311,N_8163,N_8169);
nand U8312 (N_8312,N_8002,N_8181);
and U8313 (N_8313,N_8004,N_8033);
nor U8314 (N_8314,N_8198,N_8063);
and U8315 (N_8315,N_8036,N_8044);
nand U8316 (N_8316,N_8048,N_8042);
or U8317 (N_8317,N_8153,N_8187);
nand U8318 (N_8318,N_8059,N_8024);
and U8319 (N_8319,N_8040,N_8149);
xor U8320 (N_8320,N_8167,N_8198);
or U8321 (N_8321,N_8132,N_8061);
nand U8322 (N_8322,N_8001,N_8095);
or U8323 (N_8323,N_8136,N_8060);
and U8324 (N_8324,N_8169,N_8160);
nand U8325 (N_8325,N_8183,N_8058);
and U8326 (N_8326,N_8171,N_8115);
or U8327 (N_8327,N_8024,N_8080);
or U8328 (N_8328,N_8027,N_8174);
and U8329 (N_8329,N_8023,N_8050);
and U8330 (N_8330,N_8080,N_8197);
or U8331 (N_8331,N_8007,N_8029);
nand U8332 (N_8332,N_8002,N_8035);
and U8333 (N_8333,N_8121,N_8088);
and U8334 (N_8334,N_8160,N_8147);
nor U8335 (N_8335,N_8157,N_8156);
or U8336 (N_8336,N_8143,N_8122);
and U8337 (N_8337,N_8028,N_8030);
or U8338 (N_8338,N_8037,N_8178);
nand U8339 (N_8339,N_8114,N_8005);
and U8340 (N_8340,N_8082,N_8155);
nand U8341 (N_8341,N_8166,N_8055);
and U8342 (N_8342,N_8041,N_8150);
or U8343 (N_8343,N_8109,N_8147);
nor U8344 (N_8344,N_8150,N_8013);
and U8345 (N_8345,N_8025,N_8169);
nor U8346 (N_8346,N_8138,N_8059);
and U8347 (N_8347,N_8035,N_8123);
nor U8348 (N_8348,N_8138,N_8053);
xnor U8349 (N_8349,N_8066,N_8198);
nor U8350 (N_8350,N_8045,N_8049);
or U8351 (N_8351,N_8118,N_8087);
nand U8352 (N_8352,N_8132,N_8052);
nand U8353 (N_8353,N_8091,N_8049);
or U8354 (N_8354,N_8150,N_8040);
nor U8355 (N_8355,N_8186,N_8009);
or U8356 (N_8356,N_8140,N_8088);
nand U8357 (N_8357,N_8199,N_8006);
and U8358 (N_8358,N_8127,N_8070);
nor U8359 (N_8359,N_8171,N_8151);
or U8360 (N_8360,N_8175,N_8152);
and U8361 (N_8361,N_8168,N_8116);
nand U8362 (N_8362,N_8033,N_8120);
nand U8363 (N_8363,N_8163,N_8034);
or U8364 (N_8364,N_8027,N_8097);
nand U8365 (N_8365,N_8014,N_8152);
nor U8366 (N_8366,N_8036,N_8020);
nand U8367 (N_8367,N_8017,N_8122);
or U8368 (N_8368,N_8027,N_8004);
xor U8369 (N_8369,N_8146,N_8151);
nor U8370 (N_8370,N_8160,N_8053);
or U8371 (N_8371,N_8091,N_8080);
nor U8372 (N_8372,N_8123,N_8139);
or U8373 (N_8373,N_8160,N_8063);
or U8374 (N_8374,N_8130,N_8072);
nand U8375 (N_8375,N_8110,N_8176);
and U8376 (N_8376,N_8112,N_8026);
and U8377 (N_8377,N_8067,N_8192);
and U8378 (N_8378,N_8116,N_8124);
xor U8379 (N_8379,N_8194,N_8080);
nand U8380 (N_8380,N_8029,N_8161);
xor U8381 (N_8381,N_8127,N_8055);
and U8382 (N_8382,N_8032,N_8033);
and U8383 (N_8383,N_8008,N_8187);
xor U8384 (N_8384,N_8162,N_8149);
and U8385 (N_8385,N_8178,N_8014);
or U8386 (N_8386,N_8175,N_8094);
nor U8387 (N_8387,N_8147,N_8190);
and U8388 (N_8388,N_8006,N_8130);
and U8389 (N_8389,N_8023,N_8074);
nor U8390 (N_8390,N_8024,N_8017);
or U8391 (N_8391,N_8112,N_8173);
or U8392 (N_8392,N_8137,N_8064);
and U8393 (N_8393,N_8190,N_8114);
or U8394 (N_8394,N_8197,N_8171);
nor U8395 (N_8395,N_8122,N_8068);
nand U8396 (N_8396,N_8165,N_8119);
nor U8397 (N_8397,N_8098,N_8057);
nor U8398 (N_8398,N_8066,N_8188);
nor U8399 (N_8399,N_8027,N_8137);
nand U8400 (N_8400,N_8236,N_8227);
or U8401 (N_8401,N_8372,N_8315);
nand U8402 (N_8402,N_8222,N_8391);
and U8403 (N_8403,N_8240,N_8316);
or U8404 (N_8404,N_8229,N_8368);
nor U8405 (N_8405,N_8201,N_8378);
or U8406 (N_8406,N_8328,N_8350);
nand U8407 (N_8407,N_8209,N_8273);
nand U8408 (N_8408,N_8320,N_8253);
nor U8409 (N_8409,N_8305,N_8294);
or U8410 (N_8410,N_8348,N_8323);
nand U8411 (N_8411,N_8367,N_8302);
and U8412 (N_8412,N_8314,N_8325);
nor U8413 (N_8413,N_8351,N_8220);
nand U8414 (N_8414,N_8341,N_8363);
nand U8415 (N_8415,N_8242,N_8382);
nand U8416 (N_8416,N_8286,N_8274);
nor U8417 (N_8417,N_8376,N_8386);
nand U8418 (N_8418,N_8297,N_8381);
nor U8419 (N_8419,N_8392,N_8241);
nor U8420 (N_8420,N_8203,N_8244);
nand U8421 (N_8421,N_8364,N_8313);
nor U8422 (N_8422,N_8276,N_8279);
nor U8423 (N_8423,N_8280,N_8358);
nor U8424 (N_8424,N_8272,N_8377);
nand U8425 (N_8425,N_8398,N_8349);
or U8426 (N_8426,N_8371,N_8357);
nor U8427 (N_8427,N_8344,N_8234);
and U8428 (N_8428,N_8265,N_8275);
nor U8429 (N_8429,N_8232,N_8206);
and U8430 (N_8430,N_8231,N_8204);
nor U8431 (N_8431,N_8311,N_8246);
or U8432 (N_8432,N_8293,N_8312);
nand U8433 (N_8433,N_8214,N_8385);
nand U8434 (N_8434,N_8202,N_8396);
or U8435 (N_8435,N_8249,N_8251);
nand U8436 (N_8436,N_8250,N_8223);
nand U8437 (N_8437,N_8333,N_8205);
nor U8438 (N_8438,N_8211,N_8221);
or U8439 (N_8439,N_8365,N_8281);
nand U8440 (N_8440,N_8379,N_8285);
or U8441 (N_8441,N_8224,N_8258);
nand U8442 (N_8442,N_8208,N_8268);
nand U8443 (N_8443,N_8387,N_8375);
xnor U8444 (N_8444,N_8207,N_8388);
or U8445 (N_8445,N_8322,N_8393);
or U8446 (N_8446,N_8394,N_8257);
nand U8447 (N_8447,N_8370,N_8233);
and U8448 (N_8448,N_8299,N_8395);
and U8449 (N_8449,N_8304,N_8254);
and U8450 (N_8450,N_8342,N_8327);
or U8451 (N_8451,N_8397,N_8213);
and U8452 (N_8452,N_8219,N_8271);
and U8453 (N_8453,N_8252,N_8324);
or U8454 (N_8454,N_8248,N_8200);
nand U8455 (N_8455,N_8340,N_8239);
or U8456 (N_8456,N_8331,N_8283);
nand U8457 (N_8457,N_8326,N_8303);
and U8458 (N_8458,N_8212,N_8354);
nor U8459 (N_8459,N_8347,N_8278);
nand U8460 (N_8460,N_8332,N_8338);
and U8461 (N_8461,N_8399,N_8277);
nor U8462 (N_8462,N_8366,N_8245);
nor U8463 (N_8463,N_8295,N_8330);
nor U8464 (N_8464,N_8261,N_8390);
or U8465 (N_8465,N_8355,N_8290);
or U8466 (N_8466,N_8215,N_8260);
or U8467 (N_8467,N_8292,N_8237);
nand U8468 (N_8468,N_8243,N_8334);
nand U8469 (N_8469,N_8306,N_8345);
or U8470 (N_8470,N_8238,N_8289);
nand U8471 (N_8471,N_8317,N_8301);
or U8472 (N_8472,N_8337,N_8373);
or U8473 (N_8473,N_8335,N_8266);
or U8474 (N_8474,N_8339,N_8288);
nor U8475 (N_8475,N_8318,N_8346);
and U8476 (N_8476,N_8356,N_8291);
or U8477 (N_8477,N_8307,N_8296);
nor U8478 (N_8478,N_8380,N_8263);
or U8479 (N_8479,N_8230,N_8269);
and U8480 (N_8480,N_8308,N_8321);
and U8481 (N_8481,N_8247,N_8352);
and U8482 (N_8482,N_8369,N_8359);
and U8483 (N_8483,N_8256,N_8343);
and U8484 (N_8484,N_8298,N_8300);
or U8485 (N_8485,N_8262,N_8216);
and U8486 (N_8486,N_8255,N_8267);
or U8487 (N_8487,N_8228,N_8310);
or U8488 (N_8488,N_8284,N_8210);
and U8489 (N_8489,N_8384,N_8383);
nand U8490 (N_8490,N_8336,N_8329);
and U8491 (N_8491,N_8360,N_8374);
xnor U8492 (N_8492,N_8319,N_8361);
nand U8493 (N_8493,N_8225,N_8353);
nor U8494 (N_8494,N_8389,N_8226);
or U8495 (N_8495,N_8259,N_8309);
or U8496 (N_8496,N_8270,N_8287);
or U8497 (N_8497,N_8282,N_8217);
or U8498 (N_8498,N_8235,N_8264);
nor U8499 (N_8499,N_8362,N_8218);
nand U8500 (N_8500,N_8298,N_8383);
or U8501 (N_8501,N_8248,N_8307);
or U8502 (N_8502,N_8385,N_8305);
nand U8503 (N_8503,N_8302,N_8279);
nor U8504 (N_8504,N_8318,N_8293);
and U8505 (N_8505,N_8298,N_8317);
nor U8506 (N_8506,N_8277,N_8246);
or U8507 (N_8507,N_8222,N_8246);
and U8508 (N_8508,N_8361,N_8286);
or U8509 (N_8509,N_8260,N_8207);
or U8510 (N_8510,N_8268,N_8331);
nor U8511 (N_8511,N_8368,N_8349);
or U8512 (N_8512,N_8336,N_8360);
or U8513 (N_8513,N_8305,N_8323);
nand U8514 (N_8514,N_8399,N_8269);
nor U8515 (N_8515,N_8295,N_8309);
nand U8516 (N_8516,N_8330,N_8252);
or U8517 (N_8517,N_8220,N_8316);
or U8518 (N_8518,N_8335,N_8387);
or U8519 (N_8519,N_8340,N_8209);
or U8520 (N_8520,N_8238,N_8364);
or U8521 (N_8521,N_8246,N_8212);
or U8522 (N_8522,N_8272,N_8353);
nor U8523 (N_8523,N_8315,N_8210);
or U8524 (N_8524,N_8316,N_8217);
or U8525 (N_8525,N_8221,N_8324);
and U8526 (N_8526,N_8241,N_8268);
nand U8527 (N_8527,N_8343,N_8349);
nand U8528 (N_8528,N_8392,N_8200);
and U8529 (N_8529,N_8386,N_8285);
or U8530 (N_8530,N_8271,N_8233);
nand U8531 (N_8531,N_8348,N_8336);
and U8532 (N_8532,N_8386,N_8332);
and U8533 (N_8533,N_8231,N_8396);
nand U8534 (N_8534,N_8258,N_8285);
or U8535 (N_8535,N_8222,N_8226);
nand U8536 (N_8536,N_8204,N_8235);
or U8537 (N_8537,N_8295,N_8340);
or U8538 (N_8538,N_8321,N_8326);
and U8539 (N_8539,N_8256,N_8398);
and U8540 (N_8540,N_8200,N_8388);
nor U8541 (N_8541,N_8233,N_8393);
and U8542 (N_8542,N_8282,N_8398);
or U8543 (N_8543,N_8267,N_8329);
nand U8544 (N_8544,N_8243,N_8322);
nand U8545 (N_8545,N_8235,N_8381);
and U8546 (N_8546,N_8230,N_8244);
or U8547 (N_8547,N_8345,N_8341);
nand U8548 (N_8548,N_8332,N_8272);
nor U8549 (N_8549,N_8313,N_8274);
and U8550 (N_8550,N_8374,N_8352);
or U8551 (N_8551,N_8258,N_8326);
and U8552 (N_8552,N_8361,N_8234);
nor U8553 (N_8553,N_8389,N_8377);
or U8554 (N_8554,N_8264,N_8394);
or U8555 (N_8555,N_8244,N_8360);
nor U8556 (N_8556,N_8351,N_8213);
nor U8557 (N_8557,N_8365,N_8388);
nand U8558 (N_8558,N_8379,N_8263);
nand U8559 (N_8559,N_8348,N_8207);
and U8560 (N_8560,N_8205,N_8358);
and U8561 (N_8561,N_8285,N_8358);
or U8562 (N_8562,N_8284,N_8387);
or U8563 (N_8563,N_8214,N_8375);
or U8564 (N_8564,N_8267,N_8397);
nor U8565 (N_8565,N_8339,N_8245);
and U8566 (N_8566,N_8344,N_8322);
and U8567 (N_8567,N_8332,N_8249);
and U8568 (N_8568,N_8216,N_8351);
xnor U8569 (N_8569,N_8329,N_8307);
or U8570 (N_8570,N_8376,N_8377);
or U8571 (N_8571,N_8270,N_8257);
and U8572 (N_8572,N_8281,N_8339);
nor U8573 (N_8573,N_8221,N_8267);
or U8574 (N_8574,N_8270,N_8334);
and U8575 (N_8575,N_8331,N_8379);
or U8576 (N_8576,N_8353,N_8274);
xor U8577 (N_8577,N_8307,N_8392);
nand U8578 (N_8578,N_8399,N_8356);
nand U8579 (N_8579,N_8313,N_8251);
nor U8580 (N_8580,N_8321,N_8333);
nand U8581 (N_8581,N_8264,N_8367);
and U8582 (N_8582,N_8387,N_8241);
nor U8583 (N_8583,N_8330,N_8374);
or U8584 (N_8584,N_8256,N_8359);
nand U8585 (N_8585,N_8223,N_8303);
xnor U8586 (N_8586,N_8233,N_8301);
nand U8587 (N_8587,N_8363,N_8309);
and U8588 (N_8588,N_8320,N_8351);
or U8589 (N_8589,N_8395,N_8309);
and U8590 (N_8590,N_8247,N_8290);
nand U8591 (N_8591,N_8359,N_8226);
or U8592 (N_8592,N_8294,N_8391);
or U8593 (N_8593,N_8360,N_8362);
and U8594 (N_8594,N_8287,N_8316);
nand U8595 (N_8595,N_8372,N_8209);
and U8596 (N_8596,N_8263,N_8252);
and U8597 (N_8597,N_8393,N_8328);
or U8598 (N_8598,N_8222,N_8244);
or U8599 (N_8599,N_8319,N_8373);
or U8600 (N_8600,N_8412,N_8529);
and U8601 (N_8601,N_8509,N_8592);
nor U8602 (N_8602,N_8425,N_8515);
nor U8603 (N_8603,N_8462,N_8586);
or U8604 (N_8604,N_8476,N_8545);
nor U8605 (N_8605,N_8418,N_8439);
nor U8606 (N_8606,N_8491,N_8402);
nor U8607 (N_8607,N_8411,N_8488);
nand U8608 (N_8608,N_8578,N_8449);
nor U8609 (N_8609,N_8516,N_8557);
or U8610 (N_8610,N_8581,N_8489);
and U8611 (N_8611,N_8480,N_8599);
and U8612 (N_8612,N_8558,N_8417);
or U8613 (N_8613,N_8421,N_8452);
nand U8614 (N_8614,N_8467,N_8466);
and U8615 (N_8615,N_8503,N_8526);
and U8616 (N_8616,N_8584,N_8474);
nor U8617 (N_8617,N_8546,N_8431);
or U8618 (N_8618,N_8541,N_8407);
or U8619 (N_8619,N_8475,N_8420);
and U8620 (N_8620,N_8519,N_8443);
and U8621 (N_8621,N_8543,N_8561);
or U8622 (N_8622,N_8571,N_8448);
nor U8623 (N_8623,N_8442,N_8416);
nand U8624 (N_8624,N_8446,N_8508);
xor U8625 (N_8625,N_8424,N_8595);
and U8626 (N_8626,N_8485,N_8594);
or U8627 (N_8627,N_8512,N_8479);
or U8628 (N_8628,N_8441,N_8413);
nand U8629 (N_8629,N_8538,N_8477);
nand U8630 (N_8630,N_8597,N_8497);
nor U8631 (N_8631,N_8401,N_8569);
and U8632 (N_8632,N_8455,N_8481);
and U8633 (N_8633,N_8579,N_8560);
or U8634 (N_8634,N_8428,N_8507);
or U8635 (N_8635,N_8457,N_8494);
nor U8636 (N_8636,N_8473,N_8451);
nor U8637 (N_8637,N_8499,N_8582);
nor U8638 (N_8638,N_8530,N_8565);
nand U8639 (N_8639,N_8570,N_8486);
xnor U8640 (N_8640,N_8589,N_8470);
nand U8641 (N_8641,N_8534,N_8506);
and U8642 (N_8642,N_8437,N_8504);
and U8643 (N_8643,N_8400,N_8495);
and U8644 (N_8644,N_8572,N_8568);
or U8645 (N_8645,N_8583,N_8542);
and U8646 (N_8646,N_8454,N_8461);
and U8647 (N_8647,N_8426,N_8471);
and U8648 (N_8648,N_8410,N_8520);
nand U8649 (N_8649,N_8478,N_8422);
and U8650 (N_8650,N_8405,N_8434);
and U8651 (N_8651,N_8567,N_8464);
or U8652 (N_8652,N_8468,N_8593);
and U8653 (N_8653,N_8552,N_8587);
or U8654 (N_8654,N_8414,N_8450);
nand U8655 (N_8655,N_8433,N_8563);
nor U8656 (N_8656,N_8566,N_8493);
nor U8657 (N_8657,N_8596,N_8460);
and U8658 (N_8658,N_8598,N_8456);
or U8659 (N_8659,N_8531,N_8429);
nor U8660 (N_8660,N_8430,N_8528);
or U8661 (N_8661,N_8403,N_8440);
and U8662 (N_8662,N_8463,N_8532);
nor U8663 (N_8663,N_8436,N_8573);
nand U8664 (N_8664,N_8524,N_8444);
and U8665 (N_8665,N_8537,N_8585);
nand U8666 (N_8666,N_8547,N_8591);
nor U8667 (N_8667,N_8510,N_8408);
xor U8668 (N_8668,N_8551,N_8580);
nor U8669 (N_8669,N_8555,N_8590);
nor U8670 (N_8670,N_8423,N_8458);
or U8671 (N_8671,N_8501,N_8505);
nor U8672 (N_8672,N_8406,N_8535);
nand U8673 (N_8673,N_8518,N_8484);
nand U8674 (N_8674,N_8554,N_8523);
and U8675 (N_8675,N_8522,N_8559);
nor U8676 (N_8676,N_8472,N_8577);
nand U8677 (N_8677,N_8548,N_8540);
nor U8678 (N_8678,N_8438,N_8482);
and U8679 (N_8679,N_8483,N_8500);
and U8680 (N_8680,N_8447,N_8574);
or U8681 (N_8681,N_8588,N_8576);
and U8682 (N_8682,N_8511,N_8453);
nand U8683 (N_8683,N_8487,N_8432);
and U8684 (N_8684,N_8490,N_8492);
and U8685 (N_8685,N_8496,N_8435);
or U8686 (N_8686,N_8459,N_8498);
nand U8687 (N_8687,N_8539,N_8521);
or U8688 (N_8688,N_8575,N_8514);
nand U8689 (N_8689,N_8419,N_8404);
and U8690 (N_8690,N_8527,N_8533);
nor U8691 (N_8691,N_8549,N_8445);
and U8692 (N_8692,N_8562,N_8513);
nor U8693 (N_8693,N_8415,N_8550);
or U8694 (N_8694,N_8556,N_8427);
nor U8695 (N_8695,N_8536,N_8409);
xor U8696 (N_8696,N_8553,N_8502);
and U8697 (N_8697,N_8525,N_8544);
nand U8698 (N_8698,N_8469,N_8465);
nor U8699 (N_8699,N_8564,N_8517);
nor U8700 (N_8700,N_8583,N_8487);
nand U8701 (N_8701,N_8441,N_8520);
nor U8702 (N_8702,N_8570,N_8585);
and U8703 (N_8703,N_8463,N_8405);
and U8704 (N_8704,N_8563,N_8589);
or U8705 (N_8705,N_8411,N_8479);
or U8706 (N_8706,N_8433,N_8489);
xnor U8707 (N_8707,N_8460,N_8534);
or U8708 (N_8708,N_8561,N_8562);
or U8709 (N_8709,N_8487,N_8594);
nand U8710 (N_8710,N_8553,N_8404);
nand U8711 (N_8711,N_8593,N_8583);
and U8712 (N_8712,N_8527,N_8414);
nor U8713 (N_8713,N_8584,N_8488);
or U8714 (N_8714,N_8422,N_8433);
nand U8715 (N_8715,N_8444,N_8474);
and U8716 (N_8716,N_8583,N_8539);
or U8717 (N_8717,N_8463,N_8444);
and U8718 (N_8718,N_8571,N_8526);
or U8719 (N_8719,N_8581,N_8450);
and U8720 (N_8720,N_8407,N_8422);
nand U8721 (N_8721,N_8459,N_8456);
and U8722 (N_8722,N_8447,N_8545);
and U8723 (N_8723,N_8463,N_8456);
nor U8724 (N_8724,N_8430,N_8405);
or U8725 (N_8725,N_8443,N_8538);
nor U8726 (N_8726,N_8557,N_8507);
xnor U8727 (N_8727,N_8588,N_8520);
and U8728 (N_8728,N_8580,N_8404);
and U8729 (N_8729,N_8513,N_8483);
and U8730 (N_8730,N_8599,N_8592);
or U8731 (N_8731,N_8554,N_8436);
nor U8732 (N_8732,N_8576,N_8426);
or U8733 (N_8733,N_8418,N_8522);
or U8734 (N_8734,N_8465,N_8517);
nor U8735 (N_8735,N_8582,N_8482);
nand U8736 (N_8736,N_8411,N_8487);
xor U8737 (N_8737,N_8587,N_8503);
and U8738 (N_8738,N_8506,N_8532);
or U8739 (N_8739,N_8553,N_8401);
and U8740 (N_8740,N_8586,N_8558);
or U8741 (N_8741,N_8442,N_8578);
and U8742 (N_8742,N_8472,N_8557);
or U8743 (N_8743,N_8421,N_8519);
or U8744 (N_8744,N_8478,N_8530);
and U8745 (N_8745,N_8549,N_8468);
or U8746 (N_8746,N_8501,N_8553);
or U8747 (N_8747,N_8590,N_8548);
nor U8748 (N_8748,N_8509,N_8449);
and U8749 (N_8749,N_8572,N_8503);
nand U8750 (N_8750,N_8471,N_8465);
nor U8751 (N_8751,N_8457,N_8478);
nand U8752 (N_8752,N_8452,N_8410);
and U8753 (N_8753,N_8460,N_8430);
and U8754 (N_8754,N_8534,N_8555);
nand U8755 (N_8755,N_8477,N_8589);
nor U8756 (N_8756,N_8510,N_8502);
xnor U8757 (N_8757,N_8514,N_8540);
nand U8758 (N_8758,N_8507,N_8577);
or U8759 (N_8759,N_8468,N_8464);
nor U8760 (N_8760,N_8401,N_8583);
nor U8761 (N_8761,N_8427,N_8408);
nand U8762 (N_8762,N_8453,N_8509);
or U8763 (N_8763,N_8497,N_8583);
nand U8764 (N_8764,N_8462,N_8411);
nand U8765 (N_8765,N_8446,N_8471);
or U8766 (N_8766,N_8432,N_8585);
or U8767 (N_8767,N_8560,N_8587);
nor U8768 (N_8768,N_8563,N_8497);
nor U8769 (N_8769,N_8533,N_8407);
nand U8770 (N_8770,N_8483,N_8581);
or U8771 (N_8771,N_8594,N_8591);
nor U8772 (N_8772,N_8512,N_8469);
or U8773 (N_8773,N_8593,N_8427);
nor U8774 (N_8774,N_8462,N_8454);
or U8775 (N_8775,N_8552,N_8500);
nand U8776 (N_8776,N_8410,N_8575);
nand U8777 (N_8777,N_8499,N_8469);
xnor U8778 (N_8778,N_8502,N_8507);
and U8779 (N_8779,N_8522,N_8557);
xnor U8780 (N_8780,N_8593,N_8592);
nor U8781 (N_8781,N_8482,N_8424);
and U8782 (N_8782,N_8528,N_8537);
and U8783 (N_8783,N_8489,N_8446);
nand U8784 (N_8784,N_8490,N_8469);
and U8785 (N_8785,N_8403,N_8470);
nor U8786 (N_8786,N_8442,N_8577);
nand U8787 (N_8787,N_8453,N_8494);
nor U8788 (N_8788,N_8519,N_8459);
nand U8789 (N_8789,N_8408,N_8582);
nor U8790 (N_8790,N_8424,N_8407);
or U8791 (N_8791,N_8505,N_8538);
nor U8792 (N_8792,N_8496,N_8459);
nor U8793 (N_8793,N_8467,N_8576);
nand U8794 (N_8794,N_8413,N_8488);
nand U8795 (N_8795,N_8483,N_8479);
or U8796 (N_8796,N_8404,N_8416);
nand U8797 (N_8797,N_8557,N_8532);
nand U8798 (N_8798,N_8409,N_8484);
and U8799 (N_8799,N_8563,N_8495);
and U8800 (N_8800,N_8737,N_8640);
and U8801 (N_8801,N_8632,N_8783);
or U8802 (N_8802,N_8774,N_8793);
and U8803 (N_8803,N_8655,N_8784);
nand U8804 (N_8804,N_8795,N_8671);
or U8805 (N_8805,N_8647,N_8704);
nand U8806 (N_8806,N_8615,N_8780);
or U8807 (N_8807,N_8680,N_8638);
or U8808 (N_8808,N_8715,N_8688);
nand U8809 (N_8809,N_8686,N_8631);
or U8810 (N_8810,N_8687,N_8781);
nand U8811 (N_8811,N_8667,N_8726);
nand U8812 (N_8812,N_8619,N_8603);
or U8813 (N_8813,N_8744,N_8718);
or U8814 (N_8814,N_8728,N_8751);
nand U8815 (N_8815,N_8652,N_8646);
nor U8816 (N_8816,N_8643,N_8653);
and U8817 (N_8817,N_8636,N_8778);
and U8818 (N_8818,N_8790,N_8637);
nor U8819 (N_8819,N_8729,N_8607);
and U8820 (N_8820,N_8634,N_8730);
or U8821 (N_8821,N_8714,N_8733);
nor U8822 (N_8822,N_8685,N_8771);
or U8823 (N_8823,N_8734,N_8650);
nor U8824 (N_8824,N_8604,N_8639);
nand U8825 (N_8825,N_8757,N_8738);
and U8826 (N_8826,N_8689,N_8662);
nand U8827 (N_8827,N_8661,N_8775);
nor U8828 (N_8828,N_8788,N_8705);
nand U8829 (N_8829,N_8684,N_8766);
and U8830 (N_8830,N_8796,N_8675);
or U8831 (N_8831,N_8611,N_8747);
nor U8832 (N_8832,N_8679,N_8641);
or U8833 (N_8833,N_8756,N_8697);
or U8834 (N_8834,N_8617,N_8772);
nand U8835 (N_8835,N_8659,N_8713);
or U8836 (N_8836,N_8782,N_8707);
nand U8837 (N_8837,N_8798,N_8703);
or U8838 (N_8838,N_8725,N_8630);
nor U8839 (N_8839,N_8602,N_8765);
or U8840 (N_8840,N_8799,N_8678);
nor U8841 (N_8841,N_8777,N_8609);
nor U8842 (N_8842,N_8700,N_8642);
or U8843 (N_8843,N_8721,N_8649);
or U8844 (N_8844,N_8656,N_8768);
nor U8845 (N_8845,N_8758,N_8690);
nand U8846 (N_8846,N_8746,N_8731);
xnor U8847 (N_8847,N_8742,N_8614);
and U8848 (N_8848,N_8706,N_8691);
nor U8849 (N_8849,N_8717,N_8606);
nor U8850 (N_8850,N_8722,N_8753);
nor U8851 (N_8851,N_8792,N_8754);
nor U8852 (N_8852,N_8702,N_8748);
and U8853 (N_8853,N_8712,N_8767);
or U8854 (N_8854,N_8668,N_8727);
or U8855 (N_8855,N_8769,N_8708);
nand U8856 (N_8856,N_8618,N_8695);
or U8857 (N_8857,N_8786,N_8785);
and U8858 (N_8858,N_8664,N_8683);
and U8859 (N_8859,N_8770,N_8626);
nor U8860 (N_8860,N_8677,N_8791);
or U8861 (N_8861,N_8797,N_8629);
nor U8862 (N_8862,N_8670,N_8622);
nand U8863 (N_8863,N_8660,N_8710);
nand U8864 (N_8864,N_8613,N_8628);
nand U8865 (N_8865,N_8709,N_8635);
nand U8866 (N_8866,N_8681,N_8755);
and U8867 (N_8867,N_8764,N_8610);
nor U8868 (N_8868,N_8720,N_8612);
nand U8869 (N_8869,N_8648,N_8739);
or U8870 (N_8870,N_8787,N_8749);
and U8871 (N_8871,N_8760,N_8724);
and U8872 (N_8872,N_8625,N_8651);
and U8873 (N_8873,N_8608,N_8743);
nand U8874 (N_8874,N_8735,N_8654);
or U8875 (N_8875,N_8669,N_8716);
nand U8876 (N_8876,N_8673,N_8696);
nand U8877 (N_8877,N_8601,N_8741);
or U8878 (N_8878,N_8719,N_8773);
or U8879 (N_8879,N_8657,N_8658);
nand U8880 (N_8880,N_8644,N_8645);
nand U8881 (N_8881,N_8674,N_8605);
xnor U8882 (N_8882,N_8701,N_8676);
and U8883 (N_8883,N_8621,N_8682);
or U8884 (N_8884,N_8763,N_8732);
nor U8885 (N_8885,N_8698,N_8620);
and U8886 (N_8886,N_8736,N_8745);
nand U8887 (N_8887,N_8752,N_8627);
nor U8888 (N_8888,N_8600,N_8794);
or U8889 (N_8889,N_8759,N_8711);
or U8890 (N_8890,N_8663,N_8750);
xor U8891 (N_8891,N_8624,N_8779);
and U8892 (N_8892,N_8776,N_8762);
or U8893 (N_8893,N_8761,N_8666);
or U8894 (N_8894,N_8665,N_8699);
and U8895 (N_8895,N_8672,N_8694);
or U8896 (N_8896,N_8693,N_8789);
nand U8897 (N_8897,N_8723,N_8616);
or U8898 (N_8898,N_8623,N_8740);
nand U8899 (N_8899,N_8692,N_8633);
or U8900 (N_8900,N_8774,N_8635);
nand U8901 (N_8901,N_8628,N_8738);
nand U8902 (N_8902,N_8733,N_8650);
or U8903 (N_8903,N_8600,N_8729);
and U8904 (N_8904,N_8712,N_8737);
or U8905 (N_8905,N_8749,N_8741);
and U8906 (N_8906,N_8693,N_8656);
and U8907 (N_8907,N_8620,N_8728);
nor U8908 (N_8908,N_8722,N_8612);
nand U8909 (N_8909,N_8650,N_8795);
and U8910 (N_8910,N_8645,N_8636);
nand U8911 (N_8911,N_8753,N_8741);
nor U8912 (N_8912,N_8717,N_8615);
nor U8913 (N_8913,N_8746,N_8641);
or U8914 (N_8914,N_8773,N_8734);
nand U8915 (N_8915,N_8713,N_8634);
nand U8916 (N_8916,N_8722,N_8763);
nor U8917 (N_8917,N_8712,N_8659);
or U8918 (N_8918,N_8731,N_8707);
nand U8919 (N_8919,N_8779,N_8620);
and U8920 (N_8920,N_8658,N_8704);
or U8921 (N_8921,N_8778,N_8721);
nor U8922 (N_8922,N_8630,N_8793);
nand U8923 (N_8923,N_8604,N_8756);
nor U8924 (N_8924,N_8648,N_8799);
nand U8925 (N_8925,N_8661,N_8679);
nand U8926 (N_8926,N_8686,N_8754);
and U8927 (N_8927,N_8689,N_8760);
nand U8928 (N_8928,N_8746,N_8791);
or U8929 (N_8929,N_8774,N_8794);
and U8930 (N_8930,N_8738,N_8763);
nor U8931 (N_8931,N_8742,N_8636);
or U8932 (N_8932,N_8649,N_8761);
nand U8933 (N_8933,N_8750,N_8738);
or U8934 (N_8934,N_8738,N_8669);
nand U8935 (N_8935,N_8772,N_8670);
nor U8936 (N_8936,N_8604,N_8730);
or U8937 (N_8937,N_8731,N_8674);
nor U8938 (N_8938,N_8703,N_8627);
and U8939 (N_8939,N_8669,N_8685);
or U8940 (N_8940,N_8718,N_8629);
nand U8941 (N_8941,N_8733,N_8656);
or U8942 (N_8942,N_8678,N_8785);
and U8943 (N_8943,N_8608,N_8712);
or U8944 (N_8944,N_8756,N_8605);
nand U8945 (N_8945,N_8795,N_8657);
nor U8946 (N_8946,N_8761,N_8741);
or U8947 (N_8947,N_8769,N_8653);
nand U8948 (N_8948,N_8663,N_8647);
and U8949 (N_8949,N_8755,N_8645);
and U8950 (N_8950,N_8772,N_8718);
or U8951 (N_8951,N_8651,N_8653);
nand U8952 (N_8952,N_8652,N_8721);
or U8953 (N_8953,N_8660,N_8626);
and U8954 (N_8954,N_8672,N_8788);
or U8955 (N_8955,N_8685,N_8601);
or U8956 (N_8956,N_8662,N_8711);
and U8957 (N_8957,N_8749,N_8746);
and U8958 (N_8958,N_8640,N_8624);
nor U8959 (N_8959,N_8698,N_8689);
or U8960 (N_8960,N_8691,N_8714);
nand U8961 (N_8961,N_8689,N_8737);
nor U8962 (N_8962,N_8746,N_8795);
and U8963 (N_8963,N_8639,N_8606);
or U8964 (N_8964,N_8614,N_8700);
nor U8965 (N_8965,N_8665,N_8680);
and U8966 (N_8966,N_8732,N_8745);
and U8967 (N_8967,N_8612,N_8717);
nor U8968 (N_8968,N_8643,N_8748);
nand U8969 (N_8969,N_8712,N_8730);
or U8970 (N_8970,N_8676,N_8667);
and U8971 (N_8971,N_8716,N_8717);
nand U8972 (N_8972,N_8729,N_8759);
and U8973 (N_8973,N_8641,N_8708);
or U8974 (N_8974,N_8677,N_8678);
and U8975 (N_8975,N_8709,N_8708);
or U8976 (N_8976,N_8604,N_8746);
or U8977 (N_8977,N_8732,N_8706);
or U8978 (N_8978,N_8642,N_8629);
nand U8979 (N_8979,N_8775,N_8638);
and U8980 (N_8980,N_8628,N_8755);
and U8981 (N_8981,N_8635,N_8637);
or U8982 (N_8982,N_8628,N_8601);
or U8983 (N_8983,N_8724,N_8705);
nand U8984 (N_8984,N_8666,N_8773);
or U8985 (N_8985,N_8792,N_8682);
nand U8986 (N_8986,N_8663,N_8713);
nand U8987 (N_8987,N_8727,N_8665);
nand U8988 (N_8988,N_8778,N_8672);
nand U8989 (N_8989,N_8603,N_8687);
nand U8990 (N_8990,N_8781,N_8706);
nand U8991 (N_8991,N_8769,N_8779);
nor U8992 (N_8992,N_8704,N_8600);
nand U8993 (N_8993,N_8716,N_8774);
nand U8994 (N_8994,N_8600,N_8747);
or U8995 (N_8995,N_8713,N_8720);
nor U8996 (N_8996,N_8630,N_8680);
or U8997 (N_8997,N_8770,N_8701);
nor U8998 (N_8998,N_8658,N_8710);
or U8999 (N_8999,N_8732,N_8615);
nand U9000 (N_9000,N_8951,N_8831);
or U9001 (N_9001,N_8892,N_8982);
nand U9002 (N_9002,N_8991,N_8966);
nand U9003 (N_9003,N_8935,N_8849);
and U9004 (N_9004,N_8806,N_8960);
or U9005 (N_9005,N_8927,N_8979);
nand U9006 (N_9006,N_8915,N_8977);
nand U9007 (N_9007,N_8888,N_8906);
or U9008 (N_9008,N_8993,N_8998);
nand U9009 (N_9009,N_8808,N_8872);
nand U9010 (N_9010,N_8859,N_8827);
or U9011 (N_9011,N_8830,N_8968);
or U9012 (N_9012,N_8832,N_8867);
and U9013 (N_9013,N_8976,N_8862);
or U9014 (N_9014,N_8876,N_8852);
or U9015 (N_9015,N_8889,N_8987);
or U9016 (N_9016,N_8962,N_8978);
and U9017 (N_9017,N_8874,N_8890);
nor U9018 (N_9018,N_8948,N_8885);
nand U9019 (N_9019,N_8999,N_8916);
or U9020 (N_9020,N_8802,N_8850);
xnor U9021 (N_9021,N_8924,N_8981);
or U9022 (N_9022,N_8923,N_8946);
and U9023 (N_9023,N_8819,N_8828);
nor U9024 (N_9024,N_8837,N_8917);
nor U9025 (N_9025,N_8818,N_8878);
nand U9026 (N_9026,N_8914,N_8857);
or U9027 (N_9027,N_8980,N_8866);
nor U9028 (N_9028,N_8975,N_8858);
nand U9029 (N_9029,N_8861,N_8825);
and U9030 (N_9030,N_8816,N_8971);
nor U9031 (N_9031,N_8992,N_8944);
nor U9032 (N_9032,N_8809,N_8891);
nand U9033 (N_9033,N_8942,N_8938);
nor U9034 (N_9034,N_8899,N_8921);
or U9035 (N_9035,N_8961,N_8901);
and U9036 (N_9036,N_8860,N_8985);
nand U9037 (N_9037,N_8972,N_8879);
and U9038 (N_9038,N_8940,N_8936);
and U9039 (N_9039,N_8957,N_8912);
or U9040 (N_9040,N_8817,N_8884);
nand U9041 (N_9041,N_8814,N_8834);
nand U9042 (N_9042,N_8969,N_8897);
nand U9043 (N_9043,N_8974,N_8848);
nand U9044 (N_9044,N_8886,N_8931);
nand U9045 (N_9045,N_8911,N_8933);
nand U9046 (N_9046,N_8820,N_8868);
nor U9047 (N_9047,N_8856,N_8869);
and U9048 (N_9048,N_8918,N_8882);
nor U9049 (N_9049,N_8800,N_8929);
and U9050 (N_9050,N_8836,N_8810);
nand U9051 (N_9051,N_8967,N_8840);
and U9052 (N_9052,N_8907,N_8947);
and U9053 (N_9053,N_8845,N_8871);
nand U9054 (N_9054,N_8956,N_8887);
xor U9055 (N_9055,N_8903,N_8863);
nor U9056 (N_9056,N_8953,N_8804);
nand U9057 (N_9057,N_8986,N_8846);
or U9058 (N_9058,N_8815,N_8943);
or U9059 (N_9059,N_8988,N_8841);
xnor U9060 (N_9060,N_8877,N_8824);
or U9061 (N_9061,N_8955,N_8829);
nand U9062 (N_9062,N_8880,N_8913);
nand U9063 (N_9063,N_8811,N_8904);
and U9064 (N_9064,N_8894,N_8842);
nand U9065 (N_9065,N_8821,N_8995);
nand U9066 (N_9066,N_8870,N_8996);
nor U9067 (N_9067,N_8939,N_8941);
nor U9068 (N_9068,N_8984,N_8847);
or U9069 (N_9069,N_8952,N_8839);
nand U9070 (N_9070,N_8805,N_8902);
nand U9071 (N_9071,N_8959,N_8838);
or U9072 (N_9072,N_8803,N_8950);
or U9073 (N_9073,N_8922,N_8865);
or U9074 (N_9074,N_8965,N_8812);
nor U9075 (N_9075,N_8908,N_8997);
and U9076 (N_9076,N_8949,N_8881);
or U9077 (N_9077,N_8807,N_8919);
and U9078 (N_9078,N_8864,N_8964);
nand U9079 (N_9079,N_8934,N_8963);
nor U9080 (N_9080,N_8898,N_8826);
nor U9081 (N_9081,N_8990,N_8926);
or U9082 (N_9082,N_8873,N_8932);
nor U9083 (N_9083,N_8853,N_8813);
nor U9084 (N_9084,N_8843,N_8994);
and U9085 (N_9085,N_8954,N_8900);
and U9086 (N_9086,N_8895,N_8854);
nor U9087 (N_9087,N_8833,N_8989);
nor U9088 (N_9088,N_8937,N_8896);
and U9089 (N_9089,N_8835,N_8930);
and U9090 (N_9090,N_8910,N_8925);
nand U9091 (N_9091,N_8883,N_8945);
or U9092 (N_9092,N_8875,N_8970);
nand U9093 (N_9093,N_8983,N_8893);
or U9094 (N_9094,N_8909,N_8958);
nor U9095 (N_9095,N_8973,N_8844);
or U9096 (N_9096,N_8823,N_8855);
nand U9097 (N_9097,N_8928,N_8822);
nand U9098 (N_9098,N_8905,N_8851);
nor U9099 (N_9099,N_8801,N_8920);
nand U9100 (N_9100,N_8976,N_8901);
nor U9101 (N_9101,N_8992,N_8919);
nor U9102 (N_9102,N_8905,N_8945);
nor U9103 (N_9103,N_8923,N_8882);
or U9104 (N_9104,N_8802,N_8918);
nand U9105 (N_9105,N_8909,N_8984);
or U9106 (N_9106,N_8905,N_8943);
or U9107 (N_9107,N_8876,N_8988);
nor U9108 (N_9108,N_8810,N_8850);
nand U9109 (N_9109,N_8847,N_8869);
or U9110 (N_9110,N_8847,N_8866);
nor U9111 (N_9111,N_8909,N_8877);
and U9112 (N_9112,N_8951,N_8832);
or U9113 (N_9113,N_8965,N_8970);
nand U9114 (N_9114,N_8828,N_8920);
nand U9115 (N_9115,N_8879,N_8937);
or U9116 (N_9116,N_8949,N_8987);
nand U9117 (N_9117,N_8832,N_8849);
nand U9118 (N_9118,N_8842,N_8973);
or U9119 (N_9119,N_8871,N_8812);
or U9120 (N_9120,N_8951,N_8948);
or U9121 (N_9121,N_8851,N_8993);
nor U9122 (N_9122,N_8975,N_8841);
xnor U9123 (N_9123,N_8960,N_8867);
or U9124 (N_9124,N_8912,N_8868);
and U9125 (N_9125,N_8938,N_8889);
or U9126 (N_9126,N_8941,N_8874);
nand U9127 (N_9127,N_8877,N_8985);
nand U9128 (N_9128,N_8983,N_8884);
nand U9129 (N_9129,N_8927,N_8858);
xor U9130 (N_9130,N_8815,N_8803);
nor U9131 (N_9131,N_8801,N_8872);
nor U9132 (N_9132,N_8960,N_8900);
and U9133 (N_9133,N_8967,N_8897);
nor U9134 (N_9134,N_8981,N_8990);
and U9135 (N_9135,N_8914,N_8835);
xor U9136 (N_9136,N_8883,N_8804);
nand U9137 (N_9137,N_8995,N_8940);
and U9138 (N_9138,N_8991,N_8812);
nor U9139 (N_9139,N_8994,N_8916);
nand U9140 (N_9140,N_8822,N_8882);
nor U9141 (N_9141,N_8870,N_8937);
and U9142 (N_9142,N_8932,N_8867);
and U9143 (N_9143,N_8805,N_8868);
nor U9144 (N_9144,N_8839,N_8947);
nand U9145 (N_9145,N_8877,N_8912);
or U9146 (N_9146,N_8927,N_8802);
and U9147 (N_9147,N_8971,N_8924);
nor U9148 (N_9148,N_8802,N_8848);
nand U9149 (N_9149,N_8886,N_8817);
or U9150 (N_9150,N_8869,N_8813);
or U9151 (N_9151,N_8976,N_8879);
or U9152 (N_9152,N_8978,N_8968);
or U9153 (N_9153,N_8940,N_8913);
or U9154 (N_9154,N_8907,N_8971);
nor U9155 (N_9155,N_8839,N_8879);
nand U9156 (N_9156,N_8869,N_8928);
nand U9157 (N_9157,N_8831,N_8817);
nor U9158 (N_9158,N_8824,N_8848);
or U9159 (N_9159,N_8846,N_8909);
nor U9160 (N_9160,N_8999,N_8809);
or U9161 (N_9161,N_8867,N_8983);
nand U9162 (N_9162,N_8845,N_8870);
nand U9163 (N_9163,N_8930,N_8953);
nor U9164 (N_9164,N_8814,N_8807);
nor U9165 (N_9165,N_8899,N_8843);
and U9166 (N_9166,N_8897,N_8975);
nand U9167 (N_9167,N_8967,N_8983);
nand U9168 (N_9168,N_8983,N_8848);
nor U9169 (N_9169,N_8802,N_8905);
nand U9170 (N_9170,N_8966,N_8815);
or U9171 (N_9171,N_8885,N_8882);
and U9172 (N_9172,N_8908,N_8984);
nor U9173 (N_9173,N_8815,N_8971);
nand U9174 (N_9174,N_8960,N_8956);
and U9175 (N_9175,N_8976,N_8964);
and U9176 (N_9176,N_8978,N_8866);
or U9177 (N_9177,N_8926,N_8883);
or U9178 (N_9178,N_8994,N_8945);
or U9179 (N_9179,N_8885,N_8831);
nor U9180 (N_9180,N_8987,N_8836);
nand U9181 (N_9181,N_8990,N_8865);
nor U9182 (N_9182,N_8886,N_8959);
nor U9183 (N_9183,N_8802,N_8877);
and U9184 (N_9184,N_8971,N_8947);
nor U9185 (N_9185,N_8857,N_8843);
or U9186 (N_9186,N_8867,N_8988);
nand U9187 (N_9187,N_8999,N_8801);
nand U9188 (N_9188,N_8815,N_8890);
nor U9189 (N_9189,N_8982,N_8840);
nor U9190 (N_9190,N_8803,N_8944);
or U9191 (N_9191,N_8944,N_8850);
and U9192 (N_9192,N_8840,N_8812);
nor U9193 (N_9193,N_8924,N_8880);
nand U9194 (N_9194,N_8872,N_8991);
nor U9195 (N_9195,N_8880,N_8989);
nor U9196 (N_9196,N_8902,N_8916);
nand U9197 (N_9197,N_8867,N_8821);
and U9198 (N_9198,N_8845,N_8998);
and U9199 (N_9199,N_8951,N_8973);
and U9200 (N_9200,N_9110,N_9057);
or U9201 (N_9201,N_9124,N_9022);
nand U9202 (N_9202,N_9128,N_9180);
and U9203 (N_9203,N_9147,N_9139);
nor U9204 (N_9204,N_9121,N_9199);
and U9205 (N_9205,N_9053,N_9035);
nand U9206 (N_9206,N_9096,N_9186);
nand U9207 (N_9207,N_9137,N_9101);
and U9208 (N_9208,N_9135,N_9009);
and U9209 (N_9209,N_9193,N_9127);
nand U9210 (N_9210,N_9075,N_9082);
and U9211 (N_9211,N_9158,N_9189);
nor U9212 (N_9212,N_9145,N_9175);
nor U9213 (N_9213,N_9182,N_9046);
and U9214 (N_9214,N_9078,N_9054);
nand U9215 (N_9215,N_9143,N_9157);
nor U9216 (N_9216,N_9045,N_9120);
nand U9217 (N_9217,N_9034,N_9042);
and U9218 (N_9218,N_9171,N_9134);
nor U9219 (N_9219,N_9015,N_9181);
nor U9220 (N_9220,N_9064,N_9055);
or U9221 (N_9221,N_9125,N_9163);
or U9222 (N_9222,N_9049,N_9081);
nand U9223 (N_9223,N_9018,N_9149);
and U9224 (N_9224,N_9178,N_9197);
nand U9225 (N_9225,N_9154,N_9152);
nor U9226 (N_9226,N_9080,N_9177);
and U9227 (N_9227,N_9047,N_9192);
nor U9228 (N_9228,N_9028,N_9040);
or U9229 (N_9229,N_9169,N_9109);
nand U9230 (N_9230,N_9108,N_9138);
and U9231 (N_9231,N_9179,N_9160);
and U9232 (N_9232,N_9170,N_9033);
or U9233 (N_9233,N_9039,N_9031);
and U9234 (N_9234,N_9103,N_9062);
nand U9235 (N_9235,N_9017,N_9194);
nor U9236 (N_9236,N_9013,N_9097);
and U9237 (N_9237,N_9073,N_9164);
nand U9238 (N_9238,N_9100,N_9059);
nor U9239 (N_9239,N_9020,N_9184);
or U9240 (N_9240,N_9113,N_9117);
or U9241 (N_9241,N_9130,N_9112);
and U9242 (N_9242,N_9027,N_9038);
nand U9243 (N_9243,N_9001,N_9026);
nand U9244 (N_9244,N_9068,N_9111);
or U9245 (N_9245,N_9076,N_9014);
nor U9246 (N_9246,N_9056,N_9183);
nand U9247 (N_9247,N_9048,N_9041);
or U9248 (N_9248,N_9063,N_9070);
or U9249 (N_9249,N_9168,N_9187);
and U9250 (N_9250,N_9066,N_9131);
or U9251 (N_9251,N_9190,N_9092);
nor U9252 (N_9252,N_9016,N_9141);
nand U9253 (N_9253,N_9051,N_9052);
or U9254 (N_9254,N_9185,N_9174);
nor U9255 (N_9255,N_9029,N_9165);
nand U9256 (N_9256,N_9044,N_9133);
xor U9257 (N_9257,N_9161,N_9024);
and U9258 (N_9258,N_9071,N_9146);
and U9259 (N_9259,N_9000,N_9104);
or U9260 (N_9260,N_9116,N_9087);
and U9261 (N_9261,N_9072,N_9167);
nor U9262 (N_9262,N_9151,N_9106);
and U9263 (N_9263,N_9093,N_9030);
nand U9264 (N_9264,N_9008,N_9065);
nand U9265 (N_9265,N_9119,N_9150);
nor U9266 (N_9266,N_9090,N_9156);
or U9267 (N_9267,N_9136,N_9155);
nor U9268 (N_9268,N_9188,N_9098);
or U9269 (N_9269,N_9077,N_9037);
nand U9270 (N_9270,N_9105,N_9198);
nor U9271 (N_9271,N_9142,N_9148);
nor U9272 (N_9272,N_9067,N_9032);
or U9273 (N_9273,N_9021,N_9088);
or U9274 (N_9274,N_9083,N_9159);
and U9275 (N_9275,N_9007,N_9019);
or U9276 (N_9276,N_9079,N_9089);
nor U9277 (N_9277,N_9196,N_9061);
nor U9278 (N_9278,N_9166,N_9173);
and U9279 (N_9279,N_9050,N_9102);
or U9280 (N_9280,N_9191,N_9025);
nand U9281 (N_9281,N_9005,N_9132);
or U9282 (N_9282,N_9129,N_9085);
nand U9283 (N_9283,N_9002,N_9195);
nor U9284 (N_9284,N_9086,N_9058);
nor U9285 (N_9285,N_9107,N_9144);
and U9286 (N_9286,N_9114,N_9094);
and U9287 (N_9287,N_9023,N_9010);
and U9288 (N_9288,N_9140,N_9074);
xnor U9289 (N_9289,N_9172,N_9162);
and U9290 (N_9290,N_9012,N_9004);
nor U9291 (N_9291,N_9091,N_9153);
nor U9292 (N_9292,N_9003,N_9122);
and U9293 (N_9293,N_9036,N_9115);
or U9294 (N_9294,N_9118,N_9126);
or U9295 (N_9295,N_9060,N_9095);
nor U9296 (N_9296,N_9099,N_9123);
nor U9297 (N_9297,N_9176,N_9011);
or U9298 (N_9298,N_9006,N_9084);
and U9299 (N_9299,N_9043,N_9069);
and U9300 (N_9300,N_9086,N_9031);
nand U9301 (N_9301,N_9041,N_9104);
nand U9302 (N_9302,N_9175,N_9026);
and U9303 (N_9303,N_9191,N_9033);
nand U9304 (N_9304,N_9141,N_9019);
nor U9305 (N_9305,N_9193,N_9072);
or U9306 (N_9306,N_9030,N_9197);
and U9307 (N_9307,N_9033,N_9019);
nor U9308 (N_9308,N_9154,N_9192);
nand U9309 (N_9309,N_9083,N_9133);
nand U9310 (N_9310,N_9038,N_9151);
or U9311 (N_9311,N_9056,N_9132);
nand U9312 (N_9312,N_9175,N_9004);
or U9313 (N_9313,N_9127,N_9160);
nand U9314 (N_9314,N_9022,N_9080);
or U9315 (N_9315,N_9135,N_9131);
and U9316 (N_9316,N_9131,N_9138);
or U9317 (N_9317,N_9026,N_9012);
and U9318 (N_9318,N_9155,N_9070);
or U9319 (N_9319,N_9042,N_9082);
and U9320 (N_9320,N_9135,N_9060);
and U9321 (N_9321,N_9125,N_9085);
nand U9322 (N_9322,N_9027,N_9167);
or U9323 (N_9323,N_9096,N_9030);
or U9324 (N_9324,N_9020,N_9132);
or U9325 (N_9325,N_9015,N_9103);
nand U9326 (N_9326,N_9114,N_9172);
or U9327 (N_9327,N_9130,N_9104);
nor U9328 (N_9328,N_9156,N_9176);
nor U9329 (N_9329,N_9153,N_9109);
nor U9330 (N_9330,N_9188,N_9025);
nor U9331 (N_9331,N_9039,N_9119);
and U9332 (N_9332,N_9032,N_9197);
nand U9333 (N_9333,N_9187,N_9027);
nor U9334 (N_9334,N_9068,N_9137);
and U9335 (N_9335,N_9052,N_9081);
and U9336 (N_9336,N_9078,N_9125);
xnor U9337 (N_9337,N_9066,N_9068);
xor U9338 (N_9338,N_9176,N_9071);
nor U9339 (N_9339,N_9047,N_9012);
and U9340 (N_9340,N_9175,N_9131);
or U9341 (N_9341,N_9033,N_9140);
and U9342 (N_9342,N_9167,N_9061);
or U9343 (N_9343,N_9067,N_9147);
nor U9344 (N_9344,N_9139,N_9184);
or U9345 (N_9345,N_9066,N_9082);
nor U9346 (N_9346,N_9106,N_9192);
and U9347 (N_9347,N_9005,N_9186);
nor U9348 (N_9348,N_9112,N_9094);
xor U9349 (N_9349,N_9169,N_9067);
nor U9350 (N_9350,N_9000,N_9134);
nor U9351 (N_9351,N_9019,N_9079);
nand U9352 (N_9352,N_9194,N_9138);
and U9353 (N_9353,N_9008,N_9060);
nor U9354 (N_9354,N_9129,N_9015);
nand U9355 (N_9355,N_9088,N_9118);
and U9356 (N_9356,N_9070,N_9041);
nand U9357 (N_9357,N_9056,N_9146);
or U9358 (N_9358,N_9012,N_9143);
or U9359 (N_9359,N_9172,N_9119);
nor U9360 (N_9360,N_9052,N_9131);
and U9361 (N_9361,N_9160,N_9090);
and U9362 (N_9362,N_9048,N_9089);
nand U9363 (N_9363,N_9066,N_9199);
or U9364 (N_9364,N_9099,N_9108);
nand U9365 (N_9365,N_9175,N_9105);
nand U9366 (N_9366,N_9186,N_9164);
nand U9367 (N_9367,N_9078,N_9066);
or U9368 (N_9368,N_9129,N_9051);
nor U9369 (N_9369,N_9179,N_9129);
nor U9370 (N_9370,N_9159,N_9161);
or U9371 (N_9371,N_9188,N_9195);
nor U9372 (N_9372,N_9025,N_9119);
nand U9373 (N_9373,N_9086,N_9155);
or U9374 (N_9374,N_9161,N_9074);
and U9375 (N_9375,N_9116,N_9018);
and U9376 (N_9376,N_9050,N_9033);
or U9377 (N_9377,N_9041,N_9164);
and U9378 (N_9378,N_9134,N_9180);
and U9379 (N_9379,N_9199,N_9072);
nand U9380 (N_9380,N_9181,N_9138);
and U9381 (N_9381,N_9041,N_9014);
or U9382 (N_9382,N_9120,N_9195);
nor U9383 (N_9383,N_9148,N_9141);
nor U9384 (N_9384,N_9177,N_9006);
nand U9385 (N_9385,N_9011,N_9033);
nand U9386 (N_9386,N_9149,N_9093);
or U9387 (N_9387,N_9196,N_9020);
nor U9388 (N_9388,N_9066,N_9137);
nor U9389 (N_9389,N_9017,N_9047);
or U9390 (N_9390,N_9023,N_9053);
nor U9391 (N_9391,N_9136,N_9184);
or U9392 (N_9392,N_9070,N_9077);
nor U9393 (N_9393,N_9152,N_9094);
nor U9394 (N_9394,N_9141,N_9084);
and U9395 (N_9395,N_9071,N_9177);
nand U9396 (N_9396,N_9154,N_9036);
or U9397 (N_9397,N_9004,N_9015);
nand U9398 (N_9398,N_9113,N_9180);
nor U9399 (N_9399,N_9060,N_9005);
nand U9400 (N_9400,N_9375,N_9233);
xnor U9401 (N_9401,N_9344,N_9225);
and U9402 (N_9402,N_9252,N_9213);
and U9403 (N_9403,N_9307,N_9351);
or U9404 (N_9404,N_9378,N_9244);
or U9405 (N_9405,N_9303,N_9325);
nor U9406 (N_9406,N_9216,N_9289);
and U9407 (N_9407,N_9269,N_9238);
or U9408 (N_9408,N_9354,N_9258);
nand U9409 (N_9409,N_9396,N_9353);
nand U9410 (N_9410,N_9217,N_9251);
xor U9411 (N_9411,N_9320,N_9223);
or U9412 (N_9412,N_9279,N_9308);
nor U9413 (N_9413,N_9345,N_9265);
and U9414 (N_9414,N_9367,N_9256);
nand U9415 (N_9415,N_9209,N_9397);
nand U9416 (N_9416,N_9337,N_9359);
or U9417 (N_9417,N_9394,N_9310);
nand U9418 (N_9418,N_9296,N_9263);
nor U9419 (N_9419,N_9366,N_9348);
nand U9420 (N_9420,N_9387,N_9379);
and U9421 (N_9421,N_9262,N_9364);
and U9422 (N_9422,N_9336,N_9319);
nand U9423 (N_9423,N_9365,N_9290);
and U9424 (N_9424,N_9340,N_9241);
nor U9425 (N_9425,N_9287,N_9376);
and U9426 (N_9426,N_9204,N_9304);
or U9427 (N_9427,N_9382,N_9285);
nor U9428 (N_9428,N_9395,N_9257);
nor U9429 (N_9429,N_9212,N_9264);
or U9430 (N_9430,N_9361,N_9322);
and U9431 (N_9431,N_9329,N_9250);
or U9432 (N_9432,N_9346,N_9356);
nor U9433 (N_9433,N_9371,N_9274);
and U9434 (N_9434,N_9318,N_9277);
nor U9435 (N_9435,N_9231,N_9243);
nor U9436 (N_9436,N_9278,N_9254);
nor U9437 (N_9437,N_9239,N_9305);
nand U9438 (N_9438,N_9328,N_9342);
and U9439 (N_9439,N_9343,N_9358);
nor U9440 (N_9440,N_9333,N_9245);
nor U9441 (N_9441,N_9202,N_9339);
and U9442 (N_9442,N_9219,N_9324);
nor U9443 (N_9443,N_9293,N_9386);
nor U9444 (N_9444,N_9334,N_9282);
and U9445 (N_9445,N_9388,N_9363);
and U9446 (N_9446,N_9276,N_9220);
nor U9447 (N_9447,N_9393,N_9315);
nand U9448 (N_9448,N_9321,N_9255);
and U9449 (N_9449,N_9377,N_9399);
or U9450 (N_9450,N_9327,N_9338);
xnor U9451 (N_9451,N_9208,N_9384);
or U9452 (N_9452,N_9229,N_9272);
nor U9453 (N_9453,N_9326,N_9349);
or U9454 (N_9454,N_9299,N_9341);
or U9455 (N_9455,N_9283,N_9281);
nor U9456 (N_9456,N_9226,N_9301);
and U9457 (N_9457,N_9373,N_9398);
nor U9458 (N_9458,N_9357,N_9235);
and U9459 (N_9459,N_9267,N_9275);
nand U9460 (N_9460,N_9370,N_9331);
and U9461 (N_9461,N_9311,N_9215);
or U9462 (N_9462,N_9224,N_9237);
or U9463 (N_9463,N_9368,N_9313);
or U9464 (N_9464,N_9205,N_9242);
nand U9465 (N_9465,N_9309,N_9240);
or U9466 (N_9466,N_9230,N_9317);
or U9467 (N_9467,N_9291,N_9374);
nand U9468 (N_9468,N_9228,N_9350);
and U9469 (N_9469,N_9391,N_9210);
xor U9470 (N_9470,N_9369,N_9335);
or U9471 (N_9471,N_9298,N_9284);
nand U9472 (N_9472,N_9261,N_9389);
or U9473 (N_9473,N_9280,N_9271);
nor U9474 (N_9474,N_9314,N_9372);
or U9475 (N_9475,N_9246,N_9297);
or U9476 (N_9476,N_9306,N_9392);
and U9477 (N_9477,N_9248,N_9312);
nand U9478 (N_9478,N_9286,N_9270);
nor U9479 (N_9479,N_9380,N_9222);
or U9480 (N_9480,N_9249,N_9294);
and U9481 (N_9481,N_9316,N_9352);
and U9482 (N_9482,N_9214,N_9232);
nor U9483 (N_9483,N_9300,N_9236);
nor U9484 (N_9484,N_9206,N_9292);
nand U9485 (N_9485,N_9360,N_9207);
nor U9486 (N_9486,N_9323,N_9260);
nand U9487 (N_9487,N_9227,N_9203);
nor U9488 (N_9488,N_9385,N_9218);
or U9489 (N_9489,N_9247,N_9211);
nor U9490 (N_9490,N_9259,N_9268);
and U9491 (N_9491,N_9383,N_9381);
nand U9492 (N_9492,N_9273,N_9330);
nor U9493 (N_9493,N_9200,N_9302);
nand U9494 (N_9494,N_9390,N_9295);
and U9495 (N_9495,N_9253,N_9266);
nor U9496 (N_9496,N_9201,N_9288);
nand U9497 (N_9497,N_9362,N_9355);
nor U9498 (N_9498,N_9221,N_9234);
or U9499 (N_9499,N_9347,N_9332);
nor U9500 (N_9500,N_9246,N_9285);
or U9501 (N_9501,N_9286,N_9294);
xnor U9502 (N_9502,N_9320,N_9244);
nand U9503 (N_9503,N_9345,N_9321);
and U9504 (N_9504,N_9389,N_9275);
nand U9505 (N_9505,N_9200,N_9366);
nand U9506 (N_9506,N_9269,N_9230);
or U9507 (N_9507,N_9235,N_9248);
or U9508 (N_9508,N_9332,N_9380);
nand U9509 (N_9509,N_9356,N_9256);
and U9510 (N_9510,N_9254,N_9305);
nor U9511 (N_9511,N_9266,N_9303);
nor U9512 (N_9512,N_9347,N_9311);
and U9513 (N_9513,N_9338,N_9265);
or U9514 (N_9514,N_9322,N_9209);
and U9515 (N_9515,N_9260,N_9353);
or U9516 (N_9516,N_9381,N_9236);
or U9517 (N_9517,N_9330,N_9388);
and U9518 (N_9518,N_9341,N_9212);
or U9519 (N_9519,N_9306,N_9334);
and U9520 (N_9520,N_9262,N_9392);
nand U9521 (N_9521,N_9338,N_9328);
or U9522 (N_9522,N_9349,N_9297);
nor U9523 (N_9523,N_9368,N_9320);
xor U9524 (N_9524,N_9211,N_9339);
nand U9525 (N_9525,N_9346,N_9377);
and U9526 (N_9526,N_9317,N_9371);
nor U9527 (N_9527,N_9321,N_9359);
nor U9528 (N_9528,N_9281,N_9372);
nand U9529 (N_9529,N_9383,N_9272);
xnor U9530 (N_9530,N_9346,N_9360);
and U9531 (N_9531,N_9228,N_9324);
nor U9532 (N_9532,N_9361,N_9235);
nand U9533 (N_9533,N_9326,N_9264);
nand U9534 (N_9534,N_9265,N_9282);
nand U9535 (N_9535,N_9310,N_9368);
nor U9536 (N_9536,N_9226,N_9380);
and U9537 (N_9537,N_9290,N_9237);
nor U9538 (N_9538,N_9214,N_9395);
nand U9539 (N_9539,N_9313,N_9317);
nand U9540 (N_9540,N_9374,N_9307);
and U9541 (N_9541,N_9267,N_9385);
nand U9542 (N_9542,N_9345,N_9278);
nand U9543 (N_9543,N_9393,N_9273);
or U9544 (N_9544,N_9313,N_9238);
nand U9545 (N_9545,N_9316,N_9379);
nand U9546 (N_9546,N_9380,N_9342);
nor U9547 (N_9547,N_9233,N_9308);
and U9548 (N_9548,N_9300,N_9269);
and U9549 (N_9549,N_9214,N_9258);
nand U9550 (N_9550,N_9218,N_9258);
nor U9551 (N_9551,N_9370,N_9204);
nand U9552 (N_9552,N_9395,N_9265);
nand U9553 (N_9553,N_9236,N_9259);
and U9554 (N_9554,N_9370,N_9276);
xor U9555 (N_9555,N_9228,N_9360);
nor U9556 (N_9556,N_9362,N_9319);
nor U9557 (N_9557,N_9295,N_9214);
or U9558 (N_9558,N_9255,N_9212);
nor U9559 (N_9559,N_9305,N_9261);
nand U9560 (N_9560,N_9276,N_9231);
and U9561 (N_9561,N_9223,N_9339);
or U9562 (N_9562,N_9238,N_9363);
and U9563 (N_9563,N_9243,N_9384);
or U9564 (N_9564,N_9238,N_9343);
or U9565 (N_9565,N_9266,N_9260);
nand U9566 (N_9566,N_9368,N_9216);
nor U9567 (N_9567,N_9349,N_9315);
and U9568 (N_9568,N_9210,N_9298);
nor U9569 (N_9569,N_9330,N_9274);
nand U9570 (N_9570,N_9388,N_9373);
nor U9571 (N_9571,N_9336,N_9257);
or U9572 (N_9572,N_9367,N_9333);
nand U9573 (N_9573,N_9384,N_9399);
and U9574 (N_9574,N_9263,N_9345);
nand U9575 (N_9575,N_9286,N_9228);
nand U9576 (N_9576,N_9357,N_9286);
nor U9577 (N_9577,N_9281,N_9319);
nor U9578 (N_9578,N_9381,N_9362);
nand U9579 (N_9579,N_9390,N_9320);
and U9580 (N_9580,N_9379,N_9344);
nand U9581 (N_9581,N_9219,N_9238);
or U9582 (N_9582,N_9300,N_9336);
or U9583 (N_9583,N_9369,N_9285);
and U9584 (N_9584,N_9240,N_9317);
nand U9585 (N_9585,N_9389,N_9270);
or U9586 (N_9586,N_9319,N_9213);
nand U9587 (N_9587,N_9249,N_9266);
nand U9588 (N_9588,N_9217,N_9328);
or U9589 (N_9589,N_9226,N_9377);
and U9590 (N_9590,N_9238,N_9280);
nor U9591 (N_9591,N_9224,N_9234);
nor U9592 (N_9592,N_9289,N_9312);
or U9593 (N_9593,N_9277,N_9348);
or U9594 (N_9594,N_9378,N_9334);
or U9595 (N_9595,N_9345,N_9214);
nor U9596 (N_9596,N_9391,N_9276);
xnor U9597 (N_9597,N_9244,N_9344);
or U9598 (N_9598,N_9365,N_9325);
nor U9599 (N_9599,N_9268,N_9249);
or U9600 (N_9600,N_9554,N_9481);
nand U9601 (N_9601,N_9449,N_9452);
xnor U9602 (N_9602,N_9473,N_9535);
nor U9603 (N_9603,N_9450,N_9444);
or U9604 (N_9604,N_9494,N_9570);
and U9605 (N_9605,N_9490,N_9423);
nor U9606 (N_9606,N_9409,N_9577);
nor U9607 (N_9607,N_9595,N_9443);
nor U9608 (N_9608,N_9491,N_9511);
nor U9609 (N_9609,N_9573,N_9442);
and U9610 (N_9610,N_9582,N_9402);
or U9611 (N_9611,N_9411,N_9406);
nor U9612 (N_9612,N_9550,N_9558);
and U9613 (N_9613,N_9469,N_9598);
nor U9614 (N_9614,N_9540,N_9427);
or U9615 (N_9615,N_9506,N_9581);
nand U9616 (N_9616,N_9401,N_9532);
nand U9617 (N_9617,N_9584,N_9571);
or U9618 (N_9618,N_9586,N_9526);
nand U9619 (N_9619,N_9456,N_9588);
nor U9620 (N_9620,N_9447,N_9487);
and U9621 (N_9621,N_9422,N_9563);
and U9622 (N_9622,N_9551,N_9478);
nand U9623 (N_9623,N_9508,N_9549);
nand U9624 (N_9624,N_9597,N_9421);
nand U9625 (N_9625,N_9589,N_9400);
and U9626 (N_9626,N_9465,N_9455);
and U9627 (N_9627,N_9419,N_9504);
nor U9628 (N_9628,N_9579,N_9403);
nand U9629 (N_9629,N_9561,N_9440);
and U9630 (N_9630,N_9566,N_9559);
nor U9631 (N_9631,N_9430,N_9509);
and U9632 (N_9632,N_9435,N_9591);
and U9633 (N_9633,N_9521,N_9461);
nand U9634 (N_9634,N_9546,N_9416);
or U9635 (N_9635,N_9545,N_9585);
and U9636 (N_9636,N_9553,N_9433);
and U9637 (N_9637,N_9594,N_9468);
nor U9638 (N_9638,N_9458,N_9434);
nor U9639 (N_9639,N_9441,N_9425);
nor U9640 (N_9640,N_9474,N_9544);
nand U9641 (N_9641,N_9569,N_9459);
and U9642 (N_9642,N_9480,N_9492);
nand U9643 (N_9643,N_9483,N_9596);
xor U9644 (N_9644,N_9412,N_9572);
nor U9645 (N_9645,N_9445,N_9576);
and U9646 (N_9646,N_9524,N_9417);
nand U9647 (N_9647,N_9470,N_9583);
and U9648 (N_9648,N_9493,N_9439);
nor U9649 (N_9649,N_9479,N_9472);
and U9650 (N_9650,N_9533,N_9556);
or U9651 (N_9651,N_9488,N_9527);
nand U9652 (N_9652,N_9414,N_9438);
nor U9653 (N_9653,N_9529,N_9518);
or U9654 (N_9654,N_9503,N_9574);
nor U9655 (N_9655,N_9463,N_9537);
nor U9656 (N_9656,N_9505,N_9536);
nor U9657 (N_9657,N_9530,N_9500);
nand U9658 (N_9658,N_9405,N_9547);
nor U9659 (N_9659,N_9486,N_9523);
and U9660 (N_9660,N_9471,N_9462);
nor U9661 (N_9661,N_9415,N_9484);
nor U9662 (N_9662,N_9512,N_9567);
nor U9663 (N_9663,N_9542,N_9539);
and U9664 (N_9664,N_9498,N_9457);
nor U9665 (N_9665,N_9429,N_9510);
nor U9666 (N_9666,N_9410,N_9513);
nor U9667 (N_9667,N_9564,N_9575);
and U9668 (N_9668,N_9436,N_9460);
or U9669 (N_9669,N_9568,N_9424);
nand U9670 (N_9670,N_9590,N_9507);
or U9671 (N_9671,N_9404,N_9514);
nand U9672 (N_9672,N_9534,N_9496);
nor U9673 (N_9673,N_9413,N_9431);
and U9674 (N_9674,N_9420,N_9489);
and U9675 (N_9675,N_9451,N_9516);
xor U9676 (N_9676,N_9464,N_9466);
and U9677 (N_9677,N_9557,N_9448);
nand U9678 (N_9678,N_9552,N_9495);
or U9679 (N_9679,N_9499,N_9446);
nor U9680 (N_9680,N_9476,N_9485);
and U9681 (N_9681,N_9528,N_9593);
nor U9682 (N_9682,N_9531,N_9497);
and U9683 (N_9683,N_9437,N_9565);
nand U9684 (N_9684,N_9587,N_9408);
nand U9685 (N_9685,N_9519,N_9482);
or U9686 (N_9686,N_9538,N_9517);
nor U9687 (N_9687,N_9467,N_9592);
and U9688 (N_9688,N_9520,N_9555);
nor U9689 (N_9689,N_9426,N_9502);
nor U9690 (N_9690,N_9522,N_9407);
nor U9691 (N_9691,N_9477,N_9543);
or U9692 (N_9692,N_9541,N_9428);
nor U9693 (N_9693,N_9418,N_9599);
nor U9694 (N_9694,N_9562,N_9548);
and U9695 (N_9695,N_9501,N_9475);
and U9696 (N_9696,N_9453,N_9432);
or U9697 (N_9697,N_9578,N_9580);
or U9698 (N_9698,N_9454,N_9560);
nand U9699 (N_9699,N_9515,N_9525);
nor U9700 (N_9700,N_9440,N_9469);
nand U9701 (N_9701,N_9484,N_9551);
nand U9702 (N_9702,N_9476,N_9537);
or U9703 (N_9703,N_9570,N_9577);
nand U9704 (N_9704,N_9589,N_9596);
and U9705 (N_9705,N_9413,N_9574);
or U9706 (N_9706,N_9441,N_9537);
and U9707 (N_9707,N_9510,N_9512);
xnor U9708 (N_9708,N_9581,N_9418);
or U9709 (N_9709,N_9453,N_9535);
nand U9710 (N_9710,N_9426,N_9410);
and U9711 (N_9711,N_9416,N_9475);
or U9712 (N_9712,N_9572,N_9573);
and U9713 (N_9713,N_9458,N_9482);
nand U9714 (N_9714,N_9563,N_9417);
or U9715 (N_9715,N_9429,N_9465);
nand U9716 (N_9716,N_9581,N_9484);
and U9717 (N_9717,N_9461,N_9599);
nand U9718 (N_9718,N_9528,N_9437);
and U9719 (N_9719,N_9472,N_9580);
or U9720 (N_9720,N_9447,N_9421);
nor U9721 (N_9721,N_9445,N_9450);
or U9722 (N_9722,N_9414,N_9431);
nor U9723 (N_9723,N_9526,N_9567);
nor U9724 (N_9724,N_9443,N_9478);
or U9725 (N_9725,N_9489,N_9504);
and U9726 (N_9726,N_9432,N_9480);
or U9727 (N_9727,N_9436,N_9475);
nand U9728 (N_9728,N_9507,N_9472);
and U9729 (N_9729,N_9516,N_9483);
or U9730 (N_9730,N_9413,N_9598);
nand U9731 (N_9731,N_9431,N_9577);
nand U9732 (N_9732,N_9445,N_9427);
xor U9733 (N_9733,N_9598,N_9593);
nor U9734 (N_9734,N_9424,N_9548);
or U9735 (N_9735,N_9503,N_9562);
nor U9736 (N_9736,N_9493,N_9424);
nor U9737 (N_9737,N_9571,N_9455);
and U9738 (N_9738,N_9526,N_9544);
nand U9739 (N_9739,N_9466,N_9412);
nand U9740 (N_9740,N_9418,N_9419);
or U9741 (N_9741,N_9470,N_9522);
or U9742 (N_9742,N_9491,N_9559);
or U9743 (N_9743,N_9502,N_9493);
nor U9744 (N_9744,N_9568,N_9471);
nand U9745 (N_9745,N_9478,N_9460);
or U9746 (N_9746,N_9551,N_9431);
nor U9747 (N_9747,N_9410,N_9555);
and U9748 (N_9748,N_9568,N_9518);
and U9749 (N_9749,N_9436,N_9430);
nand U9750 (N_9750,N_9403,N_9440);
nand U9751 (N_9751,N_9438,N_9424);
nor U9752 (N_9752,N_9420,N_9586);
nor U9753 (N_9753,N_9573,N_9411);
nor U9754 (N_9754,N_9486,N_9409);
and U9755 (N_9755,N_9584,N_9503);
or U9756 (N_9756,N_9590,N_9426);
nand U9757 (N_9757,N_9509,N_9455);
nand U9758 (N_9758,N_9480,N_9420);
nand U9759 (N_9759,N_9568,N_9419);
nand U9760 (N_9760,N_9590,N_9438);
and U9761 (N_9761,N_9549,N_9484);
xnor U9762 (N_9762,N_9511,N_9540);
nor U9763 (N_9763,N_9480,N_9486);
or U9764 (N_9764,N_9530,N_9529);
nor U9765 (N_9765,N_9592,N_9565);
nor U9766 (N_9766,N_9501,N_9530);
nand U9767 (N_9767,N_9471,N_9411);
nor U9768 (N_9768,N_9414,N_9547);
nor U9769 (N_9769,N_9584,N_9510);
or U9770 (N_9770,N_9427,N_9468);
nand U9771 (N_9771,N_9559,N_9450);
or U9772 (N_9772,N_9560,N_9577);
and U9773 (N_9773,N_9403,N_9415);
nor U9774 (N_9774,N_9582,N_9509);
xor U9775 (N_9775,N_9447,N_9488);
xnor U9776 (N_9776,N_9447,N_9449);
or U9777 (N_9777,N_9429,N_9574);
or U9778 (N_9778,N_9569,N_9447);
and U9779 (N_9779,N_9492,N_9470);
or U9780 (N_9780,N_9463,N_9515);
nand U9781 (N_9781,N_9490,N_9584);
nand U9782 (N_9782,N_9489,N_9438);
xnor U9783 (N_9783,N_9407,N_9540);
or U9784 (N_9784,N_9587,N_9438);
and U9785 (N_9785,N_9401,N_9521);
and U9786 (N_9786,N_9597,N_9472);
nor U9787 (N_9787,N_9434,N_9531);
nor U9788 (N_9788,N_9419,N_9593);
nand U9789 (N_9789,N_9543,N_9485);
or U9790 (N_9790,N_9478,N_9585);
and U9791 (N_9791,N_9497,N_9506);
nand U9792 (N_9792,N_9484,N_9469);
nand U9793 (N_9793,N_9511,N_9487);
and U9794 (N_9794,N_9572,N_9456);
nor U9795 (N_9795,N_9550,N_9426);
nor U9796 (N_9796,N_9580,N_9551);
nor U9797 (N_9797,N_9505,N_9485);
nor U9798 (N_9798,N_9530,N_9553);
nand U9799 (N_9799,N_9435,N_9411);
nand U9800 (N_9800,N_9643,N_9600);
nand U9801 (N_9801,N_9691,N_9785);
nor U9802 (N_9802,N_9707,N_9670);
or U9803 (N_9803,N_9769,N_9748);
nand U9804 (N_9804,N_9612,N_9662);
nand U9805 (N_9805,N_9796,N_9782);
and U9806 (N_9806,N_9633,N_9686);
xor U9807 (N_9807,N_9618,N_9710);
and U9808 (N_9808,N_9665,N_9716);
or U9809 (N_9809,N_9698,N_9774);
nand U9810 (N_9810,N_9619,N_9630);
nand U9811 (N_9811,N_9765,N_9627);
nand U9812 (N_9812,N_9683,N_9671);
nor U9813 (N_9813,N_9731,N_9734);
nand U9814 (N_9814,N_9628,N_9615);
and U9815 (N_9815,N_9764,N_9678);
and U9816 (N_9816,N_9742,N_9778);
and U9817 (N_9817,N_9791,N_9732);
and U9818 (N_9818,N_9660,N_9684);
or U9819 (N_9819,N_9621,N_9755);
nor U9820 (N_9820,N_9724,N_9733);
or U9821 (N_9821,N_9607,N_9620);
or U9822 (N_9822,N_9746,N_9702);
or U9823 (N_9823,N_9721,N_9792);
xor U9824 (N_9824,N_9690,N_9728);
and U9825 (N_9825,N_9653,N_9753);
nor U9826 (N_9826,N_9750,N_9737);
nor U9827 (N_9827,N_9705,N_9756);
and U9828 (N_9828,N_9757,N_9719);
and U9829 (N_9829,N_9712,N_9609);
and U9830 (N_9830,N_9648,N_9752);
and U9831 (N_9831,N_9727,N_9775);
nor U9832 (N_9832,N_9606,N_9651);
nand U9833 (N_9833,N_9739,N_9623);
or U9834 (N_9834,N_9789,N_9700);
nand U9835 (N_9835,N_9685,N_9767);
and U9836 (N_9836,N_9706,N_9629);
nor U9837 (N_9837,N_9770,N_9637);
or U9838 (N_9838,N_9672,N_9656);
nor U9839 (N_9839,N_9632,N_9749);
and U9840 (N_9840,N_9772,N_9661);
and U9841 (N_9841,N_9795,N_9645);
nor U9842 (N_9842,N_9622,N_9675);
nand U9843 (N_9843,N_9608,N_9655);
or U9844 (N_9844,N_9713,N_9725);
and U9845 (N_9845,N_9701,N_9649);
or U9846 (N_9846,N_9704,N_9694);
and U9847 (N_9847,N_9718,N_9642);
and U9848 (N_9848,N_9664,N_9693);
and U9849 (N_9849,N_9740,N_9761);
nor U9850 (N_9850,N_9614,N_9797);
or U9851 (N_9851,N_9681,N_9639);
and U9852 (N_9852,N_9673,N_9603);
and U9853 (N_9853,N_9784,N_9604);
nor U9854 (N_9854,N_9626,N_9758);
or U9855 (N_9855,N_9692,N_9687);
or U9856 (N_9856,N_9650,N_9735);
and U9857 (N_9857,N_9715,N_9605);
nand U9858 (N_9858,N_9745,N_9647);
nand U9859 (N_9859,N_9790,N_9788);
and U9860 (N_9860,N_9635,N_9658);
nor U9861 (N_9861,N_9625,N_9760);
and U9862 (N_9862,N_9668,N_9730);
and U9863 (N_9863,N_9747,N_9709);
and U9864 (N_9864,N_9624,N_9674);
and U9865 (N_9865,N_9697,N_9667);
nor U9866 (N_9866,N_9741,N_9652);
and U9867 (N_9867,N_9663,N_9714);
nand U9868 (N_9868,N_9766,N_9617);
nor U9869 (N_9869,N_9708,N_9679);
nor U9870 (N_9870,N_9657,N_9763);
or U9871 (N_9871,N_9654,N_9754);
nand U9872 (N_9872,N_9680,N_9689);
and U9873 (N_9873,N_9794,N_9777);
and U9874 (N_9874,N_9786,N_9773);
nor U9875 (N_9875,N_9771,N_9726);
and U9876 (N_9876,N_9616,N_9676);
and U9877 (N_9877,N_9738,N_9783);
or U9878 (N_9878,N_9717,N_9677);
and U9879 (N_9879,N_9781,N_9610);
nor U9880 (N_9880,N_9779,N_9682);
nor U9881 (N_9881,N_9762,N_9723);
nand U9882 (N_9882,N_9759,N_9720);
nor U9883 (N_9883,N_9711,N_9669);
nand U9884 (N_9884,N_9722,N_9751);
xnor U9885 (N_9885,N_9768,N_9613);
and U9886 (N_9886,N_9798,N_9729);
or U9887 (N_9887,N_9601,N_9703);
nor U9888 (N_9888,N_9799,N_9688);
and U9889 (N_9889,N_9666,N_9696);
or U9890 (N_9890,N_9787,N_9634);
nor U9891 (N_9891,N_9736,N_9659);
nor U9892 (N_9892,N_9744,N_9793);
or U9893 (N_9893,N_9743,N_9641);
or U9894 (N_9894,N_9640,N_9780);
nor U9895 (N_9895,N_9611,N_9638);
and U9896 (N_9896,N_9776,N_9644);
nand U9897 (N_9897,N_9631,N_9695);
nand U9898 (N_9898,N_9636,N_9699);
nor U9899 (N_9899,N_9602,N_9646);
or U9900 (N_9900,N_9785,N_9614);
nor U9901 (N_9901,N_9641,N_9765);
nand U9902 (N_9902,N_9709,N_9794);
nor U9903 (N_9903,N_9637,N_9641);
and U9904 (N_9904,N_9775,N_9705);
nand U9905 (N_9905,N_9678,N_9728);
or U9906 (N_9906,N_9735,N_9739);
or U9907 (N_9907,N_9731,N_9714);
and U9908 (N_9908,N_9786,N_9714);
and U9909 (N_9909,N_9775,N_9696);
nand U9910 (N_9910,N_9785,N_9667);
nand U9911 (N_9911,N_9615,N_9665);
or U9912 (N_9912,N_9625,N_9706);
and U9913 (N_9913,N_9624,N_9625);
or U9914 (N_9914,N_9748,N_9630);
or U9915 (N_9915,N_9782,N_9734);
and U9916 (N_9916,N_9650,N_9729);
and U9917 (N_9917,N_9641,N_9601);
nand U9918 (N_9918,N_9709,N_9722);
and U9919 (N_9919,N_9662,N_9731);
nor U9920 (N_9920,N_9601,N_9704);
and U9921 (N_9921,N_9715,N_9726);
nand U9922 (N_9922,N_9772,N_9755);
or U9923 (N_9923,N_9790,N_9623);
nand U9924 (N_9924,N_9605,N_9752);
nor U9925 (N_9925,N_9642,N_9793);
or U9926 (N_9926,N_9691,N_9779);
and U9927 (N_9927,N_9674,N_9752);
and U9928 (N_9928,N_9742,N_9766);
and U9929 (N_9929,N_9762,N_9615);
and U9930 (N_9930,N_9773,N_9737);
and U9931 (N_9931,N_9668,N_9723);
and U9932 (N_9932,N_9642,N_9603);
nand U9933 (N_9933,N_9672,N_9677);
or U9934 (N_9934,N_9764,N_9613);
and U9935 (N_9935,N_9781,N_9663);
nor U9936 (N_9936,N_9772,N_9757);
and U9937 (N_9937,N_9787,N_9676);
nand U9938 (N_9938,N_9722,N_9628);
and U9939 (N_9939,N_9678,N_9775);
or U9940 (N_9940,N_9729,N_9747);
nor U9941 (N_9941,N_9755,N_9752);
nand U9942 (N_9942,N_9662,N_9720);
and U9943 (N_9943,N_9675,N_9696);
and U9944 (N_9944,N_9622,N_9773);
or U9945 (N_9945,N_9600,N_9622);
or U9946 (N_9946,N_9785,N_9670);
and U9947 (N_9947,N_9606,N_9646);
nor U9948 (N_9948,N_9612,N_9624);
and U9949 (N_9949,N_9666,N_9704);
nand U9950 (N_9950,N_9681,N_9698);
and U9951 (N_9951,N_9737,N_9649);
or U9952 (N_9952,N_9634,N_9638);
or U9953 (N_9953,N_9618,N_9783);
xor U9954 (N_9954,N_9653,N_9751);
nand U9955 (N_9955,N_9720,N_9644);
and U9956 (N_9956,N_9786,N_9797);
or U9957 (N_9957,N_9724,N_9739);
nor U9958 (N_9958,N_9752,N_9600);
xnor U9959 (N_9959,N_9657,N_9661);
nand U9960 (N_9960,N_9642,N_9659);
and U9961 (N_9961,N_9668,N_9680);
and U9962 (N_9962,N_9751,N_9624);
or U9963 (N_9963,N_9774,N_9718);
xor U9964 (N_9964,N_9732,N_9735);
and U9965 (N_9965,N_9691,N_9754);
and U9966 (N_9966,N_9760,N_9671);
nand U9967 (N_9967,N_9766,N_9759);
and U9968 (N_9968,N_9752,N_9693);
or U9969 (N_9969,N_9657,N_9796);
nand U9970 (N_9970,N_9677,N_9673);
nand U9971 (N_9971,N_9723,N_9665);
nor U9972 (N_9972,N_9627,N_9651);
and U9973 (N_9973,N_9745,N_9711);
nor U9974 (N_9974,N_9668,N_9675);
and U9975 (N_9975,N_9799,N_9746);
nor U9976 (N_9976,N_9690,N_9745);
or U9977 (N_9977,N_9783,N_9754);
and U9978 (N_9978,N_9788,N_9762);
nor U9979 (N_9979,N_9776,N_9708);
xor U9980 (N_9980,N_9774,N_9666);
and U9981 (N_9981,N_9741,N_9796);
nor U9982 (N_9982,N_9709,N_9675);
nand U9983 (N_9983,N_9675,N_9654);
or U9984 (N_9984,N_9794,N_9733);
nand U9985 (N_9985,N_9644,N_9610);
nand U9986 (N_9986,N_9638,N_9689);
nand U9987 (N_9987,N_9657,N_9757);
nor U9988 (N_9988,N_9741,N_9775);
nor U9989 (N_9989,N_9652,N_9754);
nor U9990 (N_9990,N_9756,N_9659);
or U9991 (N_9991,N_9613,N_9707);
nand U9992 (N_9992,N_9769,N_9731);
and U9993 (N_9993,N_9746,N_9641);
and U9994 (N_9994,N_9764,N_9765);
nand U9995 (N_9995,N_9619,N_9723);
and U9996 (N_9996,N_9639,N_9697);
or U9997 (N_9997,N_9741,N_9650);
nand U9998 (N_9998,N_9647,N_9736);
or U9999 (N_9999,N_9792,N_9624);
or UO_0 (O_0,N_9980,N_9966);
or UO_1 (O_1,N_9876,N_9865);
nor UO_2 (O_2,N_9873,N_9904);
nor UO_3 (O_3,N_9956,N_9988);
and UO_4 (O_4,N_9998,N_9809);
and UO_5 (O_5,N_9983,N_9859);
or UO_6 (O_6,N_9926,N_9902);
and UO_7 (O_7,N_9829,N_9855);
or UO_8 (O_8,N_9977,N_9805);
nand UO_9 (O_9,N_9828,N_9995);
and UO_10 (O_10,N_9823,N_9981);
or UO_11 (O_11,N_9924,N_9950);
nand UO_12 (O_12,N_9802,N_9927);
nand UO_13 (O_13,N_9844,N_9922);
nor UO_14 (O_14,N_9882,N_9866);
or UO_15 (O_15,N_9960,N_9965);
nor UO_16 (O_16,N_9850,N_9817);
nand UO_17 (O_17,N_9948,N_9848);
and UO_18 (O_18,N_9888,N_9837);
nor UO_19 (O_19,N_9897,N_9812);
and UO_20 (O_20,N_9830,N_9874);
or UO_21 (O_21,N_9853,N_9991);
or UO_22 (O_22,N_9803,N_9879);
nand UO_23 (O_23,N_9908,N_9824);
nor UO_24 (O_24,N_9920,N_9916);
or UO_25 (O_25,N_9818,N_9893);
nor UO_26 (O_26,N_9861,N_9909);
nand UO_27 (O_27,N_9935,N_9880);
and UO_28 (O_28,N_9932,N_9834);
nor UO_29 (O_29,N_9886,N_9871);
and UO_30 (O_30,N_9870,N_9963);
nand UO_31 (O_31,N_9894,N_9890);
nand UO_32 (O_32,N_9964,N_9840);
and UO_33 (O_33,N_9816,N_9990);
or UO_34 (O_34,N_9936,N_9970);
nor UO_35 (O_35,N_9947,N_9934);
nand UO_36 (O_36,N_9946,N_9933);
nor UO_37 (O_37,N_9857,N_9978);
nand UO_38 (O_38,N_9962,N_9852);
nor UO_39 (O_39,N_9900,N_9898);
nor UO_40 (O_40,N_9953,N_9972);
nand UO_41 (O_41,N_9940,N_9910);
nand UO_42 (O_42,N_9832,N_9907);
nor UO_43 (O_43,N_9849,N_9942);
or UO_44 (O_44,N_9868,N_9842);
nor UO_45 (O_45,N_9919,N_9884);
and UO_46 (O_46,N_9811,N_9891);
and UO_47 (O_47,N_9961,N_9941);
nand UO_48 (O_48,N_9915,N_9808);
nand UO_49 (O_49,N_9885,N_9869);
xnor UO_50 (O_50,N_9913,N_9992);
or UO_51 (O_51,N_9839,N_9982);
and UO_52 (O_52,N_9826,N_9949);
or UO_53 (O_53,N_9958,N_9821);
and UO_54 (O_54,N_9863,N_9994);
nand UO_55 (O_55,N_9833,N_9892);
nor UO_56 (O_56,N_9928,N_9860);
and UO_57 (O_57,N_9917,N_9806);
nor UO_58 (O_58,N_9877,N_9971);
nand UO_59 (O_59,N_9820,N_9945);
nand UO_60 (O_60,N_9929,N_9836);
nand UO_61 (O_61,N_9923,N_9827);
or UO_62 (O_62,N_9896,N_9944);
or UO_63 (O_63,N_9867,N_9939);
xor UO_64 (O_64,N_9967,N_9810);
or UO_65 (O_65,N_9996,N_9841);
and UO_66 (O_66,N_9875,N_9957);
nand UO_67 (O_67,N_9921,N_9968);
or UO_68 (O_68,N_9985,N_9815);
and UO_69 (O_69,N_9851,N_9993);
or UO_70 (O_70,N_9847,N_9822);
nor UO_71 (O_71,N_9903,N_9911);
and UO_72 (O_72,N_9955,N_9872);
or UO_73 (O_73,N_9997,N_9952);
nand UO_74 (O_74,N_9987,N_9969);
nand UO_75 (O_75,N_9804,N_9835);
nor UO_76 (O_76,N_9856,N_9889);
nand UO_77 (O_77,N_9862,N_9846);
nand UO_78 (O_78,N_9979,N_9887);
or UO_79 (O_79,N_9954,N_9901);
nand UO_80 (O_80,N_9895,N_9925);
or UO_81 (O_81,N_9984,N_9864);
or UO_82 (O_82,N_9930,N_9831);
nand UO_83 (O_83,N_9906,N_9959);
and UO_84 (O_84,N_9905,N_9881);
nor UO_85 (O_85,N_9801,N_9899);
and UO_86 (O_86,N_9999,N_9813);
or UO_87 (O_87,N_9858,N_9974);
nand UO_88 (O_88,N_9800,N_9854);
or UO_89 (O_89,N_9937,N_9878);
nand UO_90 (O_90,N_9976,N_9918);
and UO_91 (O_91,N_9975,N_9914);
or UO_92 (O_92,N_9845,N_9825);
and UO_93 (O_93,N_9931,N_9938);
nor UO_94 (O_94,N_9989,N_9807);
nand UO_95 (O_95,N_9943,N_9883);
or UO_96 (O_96,N_9819,N_9838);
nand UO_97 (O_97,N_9814,N_9951);
nand UO_98 (O_98,N_9986,N_9912);
and UO_99 (O_99,N_9843,N_9973);
nand UO_100 (O_100,N_9931,N_9840);
or UO_101 (O_101,N_9951,N_9972);
nor UO_102 (O_102,N_9835,N_9855);
and UO_103 (O_103,N_9855,N_9867);
and UO_104 (O_104,N_9917,N_9847);
and UO_105 (O_105,N_9998,N_9859);
or UO_106 (O_106,N_9884,N_9956);
or UO_107 (O_107,N_9972,N_9913);
or UO_108 (O_108,N_9948,N_9995);
nor UO_109 (O_109,N_9924,N_9887);
nand UO_110 (O_110,N_9945,N_9808);
nand UO_111 (O_111,N_9936,N_9834);
nor UO_112 (O_112,N_9887,N_9850);
or UO_113 (O_113,N_9998,N_9866);
nand UO_114 (O_114,N_9826,N_9891);
and UO_115 (O_115,N_9817,N_9981);
nand UO_116 (O_116,N_9859,N_9825);
and UO_117 (O_117,N_9801,N_9900);
and UO_118 (O_118,N_9916,N_9931);
nand UO_119 (O_119,N_9868,N_9964);
nor UO_120 (O_120,N_9898,N_9928);
nor UO_121 (O_121,N_9882,N_9863);
nand UO_122 (O_122,N_9901,N_9988);
or UO_123 (O_123,N_9823,N_9987);
or UO_124 (O_124,N_9948,N_9917);
nor UO_125 (O_125,N_9834,N_9858);
nand UO_126 (O_126,N_9951,N_9829);
nand UO_127 (O_127,N_9834,N_9954);
or UO_128 (O_128,N_9925,N_9970);
nand UO_129 (O_129,N_9922,N_9927);
nor UO_130 (O_130,N_9952,N_9945);
and UO_131 (O_131,N_9843,N_9941);
nand UO_132 (O_132,N_9815,N_9875);
nor UO_133 (O_133,N_9984,N_9883);
nand UO_134 (O_134,N_9908,N_9812);
nor UO_135 (O_135,N_9922,N_9984);
nor UO_136 (O_136,N_9894,N_9980);
or UO_137 (O_137,N_9925,N_9933);
or UO_138 (O_138,N_9807,N_9927);
nand UO_139 (O_139,N_9911,N_9985);
nand UO_140 (O_140,N_9888,N_9882);
nor UO_141 (O_141,N_9875,N_9956);
nor UO_142 (O_142,N_9972,N_9987);
nor UO_143 (O_143,N_9999,N_9920);
or UO_144 (O_144,N_9845,N_9880);
xnor UO_145 (O_145,N_9913,N_9885);
or UO_146 (O_146,N_9926,N_9999);
nor UO_147 (O_147,N_9928,N_9960);
nand UO_148 (O_148,N_9988,N_9930);
nand UO_149 (O_149,N_9922,N_9924);
nor UO_150 (O_150,N_9901,N_9919);
or UO_151 (O_151,N_9901,N_9949);
or UO_152 (O_152,N_9846,N_9931);
nand UO_153 (O_153,N_9983,N_9933);
nand UO_154 (O_154,N_9909,N_9862);
and UO_155 (O_155,N_9853,N_9875);
nor UO_156 (O_156,N_9932,N_9990);
or UO_157 (O_157,N_9802,N_9839);
and UO_158 (O_158,N_9943,N_9925);
and UO_159 (O_159,N_9857,N_9975);
or UO_160 (O_160,N_9931,N_9920);
or UO_161 (O_161,N_9973,N_9808);
or UO_162 (O_162,N_9862,N_9885);
nand UO_163 (O_163,N_9958,N_9814);
or UO_164 (O_164,N_9909,N_9807);
nor UO_165 (O_165,N_9890,N_9972);
and UO_166 (O_166,N_9873,N_9815);
nor UO_167 (O_167,N_9939,N_9855);
or UO_168 (O_168,N_9997,N_9831);
or UO_169 (O_169,N_9980,N_9814);
nor UO_170 (O_170,N_9921,N_9991);
or UO_171 (O_171,N_9995,N_9912);
nand UO_172 (O_172,N_9941,N_9818);
nand UO_173 (O_173,N_9978,N_9841);
or UO_174 (O_174,N_9956,N_9849);
or UO_175 (O_175,N_9919,N_9922);
or UO_176 (O_176,N_9876,N_9908);
nand UO_177 (O_177,N_9962,N_9936);
or UO_178 (O_178,N_9864,N_9970);
and UO_179 (O_179,N_9974,N_9825);
and UO_180 (O_180,N_9994,N_9933);
or UO_181 (O_181,N_9844,N_9807);
xor UO_182 (O_182,N_9965,N_9913);
nor UO_183 (O_183,N_9860,N_9872);
or UO_184 (O_184,N_9855,N_9891);
xor UO_185 (O_185,N_9856,N_9914);
nor UO_186 (O_186,N_9815,N_9929);
nor UO_187 (O_187,N_9936,N_9906);
nand UO_188 (O_188,N_9986,N_9859);
nor UO_189 (O_189,N_9950,N_9965);
nor UO_190 (O_190,N_9977,N_9855);
nor UO_191 (O_191,N_9827,N_9844);
or UO_192 (O_192,N_9902,N_9889);
nor UO_193 (O_193,N_9819,N_9843);
or UO_194 (O_194,N_9985,N_9972);
nor UO_195 (O_195,N_9842,N_9800);
xnor UO_196 (O_196,N_9959,N_9810);
or UO_197 (O_197,N_9998,N_9967);
nor UO_198 (O_198,N_9848,N_9844);
nor UO_199 (O_199,N_9886,N_9922);
and UO_200 (O_200,N_9800,N_9869);
nor UO_201 (O_201,N_9804,N_9915);
and UO_202 (O_202,N_9860,N_9974);
nand UO_203 (O_203,N_9992,N_9971);
and UO_204 (O_204,N_9970,N_9861);
or UO_205 (O_205,N_9966,N_9914);
nor UO_206 (O_206,N_9808,N_9900);
nor UO_207 (O_207,N_9859,N_9995);
or UO_208 (O_208,N_9915,N_9975);
or UO_209 (O_209,N_9976,N_9925);
and UO_210 (O_210,N_9818,N_9957);
nand UO_211 (O_211,N_9853,N_9813);
and UO_212 (O_212,N_9957,N_9933);
nand UO_213 (O_213,N_9835,N_9935);
nor UO_214 (O_214,N_9915,N_9887);
or UO_215 (O_215,N_9901,N_9909);
nor UO_216 (O_216,N_9988,N_9923);
nand UO_217 (O_217,N_9993,N_9859);
and UO_218 (O_218,N_9943,N_9899);
or UO_219 (O_219,N_9953,N_9906);
and UO_220 (O_220,N_9833,N_9812);
and UO_221 (O_221,N_9902,N_9936);
nand UO_222 (O_222,N_9959,N_9964);
or UO_223 (O_223,N_9946,N_9853);
and UO_224 (O_224,N_9996,N_9842);
and UO_225 (O_225,N_9911,N_9842);
and UO_226 (O_226,N_9930,N_9961);
and UO_227 (O_227,N_9916,N_9977);
nor UO_228 (O_228,N_9885,N_9802);
or UO_229 (O_229,N_9952,N_9924);
xnor UO_230 (O_230,N_9942,N_9897);
nand UO_231 (O_231,N_9945,N_9965);
nand UO_232 (O_232,N_9838,N_9840);
nand UO_233 (O_233,N_9877,N_9960);
nand UO_234 (O_234,N_9905,N_9810);
and UO_235 (O_235,N_9930,N_9888);
or UO_236 (O_236,N_9904,N_9853);
nor UO_237 (O_237,N_9938,N_9851);
nor UO_238 (O_238,N_9826,N_9860);
and UO_239 (O_239,N_9956,N_9864);
nand UO_240 (O_240,N_9923,N_9899);
and UO_241 (O_241,N_9907,N_9897);
nor UO_242 (O_242,N_9939,N_9804);
nand UO_243 (O_243,N_9859,N_9942);
or UO_244 (O_244,N_9824,N_9815);
xnor UO_245 (O_245,N_9895,N_9911);
and UO_246 (O_246,N_9989,N_9980);
nand UO_247 (O_247,N_9894,N_9891);
or UO_248 (O_248,N_9825,N_9875);
and UO_249 (O_249,N_9925,N_9991);
nor UO_250 (O_250,N_9962,N_9801);
nor UO_251 (O_251,N_9849,N_9902);
nor UO_252 (O_252,N_9874,N_9905);
and UO_253 (O_253,N_9853,N_9997);
xor UO_254 (O_254,N_9830,N_9960);
nor UO_255 (O_255,N_9961,N_9900);
or UO_256 (O_256,N_9866,N_9847);
nand UO_257 (O_257,N_9909,N_9975);
nand UO_258 (O_258,N_9817,N_9920);
nor UO_259 (O_259,N_9824,N_9894);
xor UO_260 (O_260,N_9823,N_9906);
and UO_261 (O_261,N_9900,N_9890);
or UO_262 (O_262,N_9894,N_9991);
or UO_263 (O_263,N_9908,N_9954);
nand UO_264 (O_264,N_9875,N_9939);
xor UO_265 (O_265,N_9955,N_9927);
or UO_266 (O_266,N_9893,N_9947);
or UO_267 (O_267,N_9916,N_9893);
or UO_268 (O_268,N_9977,N_9981);
nor UO_269 (O_269,N_9946,N_9874);
and UO_270 (O_270,N_9835,N_9924);
nor UO_271 (O_271,N_9898,N_9902);
nand UO_272 (O_272,N_9920,N_9815);
nand UO_273 (O_273,N_9856,N_9967);
nand UO_274 (O_274,N_9825,N_9887);
nand UO_275 (O_275,N_9866,N_9912);
nor UO_276 (O_276,N_9894,N_9858);
and UO_277 (O_277,N_9907,N_9823);
nor UO_278 (O_278,N_9921,N_9910);
nand UO_279 (O_279,N_9833,N_9806);
nand UO_280 (O_280,N_9895,N_9897);
or UO_281 (O_281,N_9845,N_9964);
or UO_282 (O_282,N_9815,N_9934);
and UO_283 (O_283,N_9958,N_9818);
or UO_284 (O_284,N_9811,N_9969);
and UO_285 (O_285,N_9887,N_9912);
and UO_286 (O_286,N_9961,N_9989);
nand UO_287 (O_287,N_9914,N_9989);
nor UO_288 (O_288,N_9817,N_9990);
nand UO_289 (O_289,N_9999,N_9832);
nor UO_290 (O_290,N_9889,N_9996);
or UO_291 (O_291,N_9974,N_9947);
and UO_292 (O_292,N_9987,N_9912);
and UO_293 (O_293,N_9925,N_9876);
nor UO_294 (O_294,N_9979,N_9800);
and UO_295 (O_295,N_9846,N_9888);
and UO_296 (O_296,N_9901,N_9911);
or UO_297 (O_297,N_9915,N_9861);
and UO_298 (O_298,N_9938,N_9926);
or UO_299 (O_299,N_9959,N_9897);
nand UO_300 (O_300,N_9842,N_9856);
or UO_301 (O_301,N_9880,N_9849);
nand UO_302 (O_302,N_9925,N_9832);
nand UO_303 (O_303,N_9834,N_9920);
nor UO_304 (O_304,N_9956,N_9995);
nand UO_305 (O_305,N_9806,N_9995);
or UO_306 (O_306,N_9821,N_9890);
nor UO_307 (O_307,N_9989,N_9947);
nor UO_308 (O_308,N_9843,N_9806);
xnor UO_309 (O_309,N_9824,N_9922);
or UO_310 (O_310,N_9966,N_9863);
nand UO_311 (O_311,N_9808,N_9920);
and UO_312 (O_312,N_9956,N_9899);
nand UO_313 (O_313,N_9899,N_9807);
and UO_314 (O_314,N_9819,N_9903);
or UO_315 (O_315,N_9838,N_9994);
nand UO_316 (O_316,N_9969,N_9865);
nand UO_317 (O_317,N_9977,N_9820);
nand UO_318 (O_318,N_9985,N_9977);
nor UO_319 (O_319,N_9817,N_9993);
nor UO_320 (O_320,N_9808,N_9851);
or UO_321 (O_321,N_9876,N_9898);
and UO_322 (O_322,N_9964,N_9848);
and UO_323 (O_323,N_9856,N_9890);
and UO_324 (O_324,N_9826,N_9917);
xor UO_325 (O_325,N_9955,N_9928);
nor UO_326 (O_326,N_9956,N_9920);
and UO_327 (O_327,N_9929,N_9976);
nand UO_328 (O_328,N_9816,N_9995);
and UO_329 (O_329,N_9836,N_9810);
and UO_330 (O_330,N_9818,N_9919);
and UO_331 (O_331,N_9925,N_9926);
nand UO_332 (O_332,N_9912,N_9844);
or UO_333 (O_333,N_9886,N_9931);
and UO_334 (O_334,N_9842,N_9907);
nor UO_335 (O_335,N_9818,N_9948);
and UO_336 (O_336,N_9878,N_9858);
nand UO_337 (O_337,N_9950,N_9840);
nand UO_338 (O_338,N_9945,N_9887);
or UO_339 (O_339,N_9980,N_9905);
or UO_340 (O_340,N_9822,N_9824);
nor UO_341 (O_341,N_9906,N_9885);
nand UO_342 (O_342,N_9820,N_9902);
nand UO_343 (O_343,N_9896,N_9877);
and UO_344 (O_344,N_9887,N_9866);
nand UO_345 (O_345,N_9899,N_9959);
nor UO_346 (O_346,N_9971,N_9825);
nand UO_347 (O_347,N_9888,N_9898);
nand UO_348 (O_348,N_9969,N_9983);
and UO_349 (O_349,N_9895,N_9918);
or UO_350 (O_350,N_9870,N_9880);
nor UO_351 (O_351,N_9883,N_9895);
and UO_352 (O_352,N_9867,N_9844);
or UO_353 (O_353,N_9953,N_9934);
or UO_354 (O_354,N_9987,N_9898);
or UO_355 (O_355,N_9800,N_9927);
nand UO_356 (O_356,N_9891,N_9902);
nand UO_357 (O_357,N_9874,N_9863);
nand UO_358 (O_358,N_9994,N_9964);
and UO_359 (O_359,N_9851,N_9831);
nor UO_360 (O_360,N_9828,N_9980);
nor UO_361 (O_361,N_9845,N_9978);
or UO_362 (O_362,N_9828,N_9866);
and UO_363 (O_363,N_9804,N_9894);
or UO_364 (O_364,N_9970,N_9836);
or UO_365 (O_365,N_9984,N_9865);
or UO_366 (O_366,N_9938,N_9836);
nor UO_367 (O_367,N_9811,N_9876);
nor UO_368 (O_368,N_9830,N_9912);
nor UO_369 (O_369,N_9941,N_9884);
and UO_370 (O_370,N_9958,N_9890);
nor UO_371 (O_371,N_9848,N_9857);
and UO_372 (O_372,N_9814,N_9983);
and UO_373 (O_373,N_9830,N_9931);
nor UO_374 (O_374,N_9930,N_9876);
nor UO_375 (O_375,N_9930,N_9921);
nor UO_376 (O_376,N_9982,N_9860);
or UO_377 (O_377,N_9862,N_9933);
or UO_378 (O_378,N_9907,N_9997);
nor UO_379 (O_379,N_9870,N_9876);
or UO_380 (O_380,N_9961,N_9892);
or UO_381 (O_381,N_9861,N_9964);
xnor UO_382 (O_382,N_9871,N_9907);
xnor UO_383 (O_383,N_9855,N_9857);
and UO_384 (O_384,N_9975,N_9953);
nand UO_385 (O_385,N_9986,N_9867);
or UO_386 (O_386,N_9941,N_9812);
nor UO_387 (O_387,N_9963,N_9936);
and UO_388 (O_388,N_9802,N_9877);
nand UO_389 (O_389,N_9923,N_9998);
nor UO_390 (O_390,N_9918,N_9887);
or UO_391 (O_391,N_9961,N_9927);
and UO_392 (O_392,N_9986,N_9994);
nand UO_393 (O_393,N_9916,N_9824);
and UO_394 (O_394,N_9896,N_9851);
nor UO_395 (O_395,N_9831,N_9954);
nor UO_396 (O_396,N_9947,N_9982);
nand UO_397 (O_397,N_9911,N_9992);
nor UO_398 (O_398,N_9901,N_9972);
nor UO_399 (O_399,N_9861,N_9932);
and UO_400 (O_400,N_9889,N_9813);
nor UO_401 (O_401,N_9988,N_9995);
and UO_402 (O_402,N_9916,N_9868);
or UO_403 (O_403,N_9992,N_9866);
nor UO_404 (O_404,N_9966,N_9906);
nor UO_405 (O_405,N_9901,N_9817);
or UO_406 (O_406,N_9807,N_9963);
or UO_407 (O_407,N_9893,N_9869);
xor UO_408 (O_408,N_9917,N_9844);
and UO_409 (O_409,N_9919,N_9971);
and UO_410 (O_410,N_9825,N_9929);
nor UO_411 (O_411,N_9865,N_9899);
nor UO_412 (O_412,N_9878,N_9821);
or UO_413 (O_413,N_9894,N_9854);
or UO_414 (O_414,N_9958,N_9995);
nor UO_415 (O_415,N_9902,N_9811);
nand UO_416 (O_416,N_9908,N_9936);
or UO_417 (O_417,N_9864,N_9965);
nor UO_418 (O_418,N_9927,N_9935);
and UO_419 (O_419,N_9879,N_9980);
nor UO_420 (O_420,N_9919,N_9940);
and UO_421 (O_421,N_9918,N_9995);
nand UO_422 (O_422,N_9897,N_9988);
nor UO_423 (O_423,N_9824,N_9973);
and UO_424 (O_424,N_9938,N_9829);
or UO_425 (O_425,N_9823,N_9811);
or UO_426 (O_426,N_9996,N_9959);
nand UO_427 (O_427,N_9920,N_9986);
or UO_428 (O_428,N_9892,N_9970);
nor UO_429 (O_429,N_9967,N_9994);
nor UO_430 (O_430,N_9806,N_9994);
nand UO_431 (O_431,N_9952,N_9963);
nor UO_432 (O_432,N_9975,N_9965);
nand UO_433 (O_433,N_9984,N_9923);
xor UO_434 (O_434,N_9998,N_9810);
or UO_435 (O_435,N_9884,N_9966);
nand UO_436 (O_436,N_9919,N_9923);
nor UO_437 (O_437,N_9877,N_9911);
nand UO_438 (O_438,N_9843,N_9839);
nor UO_439 (O_439,N_9852,N_9858);
and UO_440 (O_440,N_9896,N_9823);
or UO_441 (O_441,N_9801,N_9844);
nand UO_442 (O_442,N_9897,N_9801);
and UO_443 (O_443,N_9803,N_9947);
or UO_444 (O_444,N_9811,N_9806);
and UO_445 (O_445,N_9949,N_9945);
or UO_446 (O_446,N_9913,N_9906);
nor UO_447 (O_447,N_9866,N_9853);
and UO_448 (O_448,N_9933,N_9936);
or UO_449 (O_449,N_9931,N_9974);
nand UO_450 (O_450,N_9861,N_9917);
or UO_451 (O_451,N_9918,N_9916);
nand UO_452 (O_452,N_9974,N_9927);
nand UO_453 (O_453,N_9911,N_9821);
nor UO_454 (O_454,N_9969,N_9830);
or UO_455 (O_455,N_9901,N_9850);
nand UO_456 (O_456,N_9968,N_9974);
nand UO_457 (O_457,N_9971,N_9842);
or UO_458 (O_458,N_9931,N_9885);
xnor UO_459 (O_459,N_9979,N_9995);
xnor UO_460 (O_460,N_9967,N_9861);
nor UO_461 (O_461,N_9876,N_9996);
and UO_462 (O_462,N_9810,N_9918);
or UO_463 (O_463,N_9874,N_9913);
or UO_464 (O_464,N_9835,N_9919);
or UO_465 (O_465,N_9847,N_9900);
nor UO_466 (O_466,N_9927,N_9933);
nor UO_467 (O_467,N_9971,N_9918);
nor UO_468 (O_468,N_9883,N_9967);
nor UO_469 (O_469,N_9924,N_9847);
nor UO_470 (O_470,N_9806,N_9830);
nor UO_471 (O_471,N_9965,N_9955);
nor UO_472 (O_472,N_9800,N_9817);
or UO_473 (O_473,N_9801,N_9949);
and UO_474 (O_474,N_9895,N_9888);
nand UO_475 (O_475,N_9817,N_9825);
nand UO_476 (O_476,N_9865,N_9944);
or UO_477 (O_477,N_9894,N_9992);
nor UO_478 (O_478,N_9885,N_9809);
xor UO_479 (O_479,N_9887,N_9910);
and UO_480 (O_480,N_9923,N_9973);
or UO_481 (O_481,N_9800,N_9845);
nor UO_482 (O_482,N_9826,N_9946);
nor UO_483 (O_483,N_9806,N_9867);
nand UO_484 (O_484,N_9982,N_9995);
nor UO_485 (O_485,N_9987,N_9834);
nand UO_486 (O_486,N_9939,N_9868);
or UO_487 (O_487,N_9970,N_9878);
nand UO_488 (O_488,N_9951,N_9908);
nand UO_489 (O_489,N_9850,N_9835);
or UO_490 (O_490,N_9822,N_9919);
and UO_491 (O_491,N_9859,N_9934);
and UO_492 (O_492,N_9978,N_9862);
and UO_493 (O_493,N_9905,N_9871);
nor UO_494 (O_494,N_9958,N_9893);
or UO_495 (O_495,N_9938,N_9868);
or UO_496 (O_496,N_9947,N_9858);
or UO_497 (O_497,N_9830,N_9937);
and UO_498 (O_498,N_9916,N_9961);
or UO_499 (O_499,N_9837,N_9824);
and UO_500 (O_500,N_9816,N_9964);
and UO_501 (O_501,N_9977,N_9897);
or UO_502 (O_502,N_9998,N_9834);
or UO_503 (O_503,N_9821,N_9809);
or UO_504 (O_504,N_9816,N_9803);
and UO_505 (O_505,N_9923,N_9954);
or UO_506 (O_506,N_9922,N_9997);
or UO_507 (O_507,N_9991,N_9899);
nor UO_508 (O_508,N_9973,N_9888);
nand UO_509 (O_509,N_9800,N_9823);
or UO_510 (O_510,N_9972,N_9962);
and UO_511 (O_511,N_9817,N_9942);
or UO_512 (O_512,N_9934,N_9862);
and UO_513 (O_513,N_9886,N_9918);
nor UO_514 (O_514,N_9881,N_9999);
or UO_515 (O_515,N_9998,N_9840);
or UO_516 (O_516,N_9830,N_9837);
nand UO_517 (O_517,N_9875,N_9864);
nor UO_518 (O_518,N_9960,N_9936);
and UO_519 (O_519,N_9895,N_9942);
or UO_520 (O_520,N_9824,N_9899);
nor UO_521 (O_521,N_9897,N_9800);
and UO_522 (O_522,N_9893,N_9812);
nor UO_523 (O_523,N_9913,N_9899);
nand UO_524 (O_524,N_9808,N_9977);
or UO_525 (O_525,N_9992,N_9897);
and UO_526 (O_526,N_9807,N_9920);
nand UO_527 (O_527,N_9930,N_9919);
nor UO_528 (O_528,N_9831,N_9818);
and UO_529 (O_529,N_9895,N_9877);
nand UO_530 (O_530,N_9998,N_9885);
nor UO_531 (O_531,N_9845,N_9885);
or UO_532 (O_532,N_9841,N_9808);
nor UO_533 (O_533,N_9838,N_9959);
or UO_534 (O_534,N_9902,N_9860);
nand UO_535 (O_535,N_9902,N_9966);
and UO_536 (O_536,N_9883,N_9985);
nand UO_537 (O_537,N_9824,N_9811);
nor UO_538 (O_538,N_9920,N_9801);
nor UO_539 (O_539,N_9925,N_9808);
and UO_540 (O_540,N_9826,N_9838);
and UO_541 (O_541,N_9915,N_9899);
and UO_542 (O_542,N_9995,N_9889);
nor UO_543 (O_543,N_9960,N_9875);
nand UO_544 (O_544,N_9915,N_9916);
or UO_545 (O_545,N_9899,N_9908);
and UO_546 (O_546,N_9881,N_9810);
nand UO_547 (O_547,N_9892,N_9995);
or UO_548 (O_548,N_9890,N_9839);
and UO_549 (O_549,N_9941,N_9943);
or UO_550 (O_550,N_9895,N_9858);
nand UO_551 (O_551,N_9996,N_9948);
or UO_552 (O_552,N_9842,N_9865);
or UO_553 (O_553,N_9880,N_9906);
or UO_554 (O_554,N_9876,N_9992);
or UO_555 (O_555,N_9888,N_9901);
and UO_556 (O_556,N_9820,N_9803);
nor UO_557 (O_557,N_9901,N_9940);
nand UO_558 (O_558,N_9848,N_9831);
nand UO_559 (O_559,N_9960,N_9825);
nor UO_560 (O_560,N_9860,N_9856);
nand UO_561 (O_561,N_9905,N_9828);
and UO_562 (O_562,N_9800,N_9838);
nand UO_563 (O_563,N_9869,N_9803);
and UO_564 (O_564,N_9820,N_9859);
and UO_565 (O_565,N_9863,N_9922);
xor UO_566 (O_566,N_9881,N_9990);
and UO_567 (O_567,N_9874,N_9964);
or UO_568 (O_568,N_9811,N_9914);
nand UO_569 (O_569,N_9813,N_9850);
nand UO_570 (O_570,N_9859,N_9856);
nor UO_571 (O_571,N_9985,N_9865);
and UO_572 (O_572,N_9828,N_9805);
nor UO_573 (O_573,N_9883,N_9899);
and UO_574 (O_574,N_9887,N_9953);
nand UO_575 (O_575,N_9988,N_9816);
nand UO_576 (O_576,N_9876,N_9887);
or UO_577 (O_577,N_9971,N_9928);
nand UO_578 (O_578,N_9882,N_9871);
nor UO_579 (O_579,N_9845,N_9884);
nand UO_580 (O_580,N_9837,N_9863);
nor UO_581 (O_581,N_9832,N_9885);
nand UO_582 (O_582,N_9973,N_9906);
or UO_583 (O_583,N_9932,N_9997);
and UO_584 (O_584,N_9849,N_9802);
nor UO_585 (O_585,N_9981,N_9805);
or UO_586 (O_586,N_9806,N_9844);
nor UO_587 (O_587,N_9828,N_9983);
or UO_588 (O_588,N_9947,N_9907);
or UO_589 (O_589,N_9875,N_9897);
and UO_590 (O_590,N_9985,N_9819);
or UO_591 (O_591,N_9864,N_9975);
nand UO_592 (O_592,N_9808,N_9850);
or UO_593 (O_593,N_9977,N_9803);
nand UO_594 (O_594,N_9871,N_9857);
nand UO_595 (O_595,N_9966,N_9888);
nor UO_596 (O_596,N_9889,N_9924);
nand UO_597 (O_597,N_9889,N_9820);
and UO_598 (O_598,N_9866,N_9818);
or UO_599 (O_599,N_9912,N_9875);
and UO_600 (O_600,N_9938,N_9974);
nor UO_601 (O_601,N_9917,N_9918);
nor UO_602 (O_602,N_9880,N_9946);
and UO_603 (O_603,N_9801,N_9979);
or UO_604 (O_604,N_9922,N_9973);
or UO_605 (O_605,N_9959,N_9910);
and UO_606 (O_606,N_9875,N_9996);
nor UO_607 (O_607,N_9901,N_9945);
nand UO_608 (O_608,N_9899,N_9988);
and UO_609 (O_609,N_9906,N_9905);
nand UO_610 (O_610,N_9960,N_9887);
nand UO_611 (O_611,N_9895,N_9868);
nor UO_612 (O_612,N_9930,N_9947);
nand UO_613 (O_613,N_9884,N_9852);
nand UO_614 (O_614,N_9972,N_9970);
or UO_615 (O_615,N_9821,N_9981);
or UO_616 (O_616,N_9967,N_9836);
or UO_617 (O_617,N_9872,N_9896);
nor UO_618 (O_618,N_9975,N_9940);
nor UO_619 (O_619,N_9937,N_9875);
or UO_620 (O_620,N_9839,N_9966);
nand UO_621 (O_621,N_9853,N_9871);
nor UO_622 (O_622,N_9864,N_9947);
or UO_623 (O_623,N_9968,N_9884);
and UO_624 (O_624,N_9958,N_9956);
or UO_625 (O_625,N_9893,N_9976);
nand UO_626 (O_626,N_9971,N_9935);
xnor UO_627 (O_627,N_9851,N_9992);
nand UO_628 (O_628,N_9877,N_9934);
xnor UO_629 (O_629,N_9968,N_9965);
nand UO_630 (O_630,N_9980,N_9854);
nor UO_631 (O_631,N_9930,N_9972);
and UO_632 (O_632,N_9917,N_9800);
nor UO_633 (O_633,N_9891,N_9883);
nand UO_634 (O_634,N_9803,N_9969);
or UO_635 (O_635,N_9897,N_9955);
or UO_636 (O_636,N_9830,N_9917);
nand UO_637 (O_637,N_9957,N_9913);
and UO_638 (O_638,N_9873,N_9925);
and UO_639 (O_639,N_9903,N_9901);
nor UO_640 (O_640,N_9834,N_9964);
nor UO_641 (O_641,N_9915,N_9983);
and UO_642 (O_642,N_9878,N_9945);
nand UO_643 (O_643,N_9975,N_9937);
nor UO_644 (O_644,N_9807,N_9992);
nor UO_645 (O_645,N_9871,N_9912);
nor UO_646 (O_646,N_9917,N_9933);
nand UO_647 (O_647,N_9956,N_9972);
and UO_648 (O_648,N_9931,N_9991);
nand UO_649 (O_649,N_9877,N_9853);
nor UO_650 (O_650,N_9934,N_9955);
and UO_651 (O_651,N_9892,N_9907);
or UO_652 (O_652,N_9895,N_9853);
or UO_653 (O_653,N_9942,N_9827);
nand UO_654 (O_654,N_9909,N_9911);
or UO_655 (O_655,N_9865,N_9868);
or UO_656 (O_656,N_9821,N_9889);
nand UO_657 (O_657,N_9916,N_9983);
or UO_658 (O_658,N_9976,N_9803);
or UO_659 (O_659,N_9910,N_9954);
nand UO_660 (O_660,N_9885,N_9841);
or UO_661 (O_661,N_9803,N_9861);
xnor UO_662 (O_662,N_9994,N_9962);
and UO_663 (O_663,N_9942,N_9909);
nor UO_664 (O_664,N_9820,N_9986);
or UO_665 (O_665,N_9960,N_9998);
or UO_666 (O_666,N_9971,N_9941);
nor UO_667 (O_667,N_9916,N_9946);
nor UO_668 (O_668,N_9844,N_9940);
and UO_669 (O_669,N_9837,N_9991);
and UO_670 (O_670,N_9929,N_9834);
and UO_671 (O_671,N_9835,N_9831);
and UO_672 (O_672,N_9873,N_9907);
nor UO_673 (O_673,N_9900,N_9838);
nor UO_674 (O_674,N_9929,N_9995);
nor UO_675 (O_675,N_9936,N_9914);
or UO_676 (O_676,N_9815,N_9836);
nor UO_677 (O_677,N_9895,N_9983);
nand UO_678 (O_678,N_9966,N_9866);
nand UO_679 (O_679,N_9848,N_9835);
or UO_680 (O_680,N_9931,N_9936);
nor UO_681 (O_681,N_9960,N_9994);
or UO_682 (O_682,N_9844,N_9838);
nand UO_683 (O_683,N_9847,N_9857);
nand UO_684 (O_684,N_9977,N_9813);
nand UO_685 (O_685,N_9966,N_9996);
and UO_686 (O_686,N_9868,N_9830);
or UO_687 (O_687,N_9844,N_9953);
nand UO_688 (O_688,N_9800,N_9989);
and UO_689 (O_689,N_9962,N_9842);
and UO_690 (O_690,N_9897,N_9888);
nand UO_691 (O_691,N_9912,N_9894);
and UO_692 (O_692,N_9858,N_9840);
nand UO_693 (O_693,N_9896,N_9866);
and UO_694 (O_694,N_9897,N_9813);
or UO_695 (O_695,N_9960,N_9811);
nor UO_696 (O_696,N_9941,N_9860);
nor UO_697 (O_697,N_9908,N_9804);
nor UO_698 (O_698,N_9889,N_9842);
nor UO_699 (O_699,N_9968,N_9817);
and UO_700 (O_700,N_9902,N_9912);
and UO_701 (O_701,N_9825,N_9864);
nand UO_702 (O_702,N_9855,N_9944);
nor UO_703 (O_703,N_9968,N_9843);
or UO_704 (O_704,N_9984,N_9829);
and UO_705 (O_705,N_9837,N_9879);
nor UO_706 (O_706,N_9831,N_9948);
and UO_707 (O_707,N_9855,N_9842);
nand UO_708 (O_708,N_9934,N_9838);
nand UO_709 (O_709,N_9906,N_9979);
or UO_710 (O_710,N_9995,N_9921);
nor UO_711 (O_711,N_9857,N_9832);
nand UO_712 (O_712,N_9882,N_9927);
and UO_713 (O_713,N_9810,N_9896);
and UO_714 (O_714,N_9953,N_9952);
nand UO_715 (O_715,N_9986,N_9913);
nor UO_716 (O_716,N_9821,N_9935);
and UO_717 (O_717,N_9939,N_9935);
and UO_718 (O_718,N_9924,N_9911);
nand UO_719 (O_719,N_9887,N_9984);
nand UO_720 (O_720,N_9957,N_9953);
nand UO_721 (O_721,N_9857,N_9854);
or UO_722 (O_722,N_9857,N_9809);
nand UO_723 (O_723,N_9868,N_9941);
nor UO_724 (O_724,N_9812,N_9854);
or UO_725 (O_725,N_9800,N_9950);
and UO_726 (O_726,N_9940,N_9921);
or UO_727 (O_727,N_9871,N_9838);
or UO_728 (O_728,N_9989,N_9885);
and UO_729 (O_729,N_9955,N_9960);
or UO_730 (O_730,N_9823,N_9850);
and UO_731 (O_731,N_9878,N_9814);
nor UO_732 (O_732,N_9821,N_9859);
or UO_733 (O_733,N_9964,N_9893);
nor UO_734 (O_734,N_9926,N_9874);
nand UO_735 (O_735,N_9978,N_9901);
and UO_736 (O_736,N_9817,N_9962);
nor UO_737 (O_737,N_9834,N_9940);
nand UO_738 (O_738,N_9832,N_9892);
and UO_739 (O_739,N_9897,N_9823);
xor UO_740 (O_740,N_9978,N_9813);
nor UO_741 (O_741,N_9947,N_9938);
nor UO_742 (O_742,N_9966,N_9986);
and UO_743 (O_743,N_9879,N_9801);
and UO_744 (O_744,N_9805,N_9903);
nand UO_745 (O_745,N_9957,N_9934);
or UO_746 (O_746,N_9937,N_9802);
nand UO_747 (O_747,N_9895,N_9826);
nand UO_748 (O_748,N_9867,N_9858);
and UO_749 (O_749,N_9847,N_9915);
nand UO_750 (O_750,N_9848,N_9893);
and UO_751 (O_751,N_9838,N_9842);
or UO_752 (O_752,N_9999,N_9960);
nor UO_753 (O_753,N_9931,N_9898);
or UO_754 (O_754,N_9812,N_9832);
or UO_755 (O_755,N_9834,N_9826);
nand UO_756 (O_756,N_9830,N_9982);
xor UO_757 (O_757,N_9816,N_9920);
nor UO_758 (O_758,N_9987,N_9917);
nand UO_759 (O_759,N_9865,N_9979);
and UO_760 (O_760,N_9824,N_9979);
nand UO_761 (O_761,N_9872,N_9969);
nand UO_762 (O_762,N_9833,N_9858);
nor UO_763 (O_763,N_9854,N_9865);
nor UO_764 (O_764,N_9836,N_9971);
and UO_765 (O_765,N_9974,N_9964);
nor UO_766 (O_766,N_9836,N_9904);
nor UO_767 (O_767,N_9979,N_9805);
or UO_768 (O_768,N_9830,N_9926);
or UO_769 (O_769,N_9860,N_9948);
and UO_770 (O_770,N_9989,N_9970);
and UO_771 (O_771,N_9804,N_9861);
and UO_772 (O_772,N_9915,N_9935);
and UO_773 (O_773,N_9939,N_9852);
or UO_774 (O_774,N_9847,N_9853);
nand UO_775 (O_775,N_9976,N_9938);
nand UO_776 (O_776,N_9980,N_9895);
nand UO_777 (O_777,N_9942,N_9978);
xnor UO_778 (O_778,N_9909,N_9823);
and UO_779 (O_779,N_9810,N_9909);
nand UO_780 (O_780,N_9924,N_9918);
or UO_781 (O_781,N_9822,N_9961);
nor UO_782 (O_782,N_9993,N_9952);
nor UO_783 (O_783,N_9816,N_9922);
xor UO_784 (O_784,N_9859,N_9915);
and UO_785 (O_785,N_9918,N_9932);
nor UO_786 (O_786,N_9935,N_9954);
or UO_787 (O_787,N_9969,N_9933);
or UO_788 (O_788,N_9829,N_9843);
and UO_789 (O_789,N_9977,N_9943);
or UO_790 (O_790,N_9813,N_9854);
nor UO_791 (O_791,N_9860,N_9838);
and UO_792 (O_792,N_9904,N_9857);
or UO_793 (O_793,N_9972,N_9875);
and UO_794 (O_794,N_9976,N_9826);
nor UO_795 (O_795,N_9890,N_9955);
nor UO_796 (O_796,N_9999,N_9847);
nand UO_797 (O_797,N_9919,N_9910);
nor UO_798 (O_798,N_9874,N_9930);
nand UO_799 (O_799,N_9854,N_9900);
nor UO_800 (O_800,N_9809,N_9853);
and UO_801 (O_801,N_9949,N_9815);
and UO_802 (O_802,N_9859,N_9956);
nor UO_803 (O_803,N_9886,N_9961);
and UO_804 (O_804,N_9898,N_9843);
nor UO_805 (O_805,N_9803,N_9986);
or UO_806 (O_806,N_9985,N_9807);
or UO_807 (O_807,N_9862,N_9929);
and UO_808 (O_808,N_9943,N_9948);
or UO_809 (O_809,N_9872,N_9808);
nor UO_810 (O_810,N_9867,N_9843);
and UO_811 (O_811,N_9828,N_9998);
or UO_812 (O_812,N_9801,N_9973);
nand UO_813 (O_813,N_9987,N_9843);
nand UO_814 (O_814,N_9846,N_9803);
and UO_815 (O_815,N_9952,N_9916);
or UO_816 (O_816,N_9840,N_9859);
nor UO_817 (O_817,N_9825,N_9861);
nor UO_818 (O_818,N_9846,N_9896);
nand UO_819 (O_819,N_9941,N_9875);
nor UO_820 (O_820,N_9873,N_9960);
xor UO_821 (O_821,N_9950,N_9887);
nand UO_822 (O_822,N_9821,N_9954);
and UO_823 (O_823,N_9962,N_9952);
and UO_824 (O_824,N_9819,N_9883);
or UO_825 (O_825,N_9945,N_9847);
xnor UO_826 (O_826,N_9895,N_9863);
and UO_827 (O_827,N_9897,N_9844);
nand UO_828 (O_828,N_9825,N_9936);
or UO_829 (O_829,N_9808,N_9958);
and UO_830 (O_830,N_9882,N_9941);
nand UO_831 (O_831,N_9818,N_9965);
nor UO_832 (O_832,N_9945,N_9953);
nand UO_833 (O_833,N_9840,N_9817);
and UO_834 (O_834,N_9993,N_9867);
nand UO_835 (O_835,N_9826,N_9958);
nand UO_836 (O_836,N_9922,N_9831);
nand UO_837 (O_837,N_9953,N_9940);
nor UO_838 (O_838,N_9985,N_9917);
or UO_839 (O_839,N_9907,N_9992);
xnor UO_840 (O_840,N_9921,N_9858);
and UO_841 (O_841,N_9951,N_9983);
nor UO_842 (O_842,N_9834,N_9825);
nor UO_843 (O_843,N_9978,N_9816);
or UO_844 (O_844,N_9838,N_9912);
nand UO_845 (O_845,N_9992,N_9944);
nor UO_846 (O_846,N_9869,N_9892);
and UO_847 (O_847,N_9896,N_9928);
and UO_848 (O_848,N_9967,N_9893);
nor UO_849 (O_849,N_9862,N_9942);
and UO_850 (O_850,N_9873,N_9924);
and UO_851 (O_851,N_9816,N_9818);
and UO_852 (O_852,N_9950,N_9830);
and UO_853 (O_853,N_9861,N_9939);
and UO_854 (O_854,N_9976,N_9984);
and UO_855 (O_855,N_9878,N_9823);
or UO_856 (O_856,N_9979,N_9996);
and UO_857 (O_857,N_9850,N_9934);
nand UO_858 (O_858,N_9886,N_9809);
nor UO_859 (O_859,N_9824,N_9888);
and UO_860 (O_860,N_9957,N_9805);
or UO_861 (O_861,N_9855,N_9859);
and UO_862 (O_862,N_9906,N_9927);
nor UO_863 (O_863,N_9990,N_9902);
nor UO_864 (O_864,N_9925,N_9807);
xnor UO_865 (O_865,N_9983,N_9922);
and UO_866 (O_866,N_9986,N_9985);
and UO_867 (O_867,N_9835,N_9922);
and UO_868 (O_868,N_9813,N_9965);
nand UO_869 (O_869,N_9812,N_9903);
nor UO_870 (O_870,N_9961,N_9840);
and UO_871 (O_871,N_9990,N_9950);
or UO_872 (O_872,N_9928,N_9825);
xor UO_873 (O_873,N_9992,N_9808);
and UO_874 (O_874,N_9899,N_9955);
nor UO_875 (O_875,N_9827,N_9852);
nor UO_876 (O_876,N_9865,N_9947);
and UO_877 (O_877,N_9933,N_9801);
or UO_878 (O_878,N_9858,N_9935);
nor UO_879 (O_879,N_9895,N_9805);
xnor UO_880 (O_880,N_9960,N_9874);
nor UO_881 (O_881,N_9981,N_9972);
or UO_882 (O_882,N_9954,N_9941);
nand UO_883 (O_883,N_9830,N_9855);
or UO_884 (O_884,N_9909,N_9924);
nand UO_885 (O_885,N_9904,N_9833);
nor UO_886 (O_886,N_9942,N_9858);
xnor UO_887 (O_887,N_9802,N_9998);
or UO_888 (O_888,N_9853,N_9876);
or UO_889 (O_889,N_9894,N_9870);
or UO_890 (O_890,N_9977,N_9889);
nand UO_891 (O_891,N_9981,N_9964);
or UO_892 (O_892,N_9954,N_9944);
and UO_893 (O_893,N_9987,N_9857);
and UO_894 (O_894,N_9845,N_9986);
or UO_895 (O_895,N_9908,N_9997);
nor UO_896 (O_896,N_9808,N_9939);
or UO_897 (O_897,N_9867,N_9950);
nor UO_898 (O_898,N_9867,N_9906);
nand UO_899 (O_899,N_9823,N_9864);
and UO_900 (O_900,N_9810,N_9996);
or UO_901 (O_901,N_9898,N_9882);
nand UO_902 (O_902,N_9994,N_9860);
nor UO_903 (O_903,N_9906,N_9816);
or UO_904 (O_904,N_9987,N_9955);
nor UO_905 (O_905,N_9940,N_9895);
nor UO_906 (O_906,N_9803,N_9953);
and UO_907 (O_907,N_9876,N_9816);
xnor UO_908 (O_908,N_9933,N_9845);
nor UO_909 (O_909,N_9841,N_9999);
nor UO_910 (O_910,N_9954,N_9925);
and UO_911 (O_911,N_9971,N_9872);
and UO_912 (O_912,N_9904,N_9985);
nand UO_913 (O_913,N_9867,N_9946);
nand UO_914 (O_914,N_9875,N_9834);
nand UO_915 (O_915,N_9841,N_9835);
nor UO_916 (O_916,N_9834,N_9949);
or UO_917 (O_917,N_9987,N_9991);
nand UO_918 (O_918,N_9891,N_9906);
and UO_919 (O_919,N_9819,N_9900);
nand UO_920 (O_920,N_9958,N_9915);
nor UO_921 (O_921,N_9854,N_9952);
and UO_922 (O_922,N_9815,N_9901);
or UO_923 (O_923,N_9877,N_9968);
nand UO_924 (O_924,N_9807,N_9843);
or UO_925 (O_925,N_9959,N_9876);
and UO_926 (O_926,N_9808,N_9950);
nor UO_927 (O_927,N_9817,N_9890);
nor UO_928 (O_928,N_9824,N_9910);
nand UO_929 (O_929,N_9817,N_9999);
or UO_930 (O_930,N_9966,N_9832);
or UO_931 (O_931,N_9831,N_9896);
and UO_932 (O_932,N_9850,N_9909);
nor UO_933 (O_933,N_9981,N_9973);
and UO_934 (O_934,N_9880,N_9812);
and UO_935 (O_935,N_9921,N_9848);
or UO_936 (O_936,N_9983,N_9942);
and UO_937 (O_937,N_9890,N_9995);
or UO_938 (O_938,N_9973,N_9900);
nor UO_939 (O_939,N_9961,N_9803);
nand UO_940 (O_940,N_9804,N_9906);
and UO_941 (O_941,N_9974,N_9826);
or UO_942 (O_942,N_9933,N_9968);
or UO_943 (O_943,N_9930,N_9875);
nand UO_944 (O_944,N_9830,N_9983);
nand UO_945 (O_945,N_9944,N_9829);
nor UO_946 (O_946,N_9932,N_9902);
or UO_947 (O_947,N_9879,N_9884);
nand UO_948 (O_948,N_9959,N_9940);
or UO_949 (O_949,N_9950,N_9847);
nand UO_950 (O_950,N_9923,N_9947);
or UO_951 (O_951,N_9809,N_9831);
or UO_952 (O_952,N_9913,N_9970);
nand UO_953 (O_953,N_9953,N_9810);
and UO_954 (O_954,N_9957,N_9937);
or UO_955 (O_955,N_9874,N_9851);
and UO_956 (O_956,N_9934,N_9840);
nand UO_957 (O_957,N_9845,N_9996);
or UO_958 (O_958,N_9923,N_9862);
or UO_959 (O_959,N_9960,N_9946);
nor UO_960 (O_960,N_9983,N_9882);
and UO_961 (O_961,N_9857,N_9914);
xor UO_962 (O_962,N_9851,N_9823);
nor UO_963 (O_963,N_9906,N_9978);
and UO_964 (O_964,N_9977,N_9915);
or UO_965 (O_965,N_9879,N_9896);
xnor UO_966 (O_966,N_9868,N_9972);
and UO_967 (O_967,N_9951,N_9870);
and UO_968 (O_968,N_9930,N_9827);
or UO_969 (O_969,N_9882,N_9935);
nor UO_970 (O_970,N_9835,N_9878);
or UO_971 (O_971,N_9952,N_9886);
xor UO_972 (O_972,N_9893,N_9969);
nand UO_973 (O_973,N_9817,N_9913);
nor UO_974 (O_974,N_9808,N_9984);
nor UO_975 (O_975,N_9989,N_9933);
and UO_976 (O_976,N_9851,N_9862);
nor UO_977 (O_977,N_9941,N_9847);
nor UO_978 (O_978,N_9868,N_9912);
or UO_979 (O_979,N_9921,N_9955);
nand UO_980 (O_980,N_9974,N_9892);
nor UO_981 (O_981,N_9968,N_9981);
and UO_982 (O_982,N_9965,N_9966);
nand UO_983 (O_983,N_9841,N_9993);
nand UO_984 (O_984,N_9801,N_9970);
or UO_985 (O_985,N_9976,N_9935);
nor UO_986 (O_986,N_9889,N_9808);
and UO_987 (O_987,N_9828,N_9945);
and UO_988 (O_988,N_9903,N_9942);
nor UO_989 (O_989,N_9970,N_9879);
nand UO_990 (O_990,N_9924,N_9994);
or UO_991 (O_991,N_9991,N_9936);
and UO_992 (O_992,N_9835,N_9946);
or UO_993 (O_993,N_9961,N_9893);
nand UO_994 (O_994,N_9981,N_9914);
nand UO_995 (O_995,N_9857,N_9852);
nand UO_996 (O_996,N_9946,N_9923);
or UO_997 (O_997,N_9850,N_9871);
and UO_998 (O_998,N_9910,N_9833);
nand UO_999 (O_999,N_9891,N_9805);
nor UO_1000 (O_1000,N_9868,N_9881);
or UO_1001 (O_1001,N_9901,N_9933);
nand UO_1002 (O_1002,N_9974,N_9875);
or UO_1003 (O_1003,N_9916,N_9996);
nand UO_1004 (O_1004,N_9922,N_9956);
xnor UO_1005 (O_1005,N_9932,N_9842);
or UO_1006 (O_1006,N_9804,N_9985);
nor UO_1007 (O_1007,N_9981,N_9988);
and UO_1008 (O_1008,N_9822,N_9907);
and UO_1009 (O_1009,N_9809,N_9812);
and UO_1010 (O_1010,N_9982,N_9840);
nand UO_1011 (O_1011,N_9850,N_9869);
or UO_1012 (O_1012,N_9886,N_9905);
and UO_1013 (O_1013,N_9894,N_9977);
and UO_1014 (O_1014,N_9819,N_9984);
and UO_1015 (O_1015,N_9854,N_9885);
nor UO_1016 (O_1016,N_9955,N_9910);
nor UO_1017 (O_1017,N_9952,N_9865);
or UO_1018 (O_1018,N_9804,N_9812);
xor UO_1019 (O_1019,N_9977,N_9882);
or UO_1020 (O_1020,N_9855,N_9930);
and UO_1021 (O_1021,N_9870,N_9935);
nand UO_1022 (O_1022,N_9974,N_9948);
nand UO_1023 (O_1023,N_9923,N_9913);
and UO_1024 (O_1024,N_9944,N_9976);
nand UO_1025 (O_1025,N_9833,N_9813);
or UO_1026 (O_1026,N_9807,N_9993);
xnor UO_1027 (O_1027,N_9826,N_9948);
nor UO_1028 (O_1028,N_9880,N_9892);
nor UO_1029 (O_1029,N_9837,N_9827);
nand UO_1030 (O_1030,N_9933,N_9920);
and UO_1031 (O_1031,N_9844,N_9982);
or UO_1032 (O_1032,N_9800,N_9884);
nand UO_1033 (O_1033,N_9948,N_9939);
nor UO_1034 (O_1034,N_9871,N_9898);
or UO_1035 (O_1035,N_9831,N_9931);
nand UO_1036 (O_1036,N_9874,N_9823);
nor UO_1037 (O_1037,N_9976,N_9910);
or UO_1038 (O_1038,N_9852,N_9854);
or UO_1039 (O_1039,N_9991,N_9829);
nor UO_1040 (O_1040,N_9815,N_9807);
nand UO_1041 (O_1041,N_9967,N_9925);
and UO_1042 (O_1042,N_9964,N_9886);
and UO_1043 (O_1043,N_9886,N_9916);
xnor UO_1044 (O_1044,N_9828,N_9811);
xnor UO_1045 (O_1045,N_9956,N_9919);
nor UO_1046 (O_1046,N_9937,N_9846);
and UO_1047 (O_1047,N_9843,N_9873);
or UO_1048 (O_1048,N_9859,N_9931);
nand UO_1049 (O_1049,N_9925,N_9921);
nand UO_1050 (O_1050,N_9989,N_9917);
or UO_1051 (O_1051,N_9889,N_9838);
nor UO_1052 (O_1052,N_9849,N_9906);
and UO_1053 (O_1053,N_9804,N_9994);
nand UO_1054 (O_1054,N_9952,N_9819);
nand UO_1055 (O_1055,N_9974,N_9943);
nor UO_1056 (O_1056,N_9960,N_9986);
nor UO_1057 (O_1057,N_9976,N_9850);
nor UO_1058 (O_1058,N_9819,N_9893);
and UO_1059 (O_1059,N_9946,N_9882);
or UO_1060 (O_1060,N_9842,N_9903);
nand UO_1061 (O_1061,N_9991,N_9957);
nor UO_1062 (O_1062,N_9820,N_9885);
and UO_1063 (O_1063,N_9834,N_9867);
and UO_1064 (O_1064,N_9839,N_9901);
or UO_1065 (O_1065,N_9931,N_9998);
nor UO_1066 (O_1066,N_9909,N_9951);
and UO_1067 (O_1067,N_9825,N_9956);
nand UO_1068 (O_1068,N_9918,N_9967);
nor UO_1069 (O_1069,N_9991,N_9860);
nor UO_1070 (O_1070,N_9857,N_9922);
nand UO_1071 (O_1071,N_9878,N_9803);
nand UO_1072 (O_1072,N_9824,N_9991);
or UO_1073 (O_1073,N_9906,N_9859);
nand UO_1074 (O_1074,N_9942,N_9876);
nor UO_1075 (O_1075,N_9901,N_9830);
xnor UO_1076 (O_1076,N_9937,N_9868);
or UO_1077 (O_1077,N_9962,N_9935);
nor UO_1078 (O_1078,N_9813,N_9950);
or UO_1079 (O_1079,N_9876,N_9845);
nor UO_1080 (O_1080,N_9980,N_9833);
or UO_1081 (O_1081,N_9830,N_9872);
and UO_1082 (O_1082,N_9994,N_9854);
nand UO_1083 (O_1083,N_9948,N_9897);
nor UO_1084 (O_1084,N_9974,N_9862);
nor UO_1085 (O_1085,N_9973,N_9949);
or UO_1086 (O_1086,N_9888,N_9871);
or UO_1087 (O_1087,N_9818,N_9987);
or UO_1088 (O_1088,N_9943,N_9944);
nand UO_1089 (O_1089,N_9921,N_9817);
and UO_1090 (O_1090,N_9825,N_9901);
or UO_1091 (O_1091,N_9939,N_9862);
or UO_1092 (O_1092,N_9959,N_9977);
nor UO_1093 (O_1093,N_9980,N_9957);
or UO_1094 (O_1094,N_9872,N_9864);
nand UO_1095 (O_1095,N_9820,N_9879);
nand UO_1096 (O_1096,N_9902,N_9807);
nand UO_1097 (O_1097,N_9963,N_9964);
or UO_1098 (O_1098,N_9943,N_9814);
nand UO_1099 (O_1099,N_9915,N_9948);
or UO_1100 (O_1100,N_9941,N_9811);
or UO_1101 (O_1101,N_9993,N_9911);
nor UO_1102 (O_1102,N_9943,N_9914);
and UO_1103 (O_1103,N_9818,N_9819);
and UO_1104 (O_1104,N_9873,N_9867);
or UO_1105 (O_1105,N_9887,N_9803);
or UO_1106 (O_1106,N_9979,N_9891);
nor UO_1107 (O_1107,N_9961,N_9824);
and UO_1108 (O_1108,N_9865,N_9975);
nor UO_1109 (O_1109,N_9824,N_9997);
or UO_1110 (O_1110,N_9930,N_9860);
nor UO_1111 (O_1111,N_9811,N_9843);
or UO_1112 (O_1112,N_9941,N_9824);
nor UO_1113 (O_1113,N_9907,N_9923);
xnor UO_1114 (O_1114,N_9852,N_9859);
or UO_1115 (O_1115,N_9906,N_9916);
nor UO_1116 (O_1116,N_9868,N_9949);
nand UO_1117 (O_1117,N_9895,N_9993);
and UO_1118 (O_1118,N_9873,N_9998);
nand UO_1119 (O_1119,N_9846,N_9910);
nor UO_1120 (O_1120,N_9803,N_9902);
nand UO_1121 (O_1121,N_9925,N_9946);
nand UO_1122 (O_1122,N_9906,N_9819);
nor UO_1123 (O_1123,N_9885,N_9953);
nor UO_1124 (O_1124,N_9881,N_9960);
and UO_1125 (O_1125,N_9847,N_9888);
and UO_1126 (O_1126,N_9890,N_9872);
nor UO_1127 (O_1127,N_9924,N_9812);
and UO_1128 (O_1128,N_9840,N_9906);
nand UO_1129 (O_1129,N_9968,N_9837);
and UO_1130 (O_1130,N_9845,N_9889);
and UO_1131 (O_1131,N_9983,N_9907);
nand UO_1132 (O_1132,N_9884,N_9907);
or UO_1133 (O_1133,N_9951,N_9887);
and UO_1134 (O_1134,N_9955,N_9905);
nor UO_1135 (O_1135,N_9983,N_9879);
or UO_1136 (O_1136,N_9986,N_9878);
and UO_1137 (O_1137,N_9999,N_9825);
and UO_1138 (O_1138,N_9903,N_9948);
nand UO_1139 (O_1139,N_9831,N_9871);
or UO_1140 (O_1140,N_9970,N_9960);
and UO_1141 (O_1141,N_9996,N_9906);
or UO_1142 (O_1142,N_9835,N_9808);
and UO_1143 (O_1143,N_9977,N_9844);
nand UO_1144 (O_1144,N_9928,N_9808);
nand UO_1145 (O_1145,N_9943,N_9884);
and UO_1146 (O_1146,N_9901,N_9977);
nor UO_1147 (O_1147,N_9959,N_9911);
nor UO_1148 (O_1148,N_9899,N_9861);
nand UO_1149 (O_1149,N_9822,N_9834);
nor UO_1150 (O_1150,N_9907,N_9961);
and UO_1151 (O_1151,N_9807,N_9867);
nand UO_1152 (O_1152,N_9953,N_9834);
and UO_1153 (O_1153,N_9836,N_9903);
nor UO_1154 (O_1154,N_9803,N_9892);
or UO_1155 (O_1155,N_9946,N_9849);
nand UO_1156 (O_1156,N_9846,N_9879);
nand UO_1157 (O_1157,N_9997,N_9840);
or UO_1158 (O_1158,N_9987,N_9968);
or UO_1159 (O_1159,N_9849,N_9853);
xor UO_1160 (O_1160,N_9990,N_9850);
and UO_1161 (O_1161,N_9874,N_9885);
and UO_1162 (O_1162,N_9809,N_9901);
or UO_1163 (O_1163,N_9974,N_9807);
nand UO_1164 (O_1164,N_9919,N_9900);
or UO_1165 (O_1165,N_9952,N_9870);
nand UO_1166 (O_1166,N_9944,N_9994);
nand UO_1167 (O_1167,N_9974,N_9856);
nor UO_1168 (O_1168,N_9921,N_9971);
and UO_1169 (O_1169,N_9840,N_9864);
xnor UO_1170 (O_1170,N_9975,N_9845);
nand UO_1171 (O_1171,N_9914,N_9992);
xnor UO_1172 (O_1172,N_9928,N_9804);
nand UO_1173 (O_1173,N_9984,N_9965);
nor UO_1174 (O_1174,N_9904,N_9882);
nor UO_1175 (O_1175,N_9895,N_9981);
or UO_1176 (O_1176,N_9827,N_9976);
or UO_1177 (O_1177,N_9957,N_9876);
or UO_1178 (O_1178,N_9896,N_9939);
xnor UO_1179 (O_1179,N_9960,N_9990);
or UO_1180 (O_1180,N_9846,N_9933);
nand UO_1181 (O_1181,N_9867,N_9869);
nor UO_1182 (O_1182,N_9997,N_9998);
or UO_1183 (O_1183,N_9828,N_9935);
or UO_1184 (O_1184,N_9890,N_9994);
nand UO_1185 (O_1185,N_9947,N_9976);
nor UO_1186 (O_1186,N_9815,N_9904);
nor UO_1187 (O_1187,N_9889,N_9839);
or UO_1188 (O_1188,N_9906,N_9990);
nor UO_1189 (O_1189,N_9871,N_9887);
nand UO_1190 (O_1190,N_9807,N_9869);
and UO_1191 (O_1191,N_9836,N_9956);
nand UO_1192 (O_1192,N_9991,N_9923);
xor UO_1193 (O_1193,N_9942,N_9965);
nand UO_1194 (O_1194,N_9842,N_9915);
and UO_1195 (O_1195,N_9965,N_9919);
and UO_1196 (O_1196,N_9886,N_9858);
nand UO_1197 (O_1197,N_9845,N_9997);
nor UO_1198 (O_1198,N_9807,N_9850);
nor UO_1199 (O_1199,N_9948,N_9913);
nor UO_1200 (O_1200,N_9856,N_9987);
nand UO_1201 (O_1201,N_9891,N_9825);
nand UO_1202 (O_1202,N_9946,N_9857);
and UO_1203 (O_1203,N_9978,N_9833);
or UO_1204 (O_1204,N_9899,N_9997);
and UO_1205 (O_1205,N_9863,N_9886);
or UO_1206 (O_1206,N_9805,N_9807);
or UO_1207 (O_1207,N_9991,N_9963);
and UO_1208 (O_1208,N_9949,N_9861);
nor UO_1209 (O_1209,N_9858,N_9855);
nor UO_1210 (O_1210,N_9804,N_9963);
or UO_1211 (O_1211,N_9895,N_9977);
nor UO_1212 (O_1212,N_9965,N_9837);
nor UO_1213 (O_1213,N_9915,N_9942);
and UO_1214 (O_1214,N_9930,N_9868);
and UO_1215 (O_1215,N_9856,N_9803);
nand UO_1216 (O_1216,N_9808,N_9810);
nor UO_1217 (O_1217,N_9930,N_9820);
and UO_1218 (O_1218,N_9908,N_9872);
nand UO_1219 (O_1219,N_9803,N_9801);
and UO_1220 (O_1220,N_9833,N_9869);
nand UO_1221 (O_1221,N_9984,N_9924);
or UO_1222 (O_1222,N_9979,N_9859);
and UO_1223 (O_1223,N_9893,N_9822);
nand UO_1224 (O_1224,N_9903,N_9861);
and UO_1225 (O_1225,N_9984,N_9988);
and UO_1226 (O_1226,N_9872,N_9853);
xor UO_1227 (O_1227,N_9897,N_9896);
nand UO_1228 (O_1228,N_9940,N_9813);
nand UO_1229 (O_1229,N_9843,N_9840);
or UO_1230 (O_1230,N_9992,N_9859);
or UO_1231 (O_1231,N_9986,N_9962);
or UO_1232 (O_1232,N_9835,N_9802);
or UO_1233 (O_1233,N_9829,N_9839);
and UO_1234 (O_1234,N_9954,N_9911);
or UO_1235 (O_1235,N_9963,N_9962);
and UO_1236 (O_1236,N_9951,N_9845);
nor UO_1237 (O_1237,N_9804,N_9909);
nor UO_1238 (O_1238,N_9928,N_9840);
or UO_1239 (O_1239,N_9853,N_9824);
or UO_1240 (O_1240,N_9818,N_9875);
nor UO_1241 (O_1241,N_9841,N_9907);
nor UO_1242 (O_1242,N_9968,N_9984);
or UO_1243 (O_1243,N_9840,N_9813);
or UO_1244 (O_1244,N_9845,N_9871);
nand UO_1245 (O_1245,N_9874,N_9846);
and UO_1246 (O_1246,N_9985,N_9839);
or UO_1247 (O_1247,N_9839,N_9879);
or UO_1248 (O_1248,N_9891,N_9820);
and UO_1249 (O_1249,N_9922,N_9803);
nor UO_1250 (O_1250,N_9933,N_9826);
nand UO_1251 (O_1251,N_9991,N_9989);
nor UO_1252 (O_1252,N_9948,N_9924);
nor UO_1253 (O_1253,N_9983,N_9949);
nand UO_1254 (O_1254,N_9935,N_9904);
and UO_1255 (O_1255,N_9946,N_9962);
nand UO_1256 (O_1256,N_9937,N_9814);
or UO_1257 (O_1257,N_9962,N_9881);
and UO_1258 (O_1258,N_9815,N_9965);
nand UO_1259 (O_1259,N_9886,N_9932);
nor UO_1260 (O_1260,N_9889,N_9876);
or UO_1261 (O_1261,N_9870,N_9989);
or UO_1262 (O_1262,N_9890,N_9928);
nor UO_1263 (O_1263,N_9981,N_9948);
or UO_1264 (O_1264,N_9937,N_9982);
and UO_1265 (O_1265,N_9802,N_9931);
and UO_1266 (O_1266,N_9886,N_9941);
nor UO_1267 (O_1267,N_9862,N_9832);
nor UO_1268 (O_1268,N_9973,N_9915);
nand UO_1269 (O_1269,N_9990,N_9863);
nand UO_1270 (O_1270,N_9903,N_9810);
and UO_1271 (O_1271,N_9888,N_9935);
and UO_1272 (O_1272,N_9851,N_9976);
or UO_1273 (O_1273,N_9944,N_9840);
nor UO_1274 (O_1274,N_9996,N_9809);
xor UO_1275 (O_1275,N_9973,N_9892);
and UO_1276 (O_1276,N_9948,N_9845);
nand UO_1277 (O_1277,N_9897,N_9825);
and UO_1278 (O_1278,N_9937,N_9935);
and UO_1279 (O_1279,N_9856,N_9988);
and UO_1280 (O_1280,N_9812,N_9830);
and UO_1281 (O_1281,N_9854,N_9833);
nand UO_1282 (O_1282,N_9924,N_9825);
nand UO_1283 (O_1283,N_9920,N_9811);
nand UO_1284 (O_1284,N_9983,N_9937);
nand UO_1285 (O_1285,N_9943,N_9953);
and UO_1286 (O_1286,N_9896,N_9828);
or UO_1287 (O_1287,N_9909,N_9837);
or UO_1288 (O_1288,N_9802,N_9971);
xnor UO_1289 (O_1289,N_9832,N_9995);
nor UO_1290 (O_1290,N_9876,N_9938);
nor UO_1291 (O_1291,N_9830,N_9857);
nand UO_1292 (O_1292,N_9826,N_9981);
and UO_1293 (O_1293,N_9959,N_9819);
or UO_1294 (O_1294,N_9939,N_9837);
nand UO_1295 (O_1295,N_9996,N_9998);
and UO_1296 (O_1296,N_9864,N_9971);
and UO_1297 (O_1297,N_9948,N_9837);
nor UO_1298 (O_1298,N_9931,N_9842);
or UO_1299 (O_1299,N_9800,N_9878);
and UO_1300 (O_1300,N_9911,N_9814);
or UO_1301 (O_1301,N_9907,N_9910);
and UO_1302 (O_1302,N_9975,N_9907);
nor UO_1303 (O_1303,N_9991,N_9846);
nor UO_1304 (O_1304,N_9970,N_9933);
or UO_1305 (O_1305,N_9828,N_9962);
or UO_1306 (O_1306,N_9852,N_9824);
and UO_1307 (O_1307,N_9806,N_9899);
and UO_1308 (O_1308,N_9893,N_9931);
or UO_1309 (O_1309,N_9952,N_9983);
or UO_1310 (O_1310,N_9820,N_9873);
and UO_1311 (O_1311,N_9916,N_9841);
and UO_1312 (O_1312,N_9943,N_9999);
nand UO_1313 (O_1313,N_9925,N_9846);
or UO_1314 (O_1314,N_9966,N_9991);
and UO_1315 (O_1315,N_9946,N_9956);
and UO_1316 (O_1316,N_9933,N_9990);
nor UO_1317 (O_1317,N_9804,N_9967);
or UO_1318 (O_1318,N_9901,N_9931);
and UO_1319 (O_1319,N_9994,N_9905);
and UO_1320 (O_1320,N_9963,N_9981);
nand UO_1321 (O_1321,N_9870,N_9904);
or UO_1322 (O_1322,N_9893,N_9908);
and UO_1323 (O_1323,N_9920,N_9804);
and UO_1324 (O_1324,N_9815,N_9941);
nor UO_1325 (O_1325,N_9995,N_9999);
or UO_1326 (O_1326,N_9892,N_9905);
nor UO_1327 (O_1327,N_9963,N_9833);
and UO_1328 (O_1328,N_9829,N_9817);
nor UO_1329 (O_1329,N_9975,N_9826);
nor UO_1330 (O_1330,N_9826,N_9961);
nor UO_1331 (O_1331,N_9895,N_9893);
nor UO_1332 (O_1332,N_9958,N_9820);
nand UO_1333 (O_1333,N_9805,N_9800);
and UO_1334 (O_1334,N_9922,N_9992);
or UO_1335 (O_1335,N_9909,N_9867);
or UO_1336 (O_1336,N_9964,N_9927);
and UO_1337 (O_1337,N_9863,N_9936);
nand UO_1338 (O_1338,N_9916,N_9962);
nand UO_1339 (O_1339,N_9873,N_9916);
nand UO_1340 (O_1340,N_9952,N_9808);
or UO_1341 (O_1341,N_9919,N_9856);
nand UO_1342 (O_1342,N_9837,N_9853);
nand UO_1343 (O_1343,N_9892,N_9990);
or UO_1344 (O_1344,N_9813,N_9959);
or UO_1345 (O_1345,N_9918,N_9992);
or UO_1346 (O_1346,N_9861,N_9806);
and UO_1347 (O_1347,N_9954,N_9818);
and UO_1348 (O_1348,N_9854,N_9991);
nand UO_1349 (O_1349,N_9833,N_9952);
and UO_1350 (O_1350,N_9963,N_9907);
and UO_1351 (O_1351,N_9889,N_9841);
nor UO_1352 (O_1352,N_9968,N_9948);
and UO_1353 (O_1353,N_9875,N_9848);
nand UO_1354 (O_1354,N_9882,N_9963);
nor UO_1355 (O_1355,N_9849,N_9976);
nor UO_1356 (O_1356,N_9937,N_9995);
or UO_1357 (O_1357,N_9988,N_9918);
nor UO_1358 (O_1358,N_9906,N_9948);
nor UO_1359 (O_1359,N_9892,N_9986);
nor UO_1360 (O_1360,N_9935,N_9855);
or UO_1361 (O_1361,N_9931,N_9935);
or UO_1362 (O_1362,N_9801,N_9866);
xor UO_1363 (O_1363,N_9803,N_9931);
nand UO_1364 (O_1364,N_9971,N_9947);
or UO_1365 (O_1365,N_9866,N_9854);
nand UO_1366 (O_1366,N_9894,N_9947);
nand UO_1367 (O_1367,N_9992,N_9804);
or UO_1368 (O_1368,N_9852,N_9957);
or UO_1369 (O_1369,N_9990,N_9948);
nor UO_1370 (O_1370,N_9918,N_9893);
nand UO_1371 (O_1371,N_9911,N_9945);
nor UO_1372 (O_1372,N_9860,N_9980);
and UO_1373 (O_1373,N_9918,N_9884);
and UO_1374 (O_1374,N_9866,N_9990);
nand UO_1375 (O_1375,N_9876,N_9842);
nor UO_1376 (O_1376,N_9953,N_9910);
and UO_1377 (O_1377,N_9928,N_9931);
nor UO_1378 (O_1378,N_9995,N_9866);
nand UO_1379 (O_1379,N_9957,N_9918);
nand UO_1380 (O_1380,N_9808,N_9870);
and UO_1381 (O_1381,N_9810,N_9898);
nand UO_1382 (O_1382,N_9966,N_9967);
or UO_1383 (O_1383,N_9808,N_9974);
nand UO_1384 (O_1384,N_9936,N_9955);
nand UO_1385 (O_1385,N_9934,N_9951);
and UO_1386 (O_1386,N_9897,N_9984);
nand UO_1387 (O_1387,N_9929,N_9997);
and UO_1388 (O_1388,N_9887,N_9939);
and UO_1389 (O_1389,N_9999,N_9846);
nor UO_1390 (O_1390,N_9959,N_9891);
and UO_1391 (O_1391,N_9988,N_9966);
nor UO_1392 (O_1392,N_9904,N_9866);
and UO_1393 (O_1393,N_9815,N_9980);
and UO_1394 (O_1394,N_9864,N_9815);
nor UO_1395 (O_1395,N_9844,N_9966);
and UO_1396 (O_1396,N_9868,N_9953);
nand UO_1397 (O_1397,N_9843,N_9912);
and UO_1398 (O_1398,N_9899,N_9860);
nor UO_1399 (O_1399,N_9973,N_9952);
xor UO_1400 (O_1400,N_9995,N_9980);
nand UO_1401 (O_1401,N_9888,N_9972);
nor UO_1402 (O_1402,N_9867,N_9809);
xor UO_1403 (O_1403,N_9931,N_9940);
or UO_1404 (O_1404,N_9934,N_9845);
nand UO_1405 (O_1405,N_9995,N_9839);
or UO_1406 (O_1406,N_9880,N_9890);
and UO_1407 (O_1407,N_9919,N_9937);
nand UO_1408 (O_1408,N_9883,N_9848);
or UO_1409 (O_1409,N_9805,N_9993);
and UO_1410 (O_1410,N_9904,N_9980);
xor UO_1411 (O_1411,N_9890,N_9963);
nor UO_1412 (O_1412,N_9992,N_9828);
nor UO_1413 (O_1413,N_9863,N_9811);
nand UO_1414 (O_1414,N_9821,N_9905);
nor UO_1415 (O_1415,N_9853,N_9882);
and UO_1416 (O_1416,N_9937,N_9968);
xnor UO_1417 (O_1417,N_9996,N_9951);
nand UO_1418 (O_1418,N_9972,N_9855);
and UO_1419 (O_1419,N_9976,N_9913);
nand UO_1420 (O_1420,N_9945,N_9841);
and UO_1421 (O_1421,N_9949,N_9911);
or UO_1422 (O_1422,N_9911,N_9860);
or UO_1423 (O_1423,N_9874,N_9940);
nor UO_1424 (O_1424,N_9947,N_9935);
or UO_1425 (O_1425,N_9901,N_9844);
and UO_1426 (O_1426,N_9929,N_9925);
or UO_1427 (O_1427,N_9998,N_9932);
or UO_1428 (O_1428,N_9849,N_9848);
and UO_1429 (O_1429,N_9853,N_9998);
nor UO_1430 (O_1430,N_9855,N_9929);
and UO_1431 (O_1431,N_9922,N_9802);
or UO_1432 (O_1432,N_9859,N_9949);
or UO_1433 (O_1433,N_9887,N_9891);
nor UO_1434 (O_1434,N_9988,N_9886);
nor UO_1435 (O_1435,N_9947,N_9942);
nand UO_1436 (O_1436,N_9925,N_9999);
or UO_1437 (O_1437,N_9979,N_9982);
or UO_1438 (O_1438,N_9850,N_9928);
nor UO_1439 (O_1439,N_9813,N_9812);
nand UO_1440 (O_1440,N_9958,N_9973);
nor UO_1441 (O_1441,N_9954,N_9960);
nand UO_1442 (O_1442,N_9900,N_9817);
nor UO_1443 (O_1443,N_9917,N_9897);
nand UO_1444 (O_1444,N_9945,N_9874);
nand UO_1445 (O_1445,N_9959,N_9979);
xor UO_1446 (O_1446,N_9935,N_9973);
nor UO_1447 (O_1447,N_9985,N_9929);
nor UO_1448 (O_1448,N_9824,N_9912);
nand UO_1449 (O_1449,N_9971,N_9900);
nand UO_1450 (O_1450,N_9836,N_9880);
nand UO_1451 (O_1451,N_9814,N_9925);
nor UO_1452 (O_1452,N_9979,N_9991);
nor UO_1453 (O_1453,N_9827,N_9846);
or UO_1454 (O_1454,N_9990,N_9997);
or UO_1455 (O_1455,N_9886,N_9956);
nor UO_1456 (O_1456,N_9881,N_9923);
nor UO_1457 (O_1457,N_9945,N_9854);
or UO_1458 (O_1458,N_9944,N_9975);
and UO_1459 (O_1459,N_9856,N_9847);
nand UO_1460 (O_1460,N_9830,N_9865);
nand UO_1461 (O_1461,N_9875,N_9807);
and UO_1462 (O_1462,N_9905,N_9904);
nand UO_1463 (O_1463,N_9944,N_9958);
nand UO_1464 (O_1464,N_9948,N_9994);
or UO_1465 (O_1465,N_9972,N_9945);
or UO_1466 (O_1466,N_9829,N_9877);
nand UO_1467 (O_1467,N_9873,N_9866);
nand UO_1468 (O_1468,N_9890,N_9990);
or UO_1469 (O_1469,N_9887,N_9807);
nand UO_1470 (O_1470,N_9860,N_9999);
nand UO_1471 (O_1471,N_9915,N_9986);
nand UO_1472 (O_1472,N_9827,N_9896);
and UO_1473 (O_1473,N_9952,N_9842);
nor UO_1474 (O_1474,N_9916,N_9970);
nor UO_1475 (O_1475,N_9848,N_9815);
nand UO_1476 (O_1476,N_9857,N_9862);
or UO_1477 (O_1477,N_9816,N_9817);
or UO_1478 (O_1478,N_9964,N_9902);
or UO_1479 (O_1479,N_9934,N_9839);
or UO_1480 (O_1480,N_9800,N_9987);
nor UO_1481 (O_1481,N_9929,N_9921);
and UO_1482 (O_1482,N_9874,N_9898);
or UO_1483 (O_1483,N_9910,N_9963);
and UO_1484 (O_1484,N_9854,N_9909);
nand UO_1485 (O_1485,N_9854,N_9976);
nand UO_1486 (O_1486,N_9875,N_9860);
or UO_1487 (O_1487,N_9827,N_9851);
nand UO_1488 (O_1488,N_9993,N_9842);
nor UO_1489 (O_1489,N_9802,N_9840);
nor UO_1490 (O_1490,N_9891,N_9900);
nor UO_1491 (O_1491,N_9841,N_9844);
and UO_1492 (O_1492,N_9910,N_9890);
and UO_1493 (O_1493,N_9927,N_9862);
and UO_1494 (O_1494,N_9955,N_9861);
nor UO_1495 (O_1495,N_9889,N_9907);
and UO_1496 (O_1496,N_9859,N_9830);
nor UO_1497 (O_1497,N_9836,N_9855);
or UO_1498 (O_1498,N_9932,N_9991);
and UO_1499 (O_1499,N_9836,N_9928);
endmodule