module basic_1500_15000_2000_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_484,In_850);
or U1 (N_1,In_849,In_483);
xor U2 (N_2,In_187,In_352);
and U3 (N_3,In_122,In_1368);
and U4 (N_4,In_1339,In_926);
or U5 (N_5,In_101,In_92);
or U6 (N_6,In_1055,In_138);
xnor U7 (N_7,In_1344,In_722);
and U8 (N_8,In_1467,In_504);
nor U9 (N_9,In_1353,In_884);
and U10 (N_10,In_1214,In_901);
xor U11 (N_11,In_1453,In_1281);
and U12 (N_12,In_235,In_918);
or U13 (N_13,In_40,In_1020);
nand U14 (N_14,In_252,In_410);
nand U15 (N_15,In_1401,In_4);
xnor U16 (N_16,In_1006,In_370);
xnor U17 (N_17,In_408,In_213);
and U18 (N_18,In_693,In_100);
xor U19 (N_19,In_1324,In_1316);
nand U20 (N_20,In_71,In_1280);
xor U21 (N_21,In_1327,In_378);
or U22 (N_22,In_321,In_393);
xor U23 (N_23,In_908,In_1358);
or U24 (N_24,In_423,In_512);
xor U25 (N_25,In_1473,In_748);
nor U26 (N_26,In_599,In_1011);
xnor U27 (N_27,In_1262,In_342);
nor U28 (N_28,In_1066,In_547);
or U29 (N_29,In_622,In_583);
nand U30 (N_30,In_1212,In_470);
nor U31 (N_31,In_320,In_473);
or U32 (N_32,In_310,In_604);
nand U33 (N_33,In_1135,In_889);
nand U34 (N_34,In_692,In_660);
nor U35 (N_35,In_1164,In_1365);
nand U36 (N_36,In_480,In_155);
nor U37 (N_37,In_1152,In_734);
nor U38 (N_38,In_1375,In_1411);
and U39 (N_39,In_1478,In_1095);
and U40 (N_40,In_109,In_97);
xnor U41 (N_41,In_518,In_39);
or U42 (N_42,In_335,In_980);
nor U43 (N_43,In_615,In_308);
nand U44 (N_44,In_338,In_1201);
xor U45 (N_45,In_834,In_979);
or U46 (N_46,In_825,In_616);
and U47 (N_47,In_649,In_987);
and U48 (N_48,In_330,In_1471);
xnor U49 (N_49,In_1009,In_632);
and U50 (N_50,In_922,In_265);
nor U51 (N_51,In_142,In_1074);
nand U52 (N_52,In_10,In_520);
and U53 (N_53,In_529,In_1179);
and U54 (N_54,In_1499,In_1014);
xnor U55 (N_55,In_497,In_774);
or U56 (N_56,In_1441,In_791);
xnor U57 (N_57,In_1037,In_1308);
nand U58 (N_58,In_356,In_1078);
nand U59 (N_59,In_459,In_822);
nor U60 (N_60,In_301,In_1312);
and U61 (N_61,In_837,In_535);
nand U62 (N_62,In_650,In_680);
and U63 (N_63,In_509,In_984);
nand U64 (N_64,In_695,In_91);
and U65 (N_65,In_726,In_33);
nand U66 (N_66,In_1309,In_1422);
and U67 (N_67,In_221,In_1121);
nor U68 (N_68,In_812,In_211);
and U69 (N_69,In_396,In_415);
nor U70 (N_70,In_847,In_148);
nor U71 (N_71,In_860,In_1050);
or U72 (N_72,In_545,In_823);
or U73 (N_73,In_648,In_465);
nand U74 (N_74,In_781,In_279);
nand U75 (N_75,In_216,In_1379);
nand U76 (N_76,In_565,In_269);
nor U77 (N_77,In_1130,In_1349);
nor U78 (N_78,In_372,In_290);
xor U79 (N_79,In_1053,In_248);
xnor U80 (N_80,In_1176,In_499);
xnor U81 (N_81,In_1091,In_331);
xor U82 (N_82,In_319,In_618);
nand U83 (N_83,In_1028,In_51);
or U84 (N_84,In_1013,In_1223);
or U85 (N_85,In_461,In_741);
nand U86 (N_86,In_762,In_492);
or U87 (N_87,In_694,In_1477);
nand U88 (N_88,In_1167,In_1032);
nor U89 (N_89,In_43,In_52);
and U90 (N_90,In_688,In_427);
xor U91 (N_91,In_619,In_519);
or U92 (N_92,In_28,In_687);
and U93 (N_93,In_214,In_838);
or U94 (N_94,In_1369,In_833);
xor U95 (N_95,In_53,In_747);
nor U96 (N_96,In_627,In_14);
and U97 (N_97,In_1277,In_1105);
and U98 (N_98,In_452,In_260);
and U99 (N_99,In_686,In_585);
xnor U100 (N_100,In_18,In_324);
or U101 (N_101,In_25,In_1094);
and U102 (N_102,In_112,In_366);
and U103 (N_103,In_536,In_1360);
nor U104 (N_104,In_1274,In_963);
nand U105 (N_105,In_1313,In_1483);
xor U106 (N_106,In_1123,In_116);
nor U107 (N_107,In_96,In_1295);
nand U108 (N_108,In_815,In_871);
or U109 (N_109,In_986,In_78);
nor U110 (N_110,In_159,In_771);
and U111 (N_111,In_1355,In_11);
xor U112 (N_112,In_1498,In_1407);
xnor U113 (N_113,In_173,In_232);
and U114 (N_114,In_107,In_608);
xor U115 (N_115,In_1122,In_259);
and U116 (N_116,In_1241,In_906);
nor U117 (N_117,In_668,In_337);
xnor U118 (N_118,In_1062,In_931);
xnor U119 (N_119,In_1323,In_433);
nor U120 (N_120,In_68,In_550);
or U121 (N_121,In_1197,In_441);
and U122 (N_122,In_915,In_1104);
and U123 (N_123,In_806,In_66);
or U124 (N_124,In_885,In_992);
nand U125 (N_125,In_489,In_1373);
xor U126 (N_126,In_1366,In_600);
xnor U127 (N_127,In_939,In_1480);
or U128 (N_128,In_606,In_117);
nand U129 (N_129,In_7,In_88);
and U130 (N_130,In_919,In_1261);
nand U131 (N_131,In_1227,In_391);
xnor U132 (N_132,In_620,In_1188);
and U133 (N_133,In_1269,In_405);
or U134 (N_134,In_1007,In_323);
xnor U135 (N_135,In_1046,In_1452);
and U136 (N_136,In_130,In_970);
and U137 (N_137,In_1131,In_62);
or U138 (N_138,In_165,In_683);
and U139 (N_139,In_1033,In_298);
and U140 (N_140,In_170,In_1082);
and U141 (N_141,In_297,In_1421);
and U142 (N_142,In_1402,In_172);
xor U143 (N_143,In_233,In_240);
nor U144 (N_144,In_1015,In_540);
xor U145 (N_145,In_866,In_1326);
and U146 (N_146,In_700,In_942);
or U147 (N_147,In_1085,In_647);
xor U148 (N_148,In_1204,In_75);
and U149 (N_149,In_720,In_1127);
xor U150 (N_150,In_750,In_736);
nand U151 (N_151,In_1457,In_460);
or U152 (N_152,In_883,In_528);
and U153 (N_153,In_1116,In_176);
nand U154 (N_154,In_578,In_1034);
xnor U155 (N_155,In_8,In_554);
and U156 (N_156,In_1259,In_882);
nor U157 (N_157,In_785,In_887);
nand U158 (N_158,In_322,In_12);
nand U159 (N_159,In_1454,In_803);
nor U160 (N_160,In_892,In_880);
nand U161 (N_161,In_894,In_955);
nor U162 (N_162,In_90,In_1240);
xor U163 (N_163,In_1479,In_238);
or U164 (N_164,In_556,In_810);
nor U165 (N_165,In_663,In_777);
and U166 (N_166,In_1417,In_945);
xnor U167 (N_167,In_1184,In_898);
and U168 (N_168,In_1415,In_386);
nand U169 (N_169,In_203,In_798);
or U170 (N_170,In_1010,In_1089);
nand U171 (N_171,In_194,In_653);
nand U172 (N_172,In_429,In_1388);
xnor U173 (N_173,In_126,In_829);
xor U174 (N_174,In_525,In_1106);
or U175 (N_175,In_488,In_1093);
nand U176 (N_176,In_42,In_478);
nand U177 (N_177,In_1113,In_1146);
xor U178 (N_178,In_689,In_468);
or U179 (N_179,In_1294,In_35);
and U180 (N_180,In_394,In_510);
nand U181 (N_181,In_463,In_998);
xnor U182 (N_182,In_185,In_450);
and U183 (N_183,In_878,In_482);
xor U184 (N_184,In_891,In_250);
or U185 (N_185,In_458,In_1254);
and U186 (N_186,In_1160,In_666);
and U187 (N_187,In_1215,In_1035);
xor U188 (N_188,In_1128,In_362);
and U189 (N_189,In_1056,In_1079);
or U190 (N_190,In_895,In_1148);
and U191 (N_191,In_1057,In_703);
nor U192 (N_192,In_196,In_443);
nand U193 (N_193,In_1427,In_1352);
and U194 (N_194,In_793,In_285);
xnor U195 (N_195,In_169,In_1403);
or U196 (N_196,In_178,In_346);
nand U197 (N_197,In_1111,In_868);
nor U198 (N_198,In_655,In_739);
nor U199 (N_199,In_36,In_743);
nand U200 (N_200,In_485,In_1124);
xnor U201 (N_201,In_186,In_588);
or U202 (N_202,In_1042,In_682);
xnor U203 (N_203,In_641,In_580);
nor U204 (N_204,In_462,In_1137);
nor U205 (N_205,In_1486,In_1172);
and U206 (N_206,In_1354,In_226);
and U207 (N_207,In_139,In_1335);
xnor U208 (N_208,In_153,In_1192);
or U209 (N_209,In_576,In_80);
and U210 (N_210,In_59,In_1383);
and U211 (N_211,In_1086,In_137);
nand U212 (N_212,In_29,In_1359);
or U213 (N_213,In_735,In_1439);
or U214 (N_214,In_674,In_839);
nor U215 (N_215,In_1458,In_1474);
and U216 (N_216,In_1302,In_86);
nor U217 (N_217,In_1145,In_145);
and U218 (N_218,In_664,In_1455);
nand U219 (N_219,In_786,In_755);
xor U220 (N_220,In_1249,In_765);
nor U221 (N_221,In_1251,In_1385);
nor U222 (N_222,In_907,In_1238);
and U223 (N_223,In_418,In_445);
nor U224 (N_224,In_1213,In_768);
nor U225 (N_225,In_698,In_193);
nand U226 (N_226,In_862,In_1409);
and U227 (N_227,In_727,In_1476);
and U228 (N_228,In_1306,In_1291);
nor U229 (N_229,In_48,In_2);
xnor U230 (N_230,In_669,In_95);
or U231 (N_231,In_699,In_773);
or U232 (N_232,In_1067,In_190);
or U233 (N_233,In_354,In_1169);
xnor U234 (N_234,In_1468,In_1399);
or U235 (N_235,In_304,In_220);
xor U236 (N_236,In_560,In_709);
or U237 (N_237,In_223,In_1026);
xor U238 (N_238,In_271,In_150);
xnor U239 (N_239,In_958,In_1073);
xnor U240 (N_240,In_573,In_670);
nand U241 (N_241,In_1225,In_1058);
nor U242 (N_242,In_1207,In_779);
xor U243 (N_243,In_1198,In_523);
and U244 (N_244,In_697,In_610);
and U245 (N_245,In_951,In_347);
xor U246 (N_246,In_1177,In_344);
xor U247 (N_247,In_487,In_439);
xnor U248 (N_248,In_417,In_164);
nor U249 (N_249,In_72,In_1297);
and U250 (N_250,In_561,In_367);
nand U251 (N_251,In_311,In_38);
and U252 (N_252,In_225,In_775);
or U253 (N_253,In_934,In_180);
nand U254 (N_254,In_406,In_1210);
nand U255 (N_255,In_280,In_1278);
or U256 (N_256,In_957,In_287);
and U257 (N_257,In_179,In_132);
or U258 (N_258,In_640,In_1299);
and U259 (N_259,In_329,In_291);
xor U260 (N_260,In_769,In_1462);
nand U261 (N_261,In_0,In_1293);
nand U262 (N_262,In_645,In_913);
or U263 (N_263,In_846,In_1061);
xor U264 (N_264,In_341,In_365);
and U265 (N_265,In_21,In_728);
and U266 (N_266,In_522,In_1098);
nor U267 (N_267,In_542,In_327);
nor U268 (N_268,In_1012,In_517);
nand U269 (N_269,In_1087,In_1248);
nor U270 (N_270,In_1440,In_1024);
nand U271 (N_271,In_911,In_574);
or U272 (N_272,In_134,In_1393);
or U273 (N_273,In_123,In_654);
or U274 (N_274,In_971,In_125);
xor U275 (N_275,In_968,In_594);
nand U276 (N_276,In_359,In_814);
and U277 (N_277,In_587,In_916);
xnor U278 (N_278,In_1022,In_591);
nand U279 (N_279,In_581,In_67);
or U280 (N_280,In_275,In_1194);
xnor U281 (N_281,In_340,In_466);
and U282 (N_282,In_994,In_1395);
nand U283 (N_283,In_455,In_1038);
nor U284 (N_284,In_454,In_1163);
nand U285 (N_285,In_1495,In_1364);
nand U286 (N_286,In_792,In_1219);
or U287 (N_287,In_401,In_1456);
and U288 (N_288,In_776,In_921);
and U289 (N_289,In_1461,In_1216);
and U290 (N_290,In_229,In_1285);
or U291 (N_291,In_613,In_570);
nor U292 (N_292,In_905,In_1118);
nor U293 (N_293,In_1386,In_1224);
xor U294 (N_294,In_1150,In_538);
or U295 (N_295,In_543,In_104);
nor U296 (N_296,In_105,In_904);
and U297 (N_297,In_231,In_261);
xor U298 (N_298,In_184,In_532);
or U299 (N_299,In_79,In_224);
or U300 (N_300,In_972,In_191);
nand U301 (N_301,In_1374,In_1387);
and U302 (N_302,In_662,In_875);
and U303 (N_303,In_1406,In_472);
nand U304 (N_304,In_952,In_19);
nand U305 (N_305,In_371,In_99);
nand U306 (N_306,In_1404,In_770);
nand U307 (N_307,In_551,In_449);
or U308 (N_308,In_413,In_789);
nor U309 (N_309,In_1348,In_893);
or U310 (N_310,In_764,In_339);
and U311 (N_311,In_1263,In_1142);
xor U312 (N_312,In_1185,In_32);
nor U313 (N_313,In_577,In_592);
xor U314 (N_314,In_790,In_27);
or U315 (N_315,In_756,In_1218);
xnor U316 (N_316,In_1191,In_1202);
or U317 (N_317,In_375,In_949);
nor U318 (N_318,In_1236,In_64);
and U319 (N_319,In_421,In_938);
nor U320 (N_320,In_257,In_402);
or U321 (N_321,In_1408,In_869);
nor U322 (N_322,In_1090,In_1187);
and U323 (N_323,In_1005,In_1319);
xor U324 (N_324,In_631,In_127);
or U325 (N_325,In_886,In_1256);
nor U326 (N_326,In_412,In_114);
xnor U327 (N_327,In_1246,In_1125);
and U328 (N_328,In_171,In_133);
nand U329 (N_329,In_1064,In_1242);
xnor U330 (N_330,In_326,In_1036);
nor U331 (N_331,In_1029,In_414);
xor U332 (N_332,In_205,In_296);
xor U333 (N_333,In_827,In_842);
or U334 (N_334,In_435,In_467);
xor U335 (N_335,In_63,In_1377);
and U336 (N_336,In_853,In_1157);
nand U337 (N_337,In_270,In_719);
nand U338 (N_338,In_317,In_245);
xor U339 (N_339,In_247,In_1000);
nor U340 (N_340,In_156,In_293);
xor U341 (N_341,In_552,In_612);
nor U342 (N_342,In_83,In_993);
and U343 (N_343,In_274,In_1484);
and U344 (N_344,In_746,In_383);
and U345 (N_345,In_1490,In_309);
nand U346 (N_346,In_481,In_333);
xor U347 (N_347,In_181,In_1414);
xnor U348 (N_348,In_209,In_227);
and U349 (N_349,In_778,In_865);
nor U350 (N_350,In_586,In_479);
or U351 (N_351,In_258,In_16);
and U352 (N_352,In_672,In_58);
xor U353 (N_353,In_1027,In_124);
and U354 (N_354,In_84,In_1356);
and U355 (N_355,In_557,In_852);
nand U356 (N_356,In_1235,In_438);
and U357 (N_357,In_788,In_400);
nor U358 (N_358,In_836,In_457);
and U359 (N_359,In_246,In_1226);
or U360 (N_360,In_1083,In_749);
xor U361 (N_361,In_696,In_1258);
or U362 (N_362,In_659,In_1051);
or U363 (N_363,In_982,In_1488);
xnor U364 (N_364,In_392,In_665);
xor U365 (N_365,In_1155,In_817);
nand U366 (N_366,In_444,In_841);
nand U367 (N_367,In_589,In_1350);
nand U368 (N_368,In_947,In_685);
nand U369 (N_369,In_1229,In_300);
and U370 (N_370,In_548,In_605);
and U371 (N_371,In_1114,In_419);
or U372 (N_372,In_113,In_70);
nor U373 (N_373,In_859,In_714);
or U374 (N_374,In_767,In_679);
nor U375 (N_375,In_909,In_76);
xor U376 (N_376,In_496,In_1239);
xor U377 (N_377,In_345,In_1096);
nand U378 (N_378,In_526,In_787);
xnor U379 (N_379,In_740,In_1424);
and U380 (N_380,In_1320,In_1052);
and U381 (N_381,In_753,In_147);
nor U382 (N_382,In_1331,In_1068);
or U383 (N_383,In_1182,In_1175);
nor U384 (N_384,In_912,In_434);
or U385 (N_385,In_1442,In_446);
or U386 (N_386,In_1247,In_286);
nor U387 (N_387,In_681,In_1315);
or U388 (N_388,In_353,In_856);
and U389 (N_389,In_30,In_960);
and U390 (N_390,In_724,In_1117);
nor U391 (N_391,In_1288,In_1298);
or U392 (N_392,In_1139,In_844);
nand U393 (N_393,In_282,In_978);
nand U394 (N_394,In_22,In_956);
nand U395 (N_395,In_1436,In_1217);
nor U396 (N_396,In_168,In_349);
nand U397 (N_397,In_369,In_503);
xor U398 (N_398,In_1252,In_456);
and U399 (N_399,In_1199,In_609);
xor U400 (N_400,In_1270,In_1119);
or U401 (N_401,In_314,In_611);
nor U402 (N_402,In_721,In_1180);
or U403 (N_403,In_1231,In_6);
or U404 (N_404,In_26,In_752);
or U405 (N_405,In_218,In_1381);
xnor U406 (N_406,In_334,In_332);
and U407 (N_407,In_407,In_236);
or U408 (N_408,In_494,In_1008);
xor U409 (N_409,In_464,In_962);
and U410 (N_410,In_312,In_1054);
xor U411 (N_411,In_1300,In_189);
nand U412 (N_412,In_596,In_564);
or U413 (N_413,In_857,In_61);
or U414 (N_414,In_539,In_797);
nand U415 (N_415,In_1420,In_1178);
nor U416 (N_416,In_533,In_873);
and U417 (N_417,In_313,In_584);
nor U418 (N_418,In_380,In_13);
xor U419 (N_419,In_783,In_244);
and U420 (N_420,In_1045,In_140);
or U421 (N_421,In_381,In_707);
nor U422 (N_422,In_729,In_1289);
nor U423 (N_423,In_1072,In_328);
nand U424 (N_424,In_212,In_1413);
xor U425 (N_425,In_758,In_306);
nor U426 (N_426,In_389,In_141);
and U427 (N_427,In_1030,In_864);
xor U428 (N_428,In_969,In_1279);
or U429 (N_429,In_500,In_144);
xor U430 (N_430,In_60,In_1459);
and U431 (N_431,In_87,In_263);
nand U432 (N_432,In_1292,In_1431);
nand U433 (N_433,In_192,In_377);
nor U434 (N_434,In_1362,In_1253);
nor U435 (N_435,In_976,In_395);
nor U436 (N_436,In_1425,In_251);
xnor U437 (N_437,In_1444,In_437);
or U438 (N_438,In_56,In_1351);
or U439 (N_439,In_1001,In_974);
or U440 (N_440,In_676,In_476);
nand U441 (N_441,In_1143,In_946);
xnor U442 (N_442,In_1276,In_899);
nor U443 (N_443,In_447,In_1410);
nand U444 (N_444,In_531,In_1023);
and U445 (N_445,In_855,In_1181);
or U446 (N_446,In_1049,In_1392);
or U447 (N_447,In_1041,In_966);
xnor U448 (N_448,In_1196,In_582);
xnor U449 (N_449,In_1264,In_751);
or U450 (N_450,In_237,In_1321);
nor U451 (N_451,In_1200,In_1416);
nor U452 (N_452,In_222,In_1044);
and U453 (N_453,In_808,In_431);
nand U454 (N_454,In_404,In_1437);
xnor U455 (N_455,In_1451,In_23);
or U456 (N_456,In_1443,In_867);
nor U457 (N_457,In_200,In_398);
xnor U458 (N_458,In_731,In_870);
xnor U459 (N_459,In_646,In_1109);
xor U460 (N_460,In_1144,In_843);
nor U461 (N_461,In_409,In_1336);
nand U462 (N_462,In_940,In_416);
and U463 (N_463,In_930,In_1493);
nand U464 (N_464,In_830,In_1165);
nand U465 (N_465,In_343,In_996);
and U466 (N_466,In_630,In_1384);
xnor U467 (N_467,In_691,In_131);
and U468 (N_468,In_1161,In_831);
xnor U469 (N_469,In_325,In_964);
nor U470 (N_470,In_1136,In_119);
nor U471 (N_471,In_1400,In_835);
and U472 (N_472,In_474,In_744);
nor U473 (N_473,In_997,In_448);
nor U474 (N_474,In_1206,In_1162);
or U475 (N_475,In_914,In_712);
and U476 (N_476,In_607,In_819);
xnor U477 (N_477,In_1173,In_491);
xnor U478 (N_478,In_267,In_49);
or U479 (N_479,In_677,In_490);
xor U480 (N_480,In_382,In_903);
or U481 (N_481,In_1266,In_1390);
nor U482 (N_482,In_801,In_925);
nand U483 (N_483,In_1222,In_1154);
nand U484 (N_484,In_527,In_944);
nand U485 (N_485,In_98,In_1043);
xor U486 (N_486,In_110,In_228);
nand U487 (N_487,In_432,In_784);
and U488 (N_488,In_1019,In_1434);
or U489 (N_489,In_888,In_761);
nand U490 (N_490,In_983,In_673);
and U491 (N_491,In_425,In_937);
nand U492 (N_492,In_255,In_1070);
or U493 (N_493,In_780,In_1097);
or U494 (N_494,In_428,In_390);
nor U495 (N_495,In_1310,In_713);
xnor U496 (N_496,In_845,In_1418);
and U497 (N_497,In_420,In_935);
xor U498 (N_498,In_514,In_129);
nor U499 (N_499,In_242,In_81);
nor U500 (N_500,In_288,In_1398);
nor U501 (N_501,In_1017,In_360);
nor U502 (N_502,In_924,In_902);
or U503 (N_503,In_1435,In_502);
xor U504 (N_504,In_1296,In_93);
xor U505 (N_505,In_1485,In_1372);
nor U506 (N_506,In_1092,In_1465);
or U507 (N_507,In_234,In_1286);
or U508 (N_508,In_715,In_292);
xnor U509 (N_509,In_146,In_1449);
and U510 (N_510,In_629,In_368);
nor U511 (N_511,In_1108,In_158);
nor U512 (N_512,In_351,In_498);
nor U513 (N_513,In_628,In_278);
xnor U514 (N_514,In_1397,In_590);
nand U515 (N_515,In_284,In_920);
xor U516 (N_516,In_559,In_961);
nand U517 (N_517,In_188,In_1040);
nor U518 (N_518,In_716,In_281);
nor U519 (N_519,In_851,In_136);
nor U520 (N_520,In_1273,In_1419);
nand U521 (N_521,In_1363,In_708);
nor U522 (N_522,In_262,In_737);
or U523 (N_523,In_273,In_54);
nor U524 (N_524,In_217,In_106);
xnor U525 (N_525,In_1205,In_1343);
or U526 (N_526,In_1307,In_272);
nor U527 (N_527,In_633,In_558);
and U528 (N_528,In_73,In_861);
nand U529 (N_529,In_923,In_1311);
xnor U530 (N_530,In_1080,In_199);
or U531 (N_531,In_268,In_1048);
and U532 (N_532,In_249,In_1134);
or U533 (N_533,In_175,In_403);
nand U534 (N_534,In_544,In_475);
xnor U535 (N_535,In_802,In_374);
nand U536 (N_536,In_567,In_85);
and U537 (N_537,In_546,In_840);
or U538 (N_538,In_959,In_515);
nor U539 (N_539,In_1174,In_239);
or U540 (N_540,In_652,In_1361);
nor U541 (N_541,In_948,In_283);
nand U542 (N_542,In_121,In_1209);
or U543 (N_543,In_848,In_991);
or U544 (N_544,In_1047,In_3);
or U545 (N_545,In_1003,In_1158);
nor U546 (N_546,In_821,In_562);
nand U547 (N_547,In_1491,In_805);
nor U548 (N_548,In_877,In_1065);
xnor U549 (N_549,In_572,In_816);
or U550 (N_550,In_579,In_811);
or U551 (N_551,In_1367,In_1149);
xor U552 (N_552,In_1112,In_1031);
nand U553 (N_553,In_1211,In_1102);
nand U554 (N_554,In_1250,In_197);
and U555 (N_555,In_385,In_442);
nand U556 (N_556,In_34,In_399);
xor U557 (N_557,In_597,In_1018);
nor U558 (N_558,In_651,In_1133);
or U559 (N_559,In_206,In_254);
and U560 (N_560,In_910,In_411);
nand U561 (N_561,In_208,In_1195);
and U562 (N_562,In_1330,In_1171);
or U563 (N_563,In_41,In_757);
and U564 (N_564,In_1159,In_1303);
and U565 (N_565,In_537,In_730);
xnor U566 (N_566,In_230,In_723);
and U567 (N_567,In_1081,In_1345);
or U568 (N_568,In_1141,In_1170);
nand U569 (N_569,In_50,In_215);
nand U570 (N_570,In_174,In_1060);
or U571 (N_571,In_1221,In_1282);
nand U572 (N_572,In_495,In_953);
or U573 (N_573,In_642,In_1470);
nand U574 (N_574,In_1245,In_373);
and U575 (N_575,In_276,In_1075);
nor U576 (N_576,In_702,In_47);
or U577 (N_577,In_1426,In_941);
nand U578 (N_578,In_563,In_1328);
nand U579 (N_579,In_77,In_361);
nor U580 (N_580,In_733,In_1115);
or U581 (N_581,In_995,In_929);
and U582 (N_582,In_1487,In_644);
or U583 (N_583,In_954,In_1234);
nor U584 (N_584,In_1496,In_943);
xor U585 (N_585,In_828,In_363);
nor U586 (N_586,In_754,In_426);
nor U587 (N_587,In_355,In_1304);
nand U588 (N_588,In_508,In_671);
or U589 (N_589,In_1120,In_507);
or U590 (N_590,In_24,In_1338);
nor U591 (N_591,In_936,In_305);
or U592 (N_592,In_896,In_1107);
or U593 (N_593,In_1071,In_384);
nand U594 (N_594,In_1153,In_732);
and U595 (N_595,In_505,In_1232);
nor U596 (N_596,In_690,In_858);
and U597 (N_597,In_760,In_1088);
or U598 (N_598,In_256,In_981);
xnor U599 (N_599,In_182,In_900);
and U600 (N_600,In_928,In_167);
and U601 (N_601,In_711,In_872);
or U602 (N_602,In_1494,In_210);
nand U603 (N_603,In_989,In_854);
xnor U604 (N_604,In_307,In_1464);
or U605 (N_605,In_1275,In_1271);
or U606 (N_606,In_675,In_1140);
nand U607 (N_607,In_289,In_678);
xor U608 (N_608,In_1469,In_617);
nand U609 (N_609,In_1099,In_718);
nand U610 (N_610,In_1243,In_364);
nor U611 (N_611,In_965,In_183);
nand U612 (N_612,In_1039,In_219);
or U613 (N_613,In_453,In_1412);
or U614 (N_614,In_638,In_634);
xor U615 (N_615,In_1257,In_569);
nand U616 (N_616,In_74,In_1272);
and U617 (N_617,In_595,In_568);
nor U618 (N_618,In_807,In_69);
xnor U619 (N_619,In_1016,In_1314);
and U620 (N_620,In_824,In_977);
xor U621 (N_621,In_1084,In_725);
nor U622 (N_622,In_1432,In_661);
xor U623 (N_623,In_511,In_1260);
xnor U624 (N_624,In_9,In_493);
or U625 (N_625,In_809,In_1394);
xnor U626 (N_626,In_530,In_658);
and U627 (N_627,In_160,In_704);
xnor U628 (N_628,In_1147,In_534);
or U629 (N_629,In_31,In_706);
and U630 (N_630,In_684,In_157);
xnor U631 (N_631,In_566,In_643);
or U632 (N_632,In_243,In_818);
xor U633 (N_633,In_348,In_601);
and U634 (N_634,In_1230,In_1126);
nand U635 (N_635,In_1334,In_82);
nor U636 (N_636,In_253,In_988);
nand U637 (N_637,In_1301,In_1472);
nor U638 (N_638,In_623,In_571);
or U639 (N_639,In_151,In_705);
xor U640 (N_640,In_1371,In_1332);
and U641 (N_641,In_1357,In_745);
nand U642 (N_642,In_1168,In_624);
and U643 (N_643,In_1002,In_162);
or U644 (N_644,In_264,In_1492);
nand U645 (N_645,In_710,In_1429);
nand U646 (N_646,In_1132,In_5);
nand U647 (N_647,In_1208,In_1069);
and U648 (N_648,In_152,In_553);
and U649 (N_649,In_874,In_973);
xnor U650 (N_650,In_1103,In_1378);
nor U651 (N_651,In_1156,In_161);
nor U652 (N_652,In_477,In_598);
or U653 (N_653,In_241,In_15);
nand U654 (N_654,In_154,In_820);
or U655 (N_655,In_1244,In_863);
and U656 (N_656,In_1325,In_1475);
and U657 (N_657,In_1284,In_738);
or U658 (N_658,In_128,In_1317);
xnor U659 (N_659,In_800,In_103);
or U660 (N_660,In_379,In_1450);
nor U661 (N_661,In_795,In_1);
nor U662 (N_662,In_166,In_1220);
and U663 (N_663,In_1025,In_813);
xnor U664 (N_664,In_1380,In_516);
or U665 (N_665,In_108,In_1166);
nand U666 (N_666,In_879,In_917);
nand U667 (N_667,In_626,In_198);
nor U668 (N_668,In_299,In_1438);
nand U669 (N_669,In_46,In_471);
or U670 (N_670,In_1382,In_832);
nor U671 (N_671,In_55,In_424);
and U672 (N_672,In_1322,In_1283);
nand U673 (N_673,In_593,In_1423);
and U674 (N_674,In_1481,In_1190);
nand U675 (N_675,In_469,In_20);
nor U676 (N_676,In_118,In_1341);
or U677 (N_677,In_387,In_1228);
nand U678 (N_678,In_195,In_796);
xnor U679 (N_679,In_1193,In_350);
nor U680 (N_680,In_1340,In_303);
xnor U681 (N_681,In_1447,In_1430);
and U682 (N_682,In_1445,In_933);
nor U683 (N_683,In_927,In_506);
or U684 (N_684,In_501,In_1268);
nand U685 (N_685,In_1138,In_763);
xor U686 (N_686,In_1396,In_932);
and U687 (N_687,In_1460,In_436);
nand U688 (N_688,In_336,In_397);
and U689 (N_689,In_985,In_120);
and U690 (N_690,In_430,In_549);
and U691 (N_691,In_451,In_1189);
or U692 (N_692,In_1347,In_897);
nor U693 (N_693,In_1021,In_667);
nand U694 (N_694,In_513,In_524);
nor U695 (N_695,In_1433,In_45);
and U696 (N_696,In_804,In_1100);
nand U697 (N_697,In_163,In_316);
nand U698 (N_698,In_1389,In_575);
nand U699 (N_699,In_1077,In_639);
or U700 (N_700,In_1186,In_17);
nor U701 (N_701,In_149,In_115);
and U702 (N_702,In_1110,In_135);
nand U703 (N_703,In_202,In_1448);
xor U704 (N_704,In_177,In_357);
and U705 (N_705,In_555,In_1342);
and U706 (N_706,In_1482,In_318);
nor U707 (N_707,In_742,In_1267);
or U708 (N_708,In_315,In_657);
xor U709 (N_709,In_1376,In_1183);
xor U710 (N_710,In_89,In_1004);
and U711 (N_711,In_1329,In_201);
and U712 (N_712,In_890,In_1255);
and U713 (N_713,In_1463,In_1287);
nor U714 (N_714,In_999,In_486);
xnor U715 (N_715,In_1489,In_1237);
and U716 (N_716,In_614,In_766);
nor U717 (N_717,In_1101,In_102);
nor U718 (N_718,In_1076,In_826);
and U719 (N_719,In_656,In_1497);
nor U720 (N_720,In_772,In_621);
xnor U721 (N_721,In_1203,In_1305);
nand U722 (N_722,In_1333,In_1318);
and U723 (N_723,In_111,In_1405);
or U724 (N_724,In_295,In_876);
nand U725 (N_725,In_1233,In_1063);
xnor U726 (N_726,In_65,In_950);
nand U727 (N_727,In_1290,In_541);
and U728 (N_728,In_1337,In_388);
nor U729 (N_729,In_625,In_635);
or U730 (N_730,In_1346,In_759);
or U731 (N_731,In_302,In_1428);
xnor U732 (N_732,In_204,In_701);
nor U733 (N_733,In_603,In_1059);
and U734 (N_734,In_637,In_57);
nand U735 (N_735,In_881,In_717);
nor U736 (N_736,In_521,In_294);
nor U737 (N_737,In_1446,In_967);
xor U738 (N_738,In_37,In_975);
or U739 (N_739,In_990,In_782);
and U740 (N_740,In_440,In_207);
xor U741 (N_741,In_1391,In_1370);
or U742 (N_742,In_94,In_358);
nor U743 (N_743,In_1265,In_602);
and U744 (N_744,In_1151,In_799);
nor U745 (N_745,In_794,In_44);
or U746 (N_746,In_422,In_376);
xor U747 (N_747,In_1129,In_143);
nand U748 (N_748,In_266,In_1466);
and U749 (N_749,In_277,In_636);
nor U750 (N_750,In_872,In_1369);
nand U751 (N_751,In_316,In_248);
nor U752 (N_752,In_1305,In_705);
nor U753 (N_753,In_1190,In_1079);
nand U754 (N_754,In_1420,In_181);
nand U755 (N_755,In_689,In_525);
nor U756 (N_756,In_1320,In_550);
xor U757 (N_757,In_1484,In_432);
or U758 (N_758,In_744,In_1459);
nand U759 (N_759,In_1203,In_271);
xor U760 (N_760,In_1184,In_676);
and U761 (N_761,In_1145,In_970);
or U762 (N_762,In_164,In_298);
nor U763 (N_763,In_1300,In_852);
nand U764 (N_764,In_1238,In_1005);
or U765 (N_765,In_1196,In_153);
or U766 (N_766,In_624,In_1193);
nand U767 (N_767,In_1191,In_474);
nand U768 (N_768,In_885,In_779);
nor U769 (N_769,In_373,In_1337);
nand U770 (N_770,In_1014,In_627);
or U771 (N_771,In_1014,In_1154);
or U772 (N_772,In_1465,In_236);
xor U773 (N_773,In_987,In_638);
nor U774 (N_774,In_20,In_280);
xnor U775 (N_775,In_365,In_835);
xor U776 (N_776,In_248,In_546);
xnor U777 (N_777,In_384,In_1198);
xnor U778 (N_778,In_1458,In_1129);
nand U779 (N_779,In_641,In_184);
and U780 (N_780,In_1185,In_37);
and U781 (N_781,In_378,In_1273);
xnor U782 (N_782,In_116,In_20);
xor U783 (N_783,In_1442,In_811);
or U784 (N_784,In_1373,In_592);
nor U785 (N_785,In_804,In_819);
or U786 (N_786,In_659,In_1058);
or U787 (N_787,In_101,In_647);
and U788 (N_788,In_1286,In_1294);
nor U789 (N_789,In_1303,In_653);
or U790 (N_790,In_146,In_264);
xnor U791 (N_791,In_900,In_782);
or U792 (N_792,In_1008,In_972);
xor U793 (N_793,In_348,In_535);
and U794 (N_794,In_300,In_17);
or U795 (N_795,In_1084,In_449);
nand U796 (N_796,In_826,In_990);
nand U797 (N_797,In_202,In_169);
xor U798 (N_798,In_706,In_852);
xnor U799 (N_799,In_1339,In_1150);
xor U800 (N_800,In_266,In_361);
nor U801 (N_801,In_180,In_1118);
or U802 (N_802,In_192,In_1275);
xnor U803 (N_803,In_789,In_349);
and U804 (N_804,In_917,In_1485);
xor U805 (N_805,In_45,In_166);
nor U806 (N_806,In_98,In_363);
and U807 (N_807,In_719,In_11);
nand U808 (N_808,In_664,In_131);
nand U809 (N_809,In_720,In_1365);
or U810 (N_810,In_986,In_1087);
xor U811 (N_811,In_1326,In_651);
or U812 (N_812,In_1408,In_123);
and U813 (N_813,In_523,In_419);
nand U814 (N_814,In_699,In_1124);
or U815 (N_815,In_700,In_28);
and U816 (N_816,In_331,In_478);
nor U817 (N_817,In_648,In_1);
nor U818 (N_818,In_1037,In_318);
and U819 (N_819,In_1447,In_1111);
or U820 (N_820,In_1298,In_165);
xnor U821 (N_821,In_116,In_465);
xor U822 (N_822,In_1041,In_1464);
nor U823 (N_823,In_1144,In_960);
or U824 (N_824,In_813,In_3);
xnor U825 (N_825,In_1156,In_1497);
or U826 (N_826,In_594,In_307);
and U827 (N_827,In_266,In_304);
nor U828 (N_828,In_564,In_1257);
or U829 (N_829,In_745,In_353);
or U830 (N_830,In_1044,In_1404);
or U831 (N_831,In_822,In_735);
nor U832 (N_832,In_246,In_494);
xnor U833 (N_833,In_878,In_1310);
nand U834 (N_834,In_563,In_95);
nor U835 (N_835,In_755,In_1194);
and U836 (N_836,In_1477,In_413);
nand U837 (N_837,In_1012,In_1100);
nor U838 (N_838,In_378,In_657);
or U839 (N_839,In_1376,In_892);
nand U840 (N_840,In_201,In_1213);
and U841 (N_841,In_117,In_315);
and U842 (N_842,In_333,In_360);
nor U843 (N_843,In_1074,In_392);
nor U844 (N_844,In_23,In_1113);
nand U845 (N_845,In_1166,In_1033);
xor U846 (N_846,In_127,In_317);
nand U847 (N_847,In_26,In_1137);
nand U848 (N_848,In_817,In_1136);
nor U849 (N_849,In_249,In_1184);
xnor U850 (N_850,In_140,In_1103);
xnor U851 (N_851,In_401,In_1492);
nand U852 (N_852,In_877,In_354);
and U853 (N_853,In_130,In_456);
nand U854 (N_854,In_1,In_152);
xnor U855 (N_855,In_847,In_202);
xnor U856 (N_856,In_375,In_468);
nor U857 (N_857,In_553,In_177);
nand U858 (N_858,In_953,In_782);
and U859 (N_859,In_1255,In_1048);
nor U860 (N_860,In_786,In_345);
and U861 (N_861,In_1004,In_1075);
nand U862 (N_862,In_1338,In_419);
or U863 (N_863,In_1483,In_1492);
and U864 (N_864,In_540,In_1020);
or U865 (N_865,In_199,In_1353);
xor U866 (N_866,In_1455,In_307);
and U867 (N_867,In_724,In_665);
or U868 (N_868,In_1245,In_173);
nand U869 (N_869,In_213,In_204);
and U870 (N_870,In_694,In_1058);
nand U871 (N_871,In_1226,In_952);
xor U872 (N_872,In_1145,In_673);
or U873 (N_873,In_536,In_564);
nand U874 (N_874,In_902,In_872);
and U875 (N_875,In_260,In_1044);
xor U876 (N_876,In_191,In_403);
nor U877 (N_877,In_1205,In_315);
or U878 (N_878,In_92,In_1202);
or U879 (N_879,In_151,In_1218);
nor U880 (N_880,In_382,In_756);
and U881 (N_881,In_760,In_1273);
nand U882 (N_882,In_971,In_1419);
nand U883 (N_883,In_1027,In_1449);
nor U884 (N_884,In_70,In_163);
and U885 (N_885,In_574,In_1475);
and U886 (N_886,In_103,In_946);
nor U887 (N_887,In_149,In_1245);
nand U888 (N_888,In_1410,In_195);
nand U889 (N_889,In_941,In_690);
xor U890 (N_890,In_839,In_998);
xor U891 (N_891,In_1106,In_1467);
or U892 (N_892,In_678,In_1269);
nand U893 (N_893,In_1471,In_7);
or U894 (N_894,In_1146,In_11);
xnor U895 (N_895,In_207,In_1490);
and U896 (N_896,In_1484,In_1378);
or U897 (N_897,In_735,In_532);
and U898 (N_898,In_1453,In_303);
and U899 (N_899,In_1321,In_1034);
and U900 (N_900,In_35,In_133);
nor U901 (N_901,In_601,In_734);
and U902 (N_902,In_569,In_240);
nand U903 (N_903,In_1308,In_633);
and U904 (N_904,In_384,In_83);
nand U905 (N_905,In_533,In_722);
xor U906 (N_906,In_1120,In_1142);
nor U907 (N_907,In_1072,In_178);
nor U908 (N_908,In_140,In_760);
and U909 (N_909,In_442,In_757);
and U910 (N_910,In_871,In_1170);
xor U911 (N_911,In_624,In_1355);
or U912 (N_912,In_171,In_1468);
or U913 (N_913,In_670,In_533);
nor U914 (N_914,In_1077,In_774);
xnor U915 (N_915,In_477,In_1222);
and U916 (N_916,In_1083,In_382);
nor U917 (N_917,In_1092,In_147);
or U918 (N_918,In_972,In_49);
nor U919 (N_919,In_1490,In_795);
and U920 (N_920,In_873,In_953);
and U921 (N_921,In_442,In_565);
or U922 (N_922,In_155,In_1297);
or U923 (N_923,In_772,In_1357);
nor U924 (N_924,In_416,In_736);
nor U925 (N_925,In_1465,In_306);
and U926 (N_926,In_861,In_56);
xnor U927 (N_927,In_200,In_261);
or U928 (N_928,In_65,In_1155);
nand U929 (N_929,In_743,In_1017);
and U930 (N_930,In_874,In_604);
nor U931 (N_931,In_747,In_388);
xor U932 (N_932,In_317,In_609);
xnor U933 (N_933,In_973,In_1100);
nor U934 (N_934,In_1387,In_1239);
or U935 (N_935,In_440,In_342);
and U936 (N_936,In_786,In_408);
nand U937 (N_937,In_1421,In_595);
and U938 (N_938,In_906,In_1186);
and U939 (N_939,In_702,In_979);
nor U940 (N_940,In_350,In_1077);
and U941 (N_941,In_751,In_802);
xor U942 (N_942,In_1439,In_886);
nor U943 (N_943,In_873,In_643);
and U944 (N_944,In_455,In_757);
xor U945 (N_945,In_838,In_924);
nand U946 (N_946,In_198,In_617);
nand U947 (N_947,In_943,In_1141);
or U948 (N_948,In_1095,In_1403);
and U949 (N_949,In_691,In_10);
and U950 (N_950,In_52,In_121);
xnor U951 (N_951,In_2,In_350);
and U952 (N_952,In_674,In_312);
and U953 (N_953,In_845,In_541);
xor U954 (N_954,In_979,In_216);
or U955 (N_955,In_529,In_182);
nand U956 (N_956,In_1206,In_408);
or U957 (N_957,In_1234,In_1369);
nand U958 (N_958,In_904,In_1033);
nand U959 (N_959,In_246,In_800);
or U960 (N_960,In_933,In_1185);
xnor U961 (N_961,In_1192,In_117);
nor U962 (N_962,In_1325,In_1197);
nor U963 (N_963,In_900,In_661);
nand U964 (N_964,In_920,In_1316);
nand U965 (N_965,In_600,In_1372);
and U966 (N_966,In_1419,In_665);
xor U967 (N_967,In_83,In_1485);
or U968 (N_968,In_936,In_323);
and U969 (N_969,In_771,In_380);
nand U970 (N_970,In_1364,In_70);
nor U971 (N_971,In_223,In_728);
nand U972 (N_972,In_63,In_1284);
nor U973 (N_973,In_420,In_1278);
or U974 (N_974,In_1159,In_1168);
or U975 (N_975,In_1456,In_290);
xnor U976 (N_976,In_641,In_33);
nor U977 (N_977,In_1299,In_1324);
and U978 (N_978,In_186,In_1419);
xnor U979 (N_979,In_1276,In_1183);
and U980 (N_980,In_745,In_181);
nand U981 (N_981,In_684,In_766);
and U982 (N_982,In_906,In_1478);
or U983 (N_983,In_275,In_295);
nand U984 (N_984,In_1369,In_114);
nand U985 (N_985,In_978,In_1302);
and U986 (N_986,In_1435,In_990);
and U987 (N_987,In_17,In_75);
or U988 (N_988,In_765,In_1057);
nand U989 (N_989,In_510,In_97);
and U990 (N_990,In_555,In_1373);
nor U991 (N_991,In_1394,In_707);
nor U992 (N_992,In_381,In_1303);
nor U993 (N_993,In_1221,In_606);
or U994 (N_994,In_537,In_590);
nor U995 (N_995,In_404,In_858);
or U996 (N_996,In_1011,In_424);
nand U997 (N_997,In_886,In_459);
nor U998 (N_998,In_1053,In_581);
xor U999 (N_999,In_983,In_670);
nand U1000 (N_1000,In_945,In_1483);
or U1001 (N_1001,In_399,In_1300);
or U1002 (N_1002,In_1289,In_848);
nand U1003 (N_1003,In_224,In_945);
nor U1004 (N_1004,In_393,In_1342);
nor U1005 (N_1005,In_500,In_1099);
nand U1006 (N_1006,In_1412,In_627);
nor U1007 (N_1007,In_1084,In_1374);
or U1008 (N_1008,In_472,In_263);
nor U1009 (N_1009,In_132,In_1428);
or U1010 (N_1010,In_687,In_1155);
nor U1011 (N_1011,In_686,In_384);
nand U1012 (N_1012,In_125,In_1473);
nand U1013 (N_1013,In_426,In_1141);
nand U1014 (N_1014,In_119,In_129);
xor U1015 (N_1015,In_1137,In_652);
or U1016 (N_1016,In_1034,In_950);
xnor U1017 (N_1017,In_999,In_69);
xnor U1018 (N_1018,In_580,In_1244);
and U1019 (N_1019,In_940,In_1409);
xnor U1020 (N_1020,In_998,In_468);
or U1021 (N_1021,In_1223,In_760);
xnor U1022 (N_1022,In_2,In_492);
or U1023 (N_1023,In_316,In_1070);
or U1024 (N_1024,In_651,In_284);
xnor U1025 (N_1025,In_221,In_1306);
and U1026 (N_1026,In_146,In_159);
or U1027 (N_1027,In_1397,In_31);
nand U1028 (N_1028,In_905,In_161);
nor U1029 (N_1029,In_779,In_1132);
nand U1030 (N_1030,In_1342,In_480);
nor U1031 (N_1031,In_883,In_654);
and U1032 (N_1032,In_626,In_966);
nor U1033 (N_1033,In_220,In_525);
and U1034 (N_1034,In_78,In_866);
nand U1035 (N_1035,In_501,In_11);
or U1036 (N_1036,In_17,In_763);
xnor U1037 (N_1037,In_1399,In_708);
nor U1038 (N_1038,In_1489,In_216);
xnor U1039 (N_1039,In_374,In_652);
and U1040 (N_1040,In_1131,In_952);
or U1041 (N_1041,In_302,In_605);
nor U1042 (N_1042,In_429,In_875);
and U1043 (N_1043,In_1261,In_1491);
nor U1044 (N_1044,In_429,In_496);
and U1045 (N_1045,In_1074,In_28);
nand U1046 (N_1046,In_1052,In_297);
nor U1047 (N_1047,In_619,In_338);
nand U1048 (N_1048,In_415,In_1047);
or U1049 (N_1049,In_1349,In_435);
nor U1050 (N_1050,In_1326,In_654);
nand U1051 (N_1051,In_1446,In_266);
and U1052 (N_1052,In_1315,In_718);
nand U1053 (N_1053,In_782,In_1421);
xnor U1054 (N_1054,In_766,In_1135);
xnor U1055 (N_1055,In_271,In_263);
nor U1056 (N_1056,In_843,In_538);
and U1057 (N_1057,In_995,In_560);
or U1058 (N_1058,In_375,In_929);
xor U1059 (N_1059,In_1012,In_165);
nor U1060 (N_1060,In_1257,In_521);
and U1061 (N_1061,In_620,In_805);
xnor U1062 (N_1062,In_7,In_517);
nand U1063 (N_1063,In_222,In_331);
and U1064 (N_1064,In_401,In_493);
nor U1065 (N_1065,In_865,In_692);
nor U1066 (N_1066,In_1063,In_511);
or U1067 (N_1067,In_298,In_606);
nor U1068 (N_1068,In_1231,In_1386);
nor U1069 (N_1069,In_870,In_184);
nor U1070 (N_1070,In_1214,In_448);
xnor U1071 (N_1071,In_1360,In_565);
xnor U1072 (N_1072,In_301,In_239);
xnor U1073 (N_1073,In_1066,In_1232);
xor U1074 (N_1074,In_10,In_1009);
and U1075 (N_1075,In_1334,In_1296);
or U1076 (N_1076,In_90,In_510);
xnor U1077 (N_1077,In_331,In_793);
or U1078 (N_1078,In_572,In_70);
nand U1079 (N_1079,In_747,In_482);
or U1080 (N_1080,In_588,In_1371);
nand U1081 (N_1081,In_1384,In_474);
nand U1082 (N_1082,In_576,In_150);
or U1083 (N_1083,In_1079,In_257);
and U1084 (N_1084,In_907,In_1396);
or U1085 (N_1085,In_1461,In_384);
or U1086 (N_1086,In_533,In_1473);
or U1087 (N_1087,In_432,In_1114);
and U1088 (N_1088,In_585,In_114);
nor U1089 (N_1089,In_1380,In_187);
and U1090 (N_1090,In_188,In_328);
nand U1091 (N_1091,In_670,In_1159);
and U1092 (N_1092,In_656,In_362);
nand U1093 (N_1093,In_1022,In_881);
or U1094 (N_1094,In_36,In_1359);
or U1095 (N_1095,In_1077,In_706);
nor U1096 (N_1096,In_762,In_719);
and U1097 (N_1097,In_389,In_517);
nand U1098 (N_1098,In_752,In_1373);
and U1099 (N_1099,In_1397,In_810);
xor U1100 (N_1100,In_1428,In_1033);
xnor U1101 (N_1101,In_36,In_569);
nor U1102 (N_1102,In_51,In_1104);
nand U1103 (N_1103,In_976,In_781);
or U1104 (N_1104,In_705,In_1273);
nor U1105 (N_1105,In_1364,In_925);
xor U1106 (N_1106,In_1014,In_1236);
xor U1107 (N_1107,In_364,In_993);
nor U1108 (N_1108,In_211,In_1272);
or U1109 (N_1109,In_676,In_554);
xnor U1110 (N_1110,In_611,In_690);
or U1111 (N_1111,In_825,In_603);
xnor U1112 (N_1112,In_1268,In_256);
nand U1113 (N_1113,In_1108,In_817);
nand U1114 (N_1114,In_531,In_1062);
nand U1115 (N_1115,In_872,In_247);
and U1116 (N_1116,In_12,In_171);
nand U1117 (N_1117,In_135,In_928);
nand U1118 (N_1118,In_195,In_1180);
and U1119 (N_1119,In_460,In_1262);
and U1120 (N_1120,In_1127,In_1126);
nor U1121 (N_1121,In_1343,In_249);
and U1122 (N_1122,In_466,In_645);
nor U1123 (N_1123,In_154,In_1235);
or U1124 (N_1124,In_69,In_121);
nand U1125 (N_1125,In_1150,In_962);
and U1126 (N_1126,In_346,In_47);
or U1127 (N_1127,In_1017,In_1243);
xnor U1128 (N_1128,In_1302,In_1020);
nor U1129 (N_1129,In_1244,In_1446);
xnor U1130 (N_1130,In_613,In_112);
nor U1131 (N_1131,In_604,In_1460);
and U1132 (N_1132,In_206,In_857);
and U1133 (N_1133,In_1345,In_1266);
xnor U1134 (N_1134,In_867,In_840);
or U1135 (N_1135,In_1342,In_509);
or U1136 (N_1136,In_1001,In_696);
or U1137 (N_1137,In_1456,In_1253);
or U1138 (N_1138,In_559,In_426);
xor U1139 (N_1139,In_620,In_1231);
and U1140 (N_1140,In_1299,In_247);
nor U1141 (N_1141,In_408,In_316);
and U1142 (N_1142,In_437,In_184);
nand U1143 (N_1143,In_146,In_305);
and U1144 (N_1144,In_1159,In_184);
nand U1145 (N_1145,In_388,In_879);
nor U1146 (N_1146,In_1064,In_1106);
nand U1147 (N_1147,In_1394,In_512);
nor U1148 (N_1148,In_1412,In_944);
nand U1149 (N_1149,In_464,In_208);
nor U1150 (N_1150,In_127,In_531);
or U1151 (N_1151,In_1457,In_554);
and U1152 (N_1152,In_1234,In_538);
nand U1153 (N_1153,In_1232,In_119);
nand U1154 (N_1154,In_1399,In_14);
xor U1155 (N_1155,In_877,In_349);
and U1156 (N_1156,In_1379,In_1405);
nor U1157 (N_1157,In_296,In_1303);
or U1158 (N_1158,In_549,In_1320);
xnor U1159 (N_1159,In_1456,In_125);
nand U1160 (N_1160,In_36,In_594);
xor U1161 (N_1161,In_545,In_903);
or U1162 (N_1162,In_812,In_627);
and U1163 (N_1163,In_534,In_726);
and U1164 (N_1164,In_1353,In_455);
xnor U1165 (N_1165,In_1139,In_319);
xor U1166 (N_1166,In_1301,In_1086);
and U1167 (N_1167,In_343,In_158);
xor U1168 (N_1168,In_850,In_403);
nand U1169 (N_1169,In_1335,In_707);
xnor U1170 (N_1170,In_432,In_198);
xnor U1171 (N_1171,In_444,In_55);
xor U1172 (N_1172,In_950,In_833);
nor U1173 (N_1173,In_906,In_175);
or U1174 (N_1174,In_1309,In_563);
or U1175 (N_1175,In_1328,In_211);
xnor U1176 (N_1176,In_55,In_682);
or U1177 (N_1177,In_1467,In_526);
or U1178 (N_1178,In_28,In_367);
or U1179 (N_1179,In_725,In_1238);
xor U1180 (N_1180,In_1399,In_247);
and U1181 (N_1181,In_1112,In_680);
nor U1182 (N_1182,In_568,In_1032);
or U1183 (N_1183,In_1212,In_891);
nand U1184 (N_1184,In_417,In_857);
xor U1185 (N_1185,In_656,In_401);
or U1186 (N_1186,In_1241,In_1126);
nor U1187 (N_1187,In_1478,In_1108);
nor U1188 (N_1188,In_396,In_237);
xor U1189 (N_1189,In_1111,In_497);
nand U1190 (N_1190,In_341,In_876);
nor U1191 (N_1191,In_66,In_323);
nor U1192 (N_1192,In_992,In_1409);
nand U1193 (N_1193,In_1181,In_618);
or U1194 (N_1194,In_97,In_17);
nand U1195 (N_1195,In_406,In_942);
and U1196 (N_1196,In_426,In_1090);
nand U1197 (N_1197,In_1340,In_645);
nor U1198 (N_1198,In_17,In_1325);
nor U1199 (N_1199,In_722,In_496);
nor U1200 (N_1200,In_22,In_484);
and U1201 (N_1201,In_318,In_359);
xnor U1202 (N_1202,In_491,In_152);
and U1203 (N_1203,In_332,In_79);
nor U1204 (N_1204,In_399,In_268);
nand U1205 (N_1205,In_615,In_1361);
xor U1206 (N_1206,In_1184,In_1385);
nand U1207 (N_1207,In_32,In_1354);
xor U1208 (N_1208,In_688,In_660);
or U1209 (N_1209,In_364,In_740);
xor U1210 (N_1210,In_164,In_1231);
and U1211 (N_1211,In_931,In_237);
and U1212 (N_1212,In_737,In_452);
xor U1213 (N_1213,In_436,In_486);
nor U1214 (N_1214,In_153,In_465);
or U1215 (N_1215,In_968,In_483);
and U1216 (N_1216,In_109,In_451);
or U1217 (N_1217,In_30,In_807);
or U1218 (N_1218,In_322,In_153);
nand U1219 (N_1219,In_397,In_876);
and U1220 (N_1220,In_1077,In_609);
nand U1221 (N_1221,In_223,In_654);
nor U1222 (N_1222,In_467,In_1323);
nor U1223 (N_1223,In_421,In_1077);
nand U1224 (N_1224,In_155,In_620);
xor U1225 (N_1225,In_1334,In_702);
and U1226 (N_1226,In_597,In_217);
and U1227 (N_1227,In_1232,In_1160);
nor U1228 (N_1228,In_820,In_51);
nor U1229 (N_1229,In_486,In_952);
nand U1230 (N_1230,In_350,In_394);
nand U1231 (N_1231,In_290,In_481);
nand U1232 (N_1232,In_1339,In_389);
nor U1233 (N_1233,In_83,In_441);
nor U1234 (N_1234,In_782,In_1151);
and U1235 (N_1235,In_208,In_1438);
and U1236 (N_1236,In_1224,In_1006);
nor U1237 (N_1237,In_834,In_372);
nor U1238 (N_1238,In_546,In_1180);
nand U1239 (N_1239,In_465,In_850);
or U1240 (N_1240,In_1195,In_1270);
and U1241 (N_1241,In_113,In_57);
nor U1242 (N_1242,In_24,In_867);
nand U1243 (N_1243,In_1428,In_1082);
xnor U1244 (N_1244,In_446,In_857);
and U1245 (N_1245,In_568,In_2);
xor U1246 (N_1246,In_100,In_633);
nor U1247 (N_1247,In_844,In_557);
nand U1248 (N_1248,In_823,In_654);
nand U1249 (N_1249,In_1279,In_208);
or U1250 (N_1250,In_1364,In_1300);
nand U1251 (N_1251,In_956,In_1040);
or U1252 (N_1252,In_820,In_1017);
and U1253 (N_1253,In_829,In_1023);
nor U1254 (N_1254,In_970,In_1137);
xnor U1255 (N_1255,In_1365,In_639);
nand U1256 (N_1256,In_1197,In_142);
and U1257 (N_1257,In_1145,In_14);
xor U1258 (N_1258,In_1048,In_920);
nand U1259 (N_1259,In_1383,In_382);
nand U1260 (N_1260,In_661,In_94);
and U1261 (N_1261,In_487,In_805);
nand U1262 (N_1262,In_550,In_495);
or U1263 (N_1263,In_151,In_172);
nor U1264 (N_1264,In_258,In_870);
and U1265 (N_1265,In_380,In_309);
nor U1266 (N_1266,In_30,In_1154);
xor U1267 (N_1267,In_718,In_646);
xor U1268 (N_1268,In_1226,In_1116);
nand U1269 (N_1269,In_894,In_720);
xor U1270 (N_1270,In_790,In_84);
nor U1271 (N_1271,In_832,In_37);
or U1272 (N_1272,In_688,In_735);
nand U1273 (N_1273,In_981,In_982);
and U1274 (N_1274,In_436,In_531);
or U1275 (N_1275,In_775,In_373);
and U1276 (N_1276,In_1317,In_64);
xor U1277 (N_1277,In_1202,In_711);
and U1278 (N_1278,In_1055,In_132);
or U1279 (N_1279,In_69,In_176);
and U1280 (N_1280,In_773,In_1216);
nand U1281 (N_1281,In_129,In_1475);
or U1282 (N_1282,In_919,In_794);
nor U1283 (N_1283,In_165,In_455);
or U1284 (N_1284,In_709,In_1120);
nor U1285 (N_1285,In_200,In_241);
or U1286 (N_1286,In_853,In_255);
xor U1287 (N_1287,In_791,In_512);
nor U1288 (N_1288,In_1101,In_1263);
or U1289 (N_1289,In_582,In_1194);
nand U1290 (N_1290,In_140,In_795);
and U1291 (N_1291,In_1060,In_730);
xor U1292 (N_1292,In_39,In_906);
nand U1293 (N_1293,In_420,In_314);
or U1294 (N_1294,In_1253,In_1373);
nand U1295 (N_1295,In_766,In_302);
xor U1296 (N_1296,In_80,In_1443);
nand U1297 (N_1297,In_1070,In_250);
xnor U1298 (N_1298,In_821,In_1165);
nor U1299 (N_1299,In_919,In_1241);
and U1300 (N_1300,In_1195,In_293);
nand U1301 (N_1301,In_1347,In_1293);
and U1302 (N_1302,In_971,In_1018);
or U1303 (N_1303,In_228,In_1444);
and U1304 (N_1304,In_1412,In_133);
xor U1305 (N_1305,In_478,In_454);
or U1306 (N_1306,In_972,In_444);
xnor U1307 (N_1307,In_844,In_1101);
nor U1308 (N_1308,In_643,In_416);
nor U1309 (N_1309,In_1108,In_1061);
nor U1310 (N_1310,In_1176,In_4);
nand U1311 (N_1311,In_479,In_25);
and U1312 (N_1312,In_1195,In_549);
nand U1313 (N_1313,In_0,In_193);
nor U1314 (N_1314,In_198,In_543);
xnor U1315 (N_1315,In_1436,In_1003);
or U1316 (N_1316,In_212,In_538);
and U1317 (N_1317,In_434,In_131);
nand U1318 (N_1318,In_349,In_709);
nand U1319 (N_1319,In_36,In_683);
or U1320 (N_1320,In_344,In_225);
nor U1321 (N_1321,In_284,In_1200);
xor U1322 (N_1322,In_142,In_1100);
xnor U1323 (N_1323,In_541,In_938);
nor U1324 (N_1324,In_996,In_994);
xnor U1325 (N_1325,In_645,In_691);
or U1326 (N_1326,In_305,In_518);
nand U1327 (N_1327,In_344,In_332);
nor U1328 (N_1328,In_486,In_1214);
nand U1329 (N_1329,In_770,In_257);
xor U1330 (N_1330,In_764,In_123);
or U1331 (N_1331,In_1471,In_8);
or U1332 (N_1332,In_1272,In_762);
xor U1333 (N_1333,In_172,In_958);
nor U1334 (N_1334,In_1332,In_936);
nand U1335 (N_1335,In_215,In_717);
xnor U1336 (N_1336,In_334,In_972);
nor U1337 (N_1337,In_985,In_263);
nor U1338 (N_1338,In_270,In_682);
xnor U1339 (N_1339,In_273,In_337);
nand U1340 (N_1340,In_646,In_182);
and U1341 (N_1341,In_355,In_857);
nor U1342 (N_1342,In_932,In_893);
nor U1343 (N_1343,In_551,In_1154);
xnor U1344 (N_1344,In_1157,In_485);
or U1345 (N_1345,In_503,In_643);
xor U1346 (N_1346,In_1355,In_1123);
or U1347 (N_1347,In_408,In_1408);
and U1348 (N_1348,In_1237,In_1002);
nor U1349 (N_1349,In_98,In_140);
or U1350 (N_1350,In_661,In_54);
nor U1351 (N_1351,In_1212,In_196);
or U1352 (N_1352,In_1323,In_385);
nor U1353 (N_1353,In_1425,In_1207);
nor U1354 (N_1354,In_1323,In_679);
nor U1355 (N_1355,In_764,In_1121);
nor U1356 (N_1356,In_1364,In_686);
xnor U1357 (N_1357,In_1241,In_901);
nor U1358 (N_1358,In_776,In_541);
or U1359 (N_1359,In_804,In_313);
nor U1360 (N_1360,In_192,In_753);
nand U1361 (N_1361,In_922,In_334);
xor U1362 (N_1362,In_1207,In_986);
and U1363 (N_1363,In_327,In_883);
nand U1364 (N_1364,In_379,In_438);
or U1365 (N_1365,In_524,In_335);
and U1366 (N_1366,In_1260,In_999);
and U1367 (N_1367,In_1294,In_169);
xnor U1368 (N_1368,In_1106,In_1436);
nor U1369 (N_1369,In_1085,In_1480);
xor U1370 (N_1370,In_1005,In_267);
or U1371 (N_1371,In_105,In_960);
xnor U1372 (N_1372,In_537,In_318);
and U1373 (N_1373,In_437,In_748);
nand U1374 (N_1374,In_355,In_1448);
nor U1375 (N_1375,In_303,In_281);
nand U1376 (N_1376,In_669,In_23);
and U1377 (N_1377,In_1087,In_957);
nand U1378 (N_1378,In_371,In_285);
and U1379 (N_1379,In_19,In_1337);
nand U1380 (N_1380,In_351,In_590);
nor U1381 (N_1381,In_283,In_176);
nand U1382 (N_1382,In_375,In_1257);
nor U1383 (N_1383,In_1125,In_732);
and U1384 (N_1384,In_1265,In_291);
nor U1385 (N_1385,In_36,In_1353);
and U1386 (N_1386,In_269,In_488);
nand U1387 (N_1387,In_1293,In_1035);
nand U1388 (N_1388,In_689,In_27);
or U1389 (N_1389,In_865,In_415);
nand U1390 (N_1390,In_1225,In_208);
nand U1391 (N_1391,In_1285,In_1413);
nor U1392 (N_1392,In_1233,In_924);
and U1393 (N_1393,In_8,In_720);
and U1394 (N_1394,In_358,In_6);
xnor U1395 (N_1395,In_896,In_654);
or U1396 (N_1396,In_535,In_1361);
xnor U1397 (N_1397,In_998,In_244);
or U1398 (N_1398,In_542,In_1294);
nand U1399 (N_1399,In_871,In_519);
and U1400 (N_1400,In_1470,In_644);
nor U1401 (N_1401,In_796,In_1187);
or U1402 (N_1402,In_44,In_40);
and U1403 (N_1403,In_345,In_698);
nor U1404 (N_1404,In_500,In_869);
nor U1405 (N_1405,In_938,In_586);
nor U1406 (N_1406,In_678,In_176);
nor U1407 (N_1407,In_851,In_1314);
and U1408 (N_1408,In_1305,In_288);
nor U1409 (N_1409,In_554,In_1258);
nor U1410 (N_1410,In_394,In_1039);
or U1411 (N_1411,In_1233,In_9);
nand U1412 (N_1412,In_1218,In_955);
and U1413 (N_1413,In_1043,In_1212);
xnor U1414 (N_1414,In_798,In_500);
nor U1415 (N_1415,In_830,In_1495);
or U1416 (N_1416,In_982,In_1137);
or U1417 (N_1417,In_391,In_1443);
and U1418 (N_1418,In_1184,In_1353);
nand U1419 (N_1419,In_1391,In_1380);
or U1420 (N_1420,In_1329,In_325);
nor U1421 (N_1421,In_984,In_840);
nand U1422 (N_1422,In_1043,In_1249);
and U1423 (N_1423,In_1014,In_425);
nand U1424 (N_1424,In_639,In_640);
and U1425 (N_1425,In_1049,In_742);
nand U1426 (N_1426,In_36,In_1326);
or U1427 (N_1427,In_1158,In_1100);
or U1428 (N_1428,In_739,In_439);
xnor U1429 (N_1429,In_289,In_208);
and U1430 (N_1430,In_439,In_922);
and U1431 (N_1431,In_461,In_960);
nor U1432 (N_1432,In_1191,In_500);
nand U1433 (N_1433,In_47,In_729);
nor U1434 (N_1434,In_399,In_645);
xnor U1435 (N_1435,In_1377,In_1288);
xor U1436 (N_1436,In_167,In_1473);
and U1437 (N_1437,In_472,In_506);
xnor U1438 (N_1438,In_456,In_580);
nand U1439 (N_1439,In_70,In_1374);
nor U1440 (N_1440,In_669,In_218);
xor U1441 (N_1441,In_1008,In_1364);
nand U1442 (N_1442,In_91,In_184);
nand U1443 (N_1443,In_1498,In_343);
or U1444 (N_1444,In_200,In_755);
or U1445 (N_1445,In_543,In_1029);
and U1446 (N_1446,In_853,In_67);
and U1447 (N_1447,In_1218,In_578);
nor U1448 (N_1448,In_703,In_419);
or U1449 (N_1449,In_1447,In_70);
xor U1450 (N_1450,In_149,In_677);
xor U1451 (N_1451,In_314,In_1220);
nor U1452 (N_1452,In_1230,In_412);
nand U1453 (N_1453,In_423,In_504);
or U1454 (N_1454,In_460,In_397);
nor U1455 (N_1455,In_1157,In_1266);
nand U1456 (N_1456,In_745,In_200);
and U1457 (N_1457,In_432,In_188);
xnor U1458 (N_1458,In_891,In_1408);
nand U1459 (N_1459,In_1273,In_899);
or U1460 (N_1460,In_1352,In_27);
xor U1461 (N_1461,In_603,In_809);
nand U1462 (N_1462,In_13,In_1023);
or U1463 (N_1463,In_90,In_1446);
or U1464 (N_1464,In_439,In_699);
or U1465 (N_1465,In_80,In_1103);
or U1466 (N_1466,In_144,In_6);
nor U1467 (N_1467,In_142,In_1437);
nand U1468 (N_1468,In_840,In_454);
xor U1469 (N_1469,In_1370,In_66);
or U1470 (N_1470,In_1165,In_1044);
nand U1471 (N_1471,In_416,In_198);
nand U1472 (N_1472,In_528,In_664);
nor U1473 (N_1473,In_792,In_1245);
xnor U1474 (N_1474,In_813,In_86);
nor U1475 (N_1475,In_864,In_1225);
or U1476 (N_1476,In_306,In_1295);
nor U1477 (N_1477,In_68,In_813);
xnor U1478 (N_1478,In_209,In_253);
nand U1479 (N_1479,In_1438,In_839);
or U1480 (N_1480,In_273,In_1282);
and U1481 (N_1481,In_1377,In_85);
nor U1482 (N_1482,In_859,In_903);
nand U1483 (N_1483,In_727,In_831);
nor U1484 (N_1484,In_103,In_778);
or U1485 (N_1485,In_1277,In_183);
nor U1486 (N_1486,In_1449,In_193);
nor U1487 (N_1487,In_763,In_1393);
and U1488 (N_1488,In_1466,In_1441);
or U1489 (N_1489,In_524,In_519);
or U1490 (N_1490,In_886,In_64);
and U1491 (N_1491,In_907,In_236);
nand U1492 (N_1492,In_1432,In_733);
or U1493 (N_1493,In_910,In_749);
xnor U1494 (N_1494,In_558,In_830);
nand U1495 (N_1495,In_672,In_806);
nand U1496 (N_1496,In_116,In_646);
xor U1497 (N_1497,In_932,In_692);
or U1498 (N_1498,In_449,In_192);
nand U1499 (N_1499,In_1257,In_850);
and U1500 (N_1500,N_954,N_715);
nand U1501 (N_1501,N_595,N_10);
nor U1502 (N_1502,N_1238,N_94);
or U1503 (N_1503,N_1440,N_368);
xnor U1504 (N_1504,N_525,N_1373);
nand U1505 (N_1505,N_786,N_680);
nor U1506 (N_1506,N_571,N_1076);
xnor U1507 (N_1507,N_1199,N_235);
nor U1508 (N_1508,N_1309,N_1446);
nand U1509 (N_1509,N_1251,N_1073);
nand U1510 (N_1510,N_1051,N_666);
or U1511 (N_1511,N_874,N_805);
nor U1512 (N_1512,N_176,N_32);
and U1513 (N_1513,N_1335,N_1019);
or U1514 (N_1514,N_110,N_672);
nor U1515 (N_1515,N_1496,N_823);
or U1516 (N_1516,N_1148,N_1329);
xor U1517 (N_1517,N_378,N_1307);
and U1518 (N_1518,N_132,N_162);
and U1519 (N_1519,N_733,N_732);
nor U1520 (N_1520,N_1092,N_758);
and U1521 (N_1521,N_409,N_866);
or U1522 (N_1522,N_1404,N_726);
and U1523 (N_1523,N_41,N_926);
or U1524 (N_1524,N_834,N_438);
or U1525 (N_1525,N_1455,N_1003);
nand U1526 (N_1526,N_170,N_352);
or U1527 (N_1527,N_411,N_1105);
nor U1528 (N_1528,N_62,N_948);
xnor U1529 (N_1529,N_1120,N_268);
or U1530 (N_1530,N_965,N_429);
and U1531 (N_1531,N_166,N_727);
nand U1532 (N_1532,N_45,N_709);
nor U1533 (N_1533,N_433,N_300);
nor U1534 (N_1534,N_1012,N_473);
xor U1535 (N_1535,N_314,N_57);
or U1536 (N_1536,N_1421,N_1465);
or U1537 (N_1537,N_104,N_1395);
nor U1538 (N_1538,N_1220,N_1483);
nor U1539 (N_1539,N_426,N_1229);
xnor U1540 (N_1540,N_548,N_938);
nor U1541 (N_1541,N_212,N_1142);
nand U1542 (N_1542,N_1464,N_4);
xnor U1543 (N_1543,N_380,N_679);
nand U1544 (N_1544,N_1201,N_982);
and U1545 (N_1545,N_15,N_25);
nor U1546 (N_1546,N_784,N_161);
or U1547 (N_1547,N_1298,N_576);
or U1548 (N_1548,N_328,N_747);
xnor U1549 (N_1549,N_1346,N_1360);
xor U1550 (N_1550,N_479,N_79);
or U1551 (N_1551,N_1436,N_925);
or U1552 (N_1552,N_740,N_1417);
and U1553 (N_1553,N_1047,N_402);
nor U1554 (N_1554,N_819,N_718);
nor U1555 (N_1555,N_820,N_960);
and U1556 (N_1556,N_95,N_1406);
xor U1557 (N_1557,N_634,N_859);
nor U1558 (N_1558,N_825,N_795);
nand U1559 (N_1559,N_353,N_1333);
nand U1560 (N_1560,N_262,N_682);
and U1561 (N_1561,N_1183,N_287);
or U1562 (N_1562,N_1180,N_573);
nand U1563 (N_1563,N_1467,N_1151);
or U1564 (N_1564,N_721,N_286);
xnor U1565 (N_1565,N_205,N_1103);
and U1566 (N_1566,N_1245,N_1133);
xnor U1567 (N_1567,N_269,N_362);
or U1568 (N_1568,N_1191,N_489);
nand U1569 (N_1569,N_1001,N_937);
xor U1570 (N_1570,N_767,N_1065);
nor U1571 (N_1571,N_702,N_886);
nor U1572 (N_1572,N_1159,N_310);
or U1573 (N_1573,N_887,N_561);
and U1574 (N_1574,N_1418,N_1291);
nand U1575 (N_1575,N_307,N_1196);
xor U1576 (N_1576,N_754,N_431);
xnor U1577 (N_1577,N_652,N_686);
xnor U1578 (N_1578,N_312,N_471);
and U1579 (N_1579,N_822,N_318);
and U1580 (N_1580,N_602,N_885);
and U1581 (N_1581,N_389,N_1193);
and U1582 (N_1582,N_1218,N_164);
nor U1583 (N_1583,N_464,N_399);
xor U1584 (N_1584,N_55,N_997);
and U1585 (N_1585,N_225,N_1062);
nor U1586 (N_1586,N_500,N_29);
nand U1587 (N_1587,N_934,N_1174);
and U1588 (N_1588,N_722,N_1405);
nand U1589 (N_1589,N_1394,N_594);
nand U1590 (N_1590,N_1152,N_1212);
and U1591 (N_1591,N_1344,N_21);
or U1592 (N_1592,N_396,N_23);
or U1593 (N_1593,N_793,N_1027);
and U1594 (N_1594,N_905,N_288);
xnor U1595 (N_1595,N_1275,N_1216);
nand U1596 (N_1596,N_1023,N_851);
or U1597 (N_1597,N_853,N_1126);
xor U1598 (N_1598,N_325,N_870);
nor U1599 (N_1599,N_96,N_821);
xor U1600 (N_1600,N_1499,N_1401);
nand U1601 (N_1601,N_1271,N_1400);
nand U1602 (N_1602,N_791,N_1169);
or U1603 (N_1603,N_449,N_1338);
nand U1604 (N_1604,N_1343,N_803);
nor U1605 (N_1605,N_1241,N_1243);
nand U1606 (N_1606,N_751,N_734);
or U1607 (N_1607,N_350,N_848);
nand U1608 (N_1608,N_875,N_1319);
or U1609 (N_1609,N_285,N_942);
nand U1610 (N_1610,N_37,N_792);
nand U1611 (N_1611,N_1321,N_1119);
or U1612 (N_1612,N_901,N_536);
xor U1613 (N_1613,N_677,N_1215);
nor U1614 (N_1614,N_1137,N_1088);
xnor U1615 (N_1615,N_1443,N_668);
xnor U1616 (N_1616,N_806,N_339);
nor U1617 (N_1617,N_756,N_799);
xnor U1618 (N_1618,N_297,N_1095);
or U1619 (N_1619,N_962,N_98);
and U1620 (N_1620,N_508,N_916);
xnor U1621 (N_1621,N_476,N_1325);
xor U1622 (N_1622,N_1296,N_250);
xor U1623 (N_1623,N_1442,N_1101);
xnor U1624 (N_1624,N_949,N_1301);
or U1625 (N_1625,N_202,N_101);
and U1626 (N_1626,N_485,N_422);
nand U1627 (N_1627,N_158,N_304);
and U1628 (N_1628,N_1022,N_971);
nor U1629 (N_1629,N_1186,N_76);
and U1630 (N_1630,N_116,N_1485);
xor U1631 (N_1631,N_478,N_1078);
nand U1632 (N_1632,N_1433,N_445);
xnor U1633 (N_1633,N_619,N_1129);
xor U1634 (N_1634,N_1136,N_794);
and U1635 (N_1635,N_30,N_1263);
nor U1636 (N_1636,N_17,N_1055);
or U1637 (N_1637,N_529,N_240);
nor U1638 (N_1638,N_1388,N_507);
nor U1639 (N_1639,N_644,N_107);
or U1640 (N_1640,N_412,N_980);
nand U1641 (N_1641,N_332,N_1340);
xnor U1642 (N_1642,N_687,N_1353);
nor U1643 (N_1643,N_995,N_46);
or U1644 (N_1644,N_981,N_230);
nor U1645 (N_1645,N_67,N_81);
xor U1646 (N_1646,N_944,N_1018);
xor U1647 (N_1647,N_1213,N_706);
nor U1648 (N_1648,N_404,N_1125);
nor U1649 (N_1649,N_1057,N_1385);
or U1650 (N_1650,N_991,N_522);
and U1651 (N_1651,N_1265,N_587);
nor U1652 (N_1652,N_204,N_1497);
or U1653 (N_1653,N_1016,N_919);
nand U1654 (N_1654,N_972,N_1314);
nand U1655 (N_1655,N_222,N_810);
and U1656 (N_1656,N_920,N_480);
nand U1657 (N_1657,N_1261,N_653);
xor U1658 (N_1658,N_1117,N_1086);
xnor U1659 (N_1659,N_427,N_1163);
nor U1660 (N_1660,N_181,N_1425);
nand U1661 (N_1661,N_172,N_1020);
or U1662 (N_1662,N_208,N_557);
nand U1663 (N_1663,N_387,N_582);
or U1664 (N_1664,N_517,N_420);
nand U1665 (N_1665,N_1032,N_681);
or U1666 (N_1666,N_664,N_723);
nand U1667 (N_1667,N_1021,N_724);
xor U1668 (N_1668,N_1252,N_231);
nand U1669 (N_1669,N_259,N_103);
or U1670 (N_1670,N_598,N_743);
or U1671 (N_1671,N_629,N_929);
nor U1672 (N_1672,N_367,N_71);
or U1673 (N_1673,N_90,N_1059);
nor U1674 (N_1674,N_1121,N_60);
nor U1675 (N_1675,N_75,N_14);
nor U1676 (N_1676,N_544,N_699);
or U1677 (N_1677,N_601,N_540);
nand U1678 (N_1678,N_535,N_211);
nor U1679 (N_1679,N_125,N_1203);
or U1680 (N_1680,N_39,N_1277);
and U1681 (N_1681,N_376,N_1429);
and U1682 (N_1682,N_63,N_659);
and U1683 (N_1683,N_127,N_813);
nand U1684 (N_1684,N_1376,N_646);
nand U1685 (N_1685,N_752,N_618);
nand U1686 (N_1686,N_1334,N_1083);
xnor U1687 (N_1687,N_379,N_776);
nor U1688 (N_1688,N_1168,N_450);
nand U1689 (N_1689,N_1447,N_192);
or U1690 (N_1690,N_1378,N_191);
xnor U1691 (N_1691,N_467,N_321);
and U1692 (N_1692,N_1323,N_398);
and U1693 (N_1693,N_750,N_405);
nand U1694 (N_1694,N_203,N_1132);
xnor U1695 (N_1695,N_1204,N_145);
and U1696 (N_1696,N_979,N_940);
or U1697 (N_1697,N_624,N_1381);
nor U1698 (N_1698,N_762,N_289);
and U1699 (N_1699,N_130,N_302);
and U1700 (N_1700,N_198,N_555);
or U1701 (N_1701,N_1457,N_329);
and U1702 (N_1702,N_775,N_526);
xor U1703 (N_1703,N_860,N_725);
nor U1704 (N_1704,N_1189,N_115);
or U1705 (N_1705,N_1161,N_1289);
xor U1706 (N_1706,N_1037,N_635);
and U1707 (N_1707,N_1424,N_1317);
and U1708 (N_1708,N_961,N_1074);
and U1709 (N_1709,N_1130,N_357);
nand U1710 (N_1710,N_804,N_134);
nor U1711 (N_1711,N_61,N_407);
nor U1712 (N_1712,N_299,N_957);
xor U1713 (N_1713,N_194,N_745);
or U1714 (N_1714,N_144,N_18);
xor U1715 (N_1715,N_867,N_1480);
and U1716 (N_1716,N_1099,N_1262);
xor U1717 (N_1717,N_1112,N_854);
nand U1718 (N_1718,N_58,N_236);
nand U1719 (N_1719,N_673,N_771);
and U1720 (N_1720,N_915,N_763);
and U1721 (N_1721,N_1063,N_1068);
and U1722 (N_1722,N_88,N_779);
nor U1723 (N_1723,N_1221,N_80);
xnor U1724 (N_1724,N_220,N_1382);
nand U1725 (N_1725,N_178,N_1198);
xor U1726 (N_1726,N_1341,N_1468);
and U1727 (N_1727,N_1244,N_1115);
and U1728 (N_1728,N_520,N_632);
and U1729 (N_1729,N_351,N_364);
nand U1730 (N_1730,N_384,N_1281);
or U1731 (N_1731,N_636,N_898);
nor U1732 (N_1732,N_710,N_34);
nor U1733 (N_1733,N_1432,N_1058);
or U1734 (N_1734,N_229,N_333);
and U1735 (N_1735,N_613,N_372);
or U1736 (N_1736,N_627,N_850);
or U1737 (N_1737,N_703,N_1082);
and U1738 (N_1738,N_1386,N_559);
and U1739 (N_1739,N_1041,N_1165);
xnor U1740 (N_1740,N_373,N_24);
xnor U1741 (N_1741,N_1476,N_827);
xnor U1742 (N_1742,N_360,N_247);
xor U1743 (N_1743,N_242,N_1109);
nand U1744 (N_1744,N_1313,N_1219);
nand U1745 (N_1745,N_1164,N_1392);
xnor U1746 (N_1746,N_579,N_781);
nand U1747 (N_1747,N_1267,N_419);
nor U1748 (N_1748,N_187,N_596);
nand U1749 (N_1749,N_152,N_1403);
and U1750 (N_1750,N_1150,N_669);
nand U1751 (N_1751,N_518,N_369);
nor U1752 (N_1752,N_227,N_955);
xor U1753 (N_1753,N_1113,N_615);
nor U1754 (N_1754,N_1010,N_1416);
or U1755 (N_1755,N_1158,N_691);
and U1756 (N_1756,N_272,N_534);
xnor U1757 (N_1757,N_958,N_1458);
xor U1758 (N_1758,N_1477,N_1498);
and U1759 (N_1759,N_31,N_648);
xnor U1760 (N_1760,N_698,N_493);
nand U1761 (N_1761,N_155,N_1205);
or U1762 (N_1762,N_502,N_1106);
nor U1763 (N_1763,N_446,N_707);
nor U1764 (N_1764,N_719,N_1089);
or U1765 (N_1765,N_978,N_151);
nand U1766 (N_1766,N_501,N_833);
nand U1767 (N_1767,N_1147,N_1206);
xnor U1768 (N_1768,N_1144,N_1049);
or U1769 (N_1769,N_244,N_282);
xor U1770 (N_1770,N_1236,N_701);
xnor U1771 (N_1771,N_1084,N_1131);
nor U1772 (N_1772,N_670,N_692);
xnor U1773 (N_1773,N_946,N_296);
nor U1774 (N_1774,N_896,N_1166);
xnor U1775 (N_1775,N_1294,N_1437);
or U1776 (N_1776,N_184,N_169);
xor U1777 (N_1777,N_337,N_1258);
and U1778 (N_1778,N_910,N_527);
nor U1779 (N_1779,N_1288,N_397);
nand U1780 (N_1780,N_1038,N_403);
and U1781 (N_1781,N_108,N_1177);
or U1782 (N_1782,N_156,N_633);
or U1783 (N_1783,N_1187,N_190);
xor U1784 (N_1784,N_207,N_894);
xnor U1785 (N_1785,N_684,N_1160);
nand U1786 (N_1786,N_42,N_1028);
xor U1787 (N_1787,N_291,N_1128);
and U1788 (N_1788,N_1349,N_223);
nor U1789 (N_1789,N_1487,N_728);
xnor U1790 (N_1790,N_319,N_1450);
nand U1791 (N_1791,N_456,N_661);
and U1792 (N_1792,N_897,N_341);
and U1793 (N_1793,N_790,N_298);
nor U1794 (N_1794,N_159,N_964);
nor U1795 (N_1795,N_909,N_474);
or U1796 (N_1796,N_1175,N_461);
and U1797 (N_1797,N_443,N_678);
nor U1798 (N_1798,N_117,N_200);
or U1799 (N_1799,N_56,N_1428);
nand U1800 (N_1800,N_53,N_969);
or U1801 (N_1801,N_68,N_1045);
nor U1802 (N_1802,N_234,N_843);
or U1803 (N_1803,N_986,N_1365);
nor U1804 (N_1804,N_395,N_487);
nand U1805 (N_1805,N_1034,N_188);
and U1806 (N_1806,N_924,N_650);
xor U1807 (N_1807,N_1359,N_782);
or U1808 (N_1808,N_270,N_616);
nand U1809 (N_1809,N_283,N_584);
xor U1810 (N_1810,N_1033,N_1490);
and U1811 (N_1811,N_454,N_1188);
xor U1812 (N_1812,N_872,N_862);
or U1813 (N_1813,N_1276,N_1396);
nor U1814 (N_1814,N_1293,N_696);
nand U1815 (N_1815,N_486,N_1282);
or U1816 (N_1816,N_1134,N_2);
xor U1817 (N_1817,N_953,N_1138);
nand U1818 (N_1818,N_654,N_676);
xnor U1819 (N_1819,N_951,N_1473);
or U1820 (N_1820,N_306,N_316);
and U1821 (N_1821,N_83,N_1297);
xor U1822 (N_1822,N_324,N_550);
nand U1823 (N_1823,N_257,N_1176);
nor U1824 (N_1824,N_1014,N_1155);
nor U1825 (N_1825,N_606,N_1085);
nand U1826 (N_1826,N_835,N_1044);
and U1827 (N_1827,N_1235,N_1029);
nor U1828 (N_1828,N_943,N_439);
nand U1829 (N_1829,N_1026,N_97);
nor U1830 (N_1830,N_221,N_999);
or U1831 (N_1831,N_828,N_254);
and U1832 (N_1832,N_136,N_1207);
nand U1833 (N_1833,N_326,N_59);
and U1834 (N_1834,N_386,N_530);
and U1835 (N_1835,N_277,N_469);
xnor U1836 (N_1836,N_1361,N_906);
nor U1837 (N_1837,N_1482,N_675);
xor U1838 (N_1838,N_1460,N_1170);
nand U1839 (N_1839,N_539,N_320);
nor U1840 (N_1840,N_1355,N_742);
nor U1841 (N_1841,N_801,N_693);
xnor U1842 (N_1842,N_506,N_617);
xnor U1843 (N_1843,N_344,N_1157);
nand U1844 (N_1844,N_1124,N_1491);
xor U1845 (N_1845,N_1459,N_1452);
nand U1846 (N_1846,N_789,N_845);
or U1847 (N_1847,N_513,N_1441);
nor U1848 (N_1848,N_74,N_84);
nand U1849 (N_1849,N_142,N_1279);
nor U1850 (N_1850,N_150,N_609);
or U1851 (N_1851,N_945,N_246);
xor U1852 (N_1852,N_143,N_839);
and U1853 (N_1853,N_239,N_768);
nand U1854 (N_1854,N_163,N_1331);
nor U1855 (N_1855,N_430,N_1066);
or U1856 (N_1856,N_630,N_358);
xnor U1857 (N_1857,N_963,N_542);
xnor U1858 (N_1858,N_276,N_1179);
nor U1859 (N_1859,N_1102,N_1488);
nand U1860 (N_1860,N_537,N_499);
or U1861 (N_1861,N_241,N_363);
nor U1862 (N_1862,N_849,N_1209);
nand U1863 (N_1863,N_608,N_605);
or U1864 (N_1864,N_435,N_504);
nor U1865 (N_1865,N_1332,N_588);
and U1866 (N_1866,N_173,N_356);
nor U1867 (N_1867,N_883,N_578);
xor U1868 (N_1868,N_505,N_759);
xnor U1869 (N_1869,N_830,N_40);
and U1870 (N_1870,N_228,N_800);
xnor U1871 (N_1871,N_1339,N_711);
or U1872 (N_1872,N_1380,N_917);
and U1873 (N_1873,N_1486,N_993);
and U1874 (N_1874,N_1495,N_545);
nor U1875 (N_1875,N_189,N_102);
nor U1876 (N_1876,N_788,N_620);
nand U1877 (N_1877,N_248,N_638);
and U1878 (N_1878,N_685,N_884);
and U1879 (N_1879,N_1046,N_423);
nor U1880 (N_1880,N_893,N_284);
or U1881 (N_1881,N_253,N_416);
nand U1882 (N_1882,N_1303,N_575);
or U1883 (N_1883,N_290,N_921);
nand U1884 (N_1884,N_984,N_1197);
nand U1885 (N_1885,N_512,N_160);
nor U1886 (N_1886,N_267,N_739);
and U1887 (N_1887,N_1466,N_1270);
or U1888 (N_1888,N_1383,N_876);
and U1889 (N_1889,N_1087,N_936);
nand U1890 (N_1890,N_1153,N_106);
nand U1891 (N_1891,N_498,N_1342);
nand U1892 (N_1892,N_201,N_1108);
nand U1893 (N_1893,N_77,N_553);
and U1894 (N_1894,N_93,N_1036);
xnor U1895 (N_1895,N_1387,N_1211);
and U1896 (N_1896,N_1048,N_996);
nor U1897 (N_1897,N_123,N_581);
and U1898 (N_1898,N_1013,N_861);
nand U1899 (N_1899,N_863,N_837);
or U1900 (N_1900,N_315,N_785);
nand U1901 (N_1901,N_1031,N_1402);
or U1902 (N_1902,N_271,N_1348);
nand U1903 (N_1903,N_484,N_858);
nand U1904 (N_1904,N_251,N_64);
and U1905 (N_1905,N_524,N_349);
or U1906 (N_1906,N_1242,N_20);
nor U1907 (N_1907,N_260,N_778);
and U1908 (N_1908,N_900,N_1493);
and U1909 (N_1909,N_931,N_105);
nor U1910 (N_1910,N_857,N_1060);
or U1911 (N_1911,N_1043,N_838);
nand U1912 (N_1912,N_483,N_1273);
or U1913 (N_1913,N_361,N_54);
or U1914 (N_1914,N_1410,N_448);
and U1915 (N_1915,N_1178,N_432);
nor U1916 (N_1916,N_1326,N_35);
nor U1917 (N_1917,N_1352,N_731);
and U1918 (N_1918,N_757,N_983);
nor U1919 (N_1919,N_22,N_1463);
and U1920 (N_1920,N_528,N_1079);
nor U1921 (N_1921,N_7,N_532);
and U1922 (N_1922,N_645,N_436);
or U1923 (N_1923,N_153,N_475);
nand U1924 (N_1924,N_737,N_551);
nand U1925 (N_1925,N_994,N_565);
nand U1926 (N_1926,N_603,N_1239);
nand U1927 (N_1927,N_631,N_1266);
nor U1928 (N_1928,N_275,N_903);
xor U1929 (N_1929,N_1357,N_600);
xnor U1930 (N_1930,N_519,N_92);
nand U1931 (N_1931,N_462,N_174);
or U1932 (N_1932,N_481,N_628);
and U1933 (N_1933,N_147,N_196);
nand U1934 (N_1934,N_1324,N_496);
and U1935 (N_1935,N_1372,N_466);
nand U1936 (N_1936,N_708,N_878);
xor U1937 (N_1937,N_868,N_345);
nor U1938 (N_1938,N_817,N_78);
xor U1939 (N_1939,N_1162,N_274);
or U1940 (N_1940,N_649,N_563);
xnor U1941 (N_1941,N_658,N_1312);
and U1942 (N_1942,N_428,N_1091);
nor U1943 (N_1943,N_549,N_317);
nand U1944 (N_1944,N_932,N_245);
xnor U1945 (N_1945,N_1064,N_261);
xnor U1946 (N_1946,N_348,N_118);
nor U1947 (N_1947,N_424,N_273);
nor U1948 (N_1948,N_738,N_640);
xnor U1949 (N_1949,N_301,N_1390);
and U1950 (N_1950,N_65,N_281);
or U1951 (N_1951,N_748,N_109);
nor U1952 (N_1952,N_558,N_780);
nor U1953 (N_1953,N_1408,N_85);
nand U1954 (N_1954,N_491,N_988);
xor U1955 (N_1955,N_11,N_580);
nor U1956 (N_1956,N_1259,N_135);
nor U1957 (N_1957,N_1345,N_1407);
nor U1958 (N_1958,N_538,N_798);
or U1959 (N_1959,N_195,N_1430);
nor U1960 (N_1960,N_355,N_647);
or U1961 (N_1961,N_381,N_783);
and U1962 (N_1962,N_1143,N_712);
and U1963 (N_1963,N_87,N_354);
and U1964 (N_1964,N_1264,N_1456);
and U1965 (N_1965,N_1489,N_28);
xnor U1966 (N_1966,N_593,N_1061);
or U1967 (N_1967,N_124,N_1272);
or U1968 (N_1968,N_973,N_735);
nand U1969 (N_1969,N_468,N_1071);
nand U1970 (N_1970,N_1096,N_393);
and U1971 (N_1971,N_970,N_569);
nor U1972 (N_1972,N_546,N_847);
nand U1973 (N_1973,N_1328,N_607);
and U1974 (N_1974,N_1284,N_912);
and U1975 (N_1975,N_1200,N_490);
and U1976 (N_1976,N_186,N_82);
nand U1977 (N_1977,N_704,N_1370);
nand U1978 (N_1978,N_69,N_451);
xnor U1979 (N_1979,N_586,N_1094);
nand U1980 (N_1980,N_1194,N_610);
nor U1981 (N_1981,N_612,N_831);
or U1982 (N_1982,N_642,N_914);
or U1983 (N_1983,N_148,N_871);
nand U1984 (N_1984,N_122,N_975);
xor U1985 (N_1985,N_382,N_72);
nand U1986 (N_1986,N_1107,N_1139);
nand U1987 (N_1987,N_1004,N_902);
and U1988 (N_1988,N_1367,N_330);
nand U1989 (N_1989,N_1208,N_418);
and U1990 (N_1990,N_224,N_882);
xor U1991 (N_1991,N_639,N_1420);
and U1992 (N_1992,N_140,N_824);
nand U1993 (N_1993,N_237,N_918);
and U1994 (N_1994,N_1039,N_1434);
and U1995 (N_1995,N_213,N_891);
xnor U1996 (N_1996,N_1474,N_665);
nor U1997 (N_1997,N_0,N_892);
nor U1998 (N_1998,N_562,N_1173);
nor U1999 (N_1999,N_465,N_1248);
or U2000 (N_2000,N_1093,N_209);
nand U2001 (N_2001,N_336,N_1391);
and U2002 (N_2002,N_1250,N_674);
and U2003 (N_2003,N_1308,N_566);
and U2004 (N_2004,N_889,N_89);
nor U2005 (N_2005,N_1005,N_1070);
nor U2006 (N_2006,N_663,N_797);
or U2007 (N_2007,N_375,N_764);
nor U2008 (N_2008,N_749,N_495);
xnor U2009 (N_2009,N_452,N_911);
or U2010 (N_2010,N_770,N_966);
nand U2011 (N_2011,N_714,N_463);
and U2012 (N_2012,N_165,N_70);
or U2013 (N_2013,N_86,N_1454);
or U2014 (N_2014,N_447,N_133);
nand U2015 (N_2015,N_662,N_690);
nand U2016 (N_2016,N_370,N_1356);
nor U2017 (N_2017,N_694,N_410);
xnor U2018 (N_2018,N_131,N_1366);
or U2019 (N_2019,N_516,N_1472);
nand U2020 (N_2020,N_390,N_414);
xnor U2021 (N_2021,N_255,N_1268);
or U2022 (N_2022,N_952,N_48);
xor U2023 (N_2023,N_1327,N_590);
xnor U2024 (N_2024,N_904,N_459);
and U2025 (N_2025,N_985,N_890);
nand U2026 (N_2026,N_841,N_52);
xnor U2027 (N_2027,N_689,N_1000);
and U2028 (N_2028,N_1,N_881);
nor U2029 (N_2029,N_1190,N_217);
xor U2030 (N_2030,N_968,N_388);
nor U2031 (N_2031,N_1419,N_263);
or U2032 (N_2032,N_1067,N_455);
or U2033 (N_2033,N_1254,N_417);
nor U2034 (N_2034,N_472,N_621);
and U2035 (N_2035,N_206,N_1006);
and U2036 (N_2036,N_1439,N_1411);
or U2037 (N_2037,N_856,N_1114);
nor U2038 (N_2038,N_826,N_990);
nor U2039 (N_2039,N_1210,N_1393);
nor U2040 (N_2040,N_585,N_956);
and U2041 (N_2041,N_1494,N_560);
and U2042 (N_2042,N_171,N_1127);
nor U2043 (N_2043,N_342,N_1426);
nor U2044 (N_2044,N_729,N_457);
nor U2045 (N_2045,N_1192,N_832);
nand U2046 (N_2046,N_1336,N_120);
xor U2047 (N_2047,N_1280,N_50);
or U2048 (N_2048,N_895,N_1224);
nand U2049 (N_2049,N_308,N_26);
xnor U2050 (N_2050,N_347,N_292);
or U2051 (N_2051,N_1141,N_444);
nor U2052 (N_2052,N_1100,N_335);
nand U2053 (N_2053,N_716,N_753);
and U2054 (N_2054,N_1330,N_1304);
and U2055 (N_2055,N_1135,N_309);
nor U2056 (N_2056,N_210,N_182);
or U2057 (N_2057,N_967,N_1350);
and U2058 (N_2058,N_611,N_216);
and U2059 (N_2059,N_625,N_1462);
nor U2060 (N_2060,N_1414,N_9);
or U2061 (N_2061,N_774,N_1156);
xnor U2062 (N_2062,N_667,N_547);
and U2063 (N_2063,N_927,N_1471);
nand U2064 (N_2064,N_1409,N_947);
nor U2065 (N_2065,N_877,N_36);
and U2066 (N_2066,N_440,N_266);
xnor U2067 (N_2067,N_842,N_523);
xnor U2068 (N_2068,N_197,N_1253);
nor U2069 (N_2069,N_1484,N_836);
nor U2070 (N_2070,N_989,N_531);
or U2071 (N_2071,N_1322,N_922);
nor U2072 (N_2072,N_1318,N_279);
and U2073 (N_2073,N_1377,N_1413);
and U2074 (N_2074,N_657,N_574);
xor U2075 (N_2075,N_695,N_766);
or U2076 (N_2076,N_807,N_713);
or U2077 (N_2077,N_641,N_1315);
nor U2078 (N_2078,N_509,N_1053);
or U2079 (N_2079,N_626,N_814);
or U2080 (N_2080,N_334,N_1283);
or U2081 (N_2081,N_214,N_265);
and U2082 (N_2082,N_855,N_413);
nand U2083 (N_2083,N_408,N_503);
or U2084 (N_2084,N_415,N_1451);
nand U2085 (N_2085,N_1122,N_554);
nor U2086 (N_2086,N_744,N_383);
and U2087 (N_2087,N_1470,N_137);
xor U2088 (N_2088,N_1384,N_572);
and U2089 (N_2089,N_773,N_720);
xnor U2090 (N_2090,N_1140,N_99);
or U2091 (N_2091,N_177,N_697);
xnor U2092 (N_2092,N_346,N_185);
xnor U2093 (N_2093,N_1310,N_746);
nor U2094 (N_2094,N_243,N_13);
nand U2095 (N_2095,N_1149,N_19);
xnor U2096 (N_2096,N_180,N_138);
nor U2097 (N_2097,N_232,N_1260);
or U2098 (N_2098,N_33,N_1347);
xnor U2099 (N_2099,N_1040,N_1146);
nor U2100 (N_2100,N_614,N_913);
nor U2101 (N_2101,N_1364,N_38);
and U2102 (N_2102,N_1375,N_401);
nand U2103 (N_2103,N_908,N_846);
or U2104 (N_2104,N_73,N_1015);
or U2105 (N_2105,N_808,N_987);
nand U2106 (N_2106,N_1227,N_816);
xnor U2107 (N_2107,N_146,N_1290);
nand U2108 (N_2108,N_741,N_1222);
and U2109 (N_2109,N_1478,N_655);
or U2110 (N_2110,N_1154,N_930);
or U2111 (N_2111,N_323,N_1228);
and U2112 (N_2112,N_27,N_322);
xnor U2113 (N_2113,N_777,N_1240);
nor U2114 (N_2114,N_923,N_340);
nor U2115 (N_2115,N_888,N_844);
nand U2116 (N_2116,N_1302,N_1232);
nand U2117 (N_2117,N_5,N_91);
and U2118 (N_2118,N_1247,N_1306);
nor U2119 (N_2119,N_492,N_556);
xor U2120 (N_2120,N_939,N_141);
nand U2121 (N_2121,N_1246,N_514);
or U2122 (N_2122,N_1363,N_765);
or U2123 (N_2123,N_852,N_1295);
nor U2124 (N_2124,N_215,N_796);
xor U2125 (N_2125,N_1123,N_343);
xor U2126 (N_2126,N_772,N_998);
nand U2127 (N_2127,N_992,N_219);
nor U2128 (N_2128,N_1475,N_1011);
nor U2129 (N_2129,N_1469,N_238);
nor U2130 (N_2130,N_112,N_128);
or U2131 (N_2131,N_755,N_564);
or U2132 (N_2132,N_1492,N_1278);
nor U2133 (N_2133,N_392,N_1098);
nand U2134 (N_2134,N_51,N_366);
nor U2135 (N_2135,N_1069,N_252);
or U2136 (N_2136,N_295,N_1195);
and U2137 (N_2137,N_359,N_406);
xor U2138 (N_2138,N_1300,N_331);
and U2139 (N_2139,N_1050,N_1412);
or U2140 (N_2140,N_1368,N_1080);
or U2141 (N_2141,N_425,N_1292);
nand U2142 (N_2142,N_371,N_976);
and U2143 (N_2143,N_470,N_1427);
xnor U2144 (N_2144,N_1299,N_1171);
xor U2145 (N_2145,N_1369,N_1008);
xor U2146 (N_2146,N_494,N_338);
and U2147 (N_2147,N_865,N_477);
and U2148 (N_2148,N_1042,N_311);
nor U2149 (N_2149,N_1445,N_497);
or U2150 (N_2150,N_660,N_1230);
xnor U2151 (N_2151,N_570,N_1035);
xnor U2152 (N_2152,N_589,N_394);
or U2153 (N_2153,N_303,N_1118);
and U2154 (N_2154,N_543,N_809);
nand U2155 (N_2155,N_567,N_121);
or U2156 (N_2156,N_864,N_1444);
and U2157 (N_2157,N_1223,N_1017);
xnor U2158 (N_2158,N_1111,N_1461);
or U2159 (N_2159,N_199,N_935);
nor U2160 (N_2160,N_1249,N_717);
or U2161 (N_2161,N_1337,N_815);
xnor U2162 (N_2162,N_533,N_1255);
nand U2163 (N_2163,N_44,N_1389);
or U2164 (N_2164,N_736,N_1269);
and U2165 (N_2165,N_1202,N_280);
xor U2166 (N_2166,N_899,N_597);
and U2167 (N_2167,N_928,N_1358);
xnor U2168 (N_2168,N_592,N_1007);
or U2169 (N_2169,N_1479,N_167);
and U2170 (N_2170,N_149,N_1054);
or U2171 (N_2171,N_651,N_510);
nor U2172 (N_2172,N_1431,N_1423);
xor U2173 (N_2173,N_1481,N_113);
xnor U2174 (N_2174,N_1025,N_1231);
xnor U2175 (N_2175,N_305,N_1305);
nor U2176 (N_2176,N_933,N_385);
nor U2177 (N_2177,N_583,N_1397);
nor U2178 (N_2178,N_1311,N_1182);
nand U2179 (N_2179,N_541,N_818);
or U2180 (N_2180,N_218,N_1234);
and U2181 (N_2181,N_869,N_1052);
xnor U2182 (N_2182,N_552,N_179);
xnor U2183 (N_2183,N_1167,N_442);
or U2184 (N_2184,N_1320,N_950);
and U2185 (N_2185,N_787,N_1225);
xnor U2186 (N_2186,N_488,N_49);
nor U2187 (N_2187,N_1379,N_437);
xnor U2188 (N_2188,N_258,N_139);
nor U2189 (N_2189,N_880,N_688);
nand U2190 (N_2190,N_1354,N_730);
and U2191 (N_2191,N_879,N_278);
or U2192 (N_2192,N_974,N_293);
or U2193 (N_2193,N_705,N_760);
nand U2194 (N_2194,N_249,N_400);
or U2195 (N_2195,N_1371,N_1072);
or U2196 (N_2196,N_1181,N_1009);
xnor U2197 (N_2197,N_421,N_1214);
nand U2198 (N_2198,N_1274,N_47);
or U2199 (N_2199,N_591,N_907);
or U2200 (N_2200,N_840,N_256);
or U2201 (N_2201,N_671,N_377);
nand U2202 (N_2202,N_656,N_1233);
and U2203 (N_2203,N_1226,N_1415);
and U2204 (N_2204,N_313,N_264);
and U2205 (N_2205,N_327,N_811);
nand U2206 (N_2206,N_43,N_802);
xor U2207 (N_2207,N_873,N_511);
and U2208 (N_2208,N_458,N_8);
and U2209 (N_2209,N_1116,N_604);
nand U2210 (N_2210,N_154,N_12);
or U2211 (N_2211,N_16,N_1081);
nor U2212 (N_2212,N_482,N_700);
and U2213 (N_2213,N_1399,N_111);
nor U2214 (N_2214,N_1172,N_623);
and U2215 (N_2215,N_1056,N_183);
xor U2216 (N_2216,N_1217,N_829);
nand U2217 (N_2217,N_453,N_568);
nor U2218 (N_2218,N_1316,N_1285);
xor U2219 (N_2219,N_1090,N_577);
nor U2220 (N_2220,N_126,N_1237);
and U2221 (N_2221,N_1110,N_168);
xnor U2222 (N_2222,N_599,N_637);
and U2223 (N_2223,N_6,N_683);
xnor U2224 (N_2224,N_129,N_1374);
or U2225 (N_2225,N_391,N_1075);
and U2226 (N_2226,N_226,N_460);
xnor U2227 (N_2227,N_119,N_66);
and U2228 (N_2228,N_114,N_1002);
and U2229 (N_2229,N_193,N_1351);
nand U2230 (N_2230,N_1030,N_1097);
nand U2231 (N_2231,N_643,N_1449);
and U2232 (N_2232,N_1184,N_365);
xor U2233 (N_2233,N_374,N_1256);
or U2234 (N_2234,N_812,N_1024);
xor U2235 (N_2235,N_1145,N_434);
nor U2236 (N_2236,N_1448,N_1077);
nand U2237 (N_2237,N_1438,N_959);
xnor U2238 (N_2238,N_1257,N_1362);
and U2239 (N_2239,N_521,N_1286);
and U2240 (N_2240,N_977,N_769);
and U2241 (N_2241,N_1453,N_157);
nor U2242 (N_2242,N_175,N_441);
xor U2243 (N_2243,N_761,N_3);
nand U2244 (N_2244,N_1185,N_1104);
nor U2245 (N_2245,N_100,N_941);
xor U2246 (N_2246,N_515,N_1435);
or U2247 (N_2247,N_233,N_1422);
nor U2248 (N_2248,N_1398,N_1287);
xor U2249 (N_2249,N_294,N_622);
nor U2250 (N_2250,N_637,N_655);
nor U2251 (N_2251,N_1442,N_1239);
or U2252 (N_2252,N_943,N_992);
or U2253 (N_2253,N_389,N_1377);
and U2254 (N_2254,N_1099,N_379);
xnor U2255 (N_2255,N_369,N_665);
xor U2256 (N_2256,N_1460,N_189);
xnor U2257 (N_2257,N_201,N_884);
and U2258 (N_2258,N_527,N_49);
or U2259 (N_2259,N_1332,N_223);
and U2260 (N_2260,N_231,N_118);
or U2261 (N_2261,N_783,N_1413);
or U2262 (N_2262,N_723,N_439);
xnor U2263 (N_2263,N_1236,N_512);
or U2264 (N_2264,N_1384,N_144);
xnor U2265 (N_2265,N_741,N_274);
or U2266 (N_2266,N_1229,N_535);
or U2267 (N_2267,N_117,N_1339);
nor U2268 (N_2268,N_873,N_308);
nor U2269 (N_2269,N_264,N_1240);
nand U2270 (N_2270,N_82,N_1293);
nand U2271 (N_2271,N_624,N_911);
nor U2272 (N_2272,N_581,N_1450);
nand U2273 (N_2273,N_1326,N_237);
nor U2274 (N_2274,N_595,N_1143);
xor U2275 (N_2275,N_6,N_26);
or U2276 (N_2276,N_458,N_1136);
and U2277 (N_2277,N_633,N_326);
xor U2278 (N_2278,N_670,N_631);
or U2279 (N_2279,N_865,N_1487);
nand U2280 (N_2280,N_661,N_769);
nand U2281 (N_2281,N_181,N_1195);
xnor U2282 (N_2282,N_715,N_677);
xnor U2283 (N_2283,N_124,N_540);
and U2284 (N_2284,N_1238,N_1363);
xnor U2285 (N_2285,N_1016,N_1115);
nand U2286 (N_2286,N_1115,N_952);
nor U2287 (N_2287,N_1411,N_154);
xor U2288 (N_2288,N_1488,N_144);
xor U2289 (N_2289,N_130,N_146);
and U2290 (N_2290,N_972,N_978);
nand U2291 (N_2291,N_1151,N_1324);
nand U2292 (N_2292,N_353,N_1046);
and U2293 (N_2293,N_366,N_588);
and U2294 (N_2294,N_1457,N_1075);
and U2295 (N_2295,N_1217,N_1332);
or U2296 (N_2296,N_105,N_15);
and U2297 (N_2297,N_1136,N_496);
xor U2298 (N_2298,N_804,N_753);
or U2299 (N_2299,N_1139,N_534);
xor U2300 (N_2300,N_203,N_595);
and U2301 (N_2301,N_528,N_1290);
nand U2302 (N_2302,N_1462,N_557);
nand U2303 (N_2303,N_970,N_945);
and U2304 (N_2304,N_970,N_387);
nand U2305 (N_2305,N_1459,N_744);
nor U2306 (N_2306,N_1256,N_1067);
nor U2307 (N_2307,N_1156,N_520);
or U2308 (N_2308,N_609,N_69);
nand U2309 (N_2309,N_1131,N_613);
xor U2310 (N_2310,N_1405,N_301);
or U2311 (N_2311,N_1466,N_673);
xor U2312 (N_2312,N_420,N_684);
and U2313 (N_2313,N_417,N_962);
nor U2314 (N_2314,N_492,N_1010);
nand U2315 (N_2315,N_1052,N_1274);
nor U2316 (N_2316,N_1420,N_1113);
nand U2317 (N_2317,N_1046,N_1480);
nand U2318 (N_2318,N_1237,N_442);
and U2319 (N_2319,N_1066,N_20);
nand U2320 (N_2320,N_431,N_577);
and U2321 (N_2321,N_1097,N_284);
xor U2322 (N_2322,N_591,N_1189);
nor U2323 (N_2323,N_330,N_451);
xnor U2324 (N_2324,N_660,N_1458);
nand U2325 (N_2325,N_117,N_1109);
nor U2326 (N_2326,N_1104,N_1320);
nor U2327 (N_2327,N_551,N_921);
or U2328 (N_2328,N_523,N_151);
nor U2329 (N_2329,N_1476,N_1038);
nor U2330 (N_2330,N_985,N_742);
nand U2331 (N_2331,N_1152,N_1490);
xnor U2332 (N_2332,N_624,N_968);
or U2333 (N_2333,N_1258,N_744);
nand U2334 (N_2334,N_1200,N_707);
and U2335 (N_2335,N_103,N_466);
or U2336 (N_2336,N_1359,N_379);
nand U2337 (N_2337,N_867,N_308);
and U2338 (N_2338,N_349,N_1225);
or U2339 (N_2339,N_877,N_403);
xnor U2340 (N_2340,N_116,N_474);
nand U2341 (N_2341,N_1130,N_262);
xor U2342 (N_2342,N_495,N_1120);
nand U2343 (N_2343,N_413,N_1035);
or U2344 (N_2344,N_381,N_167);
xnor U2345 (N_2345,N_1015,N_883);
xor U2346 (N_2346,N_1020,N_523);
nand U2347 (N_2347,N_851,N_195);
and U2348 (N_2348,N_294,N_504);
nand U2349 (N_2349,N_102,N_418);
nand U2350 (N_2350,N_1245,N_511);
and U2351 (N_2351,N_1160,N_410);
and U2352 (N_2352,N_1045,N_1141);
xor U2353 (N_2353,N_576,N_223);
nor U2354 (N_2354,N_219,N_1195);
xnor U2355 (N_2355,N_851,N_227);
nand U2356 (N_2356,N_201,N_1211);
xor U2357 (N_2357,N_253,N_1162);
or U2358 (N_2358,N_1065,N_486);
nor U2359 (N_2359,N_594,N_1349);
and U2360 (N_2360,N_1153,N_772);
nor U2361 (N_2361,N_85,N_1235);
nand U2362 (N_2362,N_286,N_79);
or U2363 (N_2363,N_54,N_1455);
xnor U2364 (N_2364,N_647,N_996);
or U2365 (N_2365,N_549,N_457);
and U2366 (N_2366,N_479,N_886);
nor U2367 (N_2367,N_1495,N_1293);
nor U2368 (N_2368,N_625,N_806);
nor U2369 (N_2369,N_1157,N_561);
nor U2370 (N_2370,N_819,N_1334);
nand U2371 (N_2371,N_1420,N_301);
and U2372 (N_2372,N_293,N_1008);
xnor U2373 (N_2373,N_391,N_1024);
nand U2374 (N_2374,N_290,N_951);
nand U2375 (N_2375,N_433,N_151);
and U2376 (N_2376,N_450,N_156);
xnor U2377 (N_2377,N_362,N_1284);
nand U2378 (N_2378,N_293,N_1419);
nand U2379 (N_2379,N_1086,N_11);
and U2380 (N_2380,N_672,N_162);
nor U2381 (N_2381,N_756,N_912);
and U2382 (N_2382,N_754,N_1385);
or U2383 (N_2383,N_82,N_1024);
nand U2384 (N_2384,N_1237,N_744);
or U2385 (N_2385,N_1342,N_484);
xor U2386 (N_2386,N_1438,N_1308);
nor U2387 (N_2387,N_1366,N_206);
nand U2388 (N_2388,N_19,N_1316);
and U2389 (N_2389,N_1091,N_277);
nand U2390 (N_2390,N_652,N_327);
nand U2391 (N_2391,N_66,N_951);
nand U2392 (N_2392,N_926,N_1350);
xor U2393 (N_2393,N_742,N_1187);
or U2394 (N_2394,N_1347,N_258);
xnor U2395 (N_2395,N_841,N_444);
xnor U2396 (N_2396,N_791,N_139);
or U2397 (N_2397,N_169,N_1191);
or U2398 (N_2398,N_940,N_702);
and U2399 (N_2399,N_1021,N_783);
and U2400 (N_2400,N_760,N_530);
xnor U2401 (N_2401,N_707,N_750);
nor U2402 (N_2402,N_1002,N_1020);
or U2403 (N_2403,N_24,N_1289);
xnor U2404 (N_2404,N_450,N_750);
nand U2405 (N_2405,N_1213,N_121);
and U2406 (N_2406,N_271,N_59);
nand U2407 (N_2407,N_977,N_1366);
or U2408 (N_2408,N_1483,N_463);
xnor U2409 (N_2409,N_419,N_1322);
xor U2410 (N_2410,N_583,N_253);
xnor U2411 (N_2411,N_1045,N_1170);
nor U2412 (N_2412,N_1432,N_1451);
and U2413 (N_2413,N_960,N_85);
and U2414 (N_2414,N_990,N_1354);
and U2415 (N_2415,N_1063,N_229);
or U2416 (N_2416,N_909,N_1335);
xor U2417 (N_2417,N_1060,N_1416);
or U2418 (N_2418,N_456,N_613);
or U2419 (N_2419,N_1496,N_391);
or U2420 (N_2420,N_479,N_1497);
or U2421 (N_2421,N_2,N_105);
nor U2422 (N_2422,N_1490,N_937);
or U2423 (N_2423,N_149,N_956);
xnor U2424 (N_2424,N_277,N_1233);
nor U2425 (N_2425,N_1213,N_1362);
and U2426 (N_2426,N_675,N_576);
and U2427 (N_2427,N_1470,N_583);
and U2428 (N_2428,N_927,N_26);
nor U2429 (N_2429,N_157,N_1267);
xnor U2430 (N_2430,N_533,N_1022);
nor U2431 (N_2431,N_888,N_438);
nand U2432 (N_2432,N_964,N_562);
nor U2433 (N_2433,N_987,N_829);
nor U2434 (N_2434,N_167,N_1218);
xor U2435 (N_2435,N_953,N_1340);
or U2436 (N_2436,N_257,N_381);
nor U2437 (N_2437,N_168,N_298);
or U2438 (N_2438,N_373,N_1417);
or U2439 (N_2439,N_337,N_164);
and U2440 (N_2440,N_286,N_564);
or U2441 (N_2441,N_140,N_1219);
nor U2442 (N_2442,N_1340,N_797);
and U2443 (N_2443,N_1316,N_1294);
or U2444 (N_2444,N_328,N_752);
nand U2445 (N_2445,N_462,N_1222);
nand U2446 (N_2446,N_1173,N_824);
nand U2447 (N_2447,N_1357,N_441);
nor U2448 (N_2448,N_890,N_1013);
nor U2449 (N_2449,N_898,N_1072);
xnor U2450 (N_2450,N_1233,N_1143);
or U2451 (N_2451,N_1176,N_376);
nand U2452 (N_2452,N_1332,N_1361);
or U2453 (N_2453,N_233,N_81);
and U2454 (N_2454,N_1341,N_819);
or U2455 (N_2455,N_714,N_713);
or U2456 (N_2456,N_180,N_1293);
and U2457 (N_2457,N_423,N_451);
nor U2458 (N_2458,N_1089,N_18);
and U2459 (N_2459,N_159,N_1429);
and U2460 (N_2460,N_1344,N_526);
or U2461 (N_2461,N_1334,N_348);
or U2462 (N_2462,N_463,N_1076);
xor U2463 (N_2463,N_591,N_1331);
or U2464 (N_2464,N_712,N_738);
and U2465 (N_2465,N_398,N_1402);
nand U2466 (N_2466,N_1221,N_1168);
nor U2467 (N_2467,N_933,N_1181);
nand U2468 (N_2468,N_30,N_302);
nor U2469 (N_2469,N_1466,N_672);
and U2470 (N_2470,N_426,N_1333);
nand U2471 (N_2471,N_1310,N_99);
xnor U2472 (N_2472,N_1100,N_966);
xor U2473 (N_2473,N_1299,N_693);
or U2474 (N_2474,N_120,N_676);
or U2475 (N_2475,N_1061,N_430);
nor U2476 (N_2476,N_958,N_344);
nor U2477 (N_2477,N_685,N_432);
nor U2478 (N_2478,N_460,N_393);
and U2479 (N_2479,N_1037,N_1134);
and U2480 (N_2480,N_356,N_514);
nor U2481 (N_2481,N_247,N_808);
xor U2482 (N_2482,N_950,N_1437);
nor U2483 (N_2483,N_914,N_609);
or U2484 (N_2484,N_1179,N_509);
nand U2485 (N_2485,N_1154,N_1306);
nor U2486 (N_2486,N_1269,N_544);
and U2487 (N_2487,N_516,N_832);
or U2488 (N_2488,N_806,N_1048);
xnor U2489 (N_2489,N_406,N_249);
xnor U2490 (N_2490,N_592,N_169);
nor U2491 (N_2491,N_1051,N_1145);
and U2492 (N_2492,N_501,N_621);
nor U2493 (N_2493,N_435,N_35);
and U2494 (N_2494,N_605,N_390);
or U2495 (N_2495,N_1263,N_417);
nor U2496 (N_2496,N_320,N_534);
xor U2497 (N_2497,N_325,N_15);
nand U2498 (N_2498,N_215,N_945);
and U2499 (N_2499,N_43,N_357);
and U2500 (N_2500,N_108,N_471);
and U2501 (N_2501,N_383,N_211);
or U2502 (N_2502,N_1144,N_952);
nand U2503 (N_2503,N_1025,N_943);
and U2504 (N_2504,N_117,N_1434);
xor U2505 (N_2505,N_964,N_1058);
nand U2506 (N_2506,N_1013,N_360);
and U2507 (N_2507,N_1037,N_351);
xnor U2508 (N_2508,N_746,N_707);
nand U2509 (N_2509,N_1332,N_663);
nand U2510 (N_2510,N_1113,N_1400);
xnor U2511 (N_2511,N_307,N_613);
or U2512 (N_2512,N_1353,N_938);
or U2513 (N_2513,N_1074,N_384);
or U2514 (N_2514,N_1313,N_1127);
nor U2515 (N_2515,N_72,N_526);
xnor U2516 (N_2516,N_368,N_754);
nor U2517 (N_2517,N_1463,N_551);
xor U2518 (N_2518,N_709,N_611);
xnor U2519 (N_2519,N_608,N_454);
and U2520 (N_2520,N_1072,N_1073);
nand U2521 (N_2521,N_658,N_431);
xor U2522 (N_2522,N_824,N_598);
nor U2523 (N_2523,N_447,N_1171);
nor U2524 (N_2524,N_511,N_151);
nor U2525 (N_2525,N_457,N_538);
nor U2526 (N_2526,N_426,N_767);
nor U2527 (N_2527,N_517,N_913);
xnor U2528 (N_2528,N_1050,N_29);
and U2529 (N_2529,N_380,N_676);
or U2530 (N_2530,N_81,N_10);
xor U2531 (N_2531,N_1308,N_1400);
nor U2532 (N_2532,N_858,N_1078);
and U2533 (N_2533,N_774,N_691);
xor U2534 (N_2534,N_1312,N_1356);
nand U2535 (N_2535,N_1363,N_1131);
nand U2536 (N_2536,N_555,N_8);
or U2537 (N_2537,N_1249,N_639);
xnor U2538 (N_2538,N_1108,N_787);
xnor U2539 (N_2539,N_545,N_1483);
and U2540 (N_2540,N_1324,N_29);
nor U2541 (N_2541,N_948,N_585);
nand U2542 (N_2542,N_638,N_701);
and U2543 (N_2543,N_78,N_861);
and U2544 (N_2544,N_848,N_949);
or U2545 (N_2545,N_837,N_673);
nand U2546 (N_2546,N_1039,N_1379);
nor U2547 (N_2547,N_1057,N_1276);
or U2548 (N_2548,N_364,N_983);
or U2549 (N_2549,N_1244,N_561);
nor U2550 (N_2550,N_64,N_366);
or U2551 (N_2551,N_1498,N_108);
or U2552 (N_2552,N_402,N_819);
nor U2553 (N_2553,N_120,N_1109);
nand U2554 (N_2554,N_343,N_1486);
or U2555 (N_2555,N_1081,N_587);
nand U2556 (N_2556,N_991,N_447);
xnor U2557 (N_2557,N_976,N_924);
nand U2558 (N_2558,N_1255,N_990);
nor U2559 (N_2559,N_889,N_1183);
nand U2560 (N_2560,N_960,N_1111);
and U2561 (N_2561,N_1468,N_873);
xnor U2562 (N_2562,N_1413,N_600);
nor U2563 (N_2563,N_1468,N_415);
xor U2564 (N_2564,N_829,N_592);
and U2565 (N_2565,N_355,N_1074);
and U2566 (N_2566,N_1401,N_1459);
nor U2567 (N_2567,N_187,N_277);
nor U2568 (N_2568,N_1256,N_769);
and U2569 (N_2569,N_1366,N_269);
xor U2570 (N_2570,N_1421,N_207);
nor U2571 (N_2571,N_1251,N_454);
and U2572 (N_2572,N_965,N_762);
and U2573 (N_2573,N_48,N_654);
nand U2574 (N_2574,N_1104,N_790);
nor U2575 (N_2575,N_1439,N_171);
nand U2576 (N_2576,N_671,N_226);
or U2577 (N_2577,N_40,N_1241);
and U2578 (N_2578,N_1164,N_855);
xor U2579 (N_2579,N_872,N_226);
and U2580 (N_2580,N_225,N_658);
xor U2581 (N_2581,N_465,N_732);
nand U2582 (N_2582,N_1499,N_898);
or U2583 (N_2583,N_1325,N_655);
nor U2584 (N_2584,N_762,N_1353);
and U2585 (N_2585,N_1263,N_1087);
nor U2586 (N_2586,N_836,N_545);
xnor U2587 (N_2587,N_447,N_284);
nand U2588 (N_2588,N_517,N_1339);
xnor U2589 (N_2589,N_1405,N_772);
or U2590 (N_2590,N_1054,N_66);
nand U2591 (N_2591,N_616,N_1171);
or U2592 (N_2592,N_1002,N_921);
xnor U2593 (N_2593,N_528,N_1274);
or U2594 (N_2594,N_282,N_1478);
xor U2595 (N_2595,N_702,N_182);
or U2596 (N_2596,N_1299,N_1197);
and U2597 (N_2597,N_1426,N_309);
nand U2598 (N_2598,N_15,N_186);
xnor U2599 (N_2599,N_634,N_1455);
nand U2600 (N_2600,N_884,N_1413);
nor U2601 (N_2601,N_166,N_895);
or U2602 (N_2602,N_1212,N_561);
or U2603 (N_2603,N_567,N_445);
nand U2604 (N_2604,N_684,N_62);
nand U2605 (N_2605,N_1008,N_1437);
nand U2606 (N_2606,N_1143,N_696);
and U2607 (N_2607,N_527,N_394);
nor U2608 (N_2608,N_65,N_1401);
and U2609 (N_2609,N_1352,N_359);
nor U2610 (N_2610,N_1109,N_515);
and U2611 (N_2611,N_108,N_1441);
nand U2612 (N_2612,N_936,N_1459);
and U2613 (N_2613,N_365,N_892);
or U2614 (N_2614,N_37,N_1101);
xnor U2615 (N_2615,N_1478,N_320);
xnor U2616 (N_2616,N_191,N_241);
nand U2617 (N_2617,N_440,N_160);
and U2618 (N_2618,N_1138,N_1161);
nor U2619 (N_2619,N_651,N_1287);
nor U2620 (N_2620,N_326,N_1458);
xor U2621 (N_2621,N_386,N_820);
nand U2622 (N_2622,N_555,N_1288);
nand U2623 (N_2623,N_959,N_1467);
or U2624 (N_2624,N_1361,N_1006);
xor U2625 (N_2625,N_645,N_1316);
xnor U2626 (N_2626,N_161,N_1293);
and U2627 (N_2627,N_242,N_389);
and U2628 (N_2628,N_977,N_668);
or U2629 (N_2629,N_870,N_977);
or U2630 (N_2630,N_641,N_1484);
nor U2631 (N_2631,N_696,N_745);
or U2632 (N_2632,N_1462,N_538);
xnor U2633 (N_2633,N_990,N_929);
xnor U2634 (N_2634,N_1376,N_309);
nor U2635 (N_2635,N_1277,N_66);
or U2636 (N_2636,N_865,N_1296);
and U2637 (N_2637,N_1359,N_25);
and U2638 (N_2638,N_210,N_763);
nor U2639 (N_2639,N_1119,N_725);
and U2640 (N_2640,N_1442,N_377);
and U2641 (N_2641,N_1292,N_1477);
or U2642 (N_2642,N_108,N_1008);
xor U2643 (N_2643,N_1189,N_307);
xnor U2644 (N_2644,N_1,N_1216);
nand U2645 (N_2645,N_1308,N_1152);
and U2646 (N_2646,N_726,N_261);
and U2647 (N_2647,N_1216,N_1143);
and U2648 (N_2648,N_1413,N_609);
or U2649 (N_2649,N_427,N_47);
or U2650 (N_2650,N_524,N_1289);
nor U2651 (N_2651,N_425,N_203);
nand U2652 (N_2652,N_582,N_824);
nor U2653 (N_2653,N_1016,N_1125);
and U2654 (N_2654,N_843,N_890);
xor U2655 (N_2655,N_126,N_461);
and U2656 (N_2656,N_1129,N_782);
or U2657 (N_2657,N_1377,N_982);
nand U2658 (N_2658,N_910,N_339);
and U2659 (N_2659,N_663,N_40);
or U2660 (N_2660,N_395,N_855);
nand U2661 (N_2661,N_151,N_707);
nor U2662 (N_2662,N_960,N_542);
or U2663 (N_2663,N_1073,N_1037);
nand U2664 (N_2664,N_1069,N_1312);
or U2665 (N_2665,N_911,N_442);
nor U2666 (N_2666,N_563,N_1325);
nor U2667 (N_2667,N_269,N_423);
nor U2668 (N_2668,N_1021,N_1127);
nand U2669 (N_2669,N_645,N_229);
or U2670 (N_2670,N_173,N_447);
and U2671 (N_2671,N_162,N_1024);
nand U2672 (N_2672,N_757,N_1446);
nand U2673 (N_2673,N_499,N_1489);
xnor U2674 (N_2674,N_1231,N_1447);
nor U2675 (N_2675,N_549,N_391);
xor U2676 (N_2676,N_118,N_826);
nand U2677 (N_2677,N_308,N_706);
nand U2678 (N_2678,N_263,N_971);
or U2679 (N_2679,N_1212,N_1310);
xnor U2680 (N_2680,N_1433,N_1347);
nor U2681 (N_2681,N_17,N_1164);
xnor U2682 (N_2682,N_1101,N_646);
nand U2683 (N_2683,N_158,N_51);
or U2684 (N_2684,N_1023,N_1004);
xor U2685 (N_2685,N_1033,N_357);
nand U2686 (N_2686,N_949,N_802);
nand U2687 (N_2687,N_1499,N_1185);
or U2688 (N_2688,N_615,N_941);
nor U2689 (N_2689,N_10,N_1430);
xnor U2690 (N_2690,N_1314,N_141);
xnor U2691 (N_2691,N_680,N_452);
and U2692 (N_2692,N_836,N_650);
nor U2693 (N_2693,N_775,N_179);
xor U2694 (N_2694,N_449,N_1476);
and U2695 (N_2695,N_62,N_733);
nand U2696 (N_2696,N_253,N_457);
xnor U2697 (N_2697,N_1440,N_1479);
xor U2698 (N_2698,N_1069,N_431);
and U2699 (N_2699,N_1151,N_171);
nor U2700 (N_2700,N_1448,N_1127);
nor U2701 (N_2701,N_1277,N_236);
nor U2702 (N_2702,N_481,N_1221);
and U2703 (N_2703,N_1220,N_1427);
xor U2704 (N_2704,N_680,N_772);
and U2705 (N_2705,N_1232,N_982);
or U2706 (N_2706,N_505,N_774);
and U2707 (N_2707,N_762,N_155);
and U2708 (N_2708,N_1202,N_1434);
or U2709 (N_2709,N_266,N_807);
nand U2710 (N_2710,N_549,N_241);
xnor U2711 (N_2711,N_1088,N_300);
nor U2712 (N_2712,N_1321,N_1072);
nand U2713 (N_2713,N_1053,N_755);
and U2714 (N_2714,N_1043,N_1421);
nor U2715 (N_2715,N_864,N_371);
and U2716 (N_2716,N_754,N_451);
nand U2717 (N_2717,N_378,N_66);
nor U2718 (N_2718,N_1049,N_1091);
and U2719 (N_2719,N_1117,N_821);
nor U2720 (N_2720,N_1047,N_35);
xor U2721 (N_2721,N_1332,N_648);
and U2722 (N_2722,N_1055,N_1029);
nand U2723 (N_2723,N_120,N_292);
nor U2724 (N_2724,N_1222,N_181);
nor U2725 (N_2725,N_1176,N_875);
and U2726 (N_2726,N_1391,N_306);
xor U2727 (N_2727,N_571,N_628);
and U2728 (N_2728,N_508,N_1066);
or U2729 (N_2729,N_854,N_1142);
nand U2730 (N_2730,N_491,N_406);
nor U2731 (N_2731,N_1341,N_28);
and U2732 (N_2732,N_1255,N_676);
xnor U2733 (N_2733,N_1279,N_1251);
nand U2734 (N_2734,N_58,N_764);
nor U2735 (N_2735,N_1361,N_52);
nor U2736 (N_2736,N_792,N_795);
nand U2737 (N_2737,N_969,N_358);
nand U2738 (N_2738,N_1015,N_1084);
nor U2739 (N_2739,N_1381,N_1428);
and U2740 (N_2740,N_312,N_830);
or U2741 (N_2741,N_720,N_1300);
and U2742 (N_2742,N_43,N_1350);
nand U2743 (N_2743,N_1055,N_721);
nor U2744 (N_2744,N_371,N_1453);
and U2745 (N_2745,N_1126,N_1270);
xnor U2746 (N_2746,N_284,N_840);
xor U2747 (N_2747,N_915,N_1108);
xnor U2748 (N_2748,N_367,N_280);
xor U2749 (N_2749,N_1362,N_796);
or U2750 (N_2750,N_116,N_1311);
nand U2751 (N_2751,N_14,N_820);
nand U2752 (N_2752,N_380,N_709);
xnor U2753 (N_2753,N_1050,N_1028);
or U2754 (N_2754,N_1219,N_812);
xnor U2755 (N_2755,N_603,N_135);
or U2756 (N_2756,N_1080,N_841);
xnor U2757 (N_2757,N_895,N_514);
xnor U2758 (N_2758,N_1227,N_938);
or U2759 (N_2759,N_760,N_1153);
nand U2760 (N_2760,N_791,N_876);
nor U2761 (N_2761,N_991,N_628);
and U2762 (N_2762,N_921,N_274);
nand U2763 (N_2763,N_268,N_1042);
or U2764 (N_2764,N_1335,N_431);
nand U2765 (N_2765,N_935,N_10);
xnor U2766 (N_2766,N_1115,N_1371);
xor U2767 (N_2767,N_361,N_1092);
or U2768 (N_2768,N_242,N_486);
or U2769 (N_2769,N_1127,N_509);
or U2770 (N_2770,N_987,N_1368);
xor U2771 (N_2771,N_183,N_509);
or U2772 (N_2772,N_700,N_1095);
xor U2773 (N_2773,N_1385,N_343);
nand U2774 (N_2774,N_1129,N_1406);
and U2775 (N_2775,N_763,N_621);
nand U2776 (N_2776,N_1402,N_1363);
or U2777 (N_2777,N_616,N_41);
nor U2778 (N_2778,N_290,N_1209);
and U2779 (N_2779,N_1018,N_1246);
nand U2780 (N_2780,N_40,N_1073);
and U2781 (N_2781,N_973,N_694);
xnor U2782 (N_2782,N_1170,N_334);
and U2783 (N_2783,N_6,N_198);
or U2784 (N_2784,N_1222,N_282);
nand U2785 (N_2785,N_1060,N_1471);
and U2786 (N_2786,N_1143,N_407);
nor U2787 (N_2787,N_742,N_1155);
or U2788 (N_2788,N_487,N_1449);
or U2789 (N_2789,N_346,N_1302);
or U2790 (N_2790,N_358,N_119);
nor U2791 (N_2791,N_130,N_812);
and U2792 (N_2792,N_1427,N_44);
or U2793 (N_2793,N_246,N_293);
nand U2794 (N_2794,N_520,N_13);
and U2795 (N_2795,N_1183,N_1141);
or U2796 (N_2796,N_293,N_1241);
or U2797 (N_2797,N_626,N_563);
and U2798 (N_2798,N_1047,N_681);
or U2799 (N_2799,N_1244,N_873);
nor U2800 (N_2800,N_689,N_67);
nor U2801 (N_2801,N_619,N_229);
and U2802 (N_2802,N_32,N_1486);
xnor U2803 (N_2803,N_1354,N_101);
nor U2804 (N_2804,N_526,N_1266);
nand U2805 (N_2805,N_882,N_1400);
nand U2806 (N_2806,N_1151,N_774);
and U2807 (N_2807,N_842,N_81);
and U2808 (N_2808,N_1148,N_377);
and U2809 (N_2809,N_1412,N_1144);
and U2810 (N_2810,N_1110,N_1055);
and U2811 (N_2811,N_967,N_634);
and U2812 (N_2812,N_672,N_712);
and U2813 (N_2813,N_549,N_187);
nand U2814 (N_2814,N_1025,N_694);
or U2815 (N_2815,N_759,N_869);
nor U2816 (N_2816,N_275,N_55);
nand U2817 (N_2817,N_354,N_455);
or U2818 (N_2818,N_710,N_1326);
or U2819 (N_2819,N_744,N_1144);
xor U2820 (N_2820,N_341,N_778);
xor U2821 (N_2821,N_340,N_873);
and U2822 (N_2822,N_309,N_756);
xor U2823 (N_2823,N_140,N_1409);
and U2824 (N_2824,N_152,N_1134);
nor U2825 (N_2825,N_1270,N_891);
nor U2826 (N_2826,N_1014,N_1135);
and U2827 (N_2827,N_1499,N_588);
and U2828 (N_2828,N_945,N_783);
or U2829 (N_2829,N_30,N_1341);
and U2830 (N_2830,N_1346,N_373);
xnor U2831 (N_2831,N_1295,N_644);
or U2832 (N_2832,N_790,N_628);
nor U2833 (N_2833,N_662,N_108);
and U2834 (N_2834,N_11,N_58);
nand U2835 (N_2835,N_1181,N_308);
xnor U2836 (N_2836,N_615,N_238);
or U2837 (N_2837,N_334,N_563);
xor U2838 (N_2838,N_1451,N_468);
and U2839 (N_2839,N_552,N_662);
and U2840 (N_2840,N_607,N_1273);
and U2841 (N_2841,N_88,N_1129);
xor U2842 (N_2842,N_1206,N_41);
nor U2843 (N_2843,N_1405,N_842);
nand U2844 (N_2844,N_1187,N_609);
nor U2845 (N_2845,N_618,N_1428);
xor U2846 (N_2846,N_752,N_1046);
and U2847 (N_2847,N_420,N_84);
nand U2848 (N_2848,N_175,N_111);
nor U2849 (N_2849,N_331,N_898);
nand U2850 (N_2850,N_318,N_1119);
xor U2851 (N_2851,N_1356,N_1072);
or U2852 (N_2852,N_272,N_47);
xnor U2853 (N_2853,N_982,N_12);
xor U2854 (N_2854,N_1225,N_190);
xnor U2855 (N_2855,N_353,N_802);
nand U2856 (N_2856,N_1207,N_429);
nand U2857 (N_2857,N_1116,N_939);
and U2858 (N_2858,N_24,N_948);
nor U2859 (N_2859,N_1196,N_389);
and U2860 (N_2860,N_1485,N_478);
nor U2861 (N_2861,N_453,N_843);
nand U2862 (N_2862,N_1025,N_1156);
xnor U2863 (N_2863,N_442,N_1137);
xnor U2864 (N_2864,N_187,N_763);
xnor U2865 (N_2865,N_1259,N_357);
nand U2866 (N_2866,N_1062,N_572);
and U2867 (N_2867,N_405,N_1322);
nand U2868 (N_2868,N_124,N_573);
xor U2869 (N_2869,N_331,N_607);
nor U2870 (N_2870,N_154,N_630);
xnor U2871 (N_2871,N_638,N_129);
or U2872 (N_2872,N_1032,N_4);
and U2873 (N_2873,N_420,N_209);
nand U2874 (N_2874,N_1278,N_335);
xnor U2875 (N_2875,N_1313,N_1140);
nand U2876 (N_2876,N_511,N_568);
and U2877 (N_2877,N_443,N_989);
or U2878 (N_2878,N_751,N_784);
nor U2879 (N_2879,N_941,N_218);
xnor U2880 (N_2880,N_685,N_1156);
xnor U2881 (N_2881,N_872,N_464);
nand U2882 (N_2882,N_437,N_1193);
xor U2883 (N_2883,N_1136,N_708);
or U2884 (N_2884,N_1285,N_1071);
nand U2885 (N_2885,N_1303,N_785);
or U2886 (N_2886,N_275,N_270);
xor U2887 (N_2887,N_907,N_466);
nor U2888 (N_2888,N_948,N_1026);
nand U2889 (N_2889,N_728,N_467);
nor U2890 (N_2890,N_641,N_290);
nand U2891 (N_2891,N_899,N_768);
and U2892 (N_2892,N_1435,N_1283);
nand U2893 (N_2893,N_403,N_1114);
xor U2894 (N_2894,N_981,N_1113);
or U2895 (N_2895,N_1018,N_15);
nor U2896 (N_2896,N_824,N_862);
nand U2897 (N_2897,N_444,N_1459);
xor U2898 (N_2898,N_1182,N_338);
and U2899 (N_2899,N_253,N_559);
and U2900 (N_2900,N_1280,N_1029);
nor U2901 (N_2901,N_320,N_349);
nor U2902 (N_2902,N_1224,N_1476);
xor U2903 (N_2903,N_1261,N_1042);
or U2904 (N_2904,N_1461,N_1133);
and U2905 (N_2905,N_630,N_1079);
nor U2906 (N_2906,N_222,N_323);
nand U2907 (N_2907,N_549,N_1095);
xor U2908 (N_2908,N_1440,N_1328);
nor U2909 (N_2909,N_454,N_1300);
nand U2910 (N_2910,N_63,N_753);
or U2911 (N_2911,N_45,N_132);
xnor U2912 (N_2912,N_218,N_645);
and U2913 (N_2913,N_288,N_419);
nand U2914 (N_2914,N_605,N_1052);
xor U2915 (N_2915,N_133,N_1029);
nand U2916 (N_2916,N_1083,N_711);
and U2917 (N_2917,N_26,N_832);
or U2918 (N_2918,N_76,N_60);
nor U2919 (N_2919,N_284,N_1493);
nor U2920 (N_2920,N_792,N_111);
or U2921 (N_2921,N_978,N_894);
xor U2922 (N_2922,N_425,N_854);
nor U2923 (N_2923,N_1089,N_837);
nand U2924 (N_2924,N_0,N_885);
nand U2925 (N_2925,N_1364,N_1462);
xor U2926 (N_2926,N_163,N_340);
nor U2927 (N_2927,N_1082,N_682);
nor U2928 (N_2928,N_107,N_1029);
nand U2929 (N_2929,N_1321,N_205);
xor U2930 (N_2930,N_416,N_929);
or U2931 (N_2931,N_395,N_714);
nand U2932 (N_2932,N_659,N_1082);
nor U2933 (N_2933,N_139,N_449);
xor U2934 (N_2934,N_1078,N_230);
nor U2935 (N_2935,N_1312,N_641);
nand U2936 (N_2936,N_1450,N_405);
and U2937 (N_2937,N_662,N_851);
nand U2938 (N_2938,N_296,N_424);
xnor U2939 (N_2939,N_1244,N_651);
xor U2940 (N_2940,N_728,N_255);
or U2941 (N_2941,N_1179,N_886);
or U2942 (N_2942,N_342,N_716);
nand U2943 (N_2943,N_1477,N_20);
and U2944 (N_2944,N_1343,N_291);
or U2945 (N_2945,N_22,N_229);
nor U2946 (N_2946,N_318,N_1370);
or U2947 (N_2947,N_389,N_437);
xor U2948 (N_2948,N_402,N_1130);
nor U2949 (N_2949,N_848,N_926);
and U2950 (N_2950,N_21,N_309);
or U2951 (N_2951,N_1473,N_162);
xor U2952 (N_2952,N_526,N_39);
or U2953 (N_2953,N_1101,N_322);
or U2954 (N_2954,N_1294,N_925);
or U2955 (N_2955,N_977,N_808);
nand U2956 (N_2956,N_1403,N_415);
nor U2957 (N_2957,N_973,N_1102);
xor U2958 (N_2958,N_1471,N_710);
or U2959 (N_2959,N_789,N_899);
nand U2960 (N_2960,N_865,N_1417);
or U2961 (N_2961,N_219,N_1097);
nor U2962 (N_2962,N_1252,N_1479);
nor U2963 (N_2963,N_908,N_270);
and U2964 (N_2964,N_998,N_937);
nand U2965 (N_2965,N_17,N_1270);
xnor U2966 (N_2966,N_1379,N_286);
and U2967 (N_2967,N_810,N_727);
or U2968 (N_2968,N_157,N_810);
nor U2969 (N_2969,N_1010,N_1271);
or U2970 (N_2970,N_1353,N_951);
and U2971 (N_2971,N_679,N_694);
or U2972 (N_2972,N_742,N_1447);
nand U2973 (N_2973,N_1471,N_624);
or U2974 (N_2974,N_661,N_843);
xor U2975 (N_2975,N_1275,N_1270);
nand U2976 (N_2976,N_248,N_1391);
and U2977 (N_2977,N_1275,N_438);
and U2978 (N_2978,N_233,N_184);
and U2979 (N_2979,N_957,N_1303);
nand U2980 (N_2980,N_1382,N_1363);
nand U2981 (N_2981,N_1077,N_384);
xor U2982 (N_2982,N_703,N_1425);
nor U2983 (N_2983,N_1471,N_816);
xnor U2984 (N_2984,N_1366,N_496);
xor U2985 (N_2985,N_184,N_647);
or U2986 (N_2986,N_593,N_388);
nand U2987 (N_2987,N_985,N_549);
nor U2988 (N_2988,N_716,N_919);
nor U2989 (N_2989,N_490,N_1131);
nor U2990 (N_2990,N_410,N_70);
and U2991 (N_2991,N_1281,N_271);
or U2992 (N_2992,N_861,N_1268);
nand U2993 (N_2993,N_563,N_585);
xor U2994 (N_2994,N_1277,N_401);
xnor U2995 (N_2995,N_81,N_932);
xnor U2996 (N_2996,N_751,N_125);
nor U2997 (N_2997,N_639,N_696);
xor U2998 (N_2998,N_472,N_154);
and U2999 (N_2999,N_591,N_722);
and U3000 (N_3000,N_1728,N_2397);
nor U3001 (N_3001,N_2995,N_2669);
or U3002 (N_3002,N_2857,N_2057);
or U3003 (N_3003,N_2761,N_2383);
nor U3004 (N_3004,N_1929,N_1545);
or U3005 (N_3005,N_2897,N_1730);
nand U3006 (N_3006,N_2035,N_1660);
and U3007 (N_3007,N_2676,N_2513);
or U3008 (N_3008,N_2387,N_2329);
xnor U3009 (N_3009,N_2644,N_1788);
and U3010 (N_3010,N_1529,N_2093);
and U3011 (N_3011,N_2061,N_2620);
or U3012 (N_3012,N_1518,N_1790);
and U3013 (N_3013,N_1588,N_1973);
xnor U3014 (N_3014,N_2430,N_1990);
and U3015 (N_3015,N_2770,N_1875);
or U3016 (N_3016,N_1613,N_1893);
nand U3017 (N_3017,N_2176,N_2782);
or U3018 (N_3018,N_2352,N_2621);
nor U3019 (N_3019,N_2653,N_2660);
or U3020 (N_3020,N_1967,N_2802);
and U3021 (N_3021,N_2741,N_2269);
or U3022 (N_3022,N_2504,N_2299);
and U3023 (N_3023,N_2722,N_2168);
nor U3024 (N_3024,N_2951,N_1845);
nor U3025 (N_3025,N_2090,N_1528);
or U3026 (N_3026,N_2105,N_1558);
or U3027 (N_3027,N_2809,N_2727);
nand U3028 (N_3028,N_2272,N_1885);
nand U3029 (N_3029,N_2723,N_2393);
or U3030 (N_3030,N_1906,N_1589);
nand U3031 (N_3031,N_1810,N_2923);
xnor U3032 (N_3032,N_2816,N_2557);
nor U3033 (N_3033,N_2591,N_1646);
or U3034 (N_3034,N_2749,N_2926);
or U3035 (N_3035,N_2359,N_1880);
xor U3036 (N_3036,N_2232,N_1859);
nor U3037 (N_3037,N_2719,N_1624);
nand U3038 (N_3038,N_1826,N_1732);
xor U3039 (N_3039,N_2988,N_1566);
and U3040 (N_3040,N_2262,N_2881);
xor U3041 (N_3041,N_2473,N_2127);
or U3042 (N_3042,N_2395,N_1809);
and U3043 (N_3043,N_2935,N_2250);
nand U3044 (N_3044,N_2030,N_2706);
xor U3045 (N_3045,N_2418,N_2149);
nor U3046 (N_3046,N_1954,N_2990);
or U3047 (N_3047,N_2670,N_2293);
and U3048 (N_3048,N_2938,N_2537);
or U3049 (N_3049,N_2494,N_2140);
nor U3050 (N_3050,N_2053,N_2549);
xor U3051 (N_3051,N_1746,N_2804);
or U3052 (N_3052,N_2562,N_1656);
nor U3053 (N_3053,N_2139,N_2071);
nand U3054 (N_3054,N_2474,N_1903);
nor U3055 (N_3055,N_1742,N_2110);
xnor U3056 (N_3056,N_2983,N_2882);
xnor U3057 (N_3057,N_2225,N_2278);
or U3058 (N_3058,N_2162,N_2350);
xor U3059 (N_3059,N_2484,N_2689);
or U3060 (N_3060,N_2470,N_2080);
nand U3061 (N_3061,N_1657,N_1953);
nand U3062 (N_3062,N_2378,N_1592);
xor U3063 (N_3063,N_2345,N_2211);
nor U3064 (N_3064,N_2476,N_2825);
nand U3065 (N_3065,N_2880,N_2589);
or U3066 (N_3066,N_2478,N_2076);
nor U3067 (N_3067,N_2398,N_1808);
and U3068 (N_3068,N_2808,N_2593);
nand U3069 (N_3069,N_1543,N_2752);
and U3070 (N_3070,N_2865,N_2326);
nor U3071 (N_3071,N_1920,N_2666);
nor U3072 (N_3072,N_1756,N_1806);
and U3073 (N_3073,N_2776,N_1676);
or U3074 (N_3074,N_2353,N_1971);
xnor U3075 (N_3075,N_1787,N_2203);
nor U3076 (N_3076,N_1928,N_2347);
nand U3077 (N_3077,N_2948,N_1521);
nor U3078 (N_3078,N_2313,N_2129);
xor U3079 (N_3079,N_2910,N_1700);
nor U3080 (N_3080,N_1868,N_1598);
and U3081 (N_3081,N_2718,N_2681);
and U3082 (N_3082,N_2916,N_2863);
xor U3083 (N_3083,N_2142,N_2257);
nand U3084 (N_3084,N_2114,N_1927);
and U3085 (N_3085,N_2223,N_2254);
nand U3086 (N_3086,N_1759,N_1877);
and U3087 (N_3087,N_2416,N_2103);
or U3088 (N_3088,N_1510,N_1852);
or U3089 (N_3089,N_2156,N_1718);
xnor U3090 (N_3090,N_2289,N_2137);
nand U3091 (N_3091,N_2824,N_1502);
nor U3092 (N_3092,N_2958,N_1721);
or U3093 (N_3093,N_1937,N_2177);
and U3094 (N_3094,N_1949,N_2100);
or U3095 (N_3095,N_2524,N_2305);
nor U3096 (N_3096,N_2338,N_2304);
nor U3097 (N_3097,N_1863,N_2902);
xor U3098 (N_3098,N_1628,N_1523);
nand U3099 (N_3099,N_1586,N_2942);
xor U3100 (N_3100,N_1899,N_2402);
nand U3101 (N_3101,N_2095,N_2753);
nor U3102 (N_3102,N_2744,N_2956);
and U3103 (N_3103,N_2799,N_2945);
and U3104 (N_3104,N_2355,N_2357);
or U3105 (N_3105,N_2033,N_2607);
and U3106 (N_3106,N_2029,N_2303);
xnor U3107 (N_3107,N_2754,N_1668);
or U3108 (N_3108,N_1615,N_1948);
nor U3109 (N_3109,N_1614,N_2592);
xor U3110 (N_3110,N_2739,N_1664);
or U3111 (N_3111,N_2349,N_2993);
or U3112 (N_3112,N_2221,N_2091);
nor U3113 (N_3113,N_2427,N_2797);
xor U3114 (N_3114,N_2116,N_1602);
nor U3115 (N_3115,N_1620,N_1595);
xnor U3116 (N_3116,N_1618,N_2406);
nor U3117 (N_3117,N_2443,N_2964);
or U3118 (N_3118,N_2939,N_2889);
and U3119 (N_3119,N_2331,N_2067);
nand U3120 (N_3120,N_2113,N_2404);
nor U3121 (N_3121,N_1784,N_2256);
and U3122 (N_3122,N_2519,N_1715);
nand U3123 (N_3123,N_1508,N_2639);
xor U3124 (N_3124,N_2083,N_1716);
and U3125 (N_3125,N_2185,N_2437);
or U3126 (N_3126,N_2323,N_2320);
nor U3127 (N_3127,N_2758,N_2195);
xor U3128 (N_3128,N_1751,N_2944);
or U3129 (N_3129,N_2201,N_2700);
and U3130 (N_3130,N_2013,N_2714);
nand U3131 (N_3131,N_2340,N_2815);
nor U3132 (N_3132,N_1736,N_1524);
or U3133 (N_3133,N_2965,N_2943);
nand U3134 (N_3134,N_2370,N_2104);
nor U3135 (N_3135,N_2775,N_2844);
xnor U3136 (N_3136,N_1594,N_2521);
or U3137 (N_3137,N_2602,N_2847);
and U3138 (N_3138,N_2493,N_2704);
nor U3139 (N_3139,N_2175,N_2001);
nand U3140 (N_3140,N_2963,N_2241);
or U3141 (N_3141,N_2567,N_2438);
and U3142 (N_3142,N_2573,N_1515);
xor U3143 (N_3143,N_2544,N_2895);
nor U3144 (N_3144,N_2330,N_2052);
nand U3145 (N_3145,N_1617,N_1634);
nand U3146 (N_3146,N_1856,N_1557);
and U3147 (N_3147,N_1998,N_2624);
or U3148 (N_3148,N_1507,N_1912);
and U3149 (N_3149,N_2594,N_1822);
nand U3150 (N_3150,N_2862,N_2920);
nor U3151 (N_3151,N_2094,N_1532);
and U3152 (N_3152,N_2346,N_2003);
nand U3153 (N_3153,N_1853,N_1832);
and U3154 (N_3154,N_1977,N_2295);
xnor U3155 (N_3155,N_2580,N_2483);
and U3156 (N_3156,N_2248,N_1857);
or U3157 (N_3157,N_2255,N_2328);
nand U3158 (N_3158,N_1807,N_2198);
or U3159 (N_3159,N_2335,N_1693);
and U3160 (N_3160,N_1834,N_2343);
nand U3161 (N_3161,N_2364,N_2062);
nand U3162 (N_3162,N_2267,N_2673);
and U3163 (N_3163,N_2501,N_1750);
xor U3164 (N_3164,N_2538,N_2850);
nor U3165 (N_3165,N_1930,N_2227);
nor U3166 (N_3166,N_1780,N_2854);
nor U3167 (N_3167,N_1606,N_2022);
nand U3168 (N_3168,N_2024,N_2411);
or U3169 (N_3169,N_2431,N_2191);
and U3170 (N_3170,N_2906,N_2342);
xnor U3171 (N_3171,N_1839,N_2477);
nand U3172 (N_3172,N_2747,N_1995);
nand U3173 (N_3173,N_1737,N_2821);
xnor U3174 (N_3174,N_2587,N_1632);
xor U3175 (N_3175,N_1915,N_2870);
and U3176 (N_3176,N_2585,N_2774);
or U3177 (N_3177,N_2822,N_2365);
xor U3178 (N_3178,N_2459,N_2239);
and U3179 (N_3179,N_2977,N_1659);
nand U3180 (N_3180,N_2698,N_1804);
or U3181 (N_3181,N_2678,N_2000);
xnor U3182 (N_3182,N_2309,N_1590);
and U3183 (N_3183,N_2968,N_1797);
nor U3184 (N_3184,N_2655,N_2894);
and U3185 (N_3185,N_1637,N_1962);
xor U3186 (N_3186,N_2447,N_1886);
or U3187 (N_3187,N_2111,N_1651);
nor U3188 (N_3188,N_2980,N_1752);
nand U3189 (N_3189,N_2469,N_1582);
or U3190 (N_3190,N_1772,N_2550);
nand U3191 (N_3191,N_1887,N_2696);
xor U3192 (N_3192,N_1824,N_2075);
nand U3193 (N_3193,N_2017,N_2710);
nor U3194 (N_3194,N_2962,N_1647);
or U3195 (N_3195,N_1505,N_1520);
and U3196 (N_3196,N_2055,N_2658);
xnor U3197 (N_3197,N_1766,N_2121);
xnor U3198 (N_3198,N_2339,N_2569);
and U3199 (N_3199,N_2401,N_2745);
xor U3200 (N_3200,N_2291,N_2011);
nand U3201 (N_3201,N_1621,N_1879);
nand U3202 (N_3202,N_2066,N_2311);
and U3203 (N_3203,N_2633,N_2197);
nor U3204 (N_3204,N_2675,N_2765);
xnor U3205 (N_3205,N_1814,N_1623);
and U3206 (N_3206,N_1770,N_1849);
nand U3207 (N_3207,N_1561,N_2818);
or U3208 (N_3208,N_1734,N_1890);
or U3209 (N_3209,N_2726,N_2925);
or U3210 (N_3210,N_2007,N_2301);
nand U3211 (N_3211,N_2510,N_1677);
xnor U3212 (N_3212,N_1866,N_2764);
xnor U3213 (N_3213,N_2167,N_2834);
and U3214 (N_3214,N_2146,N_2540);
nand U3215 (N_3215,N_2648,N_1909);
nand U3216 (N_3216,N_2037,N_1688);
or U3217 (N_3217,N_2623,N_2183);
nand U3218 (N_3218,N_2118,N_2772);
nor U3219 (N_3219,N_2579,N_2612);
nand U3220 (N_3220,N_2181,N_2957);
nor U3221 (N_3221,N_2165,N_2814);
and U3222 (N_3222,N_2435,N_2192);
and U3223 (N_3223,N_2173,N_2885);
nand U3224 (N_3224,N_1947,N_2611);
xnor U3225 (N_3225,N_2020,N_2207);
and U3226 (N_3226,N_2101,N_2408);
xor U3227 (N_3227,N_2606,N_1921);
or U3228 (N_3228,N_2903,N_2832);
and U3229 (N_3229,N_1739,N_2518);
nor U3230 (N_3230,N_2683,N_2652);
nor U3231 (N_3231,N_1506,N_1980);
nor U3232 (N_3232,N_2271,N_2836);
xor U3233 (N_3233,N_2457,N_1919);
nor U3234 (N_3234,N_2279,N_1769);
nor U3235 (N_3235,N_2087,N_2608);
nor U3236 (N_3236,N_1754,N_1638);
nor U3237 (N_3237,N_2755,N_2733);
nor U3238 (N_3238,N_1554,N_2190);
nor U3239 (N_3239,N_2781,N_2725);
xnor U3240 (N_3240,N_2096,N_2552);
nor U3241 (N_3241,N_2038,N_2405);
nand U3242 (N_3242,N_2124,N_1673);
or U3243 (N_3243,N_1691,N_2574);
or U3244 (N_3244,N_1905,N_1897);
or U3245 (N_3245,N_2872,N_1976);
and U3246 (N_3246,N_1926,N_1705);
nor U3247 (N_3247,N_2498,N_2548);
xnor U3248 (N_3248,N_1710,N_1744);
nor U3249 (N_3249,N_2514,N_2229);
xor U3250 (N_3250,N_2006,N_2833);
nand U3251 (N_3251,N_1816,N_1760);
nor U3252 (N_3252,N_2245,N_2523);
nor U3253 (N_3253,N_2731,N_2936);
nand U3254 (N_3254,N_2997,N_1933);
nand U3255 (N_3255,N_2025,N_2724);
xor U3256 (N_3256,N_2171,N_2905);
xnor U3257 (N_3257,N_2702,N_1891);
and U3258 (N_3258,N_2187,N_2688);
nor U3259 (N_3259,N_2041,N_1901);
nand U3260 (N_3260,N_1560,N_2322);
or U3261 (N_3261,N_2701,N_1828);
and U3262 (N_3262,N_1763,N_2866);
and U3263 (N_3263,N_1610,N_2072);
nor U3264 (N_3264,N_2166,N_1993);
or U3265 (N_3265,N_1596,N_1530);
or U3266 (N_3266,N_2684,N_2327);
nor U3267 (N_3267,N_2974,N_1813);
nor U3268 (N_3268,N_1840,N_1740);
xnor U3269 (N_3269,N_2588,N_2302);
xor U3270 (N_3270,N_2287,N_1955);
or U3271 (N_3271,N_2216,N_2419);
and U3272 (N_3272,N_2125,N_2270);
and U3273 (N_3273,N_2039,N_2873);
or U3274 (N_3274,N_2975,N_1916);
xor U3275 (N_3275,N_1535,N_2784);
nand U3276 (N_3276,N_1685,N_1861);
or U3277 (N_3277,N_1981,N_1517);
or U3278 (N_3278,N_1513,N_2377);
or U3279 (N_3279,N_2317,N_1932);
nor U3280 (N_3280,N_2012,N_2490);
nand U3281 (N_3281,N_1717,N_1593);
nor U3282 (N_3282,N_1819,N_2202);
nor U3283 (N_3283,N_2065,N_2174);
xnor U3284 (N_3284,N_2917,N_2264);
nand U3285 (N_3285,N_1712,N_1603);
and U3286 (N_3286,N_2792,N_2662);
nor U3287 (N_3287,N_1665,N_2230);
or U3288 (N_3288,N_1662,N_2237);
and U3289 (N_3289,N_2439,N_1686);
and U3290 (N_3290,N_2650,N_2554);
xor U3291 (N_3291,N_2735,N_1925);
or U3292 (N_3292,N_2045,N_2078);
nand U3293 (N_3293,N_2511,N_2283);
or U3294 (N_3294,N_1585,N_2583);
and U3295 (N_3295,N_2034,N_2458);
or U3296 (N_3296,N_2984,N_1512);
or U3297 (N_3297,N_2839,N_1934);
or U3298 (N_3298,N_1648,N_1556);
nor U3299 (N_3299,N_2002,N_2609);
nand U3300 (N_3300,N_2743,N_2867);
and U3301 (N_3301,N_2795,N_2596);
nor U3302 (N_3302,N_1616,N_2778);
and U3303 (N_3303,N_2426,N_2144);
xnor U3304 (N_3304,N_1959,N_1773);
and U3305 (N_3305,N_2275,N_2021);
nor U3306 (N_3306,N_1550,N_2366);
and U3307 (N_3307,N_2687,N_2961);
or U3308 (N_3308,N_2848,N_2481);
and U3309 (N_3309,N_1791,N_1907);
nor U3310 (N_3310,N_2647,N_1789);
and U3311 (N_3311,N_2097,N_2172);
nor U3312 (N_3312,N_1539,N_2803);
and U3313 (N_3313,N_1992,N_1501);
xor U3314 (N_3314,N_1581,N_2300);
xor U3315 (N_3315,N_2638,N_1842);
nor U3316 (N_3316,N_1644,N_2157);
or U3317 (N_3317,N_2534,N_1549);
nand U3318 (N_3318,N_1864,N_1869);
nand U3319 (N_3319,N_2058,N_2088);
or U3320 (N_3320,N_2454,N_2659);
nand U3321 (N_3321,N_2649,N_2424);
or U3322 (N_3322,N_2170,N_2615);
or U3323 (N_3323,N_1938,N_2893);
nand U3324 (N_3324,N_1533,N_1619);
nand U3325 (N_3325,N_2251,N_2188);
and U3326 (N_3326,N_2535,N_2069);
or U3327 (N_3327,N_2692,N_2464);
xnor U3328 (N_3328,N_1972,N_2933);
xor U3329 (N_3329,N_2515,N_2486);
or U3330 (N_3330,N_2861,N_2635);
or U3331 (N_3331,N_2420,N_2122);
nor U3332 (N_3332,N_2841,N_2496);
or U3333 (N_3333,N_1838,N_1748);
nor U3334 (N_3334,N_2160,N_2138);
xnor U3335 (N_3335,N_1706,N_2399);
xnor U3336 (N_3336,N_2838,N_2009);
xor U3337 (N_3337,N_2441,N_1675);
xnor U3338 (N_3338,N_1851,N_2886);
and U3339 (N_3339,N_2645,N_2801);
and U3340 (N_3340,N_1548,N_1687);
nand U3341 (N_3341,N_2147,N_1889);
or U3342 (N_3342,N_2789,N_2373);
xnor U3343 (N_3343,N_2228,N_2713);
and U3344 (N_3344,N_2085,N_1542);
xor U3345 (N_3345,N_1743,N_1629);
and U3346 (N_3346,N_2634,N_2102);
and U3347 (N_3347,N_1611,N_2915);
nor U3348 (N_3348,N_2890,N_2828);
nor U3349 (N_3349,N_2924,N_2333);
nand U3350 (N_3350,N_2899,N_2605);
nand U3351 (N_3351,N_1666,N_1697);
xor U3352 (N_3352,N_1771,N_2699);
or U3353 (N_3353,N_2290,N_1654);
and U3354 (N_3354,N_1783,N_2855);
xor U3355 (N_3355,N_1956,N_2392);
xnor U3356 (N_3356,N_1626,N_2051);
and U3357 (N_3357,N_2463,N_1573);
and U3358 (N_3358,N_2159,N_1534);
xnor U3359 (N_3359,N_1935,N_2860);
and U3360 (N_3360,N_1764,N_2978);
nor U3361 (N_3361,N_1892,N_1862);
nor U3362 (N_3362,N_1942,N_2059);
nand U3363 (N_3363,N_2921,N_2258);
nor U3364 (N_3364,N_2604,N_2131);
nor U3365 (N_3365,N_2244,N_2864);
xnor U3366 (N_3366,N_1702,N_2497);
xnor U3367 (N_3367,N_1896,N_2672);
xnor U3368 (N_3368,N_1741,N_1690);
xor U3369 (N_3369,N_2637,N_2887);
or U3370 (N_3370,N_2152,N_1984);
xor U3371 (N_3371,N_2220,N_2716);
or U3372 (N_3372,N_2048,N_1714);
or U3373 (N_3373,N_1733,N_1562);
nand U3374 (N_3374,N_1786,N_2161);
nand U3375 (N_3375,N_1985,N_1960);
nand U3376 (N_3376,N_2372,N_2449);
nand U3377 (N_3377,N_2491,N_2217);
nand U3378 (N_3378,N_2243,N_2737);
and U3379 (N_3379,N_2891,N_2686);
xor U3380 (N_3380,N_2868,N_2112);
nand U3381 (N_3381,N_2665,N_1570);
xnor U3382 (N_3382,N_2888,N_2465);
nand U3383 (N_3383,N_2721,N_1782);
or U3384 (N_3384,N_2163,N_2005);
and U3385 (N_3385,N_1636,N_1979);
xnor U3386 (N_3386,N_1608,N_2249);
nor U3387 (N_3387,N_2617,N_2570);
nor U3388 (N_3388,N_2259,N_2614);
and U3389 (N_3389,N_2448,N_1527);
xor U3390 (N_3390,N_1767,N_2896);
nor U3391 (N_3391,N_2132,N_2467);
and U3392 (N_3392,N_2382,N_2334);
xor U3393 (N_3393,N_2641,N_2031);
or U3394 (N_3394,N_2601,N_1674);
or U3395 (N_3395,N_2189,N_2734);
and U3396 (N_3396,N_2576,N_2233);
nor U3397 (N_3397,N_2883,N_1873);
and U3398 (N_3398,N_2929,N_2695);
xor U3399 (N_3399,N_1547,N_1607);
or U3400 (N_3400,N_2973,N_2450);
nor U3401 (N_3401,N_2536,N_2664);
xnor U3402 (N_3402,N_2572,N_2158);
xnor U3403 (N_3403,N_2940,N_2509);
nand U3404 (N_3404,N_2907,N_2911);
nor U3405 (N_3405,N_1761,N_1643);
xor U3406 (N_3406,N_2779,N_2679);
xnor U3407 (N_3407,N_1639,N_2996);
nand U3408 (N_3408,N_1757,N_2503);
or U3409 (N_3409,N_1874,N_2771);
nand U3410 (N_3410,N_2199,N_2361);
nand U3411 (N_3411,N_2433,N_2643);
nand U3412 (N_3412,N_2380,N_1694);
or U3413 (N_3413,N_1671,N_1579);
xor U3414 (N_3414,N_1878,N_2810);
nor U3415 (N_3415,N_1945,N_2215);
nand U3416 (N_3416,N_2277,N_1961);
and U3417 (N_3417,N_2584,N_2506);
nand U3418 (N_3418,N_1574,N_2522);
nand U3419 (N_3419,N_2315,N_1625);
xor U3420 (N_3420,N_2742,N_2991);
nand U3421 (N_3421,N_2120,N_1831);
nand U3422 (N_3422,N_1726,N_1762);
nor U3423 (N_3423,N_2208,N_2064);
xor U3424 (N_3424,N_1951,N_2667);
xor U3425 (N_3425,N_2026,N_2798);
nor U3426 (N_3426,N_2879,N_2164);
nor U3427 (N_3427,N_2297,N_1821);
or U3428 (N_3428,N_2151,N_2812);
xnor U3429 (N_3429,N_2108,N_2590);
and U3430 (N_3430,N_2423,N_1720);
nand U3431 (N_3431,N_2581,N_1865);
nand U3432 (N_3432,N_1701,N_2180);
and U3433 (N_3433,N_2757,N_1536);
or U3434 (N_3434,N_1964,N_2321);
nand U3435 (N_3435,N_1792,N_1898);
nand U3436 (N_3436,N_1836,N_2876);
nand U3437 (N_3437,N_1738,N_2479);
and U3438 (N_3438,N_2184,N_1569);
nor U3439 (N_3439,N_1698,N_2089);
nand U3440 (N_3440,N_1709,N_1679);
and U3441 (N_3441,N_2010,N_1825);
nand U3442 (N_3442,N_2403,N_1703);
or U3443 (N_3443,N_2783,N_2843);
or U3444 (N_3444,N_1966,N_2738);
xor U3445 (N_3445,N_1655,N_2913);
nor U3446 (N_3446,N_1699,N_2830);
nor U3447 (N_3447,N_1724,N_2777);
or U3448 (N_3448,N_2488,N_2851);
nand U3449 (N_3449,N_2288,N_1994);
and U3450 (N_3450,N_2856,N_2566);
nor U3451 (N_3451,N_2414,N_1794);
or U3452 (N_3452,N_2050,N_2561);
nand U3453 (N_3453,N_2709,N_2028);
and U3454 (N_3454,N_2282,N_2119);
or U3455 (N_3455,N_2989,N_1775);
nor U3456 (N_3456,N_2610,N_2934);
nor U3457 (N_3457,N_1572,N_2205);
nor U3458 (N_3458,N_1601,N_1847);
and U3459 (N_3459,N_2912,N_2691);
and U3460 (N_3460,N_2356,N_1729);
nand U3461 (N_3461,N_1684,N_2852);
nand U3462 (N_3462,N_2413,N_1727);
xnor U3463 (N_3463,N_2853,N_1516);
nand U3464 (N_3464,N_2532,N_2200);
and U3465 (N_3465,N_1803,N_1630);
xor U3466 (N_3466,N_1917,N_2715);
nand U3467 (N_3467,N_2976,N_2461);
or U3468 (N_3468,N_2133,N_2790);
or U3469 (N_3469,N_2128,N_1895);
or U3470 (N_3470,N_2730,N_2794);
and U3471 (N_3471,N_2807,N_2375);
nor U3472 (N_3472,N_2539,N_1541);
or U3473 (N_3473,N_2407,N_2597);
or U3474 (N_3474,N_2242,N_2533);
and U3475 (N_3475,N_1996,N_2421);
nor U3476 (N_3476,N_2004,N_2348);
or U3477 (N_3477,N_2344,N_2871);
or U3478 (N_3478,N_2070,N_2316);
xnor U3479 (N_3479,N_1511,N_2694);
and U3480 (N_3480,N_1612,N_2008);
xor U3481 (N_3481,N_2791,N_2294);
or U3482 (N_3482,N_2369,N_1661);
or U3483 (N_3483,N_2657,N_2489);
and U3484 (N_3484,N_1820,N_2693);
and U3485 (N_3485,N_1719,N_2376);
and U3486 (N_3486,N_2671,N_2663);
or U3487 (N_3487,N_2261,N_2044);
xor U3488 (N_3488,N_2466,N_2236);
and U3489 (N_3489,N_1583,N_2932);
nand U3490 (N_3490,N_1777,N_1914);
or U3491 (N_3491,N_1753,N_2750);
and U3492 (N_3492,N_2226,N_2760);
nor U3493 (N_3493,N_2502,N_2214);
nand U3494 (N_3494,N_2046,N_2240);
xor U3495 (N_3495,N_2531,N_1871);
or U3496 (N_3496,N_2434,N_2768);
and U3497 (N_3497,N_2525,N_2520);
xor U3498 (N_3498,N_2042,N_2273);
nand U3499 (N_3499,N_2941,N_2442);
and U3500 (N_3500,N_2528,N_2135);
nor U3501 (N_3501,N_2577,N_2884);
and U3502 (N_3502,N_2685,N_2047);
and U3503 (N_3503,N_1894,N_2019);
and U3504 (N_3504,N_2630,N_1567);
and U3505 (N_3505,N_1640,N_2512);
xnor U3506 (N_3506,N_1982,N_1503);
or U3507 (N_3507,N_1627,N_2985);
or U3508 (N_3508,N_1778,N_2756);
nor U3509 (N_3509,N_2500,N_2440);
xor U3510 (N_3510,N_1747,N_2769);
nor U3511 (N_3511,N_2613,N_1844);
nand U3512 (N_3512,N_2224,N_2616);
or U3513 (N_3513,N_2953,N_2736);
xor U3514 (N_3514,N_2391,N_1815);
or U3515 (N_3515,N_2842,N_1600);
and U3516 (N_3516,N_1835,N_2073);
nand U3517 (N_3517,N_2559,N_2231);
and U3518 (N_3518,N_2386,N_2858);
nor U3519 (N_3519,N_1900,N_1811);
or U3520 (N_3520,N_2556,N_2460);
nand U3521 (N_3521,N_1848,N_1571);
nor U3522 (N_3522,N_1649,N_1631);
xnor U3523 (N_3523,N_2206,N_2805);
and U3524 (N_3524,N_1837,N_2829);
or U3525 (N_3525,N_2705,N_2636);
xor U3526 (N_3526,N_2456,N_2444);
or U3527 (N_3527,N_1983,N_2919);
nor U3528 (N_3528,N_1663,N_2981);
and U3529 (N_3529,N_2526,N_1683);
and U3530 (N_3530,N_2586,N_2603);
nor U3531 (N_3531,N_2928,N_2385);
and U3532 (N_3532,N_2482,N_1704);
xnor U3533 (N_3533,N_2253,N_1946);
nand U3534 (N_3534,N_1923,N_2690);
or U3535 (N_3535,N_2874,N_2196);
or U3536 (N_3536,N_2222,N_2453);
and U3537 (N_3537,N_2547,N_1989);
nand U3538 (N_3538,N_2578,N_2931);
and U3539 (N_3539,N_1696,N_2274);
or U3540 (N_3540,N_2595,N_2788);
or U3541 (N_3541,N_2543,N_2558);
and U3542 (N_3542,N_2027,N_2955);
xnor U3543 (N_3543,N_2468,N_2134);
nor U3544 (N_3544,N_2043,N_2529);
and U3545 (N_3545,N_1812,N_2987);
nand U3546 (N_3546,N_2499,N_2318);
or U3547 (N_3547,N_1584,N_2759);
and U3548 (N_3548,N_1918,N_2415);
or U3549 (N_3549,N_2703,N_2565);
or U3550 (N_3550,N_2074,N_1910);
xnor U3551 (N_3551,N_1860,N_2296);
xor U3552 (N_3552,N_2626,N_1924);
xor U3553 (N_3553,N_1870,N_1531);
and U3554 (N_3554,N_2740,N_1944);
nor U3555 (N_3555,N_2628,N_2827);
or U3556 (N_3556,N_1670,N_2485);
nor U3557 (N_3557,N_2209,N_2117);
or U3558 (N_3558,N_2126,N_2819);
and U3559 (N_3559,N_2831,N_2629);
or U3560 (N_3560,N_2651,N_2717);
or U3561 (N_3561,N_2285,N_2036);
or U3562 (N_3562,N_2452,N_2900);
or U3563 (N_3563,N_1538,N_2281);
and U3564 (N_3564,N_1604,N_2451);
nand U3565 (N_3565,N_2268,N_2390);
nand U3566 (N_3566,N_1781,N_1817);
xnor U3567 (N_3567,N_2674,N_2517);
and U3568 (N_3568,N_1708,N_2697);
or U3569 (N_3569,N_1963,N_2436);
nor U3570 (N_3570,N_2213,N_1597);
xor U3571 (N_3571,N_1519,N_2284);
nand U3572 (N_3572,N_1940,N_2235);
nand U3573 (N_3573,N_1970,N_2796);
nor U3574 (N_3574,N_1795,N_1500);
and U3575 (N_3575,N_2516,N_2182);
and U3576 (N_3576,N_1974,N_2625);
nor U3577 (N_3577,N_2212,N_1678);
or U3578 (N_3578,N_1881,N_2109);
xor U3579 (N_3579,N_1986,N_2711);
nand U3580 (N_3580,N_2492,N_2194);
nor U3581 (N_3581,N_1591,N_2969);
xor U3582 (N_3582,N_1568,N_2063);
or U3583 (N_3583,N_1559,N_1575);
or U3584 (N_3584,N_2568,N_2992);
or U3585 (N_3585,N_2542,N_2787);
and U3586 (N_3586,N_1850,N_2904);
xor U3587 (N_3587,N_2324,N_1526);
xor U3588 (N_3588,N_1941,N_2507);
or U3589 (N_3589,N_2319,N_2582);
xor U3590 (N_3590,N_2952,N_1855);
nor U3591 (N_3591,N_2763,N_1858);
or U3592 (N_3592,N_2336,N_2817);
nor U3593 (N_3593,N_2153,N_1776);
nor U3594 (N_3594,N_1689,N_1969);
and U3595 (N_3595,N_2632,N_2898);
and U3596 (N_3596,N_1802,N_1902);
xnor U3597 (N_3597,N_2555,N_2115);
or U3598 (N_3598,N_2937,N_2677);
nor U3599 (N_3599,N_2054,N_1798);
nor U3600 (N_3600,N_2927,N_2668);
nor U3601 (N_3601,N_1553,N_2247);
or U3602 (N_3602,N_1735,N_2098);
or U3603 (N_3603,N_2766,N_1599);
nand U3604 (N_3604,N_2079,N_2656);
nor U3605 (N_3605,N_2947,N_1707);
xor U3606 (N_3606,N_2762,N_1805);
nand U3607 (N_3607,N_2306,N_2367);
nand U3608 (N_3608,N_1580,N_2186);
or U3609 (N_3609,N_2471,N_1987);
and U3610 (N_3610,N_2362,N_1823);
nand U3611 (N_3611,N_1672,N_1830);
nand U3612 (N_3612,N_2619,N_1667);
xor U3613 (N_3613,N_2307,N_2148);
nor U3614 (N_3614,N_2384,N_1692);
xnor U3615 (N_3615,N_1943,N_2238);
xor U3616 (N_3616,N_2918,N_1801);
xor U3617 (N_3617,N_2445,N_1843);
nand U3618 (N_3618,N_1833,N_2820);
nand U3619 (N_3619,N_1779,N_2354);
nor U3620 (N_3620,N_2806,N_2374);
nor U3621 (N_3621,N_1537,N_2150);
or U3622 (N_3622,N_2960,N_1988);
xnor U3623 (N_3623,N_2892,N_2560);
nand U3624 (N_3624,N_2040,N_1564);
xnor U3625 (N_3625,N_2371,N_2332);
xor U3626 (N_3626,N_1711,N_2732);
nor U3627 (N_3627,N_2575,N_2835);
nor U3628 (N_3628,N_2751,N_2994);
nand U3629 (N_3629,N_2914,N_1968);
and U3630 (N_3630,N_1514,N_1587);
or U3631 (N_3631,N_2314,N_2553);
and U3632 (N_3632,N_1997,N_1578);
nor U3633 (N_3633,N_2358,N_2622);
and U3634 (N_3634,N_2967,N_1867);
or U3635 (N_3635,N_2640,N_2204);
or U3636 (N_3636,N_2508,N_2475);
or U3637 (N_3637,N_2971,N_1540);
or U3638 (N_3638,N_2368,N_1854);
xnor U3639 (N_3639,N_2959,N_1827);
and U3640 (N_3640,N_1758,N_2785);
nor U3641 (N_3641,N_2310,N_2455);
or U3642 (N_3642,N_2530,N_2495);
nor U3643 (N_3643,N_2379,N_2056);
or U3644 (N_3644,N_1609,N_2712);
and U3645 (N_3645,N_2618,N_1745);
and U3646 (N_3646,N_2136,N_1952);
nor U3647 (N_3647,N_1950,N_2014);
nor U3648 (N_3648,N_2545,N_1846);
nor U3649 (N_3649,N_2060,N_2018);
xnor U3650 (N_3650,N_1911,N_2145);
xor U3651 (N_3651,N_1723,N_1904);
xnor U3652 (N_3652,N_2986,N_1722);
nand U3653 (N_3653,N_2388,N_2826);
or U3654 (N_3654,N_2859,N_1922);
and U3655 (N_3655,N_2092,N_2954);
nand U3656 (N_3656,N_1883,N_1633);
xor U3657 (N_3657,N_2979,N_2748);
nand U3658 (N_3658,N_1713,N_2341);
xor U3659 (N_3659,N_2193,N_1658);
nor U3660 (N_3660,N_1642,N_2446);
nor U3661 (N_3661,N_1957,N_2527);
nand U3662 (N_3662,N_1525,N_2077);
nor U3663 (N_3663,N_2154,N_2082);
nor U3664 (N_3664,N_2840,N_2875);
nor U3665 (N_3665,N_2234,N_1888);
xor U3666 (N_3666,N_2396,N_2337);
or U3667 (N_3667,N_2720,N_2901);
xor U3668 (N_3668,N_2541,N_2972);
xor U3669 (N_3669,N_2462,N_1650);
or U3670 (N_3670,N_1653,N_2381);
xor U3671 (N_3671,N_1522,N_1800);
nor U3672 (N_3672,N_2908,N_1965);
xor U3673 (N_3673,N_2746,N_2930);
and U3674 (N_3674,N_2432,N_2627);
and U3675 (N_3675,N_2016,N_2246);
nor U3676 (N_3676,N_1765,N_2400);
nand U3677 (N_3677,N_2394,N_2086);
nor U3678 (N_3678,N_2422,N_1682);
nor U3679 (N_3679,N_1552,N_2546);
nor U3680 (N_3680,N_2780,N_2729);
and U3681 (N_3681,N_2298,N_1622);
nand U3682 (N_3682,N_1509,N_2429);
and U3683 (N_3683,N_1908,N_1931);
xor U3684 (N_3684,N_2260,N_2998);
and U3685 (N_3685,N_2682,N_1565);
and U3686 (N_3686,N_1796,N_1551);
xor U3687 (N_3687,N_2312,N_2107);
nor U3688 (N_3688,N_2178,N_2563);
nor U3689 (N_3689,N_2106,N_2049);
xor U3690 (N_3690,N_2571,N_1774);
xnor U3691 (N_3691,N_1768,N_1669);
xor U3692 (N_3692,N_2428,N_1818);
or U3693 (N_3693,N_1681,N_2813);
or U3694 (N_3694,N_2793,N_1793);
and U3695 (N_3695,N_1695,N_2425);
xnor U3696 (N_3696,N_1544,N_1829);
nand U3697 (N_3697,N_2410,N_2032);
or U3698 (N_3698,N_2099,N_2123);
nor U3699 (N_3699,N_2480,N_2487);
or U3700 (N_3700,N_2179,N_2869);
or U3701 (N_3701,N_1645,N_2218);
and U3702 (N_3702,N_2551,N_1576);
xor U3703 (N_3703,N_2600,N_2130);
or U3704 (N_3704,N_2786,N_1605);
nand U3705 (N_3705,N_1785,N_2707);
and U3706 (N_3706,N_1975,N_2286);
or U3707 (N_3707,N_2598,N_2642);
nor U3708 (N_3708,N_2811,N_2412);
nand U3709 (N_3709,N_2846,N_2773);
and U3710 (N_3710,N_2849,N_2564);
nor U3711 (N_3711,N_1641,N_2389);
nor U3712 (N_3712,N_2280,N_2708);
or U3713 (N_3713,N_1504,N_2946);
nand U3714 (N_3714,N_1882,N_1841);
xnor U3715 (N_3715,N_1876,N_2505);
or U3716 (N_3716,N_2068,N_2922);
xor U3717 (N_3717,N_1563,N_2015);
nand U3718 (N_3718,N_2966,N_2767);
or U3719 (N_3719,N_2823,N_2360);
xor U3720 (N_3720,N_2837,N_2308);
nand U3721 (N_3721,N_1731,N_2909);
or U3722 (N_3722,N_2265,N_2084);
or U3723 (N_3723,N_2292,N_2409);
nand U3724 (N_3724,N_2210,N_2169);
nor U3725 (N_3725,N_2845,N_2351);
and U3726 (N_3726,N_2252,N_2654);
or U3727 (N_3727,N_2800,N_2599);
xor U3728 (N_3728,N_2266,N_1999);
xor U3729 (N_3729,N_2472,N_2877);
nand U3730 (N_3730,N_2417,N_2631);
or U3731 (N_3731,N_2680,N_1652);
xnor U3732 (N_3732,N_2155,N_1884);
and U3733 (N_3733,N_2141,N_2661);
nand U3734 (N_3734,N_2263,N_2219);
nor U3735 (N_3735,N_2363,N_2950);
nor U3736 (N_3736,N_1555,N_1635);
and U3737 (N_3737,N_1991,N_1799);
and U3738 (N_3738,N_1546,N_2970);
nand U3739 (N_3739,N_2878,N_1749);
xor U3740 (N_3740,N_2728,N_1577);
or U3741 (N_3741,N_2276,N_1755);
or U3742 (N_3742,N_2325,N_2081);
nor U3743 (N_3743,N_1936,N_1939);
and U3744 (N_3744,N_2949,N_1958);
nand U3745 (N_3745,N_1978,N_2023);
xnor U3746 (N_3746,N_1680,N_1872);
nor U3747 (N_3747,N_2999,N_2143);
nand U3748 (N_3748,N_1725,N_2646);
nand U3749 (N_3749,N_2982,N_1913);
or U3750 (N_3750,N_2533,N_2163);
xor U3751 (N_3751,N_1609,N_2080);
nor U3752 (N_3752,N_1628,N_2671);
xor U3753 (N_3753,N_2008,N_2802);
nor U3754 (N_3754,N_1940,N_1857);
or U3755 (N_3755,N_2841,N_2424);
nand U3756 (N_3756,N_1616,N_2969);
and U3757 (N_3757,N_2609,N_2490);
xor U3758 (N_3758,N_2493,N_2405);
or U3759 (N_3759,N_2235,N_2830);
or U3760 (N_3760,N_1825,N_2978);
nor U3761 (N_3761,N_1867,N_2824);
nor U3762 (N_3762,N_1928,N_1856);
xnor U3763 (N_3763,N_2690,N_2062);
nand U3764 (N_3764,N_2576,N_2251);
and U3765 (N_3765,N_2134,N_2266);
and U3766 (N_3766,N_2702,N_1582);
or U3767 (N_3767,N_2385,N_1694);
nand U3768 (N_3768,N_2820,N_2415);
nor U3769 (N_3769,N_2477,N_2207);
nand U3770 (N_3770,N_2970,N_2198);
and U3771 (N_3771,N_2547,N_2761);
xnor U3772 (N_3772,N_2874,N_2117);
or U3773 (N_3773,N_2539,N_2062);
nor U3774 (N_3774,N_1857,N_2714);
and U3775 (N_3775,N_1956,N_2063);
nor U3776 (N_3776,N_1587,N_2040);
or U3777 (N_3777,N_1875,N_2296);
nor U3778 (N_3778,N_1825,N_2221);
xnor U3779 (N_3779,N_1613,N_2262);
and U3780 (N_3780,N_2547,N_2891);
nand U3781 (N_3781,N_2210,N_1534);
nand U3782 (N_3782,N_1945,N_2133);
nor U3783 (N_3783,N_2153,N_2914);
nand U3784 (N_3784,N_2930,N_2074);
xnor U3785 (N_3785,N_1775,N_1701);
or U3786 (N_3786,N_2128,N_2267);
xnor U3787 (N_3787,N_2403,N_2521);
or U3788 (N_3788,N_2206,N_2903);
or U3789 (N_3789,N_2750,N_2480);
nor U3790 (N_3790,N_2336,N_1689);
nand U3791 (N_3791,N_2733,N_1876);
nor U3792 (N_3792,N_2842,N_1909);
xnor U3793 (N_3793,N_2622,N_1884);
nor U3794 (N_3794,N_1544,N_2947);
nand U3795 (N_3795,N_2080,N_2667);
xor U3796 (N_3796,N_1961,N_2451);
nor U3797 (N_3797,N_2536,N_2932);
xor U3798 (N_3798,N_2574,N_2796);
and U3799 (N_3799,N_1601,N_1606);
and U3800 (N_3800,N_1530,N_2228);
or U3801 (N_3801,N_2829,N_2474);
or U3802 (N_3802,N_2273,N_1772);
nand U3803 (N_3803,N_2777,N_1573);
nand U3804 (N_3804,N_1686,N_1885);
or U3805 (N_3805,N_2013,N_1725);
xnor U3806 (N_3806,N_2078,N_2421);
nand U3807 (N_3807,N_2384,N_1836);
nor U3808 (N_3808,N_2913,N_1621);
nand U3809 (N_3809,N_2400,N_2885);
xnor U3810 (N_3810,N_2237,N_1767);
or U3811 (N_3811,N_1944,N_1540);
and U3812 (N_3812,N_2564,N_1719);
nand U3813 (N_3813,N_2232,N_2697);
or U3814 (N_3814,N_2744,N_2598);
nor U3815 (N_3815,N_2360,N_2276);
nor U3816 (N_3816,N_2226,N_2930);
or U3817 (N_3817,N_1547,N_2105);
nor U3818 (N_3818,N_2743,N_1883);
or U3819 (N_3819,N_2232,N_1768);
nand U3820 (N_3820,N_1898,N_2913);
nor U3821 (N_3821,N_1997,N_2108);
xnor U3822 (N_3822,N_2980,N_2850);
and U3823 (N_3823,N_2402,N_2251);
or U3824 (N_3824,N_1736,N_2374);
nor U3825 (N_3825,N_2898,N_2570);
nand U3826 (N_3826,N_2881,N_1822);
nand U3827 (N_3827,N_2644,N_2382);
nand U3828 (N_3828,N_2031,N_1862);
nor U3829 (N_3829,N_2421,N_1592);
nor U3830 (N_3830,N_2533,N_1777);
and U3831 (N_3831,N_1567,N_1632);
or U3832 (N_3832,N_1590,N_1938);
nor U3833 (N_3833,N_2435,N_2724);
or U3834 (N_3834,N_2143,N_2726);
or U3835 (N_3835,N_2773,N_1829);
xnor U3836 (N_3836,N_2977,N_1818);
and U3837 (N_3837,N_2246,N_2145);
nor U3838 (N_3838,N_2510,N_2475);
and U3839 (N_3839,N_1538,N_2558);
and U3840 (N_3840,N_2937,N_2613);
or U3841 (N_3841,N_2749,N_2849);
and U3842 (N_3842,N_2731,N_2123);
or U3843 (N_3843,N_2189,N_1539);
or U3844 (N_3844,N_2603,N_1842);
nand U3845 (N_3845,N_1863,N_2226);
or U3846 (N_3846,N_1561,N_2950);
nand U3847 (N_3847,N_2715,N_2182);
xnor U3848 (N_3848,N_2729,N_1977);
or U3849 (N_3849,N_2046,N_1850);
or U3850 (N_3850,N_2909,N_2805);
and U3851 (N_3851,N_2877,N_2580);
nor U3852 (N_3852,N_2962,N_1681);
xor U3853 (N_3853,N_1614,N_2369);
xor U3854 (N_3854,N_1595,N_1713);
nand U3855 (N_3855,N_2015,N_1960);
and U3856 (N_3856,N_2146,N_1824);
or U3857 (N_3857,N_2355,N_1656);
or U3858 (N_3858,N_1715,N_2285);
or U3859 (N_3859,N_2910,N_1644);
xnor U3860 (N_3860,N_2165,N_1605);
nor U3861 (N_3861,N_2642,N_2721);
nor U3862 (N_3862,N_1701,N_1965);
nor U3863 (N_3863,N_1573,N_2990);
and U3864 (N_3864,N_2963,N_2165);
xor U3865 (N_3865,N_1909,N_2584);
nor U3866 (N_3866,N_1521,N_2771);
nand U3867 (N_3867,N_2047,N_2061);
or U3868 (N_3868,N_1775,N_2580);
nand U3869 (N_3869,N_1883,N_2783);
nand U3870 (N_3870,N_2671,N_2774);
and U3871 (N_3871,N_2940,N_2435);
nand U3872 (N_3872,N_1768,N_1729);
xor U3873 (N_3873,N_2474,N_2233);
nor U3874 (N_3874,N_2700,N_1542);
and U3875 (N_3875,N_1733,N_2212);
nor U3876 (N_3876,N_2875,N_2516);
nor U3877 (N_3877,N_2835,N_2739);
and U3878 (N_3878,N_2186,N_2450);
xor U3879 (N_3879,N_2091,N_2766);
xnor U3880 (N_3880,N_2596,N_1823);
or U3881 (N_3881,N_1656,N_2610);
nand U3882 (N_3882,N_2581,N_2718);
nand U3883 (N_3883,N_1858,N_1775);
or U3884 (N_3884,N_1557,N_2693);
nor U3885 (N_3885,N_2349,N_1625);
or U3886 (N_3886,N_2993,N_1816);
nor U3887 (N_3887,N_2583,N_2138);
xor U3888 (N_3888,N_2854,N_2821);
xnor U3889 (N_3889,N_2963,N_2687);
or U3890 (N_3890,N_2959,N_2687);
or U3891 (N_3891,N_2718,N_1966);
nand U3892 (N_3892,N_1710,N_2045);
nor U3893 (N_3893,N_2153,N_1857);
nor U3894 (N_3894,N_2340,N_2519);
xor U3895 (N_3895,N_2189,N_2651);
nor U3896 (N_3896,N_1551,N_2062);
nor U3897 (N_3897,N_2396,N_1561);
xor U3898 (N_3898,N_1770,N_2090);
xnor U3899 (N_3899,N_1617,N_2392);
and U3900 (N_3900,N_2284,N_2849);
nor U3901 (N_3901,N_2915,N_2062);
nor U3902 (N_3902,N_2798,N_2800);
nand U3903 (N_3903,N_2091,N_2392);
xnor U3904 (N_3904,N_1990,N_2077);
or U3905 (N_3905,N_2897,N_1855);
and U3906 (N_3906,N_2770,N_2887);
or U3907 (N_3907,N_2195,N_2745);
xor U3908 (N_3908,N_2869,N_1806);
nand U3909 (N_3909,N_2416,N_1660);
xor U3910 (N_3910,N_2883,N_2688);
nor U3911 (N_3911,N_2145,N_2744);
xnor U3912 (N_3912,N_2461,N_2611);
nand U3913 (N_3913,N_2918,N_2767);
and U3914 (N_3914,N_2116,N_1621);
or U3915 (N_3915,N_2526,N_2140);
or U3916 (N_3916,N_2989,N_2282);
or U3917 (N_3917,N_2679,N_2615);
xor U3918 (N_3918,N_2976,N_2368);
and U3919 (N_3919,N_2080,N_1756);
nand U3920 (N_3920,N_2657,N_2994);
and U3921 (N_3921,N_2807,N_1629);
nand U3922 (N_3922,N_2172,N_2743);
nor U3923 (N_3923,N_1594,N_1682);
and U3924 (N_3924,N_1534,N_2490);
and U3925 (N_3925,N_1720,N_2253);
nor U3926 (N_3926,N_2754,N_2673);
nor U3927 (N_3927,N_1644,N_1770);
and U3928 (N_3928,N_2716,N_2360);
or U3929 (N_3929,N_2768,N_1561);
or U3930 (N_3930,N_2547,N_2700);
nand U3931 (N_3931,N_2365,N_1635);
and U3932 (N_3932,N_2161,N_2940);
or U3933 (N_3933,N_2410,N_2887);
nand U3934 (N_3934,N_1807,N_1603);
or U3935 (N_3935,N_1923,N_2572);
or U3936 (N_3936,N_2298,N_2556);
nand U3937 (N_3937,N_2450,N_1660);
or U3938 (N_3938,N_1732,N_2831);
and U3939 (N_3939,N_2716,N_2655);
or U3940 (N_3940,N_2283,N_1605);
nand U3941 (N_3941,N_2146,N_2794);
xnor U3942 (N_3942,N_2076,N_1502);
xor U3943 (N_3943,N_1787,N_1692);
and U3944 (N_3944,N_1934,N_1924);
nor U3945 (N_3945,N_1864,N_2363);
nand U3946 (N_3946,N_1645,N_2765);
or U3947 (N_3947,N_2271,N_1542);
nand U3948 (N_3948,N_1514,N_1833);
and U3949 (N_3949,N_2503,N_1953);
nor U3950 (N_3950,N_2367,N_2467);
and U3951 (N_3951,N_2847,N_1705);
xor U3952 (N_3952,N_2589,N_2499);
xnor U3953 (N_3953,N_2723,N_1588);
or U3954 (N_3954,N_2413,N_2042);
and U3955 (N_3955,N_2246,N_2343);
or U3956 (N_3956,N_1745,N_2291);
or U3957 (N_3957,N_2678,N_2071);
nor U3958 (N_3958,N_2777,N_2757);
nor U3959 (N_3959,N_2500,N_1802);
nor U3960 (N_3960,N_2458,N_2871);
or U3961 (N_3961,N_1841,N_1510);
nand U3962 (N_3962,N_1690,N_2657);
nor U3963 (N_3963,N_1607,N_2667);
or U3964 (N_3964,N_2274,N_1782);
or U3965 (N_3965,N_2524,N_1705);
nand U3966 (N_3966,N_2762,N_1967);
nor U3967 (N_3967,N_2783,N_2047);
nor U3968 (N_3968,N_2746,N_1719);
and U3969 (N_3969,N_2408,N_2458);
or U3970 (N_3970,N_2293,N_2831);
or U3971 (N_3971,N_2906,N_1920);
and U3972 (N_3972,N_2290,N_2718);
or U3973 (N_3973,N_2254,N_1678);
and U3974 (N_3974,N_2764,N_2556);
or U3975 (N_3975,N_1672,N_2043);
nand U3976 (N_3976,N_2039,N_1996);
and U3977 (N_3977,N_2590,N_2899);
and U3978 (N_3978,N_2131,N_1561);
xnor U3979 (N_3979,N_2036,N_1998);
xor U3980 (N_3980,N_1507,N_1729);
xor U3981 (N_3981,N_2101,N_2349);
and U3982 (N_3982,N_2555,N_2290);
and U3983 (N_3983,N_1987,N_2298);
nand U3984 (N_3984,N_2732,N_1593);
or U3985 (N_3985,N_2334,N_2806);
nand U3986 (N_3986,N_2214,N_1725);
and U3987 (N_3987,N_1938,N_2093);
and U3988 (N_3988,N_1997,N_1996);
nor U3989 (N_3989,N_1575,N_2422);
nand U3990 (N_3990,N_2079,N_2091);
and U3991 (N_3991,N_2031,N_2556);
nor U3992 (N_3992,N_2703,N_2575);
xnor U3993 (N_3993,N_1808,N_1905);
xor U3994 (N_3994,N_2658,N_2383);
and U3995 (N_3995,N_2683,N_1762);
xor U3996 (N_3996,N_1765,N_2344);
or U3997 (N_3997,N_2552,N_1531);
xor U3998 (N_3998,N_2444,N_1568);
nor U3999 (N_3999,N_2196,N_2424);
xor U4000 (N_4000,N_2313,N_2437);
nand U4001 (N_4001,N_2317,N_2563);
or U4002 (N_4002,N_2359,N_2468);
or U4003 (N_4003,N_2790,N_2791);
and U4004 (N_4004,N_2321,N_1868);
xnor U4005 (N_4005,N_2610,N_2055);
and U4006 (N_4006,N_2151,N_1968);
xnor U4007 (N_4007,N_1826,N_1601);
or U4008 (N_4008,N_2518,N_1982);
and U4009 (N_4009,N_2821,N_2570);
or U4010 (N_4010,N_2866,N_2188);
nand U4011 (N_4011,N_2750,N_2220);
and U4012 (N_4012,N_2942,N_1622);
or U4013 (N_4013,N_1528,N_2343);
xor U4014 (N_4014,N_1869,N_2529);
xnor U4015 (N_4015,N_1919,N_1822);
xnor U4016 (N_4016,N_1664,N_2491);
or U4017 (N_4017,N_2770,N_2168);
xor U4018 (N_4018,N_2732,N_2062);
nor U4019 (N_4019,N_2020,N_1937);
or U4020 (N_4020,N_2393,N_1702);
nor U4021 (N_4021,N_2288,N_1816);
nand U4022 (N_4022,N_2039,N_2320);
or U4023 (N_4023,N_2732,N_2102);
nor U4024 (N_4024,N_1911,N_1670);
nand U4025 (N_4025,N_2457,N_1744);
and U4026 (N_4026,N_2481,N_2092);
nand U4027 (N_4027,N_2939,N_2117);
and U4028 (N_4028,N_2740,N_1628);
and U4029 (N_4029,N_2394,N_1779);
nor U4030 (N_4030,N_1727,N_2999);
nor U4031 (N_4031,N_2964,N_1642);
nor U4032 (N_4032,N_2956,N_1940);
or U4033 (N_4033,N_1513,N_2058);
xnor U4034 (N_4034,N_1544,N_1934);
and U4035 (N_4035,N_2339,N_2946);
xor U4036 (N_4036,N_1960,N_1892);
nand U4037 (N_4037,N_2767,N_2094);
nand U4038 (N_4038,N_2217,N_2350);
nor U4039 (N_4039,N_2299,N_2944);
or U4040 (N_4040,N_2569,N_2915);
or U4041 (N_4041,N_2153,N_1980);
and U4042 (N_4042,N_2342,N_2433);
nand U4043 (N_4043,N_1821,N_2520);
and U4044 (N_4044,N_2637,N_2646);
nor U4045 (N_4045,N_2149,N_2892);
xnor U4046 (N_4046,N_1981,N_1934);
nand U4047 (N_4047,N_2362,N_2557);
nor U4048 (N_4048,N_2562,N_1554);
and U4049 (N_4049,N_1903,N_2307);
and U4050 (N_4050,N_1513,N_1814);
or U4051 (N_4051,N_2654,N_1592);
or U4052 (N_4052,N_2300,N_2678);
and U4053 (N_4053,N_2915,N_1848);
xor U4054 (N_4054,N_1563,N_2045);
and U4055 (N_4055,N_1528,N_2433);
or U4056 (N_4056,N_1900,N_1803);
nor U4057 (N_4057,N_1509,N_1926);
nand U4058 (N_4058,N_2902,N_2173);
or U4059 (N_4059,N_2881,N_2136);
nor U4060 (N_4060,N_2026,N_1655);
nand U4061 (N_4061,N_1610,N_1599);
nand U4062 (N_4062,N_2273,N_1744);
xor U4063 (N_4063,N_2966,N_1778);
nor U4064 (N_4064,N_2936,N_1805);
and U4065 (N_4065,N_1616,N_2942);
xnor U4066 (N_4066,N_1880,N_2119);
xor U4067 (N_4067,N_1657,N_2584);
nor U4068 (N_4068,N_2213,N_1656);
nor U4069 (N_4069,N_1783,N_1838);
nand U4070 (N_4070,N_2815,N_2867);
nand U4071 (N_4071,N_2789,N_2513);
nor U4072 (N_4072,N_2810,N_2610);
xnor U4073 (N_4073,N_2515,N_1896);
and U4074 (N_4074,N_1956,N_1695);
nand U4075 (N_4075,N_1791,N_2480);
or U4076 (N_4076,N_2507,N_2371);
xnor U4077 (N_4077,N_1946,N_1951);
nor U4078 (N_4078,N_2972,N_1575);
or U4079 (N_4079,N_1542,N_1835);
and U4080 (N_4080,N_1513,N_2695);
nor U4081 (N_4081,N_2270,N_2111);
nor U4082 (N_4082,N_1681,N_1759);
nor U4083 (N_4083,N_2665,N_1671);
and U4084 (N_4084,N_1731,N_1960);
xnor U4085 (N_4085,N_2817,N_2236);
or U4086 (N_4086,N_1540,N_1812);
nor U4087 (N_4087,N_2117,N_1872);
nand U4088 (N_4088,N_2718,N_2191);
or U4089 (N_4089,N_1840,N_1726);
nor U4090 (N_4090,N_2357,N_1604);
or U4091 (N_4091,N_2305,N_2171);
nor U4092 (N_4092,N_2235,N_1747);
or U4093 (N_4093,N_2963,N_1623);
nand U4094 (N_4094,N_2803,N_2673);
or U4095 (N_4095,N_2813,N_1933);
nand U4096 (N_4096,N_2649,N_2749);
nor U4097 (N_4097,N_2526,N_2619);
xor U4098 (N_4098,N_2903,N_2225);
or U4099 (N_4099,N_2346,N_1878);
xor U4100 (N_4100,N_1633,N_2018);
nor U4101 (N_4101,N_2162,N_2388);
nand U4102 (N_4102,N_2855,N_2047);
and U4103 (N_4103,N_2414,N_2896);
xor U4104 (N_4104,N_2094,N_2984);
nor U4105 (N_4105,N_2412,N_2786);
nand U4106 (N_4106,N_2518,N_1776);
and U4107 (N_4107,N_2249,N_2391);
nand U4108 (N_4108,N_2182,N_1834);
nor U4109 (N_4109,N_1776,N_2188);
nand U4110 (N_4110,N_1967,N_1701);
nand U4111 (N_4111,N_2901,N_2474);
nor U4112 (N_4112,N_2665,N_1939);
or U4113 (N_4113,N_2975,N_2727);
xor U4114 (N_4114,N_2198,N_1884);
or U4115 (N_4115,N_2599,N_1594);
nand U4116 (N_4116,N_2753,N_2408);
nor U4117 (N_4117,N_1930,N_1845);
xor U4118 (N_4118,N_1635,N_2003);
nand U4119 (N_4119,N_2981,N_2704);
xnor U4120 (N_4120,N_2268,N_2932);
xnor U4121 (N_4121,N_2671,N_2201);
or U4122 (N_4122,N_1943,N_1654);
xnor U4123 (N_4123,N_2046,N_1927);
nor U4124 (N_4124,N_2482,N_1609);
or U4125 (N_4125,N_1799,N_2772);
nor U4126 (N_4126,N_2356,N_2032);
xor U4127 (N_4127,N_1942,N_1838);
or U4128 (N_4128,N_2602,N_2010);
or U4129 (N_4129,N_2854,N_2564);
or U4130 (N_4130,N_2021,N_2780);
nand U4131 (N_4131,N_2767,N_1789);
or U4132 (N_4132,N_2218,N_2428);
and U4133 (N_4133,N_1899,N_2325);
nor U4134 (N_4134,N_2086,N_2996);
or U4135 (N_4135,N_2139,N_2302);
or U4136 (N_4136,N_1575,N_2705);
or U4137 (N_4137,N_1886,N_1760);
and U4138 (N_4138,N_2329,N_2030);
nand U4139 (N_4139,N_1847,N_1595);
nand U4140 (N_4140,N_1751,N_1921);
or U4141 (N_4141,N_1525,N_2166);
and U4142 (N_4142,N_2278,N_2803);
and U4143 (N_4143,N_2746,N_2234);
xor U4144 (N_4144,N_2609,N_2895);
xnor U4145 (N_4145,N_2415,N_2158);
or U4146 (N_4146,N_1632,N_2996);
nor U4147 (N_4147,N_2057,N_1557);
and U4148 (N_4148,N_2945,N_2809);
nand U4149 (N_4149,N_1929,N_2157);
nand U4150 (N_4150,N_2869,N_2996);
nand U4151 (N_4151,N_2335,N_1635);
or U4152 (N_4152,N_2997,N_2411);
xor U4153 (N_4153,N_2348,N_2845);
nor U4154 (N_4154,N_2063,N_2068);
or U4155 (N_4155,N_1908,N_1750);
nand U4156 (N_4156,N_2167,N_1837);
and U4157 (N_4157,N_1595,N_2154);
xnor U4158 (N_4158,N_2847,N_1734);
and U4159 (N_4159,N_1693,N_2397);
nor U4160 (N_4160,N_2470,N_2746);
nand U4161 (N_4161,N_2619,N_2241);
nor U4162 (N_4162,N_2838,N_1778);
or U4163 (N_4163,N_1643,N_2979);
and U4164 (N_4164,N_2592,N_2911);
or U4165 (N_4165,N_2108,N_2058);
or U4166 (N_4166,N_2369,N_1757);
or U4167 (N_4167,N_2346,N_2337);
and U4168 (N_4168,N_2365,N_2953);
nand U4169 (N_4169,N_1921,N_1957);
and U4170 (N_4170,N_2795,N_2035);
nand U4171 (N_4171,N_2743,N_2965);
and U4172 (N_4172,N_2919,N_2503);
nor U4173 (N_4173,N_2029,N_2811);
nor U4174 (N_4174,N_2777,N_2357);
nor U4175 (N_4175,N_2353,N_2303);
nor U4176 (N_4176,N_2092,N_1640);
and U4177 (N_4177,N_2417,N_2269);
nor U4178 (N_4178,N_1951,N_2483);
and U4179 (N_4179,N_2954,N_1513);
xor U4180 (N_4180,N_2286,N_2391);
nor U4181 (N_4181,N_1747,N_2294);
xnor U4182 (N_4182,N_1678,N_1662);
and U4183 (N_4183,N_2776,N_2785);
nor U4184 (N_4184,N_2136,N_1745);
nand U4185 (N_4185,N_2037,N_1732);
nor U4186 (N_4186,N_1919,N_1620);
or U4187 (N_4187,N_2981,N_2910);
or U4188 (N_4188,N_2179,N_2424);
and U4189 (N_4189,N_2121,N_2856);
nand U4190 (N_4190,N_2347,N_2758);
or U4191 (N_4191,N_2278,N_2411);
and U4192 (N_4192,N_2119,N_2765);
nor U4193 (N_4193,N_2174,N_1726);
nor U4194 (N_4194,N_2032,N_2313);
xor U4195 (N_4195,N_2676,N_1968);
nor U4196 (N_4196,N_2993,N_1723);
and U4197 (N_4197,N_2928,N_2615);
nor U4198 (N_4198,N_2051,N_1952);
xor U4199 (N_4199,N_1549,N_2231);
and U4200 (N_4200,N_2392,N_2540);
and U4201 (N_4201,N_2572,N_1560);
and U4202 (N_4202,N_2080,N_1969);
nand U4203 (N_4203,N_2066,N_2047);
and U4204 (N_4204,N_2404,N_1752);
or U4205 (N_4205,N_1967,N_2858);
or U4206 (N_4206,N_1643,N_2259);
and U4207 (N_4207,N_2614,N_1836);
nand U4208 (N_4208,N_2080,N_2612);
nor U4209 (N_4209,N_2822,N_2542);
and U4210 (N_4210,N_2915,N_2150);
and U4211 (N_4211,N_1759,N_1923);
nor U4212 (N_4212,N_2598,N_1537);
nor U4213 (N_4213,N_1681,N_2471);
xor U4214 (N_4214,N_2405,N_1717);
and U4215 (N_4215,N_2887,N_2626);
xor U4216 (N_4216,N_2255,N_2679);
nor U4217 (N_4217,N_1617,N_1697);
nand U4218 (N_4218,N_2878,N_1745);
xnor U4219 (N_4219,N_2834,N_2100);
and U4220 (N_4220,N_2478,N_2931);
nand U4221 (N_4221,N_1885,N_1967);
xnor U4222 (N_4222,N_1912,N_1528);
and U4223 (N_4223,N_1885,N_2107);
or U4224 (N_4224,N_2032,N_2458);
xnor U4225 (N_4225,N_2791,N_1529);
nand U4226 (N_4226,N_2231,N_1989);
nand U4227 (N_4227,N_2613,N_2364);
or U4228 (N_4228,N_2971,N_2435);
nand U4229 (N_4229,N_2612,N_2682);
nand U4230 (N_4230,N_2071,N_2892);
nor U4231 (N_4231,N_2385,N_2648);
xor U4232 (N_4232,N_2494,N_2924);
nor U4233 (N_4233,N_1536,N_1688);
or U4234 (N_4234,N_2328,N_1710);
nor U4235 (N_4235,N_2832,N_1648);
nor U4236 (N_4236,N_2358,N_2786);
or U4237 (N_4237,N_2415,N_2309);
and U4238 (N_4238,N_2317,N_2903);
or U4239 (N_4239,N_1751,N_2131);
nand U4240 (N_4240,N_2634,N_2835);
or U4241 (N_4241,N_2913,N_2164);
nand U4242 (N_4242,N_1861,N_2621);
nor U4243 (N_4243,N_2697,N_1635);
nor U4244 (N_4244,N_1694,N_2702);
nand U4245 (N_4245,N_2715,N_2184);
xnor U4246 (N_4246,N_2053,N_2661);
nand U4247 (N_4247,N_2812,N_1697);
xnor U4248 (N_4248,N_2047,N_1510);
nand U4249 (N_4249,N_2751,N_2158);
or U4250 (N_4250,N_1536,N_2007);
nor U4251 (N_4251,N_2191,N_2399);
or U4252 (N_4252,N_2603,N_2600);
and U4253 (N_4253,N_2786,N_2301);
nand U4254 (N_4254,N_2075,N_2141);
nand U4255 (N_4255,N_2213,N_1862);
nand U4256 (N_4256,N_2122,N_2262);
xnor U4257 (N_4257,N_1721,N_1994);
or U4258 (N_4258,N_2811,N_2327);
xnor U4259 (N_4259,N_2825,N_1864);
and U4260 (N_4260,N_2476,N_2817);
or U4261 (N_4261,N_2154,N_1917);
nand U4262 (N_4262,N_2950,N_1707);
or U4263 (N_4263,N_1844,N_2326);
and U4264 (N_4264,N_2940,N_1818);
nor U4265 (N_4265,N_2600,N_1616);
nand U4266 (N_4266,N_2848,N_1551);
nor U4267 (N_4267,N_2689,N_2974);
and U4268 (N_4268,N_2411,N_2935);
nor U4269 (N_4269,N_2324,N_1692);
nor U4270 (N_4270,N_1765,N_1856);
nor U4271 (N_4271,N_1633,N_2770);
nand U4272 (N_4272,N_1790,N_1524);
xor U4273 (N_4273,N_1974,N_2186);
xnor U4274 (N_4274,N_2298,N_2808);
or U4275 (N_4275,N_1775,N_2444);
and U4276 (N_4276,N_1792,N_2383);
and U4277 (N_4277,N_1633,N_2827);
or U4278 (N_4278,N_1684,N_2653);
nand U4279 (N_4279,N_2293,N_1500);
and U4280 (N_4280,N_2798,N_2311);
xor U4281 (N_4281,N_2007,N_2164);
nand U4282 (N_4282,N_2733,N_2677);
or U4283 (N_4283,N_2325,N_1557);
and U4284 (N_4284,N_2248,N_2227);
or U4285 (N_4285,N_2489,N_2789);
xnor U4286 (N_4286,N_2656,N_1759);
or U4287 (N_4287,N_2449,N_2526);
nand U4288 (N_4288,N_1633,N_2631);
nand U4289 (N_4289,N_2021,N_2993);
xor U4290 (N_4290,N_2975,N_2780);
and U4291 (N_4291,N_2723,N_2722);
nand U4292 (N_4292,N_2288,N_2853);
nor U4293 (N_4293,N_2347,N_2276);
nor U4294 (N_4294,N_2014,N_1747);
nor U4295 (N_4295,N_2608,N_2093);
nand U4296 (N_4296,N_2286,N_2697);
nor U4297 (N_4297,N_1720,N_1773);
or U4298 (N_4298,N_1813,N_2618);
and U4299 (N_4299,N_1715,N_2916);
and U4300 (N_4300,N_2579,N_1751);
xor U4301 (N_4301,N_2437,N_1600);
and U4302 (N_4302,N_2854,N_2231);
nor U4303 (N_4303,N_1829,N_1966);
and U4304 (N_4304,N_2663,N_1680);
and U4305 (N_4305,N_2687,N_1576);
or U4306 (N_4306,N_2274,N_1592);
nand U4307 (N_4307,N_1669,N_1818);
xor U4308 (N_4308,N_2223,N_2864);
nor U4309 (N_4309,N_2344,N_2485);
nand U4310 (N_4310,N_2487,N_1660);
xnor U4311 (N_4311,N_2127,N_2056);
and U4312 (N_4312,N_1937,N_2592);
nor U4313 (N_4313,N_1997,N_1657);
nor U4314 (N_4314,N_1800,N_2736);
or U4315 (N_4315,N_2450,N_1822);
nand U4316 (N_4316,N_2869,N_2245);
xor U4317 (N_4317,N_2207,N_1937);
nand U4318 (N_4318,N_1999,N_2702);
nor U4319 (N_4319,N_2668,N_2008);
nand U4320 (N_4320,N_2133,N_2147);
or U4321 (N_4321,N_2133,N_2252);
nor U4322 (N_4322,N_1784,N_2720);
or U4323 (N_4323,N_2879,N_2719);
or U4324 (N_4324,N_1788,N_1514);
or U4325 (N_4325,N_2096,N_1697);
or U4326 (N_4326,N_1928,N_2128);
and U4327 (N_4327,N_1950,N_1800);
nand U4328 (N_4328,N_1736,N_2785);
nand U4329 (N_4329,N_1680,N_1606);
nor U4330 (N_4330,N_1633,N_2000);
and U4331 (N_4331,N_2926,N_2486);
or U4332 (N_4332,N_2716,N_2072);
nand U4333 (N_4333,N_2521,N_2281);
xnor U4334 (N_4334,N_1818,N_2400);
and U4335 (N_4335,N_2343,N_2793);
and U4336 (N_4336,N_2371,N_2668);
xor U4337 (N_4337,N_2090,N_2235);
xnor U4338 (N_4338,N_1710,N_2321);
nor U4339 (N_4339,N_2585,N_2956);
or U4340 (N_4340,N_2457,N_2257);
and U4341 (N_4341,N_1660,N_2798);
nand U4342 (N_4342,N_1855,N_1628);
or U4343 (N_4343,N_1854,N_2580);
nand U4344 (N_4344,N_2940,N_1985);
nand U4345 (N_4345,N_2838,N_2413);
xor U4346 (N_4346,N_1509,N_1892);
and U4347 (N_4347,N_1966,N_1911);
xor U4348 (N_4348,N_2768,N_1888);
xnor U4349 (N_4349,N_1928,N_1530);
nor U4350 (N_4350,N_2838,N_2061);
or U4351 (N_4351,N_2296,N_1888);
xnor U4352 (N_4352,N_2459,N_2236);
nor U4353 (N_4353,N_1849,N_2880);
xnor U4354 (N_4354,N_1868,N_1737);
nor U4355 (N_4355,N_1625,N_1954);
and U4356 (N_4356,N_1564,N_2319);
or U4357 (N_4357,N_2350,N_2572);
xor U4358 (N_4358,N_1534,N_1863);
or U4359 (N_4359,N_1698,N_1558);
nor U4360 (N_4360,N_2866,N_1533);
or U4361 (N_4361,N_2586,N_2012);
xor U4362 (N_4362,N_2515,N_2667);
nand U4363 (N_4363,N_1516,N_2327);
nor U4364 (N_4364,N_2563,N_2960);
nand U4365 (N_4365,N_2925,N_1814);
and U4366 (N_4366,N_2724,N_2725);
nand U4367 (N_4367,N_2872,N_2131);
nor U4368 (N_4368,N_1712,N_2319);
nand U4369 (N_4369,N_2236,N_2102);
nor U4370 (N_4370,N_2427,N_1734);
or U4371 (N_4371,N_1991,N_2109);
nand U4372 (N_4372,N_1984,N_2189);
nand U4373 (N_4373,N_2718,N_1764);
xor U4374 (N_4374,N_2840,N_1561);
nand U4375 (N_4375,N_2895,N_2215);
and U4376 (N_4376,N_1690,N_2164);
xor U4377 (N_4377,N_2089,N_2325);
nand U4378 (N_4378,N_1631,N_2551);
and U4379 (N_4379,N_1739,N_1565);
nor U4380 (N_4380,N_2208,N_1556);
xor U4381 (N_4381,N_2731,N_2726);
or U4382 (N_4382,N_1812,N_1643);
nor U4383 (N_4383,N_2265,N_1699);
xor U4384 (N_4384,N_2739,N_2882);
xor U4385 (N_4385,N_1593,N_2879);
nor U4386 (N_4386,N_2634,N_2995);
nand U4387 (N_4387,N_1593,N_2062);
or U4388 (N_4388,N_1833,N_2593);
nor U4389 (N_4389,N_2832,N_1845);
and U4390 (N_4390,N_2347,N_2809);
nand U4391 (N_4391,N_2467,N_2871);
and U4392 (N_4392,N_1881,N_2634);
nand U4393 (N_4393,N_2695,N_1768);
or U4394 (N_4394,N_2338,N_1760);
nor U4395 (N_4395,N_1897,N_2808);
xnor U4396 (N_4396,N_1590,N_2006);
or U4397 (N_4397,N_2125,N_1787);
and U4398 (N_4398,N_2676,N_2703);
nor U4399 (N_4399,N_1894,N_2308);
and U4400 (N_4400,N_2998,N_2573);
xor U4401 (N_4401,N_2236,N_2098);
nand U4402 (N_4402,N_2072,N_2730);
and U4403 (N_4403,N_1769,N_2638);
xnor U4404 (N_4404,N_1881,N_2033);
and U4405 (N_4405,N_2899,N_2349);
xor U4406 (N_4406,N_2749,N_2608);
xor U4407 (N_4407,N_2543,N_2149);
nand U4408 (N_4408,N_2750,N_2434);
nand U4409 (N_4409,N_1695,N_2418);
nor U4410 (N_4410,N_2373,N_2117);
or U4411 (N_4411,N_1787,N_1888);
or U4412 (N_4412,N_1983,N_2014);
xnor U4413 (N_4413,N_2979,N_2350);
or U4414 (N_4414,N_2088,N_1633);
or U4415 (N_4415,N_2956,N_1829);
and U4416 (N_4416,N_1614,N_2847);
nor U4417 (N_4417,N_2964,N_2097);
nor U4418 (N_4418,N_2040,N_2941);
nor U4419 (N_4419,N_2415,N_2608);
or U4420 (N_4420,N_1846,N_1747);
or U4421 (N_4421,N_2491,N_1915);
nor U4422 (N_4422,N_2623,N_1819);
and U4423 (N_4423,N_1802,N_2834);
xor U4424 (N_4424,N_1678,N_2830);
nor U4425 (N_4425,N_1651,N_2489);
nand U4426 (N_4426,N_2772,N_1594);
xnor U4427 (N_4427,N_1640,N_2084);
and U4428 (N_4428,N_1658,N_2232);
nor U4429 (N_4429,N_2867,N_2933);
xnor U4430 (N_4430,N_2105,N_1543);
nand U4431 (N_4431,N_2678,N_2088);
nor U4432 (N_4432,N_2402,N_2571);
and U4433 (N_4433,N_2214,N_2532);
nor U4434 (N_4434,N_2606,N_1933);
nand U4435 (N_4435,N_2710,N_1552);
nand U4436 (N_4436,N_2058,N_2324);
nor U4437 (N_4437,N_1522,N_1546);
xor U4438 (N_4438,N_1564,N_2787);
xnor U4439 (N_4439,N_1993,N_2288);
xor U4440 (N_4440,N_1766,N_2984);
or U4441 (N_4441,N_2377,N_2693);
or U4442 (N_4442,N_1929,N_2638);
nand U4443 (N_4443,N_2171,N_2568);
xor U4444 (N_4444,N_1760,N_2584);
nor U4445 (N_4445,N_1800,N_2204);
and U4446 (N_4446,N_2629,N_1518);
and U4447 (N_4447,N_2774,N_1787);
nor U4448 (N_4448,N_2386,N_2555);
nand U4449 (N_4449,N_2683,N_1526);
nor U4450 (N_4450,N_2163,N_2387);
and U4451 (N_4451,N_1820,N_2740);
or U4452 (N_4452,N_2433,N_2088);
and U4453 (N_4453,N_1980,N_2099);
xor U4454 (N_4454,N_1997,N_2486);
nand U4455 (N_4455,N_2146,N_2364);
nor U4456 (N_4456,N_2365,N_1729);
nor U4457 (N_4457,N_2020,N_2415);
nand U4458 (N_4458,N_2798,N_1742);
and U4459 (N_4459,N_2345,N_2275);
and U4460 (N_4460,N_2470,N_1921);
and U4461 (N_4461,N_2779,N_2680);
and U4462 (N_4462,N_1758,N_1710);
or U4463 (N_4463,N_1832,N_2897);
nor U4464 (N_4464,N_2585,N_2858);
nor U4465 (N_4465,N_2789,N_2638);
xor U4466 (N_4466,N_2606,N_1874);
xnor U4467 (N_4467,N_2391,N_1805);
nor U4468 (N_4468,N_1902,N_1773);
nor U4469 (N_4469,N_1949,N_1748);
or U4470 (N_4470,N_2296,N_1842);
nor U4471 (N_4471,N_2751,N_1814);
nor U4472 (N_4472,N_2404,N_2931);
xnor U4473 (N_4473,N_1797,N_2855);
nand U4474 (N_4474,N_1966,N_1522);
and U4475 (N_4475,N_2828,N_2369);
and U4476 (N_4476,N_2634,N_2635);
xnor U4477 (N_4477,N_2578,N_2375);
nand U4478 (N_4478,N_1520,N_2227);
nand U4479 (N_4479,N_2387,N_2533);
xor U4480 (N_4480,N_2388,N_1931);
xnor U4481 (N_4481,N_2317,N_2216);
xor U4482 (N_4482,N_2863,N_2251);
xnor U4483 (N_4483,N_1843,N_2350);
or U4484 (N_4484,N_2336,N_1721);
xor U4485 (N_4485,N_1872,N_2161);
or U4486 (N_4486,N_2725,N_1666);
and U4487 (N_4487,N_2300,N_1604);
nand U4488 (N_4488,N_2801,N_2957);
and U4489 (N_4489,N_2720,N_1862);
or U4490 (N_4490,N_2591,N_2392);
or U4491 (N_4491,N_2168,N_1988);
nand U4492 (N_4492,N_2047,N_2468);
xor U4493 (N_4493,N_2777,N_2746);
and U4494 (N_4494,N_1698,N_2509);
nor U4495 (N_4495,N_2106,N_2924);
xor U4496 (N_4496,N_2167,N_1773);
xnor U4497 (N_4497,N_2911,N_1601);
nor U4498 (N_4498,N_1701,N_2281);
nor U4499 (N_4499,N_2441,N_1967);
or U4500 (N_4500,N_3598,N_3207);
nand U4501 (N_4501,N_4288,N_3625);
or U4502 (N_4502,N_3931,N_3940);
or U4503 (N_4503,N_3674,N_3681);
nand U4504 (N_4504,N_3618,N_3671);
nor U4505 (N_4505,N_3945,N_3470);
nand U4506 (N_4506,N_3045,N_4142);
and U4507 (N_4507,N_3372,N_4319);
or U4508 (N_4508,N_3528,N_4447);
nand U4509 (N_4509,N_4287,N_3172);
xnor U4510 (N_4510,N_3817,N_3428);
or U4511 (N_4511,N_3384,N_3571);
and U4512 (N_4512,N_3443,N_3461);
nand U4513 (N_4513,N_3190,N_4102);
or U4514 (N_4514,N_3371,N_3853);
and U4515 (N_4515,N_3762,N_3243);
and U4516 (N_4516,N_3125,N_4419);
nand U4517 (N_4517,N_4205,N_4093);
and U4518 (N_4518,N_4075,N_3965);
nor U4519 (N_4519,N_3078,N_3376);
or U4520 (N_4520,N_3669,N_3709);
nor U4521 (N_4521,N_3542,N_3409);
or U4522 (N_4522,N_3582,N_3502);
nor U4523 (N_4523,N_3141,N_3644);
nor U4524 (N_4524,N_3304,N_3905);
nand U4525 (N_4525,N_4403,N_3351);
and U4526 (N_4526,N_3805,N_4017);
and U4527 (N_4527,N_3562,N_3544);
xor U4528 (N_4528,N_3358,N_3918);
nor U4529 (N_4529,N_4049,N_3636);
nand U4530 (N_4530,N_3875,N_4357);
or U4531 (N_4531,N_4266,N_3235);
or U4532 (N_4532,N_4262,N_4192);
or U4533 (N_4533,N_3171,N_3742);
nor U4534 (N_4534,N_3036,N_4218);
xnor U4535 (N_4535,N_3056,N_4136);
xor U4536 (N_4536,N_3118,N_3585);
or U4537 (N_4537,N_3771,N_3793);
or U4538 (N_4538,N_3983,N_4278);
and U4539 (N_4539,N_3193,N_4253);
nor U4540 (N_4540,N_4021,N_4127);
xor U4541 (N_4541,N_4374,N_3816);
and U4542 (N_4542,N_4024,N_4100);
nor U4543 (N_4543,N_4008,N_4420);
nand U4544 (N_4544,N_3276,N_3884);
nand U4545 (N_4545,N_3885,N_3414);
and U4546 (N_4546,N_3436,N_3268);
and U4547 (N_4547,N_3898,N_4290);
nor U4548 (N_4548,N_4472,N_3237);
and U4549 (N_4549,N_3111,N_3189);
nand U4550 (N_4550,N_4281,N_3621);
nor U4551 (N_4551,N_4373,N_3719);
or U4552 (N_4552,N_4191,N_4272);
or U4553 (N_4553,N_4418,N_3240);
or U4554 (N_4554,N_4241,N_4382);
xnor U4555 (N_4555,N_3230,N_4244);
nand U4556 (N_4556,N_3480,N_4364);
nor U4557 (N_4557,N_4067,N_3002);
nor U4558 (N_4558,N_3849,N_3874);
nand U4559 (N_4559,N_3840,N_3293);
and U4560 (N_4560,N_3761,N_3900);
or U4561 (N_4561,N_3442,N_3035);
xnor U4562 (N_4562,N_3570,N_3254);
xnor U4563 (N_4563,N_3845,N_3090);
or U4564 (N_4564,N_4198,N_3511);
nor U4565 (N_4565,N_3925,N_4445);
and U4566 (N_4566,N_3296,N_3252);
nand U4567 (N_4567,N_3693,N_3920);
or U4568 (N_4568,N_3959,N_4004);
nor U4569 (N_4569,N_4026,N_4340);
or U4570 (N_4570,N_3533,N_4425);
and U4571 (N_4571,N_3386,N_3496);
nor U4572 (N_4572,N_4011,N_3370);
or U4573 (N_4573,N_3333,N_3687);
nor U4574 (N_4574,N_4482,N_4435);
nand U4575 (N_4575,N_4139,N_4269);
nor U4576 (N_4576,N_3028,N_4196);
xnor U4577 (N_4577,N_3432,N_4292);
and U4578 (N_4578,N_4280,N_3134);
or U4579 (N_4579,N_3613,N_3795);
or U4580 (N_4580,N_3234,N_3811);
nand U4581 (N_4581,N_4073,N_3128);
xnor U4582 (N_4582,N_3120,N_3173);
nand U4583 (N_4583,N_3708,N_4332);
and U4584 (N_4584,N_3679,N_4389);
xor U4585 (N_4585,N_3199,N_3756);
xor U4586 (N_4586,N_4379,N_3084);
nor U4587 (N_4587,N_4484,N_3808);
and U4588 (N_4588,N_3519,N_3383);
and U4589 (N_4589,N_4108,N_4132);
nand U4590 (N_4590,N_3359,N_3123);
and U4591 (N_4591,N_3616,N_3558);
xnor U4592 (N_4592,N_4215,N_4345);
and U4593 (N_4593,N_3408,N_3292);
nand U4594 (N_4594,N_4462,N_4346);
xor U4595 (N_4595,N_3614,N_3052);
nand U4596 (N_4596,N_3220,N_3332);
nand U4597 (N_4597,N_3773,N_3113);
nand U4598 (N_4598,N_3188,N_3534);
and U4599 (N_4599,N_3556,N_3955);
xnor U4600 (N_4600,N_3588,N_4444);
and U4601 (N_4601,N_3908,N_4053);
nor U4602 (N_4602,N_4454,N_3011);
xnor U4603 (N_4603,N_4165,N_3922);
and U4604 (N_4604,N_3159,N_3749);
nor U4605 (N_4605,N_3325,N_3704);
nand U4606 (N_4606,N_3327,N_4411);
and U4607 (N_4607,N_4044,N_4105);
xnor U4608 (N_4608,N_4200,N_3774);
xor U4609 (N_4609,N_3422,N_3656);
and U4610 (N_4610,N_3591,N_3871);
and U4611 (N_4611,N_3023,N_3835);
nor U4612 (N_4612,N_3993,N_3446);
xnor U4613 (N_4613,N_4414,N_3279);
or U4614 (N_4614,N_4117,N_4208);
xor U4615 (N_4615,N_3663,N_3601);
nand U4616 (N_4616,N_3407,N_3274);
or U4617 (N_4617,N_3569,N_4064);
or U4618 (N_4618,N_3478,N_4178);
nor U4619 (N_4619,N_3635,N_3301);
xor U4620 (N_4620,N_3716,N_4059);
nor U4621 (N_4621,N_4128,N_3798);
and U4622 (N_4622,N_4126,N_4316);
and U4623 (N_4623,N_3445,N_4172);
or U4624 (N_4624,N_3946,N_4209);
nor U4625 (N_4625,N_4333,N_3427);
and U4626 (N_4626,N_4433,N_4378);
and U4627 (N_4627,N_4002,N_4375);
nor U4628 (N_4628,N_3287,N_3144);
xnor U4629 (N_4629,N_3889,N_3072);
xor U4630 (N_4630,N_4099,N_4181);
and U4631 (N_4631,N_3610,N_3532);
and U4632 (N_4632,N_3713,N_3251);
or U4633 (N_4633,N_3291,N_3608);
nor U4634 (N_4634,N_3316,N_4104);
nand U4635 (N_4635,N_3425,N_3140);
nor U4636 (N_4636,N_3812,N_3826);
xnor U4637 (N_4637,N_3824,N_4499);
nor U4638 (N_4638,N_4304,N_3692);
nand U4639 (N_4639,N_3867,N_4167);
nor U4640 (N_4640,N_3701,N_4143);
or U4641 (N_4641,N_3145,N_4315);
nor U4642 (N_4642,N_4112,N_4342);
nor U4643 (N_4643,N_3649,N_3464);
nor U4644 (N_4644,N_4460,N_3214);
nand U4645 (N_4645,N_4271,N_3779);
nand U4646 (N_4646,N_3026,N_4412);
nor U4647 (N_4647,N_3659,N_4083);
xor U4648 (N_4648,N_3441,N_4352);
nor U4649 (N_4649,N_4461,N_4453);
and U4650 (N_4650,N_4034,N_3119);
and U4651 (N_4651,N_3364,N_3154);
or U4652 (N_4652,N_3523,N_3209);
xor U4653 (N_4653,N_4397,N_3772);
nor U4654 (N_4654,N_3334,N_3917);
nand U4655 (N_4655,N_4368,N_3273);
xnor U4656 (N_4656,N_4107,N_3205);
xor U4657 (N_4657,N_4068,N_3387);
and U4658 (N_4658,N_3116,N_4061);
and U4659 (N_4659,N_4161,N_4457);
xnor U4660 (N_4660,N_4284,N_3854);
or U4661 (N_4661,N_3168,N_3479);
nand U4662 (N_4662,N_4398,N_4358);
xor U4663 (N_4663,N_3906,N_4260);
nand U4664 (N_4664,N_4182,N_4338);
and U4665 (N_4665,N_3360,N_4122);
and U4666 (N_4666,N_3888,N_4255);
or U4667 (N_4667,N_3073,N_3328);
xor U4668 (N_4668,N_3087,N_3367);
and U4669 (N_4669,N_3926,N_4301);
nor U4670 (N_4670,N_4310,N_3121);
and U4671 (N_4671,N_4239,N_3305);
nand U4672 (N_4672,N_3633,N_4348);
and U4673 (N_4673,N_3013,N_3403);
nor U4674 (N_4674,N_4238,N_4355);
xor U4675 (N_4675,N_3832,N_3520);
or U4676 (N_4676,N_3350,N_3721);
nand U4677 (N_4677,N_3985,N_3178);
or U4678 (N_4678,N_3789,N_3738);
and U4679 (N_4679,N_4113,N_3748);
or U4680 (N_4680,N_4490,N_3074);
xor U4681 (N_4681,N_3796,N_3069);
and U4682 (N_4682,N_3275,N_3672);
nor U4683 (N_4683,N_3726,N_3280);
nor U4684 (N_4684,N_3236,N_4230);
and U4685 (N_4685,N_4261,N_3759);
nor U4686 (N_4686,N_4179,N_3883);
and U4687 (N_4687,N_3194,N_3987);
nor U4688 (N_4688,N_4109,N_3150);
nor U4689 (N_4689,N_3271,N_3720);
xnor U4690 (N_4690,N_3577,N_3008);
nand U4691 (N_4691,N_3311,N_4001);
nand U4692 (N_4692,N_3546,N_3780);
or U4693 (N_4693,N_3760,N_3213);
xnor U4694 (N_4694,N_3982,N_3994);
nor U4695 (N_4695,N_3752,N_3637);
and U4696 (N_4696,N_4148,N_4030);
or U4697 (N_4697,N_3284,N_3127);
and U4698 (N_4698,N_4050,N_3381);
xor U4699 (N_4699,N_3894,N_3818);
nand U4700 (N_4700,N_4264,N_3343);
nand U4701 (N_4701,N_4145,N_3488);
and U4702 (N_4702,N_4421,N_3054);
xor U4703 (N_4703,N_3554,N_3886);
and U4704 (N_4704,N_3103,N_4018);
or U4705 (N_4705,N_3298,N_3391);
nand U4706 (N_4706,N_4116,N_3664);
nand U4707 (N_4707,N_3083,N_4170);
nor U4708 (N_4708,N_4305,N_3337);
nor U4709 (N_4709,N_4091,N_3001);
or U4710 (N_4710,N_3958,N_3077);
nor U4711 (N_4711,N_4336,N_4121);
and U4712 (N_4712,N_4066,N_4446);
or U4713 (N_4713,N_3426,N_3016);
nor U4714 (N_4714,N_4046,N_4475);
xnor U4715 (N_4715,N_3473,N_3887);
and U4716 (N_4716,N_3952,N_4125);
xor U4717 (N_4717,N_4012,N_3552);
and U4718 (N_4718,N_3551,N_3247);
nor U4719 (N_4719,N_3494,N_3095);
xor U4720 (N_4720,N_3892,N_3318);
nor U4721 (N_4721,N_4394,N_3516);
or U4722 (N_4722,N_3865,N_4443);
xor U4723 (N_4723,N_3563,N_3201);
and U4724 (N_4724,N_4330,N_3971);
nor U4725 (N_4725,N_3498,N_3548);
nor U4726 (N_4726,N_3320,N_3878);
xnor U4727 (N_4727,N_3741,N_4434);
xor U4728 (N_4728,N_3399,N_3303);
and U4729 (N_4729,N_4283,N_3501);
xor U4730 (N_4730,N_4339,N_3718);
nand U4731 (N_4731,N_3617,N_3799);
nor U4732 (N_4732,N_4048,N_3509);
and U4733 (N_4733,N_3731,N_3310);
or U4734 (N_4734,N_3870,N_4430);
and U4735 (N_4735,N_3521,N_3418);
or U4736 (N_4736,N_4496,N_3665);
nor U4737 (N_4737,N_3829,N_3321);
or U4738 (N_4738,N_3363,N_3506);
or U4739 (N_4739,N_4331,N_3203);
and U4740 (N_4740,N_3265,N_3012);
and U4741 (N_4741,N_3629,N_3306);
nor U4742 (N_4742,N_3969,N_4401);
nand U4743 (N_4743,N_4328,N_4385);
nor U4744 (N_4744,N_3882,N_3820);
or U4745 (N_4745,N_3753,N_3264);
nand U4746 (N_4746,N_3737,N_3454);
nor U4747 (N_4747,N_4035,N_3972);
or U4748 (N_4748,N_3513,N_4483);
and U4749 (N_4749,N_3725,N_4450);
nand U4750 (N_4750,N_3338,N_3881);
nand U4751 (N_4751,N_4162,N_3981);
xnor U4752 (N_4752,N_3431,N_3702);
or U4753 (N_4753,N_3677,N_4185);
and U4754 (N_4754,N_3219,N_3819);
and U4755 (N_4755,N_3825,N_4028);
xor U4756 (N_4756,N_3104,N_3057);
nand U4757 (N_4757,N_3472,N_3339);
nor U4758 (N_4758,N_3970,N_3806);
or U4759 (N_4759,N_3248,N_3602);
or U4760 (N_4760,N_3196,N_3711);
xor U4761 (N_4761,N_3182,N_4089);
nor U4762 (N_4762,N_3575,N_3034);
nor U4763 (N_4763,N_3105,N_3091);
and U4764 (N_4764,N_3923,N_3967);
xnor U4765 (N_4765,N_4361,N_3146);
nand U4766 (N_4766,N_3323,N_3504);
nor U4767 (N_4767,N_4251,N_3560);
xor U4768 (N_4768,N_4173,N_3272);
or U4769 (N_4769,N_4497,N_3453);
and U4770 (N_4770,N_3216,N_3080);
nor U4771 (N_4771,N_4481,N_3787);
xor U4772 (N_4772,N_4219,N_4234);
and U4773 (N_4773,N_3014,N_3648);
nand U4774 (N_4774,N_4413,N_4402);
xor U4775 (N_4775,N_4118,N_4249);
nor U4776 (N_4776,N_3053,N_3675);
xor U4777 (N_4777,N_3382,N_4417);
nor U4778 (N_4778,N_3257,N_4084);
xnor U4779 (N_4779,N_3587,N_3162);
or U4780 (N_4780,N_3930,N_3076);
nor U4781 (N_4781,N_3345,N_4190);
nand U4782 (N_4782,N_4029,N_3312);
xor U4783 (N_4783,N_3195,N_4381);
nor U4784 (N_4784,N_3584,N_4452);
or U4785 (N_4785,N_4031,N_4211);
or U4786 (N_4786,N_3263,N_3661);
xor U4787 (N_4787,N_3522,N_3107);
nand U4788 (N_4788,N_3137,N_3902);
nor U4789 (N_4789,N_3262,N_3007);
or U4790 (N_4790,N_4156,N_3593);
xor U4791 (N_4791,N_3068,N_4405);
xor U4792 (N_4792,N_3973,N_4495);
nand U4793 (N_4793,N_4257,N_4221);
xnor U4794 (N_4794,N_4223,N_3754);
nor U4795 (N_4795,N_3942,N_4195);
or U4796 (N_4796,N_3149,N_4087);
nand U4797 (N_4797,N_4360,N_3932);
nor U4798 (N_4798,N_3114,N_3241);
nand U4799 (N_4799,N_4214,N_4123);
xnor U4800 (N_4800,N_4224,N_3487);
nor U4801 (N_4801,N_3491,N_4110);
and U4802 (N_4802,N_3861,N_3896);
or U4803 (N_4803,N_3775,N_3331);
xnor U4804 (N_4804,N_3109,N_4387);
nor U4805 (N_4805,N_3647,N_3206);
nand U4806 (N_4806,N_3483,N_3346);
nand U4807 (N_4807,N_3515,N_3846);
nand U4808 (N_4808,N_3943,N_4163);
xor U4809 (N_4809,N_4268,N_3065);
and U4810 (N_4810,N_3683,N_3757);
nor U4811 (N_4811,N_3654,N_3895);
nor U4812 (N_4812,N_3727,N_3911);
nor U4813 (N_4813,N_3691,N_4488);
or U4814 (N_4814,N_3463,N_3837);
nor U4815 (N_4815,N_3475,N_3336);
nor U4816 (N_4816,N_4404,N_4456);
or U4817 (N_4817,N_3486,N_4432);
or U4818 (N_4818,N_3088,N_3904);
nand U4819 (N_4819,N_4133,N_3361);
nand U4820 (N_4820,N_3995,N_3747);
xor U4821 (N_4821,N_3844,N_4370);
nand U4822 (N_4822,N_3822,N_3750);
nor U4823 (N_4823,N_4070,N_3344);
nor U4824 (N_4824,N_3549,N_3999);
xnor U4825 (N_4825,N_3100,N_3096);
xnor U4826 (N_4826,N_4273,N_4060);
or U4827 (N_4827,N_3836,N_3434);
nor U4828 (N_4828,N_3139,N_4337);
nand U4829 (N_4829,N_4036,N_3000);
or U4830 (N_4830,N_3813,N_4436);
nand U4831 (N_4831,N_3978,N_4400);
nand U4832 (N_4832,N_4039,N_4320);
or U4833 (N_4833,N_4473,N_3167);
nor U4834 (N_4834,N_3393,N_3927);
xnor U4835 (N_4835,N_4243,N_3156);
nor U4836 (N_4836,N_3031,N_3783);
xor U4837 (N_4837,N_3990,N_3245);
nand U4838 (N_4838,N_3791,N_3921);
or U4839 (N_4839,N_3842,N_4354);
xnor U4840 (N_4840,N_3015,N_3603);
and U4841 (N_4841,N_3622,N_4033);
and U4842 (N_4842,N_4151,N_4479);
or U4843 (N_4843,N_4392,N_3862);
nor U4844 (N_4844,N_4052,N_4094);
nand U4845 (N_4845,N_4303,N_3413);
nor U4846 (N_4846,N_3354,N_3180);
nor U4847 (N_4847,N_3085,N_3541);
xor U4848 (N_4848,N_4246,N_3368);
nor U4849 (N_4849,N_3619,N_4144);
nand U4850 (N_4850,N_4040,N_4476);
nor U4851 (N_4851,N_3181,N_3295);
or U4852 (N_4852,N_4265,N_3868);
nor U4853 (N_4853,N_3954,N_3379);
nor U4854 (N_4854,N_4371,N_3580);
or U4855 (N_4855,N_4146,N_4259);
xnor U4856 (N_4856,N_3531,N_3489);
or U4857 (N_4857,N_4206,N_4428);
xor U4858 (N_4858,N_3746,N_3055);
and U4859 (N_4859,N_4438,N_3075);
xnor U4860 (N_4860,N_3690,N_3147);
nand U4861 (N_4861,N_4494,N_4097);
nand U4862 (N_4862,N_3503,N_3830);
and U4863 (N_4863,N_3365,N_4359);
xnor U4864 (N_4864,N_3689,N_3565);
or U4865 (N_4865,N_4362,N_3438);
nand U4866 (N_4866,N_3872,N_3377);
or U4867 (N_4867,N_3559,N_3006);
nor U4868 (N_4868,N_3838,N_4470);
nor U4869 (N_4869,N_3153,N_4323);
nand U4870 (N_4870,N_3815,N_3948);
and U4871 (N_4871,N_3632,N_3061);
xnor U4872 (N_4872,N_3115,N_3703);
or U4873 (N_4873,N_3723,N_4171);
and U4874 (N_4874,N_3313,N_3729);
and U4875 (N_4875,N_3841,N_3583);
or U4876 (N_4876,N_3831,N_4111);
nor U4877 (N_4877,N_4376,N_3266);
or U4878 (N_4878,N_4153,N_4322);
nand U4879 (N_4879,N_3781,N_3395);
nor U4880 (N_4880,N_3916,N_3801);
and U4881 (N_4881,N_3277,N_3698);
xor U4882 (N_4882,N_3309,N_3106);
xnor U4883 (N_4883,N_3707,N_4166);
and U4884 (N_4884,N_4180,N_3020);
and U4885 (N_4885,N_3576,N_3717);
nand U4886 (N_4886,N_4065,N_3374);
or U4887 (N_4887,N_4313,N_4082);
nor U4888 (N_4888,N_4441,N_3540);
nor U4889 (N_4889,N_3050,N_4240);
nor U4890 (N_4890,N_3782,N_3545);
xnor U4891 (N_4891,N_3025,N_3152);
xor U4892 (N_4892,N_3863,N_4351);
and U4893 (N_4893,N_3929,N_3198);
xor U4894 (N_4894,N_4309,N_3200);
and U4895 (N_4895,N_4384,N_3030);
xor U4896 (N_4896,N_4212,N_3192);
and U4897 (N_4897,N_3094,N_3968);
nor U4898 (N_4898,N_3785,N_4295);
nand U4899 (N_4899,N_3640,N_3136);
xor U4900 (N_4900,N_4135,N_3224);
and U4901 (N_4901,N_3440,N_3249);
nor U4902 (N_4902,N_3324,N_4349);
and U4903 (N_4903,N_3101,N_3143);
nor U4904 (N_4904,N_3221,N_4101);
nand U4905 (N_4905,N_4367,N_3956);
and U4906 (N_4906,N_4155,N_3928);
nand U4907 (N_4907,N_3732,N_3357);
nand U4908 (N_4908,N_4194,N_4147);
or U4909 (N_4909,N_3112,N_3244);
or U4910 (N_4910,N_4286,N_4289);
nand U4911 (N_4911,N_3238,N_3300);
nor U4912 (N_4912,N_3957,N_3131);
nor U4913 (N_4913,N_4137,N_3218);
or U4914 (N_4914,N_3536,N_3398);
nor U4915 (N_4915,N_4047,N_3326);
nand U4916 (N_4916,N_3512,N_4267);
or U4917 (N_4917,N_3497,N_4321);
and U4918 (N_4918,N_3660,N_3490);
or U4919 (N_4919,N_4062,N_3535);
or U4920 (N_4920,N_3250,N_4037);
nor U4921 (N_4921,N_4159,N_3514);
nand U4922 (N_4922,N_3233,N_3634);
xnor U4923 (N_4923,N_3526,N_4335);
nor U4924 (N_4924,N_4051,N_3062);
nor U4925 (N_4925,N_3071,N_4458);
and U4926 (N_4926,N_3694,N_3261);
xnor U4927 (N_4927,N_4098,N_3110);
nor U4928 (N_4928,N_3040,N_3722);
nor U4929 (N_4929,N_4282,N_4217);
nor U4930 (N_4930,N_4324,N_3505);
nand U4931 (N_4931,N_3596,N_3079);
nand U4932 (N_4932,N_4410,N_3572);
nand U4933 (N_4933,N_3627,N_4439);
nor U4934 (N_4934,N_3089,N_4076);
or U4935 (N_4935,N_3005,N_4003);
and U4936 (N_4936,N_3856,N_3270);
nor U4937 (N_4937,N_4106,N_3643);
and U4938 (N_4938,N_3070,N_3476);
xor U4939 (N_4939,N_3185,N_3223);
xor U4940 (N_4940,N_4042,N_3017);
xor U4941 (N_4941,N_3620,N_3850);
nor U4942 (N_4942,N_4274,N_3670);
and U4943 (N_4943,N_3004,N_4467);
nor U4944 (N_4944,N_3208,N_4186);
or U4945 (N_4945,N_3047,N_4063);
xnor U4946 (N_4946,N_3495,N_3651);
xor U4947 (N_4947,N_4056,N_3439);
and U4948 (N_4948,N_3517,N_3764);
nand U4949 (N_4949,N_4485,N_3474);
nor U4950 (N_4950,N_3728,N_3124);
and U4951 (N_4951,N_4276,N_3724);
and U4952 (N_4952,N_3421,N_4248);
nand U4953 (N_4953,N_3566,N_4160);
nand U4954 (N_4954,N_3961,N_4463);
xor U4955 (N_4955,N_3373,N_4369);
and U4956 (N_4956,N_3048,N_3404);
nand U4957 (N_4957,N_4231,N_3433);
xor U4958 (N_4958,N_3657,N_4124);
nor U4959 (N_4959,N_4201,N_4055);
nor U4960 (N_4960,N_3997,N_3873);
and U4961 (N_4961,N_3067,N_4174);
nor U4962 (N_4962,N_3730,N_4079);
nor U4963 (N_4963,N_3186,N_3743);
or U4964 (N_4964,N_3288,N_4119);
xor U4965 (N_4965,N_3555,N_4471);
and U4966 (N_4966,N_3890,N_4175);
or U4967 (N_4967,N_4365,N_3527);
xnor U4968 (N_4968,N_3944,N_3163);
nor U4969 (N_4969,N_3976,N_3449);
and U4970 (N_4970,N_3462,N_3353);
nor U4971 (N_4971,N_4353,N_3392);
or U4972 (N_4972,N_3282,N_3184);
and U4973 (N_4973,N_3049,N_3966);
nor U4974 (N_4974,N_4285,N_3910);
xnor U4975 (N_4975,N_4237,N_3777);
or U4976 (N_4976,N_3744,N_4183);
and U4977 (N_4977,N_3043,N_3086);
and U4978 (N_4978,N_4210,N_3564);
and U4979 (N_4979,N_3117,N_3807);
nor U4980 (N_4980,N_3667,N_4498);
and U4981 (N_4981,N_3524,N_3860);
and U4982 (N_4982,N_4177,N_3626);
nor U4983 (N_4983,N_3739,N_3733);
nor U4984 (N_4984,N_4489,N_3477);
xnor U4985 (N_4985,N_4086,N_4297);
or U4986 (N_4986,N_3607,N_4242);
xor U4987 (N_4987,N_3022,N_3645);
or U4988 (N_4988,N_4188,N_4213);
nand U4989 (N_4989,N_3876,N_3977);
nand U4990 (N_4990,N_4427,N_3423);
nor U4991 (N_4991,N_4092,N_3385);
nor U4992 (N_4992,N_3242,N_3051);
nand U4993 (N_4993,N_4391,N_4225);
xnor U4994 (N_4994,N_3755,N_4277);
nand U4995 (N_4995,N_3388,N_3138);
or U4996 (N_4996,N_3212,N_3460);
nand U4997 (N_4997,N_4252,N_4492);
nand U4998 (N_4998,N_4422,N_3027);
and U4999 (N_4999,N_3215,N_3809);
nand U5000 (N_5000,N_3624,N_3467);
nand U5001 (N_5001,N_4074,N_4393);
nand U5002 (N_5002,N_4256,N_3864);
nand U5003 (N_5003,N_3126,N_3029);
nor U5004 (N_5004,N_3700,N_3880);
and U5005 (N_5005,N_4149,N_4329);
and U5006 (N_5006,N_3590,N_3609);
nand U5007 (N_5007,N_4306,N_3599);
or U5008 (N_5008,N_4254,N_3340);
or U5009 (N_5009,N_3988,N_4415);
and U5010 (N_5010,N_3435,N_3919);
xor U5011 (N_5011,N_3375,N_3855);
nand U5012 (N_5012,N_4408,N_3623);
nor U5013 (N_5013,N_3606,N_3529);
or U5014 (N_5014,N_3405,N_3269);
or U5015 (N_5015,N_3155,N_3823);
and U5016 (N_5016,N_3934,N_3630);
or U5017 (N_5017,N_3736,N_3851);
xor U5018 (N_5018,N_3557,N_4247);
nor U5019 (N_5019,N_4459,N_3650);
nand U5020 (N_5020,N_4383,N_3589);
or U5021 (N_5021,N_3652,N_3175);
nand U5022 (N_5022,N_4207,N_3897);
xnor U5023 (N_5023,N_4424,N_3914);
nor U5024 (N_5024,N_3989,N_3227);
xor U5025 (N_5025,N_3676,N_3401);
or U5026 (N_5026,N_3228,N_3662);
nor U5027 (N_5027,N_3776,N_3866);
and U5028 (N_5028,N_3044,N_4486);
nor U5029 (N_5029,N_3960,N_3682);
nor U5030 (N_5030,N_4130,N_3335);
nor U5031 (N_5031,N_3037,N_3539);
nand U5032 (N_5032,N_3594,N_4318);
nand U5033 (N_5033,N_4293,N_4477);
and U5034 (N_5034,N_4245,N_3493);
nor U5035 (N_5035,N_3597,N_4078);
nand U5036 (N_5036,N_4096,N_3060);
nand U5037 (N_5037,N_3009,N_3605);
xor U5038 (N_5038,N_3631,N_3869);
xor U5039 (N_5039,N_3169,N_3996);
and U5040 (N_5040,N_3903,N_3992);
nor U5041 (N_5041,N_4327,N_3794);
nand U5042 (N_5042,N_3450,N_3349);
and U5043 (N_5043,N_3686,N_4164);
nand U5044 (N_5044,N_3471,N_3567);
and U5045 (N_5045,N_3991,N_3530);
xnor U5046 (N_5046,N_3684,N_3259);
xnor U5047 (N_5047,N_3232,N_3611);
or U5048 (N_5048,N_3448,N_3191);
nand U5049 (N_5049,N_4090,N_3765);
nor U5050 (N_5050,N_4114,N_3417);
and U5051 (N_5051,N_3518,N_3802);
nor U5052 (N_5052,N_4226,N_4311);
or U5053 (N_5053,N_3745,N_3093);
xnor U5054 (N_5054,N_3455,N_3947);
or U5055 (N_5055,N_4270,N_3907);
and U5056 (N_5056,N_4493,N_3581);
or U5057 (N_5057,N_4449,N_4027);
xor U5058 (N_5058,N_3998,N_3406);
nand U5059 (N_5059,N_3941,N_4250);
or U5060 (N_5060,N_3658,N_3986);
xnor U5061 (N_5061,N_4088,N_3024);
nand U5062 (N_5062,N_3740,N_3380);
and U5063 (N_5063,N_4466,N_4474);
and U5064 (N_5064,N_3308,N_3267);
nor U5065 (N_5065,N_3937,N_3797);
nand U5066 (N_5066,N_3909,N_3456);
nand U5067 (N_5067,N_3416,N_4129);
and U5068 (N_5068,N_4298,N_4307);
or U5069 (N_5069,N_4399,N_3294);
nand U5070 (N_5070,N_3229,N_4232);
nor U5071 (N_5071,N_4396,N_3457);
nor U5072 (N_5072,N_3766,N_3314);
xor U5073 (N_5073,N_4189,N_4199);
nor U5074 (N_5074,N_4158,N_3315);
nand U5075 (N_5075,N_3166,N_3715);
or U5076 (N_5076,N_4491,N_3410);
and U5077 (N_5077,N_3019,N_4038);
and U5078 (N_5078,N_3042,N_3400);
or U5079 (N_5079,N_3366,N_3924);
xor U5080 (N_5080,N_4395,N_3839);
nand U5081 (N_5081,N_3612,N_3452);
nor U5082 (N_5082,N_3164,N_4203);
or U5083 (N_5083,N_4157,N_3177);
and U5084 (N_5084,N_4043,N_3814);
or U5085 (N_5085,N_4006,N_3933);
nand U5086 (N_5086,N_3210,N_3362);
nor U5087 (N_5087,N_4487,N_3033);
xnor U5088 (N_5088,N_3901,N_3424);
nand U5089 (N_5089,N_3289,N_4220);
nand U5090 (N_5090,N_3769,N_3891);
nor U5091 (N_5091,N_3058,N_4275);
nor U5092 (N_5092,N_4300,N_4480);
or U5093 (N_5093,N_3899,N_3507);
xor U5094 (N_5094,N_4216,N_3231);
nand U5095 (N_5095,N_4442,N_3547);
or U5096 (N_5096,N_4431,N_3678);
or U5097 (N_5097,N_3299,N_3397);
nand U5098 (N_5098,N_4347,N_3628);
or U5099 (N_5099,N_3132,N_4317);
xor U5100 (N_5100,N_3834,N_3319);
nor U5101 (N_5101,N_4258,N_4085);
nand U5102 (N_5102,N_4291,N_3459);
nor U5103 (N_5103,N_3394,N_3705);
nor U5104 (N_5104,N_3668,N_3763);
xor U5105 (N_5105,N_3187,N_4000);
nor U5106 (N_5106,N_3352,N_4071);
xor U5107 (N_5107,N_4279,N_3915);
nor U5108 (N_5108,N_3803,N_3356);
xor U5109 (N_5109,N_3396,N_3130);
or U5110 (N_5110,N_4103,N_3226);
and U5111 (N_5111,N_3500,N_3939);
nand U5112 (N_5112,N_3786,N_3032);
and U5113 (N_5113,N_3082,N_3211);
and U5114 (N_5114,N_3734,N_3165);
nand U5115 (N_5115,N_3197,N_3767);
xnor U5116 (N_5116,N_4152,N_3974);
nand U5117 (N_5117,N_3041,N_3962);
and U5118 (N_5118,N_4363,N_3142);
nand U5119 (N_5119,N_3810,N_3176);
xor U5120 (N_5120,N_4007,N_3258);
xor U5121 (N_5121,N_4154,N_4041);
xnor U5122 (N_5122,N_4372,N_4350);
nor U5123 (N_5123,N_4233,N_4228);
or U5124 (N_5124,N_3161,N_4045);
or U5125 (N_5125,N_3951,N_4197);
xor U5126 (N_5126,N_4429,N_3097);
xor U5127 (N_5127,N_4193,N_3322);
and U5128 (N_5128,N_4015,N_4140);
xnor U5129 (N_5129,N_3788,N_3317);
nor U5130 (N_5130,N_3290,N_4356);
nand U5131 (N_5131,N_4478,N_3297);
xnor U5132 (N_5132,N_4468,N_4451);
nand U5133 (N_5133,N_4344,N_4406);
nor U5134 (N_5134,N_3949,N_3821);
or U5135 (N_5135,N_3102,N_3550);
or U5136 (N_5136,N_4054,N_3174);
xor U5137 (N_5137,N_3712,N_3979);
and U5138 (N_5138,N_3792,N_3710);
or U5139 (N_5139,N_4020,N_3980);
and U5140 (N_5140,N_3278,N_3568);
and U5141 (N_5141,N_3561,N_3347);
or U5142 (N_5142,N_3225,N_3429);
nand U5143 (N_5143,N_3466,N_4023);
or U5144 (N_5144,N_3857,N_4423);
and U5145 (N_5145,N_3604,N_4058);
nor U5146 (N_5146,N_3342,N_3525);
and U5147 (N_5147,N_3646,N_4014);
nor U5148 (N_5148,N_4314,N_4263);
nor U5149 (N_5149,N_4325,N_3538);
nand U5150 (N_5150,N_4169,N_3437);
nor U5151 (N_5151,N_3447,N_3348);
nand U5152 (N_5152,N_3800,N_3064);
and U5153 (N_5153,N_4016,N_3666);
xnor U5154 (N_5154,N_3389,N_3492);
nor U5155 (N_5155,N_3615,N_4013);
or U5156 (N_5156,N_3260,N_3784);
xnor U5157 (N_5157,N_4227,N_3574);
and U5158 (N_5158,N_4005,N_3697);
or U5159 (N_5159,N_3833,N_3484);
nand U5160 (N_5160,N_3510,N_3129);
nor U5161 (N_5161,N_4077,N_4236);
or U5162 (N_5162,N_3573,N_3953);
and U5163 (N_5163,N_3444,N_3595);
xor U5164 (N_5164,N_3706,N_3655);
or U5165 (N_5165,N_3642,N_3217);
nand U5166 (N_5166,N_4377,N_4229);
and U5167 (N_5167,N_3179,N_3046);
or U5168 (N_5168,N_3688,N_3696);
xnor U5169 (N_5169,N_4390,N_4299);
nor U5170 (N_5170,N_3935,N_4388);
nor U5171 (N_5171,N_3653,N_3858);
xor U5172 (N_5172,N_4081,N_3600);
xnor U5173 (N_5173,N_3038,N_3133);
or U5174 (N_5174,N_3003,N_4312);
xnor U5175 (N_5175,N_4409,N_4334);
nand U5176 (N_5176,N_4010,N_3063);
and U5177 (N_5177,N_3283,N_3768);
nand U5178 (N_5178,N_3950,N_3092);
or U5179 (N_5179,N_4296,N_3638);
or U5180 (N_5180,N_3021,N_4202);
nor U5181 (N_5181,N_4426,N_4302);
and U5182 (N_5182,N_4069,N_3578);
xor U5183 (N_5183,N_4341,N_3255);
and U5184 (N_5184,N_4326,N_4057);
and U5185 (N_5185,N_4025,N_3010);
and U5186 (N_5186,N_4455,N_3913);
and U5187 (N_5187,N_3482,N_3804);
and U5188 (N_5188,N_3419,N_4131);
nand U5189 (N_5189,N_3081,N_4184);
and U5190 (N_5190,N_3222,N_3778);
or U5191 (N_5191,N_3770,N_4138);
nor U5192 (N_5192,N_4120,N_3469);
or U5193 (N_5193,N_3246,N_3039);
xor U5194 (N_5194,N_3893,N_4019);
xnor U5195 (N_5195,N_3695,N_3202);
nand U5196 (N_5196,N_4235,N_3170);
nor U5197 (N_5197,N_4380,N_3330);
xnor U5198 (N_5198,N_3099,N_3984);
and U5199 (N_5199,N_3256,N_3239);
xnor U5200 (N_5200,N_4440,N_3499);
nor U5201 (N_5201,N_4308,N_4009);
nor U5202 (N_5202,N_4437,N_3378);
or U5203 (N_5203,N_3098,N_3714);
and U5204 (N_5204,N_4465,N_3579);
nor U5205 (N_5205,N_3430,N_3465);
nand U5206 (N_5206,N_4080,N_4134);
nor U5207 (N_5207,N_3329,N_3828);
nor U5208 (N_5208,N_4176,N_4095);
xor U5209 (N_5209,N_3412,N_3286);
or U5210 (N_5210,N_4032,N_3018);
nand U5211 (N_5211,N_4469,N_3302);
nand U5212 (N_5212,N_3157,N_3415);
xor U5213 (N_5213,N_4294,N_3790);
nor U5214 (N_5214,N_4115,N_3843);
xnor U5215 (N_5215,N_3066,N_4187);
nor U5216 (N_5216,N_3912,N_3827);
xor U5217 (N_5217,N_4204,N_3964);
xor U5218 (N_5218,N_4168,N_4366);
or U5219 (N_5219,N_4222,N_3543);
nand U5220 (N_5220,N_3420,N_3553);
xor U5221 (N_5221,N_3281,N_4343);
xnor U5222 (N_5222,N_3285,N_3108);
xor U5223 (N_5223,N_3641,N_3485);
and U5224 (N_5224,N_3877,N_3135);
nor U5225 (N_5225,N_3879,N_4407);
nor U5226 (N_5226,N_3158,N_3699);
nor U5227 (N_5227,N_3369,N_3639);
xor U5228 (N_5228,N_3735,N_4448);
nand U5229 (N_5229,N_3963,N_3122);
or U5230 (N_5230,N_4464,N_3852);
nor U5231 (N_5231,N_4386,N_3975);
and U5232 (N_5232,N_3468,N_3183);
nand U5233 (N_5233,N_4022,N_3680);
nand U5234 (N_5234,N_3758,N_3936);
xor U5235 (N_5235,N_3537,N_3481);
nor U5236 (N_5236,N_3508,N_3938);
and U5237 (N_5237,N_3390,N_3451);
nand U5238 (N_5238,N_3685,N_3586);
nor U5239 (N_5239,N_3148,N_3341);
xor U5240 (N_5240,N_3402,N_3253);
or U5241 (N_5241,N_4072,N_3411);
xor U5242 (N_5242,N_4416,N_3592);
nand U5243 (N_5243,N_4141,N_4150);
nand U5244 (N_5244,N_3673,N_3848);
nor U5245 (N_5245,N_3160,N_3151);
or U5246 (N_5246,N_3355,N_3307);
nand U5247 (N_5247,N_3847,N_3458);
and U5248 (N_5248,N_3204,N_3859);
nand U5249 (N_5249,N_3059,N_3751);
or U5250 (N_5250,N_3653,N_3955);
and U5251 (N_5251,N_3791,N_3307);
nand U5252 (N_5252,N_4443,N_4238);
or U5253 (N_5253,N_3035,N_3175);
nor U5254 (N_5254,N_3868,N_3713);
nor U5255 (N_5255,N_3513,N_3713);
nor U5256 (N_5256,N_3603,N_4060);
or U5257 (N_5257,N_3619,N_4155);
nand U5258 (N_5258,N_3703,N_3959);
xor U5259 (N_5259,N_3380,N_4070);
nand U5260 (N_5260,N_3290,N_3603);
nand U5261 (N_5261,N_3880,N_4036);
or U5262 (N_5262,N_3654,N_3383);
and U5263 (N_5263,N_3676,N_3415);
or U5264 (N_5264,N_3837,N_3681);
and U5265 (N_5265,N_3111,N_3095);
nand U5266 (N_5266,N_3734,N_4180);
and U5267 (N_5267,N_3634,N_3770);
nor U5268 (N_5268,N_3593,N_4105);
nand U5269 (N_5269,N_3474,N_4340);
nand U5270 (N_5270,N_4213,N_3066);
or U5271 (N_5271,N_4105,N_3942);
or U5272 (N_5272,N_4175,N_3532);
and U5273 (N_5273,N_4178,N_3466);
and U5274 (N_5274,N_3529,N_3990);
nand U5275 (N_5275,N_3519,N_4291);
nand U5276 (N_5276,N_3674,N_3566);
xor U5277 (N_5277,N_3896,N_3232);
nand U5278 (N_5278,N_4316,N_4361);
nor U5279 (N_5279,N_3811,N_4213);
nand U5280 (N_5280,N_3659,N_3971);
or U5281 (N_5281,N_3932,N_3680);
and U5282 (N_5282,N_3216,N_4235);
nand U5283 (N_5283,N_3679,N_3056);
and U5284 (N_5284,N_3985,N_3843);
and U5285 (N_5285,N_3540,N_4290);
xnor U5286 (N_5286,N_3116,N_4210);
or U5287 (N_5287,N_3454,N_4428);
nand U5288 (N_5288,N_4323,N_4380);
nor U5289 (N_5289,N_3808,N_3227);
or U5290 (N_5290,N_4393,N_3191);
nand U5291 (N_5291,N_3221,N_3215);
nor U5292 (N_5292,N_3767,N_4333);
nand U5293 (N_5293,N_4335,N_3489);
and U5294 (N_5294,N_3090,N_4275);
and U5295 (N_5295,N_4333,N_3877);
nand U5296 (N_5296,N_4475,N_3250);
and U5297 (N_5297,N_3023,N_4281);
nor U5298 (N_5298,N_3460,N_3800);
xor U5299 (N_5299,N_3809,N_4354);
xor U5300 (N_5300,N_3517,N_3548);
nor U5301 (N_5301,N_4483,N_3269);
nand U5302 (N_5302,N_3139,N_3807);
nor U5303 (N_5303,N_4010,N_3716);
and U5304 (N_5304,N_3744,N_4230);
or U5305 (N_5305,N_3502,N_3211);
nand U5306 (N_5306,N_3219,N_4408);
or U5307 (N_5307,N_4062,N_3786);
or U5308 (N_5308,N_3550,N_3581);
xnor U5309 (N_5309,N_3572,N_3661);
and U5310 (N_5310,N_3109,N_4142);
and U5311 (N_5311,N_4412,N_4313);
and U5312 (N_5312,N_3694,N_4327);
xnor U5313 (N_5313,N_3028,N_3193);
or U5314 (N_5314,N_4114,N_3773);
xor U5315 (N_5315,N_3690,N_3619);
nand U5316 (N_5316,N_3834,N_4408);
nand U5317 (N_5317,N_3360,N_3743);
or U5318 (N_5318,N_3716,N_4467);
or U5319 (N_5319,N_3106,N_3939);
xor U5320 (N_5320,N_3821,N_3378);
and U5321 (N_5321,N_4378,N_3550);
nor U5322 (N_5322,N_3204,N_3513);
and U5323 (N_5323,N_3900,N_3922);
and U5324 (N_5324,N_3109,N_3478);
xor U5325 (N_5325,N_3689,N_3180);
and U5326 (N_5326,N_3068,N_3211);
nor U5327 (N_5327,N_4087,N_4392);
or U5328 (N_5328,N_4450,N_3137);
or U5329 (N_5329,N_3797,N_4437);
and U5330 (N_5330,N_3843,N_3933);
xnor U5331 (N_5331,N_3663,N_3354);
or U5332 (N_5332,N_4243,N_4042);
nand U5333 (N_5333,N_3131,N_3082);
and U5334 (N_5334,N_4168,N_3289);
or U5335 (N_5335,N_3815,N_3074);
and U5336 (N_5336,N_3967,N_3568);
xor U5337 (N_5337,N_4125,N_4154);
xor U5338 (N_5338,N_4470,N_4257);
or U5339 (N_5339,N_4132,N_3603);
nand U5340 (N_5340,N_3755,N_4332);
nor U5341 (N_5341,N_4227,N_3399);
nand U5342 (N_5342,N_4013,N_3724);
and U5343 (N_5343,N_4366,N_4492);
xnor U5344 (N_5344,N_3103,N_3208);
nand U5345 (N_5345,N_3209,N_3368);
xor U5346 (N_5346,N_4194,N_3430);
nor U5347 (N_5347,N_4281,N_3670);
or U5348 (N_5348,N_3846,N_3614);
nand U5349 (N_5349,N_4157,N_3212);
and U5350 (N_5350,N_4342,N_3562);
xnor U5351 (N_5351,N_4102,N_3986);
nor U5352 (N_5352,N_3183,N_3123);
or U5353 (N_5353,N_3751,N_4419);
xor U5354 (N_5354,N_4410,N_3089);
or U5355 (N_5355,N_4406,N_3192);
or U5356 (N_5356,N_3594,N_3164);
and U5357 (N_5357,N_3546,N_4279);
nor U5358 (N_5358,N_3202,N_3983);
nand U5359 (N_5359,N_4411,N_3317);
nand U5360 (N_5360,N_4276,N_3191);
nand U5361 (N_5361,N_4347,N_3603);
nand U5362 (N_5362,N_3800,N_3526);
or U5363 (N_5363,N_4290,N_4497);
nand U5364 (N_5364,N_4196,N_3904);
or U5365 (N_5365,N_4414,N_3036);
xnor U5366 (N_5366,N_3891,N_3648);
or U5367 (N_5367,N_3199,N_4489);
xnor U5368 (N_5368,N_4052,N_4161);
nor U5369 (N_5369,N_3742,N_3100);
and U5370 (N_5370,N_4093,N_4404);
nor U5371 (N_5371,N_3603,N_3388);
nor U5372 (N_5372,N_3887,N_3805);
nor U5373 (N_5373,N_3449,N_3469);
or U5374 (N_5374,N_4464,N_3100);
nor U5375 (N_5375,N_4393,N_3159);
nor U5376 (N_5376,N_4488,N_4118);
nand U5377 (N_5377,N_3986,N_4411);
nand U5378 (N_5378,N_3148,N_4417);
and U5379 (N_5379,N_3464,N_3690);
xnor U5380 (N_5380,N_3374,N_3173);
nor U5381 (N_5381,N_4228,N_3170);
nand U5382 (N_5382,N_4378,N_4166);
xnor U5383 (N_5383,N_3626,N_4130);
nand U5384 (N_5384,N_4235,N_3739);
xnor U5385 (N_5385,N_4233,N_3037);
xnor U5386 (N_5386,N_3622,N_3157);
xnor U5387 (N_5387,N_3448,N_4013);
nor U5388 (N_5388,N_3810,N_3718);
nor U5389 (N_5389,N_3974,N_3156);
or U5390 (N_5390,N_3143,N_4485);
and U5391 (N_5391,N_3300,N_3247);
nand U5392 (N_5392,N_4413,N_3414);
or U5393 (N_5393,N_4126,N_3257);
or U5394 (N_5394,N_3027,N_3444);
nor U5395 (N_5395,N_4059,N_3023);
and U5396 (N_5396,N_3335,N_4412);
and U5397 (N_5397,N_4275,N_3990);
xor U5398 (N_5398,N_3596,N_4063);
and U5399 (N_5399,N_4068,N_4381);
or U5400 (N_5400,N_3575,N_3453);
nand U5401 (N_5401,N_4028,N_4027);
or U5402 (N_5402,N_3195,N_3506);
and U5403 (N_5403,N_3139,N_3328);
or U5404 (N_5404,N_3803,N_3798);
or U5405 (N_5405,N_3819,N_4051);
nand U5406 (N_5406,N_3511,N_3811);
xor U5407 (N_5407,N_4189,N_3328);
and U5408 (N_5408,N_3322,N_3106);
and U5409 (N_5409,N_3311,N_4157);
or U5410 (N_5410,N_4182,N_3627);
or U5411 (N_5411,N_3383,N_3666);
xnor U5412 (N_5412,N_3262,N_3623);
nor U5413 (N_5413,N_4132,N_3195);
nor U5414 (N_5414,N_4456,N_3454);
nor U5415 (N_5415,N_4436,N_4221);
and U5416 (N_5416,N_3261,N_3165);
and U5417 (N_5417,N_3188,N_3433);
or U5418 (N_5418,N_3082,N_4227);
or U5419 (N_5419,N_3818,N_3628);
or U5420 (N_5420,N_3719,N_3243);
or U5421 (N_5421,N_3586,N_3380);
xnor U5422 (N_5422,N_3490,N_3288);
nor U5423 (N_5423,N_3500,N_3235);
nand U5424 (N_5424,N_3525,N_3798);
or U5425 (N_5425,N_4005,N_3563);
or U5426 (N_5426,N_3899,N_4198);
or U5427 (N_5427,N_3663,N_3928);
nor U5428 (N_5428,N_4425,N_3037);
nand U5429 (N_5429,N_4236,N_4451);
or U5430 (N_5430,N_3112,N_4485);
or U5431 (N_5431,N_3989,N_3535);
xor U5432 (N_5432,N_3335,N_3174);
xor U5433 (N_5433,N_3941,N_3648);
or U5434 (N_5434,N_3660,N_4206);
nand U5435 (N_5435,N_3713,N_4382);
nor U5436 (N_5436,N_3119,N_3603);
nor U5437 (N_5437,N_4499,N_4455);
and U5438 (N_5438,N_3981,N_3740);
and U5439 (N_5439,N_3495,N_3823);
xor U5440 (N_5440,N_4169,N_3723);
xnor U5441 (N_5441,N_3293,N_3070);
or U5442 (N_5442,N_3415,N_4494);
nor U5443 (N_5443,N_3967,N_3407);
nor U5444 (N_5444,N_4281,N_4042);
or U5445 (N_5445,N_4077,N_3448);
nor U5446 (N_5446,N_3473,N_4475);
nand U5447 (N_5447,N_4050,N_3580);
xor U5448 (N_5448,N_3126,N_3925);
nand U5449 (N_5449,N_4196,N_3430);
and U5450 (N_5450,N_3245,N_4337);
nand U5451 (N_5451,N_4236,N_4074);
xnor U5452 (N_5452,N_3433,N_3061);
xor U5453 (N_5453,N_3481,N_3910);
and U5454 (N_5454,N_3885,N_3558);
xor U5455 (N_5455,N_3274,N_3618);
and U5456 (N_5456,N_4467,N_3067);
xnor U5457 (N_5457,N_3490,N_3891);
and U5458 (N_5458,N_3459,N_3154);
or U5459 (N_5459,N_4195,N_3664);
nand U5460 (N_5460,N_4468,N_4384);
nand U5461 (N_5461,N_3733,N_3394);
and U5462 (N_5462,N_3386,N_4039);
and U5463 (N_5463,N_3183,N_3215);
and U5464 (N_5464,N_3503,N_3996);
or U5465 (N_5465,N_4399,N_4494);
or U5466 (N_5466,N_4355,N_3742);
nor U5467 (N_5467,N_3813,N_3169);
xor U5468 (N_5468,N_3929,N_3473);
or U5469 (N_5469,N_3262,N_4070);
nor U5470 (N_5470,N_3771,N_4100);
or U5471 (N_5471,N_4053,N_3580);
nor U5472 (N_5472,N_4429,N_4289);
nor U5473 (N_5473,N_3457,N_3493);
nand U5474 (N_5474,N_3914,N_4204);
nand U5475 (N_5475,N_3847,N_3033);
nor U5476 (N_5476,N_4495,N_3337);
or U5477 (N_5477,N_4406,N_4165);
nor U5478 (N_5478,N_3434,N_4243);
nand U5479 (N_5479,N_4468,N_3082);
nor U5480 (N_5480,N_3674,N_3220);
or U5481 (N_5481,N_3545,N_4210);
and U5482 (N_5482,N_3840,N_3676);
nor U5483 (N_5483,N_4441,N_4244);
nand U5484 (N_5484,N_4000,N_3695);
or U5485 (N_5485,N_4079,N_4441);
nor U5486 (N_5486,N_4444,N_4412);
nand U5487 (N_5487,N_3472,N_4434);
nand U5488 (N_5488,N_3983,N_3087);
xor U5489 (N_5489,N_3414,N_3741);
or U5490 (N_5490,N_3561,N_4108);
or U5491 (N_5491,N_3628,N_3253);
and U5492 (N_5492,N_3983,N_3280);
xor U5493 (N_5493,N_3786,N_4451);
and U5494 (N_5494,N_3777,N_3295);
or U5495 (N_5495,N_3376,N_4363);
and U5496 (N_5496,N_3911,N_4069);
or U5497 (N_5497,N_3562,N_3973);
xnor U5498 (N_5498,N_3062,N_4405);
or U5499 (N_5499,N_3310,N_4202);
xnor U5500 (N_5500,N_3133,N_3851);
xnor U5501 (N_5501,N_3811,N_3895);
and U5502 (N_5502,N_4017,N_3500);
and U5503 (N_5503,N_4073,N_3291);
nand U5504 (N_5504,N_3500,N_3913);
nor U5505 (N_5505,N_3895,N_4146);
or U5506 (N_5506,N_3054,N_3248);
or U5507 (N_5507,N_4472,N_4134);
xor U5508 (N_5508,N_4182,N_3550);
nor U5509 (N_5509,N_3714,N_3788);
nand U5510 (N_5510,N_3430,N_4267);
or U5511 (N_5511,N_3538,N_4253);
and U5512 (N_5512,N_3034,N_4395);
or U5513 (N_5513,N_4324,N_4055);
nor U5514 (N_5514,N_3441,N_3537);
xnor U5515 (N_5515,N_4416,N_3790);
nand U5516 (N_5516,N_4105,N_3187);
nor U5517 (N_5517,N_3950,N_4300);
and U5518 (N_5518,N_4250,N_4295);
and U5519 (N_5519,N_3887,N_3797);
nor U5520 (N_5520,N_4003,N_4145);
nand U5521 (N_5521,N_4208,N_3113);
nand U5522 (N_5522,N_3133,N_3173);
or U5523 (N_5523,N_3273,N_3134);
nand U5524 (N_5524,N_3957,N_4443);
or U5525 (N_5525,N_3618,N_3354);
nand U5526 (N_5526,N_4310,N_3877);
xnor U5527 (N_5527,N_3966,N_3810);
or U5528 (N_5528,N_4075,N_3100);
or U5529 (N_5529,N_4084,N_3423);
nor U5530 (N_5530,N_4134,N_4284);
or U5531 (N_5531,N_3624,N_3259);
and U5532 (N_5532,N_3967,N_3211);
or U5533 (N_5533,N_4313,N_4251);
nand U5534 (N_5534,N_3819,N_3727);
nand U5535 (N_5535,N_3629,N_4405);
or U5536 (N_5536,N_3669,N_4358);
nor U5537 (N_5537,N_3114,N_4471);
and U5538 (N_5538,N_3564,N_4050);
or U5539 (N_5539,N_3449,N_3242);
xor U5540 (N_5540,N_3039,N_3960);
and U5541 (N_5541,N_4145,N_3409);
nor U5542 (N_5542,N_4017,N_3483);
or U5543 (N_5543,N_3862,N_3551);
nor U5544 (N_5544,N_3047,N_3343);
or U5545 (N_5545,N_4150,N_3546);
nand U5546 (N_5546,N_3243,N_3167);
nor U5547 (N_5547,N_3147,N_3558);
and U5548 (N_5548,N_3672,N_3650);
nand U5549 (N_5549,N_3063,N_3230);
nor U5550 (N_5550,N_3778,N_4364);
nand U5551 (N_5551,N_3030,N_3569);
nand U5552 (N_5552,N_3454,N_4375);
nor U5553 (N_5553,N_3861,N_3060);
and U5554 (N_5554,N_3819,N_3222);
nor U5555 (N_5555,N_3308,N_4486);
xnor U5556 (N_5556,N_3863,N_4145);
nor U5557 (N_5557,N_3682,N_3846);
xor U5558 (N_5558,N_4304,N_4046);
xnor U5559 (N_5559,N_4048,N_4122);
or U5560 (N_5560,N_4130,N_3983);
or U5561 (N_5561,N_3037,N_3751);
nor U5562 (N_5562,N_3749,N_3478);
xor U5563 (N_5563,N_3950,N_3164);
and U5564 (N_5564,N_3713,N_3564);
xnor U5565 (N_5565,N_4311,N_4392);
nand U5566 (N_5566,N_4108,N_4008);
nor U5567 (N_5567,N_4180,N_3804);
and U5568 (N_5568,N_3721,N_3075);
nand U5569 (N_5569,N_3396,N_4311);
nand U5570 (N_5570,N_4297,N_4409);
xnor U5571 (N_5571,N_3502,N_3280);
nand U5572 (N_5572,N_4100,N_3036);
and U5573 (N_5573,N_3492,N_3400);
xnor U5574 (N_5574,N_3264,N_3652);
nor U5575 (N_5575,N_3559,N_3023);
nor U5576 (N_5576,N_3015,N_3831);
xnor U5577 (N_5577,N_3044,N_3783);
or U5578 (N_5578,N_3028,N_3658);
xor U5579 (N_5579,N_3788,N_4290);
or U5580 (N_5580,N_3749,N_3519);
nor U5581 (N_5581,N_3731,N_4137);
nand U5582 (N_5582,N_3647,N_4183);
and U5583 (N_5583,N_3558,N_3699);
xnor U5584 (N_5584,N_3132,N_3497);
or U5585 (N_5585,N_3845,N_4229);
nand U5586 (N_5586,N_4400,N_3766);
and U5587 (N_5587,N_3956,N_3690);
xor U5588 (N_5588,N_3170,N_4221);
or U5589 (N_5589,N_3219,N_3803);
xor U5590 (N_5590,N_3540,N_3860);
nor U5591 (N_5591,N_3473,N_3573);
and U5592 (N_5592,N_3869,N_4004);
and U5593 (N_5593,N_3881,N_3078);
or U5594 (N_5594,N_3456,N_3800);
nor U5595 (N_5595,N_3680,N_3186);
nor U5596 (N_5596,N_3280,N_3731);
nor U5597 (N_5597,N_3574,N_3071);
nand U5598 (N_5598,N_3777,N_3472);
xor U5599 (N_5599,N_3262,N_4173);
nand U5600 (N_5600,N_3071,N_4389);
nand U5601 (N_5601,N_4073,N_3972);
nand U5602 (N_5602,N_3577,N_4288);
and U5603 (N_5603,N_3284,N_3383);
or U5604 (N_5604,N_3906,N_3241);
nand U5605 (N_5605,N_4013,N_3286);
xor U5606 (N_5606,N_3954,N_3996);
and U5607 (N_5607,N_4498,N_3943);
nor U5608 (N_5608,N_3233,N_4072);
xnor U5609 (N_5609,N_3782,N_3762);
nand U5610 (N_5610,N_3165,N_3331);
and U5611 (N_5611,N_3088,N_4261);
and U5612 (N_5612,N_4074,N_3041);
and U5613 (N_5613,N_3086,N_4269);
xor U5614 (N_5614,N_3600,N_3768);
nand U5615 (N_5615,N_4371,N_3146);
and U5616 (N_5616,N_3550,N_3553);
nor U5617 (N_5617,N_3365,N_3138);
nand U5618 (N_5618,N_3835,N_3527);
nand U5619 (N_5619,N_3649,N_4473);
nor U5620 (N_5620,N_3903,N_4337);
and U5621 (N_5621,N_3429,N_4216);
nor U5622 (N_5622,N_3519,N_3871);
or U5623 (N_5623,N_3932,N_3452);
and U5624 (N_5624,N_4061,N_4142);
xor U5625 (N_5625,N_3443,N_3988);
nor U5626 (N_5626,N_3244,N_3598);
xnor U5627 (N_5627,N_3126,N_3936);
nand U5628 (N_5628,N_3535,N_3137);
xnor U5629 (N_5629,N_3381,N_4008);
nand U5630 (N_5630,N_4451,N_3095);
nand U5631 (N_5631,N_4367,N_3737);
xor U5632 (N_5632,N_4032,N_3560);
or U5633 (N_5633,N_4185,N_4407);
nor U5634 (N_5634,N_3814,N_3209);
nand U5635 (N_5635,N_4333,N_3144);
nand U5636 (N_5636,N_3309,N_3261);
or U5637 (N_5637,N_3182,N_3776);
and U5638 (N_5638,N_4160,N_4303);
nor U5639 (N_5639,N_3153,N_3257);
nor U5640 (N_5640,N_3336,N_3440);
nor U5641 (N_5641,N_3860,N_4446);
nand U5642 (N_5642,N_3250,N_3427);
or U5643 (N_5643,N_4431,N_4420);
nor U5644 (N_5644,N_4085,N_4132);
or U5645 (N_5645,N_4070,N_4318);
nor U5646 (N_5646,N_4202,N_3610);
or U5647 (N_5647,N_3285,N_3980);
nor U5648 (N_5648,N_3377,N_3846);
nand U5649 (N_5649,N_4103,N_4117);
or U5650 (N_5650,N_3026,N_3336);
and U5651 (N_5651,N_4004,N_3978);
and U5652 (N_5652,N_3785,N_3243);
xor U5653 (N_5653,N_3253,N_3487);
xor U5654 (N_5654,N_4285,N_3930);
or U5655 (N_5655,N_3233,N_3099);
or U5656 (N_5656,N_3380,N_3370);
or U5657 (N_5657,N_4118,N_3105);
nor U5658 (N_5658,N_3224,N_4097);
xnor U5659 (N_5659,N_4489,N_4457);
nor U5660 (N_5660,N_3583,N_3458);
nor U5661 (N_5661,N_4203,N_4379);
and U5662 (N_5662,N_3632,N_3008);
or U5663 (N_5663,N_3621,N_3128);
xor U5664 (N_5664,N_3257,N_3334);
nand U5665 (N_5665,N_3103,N_3310);
or U5666 (N_5666,N_3763,N_3735);
and U5667 (N_5667,N_3323,N_3043);
nor U5668 (N_5668,N_3070,N_4270);
or U5669 (N_5669,N_4400,N_4453);
nor U5670 (N_5670,N_4182,N_3826);
nor U5671 (N_5671,N_4451,N_4145);
nand U5672 (N_5672,N_3745,N_3811);
or U5673 (N_5673,N_3491,N_4363);
nor U5674 (N_5674,N_3715,N_4102);
and U5675 (N_5675,N_4135,N_4262);
or U5676 (N_5676,N_4011,N_3530);
and U5677 (N_5677,N_3412,N_3674);
or U5678 (N_5678,N_4204,N_3286);
xnor U5679 (N_5679,N_3086,N_3432);
and U5680 (N_5680,N_3433,N_3772);
xor U5681 (N_5681,N_3221,N_3684);
nand U5682 (N_5682,N_3461,N_4059);
nand U5683 (N_5683,N_3356,N_4193);
xnor U5684 (N_5684,N_3931,N_4160);
and U5685 (N_5685,N_3480,N_4473);
nor U5686 (N_5686,N_4110,N_3794);
or U5687 (N_5687,N_3363,N_3653);
xor U5688 (N_5688,N_3938,N_3198);
nor U5689 (N_5689,N_3835,N_3908);
or U5690 (N_5690,N_4015,N_3839);
nor U5691 (N_5691,N_3841,N_3380);
or U5692 (N_5692,N_3584,N_3697);
nor U5693 (N_5693,N_4114,N_4371);
nor U5694 (N_5694,N_3141,N_3925);
nand U5695 (N_5695,N_3797,N_3342);
xnor U5696 (N_5696,N_3774,N_3827);
nor U5697 (N_5697,N_4153,N_3609);
or U5698 (N_5698,N_4301,N_3499);
xnor U5699 (N_5699,N_3661,N_3784);
or U5700 (N_5700,N_4487,N_3943);
nor U5701 (N_5701,N_3362,N_4305);
nor U5702 (N_5702,N_3001,N_3968);
or U5703 (N_5703,N_3815,N_4307);
and U5704 (N_5704,N_4107,N_3367);
or U5705 (N_5705,N_3187,N_3132);
nor U5706 (N_5706,N_4016,N_4092);
xnor U5707 (N_5707,N_3265,N_3676);
nor U5708 (N_5708,N_3092,N_3993);
and U5709 (N_5709,N_4373,N_4169);
xor U5710 (N_5710,N_3168,N_3511);
xor U5711 (N_5711,N_3090,N_3801);
xnor U5712 (N_5712,N_4046,N_3538);
nand U5713 (N_5713,N_4375,N_3950);
nand U5714 (N_5714,N_3401,N_4464);
and U5715 (N_5715,N_3352,N_3327);
or U5716 (N_5716,N_3111,N_4403);
nand U5717 (N_5717,N_4076,N_4053);
or U5718 (N_5718,N_3036,N_3359);
xor U5719 (N_5719,N_4451,N_4212);
nor U5720 (N_5720,N_3486,N_3576);
nor U5721 (N_5721,N_3722,N_3468);
and U5722 (N_5722,N_4177,N_3180);
xnor U5723 (N_5723,N_3716,N_4233);
nor U5724 (N_5724,N_3719,N_3060);
nand U5725 (N_5725,N_4181,N_3847);
or U5726 (N_5726,N_4095,N_3741);
or U5727 (N_5727,N_3261,N_4149);
nand U5728 (N_5728,N_3479,N_3648);
nor U5729 (N_5729,N_3926,N_3058);
and U5730 (N_5730,N_3270,N_3444);
and U5731 (N_5731,N_4141,N_4280);
or U5732 (N_5732,N_3056,N_3266);
xor U5733 (N_5733,N_4041,N_4096);
and U5734 (N_5734,N_3861,N_4471);
xnor U5735 (N_5735,N_3665,N_3935);
or U5736 (N_5736,N_3829,N_3302);
or U5737 (N_5737,N_3235,N_3949);
nand U5738 (N_5738,N_3952,N_3065);
nand U5739 (N_5739,N_3695,N_3848);
nor U5740 (N_5740,N_3489,N_3625);
xnor U5741 (N_5741,N_3478,N_4342);
nor U5742 (N_5742,N_3245,N_3090);
xor U5743 (N_5743,N_3708,N_3470);
and U5744 (N_5744,N_4227,N_4329);
nand U5745 (N_5745,N_3941,N_3436);
xor U5746 (N_5746,N_3007,N_4247);
nand U5747 (N_5747,N_4156,N_4116);
and U5748 (N_5748,N_3759,N_3539);
xnor U5749 (N_5749,N_4497,N_3753);
and U5750 (N_5750,N_3905,N_3808);
xnor U5751 (N_5751,N_3988,N_3805);
and U5752 (N_5752,N_3771,N_3863);
and U5753 (N_5753,N_4028,N_4425);
and U5754 (N_5754,N_3194,N_3558);
xor U5755 (N_5755,N_4233,N_3156);
xnor U5756 (N_5756,N_3599,N_3011);
nand U5757 (N_5757,N_3624,N_4455);
nand U5758 (N_5758,N_3751,N_3573);
nor U5759 (N_5759,N_3654,N_4162);
nor U5760 (N_5760,N_4435,N_3610);
nor U5761 (N_5761,N_3932,N_3945);
and U5762 (N_5762,N_4495,N_3411);
nand U5763 (N_5763,N_3861,N_3287);
xor U5764 (N_5764,N_3699,N_3507);
nand U5765 (N_5765,N_3552,N_3104);
xnor U5766 (N_5766,N_3660,N_4036);
nand U5767 (N_5767,N_3474,N_3631);
nand U5768 (N_5768,N_3228,N_3691);
nand U5769 (N_5769,N_3888,N_3411);
or U5770 (N_5770,N_3158,N_3705);
nand U5771 (N_5771,N_3151,N_3920);
nor U5772 (N_5772,N_3774,N_4107);
and U5773 (N_5773,N_4101,N_3358);
and U5774 (N_5774,N_3908,N_3507);
and U5775 (N_5775,N_4344,N_3129);
or U5776 (N_5776,N_3045,N_4342);
nand U5777 (N_5777,N_4409,N_4327);
or U5778 (N_5778,N_3234,N_3002);
nor U5779 (N_5779,N_3311,N_3752);
xor U5780 (N_5780,N_3681,N_3981);
or U5781 (N_5781,N_3692,N_3305);
and U5782 (N_5782,N_4344,N_3861);
xor U5783 (N_5783,N_4354,N_4418);
nor U5784 (N_5784,N_3655,N_3795);
and U5785 (N_5785,N_3986,N_3071);
and U5786 (N_5786,N_3468,N_4421);
nor U5787 (N_5787,N_3513,N_3494);
nand U5788 (N_5788,N_3606,N_3279);
nand U5789 (N_5789,N_3202,N_3966);
nor U5790 (N_5790,N_3035,N_4115);
xnor U5791 (N_5791,N_4375,N_4274);
and U5792 (N_5792,N_4156,N_4404);
xnor U5793 (N_5793,N_4061,N_4475);
xor U5794 (N_5794,N_3028,N_3293);
xor U5795 (N_5795,N_3086,N_3169);
xor U5796 (N_5796,N_3989,N_3322);
or U5797 (N_5797,N_3112,N_4284);
xnor U5798 (N_5798,N_3225,N_3029);
and U5799 (N_5799,N_4311,N_3850);
or U5800 (N_5800,N_3809,N_3928);
or U5801 (N_5801,N_3171,N_3136);
and U5802 (N_5802,N_3388,N_3369);
nor U5803 (N_5803,N_4289,N_4466);
nor U5804 (N_5804,N_3677,N_4330);
nor U5805 (N_5805,N_4058,N_4165);
and U5806 (N_5806,N_4479,N_3664);
nor U5807 (N_5807,N_4472,N_3958);
xor U5808 (N_5808,N_3613,N_4050);
nand U5809 (N_5809,N_4200,N_4381);
nand U5810 (N_5810,N_3539,N_3974);
and U5811 (N_5811,N_3025,N_3900);
nor U5812 (N_5812,N_3602,N_3119);
nand U5813 (N_5813,N_3366,N_3506);
or U5814 (N_5814,N_3314,N_3215);
nor U5815 (N_5815,N_4336,N_3404);
xor U5816 (N_5816,N_3190,N_4219);
xnor U5817 (N_5817,N_4129,N_3805);
and U5818 (N_5818,N_3871,N_3334);
and U5819 (N_5819,N_4054,N_4126);
nand U5820 (N_5820,N_4345,N_3767);
nand U5821 (N_5821,N_3573,N_3532);
or U5822 (N_5822,N_3099,N_3208);
and U5823 (N_5823,N_3832,N_3006);
nand U5824 (N_5824,N_3898,N_4326);
xnor U5825 (N_5825,N_4204,N_3474);
or U5826 (N_5826,N_3957,N_4190);
xnor U5827 (N_5827,N_3410,N_3330);
nor U5828 (N_5828,N_3601,N_3993);
nor U5829 (N_5829,N_3088,N_3031);
nor U5830 (N_5830,N_3865,N_3070);
nand U5831 (N_5831,N_3358,N_4005);
and U5832 (N_5832,N_4011,N_3992);
xnor U5833 (N_5833,N_3028,N_3006);
xnor U5834 (N_5834,N_3842,N_4014);
nor U5835 (N_5835,N_3875,N_3409);
nand U5836 (N_5836,N_3192,N_3056);
or U5837 (N_5837,N_4498,N_3551);
nand U5838 (N_5838,N_3930,N_3495);
xor U5839 (N_5839,N_4059,N_3534);
nor U5840 (N_5840,N_3412,N_3208);
xnor U5841 (N_5841,N_3431,N_3182);
xnor U5842 (N_5842,N_4365,N_4444);
and U5843 (N_5843,N_3970,N_3189);
or U5844 (N_5844,N_4107,N_4263);
or U5845 (N_5845,N_3508,N_3559);
or U5846 (N_5846,N_3065,N_3343);
nor U5847 (N_5847,N_3595,N_3645);
and U5848 (N_5848,N_3398,N_3979);
and U5849 (N_5849,N_4282,N_3829);
nand U5850 (N_5850,N_4008,N_4360);
xnor U5851 (N_5851,N_4249,N_4217);
nor U5852 (N_5852,N_3809,N_3084);
nand U5853 (N_5853,N_4469,N_3525);
and U5854 (N_5854,N_3518,N_3280);
xor U5855 (N_5855,N_4448,N_4379);
xnor U5856 (N_5856,N_4171,N_3509);
nand U5857 (N_5857,N_3679,N_3610);
nor U5858 (N_5858,N_4108,N_4063);
xor U5859 (N_5859,N_3562,N_3040);
xor U5860 (N_5860,N_3887,N_4170);
xnor U5861 (N_5861,N_3730,N_3661);
xor U5862 (N_5862,N_3478,N_3381);
nor U5863 (N_5863,N_3774,N_3797);
xor U5864 (N_5864,N_3050,N_4089);
nor U5865 (N_5865,N_3328,N_3216);
xor U5866 (N_5866,N_3757,N_4489);
and U5867 (N_5867,N_3856,N_3298);
xnor U5868 (N_5868,N_3167,N_3409);
and U5869 (N_5869,N_3365,N_3855);
xor U5870 (N_5870,N_3064,N_3432);
or U5871 (N_5871,N_3207,N_3372);
xnor U5872 (N_5872,N_4235,N_4345);
nand U5873 (N_5873,N_3940,N_4201);
or U5874 (N_5874,N_3567,N_3540);
nand U5875 (N_5875,N_3837,N_4053);
or U5876 (N_5876,N_3752,N_4140);
nor U5877 (N_5877,N_4194,N_3678);
or U5878 (N_5878,N_3008,N_3535);
nor U5879 (N_5879,N_4040,N_4131);
or U5880 (N_5880,N_3706,N_3157);
xnor U5881 (N_5881,N_4171,N_3536);
or U5882 (N_5882,N_3993,N_3687);
nand U5883 (N_5883,N_3746,N_3991);
or U5884 (N_5884,N_3776,N_3868);
and U5885 (N_5885,N_3295,N_3676);
or U5886 (N_5886,N_3440,N_3285);
xnor U5887 (N_5887,N_3470,N_3431);
xor U5888 (N_5888,N_4182,N_4439);
nand U5889 (N_5889,N_3004,N_3469);
or U5890 (N_5890,N_4067,N_3422);
xor U5891 (N_5891,N_3605,N_3602);
nand U5892 (N_5892,N_4234,N_3499);
nor U5893 (N_5893,N_4125,N_3377);
xor U5894 (N_5894,N_4168,N_3148);
nor U5895 (N_5895,N_3116,N_3197);
and U5896 (N_5896,N_3179,N_4314);
xnor U5897 (N_5897,N_4195,N_4071);
nand U5898 (N_5898,N_3451,N_4483);
xor U5899 (N_5899,N_4058,N_4200);
xor U5900 (N_5900,N_3968,N_4357);
nor U5901 (N_5901,N_3565,N_3065);
and U5902 (N_5902,N_3213,N_4088);
or U5903 (N_5903,N_4159,N_3038);
and U5904 (N_5904,N_3722,N_3872);
nor U5905 (N_5905,N_3420,N_3162);
and U5906 (N_5906,N_3244,N_3187);
nor U5907 (N_5907,N_4466,N_3234);
or U5908 (N_5908,N_3992,N_4401);
or U5909 (N_5909,N_3748,N_3031);
or U5910 (N_5910,N_3561,N_3198);
xor U5911 (N_5911,N_3753,N_3170);
nor U5912 (N_5912,N_3450,N_3919);
nand U5913 (N_5913,N_3318,N_3225);
or U5914 (N_5914,N_3982,N_3190);
or U5915 (N_5915,N_4149,N_3482);
xor U5916 (N_5916,N_3267,N_3875);
or U5917 (N_5917,N_3607,N_3477);
xnor U5918 (N_5918,N_4389,N_3316);
and U5919 (N_5919,N_4019,N_4071);
xor U5920 (N_5920,N_3959,N_4452);
nand U5921 (N_5921,N_3301,N_4263);
nor U5922 (N_5922,N_4442,N_3142);
and U5923 (N_5923,N_3708,N_3519);
nor U5924 (N_5924,N_4482,N_3333);
or U5925 (N_5925,N_4136,N_3824);
and U5926 (N_5926,N_3832,N_4257);
nor U5927 (N_5927,N_4116,N_3773);
nand U5928 (N_5928,N_3666,N_3977);
and U5929 (N_5929,N_3871,N_3052);
nor U5930 (N_5930,N_4439,N_3202);
or U5931 (N_5931,N_3519,N_3807);
and U5932 (N_5932,N_3154,N_3942);
and U5933 (N_5933,N_3530,N_3367);
nand U5934 (N_5934,N_3196,N_3043);
and U5935 (N_5935,N_3922,N_3260);
and U5936 (N_5936,N_4009,N_3459);
or U5937 (N_5937,N_4295,N_3865);
xnor U5938 (N_5938,N_3402,N_3155);
or U5939 (N_5939,N_3017,N_4356);
or U5940 (N_5940,N_3638,N_3143);
nor U5941 (N_5941,N_3614,N_3092);
nor U5942 (N_5942,N_4289,N_3760);
and U5943 (N_5943,N_3471,N_3314);
nand U5944 (N_5944,N_4198,N_4475);
and U5945 (N_5945,N_3307,N_3717);
nand U5946 (N_5946,N_3960,N_4486);
xor U5947 (N_5947,N_4110,N_3739);
nor U5948 (N_5948,N_4061,N_4476);
or U5949 (N_5949,N_3022,N_4160);
xnor U5950 (N_5950,N_3190,N_4232);
or U5951 (N_5951,N_3076,N_3260);
or U5952 (N_5952,N_3429,N_3005);
nor U5953 (N_5953,N_4340,N_3747);
nor U5954 (N_5954,N_4395,N_3283);
xor U5955 (N_5955,N_3189,N_3938);
nor U5956 (N_5956,N_3177,N_3904);
or U5957 (N_5957,N_3567,N_3429);
xor U5958 (N_5958,N_3724,N_3006);
or U5959 (N_5959,N_4172,N_3019);
and U5960 (N_5960,N_3043,N_4235);
nor U5961 (N_5961,N_3788,N_4411);
nand U5962 (N_5962,N_3899,N_3690);
nand U5963 (N_5963,N_4419,N_4297);
and U5964 (N_5964,N_3674,N_3177);
xor U5965 (N_5965,N_3749,N_3251);
xor U5966 (N_5966,N_3011,N_4255);
nor U5967 (N_5967,N_3217,N_4304);
and U5968 (N_5968,N_3324,N_4325);
and U5969 (N_5969,N_3080,N_3803);
nand U5970 (N_5970,N_3498,N_3335);
nor U5971 (N_5971,N_4493,N_3606);
and U5972 (N_5972,N_3611,N_3317);
nor U5973 (N_5973,N_4288,N_3719);
or U5974 (N_5974,N_3253,N_4450);
xnor U5975 (N_5975,N_3669,N_4190);
nand U5976 (N_5976,N_4114,N_3318);
nand U5977 (N_5977,N_3905,N_4088);
or U5978 (N_5978,N_4192,N_3118);
xnor U5979 (N_5979,N_3072,N_4323);
nor U5980 (N_5980,N_4352,N_4021);
or U5981 (N_5981,N_3852,N_3830);
or U5982 (N_5982,N_3248,N_3600);
xnor U5983 (N_5983,N_3445,N_3952);
xnor U5984 (N_5984,N_4258,N_3624);
and U5985 (N_5985,N_3068,N_3108);
and U5986 (N_5986,N_4212,N_3980);
nor U5987 (N_5987,N_4115,N_3011);
and U5988 (N_5988,N_3611,N_3928);
or U5989 (N_5989,N_4314,N_4085);
nand U5990 (N_5990,N_3740,N_3629);
nand U5991 (N_5991,N_3489,N_3266);
and U5992 (N_5992,N_4479,N_3085);
or U5993 (N_5993,N_3787,N_3340);
nand U5994 (N_5994,N_3359,N_3465);
nand U5995 (N_5995,N_3290,N_3783);
and U5996 (N_5996,N_4438,N_3427);
xnor U5997 (N_5997,N_3380,N_4466);
and U5998 (N_5998,N_3533,N_4351);
or U5999 (N_5999,N_3072,N_3078);
nand U6000 (N_6000,N_5785,N_5735);
or U6001 (N_6001,N_4647,N_5061);
nand U6002 (N_6002,N_4854,N_5127);
xor U6003 (N_6003,N_5264,N_4875);
and U6004 (N_6004,N_5553,N_4994);
nand U6005 (N_6005,N_5611,N_5604);
or U6006 (N_6006,N_4701,N_5521);
or U6007 (N_6007,N_5269,N_5856);
xor U6008 (N_6008,N_5834,N_5290);
nand U6009 (N_6009,N_5598,N_5453);
xor U6010 (N_6010,N_5627,N_4956);
xnor U6011 (N_6011,N_4954,N_5647);
nand U6012 (N_6012,N_4823,N_4680);
nand U6013 (N_6013,N_5010,N_4957);
nand U6014 (N_6014,N_4975,N_4991);
and U6015 (N_6015,N_5133,N_5748);
nand U6016 (N_6016,N_4818,N_4539);
xor U6017 (N_6017,N_5797,N_5169);
or U6018 (N_6018,N_5998,N_5761);
and U6019 (N_6019,N_5201,N_5937);
nor U6020 (N_6020,N_5380,N_4677);
xnor U6021 (N_6021,N_5630,N_5037);
nand U6022 (N_6022,N_4901,N_4766);
xor U6023 (N_6023,N_5221,N_5689);
xor U6024 (N_6024,N_4800,N_5915);
and U6025 (N_6025,N_5080,N_5138);
xnor U6026 (N_6026,N_5130,N_5445);
nand U6027 (N_6027,N_4576,N_4526);
nand U6028 (N_6028,N_4670,N_5111);
or U6029 (N_6029,N_4807,N_4682);
and U6030 (N_6030,N_5999,N_5395);
nor U6031 (N_6031,N_4684,N_5262);
and U6032 (N_6032,N_5979,N_5049);
and U6033 (N_6033,N_4761,N_4666);
and U6034 (N_6034,N_4903,N_5985);
xnor U6035 (N_6035,N_5824,N_5450);
and U6036 (N_6036,N_5289,N_4668);
xor U6037 (N_6037,N_5462,N_5978);
or U6038 (N_6038,N_4507,N_4639);
xor U6039 (N_6039,N_4780,N_5132);
or U6040 (N_6040,N_5219,N_4830);
or U6041 (N_6041,N_5688,N_5493);
nor U6042 (N_6042,N_4616,N_5782);
and U6043 (N_6043,N_5796,N_4972);
and U6044 (N_6044,N_5795,N_5114);
nor U6045 (N_6045,N_5715,N_5517);
nand U6046 (N_6046,N_5905,N_5973);
xor U6047 (N_6047,N_5586,N_5704);
and U6048 (N_6048,N_5644,N_5487);
xor U6049 (N_6049,N_5543,N_4727);
nand U6050 (N_6050,N_5960,N_5027);
or U6051 (N_6051,N_5123,N_5098);
and U6052 (N_6052,N_5591,N_5071);
or U6053 (N_6053,N_5803,N_5549);
and U6054 (N_6054,N_5966,N_5105);
nand U6055 (N_6055,N_5734,N_4650);
nor U6056 (N_6056,N_5435,N_4767);
or U6057 (N_6057,N_5267,N_4833);
xor U6058 (N_6058,N_5754,N_4998);
and U6059 (N_6059,N_4728,N_4795);
nor U6060 (N_6060,N_5452,N_5760);
nand U6061 (N_6061,N_4642,N_5697);
or U6062 (N_6062,N_5625,N_4527);
and U6063 (N_6063,N_5442,N_4814);
xor U6064 (N_6064,N_5636,N_5134);
nand U6065 (N_6065,N_5840,N_5188);
nor U6066 (N_6066,N_5850,N_4704);
nand U6067 (N_6067,N_4897,N_5342);
or U6068 (N_6068,N_4758,N_4588);
nand U6069 (N_6069,N_4581,N_4838);
xnor U6070 (N_6070,N_5990,N_5969);
or U6071 (N_6071,N_4669,N_5066);
nor U6072 (N_6072,N_4909,N_5436);
or U6073 (N_6073,N_5043,N_5000);
nand U6074 (N_6074,N_5397,N_5956);
and U6075 (N_6075,N_5573,N_4715);
nor U6076 (N_6076,N_4709,N_5512);
and U6077 (N_6077,N_5935,N_5524);
xnor U6078 (N_6078,N_5550,N_5365);
and U6079 (N_6079,N_4984,N_5038);
and U6080 (N_6080,N_4651,N_5145);
nand U6081 (N_6081,N_5428,N_4686);
or U6082 (N_6082,N_4683,N_5230);
and U6083 (N_6083,N_5379,N_4829);
nor U6084 (N_6084,N_5645,N_5884);
nor U6085 (N_6085,N_5535,N_5839);
xor U6086 (N_6086,N_5895,N_4628);
and U6087 (N_6087,N_5214,N_4648);
or U6088 (N_6088,N_5794,N_5314);
or U6089 (N_6089,N_5333,N_5941);
nand U6090 (N_6090,N_5412,N_5476);
or U6091 (N_6091,N_5605,N_5853);
nor U6092 (N_6092,N_5102,N_5638);
xnor U6093 (N_6093,N_5449,N_4571);
xor U6094 (N_6094,N_5507,N_5967);
and U6095 (N_6095,N_5073,N_4679);
xnor U6096 (N_6096,N_5680,N_5574);
and U6097 (N_6097,N_5974,N_5668);
xnor U6098 (N_6098,N_5921,N_5659);
or U6099 (N_6099,N_5648,N_5628);
nor U6100 (N_6100,N_5213,N_4926);
xnor U6101 (N_6101,N_5349,N_4876);
and U6102 (N_6102,N_4721,N_5654);
and U6103 (N_6103,N_5060,N_5153);
nor U6104 (N_6104,N_5196,N_5408);
nand U6105 (N_6105,N_5661,N_5238);
nand U6106 (N_6106,N_5887,N_5370);
and U6107 (N_6107,N_4938,N_5767);
and U6108 (N_6108,N_4963,N_4871);
nand U6109 (N_6109,N_5718,N_5396);
nand U6110 (N_6110,N_4586,N_5943);
nor U6111 (N_6111,N_5983,N_4643);
xor U6112 (N_6112,N_4617,N_5708);
and U6113 (N_6113,N_4621,N_4783);
or U6114 (N_6114,N_5013,N_5218);
and U6115 (N_6115,N_5866,N_4733);
nand U6116 (N_6116,N_5805,N_5809);
or U6117 (N_6117,N_5858,N_4890);
nor U6118 (N_6118,N_5835,N_4911);
xor U6119 (N_6119,N_5300,N_5276);
nor U6120 (N_6120,N_4810,N_5890);
or U6121 (N_6121,N_5723,N_4501);
or U6122 (N_6122,N_4511,N_4559);
nand U6123 (N_6123,N_5072,N_4781);
or U6124 (N_6124,N_5666,N_4675);
and U6125 (N_6125,N_5294,N_5144);
or U6126 (N_6126,N_5929,N_5922);
nor U6127 (N_6127,N_5670,N_5067);
and U6128 (N_6128,N_5828,N_5880);
or U6129 (N_6129,N_4646,N_5728);
nand U6130 (N_6130,N_5936,N_4777);
or U6131 (N_6131,N_4601,N_5411);
nor U6132 (N_6132,N_4562,N_4736);
or U6133 (N_6133,N_5950,N_5774);
nor U6134 (N_6134,N_5942,N_5240);
nor U6135 (N_6135,N_4512,N_4558);
nor U6136 (N_6136,N_4678,N_5810);
and U6137 (N_6137,N_4593,N_5414);
xor U6138 (N_6138,N_5808,N_4917);
or U6139 (N_6139,N_5237,N_5756);
nor U6140 (N_6140,N_4707,N_5933);
or U6141 (N_6141,N_5631,N_5567);
and U6142 (N_6142,N_4550,N_5815);
nand U6143 (N_6143,N_5348,N_5215);
nand U6144 (N_6144,N_5646,N_5456);
nor U6145 (N_6145,N_5617,N_4714);
nand U6146 (N_6146,N_4713,N_5802);
and U6147 (N_6147,N_4899,N_4751);
nor U6148 (N_6148,N_5945,N_5254);
and U6149 (N_6149,N_5372,N_5316);
and U6150 (N_6150,N_5062,N_5778);
xor U6151 (N_6151,N_5731,N_5451);
or U6152 (N_6152,N_5258,N_4960);
or U6153 (N_6153,N_4867,N_4735);
and U6154 (N_6154,N_5303,N_5773);
xnor U6155 (N_6155,N_5307,N_5635);
nor U6156 (N_6156,N_5168,N_5057);
xnor U6157 (N_6157,N_5200,N_4641);
or U6158 (N_6158,N_4773,N_5682);
nor U6159 (N_6159,N_5677,N_5902);
xnor U6160 (N_6160,N_5772,N_5336);
xnor U6161 (N_6161,N_5690,N_5226);
nor U6162 (N_6162,N_5674,N_5807);
and U6163 (N_6163,N_4824,N_5361);
or U6164 (N_6164,N_5755,N_5871);
or U6165 (N_6165,N_4573,N_4784);
or U6166 (N_6166,N_5992,N_5430);
nor U6167 (N_6167,N_5357,N_5404);
or U6168 (N_6168,N_5924,N_5693);
and U6169 (N_6169,N_5401,N_4759);
xnor U6170 (N_6170,N_4635,N_4885);
nor U6171 (N_6171,N_4631,N_4508);
and U6172 (N_6172,N_5551,N_4763);
or U6173 (N_6173,N_5366,N_4729);
and U6174 (N_6174,N_5968,N_5224);
and U6175 (N_6175,N_5222,N_5533);
nor U6176 (N_6176,N_5247,N_5900);
xor U6177 (N_6177,N_4624,N_4782);
nor U6178 (N_6178,N_5955,N_5830);
and U6179 (N_6179,N_5538,N_5461);
nor U6180 (N_6180,N_5600,N_5672);
nand U6181 (N_6181,N_5135,N_5387);
nand U6182 (N_6182,N_4518,N_5384);
or U6183 (N_6183,N_5321,N_5385);
xnor U6184 (N_6184,N_5643,N_4557);
xor U6185 (N_6185,N_4583,N_5511);
and U6186 (N_6186,N_5958,N_5557);
xor U6187 (N_6187,N_5616,N_5882);
and U6188 (N_6188,N_4725,N_4861);
xnor U6189 (N_6189,N_5084,N_5679);
nand U6190 (N_6190,N_4710,N_5009);
or U6191 (N_6191,N_5022,N_4968);
or U6192 (N_6192,N_4565,N_5531);
nor U6193 (N_6193,N_5410,N_5390);
nand U6194 (N_6194,N_5018,N_5058);
or U6195 (N_6195,N_5288,N_5652);
or U6196 (N_6196,N_5005,N_5117);
and U6197 (N_6197,N_5852,N_5554);
xnor U6198 (N_6198,N_4528,N_4632);
and U6199 (N_6199,N_5716,N_5253);
and U6200 (N_6200,N_5416,N_5930);
nand U6201 (N_6201,N_5639,N_5842);
xnor U6202 (N_6202,N_5822,N_4724);
nand U6203 (N_6203,N_5028,N_5078);
or U6204 (N_6204,N_5245,N_4614);
nand U6205 (N_6205,N_4720,N_4538);
nor U6206 (N_6206,N_5425,N_5298);
or U6207 (N_6207,N_5613,N_4598);
xor U6208 (N_6208,N_5198,N_4920);
nor U6209 (N_6209,N_5403,N_5848);
nand U6210 (N_6210,N_5481,N_5788);
or U6211 (N_6211,N_5274,N_5319);
xnor U6212 (N_6212,N_5764,N_5355);
nor U6213 (N_6213,N_5128,N_5484);
nor U6214 (N_6214,N_5063,N_5136);
xnor U6215 (N_6215,N_4826,N_5182);
xor U6216 (N_6216,N_5984,N_5174);
and U6217 (N_6217,N_5140,N_5473);
xnor U6218 (N_6218,N_5934,N_5100);
or U6219 (N_6219,N_5779,N_4980);
and U6220 (N_6220,N_5369,N_4525);
nor U6221 (N_6221,N_5053,N_5440);
or U6222 (N_6222,N_5443,N_5110);
xnor U6223 (N_6223,N_5468,N_5722);
nand U6224 (N_6224,N_4966,N_5422);
nand U6225 (N_6225,N_5164,N_5373);
or U6226 (N_6226,N_5421,N_5106);
nand U6227 (N_6227,N_5318,N_5526);
nand U6228 (N_6228,N_4543,N_5125);
and U6229 (N_6229,N_4740,N_5886);
or U6230 (N_6230,N_4884,N_5516);
or U6231 (N_6231,N_5055,N_4623);
nor U6232 (N_6232,N_4664,N_5296);
nor U6233 (N_6233,N_4852,N_4915);
and U6234 (N_6234,N_5124,N_4585);
nand U6235 (N_6235,N_5352,N_5378);
and U6236 (N_6236,N_5885,N_5910);
or U6237 (N_6237,N_4804,N_5609);
nand U6238 (N_6238,N_5260,N_5223);
xor U6239 (N_6239,N_5814,N_4672);
or U6240 (N_6240,N_5712,N_4503);
xnor U6241 (N_6241,N_5919,N_5663);
xnor U6242 (N_6242,N_4500,N_4817);
xnor U6243 (N_6243,N_4914,N_5865);
xnor U6244 (N_6244,N_5726,N_5052);
nand U6245 (N_6245,N_5008,N_5841);
or U6246 (N_6246,N_5301,N_4886);
or U6247 (N_6247,N_4865,N_5892);
or U6248 (N_6248,N_5233,N_5225);
and U6249 (N_6249,N_4997,N_4513);
nand U6250 (N_6250,N_5041,N_5747);
nor U6251 (N_6251,N_5112,N_5423);
nor U6252 (N_6252,N_4907,N_5918);
xnor U6253 (N_6253,N_5137,N_5420);
nand U6254 (N_6254,N_5938,N_5669);
nand U6255 (N_6255,N_5570,N_5913);
nand U6256 (N_6256,N_5278,N_5431);
nand U6257 (N_6257,N_5741,N_4605);
nor U6258 (N_6258,N_4847,N_4630);
or U6259 (N_6259,N_5297,N_4992);
nand U6260 (N_6260,N_4948,N_4533);
nand U6261 (N_6261,N_4612,N_5495);
and U6262 (N_6262,N_5665,N_4535);
and U6263 (N_6263,N_5191,N_4711);
nand U6264 (N_6264,N_5029,N_5291);
xnor U6265 (N_6265,N_4502,N_5987);
and U6266 (N_6266,N_4816,N_5525);
xor U6267 (N_6267,N_4922,N_5867);
and U6268 (N_6268,N_5147,N_4653);
or U6269 (N_6269,N_5784,N_5522);
nand U6270 (N_6270,N_4746,N_5002);
nor U6271 (N_6271,N_4990,N_4681);
nand U6272 (N_6272,N_4792,N_5792);
nor U6273 (N_6273,N_5889,N_4629);
nand U6274 (N_6274,N_4698,N_4935);
and U6275 (N_6275,N_4765,N_5528);
or U6276 (N_6276,N_5801,N_5118);
nand U6277 (N_6277,N_4716,N_5426);
nand U6278 (N_6278,N_5662,N_4696);
or U6279 (N_6279,N_5873,N_4993);
xor U6280 (N_6280,N_4743,N_4661);
nand U6281 (N_6281,N_4843,N_5047);
nor U6282 (N_6282,N_4796,N_5515);
nand U6283 (N_6283,N_5508,N_5577);
or U6284 (N_6284,N_5211,N_4633);
and U6285 (N_6285,N_5601,N_4846);
nand U6286 (N_6286,N_5532,N_4927);
nor U6287 (N_6287,N_5304,N_4582);
xor U6288 (N_6288,N_5899,N_5012);
nand U6289 (N_6289,N_4695,N_5901);
or U6290 (N_6290,N_5738,N_4555);
or U6291 (N_6291,N_4530,N_4923);
nor U6292 (N_6292,N_4504,N_5286);
nor U6293 (N_6293,N_5499,N_5381);
or U6294 (N_6294,N_4625,N_4893);
nor U6295 (N_6295,N_4692,N_5438);
nor U6296 (N_6296,N_4554,N_5678);
nor U6297 (N_6297,N_5610,N_5657);
nand U6298 (N_6298,N_5283,N_5793);
nand U6299 (N_6299,N_5720,N_5402);
nand U6300 (N_6300,N_5376,N_4872);
xnor U6301 (N_6301,N_4553,N_5187);
nor U6302 (N_6302,N_5486,N_5199);
xnor U6303 (N_6303,N_4560,N_5090);
nor U6304 (N_6304,N_5167,N_5107);
nor U6305 (N_6305,N_4580,N_4883);
or U6306 (N_6306,N_5152,N_4798);
nor U6307 (N_6307,N_5285,N_5762);
or U6308 (N_6308,N_4982,N_5581);
or U6309 (N_6309,N_5891,N_5116);
xor U6310 (N_6310,N_5345,N_4825);
nor U6311 (N_6311,N_5743,N_5588);
and U6312 (N_6312,N_5740,N_4570);
nor U6313 (N_6313,N_5433,N_4943);
nor U6314 (N_6314,N_4941,N_5275);
or U6315 (N_6315,N_5860,N_4949);
nand U6316 (N_6316,N_5184,N_5231);
or U6317 (N_6317,N_4862,N_5914);
or U6318 (N_6318,N_5095,N_5050);
xor U6319 (N_6319,N_4793,N_4738);
nor U6320 (N_6320,N_4974,N_5454);
or U6321 (N_6321,N_5768,N_4953);
nand U6322 (N_6322,N_5439,N_4878);
nand U6323 (N_6323,N_5099,N_5539);
nor U6324 (N_6324,N_4690,N_5640);
nand U6325 (N_6325,N_5178,N_5494);
or U6326 (N_6326,N_4753,N_5505);
or U6327 (N_6327,N_4925,N_5250);
nor U6328 (N_6328,N_5541,N_5417);
or U6329 (N_6329,N_5589,N_5790);
xor U6330 (N_6330,N_5572,N_4958);
and U6331 (N_6331,N_4754,N_4834);
nor U6332 (N_6332,N_4618,N_5469);
and U6333 (N_6333,N_4659,N_5655);
and U6334 (N_6334,N_5024,N_5911);
nand U6335 (N_6335,N_4741,N_5121);
nand U6336 (N_6336,N_4895,N_5510);
nor U6337 (N_6337,N_5386,N_4951);
nand U6338 (N_6338,N_4775,N_4913);
nand U6339 (N_6339,N_5309,N_5711);
or U6340 (N_6340,N_5875,N_5419);
nand U6341 (N_6341,N_5033,N_4545);
nor U6342 (N_6342,N_4760,N_4717);
and U6343 (N_6343,N_4609,N_4851);
xor U6344 (N_6344,N_4750,N_5686);
and U6345 (N_6345,N_5328,N_5483);
xnor U6346 (N_6346,N_4626,N_5745);
and U6347 (N_6347,N_5994,N_4832);
or U6348 (N_6348,N_5963,N_5687);
nor U6349 (N_6349,N_4873,N_4850);
xnor U6350 (N_6350,N_4827,N_4572);
or U6351 (N_6351,N_4813,N_4578);
xor U6352 (N_6352,N_5959,N_4811);
nand U6353 (N_6353,N_5565,N_4542);
or U6354 (N_6354,N_5183,N_5786);
and U6355 (N_6355,N_5664,N_5500);
xnor U6356 (N_6356,N_5341,N_4607);
xnor U6357 (N_6357,N_5081,N_4812);
nor U6358 (N_6358,N_4837,N_5559);
xnor U6359 (N_6359,N_4604,N_4870);
nor U6360 (N_6360,N_5243,N_5362);
and U6361 (N_6361,N_5698,N_4842);
nor U6362 (N_6362,N_4928,N_4603);
or U6363 (N_6363,N_4772,N_5070);
or U6364 (N_6364,N_5520,N_5252);
or U6365 (N_6365,N_5079,N_5017);
xnor U6366 (N_6366,N_4594,N_5394);
nand U6367 (N_6367,N_5413,N_5236);
nor U6368 (N_6368,N_4888,N_5583);
xnor U6369 (N_6369,N_4891,N_5329);
or U6370 (N_6370,N_5925,N_5003);
and U6371 (N_6371,N_4858,N_4790);
nand U6372 (N_6372,N_5217,N_4739);
xor U6373 (N_6373,N_4552,N_5068);
or U6374 (N_6374,N_4930,N_5982);
and U6375 (N_6375,N_5504,N_4961);
xnor U6376 (N_6376,N_5157,N_5103);
and U6377 (N_6377,N_5883,N_5509);
nor U6378 (N_6378,N_4652,N_4918);
nor U6379 (N_6379,N_4602,N_5569);
nor U6380 (N_6380,N_5696,N_5713);
and U6381 (N_6381,N_5308,N_4952);
nand U6382 (N_6382,N_4799,N_4749);
or U6383 (N_6383,N_5721,N_5656);
or U6384 (N_6384,N_5703,N_5874);
nand U6385 (N_6385,N_5205,N_4522);
or U6386 (N_6386,N_4877,N_5374);
xor U6387 (N_6387,N_5523,N_4821);
nor U6388 (N_6388,N_5389,N_5470);
or U6389 (N_6389,N_5324,N_5832);
xnor U6390 (N_6390,N_4579,N_5399);
xor U6391 (N_6391,N_5823,N_5746);
xnor U6392 (N_6392,N_5806,N_5825);
or U6393 (N_6393,N_5518,N_4981);
nand U6394 (N_6394,N_5621,N_5197);
or U6395 (N_6395,N_4591,N_5739);
and U6396 (N_6396,N_5618,N_4801);
xnor U6397 (N_6397,N_4685,N_5692);
xor U6398 (N_6398,N_5650,N_4726);
nand U6399 (N_6399,N_5161,N_5878);
xnor U6400 (N_6400,N_4809,N_4745);
and U6401 (N_6401,N_4869,N_5093);
nor U6402 (N_6402,N_4764,N_5400);
nand U6403 (N_6403,N_4556,N_4929);
nand U6404 (N_6404,N_4978,N_4894);
nor U6405 (N_6405,N_5496,N_5292);
nor U6406 (N_6406,N_5463,N_4934);
and U6407 (N_6407,N_4663,N_4785);
nor U6408 (N_6408,N_5733,N_5702);
xnor U6409 (N_6409,N_4802,N_4551);
and U6410 (N_6410,N_5820,N_5299);
xnor U6411 (N_6411,N_5584,N_5326);
and U6412 (N_6412,N_4828,N_5758);
or U6413 (N_6413,N_4947,N_4924);
xor U6414 (N_6414,N_5597,N_5344);
nor U6415 (N_6415,N_5844,N_4973);
or U6416 (N_6416,N_5917,N_5685);
nor U6417 (N_6417,N_5812,N_4700);
xor U6418 (N_6418,N_5320,N_4887);
xnor U6419 (N_6419,N_4524,N_4563);
xnor U6420 (N_6420,N_4712,N_5552);
xnor U6421 (N_6421,N_5947,N_5367);
and U6422 (N_6422,N_5916,N_4731);
and U6423 (N_6423,N_5109,N_5953);
nor U6424 (N_6424,N_5530,N_5069);
nand U6425 (N_6425,N_5353,N_4840);
and U6426 (N_6426,N_5980,N_5166);
nor U6427 (N_6427,N_5971,N_4620);
nand U6428 (N_6428,N_5266,N_5489);
or U6429 (N_6429,N_5165,N_5972);
or U6430 (N_6430,N_5859,N_4622);
or U6431 (N_6431,N_5194,N_5671);
nand U6432 (N_6432,N_4892,N_4536);
xor U6433 (N_6433,N_5330,N_4776);
nand U6434 (N_6434,N_4516,N_5040);
and U6435 (N_6435,N_4962,N_4788);
or U6436 (N_6436,N_5268,N_5193);
nor U6437 (N_6437,N_5619,N_5126);
and U6438 (N_6438,N_5368,N_5241);
nand U6439 (N_6439,N_5087,N_4691);
nor U6440 (N_6440,N_5923,N_5781);
and U6441 (N_6441,N_5295,N_5113);
and U6442 (N_6442,N_5388,N_5088);
nor U6443 (N_6443,N_5596,N_4921);
or U6444 (N_6444,N_4786,N_5877);
nor U6445 (N_6445,N_5190,N_5944);
and U6446 (N_6446,N_5699,N_4989);
or U6447 (N_6447,N_5744,N_4778);
nand U6448 (N_6448,N_4882,N_5460);
or U6449 (N_6449,N_5695,N_5016);
nand U6450 (N_6450,N_5120,N_4517);
nor U6451 (N_6451,N_5939,N_5615);
or U6452 (N_6452,N_5673,N_4676);
nand U6453 (N_6453,N_4815,N_4660);
nand U6454 (N_6454,N_5846,N_5313);
nand U6455 (N_6455,N_5787,N_5228);
or U6456 (N_6456,N_5946,N_5789);
xnor U6457 (N_6457,N_5717,N_5681);
nand U6458 (N_6458,N_4919,N_5256);
nor U6459 (N_6459,N_5139,N_5054);
or U6460 (N_6460,N_5115,N_4937);
and U6461 (N_6461,N_4529,N_4905);
xor U6462 (N_6462,N_5626,N_4908);
or U6463 (N_6463,N_5466,N_5819);
or U6464 (N_6464,N_4787,N_4864);
nor U6465 (N_6465,N_5607,N_5907);
nand U6466 (N_6466,N_5325,N_4655);
xor U6467 (N_6467,N_5092,N_4644);
nand U6468 (N_6468,N_5432,N_4768);
or U6469 (N_6469,N_4587,N_5872);
nor U6470 (N_6470,N_4939,N_4656);
nor U6471 (N_6471,N_5273,N_5021);
xor U6472 (N_6472,N_4900,N_5122);
xor U6473 (N_6473,N_5281,N_5964);
nor U6474 (N_6474,N_5641,N_5246);
xnor U6475 (N_6475,N_5700,N_4613);
nand U6476 (N_6476,N_5582,N_5849);
or U6477 (N_6477,N_5065,N_5074);
nor U6478 (N_6478,N_4569,N_5143);
and U6479 (N_6479,N_5833,N_5282);
nand U6480 (N_6480,N_5044,N_5181);
and U6481 (N_6481,N_4640,N_4983);
nor U6482 (N_6482,N_5732,N_5851);
or U6483 (N_6483,N_5694,N_5602);
or U6484 (N_6484,N_5676,N_5608);
nand U6485 (N_6485,N_5444,N_5777);
nand U6486 (N_6486,N_4898,N_5392);
or U6487 (N_6487,N_5977,N_4863);
or U6488 (N_6488,N_4880,N_5263);
and U6489 (N_6489,N_5415,N_5363);
and U6490 (N_6490,N_5441,N_5497);
and U6491 (N_6491,N_4636,N_4762);
or U6492 (N_6492,N_4584,N_5561);
or U6493 (N_6493,N_5358,N_5864);
nor U6494 (N_6494,N_4705,N_5753);
or U6495 (N_6495,N_5323,N_5729);
or U6496 (N_6496,N_4848,N_5897);
or U6497 (N_6497,N_4779,N_5405);
xnor U6498 (N_6498,N_5334,N_5035);
or U6499 (N_6499,N_5467,N_4932);
nor U6500 (N_6500,N_5529,N_5270);
xnor U6501 (N_6501,N_5750,N_4561);
xor U6502 (N_6502,N_5427,N_4693);
nor U6503 (N_6503,N_5862,N_5991);
nand U6504 (N_6504,N_4568,N_5780);
and U6505 (N_6505,N_5791,N_4896);
and U6506 (N_6506,N_5579,N_5881);
and U6507 (N_6507,N_5265,N_5776);
and U6508 (N_6508,N_5042,N_5173);
nor U6509 (N_6509,N_4794,N_4860);
or U6510 (N_6510,N_5800,N_4658);
nand U6511 (N_6511,N_5547,N_5331);
xor U6512 (N_6512,N_5097,N_5089);
or U6513 (N_6513,N_5271,N_4969);
or U6514 (N_6514,N_5818,N_5926);
xnor U6515 (N_6515,N_5869,N_4857);
nor U6516 (N_6516,N_4967,N_5195);
and U6517 (N_6517,N_5513,N_5377);
or U6518 (N_6518,N_5051,N_5783);
and U6519 (N_6519,N_5354,N_5429);
or U6520 (N_6520,N_5310,N_5216);
and U6521 (N_6521,N_4755,N_4610);
xnor U6522 (N_6522,N_5339,N_4866);
or U6523 (N_6523,N_5083,N_5642);
and U6524 (N_6524,N_4534,N_5407);
or U6525 (N_6525,N_4549,N_5447);
xnor U6526 (N_6526,N_5206,N_5064);
nor U6527 (N_6527,N_4964,N_5340);
xor U6528 (N_6528,N_5940,N_5472);
nor U6529 (N_6529,N_4770,N_5085);
nor U6530 (N_6530,N_5019,N_5056);
or U6531 (N_6531,N_5838,N_5811);
xnor U6532 (N_6532,N_5475,N_5150);
and U6533 (N_6533,N_5863,N_4703);
nor U6534 (N_6534,N_4654,N_5759);
nor U6535 (N_6535,N_5160,N_5683);
nand U6536 (N_6536,N_4831,N_5480);
and U6537 (N_6537,N_5749,N_4718);
nor U6538 (N_6538,N_4940,N_5904);
nand U6539 (N_6539,N_5091,N_4548);
nand U6540 (N_6540,N_5242,N_5587);
nand U6541 (N_6541,N_5813,N_5011);
or U6542 (N_6542,N_5492,N_4606);
xnor U6543 (N_6543,N_4950,N_4541);
nand U6544 (N_6544,N_5108,N_4757);
nor U6545 (N_6545,N_4835,N_4694);
and U6546 (N_6546,N_5186,N_5478);
and U6547 (N_6547,N_5568,N_5346);
nand U6548 (N_6548,N_5879,N_5501);
xnor U6549 (N_6549,N_5360,N_4742);
and U6550 (N_6550,N_5769,N_5189);
nand U6551 (N_6551,N_5163,N_5096);
and U6552 (N_6552,N_5212,N_5203);
and U6553 (N_6553,N_4944,N_5031);
nor U6554 (N_6554,N_5261,N_5603);
xor U6555 (N_6555,N_4747,N_5564);
nor U6556 (N_6556,N_5843,N_4803);
xnor U6557 (N_6557,N_5563,N_5622);
and U6558 (N_6558,N_5082,N_5634);
nor U6559 (N_6559,N_4985,N_5076);
nand U6560 (N_6560,N_4797,N_4627);
and U6561 (N_6561,N_4931,N_5327);
nor U6562 (N_6562,N_5893,N_4976);
and U6563 (N_6563,N_5908,N_5701);
xor U6564 (N_6564,N_5146,N_5766);
and U6565 (N_6565,N_5312,N_5857);
nand U6566 (N_6566,N_4822,N_5578);
nor U6567 (N_6567,N_5383,N_5158);
xnor U6568 (N_6568,N_4996,N_5479);
and U6569 (N_6569,N_5086,N_4806);
nand U6570 (N_6570,N_4819,N_4916);
nand U6571 (N_6571,N_4595,N_4566);
nand U6572 (N_6572,N_4667,N_5948);
or U6573 (N_6573,N_5172,N_5006);
nand U6574 (N_6574,N_4902,N_5675);
or U6575 (N_6575,N_5398,N_4689);
xnor U6576 (N_6576,N_5751,N_4645);
nand U6577 (N_6577,N_4737,N_4687);
nand U6578 (N_6578,N_5651,N_5317);
or U6579 (N_6579,N_4509,N_4575);
or U6580 (N_6580,N_4986,N_4638);
xor U6581 (N_6581,N_5537,N_5406);
xnor U6582 (N_6582,N_5148,N_5046);
nand U6583 (N_6583,N_4599,N_5032);
and U6584 (N_6584,N_5826,N_5725);
or U6585 (N_6585,N_4531,N_4805);
or U6586 (N_6586,N_4844,N_5954);
nand U6587 (N_6587,N_5845,N_5706);
nand U6588 (N_6588,N_5001,N_5498);
nand U6589 (N_6589,N_5730,N_5970);
and U6590 (N_6590,N_4881,N_5371);
and U6591 (N_6591,N_5804,N_4673);
and U6592 (N_6592,N_5338,N_5465);
nor U6593 (N_6593,N_5075,N_5234);
or U6594 (N_6594,N_5997,N_5506);
xnor U6595 (N_6595,N_4988,N_5337);
xor U6596 (N_6596,N_5527,N_5322);
or U6597 (N_6597,N_5034,N_5142);
nand U6598 (N_6598,N_4671,N_5576);
xnor U6599 (N_6599,N_4959,N_5737);
nand U6600 (N_6600,N_5562,N_5556);
or U6601 (N_6601,N_5855,N_5094);
or U6602 (N_6602,N_5536,N_4849);
nor U6603 (N_6603,N_5382,N_4987);
nand U6604 (N_6604,N_5519,N_5204);
nor U6605 (N_6605,N_5770,N_4933);
or U6606 (N_6606,N_4756,N_5350);
nor U6607 (N_6607,N_4730,N_5714);
nand U6608 (N_6608,N_4965,N_4774);
nor U6609 (N_6609,N_5004,N_4971);
xor U6610 (N_6610,N_5896,N_4702);
xnor U6611 (N_6611,N_5798,N_5920);
xnor U6612 (N_6612,N_4657,N_5077);
or U6613 (N_6613,N_5649,N_4855);
or U6614 (N_6614,N_5257,N_5149);
or U6615 (N_6615,N_4699,N_4979);
nand U6616 (N_6616,N_5141,N_5502);
nand U6617 (N_6617,N_5279,N_5209);
or U6618 (N_6618,N_5332,N_5566);
and U6619 (N_6619,N_5159,N_4906);
or U6620 (N_6620,N_5025,N_5927);
or U6621 (N_6621,N_4520,N_5446);
xnor U6622 (N_6622,N_5131,N_4505);
or U6623 (N_6623,N_5020,N_4999);
nor U6624 (N_6624,N_5594,N_5633);
xnor U6625 (N_6625,N_4611,N_5637);
nand U6626 (N_6626,N_5710,N_5059);
nor U6627 (N_6627,N_4722,N_5177);
nand U6628 (N_6628,N_5870,N_5045);
nor U6629 (N_6629,N_5464,N_4532);
and U6630 (N_6630,N_5503,N_5571);
nor U6631 (N_6631,N_5962,N_5305);
xor U6632 (N_6632,N_5039,N_5995);
nand U6633 (N_6633,N_5763,N_5391);
or U6634 (N_6634,N_5831,N_5861);
and U6635 (N_6635,N_5180,N_5015);
nand U6636 (N_6636,N_5957,N_5347);
or U6637 (N_6637,N_5248,N_5488);
or U6638 (N_6638,N_4589,N_5829);
or U6639 (N_6639,N_4955,N_5311);
nand U6640 (N_6640,N_5208,N_5548);
and U6641 (N_6641,N_4977,N_4577);
xor U6642 (N_6642,N_5903,N_5612);
xnor U6643 (N_6643,N_4769,N_5335);
xor U6644 (N_6644,N_5580,N_5284);
xor U6645 (N_6645,N_5575,N_4515);
nand U6646 (N_6646,N_5951,N_4868);
and U6647 (N_6647,N_4706,N_4506);
or U6648 (N_6648,N_5514,N_5989);
or U6649 (N_6649,N_5742,N_5709);
nand U6650 (N_6650,N_4564,N_5129);
nand U6651 (N_6651,N_4574,N_4910);
xor U6652 (N_6652,N_5757,N_5458);
and U6653 (N_6653,N_5595,N_5765);
xnor U6654 (N_6654,N_5827,N_4547);
nor U6655 (N_6655,N_5477,N_5558);
and U6656 (N_6656,N_5898,N_5707);
and U6657 (N_6657,N_4839,N_4946);
xnor U6658 (N_6658,N_4936,N_5485);
or U6659 (N_6659,N_4771,N_5629);
xnor U6660 (N_6660,N_5026,N_5457);
and U6661 (N_6661,N_5821,N_5993);
nor U6662 (N_6662,N_4521,N_5277);
and U6663 (N_6663,N_5606,N_4853);
xor U6664 (N_6664,N_5448,N_5306);
xnor U6665 (N_6665,N_5684,N_4619);
nand U6666 (N_6666,N_5986,N_5280);
nand U6667 (N_6667,N_5961,N_5599);
and U6668 (N_6668,N_5418,N_5540);
nor U6669 (N_6669,N_5119,N_5719);
xnor U6670 (N_6670,N_4748,N_5623);
xnor U6671 (N_6671,N_4732,N_5614);
and U6672 (N_6672,N_5459,N_4608);
and U6673 (N_6673,N_4615,N_4519);
nor U6674 (N_6674,N_5272,N_5315);
and U6675 (N_6675,N_5534,N_5185);
or U6676 (N_6676,N_5151,N_4841);
or U6677 (N_6677,N_4836,N_5359);
nand U6678 (N_6678,N_5544,N_5162);
or U6679 (N_6679,N_5816,N_5192);
nor U6680 (N_6680,N_4540,N_5154);
nor U6681 (N_6681,N_4546,N_5249);
and U6682 (N_6682,N_4723,N_4637);
nand U6683 (N_6683,N_5287,N_5667);
nand U6684 (N_6684,N_5210,N_5101);
and U6685 (N_6685,N_4537,N_5393);
nor U6686 (N_6686,N_5239,N_4856);
and U6687 (N_6687,N_4510,N_5437);
and U6688 (N_6688,N_5981,N_5658);
and U6689 (N_6689,N_5931,N_5724);
nand U6690 (N_6690,N_4708,N_5220);
xor U6691 (N_6691,N_5007,N_5876);
nor U6692 (N_6692,N_5727,N_5976);
nand U6693 (N_6693,N_4789,N_5232);
and U6694 (N_6694,N_4719,N_5705);
and U6695 (N_6695,N_5155,N_5351);
and U6696 (N_6696,N_5356,N_5975);
nand U6697 (N_6697,N_5179,N_4523);
nor U6698 (N_6698,N_4544,N_4634);
or U6699 (N_6699,N_5736,N_5293);
and U6700 (N_6700,N_4688,N_5894);
nand U6701 (N_6701,N_5023,N_5545);
nand U6702 (N_6702,N_4596,N_4820);
nand U6703 (N_6703,N_5175,N_5455);
nand U6704 (N_6704,N_5490,N_4752);
nor U6705 (N_6705,N_5424,N_5343);
xor U6706 (N_6706,N_5847,N_4874);
and U6707 (N_6707,N_5255,N_4567);
or U6708 (N_6708,N_4912,N_4514);
or U6709 (N_6709,N_5030,N_4889);
nor U6710 (N_6710,N_4597,N_5691);
nor U6711 (N_6711,N_5593,N_5364);
or U6712 (N_6712,N_4945,N_5227);
nand U6713 (N_6713,N_5590,N_4995);
xor U6714 (N_6714,N_4791,N_5229);
nor U6715 (N_6715,N_5928,N_4744);
nor U6716 (N_6716,N_5202,N_5932);
nor U6717 (N_6717,N_5302,N_5207);
xor U6718 (N_6718,N_5104,N_5471);
nor U6719 (N_6719,N_5949,N_5244);
nand U6720 (N_6720,N_5542,N_5235);
and U6721 (N_6721,N_5014,N_5171);
nor U6722 (N_6722,N_5817,N_5620);
xnor U6723 (N_6723,N_5906,N_4859);
or U6724 (N_6724,N_5474,N_5799);
or U6725 (N_6725,N_5048,N_5912);
and U6726 (N_6726,N_4904,N_5156);
and U6727 (N_6727,N_4600,N_5660);
xnor U6728 (N_6728,N_4662,N_5170);
and U6729 (N_6729,N_5988,N_5868);
nand U6730 (N_6730,N_5434,N_5546);
nand U6731 (N_6731,N_5632,N_5036);
or U6732 (N_6732,N_5259,N_5491);
or U6733 (N_6733,N_5409,N_5176);
or U6734 (N_6734,N_5624,N_5752);
nor U6735 (N_6735,N_5653,N_4592);
and U6736 (N_6736,N_5965,N_4808);
xor U6737 (N_6737,N_5251,N_4649);
nand U6738 (N_6738,N_4697,N_5585);
and U6739 (N_6739,N_5555,N_5952);
or U6740 (N_6740,N_4942,N_4590);
xor U6741 (N_6741,N_5775,N_5375);
or U6742 (N_6742,N_5854,N_5836);
nand U6743 (N_6743,N_4734,N_5996);
nand U6744 (N_6744,N_5771,N_5482);
and U6745 (N_6745,N_5592,N_4665);
xor U6746 (N_6746,N_4674,N_5909);
xnor U6747 (N_6747,N_4879,N_5560);
nand U6748 (N_6748,N_4970,N_4845);
xnor U6749 (N_6749,N_5837,N_5888);
nor U6750 (N_6750,N_5616,N_5640);
and U6751 (N_6751,N_4742,N_5364);
nor U6752 (N_6752,N_4520,N_4870);
nand U6753 (N_6753,N_5700,N_5561);
nor U6754 (N_6754,N_5540,N_5690);
nand U6755 (N_6755,N_5877,N_4828);
xor U6756 (N_6756,N_5958,N_5797);
and U6757 (N_6757,N_5017,N_5434);
or U6758 (N_6758,N_5972,N_5910);
and U6759 (N_6759,N_5590,N_5195);
xnor U6760 (N_6760,N_4634,N_4664);
nand U6761 (N_6761,N_4715,N_4588);
nand U6762 (N_6762,N_4630,N_5088);
and U6763 (N_6763,N_4731,N_4883);
xor U6764 (N_6764,N_4663,N_5599);
nand U6765 (N_6765,N_5622,N_5030);
or U6766 (N_6766,N_5917,N_4738);
nor U6767 (N_6767,N_5813,N_4856);
nand U6768 (N_6768,N_5241,N_5377);
and U6769 (N_6769,N_5360,N_4947);
xnor U6770 (N_6770,N_4692,N_4832);
nand U6771 (N_6771,N_4530,N_5486);
or U6772 (N_6772,N_4890,N_4506);
and U6773 (N_6773,N_5937,N_5809);
and U6774 (N_6774,N_5378,N_4685);
or U6775 (N_6775,N_5319,N_5206);
nor U6776 (N_6776,N_5403,N_4849);
or U6777 (N_6777,N_4805,N_4774);
xor U6778 (N_6778,N_5433,N_5286);
and U6779 (N_6779,N_5720,N_5198);
or U6780 (N_6780,N_5130,N_5700);
nor U6781 (N_6781,N_5701,N_4604);
xnor U6782 (N_6782,N_5475,N_5409);
nand U6783 (N_6783,N_5938,N_4589);
nand U6784 (N_6784,N_5192,N_5284);
and U6785 (N_6785,N_5895,N_5767);
nor U6786 (N_6786,N_4704,N_5421);
nand U6787 (N_6787,N_4999,N_4577);
xor U6788 (N_6788,N_5639,N_5701);
xnor U6789 (N_6789,N_4614,N_4758);
or U6790 (N_6790,N_4797,N_5041);
nor U6791 (N_6791,N_4925,N_4642);
and U6792 (N_6792,N_4764,N_5180);
nor U6793 (N_6793,N_5245,N_5885);
or U6794 (N_6794,N_5829,N_5925);
and U6795 (N_6795,N_4825,N_5180);
nand U6796 (N_6796,N_4562,N_5772);
xor U6797 (N_6797,N_5500,N_4580);
xnor U6798 (N_6798,N_4518,N_5012);
xnor U6799 (N_6799,N_4885,N_4628);
or U6800 (N_6800,N_5671,N_4932);
xor U6801 (N_6801,N_4938,N_5380);
nor U6802 (N_6802,N_5256,N_4806);
and U6803 (N_6803,N_5968,N_4541);
nor U6804 (N_6804,N_5226,N_4884);
nand U6805 (N_6805,N_5594,N_5580);
nor U6806 (N_6806,N_5437,N_5273);
xor U6807 (N_6807,N_5530,N_5522);
xnor U6808 (N_6808,N_5410,N_4789);
nand U6809 (N_6809,N_5653,N_5982);
xnor U6810 (N_6810,N_5021,N_4729);
and U6811 (N_6811,N_4597,N_5019);
nand U6812 (N_6812,N_5288,N_5947);
nand U6813 (N_6813,N_4956,N_5174);
nor U6814 (N_6814,N_5120,N_5056);
nor U6815 (N_6815,N_5813,N_5298);
nand U6816 (N_6816,N_4666,N_5869);
xor U6817 (N_6817,N_4786,N_5100);
nand U6818 (N_6818,N_5117,N_5414);
xnor U6819 (N_6819,N_5869,N_5971);
xnor U6820 (N_6820,N_4626,N_4953);
or U6821 (N_6821,N_4848,N_5501);
and U6822 (N_6822,N_5183,N_5923);
and U6823 (N_6823,N_5450,N_5348);
or U6824 (N_6824,N_4566,N_5711);
or U6825 (N_6825,N_5194,N_4633);
xnor U6826 (N_6826,N_5544,N_4955);
nand U6827 (N_6827,N_4647,N_4681);
nand U6828 (N_6828,N_5952,N_5229);
and U6829 (N_6829,N_5399,N_4613);
or U6830 (N_6830,N_4642,N_5742);
xor U6831 (N_6831,N_4560,N_5845);
or U6832 (N_6832,N_5547,N_4541);
nor U6833 (N_6833,N_4795,N_5576);
and U6834 (N_6834,N_4868,N_5539);
and U6835 (N_6835,N_5539,N_4986);
xor U6836 (N_6836,N_5188,N_5618);
or U6837 (N_6837,N_5704,N_4967);
nor U6838 (N_6838,N_4612,N_5325);
nand U6839 (N_6839,N_5926,N_5551);
and U6840 (N_6840,N_4669,N_4836);
or U6841 (N_6841,N_5291,N_5255);
nand U6842 (N_6842,N_5117,N_5041);
and U6843 (N_6843,N_4992,N_4839);
or U6844 (N_6844,N_5570,N_5132);
xnor U6845 (N_6845,N_4726,N_4577);
nor U6846 (N_6846,N_5593,N_5500);
and U6847 (N_6847,N_5412,N_5438);
nand U6848 (N_6848,N_5289,N_5926);
nand U6849 (N_6849,N_5340,N_4722);
xnor U6850 (N_6850,N_5554,N_5911);
or U6851 (N_6851,N_5708,N_4674);
nor U6852 (N_6852,N_5146,N_4786);
nor U6853 (N_6853,N_5037,N_5501);
nor U6854 (N_6854,N_5333,N_5764);
nor U6855 (N_6855,N_4734,N_5845);
nand U6856 (N_6856,N_5364,N_5949);
or U6857 (N_6857,N_5160,N_4527);
or U6858 (N_6858,N_5083,N_5561);
or U6859 (N_6859,N_5431,N_5847);
or U6860 (N_6860,N_5372,N_4866);
or U6861 (N_6861,N_5146,N_5412);
nor U6862 (N_6862,N_4511,N_5503);
nand U6863 (N_6863,N_5843,N_5677);
nor U6864 (N_6864,N_5737,N_4842);
and U6865 (N_6865,N_4630,N_5543);
or U6866 (N_6866,N_4890,N_5623);
xnor U6867 (N_6867,N_4822,N_4954);
xnor U6868 (N_6868,N_5022,N_5903);
xor U6869 (N_6869,N_5976,N_4501);
and U6870 (N_6870,N_5656,N_5254);
nor U6871 (N_6871,N_5609,N_4714);
or U6872 (N_6872,N_5226,N_4608);
nand U6873 (N_6873,N_4916,N_5070);
and U6874 (N_6874,N_4705,N_5849);
nor U6875 (N_6875,N_5938,N_5721);
xnor U6876 (N_6876,N_4830,N_5669);
or U6877 (N_6877,N_5593,N_5759);
xor U6878 (N_6878,N_5775,N_4677);
or U6879 (N_6879,N_4637,N_4771);
and U6880 (N_6880,N_5756,N_5180);
and U6881 (N_6881,N_5971,N_5528);
or U6882 (N_6882,N_4670,N_4825);
or U6883 (N_6883,N_5962,N_4976);
or U6884 (N_6884,N_4743,N_5711);
or U6885 (N_6885,N_5428,N_4897);
or U6886 (N_6886,N_5213,N_4616);
nor U6887 (N_6887,N_5294,N_4662);
and U6888 (N_6888,N_4787,N_5414);
nand U6889 (N_6889,N_5005,N_5833);
or U6890 (N_6890,N_5547,N_5091);
and U6891 (N_6891,N_5357,N_5154);
nor U6892 (N_6892,N_4773,N_5363);
or U6893 (N_6893,N_4947,N_5902);
nor U6894 (N_6894,N_5230,N_4989);
and U6895 (N_6895,N_5592,N_5497);
nand U6896 (N_6896,N_4562,N_5790);
or U6897 (N_6897,N_5581,N_5077);
or U6898 (N_6898,N_5880,N_5878);
nor U6899 (N_6899,N_5491,N_5983);
nor U6900 (N_6900,N_5264,N_4935);
nand U6901 (N_6901,N_5501,N_5042);
or U6902 (N_6902,N_4528,N_5109);
xnor U6903 (N_6903,N_5068,N_5441);
or U6904 (N_6904,N_5860,N_5278);
and U6905 (N_6905,N_5926,N_5782);
nand U6906 (N_6906,N_5833,N_5665);
or U6907 (N_6907,N_5870,N_5604);
xnor U6908 (N_6908,N_5602,N_5981);
nand U6909 (N_6909,N_5990,N_5384);
nand U6910 (N_6910,N_4746,N_4743);
or U6911 (N_6911,N_5863,N_5039);
or U6912 (N_6912,N_5796,N_5018);
or U6913 (N_6913,N_5074,N_4612);
xnor U6914 (N_6914,N_5202,N_4881);
nor U6915 (N_6915,N_5009,N_5096);
nand U6916 (N_6916,N_5974,N_5813);
nor U6917 (N_6917,N_5405,N_5533);
or U6918 (N_6918,N_5292,N_4737);
or U6919 (N_6919,N_5644,N_5902);
xnor U6920 (N_6920,N_5465,N_5920);
nor U6921 (N_6921,N_4867,N_5083);
nor U6922 (N_6922,N_5699,N_4860);
or U6923 (N_6923,N_5488,N_5859);
xor U6924 (N_6924,N_4854,N_4641);
or U6925 (N_6925,N_4594,N_5360);
nor U6926 (N_6926,N_4942,N_5534);
xor U6927 (N_6927,N_4857,N_5824);
nor U6928 (N_6928,N_5223,N_5203);
xnor U6929 (N_6929,N_5303,N_5563);
or U6930 (N_6930,N_5034,N_5777);
or U6931 (N_6931,N_5823,N_5702);
nand U6932 (N_6932,N_5382,N_5846);
nor U6933 (N_6933,N_4875,N_5520);
xnor U6934 (N_6934,N_5693,N_4613);
nand U6935 (N_6935,N_5088,N_4976);
xor U6936 (N_6936,N_4563,N_4560);
nor U6937 (N_6937,N_4978,N_5794);
nor U6938 (N_6938,N_5462,N_5011);
and U6939 (N_6939,N_4862,N_5578);
nand U6940 (N_6940,N_5686,N_5353);
or U6941 (N_6941,N_5643,N_5257);
nor U6942 (N_6942,N_5219,N_5020);
nand U6943 (N_6943,N_5628,N_4692);
xor U6944 (N_6944,N_5963,N_5514);
or U6945 (N_6945,N_4608,N_5379);
or U6946 (N_6946,N_5050,N_5101);
xnor U6947 (N_6947,N_5607,N_5887);
xor U6948 (N_6948,N_5298,N_5337);
or U6949 (N_6949,N_5065,N_5036);
nor U6950 (N_6950,N_5153,N_5359);
xor U6951 (N_6951,N_5119,N_4826);
or U6952 (N_6952,N_5290,N_4640);
nor U6953 (N_6953,N_5914,N_5825);
nand U6954 (N_6954,N_5315,N_4589);
xnor U6955 (N_6955,N_5421,N_5203);
xor U6956 (N_6956,N_5753,N_4632);
nor U6957 (N_6957,N_5082,N_5425);
or U6958 (N_6958,N_5698,N_5396);
nor U6959 (N_6959,N_4935,N_5790);
xnor U6960 (N_6960,N_5573,N_5323);
or U6961 (N_6961,N_5326,N_5771);
or U6962 (N_6962,N_5634,N_4598);
xor U6963 (N_6963,N_4537,N_5519);
or U6964 (N_6964,N_4784,N_5526);
or U6965 (N_6965,N_5747,N_5161);
xnor U6966 (N_6966,N_5762,N_4951);
or U6967 (N_6967,N_4522,N_4792);
or U6968 (N_6968,N_4809,N_4688);
xor U6969 (N_6969,N_5764,N_5776);
and U6970 (N_6970,N_5165,N_5085);
nand U6971 (N_6971,N_5546,N_5416);
nor U6972 (N_6972,N_5954,N_5986);
nand U6973 (N_6973,N_4990,N_5140);
xor U6974 (N_6974,N_5041,N_5250);
nor U6975 (N_6975,N_4734,N_5085);
xor U6976 (N_6976,N_5300,N_4682);
and U6977 (N_6977,N_4839,N_5686);
nor U6978 (N_6978,N_4643,N_5108);
or U6979 (N_6979,N_5777,N_4565);
or U6980 (N_6980,N_5106,N_4822);
xnor U6981 (N_6981,N_5493,N_5036);
nand U6982 (N_6982,N_5567,N_5104);
or U6983 (N_6983,N_4787,N_4823);
and U6984 (N_6984,N_4554,N_5876);
xnor U6985 (N_6985,N_5528,N_4564);
nand U6986 (N_6986,N_5734,N_5809);
or U6987 (N_6987,N_4515,N_4880);
and U6988 (N_6988,N_5260,N_4688);
xor U6989 (N_6989,N_5743,N_5908);
or U6990 (N_6990,N_4558,N_4744);
xnor U6991 (N_6991,N_5775,N_4509);
xnor U6992 (N_6992,N_4822,N_5593);
xnor U6993 (N_6993,N_5701,N_4737);
and U6994 (N_6994,N_5670,N_4778);
xor U6995 (N_6995,N_5014,N_4665);
or U6996 (N_6996,N_5190,N_4788);
or U6997 (N_6997,N_5511,N_5413);
nor U6998 (N_6998,N_5985,N_5169);
and U6999 (N_6999,N_4680,N_4781);
nor U7000 (N_7000,N_4934,N_5044);
xor U7001 (N_7001,N_5839,N_4864);
and U7002 (N_7002,N_5797,N_5306);
or U7003 (N_7003,N_4905,N_4808);
nor U7004 (N_7004,N_4666,N_5078);
nor U7005 (N_7005,N_5446,N_5028);
nor U7006 (N_7006,N_5230,N_5709);
nand U7007 (N_7007,N_5604,N_4900);
nand U7008 (N_7008,N_5959,N_5000);
and U7009 (N_7009,N_5238,N_4720);
and U7010 (N_7010,N_5726,N_5707);
xnor U7011 (N_7011,N_4969,N_5428);
and U7012 (N_7012,N_5437,N_5484);
nor U7013 (N_7013,N_5889,N_4506);
xor U7014 (N_7014,N_4798,N_5707);
or U7015 (N_7015,N_5827,N_5581);
xor U7016 (N_7016,N_4934,N_5617);
nor U7017 (N_7017,N_5568,N_5213);
and U7018 (N_7018,N_4527,N_4869);
or U7019 (N_7019,N_5487,N_4747);
or U7020 (N_7020,N_5651,N_5974);
nor U7021 (N_7021,N_4846,N_5518);
nor U7022 (N_7022,N_5456,N_5606);
nand U7023 (N_7023,N_5780,N_5169);
nor U7024 (N_7024,N_5744,N_4528);
nor U7025 (N_7025,N_5262,N_5301);
and U7026 (N_7026,N_5796,N_4777);
nor U7027 (N_7027,N_5389,N_5472);
and U7028 (N_7028,N_4856,N_5405);
or U7029 (N_7029,N_5751,N_5414);
nor U7030 (N_7030,N_5423,N_4625);
nand U7031 (N_7031,N_4669,N_5576);
nand U7032 (N_7032,N_5460,N_4749);
and U7033 (N_7033,N_5554,N_5613);
or U7034 (N_7034,N_5745,N_5903);
xnor U7035 (N_7035,N_5481,N_5770);
xor U7036 (N_7036,N_4897,N_5736);
nand U7037 (N_7037,N_4833,N_4920);
nand U7038 (N_7038,N_5872,N_4705);
or U7039 (N_7039,N_5046,N_4617);
and U7040 (N_7040,N_4807,N_5394);
nand U7041 (N_7041,N_4656,N_5215);
nand U7042 (N_7042,N_5970,N_4693);
xnor U7043 (N_7043,N_5762,N_5698);
and U7044 (N_7044,N_4578,N_4545);
nor U7045 (N_7045,N_5711,N_4568);
or U7046 (N_7046,N_5870,N_5838);
nor U7047 (N_7047,N_5722,N_4509);
or U7048 (N_7048,N_4770,N_5124);
nand U7049 (N_7049,N_5492,N_4770);
or U7050 (N_7050,N_4801,N_5059);
or U7051 (N_7051,N_5216,N_4600);
nor U7052 (N_7052,N_5086,N_4723);
or U7053 (N_7053,N_4906,N_5531);
nand U7054 (N_7054,N_4805,N_5587);
xor U7055 (N_7055,N_5290,N_5704);
nor U7056 (N_7056,N_4700,N_4907);
or U7057 (N_7057,N_5791,N_5612);
nand U7058 (N_7058,N_4986,N_5490);
and U7059 (N_7059,N_5105,N_4622);
nand U7060 (N_7060,N_5528,N_4585);
nand U7061 (N_7061,N_4814,N_5992);
nand U7062 (N_7062,N_5529,N_5048);
or U7063 (N_7063,N_5482,N_5661);
or U7064 (N_7064,N_4824,N_4938);
and U7065 (N_7065,N_4873,N_4916);
and U7066 (N_7066,N_5616,N_5199);
nand U7067 (N_7067,N_5045,N_5711);
or U7068 (N_7068,N_5555,N_5766);
nor U7069 (N_7069,N_5239,N_5600);
and U7070 (N_7070,N_4957,N_5810);
nand U7071 (N_7071,N_4712,N_5193);
and U7072 (N_7072,N_5606,N_5394);
nor U7073 (N_7073,N_5252,N_5949);
or U7074 (N_7074,N_4943,N_5543);
and U7075 (N_7075,N_5791,N_5831);
nand U7076 (N_7076,N_5654,N_5474);
xnor U7077 (N_7077,N_5700,N_4720);
nor U7078 (N_7078,N_5959,N_5954);
or U7079 (N_7079,N_4947,N_5383);
xnor U7080 (N_7080,N_4606,N_4641);
nor U7081 (N_7081,N_5696,N_5100);
or U7082 (N_7082,N_5229,N_5839);
xnor U7083 (N_7083,N_4919,N_4967);
nand U7084 (N_7084,N_5284,N_5208);
nor U7085 (N_7085,N_5401,N_5169);
nor U7086 (N_7086,N_5959,N_5234);
nor U7087 (N_7087,N_5866,N_4684);
nor U7088 (N_7088,N_4821,N_5267);
nand U7089 (N_7089,N_5154,N_5099);
nor U7090 (N_7090,N_5172,N_4833);
and U7091 (N_7091,N_4615,N_5640);
nor U7092 (N_7092,N_5533,N_4771);
nor U7093 (N_7093,N_4574,N_5330);
xnor U7094 (N_7094,N_5820,N_5744);
nand U7095 (N_7095,N_5104,N_5089);
nor U7096 (N_7096,N_5351,N_5890);
or U7097 (N_7097,N_5297,N_5317);
nor U7098 (N_7098,N_5531,N_4521);
and U7099 (N_7099,N_4888,N_5922);
nor U7100 (N_7100,N_5702,N_5755);
nor U7101 (N_7101,N_4532,N_5070);
or U7102 (N_7102,N_5554,N_5960);
nor U7103 (N_7103,N_5506,N_5939);
nand U7104 (N_7104,N_5016,N_5264);
or U7105 (N_7105,N_5195,N_4740);
xor U7106 (N_7106,N_5030,N_5292);
nor U7107 (N_7107,N_5823,N_4705);
and U7108 (N_7108,N_4805,N_5405);
and U7109 (N_7109,N_5365,N_5471);
or U7110 (N_7110,N_5465,N_4957);
and U7111 (N_7111,N_4725,N_5174);
nor U7112 (N_7112,N_5035,N_4751);
or U7113 (N_7113,N_5239,N_5034);
nor U7114 (N_7114,N_4691,N_5450);
and U7115 (N_7115,N_5024,N_5691);
nand U7116 (N_7116,N_5136,N_5817);
and U7117 (N_7117,N_5125,N_5051);
nand U7118 (N_7118,N_5006,N_4773);
nor U7119 (N_7119,N_5882,N_5533);
nand U7120 (N_7120,N_5210,N_5829);
and U7121 (N_7121,N_5654,N_5238);
and U7122 (N_7122,N_4874,N_5544);
and U7123 (N_7123,N_5947,N_5152);
xnor U7124 (N_7124,N_5660,N_4994);
or U7125 (N_7125,N_4895,N_4512);
and U7126 (N_7126,N_5221,N_5590);
or U7127 (N_7127,N_4840,N_5203);
and U7128 (N_7128,N_5354,N_4516);
or U7129 (N_7129,N_4653,N_5120);
nand U7130 (N_7130,N_4515,N_5739);
or U7131 (N_7131,N_5116,N_5134);
and U7132 (N_7132,N_5866,N_5291);
or U7133 (N_7133,N_4655,N_5277);
nor U7134 (N_7134,N_5314,N_4613);
xnor U7135 (N_7135,N_4944,N_5766);
nor U7136 (N_7136,N_4777,N_4903);
xor U7137 (N_7137,N_5705,N_4729);
nor U7138 (N_7138,N_5837,N_5613);
and U7139 (N_7139,N_4916,N_5762);
nand U7140 (N_7140,N_5982,N_5768);
nor U7141 (N_7141,N_5551,N_5378);
nor U7142 (N_7142,N_5902,N_4996);
nor U7143 (N_7143,N_5538,N_4773);
or U7144 (N_7144,N_4837,N_5054);
and U7145 (N_7145,N_5306,N_5341);
and U7146 (N_7146,N_5736,N_4771);
nor U7147 (N_7147,N_5382,N_5499);
and U7148 (N_7148,N_5991,N_5423);
and U7149 (N_7149,N_5340,N_4825);
or U7150 (N_7150,N_4618,N_5007);
nor U7151 (N_7151,N_5320,N_4912);
nand U7152 (N_7152,N_5372,N_5738);
nor U7153 (N_7153,N_5552,N_5575);
xor U7154 (N_7154,N_4653,N_5810);
or U7155 (N_7155,N_5973,N_5728);
nand U7156 (N_7156,N_5488,N_5291);
nor U7157 (N_7157,N_5855,N_5558);
or U7158 (N_7158,N_5893,N_5189);
and U7159 (N_7159,N_5230,N_5701);
nand U7160 (N_7160,N_5641,N_5323);
xor U7161 (N_7161,N_5753,N_5128);
and U7162 (N_7162,N_4915,N_5465);
nand U7163 (N_7163,N_5985,N_4587);
or U7164 (N_7164,N_5060,N_5339);
nand U7165 (N_7165,N_5903,N_4938);
xor U7166 (N_7166,N_4843,N_5212);
xnor U7167 (N_7167,N_5256,N_5286);
xnor U7168 (N_7168,N_5817,N_4948);
and U7169 (N_7169,N_4918,N_5271);
or U7170 (N_7170,N_5552,N_4578);
and U7171 (N_7171,N_4657,N_5033);
or U7172 (N_7172,N_5919,N_5648);
and U7173 (N_7173,N_5761,N_4725);
nand U7174 (N_7174,N_4652,N_5325);
nand U7175 (N_7175,N_5634,N_5357);
and U7176 (N_7176,N_5605,N_5937);
and U7177 (N_7177,N_5108,N_5700);
xnor U7178 (N_7178,N_5795,N_5665);
and U7179 (N_7179,N_5231,N_5877);
or U7180 (N_7180,N_5930,N_5422);
nor U7181 (N_7181,N_4738,N_4916);
xor U7182 (N_7182,N_5660,N_5444);
nand U7183 (N_7183,N_5043,N_4599);
xor U7184 (N_7184,N_5968,N_5392);
nor U7185 (N_7185,N_5172,N_4932);
nor U7186 (N_7186,N_5103,N_5194);
nor U7187 (N_7187,N_4731,N_4970);
or U7188 (N_7188,N_5174,N_5395);
xnor U7189 (N_7189,N_4599,N_4606);
nand U7190 (N_7190,N_5838,N_4907);
and U7191 (N_7191,N_5726,N_5805);
nand U7192 (N_7192,N_5045,N_5524);
or U7193 (N_7193,N_5904,N_4707);
nand U7194 (N_7194,N_5706,N_5925);
nand U7195 (N_7195,N_5957,N_5976);
or U7196 (N_7196,N_4961,N_5341);
or U7197 (N_7197,N_4510,N_5949);
and U7198 (N_7198,N_5011,N_4790);
or U7199 (N_7199,N_5428,N_5298);
and U7200 (N_7200,N_5037,N_4685);
or U7201 (N_7201,N_5246,N_5494);
or U7202 (N_7202,N_4764,N_5402);
and U7203 (N_7203,N_4744,N_5965);
nand U7204 (N_7204,N_5470,N_5531);
nand U7205 (N_7205,N_5385,N_5931);
or U7206 (N_7206,N_5056,N_4850);
or U7207 (N_7207,N_4986,N_5312);
and U7208 (N_7208,N_5121,N_5350);
nor U7209 (N_7209,N_5274,N_4842);
and U7210 (N_7210,N_4866,N_4629);
and U7211 (N_7211,N_5323,N_5881);
nand U7212 (N_7212,N_4611,N_5826);
nand U7213 (N_7213,N_5247,N_5022);
nor U7214 (N_7214,N_5267,N_5348);
xnor U7215 (N_7215,N_5083,N_4641);
nor U7216 (N_7216,N_5806,N_4632);
nand U7217 (N_7217,N_5153,N_5884);
xnor U7218 (N_7218,N_5707,N_5635);
and U7219 (N_7219,N_4751,N_5702);
nand U7220 (N_7220,N_5066,N_5591);
nand U7221 (N_7221,N_4828,N_5238);
nand U7222 (N_7222,N_5942,N_5258);
nand U7223 (N_7223,N_5106,N_5329);
or U7224 (N_7224,N_5093,N_4614);
nand U7225 (N_7225,N_5340,N_5825);
and U7226 (N_7226,N_5612,N_5689);
xnor U7227 (N_7227,N_4645,N_5106);
nand U7228 (N_7228,N_5435,N_5408);
xor U7229 (N_7229,N_5182,N_5450);
nand U7230 (N_7230,N_5357,N_4637);
or U7231 (N_7231,N_5702,N_5573);
nor U7232 (N_7232,N_5865,N_4710);
nor U7233 (N_7233,N_5583,N_5676);
xnor U7234 (N_7234,N_4815,N_4824);
xnor U7235 (N_7235,N_4831,N_5576);
or U7236 (N_7236,N_5442,N_4853);
and U7237 (N_7237,N_5138,N_5615);
or U7238 (N_7238,N_5421,N_5967);
nand U7239 (N_7239,N_5067,N_5683);
xor U7240 (N_7240,N_4572,N_5613);
nand U7241 (N_7241,N_4503,N_5475);
nand U7242 (N_7242,N_5249,N_5286);
or U7243 (N_7243,N_5427,N_5975);
and U7244 (N_7244,N_4957,N_4620);
xnor U7245 (N_7245,N_5224,N_5861);
or U7246 (N_7246,N_5562,N_4624);
nand U7247 (N_7247,N_4846,N_4976);
and U7248 (N_7248,N_4764,N_5350);
nand U7249 (N_7249,N_5630,N_5621);
or U7250 (N_7250,N_4560,N_5237);
nor U7251 (N_7251,N_4677,N_5037);
xor U7252 (N_7252,N_5353,N_4965);
xnor U7253 (N_7253,N_5633,N_5388);
or U7254 (N_7254,N_4765,N_5752);
nor U7255 (N_7255,N_4510,N_4554);
nor U7256 (N_7256,N_5131,N_4565);
xor U7257 (N_7257,N_4777,N_4523);
and U7258 (N_7258,N_4986,N_5578);
nand U7259 (N_7259,N_5485,N_5642);
or U7260 (N_7260,N_5719,N_5137);
or U7261 (N_7261,N_5044,N_4703);
nor U7262 (N_7262,N_4780,N_5153);
xor U7263 (N_7263,N_4745,N_5252);
nand U7264 (N_7264,N_5277,N_4664);
xor U7265 (N_7265,N_4952,N_5574);
or U7266 (N_7266,N_4836,N_5332);
xnor U7267 (N_7267,N_5127,N_5896);
nand U7268 (N_7268,N_4810,N_4630);
xnor U7269 (N_7269,N_4841,N_4671);
xor U7270 (N_7270,N_4651,N_5642);
and U7271 (N_7271,N_4796,N_4745);
and U7272 (N_7272,N_4662,N_4812);
and U7273 (N_7273,N_5090,N_4603);
nor U7274 (N_7274,N_5352,N_4594);
and U7275 (N_7275,N_5104,N_5597);
and U7276 (N_7276,N_5036,N_4765);
nand U7277 (N_7277,N_5362,N_4853);
nand U7278 (N_7278,N_5789,N_4543);
and U7279 (N_7279,N_4520,N_5889);
nand U7280 (N_7280,N_5470,N_5848);
or U7281 (N_7281,N_5727,N_5556);
nand U7282 (N_7282,N_5166,N_4542);
and U7283 (N_7283,N_5621,N_5200);
and U7284 (N_7284,N_5890,N_5552);
nand U7285 (N_7285,N_4917,N_5037);
nor U7286 (N_7286,N_5736,N_5709);
nor U7287 (N_7287,N_5679,N_4813);
xor U7288 (N_7288,N_4882,N_5450);
and U7289 (N_7289,N_5467,N_5323);
nand U7290 (N_7290,N_5422,N_4892);
and U7291 (N_7291,N_4729,N_5940);
nand U7292 (N_7292,N_5662,N_5584);
or U7293 (N_7293,N_5942,N_4917);
nand U7294 (N_7294,N_4692,N_4864);
or U7295 (N_7295,N_5839,N_5005);
and U7296 (N_7296,N_5061,N_5833);
nand U7297 (N_7297,N_5109,N_4569);
nand U7298 (N_7298,N_5430,N_5136);
xor U7299 (N_7299,N_5042,N_5651);
nor U7300 (N_7300,N_5588,N_4503);
and U7301 (N_7301,N_5901,N_5491);
xor U7302 (N_7302,N_5220,N_4887);
xor U7303 (N_7303,N_4668,N_5537);
nand U7304 (N_7304,N_4886,N_4744);
nor U7305 (N_7305,N_5523,N_5231);
nand U7306 (N_7306,N_5358,N_5681);
nor U7307 (N_7307,N_5620,N_5909);
xnor U7308 (N_7308,N_4550,N_5613);
xnor U7309 (N_7309,N_4980,N_5213);
or U7310 (N_7310,N_5197,N_5605);
or U7311 (N_7311,N_4782,N_5076);
nand U7312 (N_7312,N_5697,N_4678);
nor U7313 (N_7313,N_5143,N_5121);
nor U7314 (N_7314,N_4808,N_5907);
and U7315 (N_7315,N_5690,N_4936);
nor U7316 (N_7316,N_5989,N_4567);
nor U7317 (N_7317,N_5222,N_4501);
and U7318 (N_7318,N_4877,N_5559);
or U7319 (N_7319,N_5673,N_5026);
or U7320 (N_7320,N_5174,N_5253);
or U7321 (N_7321,N_5173,N_4968);
xor U7322 (N_7322,N_5716,N_4815);
nor U7323 (N_7323,N_5187,N_4574);
nor U7324 (N_7324,N_5266,N_4916);
and U7325 (N_7325,N_5573,N_5530);
nor U7326 (N_7326,N_4974,N_4919);
and U7327 (N_7327,N_5082,N_5959);
nand U7328 (N_7328,N_5326,N_5586);
xor U7329 (N_7329,N_4808,N_5169);
or U7330 (N_7330,N_5729,N_4669);
nor U7331 (N_7331,N_5564,N_5245);
nand U7332 (N_7332,N_5966,N_5054);
nand U7333 (N_7333,N_5419,N_4962);
xnor U7334 (N_7334,N_4501,N_5915);
and U7335 (N_7335,N_5641,N_5530);
xor U7336 (N_7336,N_4508,N_4932);
nor U7337 (N_7337,N_5545,N_5488);
or U7338 (N_7338,N_5903,N_5668);
and U7339 (N_7339,N_5767,N_5317);
and U7340 (N_7340,N_5578,N_4884);
nor U7341 (N_7341,N_5977,N_5217);
or U7342 (N_7342,N_5953,N_4502);
nand U7343 (N_7343,N_5259,N_5323);
and U7344 (N_7344,N_5509,N_4580);
or U7345 (N_7345,N_5114,N_5513);
or U7346 (N_7346,N_4706,N_4771);
or U7347 (N_7347,N_4713,N_5793);
xnor U7348 (N_7348,N_5595,N_5014);
nand U7349 (N_7349,N_5771,N_4787);
and U7350 (N_7350,N_4851,N_5544);
xor U7351 (N_7351,N_4868,N_4978);
and U7352 (N_7352,N_5670,N_5192);
nor U7353 (N_7353,N_5158,N_5606);
nand U7354 (N_7354,N_5931,N_5026);
nand U7355 (N_7355,N_5724,N_5991);
and U7356 (N_7356,N_5425,N_5523);
nand U7357 (N_7357,N_5902,N_4908);
and U7358 (N_7358,N_5749,N_4543);
xnor U7359 (N_7359,N_5810,N_5905);
nor U7360 (N_7360,N_5080,N_4509);
nor U7361 (N_7361,N_4829,N_5354);
xor U7362 (N_7362,N_4674,N_4506);
nor U7363 (N_7363,N_5716,N_4905);
or U7364 (N_7364,N_5078,N_5297);
xnor U7365 (N_7365,N_4781,N_4623);
xor U7366 (N_7366,N_4542,N_5324);
xor U7367 (N_7367,N_4827,N_4970);
nand U7368 (N_7368,N_5385,N_5945);
nand U7369 (N_7369,N_5190,N_4865);
nor U7370 (N_7370,N_5690,N_5119);
or U7371 (N_7371,N_4973,N_5917);
nor U7372 (N_7372,N_5809,N_5983);
or U7373 (N_7373,N_4673,N_5409);
nand U7374 (N_7374,N_5652,N_5715);
or U7375 (N_7375,N_5824,N_5019);
and U7376 (N_7376,N_5346,N_5583);
xnor U7377 (N_7377,N_5093,N_5937);
or U7378 (N_7378,N_5496,N_4819);
nor U7379 (N_7379,N_5134,N_4611);
or U7380 (N_7380,N_4654,N_5877);
or U7381 (N_7381,N_5647,N_4971);
and U7382 (N_7382,N_5829,N_5275);
or U7383 (N_7383,N_5975,N_5419);
nand U7384 (N_7384,N_5973,N_4673);
xor U7385 (N_7385,N_5739,N_4821);
or U7386 (N_7386,N_5939,N_4504);
xnor U7387 (N_7387,N_5353,N_4857);
nor U7388 (N_7388,N_5510,N_4572);
nand U7389 (N_7389,N_5953,N_4650);
xor U7390 (N_7390,N_5834,N_5009);
or U7391 (N_7391,N_5911,N_4974);
xor U7392 (N_7392,N_5251,N_5716);
nand U7393 (N_7393,N_5171,N_5554);
or U7394 (N_7394,N_5754,N_4756);
nor U7395 (N_7395,N_4707,N_4590);
and U7396 (N_7396,N_5435,N_5635);
xor U7397 (N_7397,N_4556,N_5635);
or U7398 (N_7398,N_5437,N_5129);
nand U7399 (N_7399,N_4846,N_4948);
and U7400 (N_7400,N_5811,N_4636);
and U7401 (N_7401,N_5177,N_5999);
and U7402 (N_7402,N_4726,N_5830);
nand U7403 (N_7403,N_5351,N_5398);
and U7404 (N_7404,N_4991,N_4649);
and U7405 (N_7405,N_5978,N_4934);
and U7406 (N_7406,N_4764,N_5291);
nand U7407 (N_7407,N_5564,N_5109);
or U7408 (N_7408,N_5696,N_5077);
nor U7409 (N_7409,N_5237,N_5108);
and U7410 (N_7410,N_4872,N_4813);
nand U7411 (N_7411,N_5930,N_5871);
and U7412 (N_7412,N_4672,N_4762);
nor U7413 (N_7413,N_5793,N_5338);
xnor U7414 (N_7414,N_5731,N_5479);
nand U7415 (N_7415,N_5853,N_5032);
nor U7416 (N_7416,N_5288,N_5201);
or U7417 (N_7417,N_5057,N_4546);
or U7418 (N_7418,N_4857,N_5957);
nor U7419 (N_7419,N_5576,N_5575);
or U7420 (N_7420,N_4671,N_4585);
nor U7421 (N_7421,N_5010,N_5094);
xor U7422 (N_7422,N_4506,N_5682);
nor U7423 (N_7423,N_5986,N_5099);
nand U7424 (N_7424,N_5801,N_5791);
nand U7425 (N_7425,N_5426,N_5241);
nor U7426 (N_7426,N_4721,N_4838);
nor U7427 (N_7427,N_5736,N_4578);
nor U7428 (N_7428,N_5386,N_5493);
xnor U7429 (N_7429,N_5194,N_5981);
nand U7430 (N_7430,N_5638,N_5145);
or U7431 (N_7431,N_4543,N_5618);
or U7432 (N_7432,N_5818,N_5823);
and U7433 (N_7433,N_4612,N_5000);
xnor U7434 (N_7434,N_4938,N_4841);
nand U7435 (N_7435,N_5167,N_4877);
and U7436 (N_7436,N_5748,N_5362);
and U7437 (N_7437,N_5054,N_5847);
nand U7438 (N_7438,N_5287,N_5235);
or U7439 (N_7439,N_4852,N_5615);
nand U7440 (N_7440,N_5658,N_5788);
nor U7441 (N_7441,N_5491,N_5482);
nand U7442 (N_7442,N_5130,N_4595);
nor U7443 (N_7443,N_5037,N_5323);
and U7444 (N_7444,N_4551,N_5583);
nor U7445 (N_7445,N_5845,N_5636);
xor U7446 (N_7446,N_5183,N_5456);
or U7447 (N_7447,N_5253,N_5326);
xor U7448 (N_7448,N_5037,N_4965);
or U7449 (N_7449,N_5582,N_4945);
and U7450 (N_7450,N_5487,N_5163);
nor U7451 (N_7451,N_5501,N_5365);
or U7452 (N_7452,N_5727,N_5668);
xor U7453 (N_7453,N_5114,N_5873);
or U7454 (N_7454,N_4815,N_4568);
xnor U7455 (N_7455,N_5137,N_4689);
xnor U7456 (N_7456,N_4857,N_5341);
and U7457 (N_7457,N_5634,N_5761);
nor U7458 (N_7458,N_4701,N_5100);
nor U7459 (N_7459,N_4926,N_5210);
or U7460 (N_7460,N_4823,N_5535);
xnor U7461 (N_7461,N_4623,N_5100);
and U7462 (N_7462,N_5223,N_5682);
xor U7463 (N_7463,N_4585,N_4784);
nor U7464 (N_7464,N_5825,N_4602);
nand U7465 (N_7465,N_5248,N_5497);
or U7466 (N_7466,N_5473,N_5318);
and U7467 (N_7467,N_5601,N_4783);
or U7468 (N_7468,N_5456,N_5625);
or U7469 (N_7469,N_5063,N_5546);
and U7470 (N_7470,N_4570,N_5768);
nor U7471 (N_7471,N_5999,N_5970);
xor U7472 (N_7472,N_5109,N_5852);
nand U7473 (N_7473,N_5959,N_5320);
or U7474 (N_7474,N_5485,N_5916);
nand U7475 (N_7475,N_5311,N_5011);
nand U7476 (N_7476,N_5619,N_5071);
or U7477 (N_7477,N_4552,N_5165);
and U7478 (N_7478,N_5245,N_5021);
nor U7479 (N_7479,N_5164,N_5473);
xor U7480 (N_7480,N_5402,N_5263);
or U7481 (N_7481,N_5100,N_4947);
xor U7482 (N_7482,N_5296,N_4814);
or U7483 (N_7483,N_5941,N_4528);
or U7484 (N_7484,N_5831,N_4525);
or U7485 (N_7485,N_5499,N_5605);
nor U7486 (N_7486,N_4649,N_4667);
and U7487 (N_7487,N_5853,N_4679);
nand U7488 (N_7488,N_5064,N_5454);
nor U7489 (N_7489,N_4922,N_5753);
and U7490 (N_7490,N_5324,N_5033);
or U7491 (N_7491,N_5678,N_5460);
nor U7492 (N_7492,N_5169,N_5951);
or U7493 (N_7493,N_4896,N_5084);
nor U7494 (N_7494,N_5410,N_4709);
or U7495 (N_7495,N_5554,N_4658);
nor U7496 (N_7496,N_4944,N_5650);
or U7497 (N_7497,N_5674,N_5107);
and U7498 (N_7498,N_5366,N_5245);
nand U7499 (N_7499,N_5374,N_4646);
nor U7500 (N_7500,N_6308,N_7126);
xor U7501 (N_7501,N_6521,N_7132);
and U7502 (N_7502,N_6944,N_6495);
nand U7503 (N_7503,N_6823,N_6479);
xor U7504 (N_7504,N_6474,N_7210);
and U7505 (N_7505,N_7227,N_6936);
and U7506 (N_7506,N_6703,N_6131);
and U7507 (N_7507,N_6425,N_7116);
and U7508 (N_7508,N_6814,N_6824);
nand U7509 (N_7509,N_6300,N_6546);
nand U7510 (N_7510,N_6890,N_7193);
or U7511 (N_7511,N_6625,N_7347);
xnor U7512 (N_7512,N_7389,N_6203);
nand U7513 (N_7513,N_6607,N_7283);
xor U7514 (N_7514,N_6841,N_6340);
or U7515 (N_7515,N_7084,N_6385);
or U7516 (N_7516,N_7370,N_6424);
nand U7517 (N_7517,N_7120,N_7329);
nand U7518 (N_7518,N_6247,N_6181);
nand U7519 (N_7519,N_6827,N_6342);
nor U7520 (N_7520,N_6820,N_6948);
and U7521 (N_7521,N_7432,N_6293);
xor U7522 (N_7522,N_6929,N_6579);
nor U7523 (N_7523,N_7065,N_7266);
xor U7524 (N_7524,N_7160,N_7056);
xor U7525 (N_7525,N_6162,N_6576);
xor U7526 (N_7526,N_6624,N_7268);
nor U7527 (N_7527,N_6485,N_6160);
xor U7528 (N_7528,N_6808,N_7143);
xnor U7529 (N_7529,N_7038,N_7427);
nand U7530 (N_7530,N_7294,N_6518);
or U7531 (N_7531,N_6063,N_6784);
xnor U7532 (N_7532,N_7484,N_7149);
nor U7533 (N_7533,N_6013,N_6436);
xnor U7534 (N_7534,N_7040,N_7241);
nand U7535 (N_7535,N_6403,N_6573);
nand U7536 (N_7536,N_6834,N_6122);
nand U7537 (N_7537,N_6646,N_6561);
xnor U7538 (N_7538,N_6431,N_6962);
and U7539 (N_7539,N_6807,N_6527);
nor U7540 (N_7540,N_6652,N_6678);
nand U7541 (N_7541,N_7097,N_7032);
or U7542 (N_7542,N_7343,N_6075);
and U7543 (N_7543,N_6639,N_7360);
and U7544 (N_7544,N_6269,N_6898);
nand U7545 (N_7545,N_6391,N_7248);
nor U7546 (N_7546,N_6679,N_6006);
nor U7547 (N_7547,N_6360,N_7047);
nor U7548 (N_7548,N_6884,N_7170);
nor U7549 (N_7549,N_6701,N_7220);
nand U7550 (N_7550,N_6610,N_7141);
and U7551 (N_7551,N_7224,N_7453);
nor U7552 (N_7552,N_6535,N_7437);
nor U7553 (N_7553,N_6438,N_6531);
and U7554 (N_7554,N_6344,N_6888);
and U7555 (N_7555,N_6174,N_7277);
nor U7556 (N_7556,N_7489,N_6037);
or U7557 (N_7557,N_7014,N_6088);
xnor U7558 (N_7558,N_6106,N_6294);
nand U7559 (N_7559,N_7113,N_6314);
xnor U7560 (N_7560,N_7420,N_6484);
or U7561 (N_7561,N_7273,N_6802);
and U7562 (N_7562,N_6583,N_6178);
xor U7563 (N_7563,N_6341,N_6675);
nand U7564 (N_7564,N_7192,N_6567);
nand U7565 (N_7565,N_6502,N_7185);
or U7566 (N_7566,N_6614,N_7336);
or U7567 (N_7567,N_7001,N_7302);
and U7568 (N_7568,N_7445,N_6722);
or U7569 (N_7569,N_7181,N_6061);
or U7570 (N_7570,N_6907,N_7184);
nor U7571 (N_7571,N_7304,N_6992);
xor U7572 (N_7572,N_7042,N_7150);
or U7573 (N_7573,N_7317,N_6249);
or U7574 (N_7574,N_7234,N_6477);
xnor U7575 (N_7575,N_6400,N_7109);
xnor U7576 (N_7576,N_6872,N_6040);
nor U7577 (N_7577,N_6685,N_7173);
nor U7578 (N_7578,N_6121,N_7371);
and U7579 (N_7579,N_7095,N_6497);
xor U7580 (N_7580,N_6971,N_7121);
xor U7581 (N_7581,N_6961,N_6564);
or U7582 (N_7582,N_6533,N_6970);
nor U7583 (N_7583,N_7478,N_6832);
and U7584 (N_7584,N_7088,N_6292);
xnor U7585 (N_7585,N_6669,N_6661);
or U7586 (N_7586,N_6470,N_6141);
nand U7587 (N_7587,N_6592,N_7286);
nand U7588 (N_7588,N_6738,N_7275);
nand U7589 (N_7589,N_6829,N_6411);
nand U7590 (N_7590,N_7418,N_6838);
nand U7591 (N_7591,N_6885,N_7467);
and U7592 (N_7592,N_6705,N_6361);
or U7593 (N_7593,N_7493,N_6167);
xnor U7594 (N_7594,N_6440,N_6598);
nor U7595 (N_7595,N_7009,N_6241);
or U7596 (N_7596,N_6966,N_6672);
nor U7597 (N_7597,N_6018,N_7479);
nor U7598 (N_7598,N_6983,N_6645);
nand U7599 (N_7599,N_6336,N_6822);
xnor U7600 (N_7600,N_6761,N_6316);
or U7601 (N_7601,N_6654,N_6156);
nand U7602 (N_7602,N_6605,N_6151);
and U7603 (N_7603,N_6083,N_6111);
nor U7604 (N_7604,N_6955,N_6641);
and U7605 (N_7605,N_7069,N_6007);
or U7606 (N_7606,N_6041,N_6472);
or U7607 (N_7607,N_6124,N_6954);
or U7608 (N_7608,N_6956,N_6878);
and U7609 (N_7609,N_6916,N_7450);
nor U7610 (N_7610,N_6544,N_7213);
and U7611 (N_7611,N_6603,N_6370);
or U7612 (N_7612,N_6519,N_7378);
or U7613 (N_7613,N_6109,N_6259);
nand U7614 (N_7614,N_6875,N_6305);
nor U7615 (N_7615,N_6159,N_6500);
and U7616 (N_7616,N_6777,N_6723);
and U7617 (N_7617,N_6538,N_7357);
nand U7618 (N_7618,N_7481,N_6800);
and U7619 (N_7619,N_6771,N_6132);
and U7620 (N_7620,N_6831,N_7480);
nor U7621 (N_7621,N_6504,N_6190);
and U7622 (N_7622,N_6825,N_7298);
nand U7623 (N_7623,N_7147,N_6959);
nand U7624 (N_7624,N_6127,N_6999);
or U7625 (N_7625,N_6346,N_6200);
xor U7626 (N_7626,N_6317,N_6067);
nor U7627 (N_7627,N_6450,N_7279);
and U7628 (N_7628,N_6096,N_6478);
or U7629 (N_7629,N_7183,N_6804);
or U7630 (N_7630,N_6599,N_6666);
and U7631 (N_7631,N_7233,N_7440);
and U7632 (N_7632,N_6756,N_7247);
xor U7633 (N_7633,N_6942,N_6819);
nand U7634 (N_7634,N_6523,N_6307);
or U7635 (N_7635,N_7071,N_6996);
and U7636 (N_7636,N_6322,N_7319);
and U7637 (N_7637,N_6560,N_6941);
nor U7638 (N_7638,N_6285,N_7171);
nand U7639 (N_7639,N_6489,N_6882);
nor U7640 (N_7640,N_6731,N_6613);
nor U7641 (N_7641,N_7444,N_6860);
and U7642 (N_7642,N_7242,N_6036);
nor U7643 (N_7643,N_6866,N_7118);
nand U7644 (N_7644,N_7216,N_6301);
nor U7645 (N_7645,N_6099,N_7020);
nand U7646 (N_7646,N_6422,N_6304);
nand U7647 (N_7647,N_6023,N_7383);
and U7648 (N_7648,N_6806,N_6094);
or U7649 (N_7649,N_6911,N_6445);
or U7650 (N_7650,N_7063,N_6208);
and U7651 (N_7651,N_6539,N_6619);
or U7652 (N_7652,N_7498,N_6781);
xnor U7653 (N_7653,N_6228,N_6321);
xor U7654 (N_7654,N_7203,N_7293);
and U7655 (N_7655,N_6343,N_7413);
and U7656 (N_7656,N_6015,N_6278);
and U7657 (N_7657,N_7359,N_6821);
and U7658 (N_7658,N_6125,N_7259);
nand U7659 (N_7659,N_7442,N_7491);
or U7660 (N_7660,N_6656,N_6810);
and U7661 (N_7661,N_6812,N_6056);
nor U7662 (N_7662,N_7180,N_7195);
nor U7663 (N_7663,N_6998,N_6437);
xnor U7664 (N_7664,N_6967,N_6152);
xor U7665 (N_7665,N_6442,N_6380);
nor U7666 (N_7666,N_7340,N_6526);
nor U7667 (N_7667,N_7376,N_6853);
or U7668 (N_7668,N_6651,N_6997);
nor U7669 (N_7669,N_6760,N_7243);
xor U7670 (N_7670,N_6615,N_6356);
nor U7671 (N_7671,N_7494,N_7175);
or U7672 (N_7672,N_6930,N_7240);
or U7673 (N_7673,N_6862,N_6170);
nand U7674 (N_7674,N_6295,N_6648);
xor U7675 (N_7675,N_7265,N_6904);
xnor U7676 (N_7676,N_6443,N_6530);
or U7677 (N_7677,N_6662,N_6813);
or U7678 (N_7678,N_7154,N_7236);
nand U7679 (N_7679,N_6766,N_6367);
xnor U7680 (N_7680,N_6745,N_7153);
or U7681 (N_7681,N_7305,N_7096);
xor U7682 (N_7682,N_7252,N_7261);
and U7683 (N_7683,N_7198,N_6274);
and U7684 (N_7684,N_6177,N_7475);
nand U7685 (N_7685,N_7177,N_6382);
nor U7686 (N_7686,N_7139,N_7111);
nand U7687 (N_7687,N_7404,N_6076);
nor U7688 (N_7688,N_6691,N_6548);
xnor U7689 (N_7689,N_6011,N_6318);
nor U7690 (N_7690,N_7060,N_6359);
or U7691 (N_7691,N_6388,N_6226);
or U7692 (N_7692,N_6906,N_6009);
nand U7693 (N_7693,N_6782,N_6892);
or U7694 (N_7694,N_7366,N_6505);
nor U7695 (N_7695,N_7310,N_6287);
and U7696 (N_7696,N_6501,N_6010);
nand U7697 (N_7697,N_7375,N_6179);
and U7698 (N_7698,N_6569,N_6871);
xnor U7699 (N_7699,N_7300,N_6325);
xor U7700 (N_7700,N_6065,N_7140);
nor U7701 (N_7701,N_7188,N_6284);
nand U7702 (N_7702,N_6078,N_6846);
or U7703 (N_7703,N_6503,N_6237);
nor U7704 (N_7704,N_6345,N_6665);
and U7705 (N_7705,N_6951,N_6586);
or U7706 (N_7706,N_6275,N_7209);
nor U7707 (N_7707,N_6271,N_7356);
nor U7708 (N_7708,N_6401,N_6187);
nand U7709 (N_7709,N_7382,N_6323);
or U7710 (N_7710,N_6864,N_6702);
xor U7711 (N_7711,N_6138,N_6005);
or U7712 (N_7712,N_6608,N_6975);
nand U7713 (N_7713,N_6414,N_6748);
nor U7714 (N_7714,N_7422,N_6326);
nor U7715 (N_7715,N_7219,N_6577);
and U7716 (N_7716,N_6147,N_6676);
xor U7717 (N_7717,N_6606,N_7278);
xnor U7718 (N_7718,N_7023,N_6555);
and U7719 (N_7719,N_6987,N_6550);
nand U7720 (N_7720,N_6357,N_6534);
xnor U7721 (N_7721,N_7022,N_6729);
nand U7722 (N_7722,N_6462,N_7428);
nor U7723 (N_7723,N_6309,N_7411);
nand U7724 (N_7724,N_6223,N_6339);
nand U7725 (N_7725,N_6466,N_7007);
nand U7726 (N_7726,N_6260,N_6815);
or U7727 (N_7727,N_6498,N_6254);
nand U7728 (N_7728,N_6195,N_7098);
and U7729 (N_7729,N_6783,N_7030);
nor U7730 (N_7730,N_6769,N_6054);
xnor U7731 (N_7731,N_7301,N_6673);
nor U7732 (N_7732,N_6937,N_6427);
nor U7733 (N_7733,N_6115,N_6517);
nand U7734 (N_7734,N_6256,N_7064);
nor U7735 (N_7735,N_7256,N_6587);
and U7736 (N_7736,N_6158,N_6710);
and U7737 (N_7737,N_6939,N_6420);
xnor U7738 (N_7738,N_6704,N_6390);
xnor U7739 (N_7739,N_6716,N_6404);
xor U7740 (N_7740,N_7439,N_7331);
xnor U7741 (N_7741,N_6303,N_6394);
and U7742 (N_7742,N_6994,N_6488);
nand U7743 (N_7743,N_6621,N_7372);
nand U7744 (N_7744,N_6328,N_7362);
and U7745 (N_7745,N_7080,N_7441);
and U7746 (N_7746,N_6383,N_6737);
nor U7747 (N_7747,N_7018,N_6628);
xnor U7748 (N_7748,N_7401,N_6778);
and U7749 (N_7749,N_6508,N_6847);
xor U7750 (N_7750,N_6296,N_6989);
nor U7751 (N_7751,N_6407,N_6413);
nand U7752 (N_7752,N_6978,N_6507);
nand U7753 (N_7753,N_6644,N_7367);
xnor U7754 (N_7754,N_6059,N_6713);
xnor U7755 (N_7755,N_6446,N_7017);
nand U7756 (N_7756,N_7045,N_6012);
or U7757 (N_7757,N_6626,N_7206);
or U7758 (N_7758,N_7041,N_6454);
and U7759 (N_7759,N_6842,N_6135);
and U7760 (N_7760,N_6312,N_7276);
or U7761 (N_7761,N_6025,N_6331);
nand U7762 (N_7762,N_6288,N_6042);
and U7763 (N_7763,N_7267,N_6611);
and U7764 (N_7764,N_6191,N_7258);
nand U7765 (N_7765,N_7215,N_6110);
nor U7766 (N_7766,N_7464,N_6578);
xnor U7767 (N_7767,N_7090,N_6092);
or U7768 (N_7768,N_6381,N_7281);
and U7769 (N_7769,N_6168,N_6868);
xnor U7770 (N_7770,N_6212,N_7204);
or U7771 (N_7771,N_7386,N_7076);
nor U7772 (N_7772,N_6055,N_7390);
xnor U7773 (N_7773,N_6019,N_7434);
xnor U7774 (N_7774,N_7391,N_6789);
and U7775 (N_7775,N_6248,N_6492);
xnor U7776 (N_7776,N_6302,N_7159);
nor U7777 (N_7777,N_6686,N_6522);
xnor U7778 (N_7778,N_6395,N_6483);
nor U7779 (N_7779,N_6620,N_6355);
xor U7780 (N_7780,N_6140,N_7388);
or U7781 (N_7781,N_6844,N_7462);
and U7782 (N_7782,N_6974,N_6843);
nor U7783 (N_7783,N_7353,N_6683);
nand U7784 (N_7784,N_6165,N_6750);
and U7785 (N_7785,N_6245,N_6684);
or U7786 (N_7786,N_7110,N_6148);
or U7787 (N_7787,N_6799,N_6857);
nand U7788 (N_7788,N_7469,N_6034);
nand U7789 (N_7789,N_6496,N_7100);
nor U7790 (N_7790,N_6313,N_6150);
nor U7791 (N_7791,N_6351,N_6920);
and U7792 (N_7792,N_6108,N_6876);
nand U7793 (N_7793,N_6718,N_6874);
or U7794 (N_7794,N_7449,N_6246);
nand U7795 (N_7795,N_6338,N_6752);
nor U7796 (N_7796,N_6755,N_6856);
or U7797 (N_7797,N_6643,N_7324);
nand U7798 (N_7798,N_6883,N_6163);
xor U7799 (N_7799,N_6664,N_7218);
nand U7800 (N_7800,N_7237,N_7196);
or U7801 (N_7801,N_7456,N_6708);
nor U7802 (N_7802,N_7130,N_6103);
nand U7803 (N_7803,N_6044,N_6139);
or U7804 (N_7804,N_7037,N_6744);
nor U7805 (N_7805,N_7131,N_6185);
nand U7806 (N_7806,N_6243,N_6952);
xor U7807 (N_7807,N_6870,N_6696);
nand U7808 (N_7808,N_7146,N_6765);
nor U7809 (N_7809,N_7482,N_6028);
nand U7810 (N_7810,N_6933,N_6528);
xnor U7811 (N_7811,N_7158,N_6811);
xnor U7812 (N_7812,N_7322,N_6144);
xor U7813 (N_7813,N_6085,N_6353);
nand U7814 (N_7814,N_6739,N_6008);
and U7815 (N_7815,N_7054,N_6659);
nor U7816 (N_7816,N_6617,N_6213);
and U7817 (N_7817,N_6358,N_6051);
nor U7818 (N_7818,N_6238,N_6236);
and U7819 (N_7819,N_6963,N_6095);
and U7820 (N_7820,N_6764,N_7006);
or U7821 (N_7821,N_6277,N_6297);
nor U7822 (N_7822,N_6120,N_6969);
nand U7823 (N_7823,N_6255,N_6244);
nor U7824 (N_7824,N_6128,N_6430);
nor U7825 (N_7825,N_7168,N_6220);
xor U7826 (N_7826,N_6923,N_6917);
or U7827 (N_7827,N_7191,N_6889);
xor U7828 (N_7828,N_6219,N_7239);
and U7829 (N_7829,N_6362,N_6682);
nor U7830 (N_7830,N_6572,N_6197);
nor U7831 (N_7831,N_6184,N_6020);
nand U7832 (N_7832,N_7034,N_6779);
xor U7833 (N_7833,N_6230,N_7392);
or U7834 (N_7834,N_7308,N_6670);
nand U7835 (N_7835,N_6428,N_7485);
and U7836 (N_7836,N_6104,N_6973);
xnor U7837 (N_7837,N_6235,N_7472);
xor U7838 (N_7838,N_7395,N_6721);
or U7839 (N_7839,N_6393,N_7202);
and U7840 (N_7840,N_7232,N_6867);
xor U7841 (N_7841,N_7446,N_7291);
and U7842 (N_7842,N_7048,N_6218);
nor U7843 (N_7843,N_6455,N_6692);
nor U7844 (N_7844,N_6102,N_7142);
or U7845 (N_7845,N_6444,N_6833);
or U7846 (N_7846,N_6263,N_7074);
xnor U7847 (N_7847,N_6563,N_7174);
or U7848 (N_7848,N_6689,N_6227);
and U7849 (N_7849,N_6240,N_7089);
nand U7850 (N_7850,N_6082,N_6196);
and U7851 (N_7851,N_6137,N_6554);
or U7852 (N_7852,N_6986,N_6460);
and U7853 (N_7853,N_7374,N_7355);
xor U7854 (N_7854,N_7245,N_7156);
or U7855 (N_7855,N_7409,N_6946);
nand U7856 (N_7856,N_7026,N_6232);
and U7857 (N_7857,N_6928,N_6027);
or U7858 (N_7858,N_7398,N_7393);
or U7859 (N_7859,N_6902,N_6596);
or U7860 (N_7860,N_7035,N_6369);
xnor U7861 (N_7861,N_6387,N_7468);
xor U7862 (N_7862,N_7421,N_7315);
nand U7863 (N_7863,N_6283,N_7321);
nand U7864 (N_7864,N_6105,N_6189);
xor U7865 (N_7865,N_6133,N_6014);
nand U7866 (N_7866,N_6529,N_6024);
or U7867 (N_7867,N_7024,N_7194);
or U7868 (N_7868,N_7137,N_6419);
xnor U7869 (N_7869,N_6153,N_6298);
xnor U7870 (N_7870,N_6273,N_6052);
nand U7871 (N_7871,N_6582,N_6629);
and U7872 (N_7872,N_7414,N_6049);
nand U7873 (N_7873,N_6536,N_7499);
or U7874 (N_7874,N_7000,N_7410);
nand U7875 (N_7875,N_6927,N_6775);
xor U7876 (N_7876,N_6965,N_7358);
nand U7877 (N_7877,N_7086,N_6145);
xnor U7878 (N_7878,N_7263,N_6396);
and U7879 (N_7879,N_7186,N_6727);
and U7880 (N_7880,N_6861,N_6757);
nand U7881 (N_7881,N_7260,N_6788);
xor U7882 (N_7882,N_6439,N_7036);
or U7883 (N_7883,N_6215,N_7112);
nor U7884 (N_7884,N_7029,N_6638);
nand U7885 (N_7885,N_7226,N_6932);
nor U7886 (N_7886,N_7495,N_6461);
and U7887 (N_7887,N_7458,N_6524);
xor U7888 (N_7888,N_7270,N_6406);
nor U7889 (N_7889,N_6222,N_6199);
and U7890 (N_7890,N_6224,N_7309);
nand U7891 (N_7891,N_6491,N_6979);
or U7892 (N_7892,N_7162,N_6217);
xor U7893 (N_7893,N_6934,N_7429);
nor U7894 (N_7894,N_6943,N_6216);
or U7895 (N_7895,N_6402,N_6229);
nand U7896 (N_7896,N_7052,N_7062);
nand U7897 (N_7897,N_6657,N_6903);
nor U7898 (N_7898,N_6734,N_7039);
and U7899 (N_7899,N_7028,N_6711);
nand U7900 (N_7900,N_6398,N_7461);
nand U7901 (N_7901,N_6633,N_6073);
nor U7902 (N_7902,N_7083,N_7345);
or U7903 (N_7903,N_6330,N_6805);
and U7904 (N_7904,N_7323,N_6149);
or U7905 (N_7905,N_6749,N_7046);
nor U7906 (N_7906,N_7115,N_7399);
nand U7907 (N_7907,N_6763,N_6730);
nor U7908 (N_7908,N_7051,N_6901);
or U7909 (N_7909,N_7043,N_7463);
and U7910 (N_7910,N_7369,N_6677);
nor U7911 (N_7911,N_6960,N_6060);
xnor U7912 (N_7912,N_7314,N_7125);
xor U7913 (N_7913,N_7151,N_7107);
or U7914 (N_7914,N_6949,N_6801);
or U7915 (N_7915,N_6840,N_6851);
nor U7916 (N_7916,N_6604,N_6794);
nand U7917 (N_7917,N_6887,N_7405);
nand U7918 (N_7918,N_6003,N_6264);
xor U7919 (N_7919,N_7417,N_7249);
or U7920 (N_7920,N_6558,N_7246);
and U7921 (N_7921,N_6270,N_6743);
nor U7922 (N_7922,N_6706,N_7161);
nand U7923 (N_7923,N_7280,N_7471);
xor U7924 (N_7924,N_7406,N_6225);
and U7925 (N_7925,N_6335,N_7199);
nor U7926 (N_7926,N_6354,N_6627);
xnor U7927 (N_7927,N_6206,N_6129);
and U7928 (N_7928,N_7274,N_6134);
and U7929 (N_7929,N_6091,N_6242);
and U7930 (N_7930,N_7128,N_6089);
nor U7931 (N_7931,N_6707,N_7465);
nor U7932 (N_7932,N_7012,N_7403);
xnor U7933 (N_7933,N_6559,N_6035);
xor U7934 (N_7934,N_7368,N_6116);
xnor U7935 (N_7935,N_6026,N_7416);
or U7936 (N_7936,N_6276,N_6631);
and U7937 (N_7937,N_6977,N_6058);
nor U7938 (N_7938,N_6113,N_6557);
and U7939 (N_7939,N_7200,N_6421);
xnor U7940 (N_7940,N_7313,N_6568);
nor U7941 (N_7941,N_7459,N_6376);
or U7942 (N_7942,N_6033,N_6205);
or U7943 (N_7943,N_7497,N_6595);
or U7944 (N_7944,N_7033,N_6077);
nand U7945 (N_7945,N_6668,N_6057);
nand U7946 (N_7946,N_6409,N_6112);
nand U7947 (N_7947,N_6551,N_6725);
and U7948 (N_7948,N_6506,N_6623);
xnor U7949 (N_7949,N_6087,N_7373);
xor U7950 (N_7950,N_6310,N_6451);
and U7951 (N_7951,N_7238,N_6995);
and U7952 (N_7952,N_6712,N_7172);
nor U7953 (N_7953,N_7425,N_6021);
xor U7954 (N_7954,N_6173,N_6740);
nand U7955 (N_7955,N_7316,N_6570);
nor U7956 (N_7956,N_6311,N_7148);
nand U7957 (N_7957,N_7257,N_6459);
nand U7958 (N_7958,N_6597,N_6649);
nand U7959 (N_7959,N_6733,N_6982);
or U7960 (N_7960,N_7225,N_6798);
and U7961 (N_7961,N_7067,N_6251);
nor U7962 (N_7962,N_7134,N_7169);
and U7963 (N_7963,N_7282,N_7189);
nor U7964 (N_7964,N_6650,N_6981);
or U7965 (N_7965,N_7483,N_6732);
nor U7966 (N_7966,N_6791,N_6826);
or U7967 (N_7967,N_6990,N_6392);
or U7968 (N_7968,N_6365,N_7288);
xor U7969 (N_7969,N_6797,N_7307);
xor U7970 (N_7970,N_7073,N_6976);
nor U7971 (N_7971,N_7122,N_6796);
nor U7972 (N_7972,N_7338,N_6250);
or U7973 (N_7973,N_7119,N_6130);
nand U7974 (N_7974,N_7025,N_6803);
nor U7975 (N_7975,N_7106,N_6768);
nand U7976 (N_7976,N_6945,N_6588);
xor U7977 (N_7977,N_7460,N_6896);
xor U7978 (N_7978,N_6457,N_6647);
nor U7979 (N_7979,N_6787,N_6154);
nand U7980 (N_7980,N_7136,N_6584);
xnor U7981 (N_7981,N_7127,N_6327);
xor U7982 (N_7982,N_6473,N_6386);
nand U7983 (N_7983,N_6658,N_7351);
nand U7984 (N_7984,N_6537,N_6886);
or U7985 (N_7985,N_6046,N_6622);
and U7986 (N_7986,N_6281,N_6581);
and U7987 (N_7987,N_7470,N_6201);
and U7988 (N_7988,N_6741,N_7223);
xor U7989 (N_7989,N_7473,N_6449);
or U7990 (N_7990,N_6912,N_7190);
nor U7991 (N_7991,N_7443,N_6728);
nor U7992 (N_7992,N_6107,N_7474);
nand U7993 (N_7993,N_7075,N_6333);
and U7994 (N_7994,N_6532,N_7438);
and U7995 (N_7995,N_6922,N_6002);
or U7996 (N_7996,N_6183,N_6816);
nor U7997 (N_7997,N_6039,N_6332);
nand U7998 (N_7998,N_6836,N_7003);
and U7999 (N_7999,N_6835,N_6947);
nand U8000 (N_8000,N_6435,N_6265);
and U8001 (N_8001,N_6211,N_6742);
nor U8002 (N_8002,N_6074,N_7342);
or U8003 (N_8003,N_7004,N_6634);
and U8004 (N_8004,N_6324,N_6257);
nor U8005 (N_8005,N_7105,N_6467);
or U8006 (N_8006,N_7423,N_7490);
or U8007 (N_8007,N_7002,N_6786);
xnor U8008 (N_8008,N_6931,N_6510);
nand U8009 (N_8009,N_7400,N_6231);
nor U8010 (N_8010,N_7235,N_7452);
xnor U8011 (N_8011,N_7292,N_6198);
nor U8012 (N_8012,N_6695,N_7448);
nand U8013 (N_8013,N_6543,N_7320);
or U8014 (N_8014,N_7253,N_7167);
nor U8015 (N_8015,N_7212,N_6416);
nand U8016 (N_8016,N_7208,N_6900);
xor U8017 (N_8017,N_6100,N_6136);
nand U8018 (N_8018,N_7229,N_7031);
nand U8019 (N_8019,N_6958,N_7250);
and U8020 (N_8020,N_6758,N_6207);
xor U8021 (N_8021,N_6031,N_6809);
nand U8022 (N_8022,N_7070,N_6188);
nor U8023 (N_8023,N_6192,N_6594);
or U8024 (N_8024,N_6865,N_6253);
and U8025 (N_8025,N_7436,N_6566);
xnor U8026 (N_8026,N_6751,N_6378);
and U8027 (N_8027,N_7015,N_7092);
and U8028 (N_8028,N_6509,N_6935);
xor U8029 (N_8029,N_6897,N_7165);
nand U8030 (N_8030,N_6452,N_6855);
nor U8031 (N_8031,N_7197,N_7117);
xnor U8032 (N_8032,N_6291,N_7312);
or U8033 (N_8033,N_6770,N_6698);
and U8034 (N_8034,N_7059,N_7005);
nor U8035 (N_8035,N_6541,N_6098);
xnor U8036 (N_8036,N_6925,N_6379);
and U8037 (N_8037,N_7330,N_6368);
xnor U8038 (N_8038,N_6571,N_6690);
nor U8039 (N_8039,N_6363,N_6688);
and U8040 (N_8040,N_6038,N_6877);
xnor U8041 (N_8041,N_6182,N_6221);
nand U8042 (N_8042,N_7387,N_7055);
nor U8043 (N_8043,N_6166,N_6795);
nand U8044 (N_8044,N_7447,N_6540);
xnor U8045 (N_8045,N_7103,N_6146);
or U8046 (N_8046,N_6792,N_7094);
nor U8047 (N_8047,N_7454,N_6204);
nor U8048 (N_8048,N_6123,N_6893);
nand U8049 (N_8049,N_6482,N_6453);
nand U8050 (N_8050,N_6456,N_7272);
nor U8051 (N_8051,N_6352,N_6516);
or U8052 (N_8052,N_6985,N_6372);
xnor U8053 (N_8053,N_6029,N_6319);
nor U8054 (N_8054,N_6697,N_7164);
xor U8055 (N_8055,N_6016,N_6410);
or U8056 (N_8056,N_6371,N_7027);
or U8057 (N_8057,N_6556,N_6938);
nor U8058 (N_8058,N_6434,N_7102);
nor U8059 (N_8059,N_6609,N_6043);
or U8060 (N_8060,N_7157,N_7021);
nand U8061 (N_8061,N_6515,N_7211);
nor U8062 (N_8062,N_7010,N_6653);
or U8063 (N_8063,N_6774,N_7166);
or U8064 (N_8064,N_6193,N_6234);
and U8065 (N_8065,N_6412,N_7396);
nor U8066 (N_8066,N_6680,N_6417);
or U8067 (N_8067,N_6926,N_6261);
or U8068 (N_8068,N_6047,N_7214);
nand U8069 (N_8069,N_7016,N_6064);
or U8070 (N_8070,N_7299,N_7077);
or U8071 (N_8071,N_6171,N_6881);
or U8072 (N_8072,N_7486,N_6924);
and U8073 (N_8073,N_7087,N_7081);
xnor U8074 (N_8074,N_6674,N_6914);
nor U8075 (N_8075,N_6848,N_7327);
or U8076 (N_8076,N_6908,N_6289);
nand U8077 (N_8077,N_7344,N_7431);
xor U8078 (N_8078,N_6919,N_7085);
or U8079 (N_8079,N_6334,N_7101);
and U8080 (N_8080,N_7455,N_7492);
xor U8081 (N_8081,N_7496,N_6950);
and U8082 (N_8082,N_7019,N_6001);
nand U8083 (N_8083,N_6717,N_7244);
or U8084 (N_8084,N_6418,N_7044);
and U8085 (N_8085,N_6397,N_6667);
nor U8086 (N_8086,N_6180,N_6299);
xnor U8087 (N_8087,N_6616,N_6636);
or U8088 (N_8088,N_6172,N_7326);
or U8089 (N_8089,N_7104,N_6048);
nor U8090 (N_8090,N_6290,N_6004);
or U8091 (N_8091,N_6337,N_7114);
nand U8092 (N_8092,N_6348,N_6772);
nand U8093 (N_8093,N_6859,N_7361);
nor U8094 (N_8094,N_7144,N_6895);
xor U8095 (N_8095,N_6545,N_7078);
or U8096 (N_8096,N_7341,N_6030);
nand U8097 (N_8097,N_6681,N_6957);
nor U8098 (N_8098,N_6767,N_6852);
nand U8099 (N_8099,N_6066,N_6580);
nor U8100 (N_8100,N_7011,N_6441);
nor U8101 (N_8101,N_7380,N_7207);
or U8102 (N_8102,N_7108,N_6699);
and U8103 (N_8103,N_6918,N_6186);
nor U8104 (N_8104,N_6858,N_7008);
nand U8105 (N_8105,N_6854,N_6164);
or U8106 (N_8106,N_6377,N_6017);
or U8107 (N_8107,N_7384,N_6280);
nor U8108 (N_8108,N_6086,N_6547);
xnor U8109 (N_8109,N_7066,N_6475);
xnor U8110 (N_8110,N_7264,N_6693);
xor U8111 (N_8111,N_6079,N_6828);
and U8112 (N_8112,N_6873,N_6565);
nor U8113 (N_8113,N_6991,N_7337);
nand U8114 (N_8114,N_6481,N_7050);
and U8115 (N_8115,N_6214,N_6593);
xnor U8116 (N_8116,N_6081,N_7426);
or U8117 (N_8117,N_7217,N_6754);
xnor U8118 (N_8118,N_6719,N_6347);
nor U8119 (N_8119,N_6084,N_6575);
nand U8120 (N_8120,N_7093,N_6426);
xor U8121 (N_8121,N_6118,N_7350);
xnor U8122 (N_8122,N_6097,N_6562);
nor U8123 (N_8123,N_6655,N_7349);
or U8124 (N_8124,N_7295,N_7124);
or U8125 (N_8125,N_6709,N_7332);
or U8126 (N_8126,N_6252,N_6493);
and U8127 (N_8127,N_6469,N_7402);
nor U8128 (N_8128,N_6239,N_7352);
nand U8129 (N_8129,N_7364,N_7231);
and U8130 (N_8130,N_6790,N_6511);
nand U8131 (N_8131,N_6759,N_6155);
and U8132 (N_8132,N_6630,N_6433);
nor U8133 (N_8133,N_6642,N_6349);
or U8134 (N_8134,N_6793,N_7271);
nand U8135 (N_8135,N_6487,N_6818);
or U8136 (N_8136,N_6429,N_6940);
and U8137 (N_8137,N_6905,N_6589);
xor U8138 (N_8138,N_6964,N_6785);
or U8139 (N_8139,N_7289,N_6161);
nand U8140 (N_8140,N_7269,N_7079);
nor U8141 (N_8141,N_7339,N_6090);
or U8142 (N_8142,N_6458,N_6753);
xnor U8143 (N_8143,N_7487,N_7412);
nand U8144 (N_8144,N_6830,N_6069);
nand U8145 (N_8145,N_7335,N_6762);
nand U8146 (N_8146,N_6968,N_7251);
xnor U8147 (N_8147,N_6585,N_7379);
xor U8148 (N_8148,N_7049,N_6032);
nor U8149 (N_8149,N_6471,N_7287);
and U8150 (N_8150,N_6549,N_7222);
nand U8151 (N_8151,N_7285,N_7201);
or U8152 (N_8152,N_6724,N_6476);
nand U8153 (N_8153,N_6663,N_6045);
nor U8154 (N_8154,N_6415,N_6080);
nand U8155 (N_8155,N_6845,N_6817);
or U8156 (N_8156,N_7053,N_7419);
nand U8157 (N_8157,N_7397,N_7230);
nor U8158 (N_8158,N_7430,N_7178);
or U8159 (N_8159,N_7072,N_6490);
nor U8160 (N_8160,N_6700,N_6746);
nor U8161 (N_8161,N_6447,N_6542);
and U8162 (N_8162,N_6169,N_6117);
or U8163 (N_8163,N_6910,N_6175);
xnor U8164 (N_8164,N_7082,N_6715);
xnor U8165 (N_8165,N_6720,N_7433);
nor U8166 (N_8166,N_7254,N_6464);
nor U8167 (N_8167,N_6880,N_6913);
xnor U8168 (N_8168,N_6726,N_6773);
nand U8169 (N_8169,N_6574,N_6101);
xor U8170 (N_8170,N_6022,N_6465);
and U8171 (N_8171,N_6119,N_6389);
or U8172 (N_8172,N_6863,N_6590);
and U8173 (N_8173,N_6494,N_7488);
and U8174 (N_8174,N_6268,N_7290);
or U8175 (N_8175,N_7068,N_6747);
nor U8176 (N_8176,N_6513,N_6209);
or U8177 (N_8177,N_6072,N_6176);
or U8178 (N_8178,N_7091,N_6839);
xor U8179 (N_8179,N_6909,N_7182);
and U8180 (N_8180,N_7129,N_6736);
nor U8181 (N_8181,N_6000,N_6071);
nor U8182 (N_8182,N_6618,N_6448);
and U8183 (N_8183,N_6525,N_6068);
xor U8184 (N_8184,N_7328,N_7381);
xnor U8185 (N_8185,N_6694,N_7325);
and U8186 (N_8186,N_7179,N_6408);
xnor U8187 (N_8187,N_6849,N_6374);
nor U8188 (N_8188,N_6687,N_7163);
and U8189 (N_8189,N_7013,N_6921);
or U8190 (N_8190,N_6258,N_6350);
xnor U8191 (N_8191,N_6660,N_6306);
and U8192 (N_8192,N_6635,N_7407);
nand U8193 (N_8193,N_7138,N_6202);
and U8194 (N_8194,N_6062,N_6993);
nand U8195 (N_8195,N_6602,N_6267);
nor U8196 (N_8196,N_6514,N_7451);
xnor U8197 (N_8197,N_7346,N_6266);
nand U8198 (N_8198,N_7435,N_6735);
nand U8199 (N_8199,N_7123,N_6972);
nor U8200 (N_8200,N_6601,N_6480);
and U8201 (N_8201,N_7457,N_7221);
or U8202 (N_8202,N_7415,N_6591);
nor U8203 (N_8203,N_7187,N_6714);
nand U8204 (N_8204,N_7377,N_7099);
nand U8205 (N_8205,N_6315,N_6988);
or U8206 (N_8206,N_6637,N_6282);
and U8207 (N_8207,N_6114,N_7365);
nor U8208 (N_8208,N_7348,N_6612);
nand U8209 (N_8209,N_6953,N_7152);
or U8210 (N_8210,N_6375,N_6272);
and U8211 (N_8211,N_6233,N_7145);
xnor U8212 (N_8212,N_6210,N_7318);
xor U8213 (N_8213,N_7424,N_6486);
nand U8214 (N_8214,N_6142,N_7058);
nor U8215 (N_8215,N_7477,N_7297);
and U8216 (N_8216,N_6837,N_6194);
nor U8217 (N_8217,N_6405,N_6286);
or U8218 (N_8218,N_6671,N_6632);
nor U8219 (N_8219,N_6384,N_6329);
or U8220 (N_8220,N_7262,N_6423);
nand U8221 (N_8221,N_6553,N_7255);
nor U8222 (N_8222,N_6980,N_7303);
nor U8223 (N_8223,N_6869,N_6850);
and U8224 (N_8224,N_6780,N_6600);
and U8225 (N_8225,N_7155,N_6891);
nor U8226 (N_8226,N_6899,N_6552);
nand U8227 (N_8227,N_6984,N_6915);
xnor U8228 (N_8228,N_6432,N_7057);
nor U8229 (N_8229,N_7176,N_7334);
xor U8230 (N_8230,N_6050,N_7228);
and U8231 (N_8231,N_7296,N_6320);
or U8232 (N_8232,N_6640,N_7385);
or U8233 (N_8233,N_6364,N_7135);
nand U8234 (N_8234,N_6053,N_6399);
and U8235 (N_8235,N_6499,N_6512);
and U8236 (N_8236,N_6366,N_7408);
and U8237 (N_8237,N_6093,N_6070);
nor U8238 (N_8238,N_7205,N_7133);
and U8239 (N_8239,N_7306,N_6262);
xnor U8240 (N_8240,N_6143,N_6126);
or U8241 (N_8241,N_6894,N_7061);
and U8242 (N_8242,N_7466,N_7333);
nor U8243 (N_8243,N_7394,N_6879);
and U8244 (N_8244,N_6776,N_7476);
nor U8245 (N_8245,N_6463,N_6157);
or U8246 (N_8246,N_7354,N_7284);
xor U8247 (N_8247,N_6373,N_7311);
nor U8248 (N_8248,N_6279,N_6468);
xor U8249 (N_8249,N_6520,N_7363);
and U8250 (N_8250,N_6683,N_6498);
nor U8251 (N_8251,N_6934,N_6050);
xnor U8252 (N_8252,N_7256,N_7472);
and U8253 (N_8253,N_7300,N_6970);
and U8254 (N_8254,N_6173,N_6178);
nand U8255 (N_8255,N_7197,N_7428);
xnor U8256 (N_8256,N_7146,N_7280);
xnor U8257 (N_8257,N_6711,N_6308);
nand U8258 (N_8258,N_6492,N_6273);
or U8259 (N_8259,N_6292,N_6726);
nand U8260 (N_8260,N_6776,N_6278);
and U8261 (N_8261,N_6046,N_7172);
or U8262 (N_8262,N_6338,N_6989);
nor U8263 (N_8263,N_7013,N_7042);
xnor U8264 (N_8264,N_6880,N_6983);
or U8265 (N_8265,N_7426,N_6830);
nor U8266 (N_8266,N_7404,N_6588);
xor U8267 (N_8267,N_7113,N_6385);
nand U8268 (N_8268,N_6338,N_7241);
and U8269 (N_8269,N_6211,N_6899);
nor U8270 (N_8270,N_6241,N_6868);
nand U8271 (N_8271,N_6715,N_6143);
or U8272 (N_8272,N_6863,N_7165);
nor U8273 (N_8273,N_6577,N_6734);
or U8274 (N_8274,N_6198,N_6852);
and U8275 (N_8275,N_6799,N_6786);
nand U8276 (N_8276,N_6920,N_6627);
nand U8277 (N_8277,N_7386,N_6396);
or U8278 (N_8278,N_7356,N_7375);
nor U8279 (N_8279,N_6682,N_6681);
nor U8280 (N_8280,N_7345,N_6730);
nor U8281 (N_8281,N_7184,N_6977);
and U8282 (N_8282,N_6655,N_7395);
and U8283 (N_8283,N_6637,N_6343);
nor U8284 (N_8284,N_6509,N_6285);
nor U8285 (N_8285,N_6113,N_7299);
xor U8286 (N_8286,N_6288,N_6978);
nand U8287 (N_8287,N_6133,N_6168);
nor U8288 (N_8288,N_6399,N_6909);
nor U8289 (N_8289,N_6829,N_7422);
or U8290 (N_8290,N_6935,N_6519);
xor U8291 (N_8291,N_7006,N_7125);
or U8292 (N_8292,N_6690,N_7331);
nor U8293 (N_8293,N_6559,N_7087);
xor U8294 (N_8294,N_7248,N_6072);
xnor U8295 (N_8295,N_7472,N_6779);
or U8296 (N_8296,N_6326,N_6123);
xnor U8297 (N_8297,N_7218,N_6705);
xnor U8298 (N_8298,N_6271,N_7319);
xor U8299 (N_8299,N_6480,N_7251);
nor U8300 (N_8300,N_6303,N_6829);
nand U8301 (N_8301,N_7441,N_7438);
nor U8302 (N_8302,N_7313,N_6957);
xor U8303 (N_8303,N_6377,N_7371);
nor U8304 (N_8304,N_6511,N_7234);
or U8305 (N_8305,N_6331,N_6593);
or U8306 (N_8306,N_7463,N_7119);
and U8307 (N_8307,N_6425,N_7289);
nor U8308 (N_8308,N_6622,N_6946);
nand U8309 (N_8309,N_6202,N_6630);
and U8310 (N_8310,N_6980,N_7426);
and U8311 (N_8311,N_6121,N_7181);
nand U8312 (N_8312,N_6126,N_6370);
xnor U8313 (N_8313,N_6196,N_7128);
and U8314 (N_8314,N_6312,N_7110);
xor U8315 (N_8315,N_7145,N_6324);
nand U8316 (N_8316,N_6834,N_7220);
or U8317 (N_8317,N_6854,N_6217);
and U8318 (N_8318,N_6327,N_6633);
nor U8319 (N_8319,N_6063,N_6942);
and U8320 (N_8320,N_6234,N_6685);
or U8321 (N_8321,N_6887,N_7293);
or U8322 (N_8322,N_6745,N_6392);
xnor U8323 (N_8323,N_6032,N_6988);
nor U8324 (N_8324,N_6113,N_6264);
nor U8325 (N_8325,N_6615,N_6083);
nand U8326 (N_8326,N_7233,N_6697);
xor U8327 (N_8327,N_6101,N_7284);
nor U8328 (N_8328,N_6993,N_6261);
xnor U8329 (N_8329,N_7192,N_6853);
nor U8330 (N_8330,N_7268,N_7422);
and U8331 (N_8331,N_6331,N_6548);
nor U8332 (N_8332,N_6429,N_6811);
nor U8333 (N_8333,N_7131,N_6573);
nand U8334 (N_8334,N_6687,N_6118);
and U8335 (N_8335,N_6529,N_6474);
nand U8336 (N_8336,N_6194,N_7216);
nor U8337 (N_8337,N_6374,N_6696);
xor U8338 (N_8338,N_7370,N_6956);
xor U8339 (N_8339,N_7442,N_7492);
or U8340 (N_8340,N_6366,N_6813);
and U8341 (N_8341,N_6520,N_6877);
and U8342 (N_8342,N_6658,N_7478);
xnor U8343 (N_8343,N_7425,N_7383);
nand U8344 (N_8344,N_7293,N_6767);
nand U8345 (N_8345,N_6874,N_7341);
or U8346 (N_8346,N_6361,N_7137);
and U8347 (N_8347,N_6748,N_6610);
xor U8348 (N_8348,N_7208,N_6299);
nand U8349 (N_8349,N_7127,N_6201);
and U8350 (N_8350,N_6531,N_7402);
xnor U8351 (N_8351,N_7106,N_7059);
or U8352 (N_8352,N_6952,N_6608);
nor U8353 (N_8353,N_6117,N_7290);
or U8354 (N_8354,N_6138,N_6599);
nor U8355 (N_8355,N_7050,N_6483);
nor U8356 (N_8356,N_6889,N_6092);
and U8357 (N_8357,N_7160,N_6002);
and U8358 (N_8358,N_7464,N_6776);
and U8359 (N_8359,N_6677,N_7400);
nor U8360 (N_8360,N_6367,N_7155);
nand U8361 (N_8361,N_7182,N_6683);
nand U8362 (N_8362,N_6827,N_6277);
xor U8363 (N_8363,N_6285,N_7203);
nor U8364 (N_8364,N_6589,N_7205);
xnor U8365 (N_8365,N_6303,N_6211);
nor U8366 (N_8366,N_6705,N_6993);
nor U8367 (N_8367,N_7224,N_7130);
or U8368 (N_8368,N_7435,N_6484);
nand U8369 (N_8369,N_6943,N_7129);
nor U8370 (N_8370,N_6880,N_7125);
nand U8371 (N_8371,N_6839,N_6202);
xnor U8372 (N_8372,N_6793,N_7129);
xor U8373 (N_8373,N_6779,N_6869);
nand U8374 (N_8374,N_7072,N_7498);
nor U8375 (N_8375,N_7329,N_6336);
nand U8376 (N_8376,N_6718,N_6935);
and U8377 (N_8377,N_6568,N_6782);
or U8378 (N_8378,N_6901,N_6487);
nand U8379 (N_8379,N_7114,N_6914);
nand U8380 (N_8380,N_6879,N_6851);
nand U8381 (N_8381,N_7031,N_7394);
xnor U8382 (N_8382,N_7497,N_6616);
and U8383 (N_8383,N_7393,N_6992);
nand U8384 (N_8384,N_6901,N_6632);
xnor U8385 (N_8385,N_7049,N_7358);
or U8386 (N_8386,N_7311,N_6795);
xor U8387 (N_8387,N_7104,N_6481);
xor U8388 (N_8388,N_6435,N_6410);
nand U8389 (N_8389,N_6174,N_6146);
or U8390 (N_8390,N_7490,N_7165);
nor U8391 (N_8391,N_6148,N_6183);
and U8392 (N_8392,N_7043,N_6289);
nand U8393 (N_8393,N_6899,N_6637);
nor U8394 (N_8394,N_6322,N_6278);
nor U8395 (N_8395,N_7438,N_6250);
nor U8396 (N_8396,N_6185,N_6615);
nand U8397 (N_8397,N_7258,N_7467);
xnor U8398 (N_8398,N_6471,N_7354);
or U8399 (N_8399,N_6758,N_7272);
nor U8400 (N_8400,N_7022,N_6839);
and U8401 (N_8401,N_7093,N_7020);
or U8402 (N_8402,N_6066,N_6400);
or U8403 (N_8403,N_6469,N_6090);
and U8404 (N_8404,N_6734,N_6994);
xor U8405 (N_8405,N_6043,N_6856);
nand U8406 (N_8406,N_6752,N_6309);
xor U8407 (N_8407,N_6093,N_7365);
nor U8408 (N_8408,N_6676,N_6628);
or U8409 (N_8409,N_7112,N_7169);
and U8410 (N_8410,N_6393,N_6133);
nor U8411 (N_8411,N_7155,N_7033);
nand U8412 (N_8412,N_6550,N_7286);
nor U8413 (N_8413,N_6562,N_7228);
nor U8414 (N_8414,N_7210,N_7366);
and U8415 (N_8415,N_6649,N_7289);
or U8416 (N_8416,N_7474,N_7481);
nor U8417 (N_8417,N_6055,N_6394);
nor U8418 (N_8418,N_7056,N_6807);
nand U8419 (N_8419,N_7177,N_6275);
and U8420 (N_8420,N_6797,N_6360);
nand U8421 (N_8421,N_6248,N_6409);
nor U8422 (N_8422,N_7203,N_6247);
and U8423 (N_8423,N_6522,N_6600);
nor U8424 (N_8424,N_6037,N_6551);
and U8425 (N_8425,N_7322,N_7126);
and U8426 (N_8426,N_7052,N_6106);
and U8427 (N_8427,N_6730,N_6587);
or U8428 (N_8428,N_6809,N_7184);
nand U8429 (N_8429,N_6435,N_6994);
nor U8430 (N_8430,N_6369,N_6850);
xor U8431 (N_8431,N_7221,N_6945);
nand U8432 (N_8432,N_7104,N_6644);
xor U8433 (N_8433,N_6141,N_6247);
xnor U8434 (N_8434,N_7116,N_7426);
and U8435 (N_8435,N_6607,N_7180);
nor U8436 (N_8436,N_7366,N_6332);
or U8437 (N_8437,N_6477,N_6422);
nor U8438 (N_8438,N_7025,N_7033);
and U8439 (N_8439,N_7086,N_6935);
nand U8440 (N_8440,N_7446,N_7198);
nor U8441 (N_8441,N_7296,N_6518);
and U8442 (N_8442,N_7481,N_6649);
nor U8443 (N_8443,N_7270,N_6345);
or U8444 (N_8444,N_7300,N_6522);
xor U8445 (N_8445,N_6222,N_6548);
xnor U8446 (N_8446,N_7404,N_6897);
nor U8447 (N_8447,N_6561,N_6195);
nand U8448 (N_8448,N_6001,N_6486);
or U8449 (N_8449,N_6862,N_6897);
nand U8450 (N_8450,N_6656,N_6596);
xnor U8451 (N_8451,N_7095,N_7038);
or U8452 (N_8452,N_6320,N_7195);
nand U8453 (N_8453,N_6127,N_6758);
and U8454 (N_8454,N_7086,N_6901);
and U8455 (N_8455,N_6724,N_7150);
nor U8456 (N_8456,N_6722,N_6248);
or U8457 (N_8457,N_7195,N_7347);
nand U8458 (N_8458,N_7246,N_6446);
nand U8459 (N_8459,N_6351,N_7094);
xor U8460 (N_8460,N_7376,N_6791);
nor U8461 (N_8461,N_7169,N_6063);
xor U8462 (N_8462,N_6011,N_7482);
xnor U8463 (N_8463,N_6010,N_6653);
nor U8464 (N_8464,N_7407,N_7369);
or U8465 (N_8465,N_6287,N_6838);
and U8466 (N_8466,N_7143,N_6034);
and U8467 (N_8467,N_6176,N_7265);
xor U8468 (N_8468,N_6252,N_6469);
xor U8469 (N_8469,N_7331,N_7072);
nor U8470 (N_8470,N_6805,N_6848);
or U8471 (N_8471,N_6512,N_7228);
xor U8472 (N_8472,N_6630,N_6330);
or U8473 (N_8473,N_6885,N_6878);
xnor U8474 (N_8474,N_6809,N_6590);
nand U8475 (N_8475,N_6587,N_7475);
xor U8476 (N_8476,N_6027,N_7082);
nand U8477 (N_8477,N_6091,N_6477);
nand U8478 (N_8478,N_6546,N_7321);
or U8479 (N_8479,N_7424,N_7335);
and U8480 (N_8480,N_6095,N_6623);
nor U8481 (N_8481,N_6249,N_6048);
xor U8482 (N_8482,N_6110,N_6949);
and U8483 (N_8483,N_7312,N_6382);
and U8484 (N_8484,N_6689,N_6986);
nor U8485 (N_8485,N_6816,N_6176);
nand U8486 (N_8486,N_6157,N_7082);
or U8487 (N_8487,N_6651,N_7415);
nor U8488 (N_8488,N_6283,N_6737);
nor U8489 (N_8489,N_6218,N_6586);
xnor U8490 (N_8490,N_6816,N_6193);
xor U8491 (N_8491,N_6947,N_6884);
or U8492 (N_8492,N_6059,N_6564);
nand U8493 (N_8493,N_6478,N_7150);
xnor U8494 (N_8494,N_7196,N_6922);
xor U8495 (N_8495,N_6001,N_6848);
or U8496 (N_8496,N_7144,N_7054);
and U8497 (N_8497,N_7300,N_6230);
nor U8498 (N_8498,N_7348,N_6980);
nand U8499 (N_8499,N_6297,N_6465);
nor U8500 (N_8500,N_7142,N_6137);
xor U8501 (N_8501,N_6922,N_6954);
xor U8502 (N_8502,N_7417,N_7316);
or U8503 (N_8503,N_6101,N_6770);
nand U8504 (N_8504,N_6473,N_6718);
and U8505 (N_8505,N_6728,N_6962);
xor U8506 (N_8506,N_7382,N_6912);
nor U8507 (N_8507,N_6013,N_6705);
and U8508 (N_8508,N_6401,N_6928);
xor U8509 (N_8509,N_7409,N_6052);
and U8510 (N_8510,N_7045,N_6811);
nor U8511 (N_8511,N_6487,N_6760);
nand U8512 (N_8512,N_7427,N_7085);
nand U8513 (N_8513,N_6326,N_7416);
nor U8514 (N_8514,N_7109,N_7172);
nor U8515 (N_8515,N_7436,N_6662);
or U8516 (N_8516,N_6196,N_6337);
nor U8517 (N_8517,N_6286,N_6514);
xor U8518 (N_8518,N_6751,N_6859);
xnor U8519 (N_8519,N_7199,N_6371);
and U8520 (N_8520,N_7148,N_6208);
nor U8521 (N_8521,N_6780,N_6145);
nor U8522 (N_8522,N_7231,N_6693);
nand U8523 (N_8523,N_6339,N_6358);
nand U8524 (N_8524,N_7369,N_7040);
xnor U8525 (N_8525,N_6498,N_7310);
and U8526 (N_8526,N_6414,N_6117);
nor U8527 (N_8527,N_6696,N_6513);
or U8528 (N_8528,N_7146,N_6400);
nand U8529 (N_8529,N_6485,N_6230);
or U8530 (N_8530,N_6385,N_6883);
xnor U8531 (N_8531,N_6298,N_7041);
nor U8532 (N_8532,N_6768,N_6244);
or U8533 (N_8533,N_7121,N_6759);
and U8534 (N_8534,N_7192,N_7425);
nand U8535 (N_8535,N_6776,N_6746);
and U8536 (N_8536,N_6993,N_6701);
or U8537 (N_8537,N_6236,N_6992);
and U8538 (N_8538,N_6490,N_6513);
nor U8539 (N_8539,N_7449,N_6123);
and U8540 (N_8540,N_6040,N_6455);
or U8541 (N_8541,N_6328,N_7131);
and U8542 (N_8542,N_6994,N_6776);
or U8543 (N_8543,N_6923,N_7414);
and U8544 (N_8544,N_6463,N_6927);
and U8545 (N_8545,N_6939,N_6892);
or U8546 (N_8546,N_7381,N_6685);
and U8547 (N_8547,N_7081,N_6712);
xor U8548 (N_8548,N_6952,N_6422);
and U8549 (N_8549,N_6084,N_6517);
nand U8550 (N_8550,N_7010,N_6994);
xnor U8551 (N_8551,N_6944,N_6008);
and U8552 (N_8552,N_6570,N_7226);
nand U8553 (N_8553,N_6007,N_6487);
or U8554 (N_8554,N_7010,N_6615);
xnor U8555 (N_8555,N_6031,N_6294);
nand U8556 (N_8556,N_6524,N_6414);
nor U8557 (N_8557,N_6185,N_7474);
nor U8558 (N_8558,N_6477,N_6089);
and U8559 (N_8559,N_6105,N_7171);
nand U8560 (N_8560,N_6849,N_7236);
or U8561 (N_8561,N_6292,N_6082);
or U8562 (N_8562,N_7367,N_6819);
or U8563 (N_8563,N_7031,N_6110);
xnor U8564 (N_8564,N_6411,N_7255);
nand U8565 (N_8565,N_6104,N_6621);
and U8566 (N_8566,N_6542,N_6051);
or U8567 (N_8567,N_7224,N_6345);
nand U8568 (N_8568,N_7093,N_7288);
xnor U8569 (N_8569,N_6314,N_7083);
xor U8570 (N_8570,N_6862,N_6711);
nor U8571 (N_8571,N_6634,N_6217);
nor U8572 (N_8572,N_7473,N_7372);
nor U8573 (N_8573,N_7311,N_6622);
or U8574 (N_8574,N_6597,N_6688);
or U8575 (N_8575,N_7298,N_6059);
nand U8576 (N_8576,N_6754,N_6884);
nor U8577 (N_8577,N_7332,N_6017);
nand U8578 (N_8578,N_7299,N_7106);
and U8579 (N_8579,N_7205,N_6901);
or U8580 (N_8580,N_6189,N_6603);
or U8581 (N_8581,N_6406,N_6817);
and U8582 (N_8582,N_6014,N_6299);
nand U8583 (N_8583,N_7497,N_6243);
xnor U8584 (N_8584,N_6187,N_6404);
and U8585 (N_8585,N_6816,N_6391);
xor U8586 (N_8586,N_7337,N_7255);
nand U8587 (N_8587,N_7364,N_6246);
xnor U8588 (N_8588,N_6202,N_6176);
nor U8589 (N_8589,N_7219,N_6836);
xor U8590 (N_8590,N_7027,N_6223);
and U8591 (N_8591,N_6372,N_7287);
nand U8592 (N_8592,N_6427,N_6847);
xnor U8593 (N_8593,N_7214,N_6940);
or U8594 (N_8594,N_6257,N_6066);
xnor U8595 (N_8595,N_6522,N_7097);
xnor U8596 (N_8596,N_6657,N_7263);
and U8597 (N_8597,N_6612,N_7179);
nand U8598 (N_8598,N_6382,N_6777);
xnor U8599 (N_8599,N_6564,N_6318);
xnor U8600 (N_8600,N_6027,N_7319);
or U8601 (N_8601,N_6946,N_7320);
nor U8602 (N_8602,N_6297,N_7071);
nor U8603 (N_8603,N_6138,N_7137);
and U8604 (N_8604,N_6335,N_6298);
xor U8605 (N_8605,N_7266,N_6630);
or U8606 (N_8606,N_6843,N_7391);
and U8607 (N_8607,N_6917,N_6238);
xnor U8608 (N_8608,N_6589,N_6899);
and U8609 (N_8609,N_7048,N_6361);
or U8610 (N_8610,N_7145,N_6792);
or U8611 (N_8611,N_6224,N_6754);
nor U8612 (N_8612,N_6995,N_7284);
nand U8613 (N_8613,N_6723,N_6363);
xor U8614 (N_8614,N_6990,N_6019);
nand U8615 (N_8615,N_6879,N_7272);
or U8616 (N_8616,N_7201,N_7063);
nand U8617 (N_8617,N_6224,N_7194);
and U8618 (N_8618,N_7205,N_7096);
and U8619 (N_8619,N_6249,N_7457);
or U8620 (N_8620,N_6597,N_6809);
and U8621 (N_8621,N_6581,N_6380);
xor U8622 (N_8622,N_7032,N_7129);
xor U8623 (N_8623,N_6384,N_7250);
nor U8624 (N_8624,N_6354,N_6063);
nor U8625 (N_8625,N_7314,N_6296);
nand U8626 (N_8626,N_7257,N_6952);
or U8627 (N_8627,N_6124,N_6064);
or U8628 (N_8628,N_6076,N_6429);
and U8629 (N_8629,N_6437,N_6394);
or U8630 (N_8630,N_6608,N_6616);
nor U8631 (N_8631,N_6016,N_6199);
nor U8632 (N_8632,N_6956,N_6048);
or U8633 (N_8633,N_7412,N_7006);
or U8634 (N_8634,N_6927,N_7104);
nand U8635 (N_8635,N_6506,N_7362);
nand U8636 (N_8636,N_6811,N_7457);
or U8637 (N_8637,N_6945,N_6369);
xor U8638 (N_8638,N_7239,N_7037);
nand U8639 (N_8639,N_7007,N_6859);
nor U8640 (N_8640,N_6788,N_6668);
nor U8641 (N_8641,N_7050,N_6086);
nand U8642 (N_8642,N_6256,N_7392);
xor U8643 (N_8643,N_7043,N_6702);
and U8644 (N_8644,N_7270,N_6140);
xnor U8645 (N_8645,N_6562,N_7359);
nand U8646 (N_8646,N_6677,N_6348);
or U8647 (N_8647,N_6521,N_6554);
xor U8648 (N_8648,N_6101,N_7015);
nor U8649 (N_8649,N_7293,N_6047);
nor U8650 (N_8650,N_6597,N_6647);
and U8651 (N_8651,N_6730,N_6488);
nand U8652 (N_8652,N_6555,N_7440);
nor U8653 (N_8653,N_6510,N_6860);
and U8654 (N_8654,N_7034,N_6227);
or U8655 (N_8655,N_6285,N_7304);
and U8656 (N_8656,N_7280,N_6408);
and U8657 (N_8657,N_7006,N_7309);
and U8658 (N_8658,N_6497,N_6416);
nor U8659 (N_8659,N_6622,N_7149);
or U8660 (N_8660,N_7438,N_6467);
xnor U8661 (N_8661,N_6430,N_6844);
nand U8662 (N_8662,N_6255,N_6373);
and U8663 (N_8663,N_7266,N_6081);
nand U8664 (N_8664,N_7315,N_7328);
or U8665 (N_8665,N_6272,N_7335);
and U8666 (N_8666,N_6366,N_6585);
xnor U8667 (N_8667,N_6138,N_6875);
or U8668 (N_8668,N_6283,N_7315);
xnor U8669 (N_8669,N_7417,N_7455);
nand U8670 (N_8670,N_6863,N_6106);
xor U8671 (N_8671,N_7098,N_7091);
or U8672 (N_8672,N_7075,N_7009);
or U8673 (N_8673,N_7132,N_6319);
and U8674 (N_8674,N_6572,N_7155);
xnor U8675 (N_8675,N_6703,N_6905);
nor U8676 (N_8676,N_7141,N_6558);
nand U8677 (N_8677,N_6646,N_6616);
and U8678 (N_8678,N_6825,N_6632);
and U8679 (N_8679,N_6367,N_6523);
and U8680 (N_8680,N_6858,N_6084);
or U8681 (N_8681,N_7390,N_7363);
nor U8682 (N_8682,N_7193,N_7322);
xnor U8683 (N_8683,N_6063,N_6206);
nand U8684 (N_8684,N_6750,N_7209);
nand U8685 (N_8685,N_7446,N_6783);
and U8686 (N_8686,N_7035,N_6194);
and U8687 (N_8687,N_6808,N_7311);
nand U8688 (N_8688,N_7157,N_7370);
nand U8689 (N_8689,N_6754,N_6560);
and U8690 (N_8690,N_6257,N_6771);
xor U8691 (N_8691,N_6576,N_7462);
or U8692 (N_8692,N_6102,N_6772);
nor U8693 (N_8693,N_7426,N_6292);
and U8694 (N_8694,N_7391,N_6424);
nor U8695 (N_8695,N_6040,N_6653);
or U8696 (N_8696,N_6049,N_6466);
xor U8697 (N_8697,N_6555,N_6009);
nand U8698 (N_8698,N_7375,N_6710);
nor U8699 (N_8699,N_6834,N_7131);
and U8700 (N_8700,N_6325,N_6205);
or U8701 (N_8701,N_7245,N_6079);
xnor U8702 (N_8702,N_7105,N_6737);
and U8703 (N_8703,N_6069,N_7197);
nand U8704 (N_8704,N_6935,N_6422);
nand U8705 (N_8705,N_7227,N_6236);
xor U8706 (N_8706,N_6406,N_7162);
and U8707 (N_8707,N_6259,N_6540);
or U8708 (N_8708,N_7415,N_7330);
nand U8709 (N_8709,N_6553,N_6598);
or U8710 (N_8710,N_6264,N_6300);
and U8711 (N_8711,N_6089,N_7029);
or U8712 (N_8712,N_6878,N_6445);
and U8713 (N_8713,N_6403,N_6228);
or U8714 (N_8714,N_6392,N_6449);
nand U8715 (N_8715,N_6771,N_6874);
xor U8716 (N_8716,N_7283,N_6479);
nor U8717 (N_8717,N_6410,N_6682);
xor U8718 (N_8718,N_6156,N_6758);
xor U8719 (N_8719,N_7024,N_6331);
or U8720 (N_8720,N_6974,N_7436);
nor U8721 (N_8721,N_7106,N_7425);
xor U8722 (N_8722,N_7250,N_6326);
or U8723 (N_8723,N_6971,N_7379);
xor U8724 (N_8724,N_6854,N_6863);
nor U8725 (N_8725,N_7160,N_6187);
nor U8726 (N_8726,N_6549,N_7140);
or U8727 (N_8727,N_7091,N_7434);
xnor U8728 (N_8728,N_6774,N_7336);
nand U8729 (N_8729,N_6928,N_6870);
nand U8730 (N_8730,N_7218,N_6818);
xor U8731 (N_8731,N_6383,N_6903);
and U8732 (N_8732,N_6912,N_7393);
or U8733 (N_8733,N_6588,N_7168);
xnor U8734 (N_8734,N_7126,N_6934);
xnor U8735 (N_8735,N_6085,N_6434);
or U8736 (N_8736,N_6605,N_6177);
nand U8737 (N_8737,N_6696,N_6116);
nor U8738 (N_8738,N_6635,N_6650);
nand U8739 (N_8739,N_6595,N_6080);
or U8740 (N_8740,N_6864,N_6938);
nand U8741 (N_8741,N_7091,N_6604);
nand U8742 (N_8742,N_7418,N_6029);
or U8743 (N_8743,N_6045,N_6085);
nor U8744 (N_8744,N_7485,N_6727);
or U8745 (N_8745,N_6465,N_6171);
nor U8746 (N_8746,N_6431,N_7173);
and U8747 (N_8747,N_6994,N_7461);
nor U8748 (N_8748,N_6682,N_6973);
or U8749 (N_8749,N_7296,N_7322);
and U8750 (N_8750,N_6704,N_6775);
and U8751 (N_8751,N_6554,N_6861);
nor U8752 (N_8752,N_6025,N_7424);
xnor U8753 (N_8753,N_6009,N_6966);
nor U8754 (N_8754,N_7434,N_7276);
and U8755 (N_8755,N_6488,N_6335);
nor U8756 (N_8756,N_6871,N_6188);
xnor U8757 (N_8757,N_6604,N_6923);
xnor U8758 (N_8758,N_6505,N_7465);
or U8759 (N_8759,N_6275,N_6042);
nand U8760 (N_8760,N_7341,N_6048);
nor U8761 (N_8761,N_7377,N_7090);
xor U8762 (N_8762,N_6263,N_6683);
and U8763 (N_8763,N_6152,N_7083);
nand U8764 (N_8764,N_6175,N_7100);
or U8765 (N_8765,N_6777,N_7038);
nand U8766 (N_8766,N_6955,N_6827);
xnor U8767 (N_8767,N_7424,N_6221);
nand U8768 (N_8768,N_6495,N_7175);
nand U8769 (N_8769,N_6405,N_6468);
nor U8770 (N_8770,N_6487,N_6341);
nor U8771 (N_8771,N_6575,N_6202);
nor U8772 (N_8772,N_6765,N_6359);
xor U8773 (N_8773,N_6528,N_7129);
xor U8774 (N_8774,N_6599,N_7256);
nor U8775 (N_8775,N_6426,N_6533);
nor U8776 (N_8776,N_7380,N_6839);
and U8777 (N_8777,N_6613,N_6406);
xor U8778 (N_8778,N_6580,N_7331);
or U8779 (N_8779,N_7180,N_7202);
nand U8780 (N_8780,N_7151,N_6913);
or U8781 (N_8781,N_6683,N_6977);
and U8782 (N_8782,N_6088,N_7088);
nor U8783 (N_8783,N_6445,N_6154);
nand U8784 (N_8784,N_7175,N_7390);
xnor U8785 (N_8785,N_6723,N_7466);
xor U8786 (N_8786,N_6616,N_7372);
or U8787 (N_8787,N_7470,N_7306);
xor U8788 (N_8788,N_6064,N_6038);
nand U8789 (N_8789,N_7493,N_6345);
and U8790 (N_8790,N_6117,N_6712);
nand U8791 (N_8791,N_7245,N_7423);
or U8792 (N_8792,N_6699,N_6535);
and U8793 (N_8793,N_6487,N_6926);
and U8794 (N_8794,N_7366,N_6746);
nor U8795 (N_8795,N_7271,N_6247);
or U8796 (N_8796,N_6363,N_7221);
xnor U8797 (N_8797,N_6921,N_7432);
and U8798 (N_8798,N_6353,N_7205);
nand U8799 (N_8799,N_6441,N_7406);
xnor U8800 (N_8800,N_6631,N_6045);
or U8801 (N_8801,N_7403,N_6174);
and U8802 (N_8802,N_6479,N_6229);
and U8803 (N_8803,N_7237,N_7231);
nor U8804 (N_8804,N_7330,N_6524);
nand U8805 (N_8805,N_6391,N_6885);
nand U8806 (N_8806,N_6630,N_6680);
or U8807 (N_8807,N_7121,N_6058);
xnor U8808 (N_8808,N_6857,N_6234);
nor U8809 (N_8809,N_6655,N_7183);
or U8810 (N_8810,N_6670,N_6065);
and U8811 (N_8811,N_6388,N_7021);
or U8812 (N_8812,N_7370,N_7037);
or U8813 (N_8813,N_6380,N_6187);
xor U8814 (N_8814,N_6738,N_6025);
xor U8815 (N_8815,N_6651,N_6491);
nand U8816 (N_8816,N_6268,N_6806);
or U8817 (N_8817,N_6171,N_6654);
nor U8818 (N_8818,N_6008,N_6890);
xor U8819 (N_8819,N_6076,N_6983);
xnor U8820 (N_8820,N_6078,N_7135);
nand U8821 (N_8821,N_6418,N_7163);
nand U8822 (N_8822,N_7164,N_6415);
or U8823 (N_8823,N_6586,N_7116);
and U8824 (N_8824,N_6905,N_6395);
or U8825 (N_8825,N_7185,N_7329);
nand U8826 (N_8826,N_6318,N_6224);
nor U8827 (N_8827,N_7187,N_6325);
nand U8828 (N_8828,N_6218,N_7141);
and U8829 (N_8829,N_6397,N_7407);
nand U8830 (N_8830,N_6297,N_6419);
xnor U8831 (N_8831,N_6527,N_6932);
nor U8832 (N_8832,N_6220,N_6464);
xor U8833 (N_8833,N_6875,N_6280);
and U8834 (N_8834,N_6403,N_7242);
xnor U8835 (N_8835,N_6076,N_6335);
nor U8836 (N_8836,N_7149,N_7322);
nand U8837 (N_8837,N_7493,N_6711);
or U8838 (N_8838,N_6335,N_6966);
and U8839 (N_8839,N_7206,N_6629);
and U8840 (N_8840,N_6103,N_6858);
and U8841 (N_8841,N_7202,N_6646);
nand U8842 (N_8842,N_6945,N_6972);
and U8843 (N_8843,N_6655,N_7262);
nor U8844 (N_8844,N_7127,N_7223);
nand U8845 (N_8845,N_6509,N_6120);
nand U8846 (N_8846,N_6344,N_7365);
nor U8847 (N_8847,N_6713,N_6903);
and U8848 (N_8848,N_6318,N_7410);
or U8849 (N_8849,N_7248,N_6158);
nor U8850 (N_8850,N_7470,N_7368);
xnor U8851 (N_8851,N_7489,N_6559);
nor U8852 (N_8852,N_6904,N_6908);
nor U8853 (N_8853,N_6922,N_6963);
or U8854 (N_8854,N_6810,N_6652);
or U8855 (N_8855,N_7010,N_6628);
or U8856 (N_8856,N_6060,N_6601);
nand U8857 (N_8857,N_6726,N_6924);
and U8858 (N_8858,N_7436,N_6753);
xnor U8859 (N_8859,N_6370,N_6810);
nand U8860 (N_8860,N_6112,N_7170);
xnor U8861 (N_8861,N_6234,N_7131);
nand U8862 (N_8862,N_6908,N_7353);
nor U8863 (N_8863,N_6725,N_7376);
or U8864 (N_8864,N_7403,N_7101);
and U8865 (N_8865,N_7319,N_7007);
nand U8866 (N_8866,N_6461,N_7061);
and U8867 (N_8867,N_6155,N_6374);
or U8868 (N_8868,N_6848,N_7448);
nor U8869 (N_8869,N_6780,N_6601);
and U8870 (N_8870,N_7423,N_7047);
xor U8871 (N_8871,N_6274,N_6683);
xnor U8872 (N_8872,N_7441,N_7457);
nand U8873 (N_8873,N_7222,N_7368);
or U8874 (N_8874,N_6120,N_7489);
nor U8875 (N_8875,N_6236,N_7384);
or U8876 (N_8876,N_6676,N_6571);
nor U8877 (N_8877,N_6678,N_6104);
nand U8878 (N_8878,N_7250,N_7114);
nand U8879 (N_8879,N_6463,N_7223);
xor U8880 (N_8880,N_6087,N_7355);
nor U8881 (N_8881,N_6201,N_6343);
and U8882 (N_8882,N_6574,N_7486);
and U8883 (N_8883,N_6025,N_7281);
or U8884 (N_8884,N_6658,N_6120);
or U8885 (N_8885,N_6642,N_6208);
and U8886 (N_8886,N_6583,N_6333);
xnor U8887 (N_8887,N_7350,N_6815);
or U8888 (N_8888,N_7042,N_6669);
nor U8889 (N_8889,N_6658,N_6557);
xor U8890 (N_8890,N_6015,N_7424);
xnor U8891 (N_8891,N_7008,N_6654);
nor U8892 (N_8892,N_7266,N_6196);
nand U8893 (N_8893,N_6913,N_6697);
xor U8894 (N_8894,N_7372,N_6617);
nand U8895 (N_8895,N_7494,N_6293);
xnor U8896 (N_8896,N_6543,N_6638);
nor U8897 (N_8897,N_6122,N_7488);
or U8898 (N_8898,N_7212,N_7117);
nand U8899 (N_8899,N_6303,N_6873);
and U8900 (N_8900,N_7154,N_6370);
or U8901 (N_8901,N_6555,N_6097);
nor U8902 (N_8902,N_6810,N_7346);
or U8903 (N_8903,N_6762,N_7345);
nand U8904 (N_8904,N_7469,N_6640);
or U8905 (N_8905,N_6656,N_7246);
nand U8906 (N_8906,N_6965,N_7332);
nor U8907 (N_8907,N_6194,N_6735);
nand U8908 (N_8908,N_6662,N_7244);
nor U8909 (N_8909,N_6231,N_6907);
nor U8910 (N_8910,N_6863,N_6855);
or U8911 (N_8911,N_7290,N_7205);
nor U8912 (N_8912,N_6618,N_6261);
and U8913 (N_8913,N_7231,N_7315);
or U8914 (N_8914,N_6251,N_6440);
and U8915 (N_8915,N_6639,N_7161);
or U8916 (N_8916,N_6182,N_6059);
and U8917 (N_8917,N_7247,N_6541);
xor U8918 (N_8918,N_7280,N_7459);
xor U8919 (N_8919,N_7267,N_6836);
nor U8920 (N_8920,N_6378,N_6258);
and U8921 (N_8921,N_6532,N_7248);
and U8922 (N_8922,N_6193,N_6264);
nand U8923 (N_8923,N_6324,N_7323);
nor U8924 (N_8924,N_7337,N_6621);
nor U8925 (N_8925,N_6862,N_6878);
or U8926 (N_8926,N_6194,N_6789);
xnor U8927 (N_8927,N_7212,N_6823);
nor U8928 (N_8928,N_6528,N_6700);
nand U8929 (N_8929,N_6811,N_6067);
nor U8930 (N_8930,N_6984,N_6183);
nand U8931 (N_8931,N_6203,N_6969);
nor U8932 (N_8932,N_6747,N_6621);
xnor U8933 (N_8933,N_6366,N_6109);
or U8934 (N_8934,N_6931,N_6816);
nor U8935 (N_8935,N_6571,N_6288);
nor U8936 (N_8936,N_6233,N_6283);
nand U8937 (N_8937,N_7496,N_7460);
nand U8938 (N_8938,N_6903,N_6666);
xnor U8939 (N_8939,N_6760,N_7354);
xnor U8940 (N_8940,N_6896,N_6472);
nor U8941 (N_8941,N_6108,N_7315);
and U8942 (N_8942,N_7132,N_6294);
or U8943 (N_8943,N_7119,N_6595);
xnor U8944 (N_8944,N_7244,N_6060);
nor U8945 (N_8945,N_6699,N_6236);
and U8946 (N_8946,N_6069,N_6902);
and U8947 (N_8947,N_7150,N_6592);
xnor U8948 (N_8948,N_6941,N_6139);
nor U8949 (N_8949,N_6027,N_7417);
xnor U8950 (N_8950,N_6858,N_7116);
and U8951 (N_8951,N_6071,N_7446);
xor U8952 (N_8952,N_7134,N_6903);
nand U8953 (N_8953,N_7077,N_7283);
xor U8954 (N_8954,N_6448,N_7308);
and U8955 (N_8955,N_6425,N_6190);
nand U8956 (N_8956,N_7017,N_7160);
nand U8957 (N_8957,N_6750,N_6117);
and U8958 (N_8958,N_7341,N_6869);
nand U8959 (N_8959,N_7027,N_6430);
nand U8960 (N_8960,N_6819,N_7320);
and U8961 (N_8961,N_6765,N_6328);
nor U8962 (N_8962,N_7462,N_7386);
and U8963 (N_8963,N_7477,N_6707);
or U8964 (N_8964,N_6286,N_6084);
and U8965 (N_8965,N_6783,N_6465);
xor U8966 (N_8966,N_6323,N_6977);
nand U8967 (N_8967,N_6440,N_7045);
nor U8968 (N_8968,N_7060,N_7175);
nor U8969 (N_8969,N_6664,N_6247);
and U8970 (N_8970,N_6350,N_6260);
and U8971 (N_8971,N_6186,N_6423);
or U8972 (N_8972,N_7469,N_7252);
or U8973 (N_8973,N_6394,N_6104);
and U8974 (N_8974,N_7121,N_7311);
xnor U8975 (N_8975,N_6345,N_6776);
nand U8976 (N_8976,N_6445,N_7014);
nor U8977 (N_8977,N_6313,N_7362);
nand U8978 (N_8978,N_6842,N_6295);
nand U8979 (N_8979,N_6268,N_6150);
xnor U8980 (N_8980,N_6190,N_7139);
or U8981 (N_8981,N_6434,N_6729);
and U8982 (N_8982,N_7454,N_6185);
or U8983 (N_8983,N_6518,N_7047);
or U8984 (N_8984,N_7204,N_6464);
and U8985 (N_8985,N_6757,N_7229);
xor U8986 (N_8986,N_6474,N_7247);
xnor U8987 (N_8987,N_6560,N_7209);
nor U8988 (N_8988,N_6187,N_7234);
nand U8989 (N_8989,N_6011,N_6254);
xor U8990 (N_8990,N_6127,N_7111);
or U8991 (N_8991,N_6082,N_6206);
xnor U8992 (N_8992,N_6830,N_7075);
and U8993 (N_8993,N_7288,N_7360);
nor U8994 (N_8994,N_6259,N_6989);
or U8995 (N_8995,N_6734,N_6616);
and U8996 (N_8996,N_7434,N_6630);
xor U8997 (N_8997,N_7280,N_6803);
xor U8998 (N_8998,N_7337,N_6680);
nand U8999 (N_8999,N_6379,N_7105);
nor U9000 (N_9000,N_8008,N_8254);
and U9001 (N_9001,N_8895,N_8321);
and U9002 (N_9002,N_8700,N_8104);
or U9003 (N_9003,N_7608,N_8566);
nor U9004 (N_9004,N_8387,N_8375);
or U9005 (N_9005,N_7660,N_7600);
or U9006 (N_9006,N_7612,N_8453);
nand U9007 (N_9007,N_8891,N_8064);
xor U9008 (N_9008,N_8850,N_7718);
nand U9009 (N_9009,N_8780,N_8890);
or U9010 (N_9010,N_8662,N_7709);
or U9011 (N_9011,N_8930,N_7858);
or U9012 (N_9012,N_8364,N_8155);
nor U9013 (N_9013,N_8531,N_8690);
and U9014 (N_9014,N_8560,N_8846);
and U9015 (N_9015,N_7655,N_8436);
and U9016 (N_9016,N_8685,N_7755);
nor U9017 (N_9017,N_8402,N_8195);
nor U9018 (N_9018,N_7673,N_8392);
nor U9019 (N_9019,N_8694,N_8371);
and U9020 (N_9020,N_7842,N_7951);
nand U9021 (N_9021,N_7888,N_7806);
xor U9022 (N_9022,N_8206,N_8153);
nand U9023 (N_9023,N_7958,N_8989);
and U9024 (N_9024,N_8672,N_8490);
nor U9025 (N_9025,N_8553,N_8742);
or U9026 (N_9026,N_8857,N_7791);
xor U9027 (N_9027,N_8051,N_8606);
or U9028 (N_9028,N_8154,N_8594);
and U9029 (N_9029,N_8474,N_7552);
and U9030 (N_9030,N_7939,N_7730);
xnor U9031 (N_9031,N_8649,N_8109);
and U9032 (N_9032,N_8860,N_8084);
or U9033 (N_9033,N_7564,N_8894);
nor U9034 (N_9034,N_8726,N_8188);
xnor U9035 (N_9035,N_8950,N_8975);
or U9036 (N_9036,N_8452,N_8707);
xor U9037 (N_9037,N_8691,N_8476);
nand U9038 (N_9038,N_8212,N_8279);
nor U9039 (N_9039,N_7707,N_7578);
or U9040 (N_9040,N_8388,N_8249);
and U9041 (N_9041,N_8351,N_7532);
nor U9042 (N_9042,N_8259,N_8596);
or U9043 (N_9043,N_8514,N_8335);
or U9044 (N_9044,N_7903,N_8302);
nor U9045 (N_9045,N_8903,N_8372);
and U9046 (N_9046,N_8945,N_8246);
or U9047 (N_9047,N_8763,N_8512);
or U9048 (N_9048,N_8067,N_7774);
and U9049 (N_9049,N_8611,N_8519);
or U9050 (N_9050,N_8783,N_7577);
nor U9051 (N_9051,N_8532,N_8097);
and U9052 (N_9052,N_7554,N_8066);
or U9053 (N_9053,N_8712,N_7638);
or U9054 (N_9054,N_7807,N_7705);
nand U9055 (N_9055,N_8654,N_8463);
or U9056 (N_9056,N_8171,N_8396);
and U9057 (N_9057,N_7770,N_8468);
and U9058 (N_9058,N_8577,N_8541);
nand U9059 (N_9059,N_8352,N_8883);
nand U9060 (N_9060,N_7688,N_7698);
nor U9061 (N_9061,N_7780,N_8982);
or U9062 (N_9062,N_8092,N_8026);
and U9063 (N_9063,N_7777,N_7559);
xnor U9064 (N_9064,N_7759,N_8717);
or U9065 (N_9065,N_8162,N_8681);
nand U9066 (N_9066,N_8904,N_8622);
nor U9067 (N_9067,N_8349,N_8709);
nand U9068 (N_9068,N_8211,N_8922);
and U9069 (N_9069,N_8605,N_7764);
nor U9070 (N_9070,N_8477,N_7535);
and U9071 (N_9071,N_7902,N_8487);
xnor U9072 (N_9072,N_8919,N_8770);
and U9073 (N_9073,N_7666,N_7592);
xor U9074 (N_9074,N_8976,N_7675);
or U9075 (N_9075,N_8174,N_7756);
nand U9076 (N_9076,N_7889,N_8803);
and U9077 (N_9077,N_8409,N_7972);
or U9078 (N_9078,N_7845,N_8258);
xor U9079 (N_9079,N_8161,N_7974);
xnor U9080 (N_9080,N_7636,N_8908);
or U9081 (N_9081,N_8808,N_8497);
or U9082 (N_9082,N_8973,N_7996);
nand U9083 (N_9083,N_8809,N_7987);
and U9084 (N_9084,N_8695,N_7907);
and U9085 (N_9085,N_8141,N_8076);
nor U9086 (N_9086,N_7886,N_7722);
xnor U9087 (N_9087,N_8927,N_7773);
or U9088 (N_9088,N_7904,N_8277);
nor U9089 (N_9089,N_7905,N_8173);
xnor U9090 (N_9090,N_8933,N_8494);
xnor U9091 (N_9091,N_8237,N_8117);
or U9092 (N_9092,N_8492,N_8444);
and U9093 (N_9093,N_8844,N_8993);
and U9094 (N_9094,N_7884,N_7613);
nand U9095 (N_9095,N_8004,N_7644);
nand U9096 (N_9096,N_8417,N_8175);
xor U9097 (N_9097,N_8988,N_8003);
nand U9098 (N_9098,N_8242,N_7841);
nand U9099 (N_9099,N_8429,N_8106);
and U9100 (N_9100,N_8885,N_7736);
nand U9101 (N_9101,N_8193,N_8901);
nand U9102 (N_9102,N_8370,N_8458);
xnor U9103 (N_9103,N_8227,N_7910);
nor U9104 (N_9104,N_7717,N_8344);
xor U9105 (N_9105,N_7859,N_8774);
nand U9106 (N_9106,N_8621,N_8610);
and U9107 (N_9107,N_8460,N_7606);
and U9108 (N_9108,N_8368,N_8985);
nand U9109 (N_9109,N_7874,N_8493);
nand U9110 (N_9110,N_8957,N_8061);
or U9111 (N_9111,N_8473,N_8217);
nor U9112 (N_9112,N_8183,N_7618);
nand U9113 (N_9113,N_7751,N_8794);
nor U9114 (N_9114,N_8591,N_8399);
or U9115 (N_9115,N_8646,N_7594);
nor U9116 (N_9116,N_8992,N_8854);
or U9117 (N_9117,N_8401,N_8853);
or U9118 (N_9118,N_7508,N_8159);
xor U9119 (N_9119,N_8562,N_8397);
nor U9120 (N_9120,N_8789,N_8385);
xor U9121 (N_9121,N_7720,N_8521);
nand U9122 (N_9122,N_8245,N_7801);
xor U9123 (N_9123,N_8574,N_8791);
or U9124 (N_9124,N_8953,N_8815);
and U9125 (N_9125,N_7950,N_8380);
and U9126 (N_9126,N_7686,N_8379);
and U9127 (N_9127,N_7980,N_8085);
nor U9128 (N_9128,N_7569,N_8482);
nor U9129 (N_9129,N_7669,N_8329);
nor U9130 (N_9130,N_8164,N_8609);
or U9131 (N_9131,N_8810,N_8111);
or U9132 (N_9132,N_8229,N_7781);
xnor U9133 (N_9133,N_8485,N_8342);
nor U9134 (N_9134,N_8811,N_7741);
xnor U9135 (N_9135,N_8907,N_8038);
xnor U9136 (N_9136,N_8569,N_7820);
and U9137 (N_9137,N_7985,N_7919);
or U9138 (N_9138,N_8830,N_8859);
nand U9139 (N_9139,N_8074,N_8313);
or U9140 (N_9140,N_8251,N_8872);
xnor U9141 (N_9141,N_8079,N_8875);
or U9142 (N_9142,N_8197,N_8006);
xor U9143 (N_9143,N_8619,N_8420);
and U9144 (N_9144,N_8090,N_8708);
xor U9145 (N_9145,N_8101,N_8886);
nand U9146 (N_9146,N_7533,N_8880);
nor U9147 (N_9147,N_8938,N_8644);
xnor U9148 (N_9148,N_8210,N_7584);
and U9149 (N_9149,N_8878,N_7761);
nand U9150 (N_9150,N_8977,N_7656);
nand U9151 (N_9151,N_7649,N_7639);
xor U9152 (N_9152,N_7567,N_7783);
and U9153 (N_9153,N_8906,N_7527);
nand U9154 (N_9154,N_8226,N_8963);
nand U9155 (N_9155,N_8561,N_8847);
or U9156 (N_9156,N_8608,N_8295);
or U9157 (N_9157,N_8884,N_8925);
xnor U9158 (N_9158,N_7670,N_7968);
nor U9159 (N_9159,N_7786,N_7788);
nor U9160 (N_9160,N_8817,N_7620);
or U9161 (N_9161,N_8876,N_8589);
or U9162 (N_9162,N_8959,N_7802);
xor U9163 (N_9163,N_7511,N_7732);
or U9164 (N_9164,N_7938,N_7557);
and U9165 (N_9165,N_7500,N_8551);
xor U9166 (N_9166,N_8348,N_8733);
xor U9167 (N_9167,N_8432,N_8149);
nand U9168 (N_9168,N_7719,N_7760);
and U9169 (N_9169,N_7978,N_7714);
xor U9170 (N_9170,N_8238,N_7685);
and U9171 (N_9171,N_8518,N_7819);
and U9172 (N_9172,N_7862,N_8807);
nand U9173 (N_9173,N_8509,N_7892);
nand U9174 (N_9174,N_8291,N_7937);
nor U9175 (N_9175,N_7662,N_8782);
or U9176 (N_9176,N_8506,N_8105);
and U9177 (N_9177,N_8784,N_8792);
nor U9178 (N_9178,N_7723,N_7521);
nor U9179 (N_9179,N_8099,N_8033);
or U9180 (N_9180,N_8586,N_8639);
nand U9181 (N_9181,N_8260,N_8102);
xor U9182 (N_9182,N_8871,N_8032);
and U9183 (N_9183,N_7823,N_8734);
and U9184 (N_9184,N_8446,N_8350);
nand U9185 (N_9185,N_7843,N_8096);
nand U9186 (N_9186,N_7932,N_7598);
xnor U9187 (N_9187,N_7616,N_8664);
xor U9188 (N_9188,N_8526,N_8472);
nor U9189 (N_9189,N_8471,N_7810);
nand U9190 (N_9190,N_7915,N_7945);
or U9191 (N_9191,N_8016,N_8762);
or U9192 (N_9192,N_7556,N_8430);
or U9193 (N_9193,N_8145,N_8597);
nand U9194 (N_9194,N_8421,N_8580);
or U9195 (N_9195,N_8146,N_7692);
or U9196 (N_9196,N_8314,N_8336);
and U9197 (N_9197,N_8592,N_7876);
nor U9198 (N_9198,N_8383,N_8386);
nor U9199 (N_9199,N_8640,N_8579);
nor U9200 (N_9200,N_8994,N_8682);
xor U9201 (N_9201,N_8643,N_8999);
nor U9202 (N_9202,N_8942,N_8200);
nor U9203 (N_9203,N_8823,N_7796);
or U9204 (N_9204,N_7540,N_8523);
or U9205 (N_9205,N_8947,N_8582);
nand U9206 (N_9206,N_7778,N_8650);
or U9207 (N_9207,N_7966,N_8330);
nand U9208 (N_9208,N_8507,N_8852);
and U9209 (N_9209,N_8118,N_7955);
or U9210 (N_9210,N_8554,N_8483);
or U9211 (N_9211,N_7581,N_7812);
nor U9212 (N_9212,N_8669,N_8819);
nor U9213 (N_9213,N_8900,N_7952);
or U9214 (N_9214,N_8499,N_8180);
nand U9215 (N_9215,N_8310,N_7826);
or U9216 (N_9216,N_7645,N_7558);
and U9217 (N_9217,N_8040,N_8393);
xor U9218 (N_9218,N_7696,N_8728);
nor U9219 (N_9219,N_8635,N_7502);
or U9220 (N_9220,N_8533,N_7962);
nor U9221 (N_9221,N_7525,N_7694);
and U9222 (N_9222,N_8576,N_8137);
nand U9223 (N_9223,N_7961,N_8305);
nor U9224 (N_9224,N_7630,N_8858);
nor U9225 (N_9225,N_7896,N_8593);
or U9226 (N_9226,N_8658,N_7973);
nor U9227 (N_9227,N_8839,N_8012);
xor U9228 (N_9228,N_7779,N_8501);
and U9229 (N_9229,N_7772,N_8581);
nor U9230 (N_9230,N_8100,N_8108);
nor U9231 (N_9231,N_7844,N_7857);
nor U9232 (N_9232,N_7993,N_8767);
xnor U9233 (N_9233,N_8094,N_7665);
and U9234 (N_9234,N_7839,N_8828);
nand U9235 (N_9235,N_8115,N_7603);
or U9236 (N_9236,N_8165,N_8382);
xor U9237 (N_9237,N_8422,N_8618);
and U9238 (N_9238,N_7880,N_7870);
and U9239 (N_9239,N_8738,N_8949);
nand U9240 (N_9240,N_7815,N_8272);
xor U9241 (N_9241,N_8796,N_8062);
xor U9242 (N_9242,N_7659,N_8710);
nand U9243 (N_9243,N_8740,N_8882);
nand U9244 (N_9244,N_8496,N_8152);
or U9245 (N_9245,N_7800,N_7681);
or U9246 (N_9246,N_8470,N_8128);
nor U9247 (N_9247,N_8338,N_8355);
nor U9248 (N_9248,N_7731,N_8340);
or U9249 (N_9249,N_7632,N_8913);
and U9250 (N_9250,N_8737,N_8928);
nor U9251 (N_9251,N_8918,N_8686);
or U9252 (N_9252,N_8825,N_7625);
or U9253 (N_9253,N_8256,N_8018);
xnor U9254 (N_9254,N_8081,N_8046);
and U9255 (N_9255,N_7652,N_8187);
nor U9256 (N_9256,N_8119,N_8292);
and U9257 (N_9257,N_7671,N_8513);
nand U9258 (N_9258,N_8788,N_8083);
or U9259 (N_9259,N_8931,N_8011);
or U9260 (N_9260,N_8600,N_8970);
nand U9261 (N_9261,N_7804,N_8007);
nand U9262 (N_9262,N_8902,N_8270);
nor U9263 (N_9263,N_8144,N_7833);
nor U9264 (N_9264,N_8264,N_8239);
nor U9265 (N_9265,N_8620,N_8833);
xnor U9266 (N_9266,N_8773,N_8013);
or U9267 (N_9267,N_7953,N_7550);
xor U9268 (N_9268,N_8280,N_7522);
nor U9269 (N_9269,N_7768,N_7941);
and U9270 (N_9270,N_8181,N_8874);
xor U9271 (N_9271,N_8546,N_8879);
and U9272 (N_9272,N_8941,N_8345);
nand U9273 (N_9273,N_7501,N_8747);
xnor U9274 (N_9274,N_8914,N_8315);
xnor U9275 (N_9275,N_8148,N_7745);
xor U9276 (N_9276,N_8966,N_8268);
or U9277 (N_9277,N_7629,N_8278);
nor U9278 (N_9278,N_8486,N_8751);
nand U9279 (N_9279,N_8732,N_8556);
nand U9280 (N_9280,N_8539,N_7586);
xnor U9281 (N_9281,N_8398,N_7658);
or U9282 (N_9282,N_8326,N_8086);
or U9283 (N_9283,N_7512,N_8881);
nor U9284 (N_9284,N_8920,N_8758);
nand U9285 (N_9285,N_8641,N_7514);
or U9286 (N_9286,N_7726,N_7633);
xnor U9287 (N_9287,N_8534,N_8631);
xnor U9288 (N_9288,N_7808,N_8893);
or U9289 (N_9289,N_7861,N_8912);
nand U9290 (N_9290,N_8516,N_8015);
nand U9291 (N_9291,N_7589,N_8439);
nor U9292 (N_9292,N_8124,N_8199);
xnor U9293 (N_9293,N_8303,N_8495);
xor U9294 (N_9294,N_8220,N_8921);
xnor U9295 (N_9295,N_7548,N_8410);
and U9296 (N_9296,N_8836,N_7505);
xor U9297 (N_9297,N_7828,N_8755);
xnor U9298 (N_9298,N_8029,N_7999);
and U9299 (N_9299,N_8070,N_8729);
nand U9300 (N_9300,N_8065,N_7553);
nor U9301 (N_9301,N_8971,N_7882);
nand U9302 (N_9302,N_7534,N_8870);
xor U9303 (N_9303,N_8163,N_7684);
nor U9304 (N_9304,N_7537,N_7699);
or U9305 (N_9305,N_7555,N_7715);
nand U9306 (N_9306,N_8845,N_8300);
nand U9307 (N_9307,N_7957,N_7596);
xor U9308 (N_9308,N_8050,N_8488);
nor U9309 (N_9309,N_7798,N_8716);
and U9310 (N_9310,N_7852,N_8223);
and U9311 (N_9311,N_8481,N_8025);
and U9312 (N_9312,N_8759,N_8140);
nand U9313 (N_9313,N_8588,N_7942);
and U9314 (N_9314,N_8282,N_8002);
nor U9315 (N_9315,N_7960,N_8243);
or U9316 (N_9316,N_8688,N_7713);
nor U9317 (N_9317,N_8323,N_8670);
xnor U9318 (N_9318,N_8696,N_7887);
nor U9319 (N_9319,N_7847,N_8415);
or U9320 (N_9320,N_8575,N_7947);
nor U9321 (N_9321,N_7542,N_8892);
or U9322 (N_9322,N_8034,N_8739);
nand U9323 (N_9323,N_7994,N_7562);
nand U9324 (N_9324,N_8826,N_8353);
nor U9325 (N_9325,N_7752,N_7591);
nor U9326 (N_9326,N_7797,N_7579);
and U9327 (N_9327,N_8271,N_8676);
and U9328 (N_9328,N_8139,N_8343);
or U9329 (N_9329,N_7610,N_7517);
and U9330 (N_9330,N_7899,N_8311);
nand U9331 (N_9331,N_8714,N_8552);
nor U9332 (N_9332,N_7921,N_8044);
nor U9333 (N_9333,N_8435,N_7516);
xor U9334 (N_9334,N_7728,N_8235);
xnor U9335 (N_9335,N_8967,N_8812);
xor U9336 (N_9336,N_7513,N_7927);
xnor U9337 (N_9337,N_7680,N_8629);
and U9338 (N_9338,N_8517,N_7565);
nand U9339 (N_9339,N_8771,N_7871);
nand U9340 (N_9340,N_7765,N_7716);
nor U9341 (N_9341,N_8186,N_8088);
xor U9342 (N_9342,N_8655,N_8135);
nand U9343 (N_9343,N_8457,N_8121);
or U9344 (N_9344,N_7744,N_7689);
nand U9345 (N_9345,N_8730,N_8306);
nor U9346 (N_9346,N_7943,N_8851);
xor U9347 (N_9347,N_7867,N_7964);
xor U9348 (N_9348,N_8565,N_8752);
or U9349 (N_9349,N_8215,N_7747);
nor U9350 (N_9350,N_8766,N_8363);
nor U9351 (N_9351,N_8684,N_8865);
nand U9352 (N_9352,N_8142,N_7771);
nor U9353 (N_9353,N_8308,N_7743);
nor U9354 (N_9354,N_7856,N_8428);
and U9355 (N_9355,N_8598,N_8424);
or U9356 (N_9356,N_8722,N_8120);
and U9357 (N_9357,N_8339,N_7831);
nor U9358 (N_9358,N_7753,N_8951);
or U9359 (N_9359,N_7614,N_8940);
nand U9360 (N_9360,N_8361,N_7840);
and U9361 (N_9361,N_8133,N_8761);
nand U9362 (N_9362,N_8182,N_8804);
nor U9363 (N_9363,N_8341,N_8797);
nand U9364 (N_9364,N_8433,N_8301);
nand U9365 (N_9365,N_8047,N_8652);
and U9366 (N_9366,N_7750,N_8151);
xor U9367 (N_9367,N_7979,N_7519);
and U9368 (N_9368,N_8749,N_7930);
or U9369 (N_9369,N_8653,N_8800);
xnor U9370 (N_9370,N_7640,N_8571);
nor U9371 (N_9371,N_8451,N_7809);
nor U9372 (N_9372,N_8802,N_8122);
nor U9373 (N_9373,N_7650,N_8281);
nand U9374 (N_9374,N_8793,N_8461);
xnor U9375 (N_9375,N_7678,N_8630);
nor U9376 (N_9376,N_7827,N_8524);
or U9377 (N_9377,N_8412,N_8805);
or U9378 (N_9378,N_8334,N_8990);
xor U9379 (N_9379,N_8502,N_8926);
nor U9380 (N_9380,N_7997,N_7885);
nor U9381 (N_9381,N_8287,N_8359);
and U9382 (N_9382,N_7568,N_8743);
nor U9383 (N_9383,N_8244,N_8276);
xnor U9384 (N_9384,N_8842,N_8358);
xor U9385 (N_9385,N_7635,N_7883);
nand U9386 (N_9386,N_8373,N_7536);
and U9387 (N_9387,N_7695,N_8750);
and U9388 (N_9388,N_8855,N_8668);
xor U9389 (N_9389,N_7721,N_7700);
nor U9390 (N_9390,N_7712,N_8078);
nand U9391 (N_9391,N_8489,N_8357);
and U9392 (N_9392,N_8583,N_7661);
xor U9393 (N_9393,N_8877,N_8418);
xor U9394 (N_9394,N_8657,N_8331);
xor U9395 (N_9395,N_8039,N_8748);
nor U9396 (N_9396,N_8285,N_8776);
xor U9397 (N_9397,N_8756,N_7991);
xor U9398 (N_9398,N_8168,N_8602);
or U9399 (N_9399,N_7834,N_8009);
nor U9400 (N_9400,N_8515,N_7623);
nor U9401 (N_9401,N_8498,N_8230);
xor U9402 (N_9402,N_7646,N_7893);
xnor U9403 (N_9403,N_8150,N_7956);
nand U9404 (N_9404,N_8547,N_8980);
or U9405 (N_9405,N_8544,N_8005);
and U9406 (N_9406,N_7869,N_8127);
xor U9407 (N_9407,N_7787,N_8968);
xnor U9408 (N_9408,N_8563,N_8134);
nand U9409 (N_9409,N_7916,N_7836);
xnor U9410 (N_9410,N_8692,N_8715);
or U9411 (N_9411,N_8296,N_7529);
or U9412 (N_9412,N_8827,N_7729);
nor U9413 (N_9413,N_8365,N_7622);
nand U9414 (N_9414,N_7822,N_8068);
or U9415 (N_9415,N_8824,N_7549);
xnor U9416 (N_9416,N_8558,N_8645);
nor U9417 (N_9417,N_8138,N_8572);
nand U9418 (N_9418,N_8202,N_7894);
or U9419 (N_9419,N_7693,N_8636);
xnor U9420 (N_9420,N_7895,N_7510);
and U9421 (N_9421,N_8991,N_8637);
or U9422 (N_9422,N_8112,N_8427);
xor U9423 (N_9423,N_7878,N_7507);
and U9424 (N_9424,N_8022,N_8896);
and U9425 (N_9425,N_8663,N_8503);
or U9426 (N_9426,N_8219,N_7805);
nand U9427 (N_9427,N_7898,N_7573);
and U9428 (N_9428,N_7775,N_7992);
and U9429 (N_9429,N_8316,N_8969);
and U9430 (N_9430,N_7544,N_7627);
and U9431 (N_9431,N_7965,N_8848);
xnor U9432 (N_9432,N_8248,N_8213);
or U9433 (N_9433,N_7615,N_8772);
xor U9434 (N_9434,N_8275,N_8981);
nand U9435 (N_9435,N_7983,N_8419);
or U9436 (N_9436,N_7710,N_7737);
or U9437 (N_9437,N_8866,N_8167);
and U9438 (N_9438,N_7855,N_7526);
and U9439 (N_9439,N_7793,N_8376);
and U9440 (N_9440,N_8098,N_8616);
nor U9441 (N_9441,N_8987,N_7879);
and U9442 (N_9442,N_8965,N_8613);
or U9443 (N_9443,N_8262,N_7624);
or U9444 (N_9444,N_7881,N_7748);
nor U9445 (N_9445,N_8216,N_7643);
and U9446 (N_9446,N_8045,N_7817);
nor U9447 (N_9447,N_8191,N_8964);
nor U9448 (N_9448,N_7776,N_8072);
nor U9449 (N_9449,N_7541,N_8687);
and U9450 (N_9450,N_8675,N_7648);
nor U9451 (N_9451,N_7725,N_7971);
nor U9452 (N_9452,N_7724,N_7604);
nor U9453 (N_9453,N_8464,N_8110);
and U9454 (N_9454,N_8059,N_7663);
nor U9455 (N_9455,N_8190,N_7865);
and U9456 (N_9456,N_8887,N_7763);
nand U9457 (N_9457,N_7563,N_7890);
nor U9458 (N_9458,N_8944,N_8208);
xor U9459 (N_9459,N_8378,N_8704);
or U9460 (N_9460,N_8573,N_8864);
nor U9461 (N_9461,N_8821,N_8103);
nand U9462 (N_9462,N_7866,N_7990);
and U9463 (N_9463,N_8440,N_7677);
and U9464 (N_9464,N_7850,N_8448);
and U9465 (N_9465,N_8325,N_7676);
nor U9466 (N_9466,N_8147,N_7547);
and U9467 (N_9467,N_8441,N_8389);
xnor U9468 (N_9468,N_8234,N_8873);
and U9469 (N_9469,N_8036,N_8627);
xor U9470 (N_9470,N_7926,N_8327);
xor U9471 (N_9471,N_8377,N_8910);
nor U9472 (N_9472,N_8028,N_8404);
or U9473 (N_9473,N_7998,N_7935);
or U9474 (N_9474,N_8995,N_8423);
nor U9475 (N_9475,N_8307,N_8948);
nand U9476 (N_9476,N_8549,N_7621);
or U9477 (N_9477,N_8052,N_8585);
and U9478 (N_9478,N_8113,N_8027);
and U9479 (N_9479,N_7832,N_8438);
xor U9480 (N_9480,N_8706,N_7912);
xnor U9481 (N_9481,N_7575,N_8651);
or U9482 (N_9482,N_7949,N_8698);
or U9483 (N_9483,N_8293,N_7605);
nor U9484 (N_9484,N_8671,N_7642);
nor U9485 (N_9485,N_7593,N_8725);
and U9486 (N_9486,N_8466,N_8298);
or U9487 (N_9487,N_8863,N_8218);
or U9488 (N_9488,N_8087,N_8449);
nor U9489 (N_9489,N_7668,N_8731);
nand U9490 (N_9490,N_8764,N_7524);
nor U9491 (N_9491,N_8360,N_8736);
or U9492 (N_9492,N_7704,N_7545);
nor U9493 (N_9493,N_8559,N_8205);
nand U9494 (N_9494,N_8414,N_8703);
nor U9495 (N_9495,N_8954,N_8705);
nor U9496 (N_9496,N_7711,N_7561);
and U9497 (N_9497,N_8224,N_7641);
nor U9498 (N_9498,N_8932,N_8284);
or U9499 (N_9499,N_8023,N_7628);
nand U9500 (N_9500,N_8269,N_8984);
and U9501 (N_9501,N_8082,N_8286);
and U9502 (N_9502,N_8048,N_8426);
nand U9503 (N_9503,N_7891,N_8986);
and U9504 (N_9504,N_8946,N_8841);
nand U9505 (N_9505,N_8727,N_7583);
and U9506 (N_9506,N_8055,N_8693);
and U9507 (N_9507,N_8356,N_7582);
xnor U9508 (N_9508,N_7929,N_8799);
and U9509 (N_9509,N_8390,N_8384);
nor U9510 (N_9510,N_8648,N_7607);
xor U9511 (N_9511,N_8567,N_8095);
and U9512 (N_9512,N_8535,N_8790);
and U9513 (N_9513,N_8711,N_8679);
nor U9514 (N_9514,N_8661,N_8744);
nor U9515 (N_9515,N_8297,N_8937);
or U9516 (N_9516,N_8192,N_8760);
xor U9517 (N_9517,N_7749,N_7920);
or U9518 (N_9518,N_8333,N_8522);
or U9519 (N_9519,N_8058,N_8116);
nand U9520 (N_9520,N_7918,N_8035);
nor U9521 (N_9521,N_8607,N_8024);
and U9522 (N_9522,N_7868,N_8719);
nor U9523 (N_9523,N_8818,N_7813);
nand U9524 (N_9524,N_7848,N_8443);
or U9525 (N_9525,N_7687,N_8939);
or U9526 (N_9526,N_8317,N_7811);
nand U9527 (N_9527,N_7934,N_8366);
or U9528 (N_9528,N_7576,N_7984);
nand U9529 (N_9529,N_8936,N_8178);
nor U9530 (N_9530,N_8905,N_8540);
or U9531 (N_9531,N_7897,N_8974);
nand U9532 (N_9532,N_8584,N_8952);
nor U9533 (N_9533,N_8252,N_8674);
nand U9534 (N_9534,N_7674,N_8527);
and U9535 (N_9535,N_8166,N_7587);
xnor U9536 (N_9536,N_7782,N_8324);
xnor U9537 (N_9537,N_8961,N_8862);
and U9538 (N_9538,N_8247,N_8172);
and U9539 (N_9539,N_8656,N_7924);
and U9540 (N_9540,N_8626,N_7520);
and U9541 (N_9541,N_8979,N_7701);
nand U9542 (N_9542,N_8411,N_8125);
xor U9543 (N_9543,N_8322,N_8813);
nand U9544 (N_9544,N_7923,N_7585);
nand U9545 (N_9545,N_8868,N_8538);
nor U9546 (N_9546,N_7691,N_8601);
nor U9547 (N_9547,N_7509,N_7872);
and U9548 (N_9548,N_7619,N_8814);
nor U9549 (N_9549,N_8867,N_8400);
nor U9550 (N_9550,N_7672,N_8201);
and U9551 (N_9551,N_8689,N_8978);
and U9552 (N_9552,N_8126,N_7986);
nor U9553 (N_9553,N_8053,N_8604);
xor U9554 (N_9554,N_8462,N_8543);
and U9555 (N_9555,N_8049,N_8391);
or U9556 (N_9556,N_8525,N_8179);
nor U9557 (N_9557,N_7708,N_8130);
nor U9558 (N_9558,N_7864,N_8063);
or U9559 (N_9559,N_8504,N_8909);
nand U9560 (N_9560,N_7875,N_7830);
and U9561 (N_9561,N_7963,N_8263);
nor U9562 (N_9562,N_7954,N_7933);
nand U9563 (N_9563,N_7758,N_7609);
and U9564 (N_9564,N_7697,N_8779);
xor U9565 (N_9565,N_7602,N_8257);
xnor U9566 (N_9566,N_8236,N_7766);
xnor U9567 (N_9567,N_8031,N_8057);
nor U9568 (N_9568,N_8612,N_8660);
or U9569 (N_9569,N_8666,N_8888);
and U9570 (N_9570,N_8840,N_8832);
or U9571 (N_9571,N_8346,N_8683);
nor U9572 (N_9572,N_8548,N_7931);
and U9573 (N_9573,N_8713,N_8014);
xnor U9574 (N_9574,N_7975,N_8835);
or U9575 (N_9575,N_8222,N_7631);
and U9576 (N_9576,N_8701,N_7814);
xnor U9577 (N_9577,N_8071,N_7911);
or U9578 (N_9578,N_7767,N_8787);
or U9579 (N_9579,N_7531,N_7976);
nor U9580 (N_9580,N_8021,N_8283);
nand U9581 (N_9581,N_7626,N_7682);
nand U9582 (N_9582,N_7679,N_7504);
xnor U9583 (N_9583,N_8628,N_8735);
xnor U9584 (N_9584,N_7969,N_8232);
xor U9585 (N_9585,N_8442,N_7727);
or U9586 (N_9586,N_8911,N_7789);
and U9587 (N_9587,N_8362,N_7906);
nand U9588 (N_9588,N_8798,N_8638);
nand U9589 (N_9589,N_8721,N_7795);
nor U9590 (N_9590,N_8633,N_7754);
nand U9591 (N_9591,N_8114,N_8395);
xnor U9592 (N_9592,N_8929,N_7528);
or U9593 (N_9593,N_8320,N_7967);
nor U9594 (N_9594,N_7523,N_7860);
and U9595 (N_9595,N_8266,N_8233);
nor U9596 (N_9596,N_8542,N_7595);
or U9597 (N_9597,N_8590,N_8169);
nor U9598 (N_9598,N_8267,N_7946);
and U9599 (N_9599,N_7538,N_8019);
nand U9600 (N_9600,N_7803,N_8304);
nand U9601 (N_9601,N_8194,N_7739);
and U9602 (N_9602,N_8475,N_7792);
xor U9603 (N_9603,N_7818,N_8299);
and U9604 (N_9604,N_8123,N_8454);
xor U9605 (N_9605,N_8897,N_8010);
nor U9606 (N_9606,N_7539,N_8632);
and U9607 (N_9607,N_8160,N_7518);
nor U9608 (N_9608,N_8781,N_8185);
or U9609 (N_9609,N_8131,N_8176);
nand U9610 (N_9610,N_8288,N_8136);
or U9611 (N_9611,N_8843,N_8354);
and U9612 (N_9612,N_8407,N_8960);
nand U9613 (N_9613,N_8505,N_8156);
and U9614 (N_9614,N_7706,N_7913);
or U9615 (N_9615,N_8778,N_8158);
or U9616 (N_9616,N_7829,N_7944);
xor U9617 (N_9617,N_8943,N_7571);
and U9618 (N_9618,N_8754,N_8955);
or U9619 (N_9619,N_7599,N_7580);
nand U9620 (N_9620,N_8394,N_7546);
and U9621 (N_9621,N_8753,N_8775);
nor U9622 (N_9622,N_8699,N_7657);
xor U9623 (N_9623,N_7543,N_8456);
and U9624 (N_9624,N_8555,N_8467);
nand U9625 (N_9625,N_8769,N_8530);
xnor U9626 (N_9626,N_7982,N_8041);
or U9627 (N_9627,N_8129,N_8745);
nor U9628 (N_9628,N_8221,N_8091);
xor U9629 (N_9629,N_7901,N_8479);
nor U9630 (N_9630,N_8408,N_7959);
or U9631 (N_9631,N_7922,N_7909);
and U9632 (N_9632,N_8416,N_8983);
nand U9633 (N_9633,N_8484,N_8916);
xor U9634 (N_9634,N_8255,N_7988);
or U9635 (N_9635,N_7799,N_8718);
nor U9636 (N_9636,N_8723,N_8746);
xnor U9637 (N_9637,N_8757,N_8624);
xor U9638 (N_9638,N_7738,N_8537);
or U9639 (N_9639,N_8564,N_8037);
xor U9640 (N_9640,N_8587,N_8080);
xor U9641 (N_9641,N_8595,N_7877);
nand U9642 (N_9642,N_8972,N_8225);
xor U9643 (N_9643,N_8820,N_8834);
nand U9644 (N_9644,N_8557,N_8962);
xor U9645 (N_9645,N_8856,N_8849);
or U9646 (N_9646,N_8196,N_8500);
nor U9647 (N_9647,N_7566,N_8956);
or U9648 (N_9648,N_8030,N_8000);
and U9649 (N_9649,N_7940,N_7873);
nand U9650 (N_9650,N_8741,N_8347);
nor U9651 (N_9651,N_8617,N_8508);
and U9652 (N_9652,N_7824,N_7654);
nand U9653 (N_9653,N_7784,N_8831);
or U9654 (N_9654,N_8319,N_8623);
or U9655 (N_9655,N_8570,N_7854);
or U9656 (N_9656,N_8093,N_8265);
or U9657 (N_9657,N_8374,N_8204);
or U9658 (N_9658,N_7702,N_8614);
xnor U9659 (N_9659,N_7634,N_8677);
and U9660 (N_9660,N_8806,N_7936);
xor U9661 (N_9661,N_8250,N_8381);
xor U9662 (N_9662,N_8599,N_8413);
nor U9663 (N_9663,N_8231,N_7790);
xor U9664 (N_9664,N_8203,N_7846);
or U9665 (N_9665,N_7816,N_7908);
or U9666 (N_9666,N_7981,N_8132);
and U9667 (N_9667,N_7637,N_7821);
xnor U9668 (N_9668,N_8765,N_8822);
nor U9669 (N_9669,N_8642,N_8447);
xnor U9670 (N_9670,N_8437,N_7970);
nand U9671 (N_9671,N_8056,N_8511);
or U9672 (N_9672,N_7851,N_8510);
and U9673 (N_9673,N_7653,N_8917);
nand U9674 (N_9674,N_7900,N_7914);
xnor U9675 (N_9675,N_8665,N_7849);
or U9676 (N_9676,N_8170,N_8680);
nand U9677 (N_9677,N_8077,N_7651);
and U9678 (N_9678,N_8189,N_7601);
nor U9679 (N_9679,N_7503,N_8157);
and U9680 (N_9680,N_8042,N_8478);
nand U9681 (N_9681,N_7530,N_8647);
nand U9682 (N_9682,N_7733,N_8861);
nor U9683 (N_9683,N_7794,N_7757);
and U9684 (N_9684,N_8107,N_8143);
and U9685 (N_9685,N_8312,N_8724);
or U9686 (N_9686,N_8786,N_7853);
or U9687 (N_9687,N_8795,N_8228);
xnor U9688 (N_9688,N_8659,N_7683);
nand U9689 (N_9689,N_7948,N_8001);
nor U9690 (N_9690,N_8309,N_8889);
and U9691 (N_9691,N_7617,N_8214);
xnor U9692 (N_9692,N_8465,N_7588);
xnor U9693 (N_9693,N_8578,N_8274);
and U9694 (N_9694,N_8998,N_8459);
or U9695 (N_9695,N_7863,N_7703);
and U9696 (N_9696,N_8801,N_7837);
or U9697 (N_9697,N_8406,N_7551);
xor U9698 (N_9698,N_8536,N_7506);
xor U9699 (N_9699,N_7762,N_8073);
nand U9700 (N_9700,N_8043,N_8403);
nand U9701 (N_9701,N_7735,N_8520);
nor U9702 (N_9702,N_7835,N_8667);
nand U9703 (N_9703,N_7734,N_8337);
nor U9704 (N_9704,N_8768,N_7989);
or U9705 (N_9705,N_8697,N_7690);
nand U9706 (N_9706,N_8678,N_8425);
nor U9707 (N_9707,N_8996,N_7515);
and U9708 (N_9708,N_7785,N_8816);
and U9709 (N_9709,N_8958,N_7825);
and U9710 (N_9710,N_7597,N_8184);
or U9711 (N_9711,N_8777,N_8328);
xor U9712 (N_9712,N_8720,N_8060);
or U9713 (N_9713,N_8318,N_8069);
nor U9714 (N_9714,N_8369,N_8177);
and U9715 (N_9715,N_8785,N_8450);
nand U9716 (N_9716,N_8445,N_7611);
nor U9717 (N_9717,N_7742,N_8603);
and U9718 (N_9718,N_8625,N_7572);
and U9719 (N_9719,N_8528,N_8434);
nand U9720 (N_9720,N_7925,N_8550);
and U9721 (N_9721,N_8829,N_8935);
xnor U9722 (N_9722,N_8289,N_8367);
or U9723 (N_9723,N_8253,N_7838);
nand U9724 (N_9724,N_8869,N_8923);
xor U9725 (N_9725,N_8089,N_8997);
xnor U9726 (N_9726,N_8455,N_8915);
and U9727 (N_9727,N_8332,N_8898);
nor U9728 (N_9728,N_8241,N_7977);
nand U9729 (N_9729,N_8207,N_8431);
nor U9730 (N_9730,N_8568,N_8290);
xnor U9731 (N_9731,N_7928,N_8615);
nand U9732 (N_9732,N_7995,N_8934);
nand U9733 (N_9733,N_8480,N_7740);
nor U9734 (N_9734,N_8673,N_8209);
nor U9735 (N_9735,N_7746,N_8261);
nor U9736 (N_9736,N_8273,N_7664);
nor U9737 (N_9737,N_8469,N_8017);
nand U9738 (N_9738,N_8054,N_8837);
xor U9739 (N_9739,N_8529,N_8634);
or U9740 (N_9740,N_7560,N_8491);
nand U9741 (N_9741,N_7769,N_8899);
xor U9742 (N_9742,N_8405,N_7647);
or U9743 (N_9743,N_8240,N_7570);
or U9744 (N_9744,N_7667,N_8075);
nand U9745 (N_9745,N_8198,N_7917);
xnor U9746 (N_9746,N_8702,N_8294);
or U9747 (N_9747,N_8924,N_7574);
nor U9748 (N_9748,N_8545,N_8020);
nand U9749 (N_9749,N_7590,N_8838);
nor U9750 (N_9750,N_7664,N_7799);
or U9751 (N_9751,N_8205,N_7694);
xor U9752 (N_9752,N_8623,N_7825);
xor U9753 (N_9753,N_8901,N_7831);
nor U9754 (N_9754,N_8196,N_8648);
xor U9755 (N_9755,N_8798,N_8731);
xor U9756 (N_9756,N_7793,N_7855);
nor U9757 (N_9757,N_8062,N_8932);
nor U9758 (N_9758,N_8092,N_8983);
nor U9759 (N_9759,N_7638,N_7889);
and U9760 (N_9760,N_8235,N_7958);
or U9761 (N_9761,N_7811,N_8998);
or U9762 (N_9762,N_7859,N_8785);
nand U9763 (N_9763,N_8057,N_8850);
or U9764 (N_9764,N_8690,N_8618);
xor U9765 (N_9765,N_8702,N_8873);
nand U9766 (N_9766,N_8172,N_8239);
nor U9767 (N_9767,N_8972,N_8333);
nand U9768 (N_9768,N_8160,N_8393);
nor U9769 (N_9769,N_8116,N_7767);
nand U9770 (N_9770,N_7862,N_8687);
nor U9771 (N_9771,N_8208,N_8281);
nand U9772 (N_9772,N_7506,N_7708);
or U9773 (N_9773,N_7952,N_7516);
and U9774 (N_9774,N_7874,N_8544);
nor U9775 (N_9775,N_8881,N_8275);
xnor U9776 (N_9776,N_7574,N_8587);
and U9777 (N_9777,N_8688,N_8193);
xor U9778 (N_9778,N_8773,N_8020);
xnor U9779 (N_9779,N_8499,N_7930);
or U9780 (N_9780,N_7687,N_8527);
or U9781 (N_9781,N_8299,N_7810);
nand U9782 (N_9782,N_8035,N_8702);
xnor U9783 (N_9783,N_7917,N_8028);
nand U9784 (N_9784,N_8415,N_8380);
xor U9785 (N_9785,N_8153,N_8535);
nor U9786 (N_9786,N_8771,N_8370);
or U9787 (N_9787,N_8369,N_8877);
and U9788 (N_9788,N_8691,N_7515);
and U9789 (N_9789,N_8101,N_7667);
or U9790 (N_9790,N_8956,N_8718);
nor U9791 (N_9791,N_8662,N_8904);
and U9792 (N_9792,N_7858,N_8614);
and U9793 (N_9793,N_7555,N_8281);
xor U9794 (N_9794,N_8622,N_8890);
nand U9795 (N_9795,N_8219,N_8990);
xor U9796 (N_9796,N_8121,N_8162);
and U9797 (N_9797,N_8777,N_8601);
and U9798 (N_9798,N_8278,N_7936);
nand U9799 (N_9799,N_7986,N_7930);
nand U9800 (N_9800,N_7633,N_7721);
nand U9801 (N_9801,N_8631,N_8502);
xnor U9802 (N_9802,N_8487,N_7985);
nor U9803 (N_9803,N_7952,N_7636);
or U9804 (N_9804,N_8718,N_8503);
and U9805 (N_9805,N_7602,N_8572);
nor U9806 (N_9806,N_7865,N_7971);
and U9807 (N_9807,N_8824,N_7667);
and U9808 (N_9808,N_7898,N_8597);
nand U9809 (N_9809,N_8682,N_8262);
xnor U9810 (N_9810,N_8633,N_8363);
nand U9811 (N_9811,N_8504,N_8430);
and U9812 (N_9812,N_8995,N_8181);
nor U9813 (N_9813,N_8912,N_8985);
nand U9814 (N_9814,N_7839,N_8033);
and U9815 (N_9815,N_8110,N_8930);
nand U9816 (N_9816,N_7852,N_7595);
nor U9817 (N_9817,N_7653,N_7935);
and U9818 (N_9818,N_8535,N_8171);
and U9819 (N_9819,N_8510,N_7666);
nand U9820 (N_9820,N_7722,N_8526);
nor U9821 (N_9821,N_7755,N_7506);
and U9822 (N_9822,N_8196,N_7889);
or U9823 (N_9823,N_7813,N_7908);
xnor U9824 (N_9824,N_7570,N_8866);
xor U9825 (N_9825,N_8219,N_8108);
xnor U9826 (N_9826,N_8928,N_8170);
nand U9827 (N_9827,N_8903,N_8023);
nor U9828 (N_9828,N_8334,N_8140);
nor U9829 (N_9829,N_7798,N_8967);
nor U9830 (N_9830,N_8377,N_8060);
nand U9831 (N_9831,N_8643,N_8465);
nor U9832 (N_9832,N_8970,N_7931);
nand U9833 (N_9833,N_8085,N_8868);
or U9834 (N_9834,N_8736,N_7864);
or U9835 (N_9835,N_8563,N_8591);
xnor U9836 (N_9836,N_8016,N_7550);
or U9837 (N_9837,N_8223,N_8534);
nand U9838 (N_9838,N_8672,N_8284);
nand U9839 (N_9839,N_8144,N_8421);
nor U9840 (N_9840,N_8542,N_8509);
xor U9841 (N_9841,N_7897,N_8678);
and U9842 (N_9842,N_8313,N_8394);
xor U9843 (N_9843,N_8743,N_7662);
and U9844 (N_9844,N_8681,N_7856);
xnor U9845 (N_9845,N_8692,N_8741);
or U9846 (N_9846,N_8015,N_7578);
nand U9847 (N_9847,N_8714,N_8782);
nand U9848 (N_9848,N_8277,N_7987);
nor U9849 (N_9849,N_8004,N_8317);
nand U9850 (N_9850,N_8512,N_8176);
nor U9851 (N_9851,N_8548,N_7593);
nand U9852 (N_9852,N_7629,N_7568);
nand U9853 (N_9853,N_7800,N_8763);
or U9854 (N_9854,N_7512,N_8264);
nand U9855 (N_9855,N_8689,N_8156);
nor U9856 (N_9856,N_8160,N_8788);
or U9857 (N_9857,N_8634,N_8710);
xor U9858 (N_9858,N_8243,N_8972);
nand U9859 (N_9859,N_8399,N_8710);
nor U9860 (N_9860,N_7606,N_8854);
xnor U9861 (N_9861,N_7656,N_8258);
xor U9862 (N_9862,N_8237,N_8698);
nand U9863 (N_9863,N_8086,N_8943);
nor U9864 (N_9864,N_8725,N_7722);
xnor U9865 (N_9865,N_8293,N_8344);
nand U9866 (N_9866,N_8081,N_7871);
nor U9867 (N_9867,N_8831,N_8406);
and U9868 (N_9868,N_8847,N_8990);
nand U9869 (N_9869,N_8991,N_8932);
xor U9870 (N_9870,N_8421,N_8285);
xnor U9871 (N_9871,N_8575,N_8063);
and U9872 (N_9872,N_7834,N_8949);
nor U9873 (N_9873,N_8896,N_8242);
and U9874 (N_9874,N_8166,N_8216);
or U9875 (N_9875,N_8922,N_8165);
xor U9876 (N_9876,N_8939,N_8848);
and U9877 (N_9877,N_8020,N_7793);
and U9878 (N_9878,N_8206,N_8968);
and U9879 (N_9879,N_8626,N_7774);
nand U9880 (N_9880,N_8037,N_8580);
and U9881 (N_9881,N_8691,N_7667);
or U9882 (N_9882,N_7603,N_8421);
and U9883 (N_9883,N_7877,N_7631);
nand U9884 (N_9884,N_8008,N_8703);
or U9885 (N_9885,N_8059,N_8482);
and U9886 (N_9886,N_8172,N_8166);
nor U9887 (N_9887,N_7504,N_7532);
xor U9888 (N_9888,N_8267,N_8382);
nor U9889 (N_9889,N_7807,N_8420);
nand U9890 (N_9890,N_8387,N_7875);
and U9891 (N_9891,N_7609,N_8522);
nor U9892 (N_9892,N_8470,N_8371);
and U9893 (N_9893,N_8682,N_7604);
and U9894 (N_9894,N_8627,N_7879);
and U9895 (N_9895,N_8503,N_7800);
xor U9896 (N_9896,N_7534,N_7571);
and U9897 (N_9897,N_8912,N_8816);
nand U9898 (N_9898,N_8035,N_7798);
and U9899 (N_9899,N_8860,N_8911);
nor U9900 (N_9900,N_7669,N_8170);
and U9901 (N_9901,N_8372,N_8302);
nor U9902 (N_9902,N_7557,N_8853);
nor U9903 (N_9903,N_8363,N_8574);
or U9904 (N_9904,N_8560,N_7835);
or U9905 (N_9905,N_8477,N_7966);
nor U9906 (N_9906,N_8164,N_8671);
or U9907 (N_9907,N_8992,N_8961);
and U9908 (N_9908,N_8649,N_7620);
and U9909 (N_9909,N_8930,N_8293);
nor U9910 (N_9910,N_8529,N_8401);
nor U9911 (N_9911,N_7704,N_8425);
nor U9912 (N_9912,N_8295,N_7537);
nand U9913 (N_9913,N_7821,N_8192);
or U9914 (N_9914,N_8255,N_7885);
xnor U9915 (N_9915,N_7613,N_8867);
nor U9916 (N_9916,N_8419,N_8167);
or U9917 (N_9917,N_8620,N_8683);
or U9918 (N_9918,N_8916,N_8750);
and U9919 (N_9919,N_8295,N_8042);
or U9920 (N_9920,N_8050,N_7550);
nor U9921 (N_9921,N_8412,N_8300);
or U9922 (N_9922,N_7992,N_8410);
or U9923 (N_9923,N_7988,N_7834);
and U9924 (N_9924,N_8170,N_7812);
and U9925 (N_9925,N_7799,N_7964);
or U9926 (N_9926,N_8980,N_8626);
or U9927 (N_9927,N_8396,N_7983);
xor U9928 (N_9928,N_8632,N_7678);
nor U9929 (N_9929,N_7505,N_8284);
nand U9930 (N_9930,N_7718,N_8625);
or U9931 (N_9931,N_8216,N_8424);
xor U9932 (N_9932,N_8521,N_8208);
or U9933 (N_9933,N_7729,N_8159);
and U9934 (N_9934,N_8940,N_8755);
nor U9935 (N_9935,N_8289,N_8339);
xnor U9936 (N_9936,N_8639,N_8095);
nand U9937 (N_9937,N_8800,N_8817);
nor U9938 (N_9938,N_8952,N_7633);
nor U9939 (N_9939,N_7787,N_8997);
xnor U9940 (N_9940,N_8205,N_7831);
nand U9941 (N_9941,N_7969,N_8086);
or U9942 (N_9942,N_8106,N_8133);
and U9943 (N_9943,N_8318,N_7798);
nor U9944 (N_9944,N_8160,N_8879);
nor U9945 (N_9945,N_7859,N_8989);
xnor U9946 (N_9946,N_8907,N_7528);
or U9947 (N_9947,N_8406,N_7783);
and U9948 (N_9948,N_8076,N_7933);
nand U9949 (N_9949,N_8152,N_8849);
nand U9950 (N_9950,N_8398,N_8845);
or U9951 (N_9951,N_8070,N_8912);
nand U9952 (N_9952,N_8282,N_8407);
or U9953 (N_9953,N_8103,N_7712);
nor U9954 (N_9954,N_8121,N_8898);
or U9955 (N_9955,N_7685,N_8382);
or U9956 (N_9956,N_8762,N_8168);
nand U9957 (N_9957,N_7650,N_7533);
or U9958 (N_9958,N_8988,N_8025);
nand U9959 (N_9959,N_8285,N_8019);
and U9960 (N_9960,N_8778,N_8923);
xnor U9961 (N_9961,N_8286,N_8816);
nand U9962 (N_9962,N_8565,N_8938);
and U9963 (N_9963,N_7714,N_8541);
nand U9964 (N_9964,N_8848,N_7655);
nor U9965 (N_9965,N_7558,N_8161);
nand U9966 (N_9966,N_8329,N_8532);
xnor U9967 (N_9967,N_8335,N_7508);
or U9968 (N_9968,N_7812,N_8975);
and U9969 (N_9969,N_7676,N_7631);
nand U9970 (N_9970,N_8486,N_8886);
and U9971 (N_9971,N_7728,N_8621);
nand U9972 (N_9972,N_8178,N_8103);
nand U9973 (N_9973,N_7879,N_8631);
xnor U9974 (N_9974,N_8170,N_8166);
xor U9975 (N_9975,N_8835,N_8293);
xnor U9976 (N_9976,N_8628,N_7918);
nor U9977 (N_9977,N_8820,N_7866);
or U9978 (N_9978,N_8837,N_8821);
nor U9979 (N_9979,N_8395,N_8583);
nor U9980 (N_9980,N_8957,N_8894);
xnor U9981 (N_9981,N_8999,N_8907);
xor U9982 (N_9982,N_8271,N_8556);
nor U9983 (N_9983,N_8895,N_8387);
xnor U9984 (N_9984,N_7848,N_7774);
or U9985 (N_9985,N_7844,N_8318);
nand U9986 (N_9986,N_8593,N_7804);
or U9987 (N_9987,N_8019,N_7568);
and U9988 (N_9988,N_8716,N_7612);
nand U9989 (N_9989,N_7831,N_8974);
nor U9990 (N_9990,N_8326,N_8379);
xnor U9991 (N_9991,N_7565,N_7564);
and U9992 (N_9992,N_7605,N_8850);
xor U9993 (N_9993,N_8167,N_8591);
nor U9994 (N_9994,N_8800,N_7582);
nor U9995 (N_9995,N_8128,N_8256);
and U9996 (N_9996,N_7900,N_8401);
and U9997 (N_9997,N_7734,N_7711);
nor U9998 (N_9998,N_8734,N_7602);
or U9999 (N_9999,N_8303,N_8481);
nor U10000 (N_10000,N_8043,N_7556);
xnor U10001 (N_10001,N_8638,N_8320);
xnor U10002 (N_10002,N_7991,N_8503);
or U10003 (N_10003,N_8065,N_8546);
or U10004 (N_10004,N_8985,N_8251);
xor U10005 (N_10005,N_8563,N_8164);
and U10006 (N_10006,N_8431,N_8106);
xnor U10007 (N_10007,N_8853,N_8019);
xnor U10008 (N_10008,N_7972,N_8529);
nand U10009 (N_10009,N_8133,N_7594);
xnor U10010 (N_10010,N_8932,N_8257);
or U10011 (N_10011,N_7903,N_8654);
or U10012 (N_10012,N_8006,N_8801);
xnor U10013 (N_10013,N_8104,N_7896);
xor U10014 (N_10014,N_7727,N_8844);
or U10015 (N_10015,N_7599,N_8709);
nand U10016 (N_10016,N_8561,N_8651);
nand U10017 (N_10017,N_7793,N_7712);
nand U10018 (N_10018,N_8298,N_7602);
and U10019 (N_10019,N_7670,N_8582);
nor U10020 (N_10020,N_7566,N_8530);
or U10021 (N_10021,N_8304,N_7534);
or U10022 (N_10022,N_8564,N_8626);
nor U10023 (N_10023,N_7749,N_8381);
nand U10024 (N_10024,N_8073,N_8821);
xor U10025 (N_10025,N_8421,N_8615);
nand U10026 (N_10026,N_8703,N_8954);
nand U10027 (N_10027,N_8341,N_8323);
nor U10028 (N_10028,N_8872,N_8440);
xnor U10029 (N_10029,N_8663,N_8871);
nor U10030 (N_10030,N_7900,N_8360);
nor U10031 (N_10031,N_8844,N_7702);
or U10032 (N_10032,N_7939,N_8859);
and U10033 (N_10033,N_8141,N_8722);
nand U10034 (N_10034,N_8487,N_8943);
nand U10035 (N_10035,N_8823,N_8703);
nand U10036 (N_10036,N_8205,N_8119);
nand U10037 (N_10037,N_8712,N_7991);
and U10038 (N_10038,N_8912,N_8417);
and U10039 (N_10039,N_8600,N_8540);
and U10040 (N_10040,N_8458,N_8513);
and U10041 (N_10041,N_8905,N_7923);
and U10042 (N_10042,N_8335,N_8902);
or U10043 (N_10043,N_8809,N_7996);
nor U10044 (N_10044,N_8418,N_7930);
and U10045 (N_10045,N_8958,N_7753);
xnor U10046 (N_10046,N_7756,N_8031);
and U10047 (N_10047,N_7551,N_8329);
nor U10048 (N_10048,N_8723,N_7893);
nor U10049 (N_10049,N_8500,N_8431);
and U10050 (N_10050,N_8592,N_7809);
and U10051 (N_10051,N_8867,N_8376);
or U10052 (N_10052,N_8647,N_8902);
and U10053 (N_10053,N_8596,N_8392);
nand U10054 (N_10054,N_7500,N_7759);
nor U10055 (N_10055,N_7979,N_7531);
nor U10056 (N_10056,N_8190,N_8391);
or U10057 (N_10057,N_7525,N_8967);
nand U10058 (N_10058,N_8706,N_7849);
nand U10059 (N_10059,N_7543,N_8625);
or U10060 (N_10060,N_8633,N_8272);
xnor U10061 (N_10061,N_8813,N_7931);
nor U10062 (N_10062,N_7825,N_7877);
and U10063 (N_10063,N_8722,N_8369);
xnor U10064 (N_10064,N_8048,N_8296);
xnor U10065 (N_10065,N_8934,N_7923);
nand U10066 (N_10066,N_8949,N_8451);
nand U10067 (N_10067,N_8215,N_8219);
and U10068 (N_10068,N_8364,N_7691);
or U10069 (N_10069,N_7544,N_8069);
nand U10070 (N_10070,N_7589,N_7674);
nand U10071 (N_10071,N_8365,N_8191);
nand U10072 (N_10072,N_8875,N_7837);
nand U10073 (N_10073,N_8135,N_7586);
nor U10074 (N_10074,N_8291,N_8515);
nand U10075 (N_10075,N_8095,N_8807);
xor U10076 (N_10076,N_8058,N_8876);
nor U10077 (N_10077,N_7563,N_7543);
nor U10078 (N_10078,N_7791,N_8069);
or U10079 (N_10079,N_8373,N_8662);
and U10080 (N_10080,N_8008,N_7590);
nor U10081 (N_10081,N_7796,N_8648);
nand U10082 (N_10082,N_7675,N_8692);
or U10083 (N_10083,N_7645,N_8767);
xor U10084 (N_10084,N_7685,N_8254);
xnor U10085 (N_10085,N_7615,N_7889);
nand U10086 (N_10086,N_8522,N_8854);
xor U10087 (N_10087,N_7818,N_8470);
nor U10088 (N_10088,N_8052,N_7627);
nor U10089 (N_10089,N_7763,N_8083);
and U10090 (N_10090,N_8614,N_8678);
nand U10091 (N_10091,N_8710,N_7508);
and U10092 (N_10092,N_7509,N_8217);
nand U10093 (N_10093,N_8618,N_8966);
nor U10094 (N_10094,N_7539,N_7659);
nand U10095 (N_10095,N_8684,N_8553);
nand U10096 (N_10096,N_7523,N_8462);
or U10097 (N_10097,N_7604,N_8839);
xor U10098 (N_10098,N_7606,N_8659);
or U10099 (N_10099,N_7782,N_8390);
or U10100 (N_10100,N_8811,N_7742);
nor U10101 (N_10101,N_7816,N_8800);
xor U10102 (N_10102,N_8474,N_8689);
and U10103 (N_10103,N_8140,N_8944);
nor U10104 (N_10104,N_7869,N_7609);
and U10105 (N_10105,N_7806,N_8305);
and U10106 (N_10106,N_8600,N_8007);
and U10107 (N_10107,N_8800,N_8053);
and U10108 (N_10108,N_8005,N_8387);
xnor U10109 (N_10109,N_8322,N_8468);
nand U10110 (N_10110,N_8993,N_8816);
nand U10111 (N_10111,N_8347,N_8920);
and U10112 (N_10112,N_7580,N_8378);
or U10113 (N_10113,N_7693,N_8754);
or U10114 (N_10114,N_8164,N_8061);
xor U10115 (N_10115,N_8172,N_8233);
nand U10116 (N_10116,N_8617,N_8223);
nor U10117 (N_10117,N_8562,N_7530);
and U10118 (N_10118,N_7975,N_8006);
nor U10119 (N_10119,N_8326,N_7791);
and U10120 (N_10120,N_8667,N_8360);
or U10121 (N_10121,N_8431,N_8866);
and U10122 (N_10122,N_8520,N_8752);
and U10123 (N_10123,N_8559,N_7852);
nor U10124 (N_10124,N_7915,N_7797);
or U10125 (N_10125,N_8723,N_8442);
nor U10126 (N_10126,N_8469,N_8333);
or U10127 (N_10127,N_8687,N_8419);
or U10128 (N_10128,N_7942,N_8096);
xor U10129 (N_10129,N_7789,N_8686);
or U10130 (N_10130,N_8503,N_8846);
nand U10131 (N_10131,N_8690,N_8486);
or U10132 (N_10132,N_7738,N_8614);
and U10133 (N_10133,N_8664,N_8204);
nor U10134 (N_10134,N_8211,N_8181);
or U10135 (N_10135,N_8920,N_8529);
xnor U10136 (N_10136,N_8477,N_8337);
xor U10137 (N_10137,N_7750,N_7628);
nor U10138 (N_10138,N_8330,N_8813);
xor U10139 (N_10139,N_7901,N_7882);
or U10140 (N_10140,N_7826,N_8614);
and U10141 (N_10141,N_8540,N_8547);
and U10142 (N_10142,N_7645,N_8456);
nand U10143 (N_10143,N_8752,N_8580);
and U10144 (N_10144,N_8751,N_7654);
nor U10145 (N_10145,N_7556,N_8061);
xnor U10146 (N_10146,N_8300,N_7936);
xnor U10147 (N_10147,N_8227,N_8414);
or U10148 (N_10148,N_8299,N_7928);
and U10149 (N_10149,N_8873,N_8938);
xor U10150 (N_10150,N_8435,N_8803);
nor U10151 (N_10151,N_8961,N_7692);
nor U10152 (N_10152,N_7859,N_8356);
nor U10153 (N_10153,N_8060,N_8453);
nor U10154 (N_10154,N_8153,N_8425);
nand U10155 (N_10155,N_7949,N_8044);
nor U10156 (N_10156,N_7991,N_8440);
nand U10157 (N_10157,N_8569,N_8623);
nor U10158 (N_10158,N_8947,N_7546);
or U10159 (N_10159,N_8146,N_8178);
xnor U10160 (N_10160,N_8630,N_8521);
nor U10161 (N_10161,N_8506,N_8116);
xor U10162 (N_10162,N_8176,N_7572);
or U10163 (N_10163,N_8944,N_8740);
and U10164 (N_10164,N_8002,N_8692);
and U10165 (N_10165,N_7729,N_8717);
and U10166 (N_10166,N_7900,N_8531);
nor U10167 (N_10167,N_8105,N_7775);
and U10168 (N_10168,N_8802,N_8322);
nor U10169 (N_10169,N_7774,N_8325);
nor U10170 (N_10170,N_8897,N_8012);
nand U10171 (N_10171,N_8339,N_8484);
or U10172 (N_10172,N_8595,N_7832);
or U10173 (N_10173,N_8698,N_7834);
nor U10174 (N_10174,N_7783,N_7873);
nand U10175 (N_10175,N_8044,N_8427);
nand U10176 (N_10176,N_7625,N_8817);
or U10177 (N_10177,N_8794,N_7662);
xnor U10178 (N_10178,N_8924,N_8245);
xor U10179 (N_10179,N_8019,N_7509);
and U10180 (N_10180,N_8610,N_7558);
nand U10181 (N_10181,N_8727,N_8332);
xor U10182 (N_10182,N_8594,N_7977);
xnor U10183 (N_10183,N_8113,N_7605);
xor U10184 (N_10184,N_8988,N_7633);
nor U10185 (N_10185,N_7870,N_8336);
nor U10186 (N_10186,N_8324,N_7799);
or U10187 (N_10187,N_8136,N_8088);
nand U10188 (N_10188,N_7665,N_8185);
nand U10189 (N_10189,N_7775,N_8438);
xnor U10190 (N_10190,N_8969,N_8231);
or U10191 (N_10191,N_8358,N_7658);
xor U10192 (N_10192,N_8451,N_8832);
nand U10193 (N_10193,N_8158,N_8153);
nor U10194 (N_10194,N_8094,N_7922);
xor U10195 (N_10195,N_7657,N_8100);
and U10196 (N_10196,N_8567,N_8865);
nor U10197 (N_10197,N_8379,N_8222);
xor U10198 (N_10198,N_8938,N_7835);
xor U10199 (N_10199,N_8387,N_7831);
and U10200 (N_10200,N_8990,N_7840);
nand U10201 (N_10201,N_7605,N_8244);
or U10202 (N_10202,N_8670,N_8398);
nor U10203 (N_10203,N_7718,N_7662);
nor U10204 (N_10204,N_8244,N_8685);
xnor U10205 (N_10205,N_8014,N_8534);
xnor U10206 (N_10206,N_8441,N_8806);
xor U10207 (N_10207,N_8732,N_7661);
or U10208 (N_10208,N_7992,N_7610);
or U10209 (N_10209,N_7704,N_8397);
or U10210 (N_10210,N_8583,N_7763);
and U10211 (N_10211,N_8179,N_8967);
and U10212 (N_10212,N_8458,N_8564);
nand U10213 (N_10213,N_8058,N_8141);
nand U10214 (N_10214,N_7612,N_7856);
or U10215 (N_10215,N_8314,N_8055);
and U10216 (N_10216,N_8059,N_7941);
or U10217 (N_10217,N_8501,N_8831);
nand U10218 (N_10218,N_7891,N_7991);
nor U10219 (N_10219,N_7516,N_7856);
and U10220 (N_10220,N_8758,N_8544);
and U10221 (N_10221,N_8898,N_7843);
or U10222 (N_10222,N_8194,N_8479);
nor U10223 (N_10223,N_8405,N_8196);
or U10224 (N_10224,N_8172,N_7886);
or U10225 (N_10225,N_7727,N_8752);
nor U10226 (N_10226,N_8481,N_7573);
xor U10227 (N_10227,N_8699,N_8627);
nor U10228 (N_10228,N_8029,N_7528);
or U10229 (N_10229,N_8909,N_7534);
nor U10230 (N_10230,N_7965,N_8032);
or U10231 (N_10231,N_8708,N_8194);
or U10232 (N_10232,N_8801,N_8654);
nor U10233 (N_10233,N_8994,N_7603);
nand U10234 (N_10234,N_8958,N_8842);
nor U10235 (N_10235,N_8472,N_7594);
xor U10236 (N_10236,N_8427,N_8825);
xor U10237 (N_10237,N_8932,N_7803);
nor U10238 (N_10238,N_7966,N_8240);
nand U10239 (N_10239,N_7671,N_7857);
nor U10240 (N_10240,N_8082,N_8468);
or U10241 (N_10241,N_8654,N_8822);
nand U10242 (N_10242,N_8492,N_7899);
and U10243 (N_10243,N_7650,N_8467);
nor U10244 (N_10244,N_8588,N_8012);
nand U10245 (N_10245,N_7598,N_8755);
nor U10246 (N_10246,N_8335,N_8211);
and U10247 (N_10247,N_8631,N_8820);
or U10248 (N_10248,N_8854,N_7656);
nand U10249 (N_10249,N_8922,N_8659);
or U10250 (N_10250,N_8530,N_7526);
xor U10251 (N_10251,N_8196,N_7829);
xor U10252 (N_10252,N_8678,N_8189);
nand U10253 (N_10253,N_8532,N_8257);
or U10254 (N_10254,N_8400,N_8669);
nand U10255 (N_10255,N_8974,N_8006);
xor U10256 (N_10256,N_8429,N_7787);
and U10257 (N_10257,N_8927,N_8264);
xor U10258 (N_10258,N_7968,N_7831);
nor U10259 (N_10259,N_8621,N_7844);
xor U10260 (N_10260,N_7853,N_8105);
or U10261 (N_10261,N_8033,N_8460);
and U10262 (N_10262,N_7768,N_7589);
nand U10263 (N_10263,N_8650,N_8266);
and U10264 (N_10264,N_7542,N_7865);
xnor U10265 (N_10265,N_8823,N_8039);
xnor U10266 (N_10266,N_8911,N_8299);
and U10267 (N_10267,N_8882,N_8172);
xnor U10268 (N_10268,N_8766,N_7839);
nor U10269 (N_10269,N_8370,N_8502);
and U10270 (N_10270,N_8994,N_8921);
or U10271 (N_10271,N_8863,N_7773);
or U10272 (N_10272,N_7875,N_8786);
nor U10273 (N_10273,N_8363,N_7922);
and U10274 (N_10274,N_8436,N_8869);
nor U10275 (N_10275,N_7910,N_7636);
or U10276 (N_10276,N_7655,N_8798);
nor U10277 (N_10277,N_8590,N_8821);
or U10278 (N_10278,N_7561,N_7793);
and U10279 (N_10279,N_7831,N_7561);
and U10280 (N_10280,N_8108,N_8891);
xnor U10281 (N_10281,N_8417,N_8301);
and U10282 (N_10282,N_8642,N_8593);
xnor U10283 (N_10283,N_8320,N_8542);
and U10284 (N_10284,N_8287,N_8561);
or U10285 (N_10285,N_7613,N_8770);
xnor U10286 (N_10286,N_7549,N_7747);
and U10287 (N_10287,N_8225,N_7793);
nand U10288 (N_10288,N_7658,N_8534);
or U10289 (N_10289,N_7581,N_8276);
and U10290 (N_10290,N_8045,N_8849);
or U10291 (N_10291,N_8877,N_8658);
xnor U10292 (N_10292,N_7539,N_8116);
or U10293 (N_10293,N_8232,N_8130);
xnor U10294 (N_10294,N_8088,N_8138);
xnor U10295 (N_10295,N_8115,N_8191);
or U10296 (N_10296,N_8288,N_7683);
nor U10297 (N_10297,N_8518,N_8501);
nor U10298 (N_10298,N_7717,N_8299);
xor U10299 (N_10299,N_8388,N_7859);
xnor U10300 (N_10300,N_8852,N_7783);
or U10301 (N_10301,N_7510,N_7957);
or U10302 (N_10302,N_8300,N_7710);
or U10303 (N_10303,N_8878,N_7583);
xnor U10304 (N_10304,N_8528,N_7902);
or U10305 (N_10305,N_8346,N_8501);
and U10306 (N_10306,N_8867,N_7598);
and U10307 (N_10307,N_8716,N_8612);
and U10308 (N_10308,N_8018,N_8592);
xor U10309 (N_10309,N_7743,N_8715);
or U10310 (N_10310,N_8287,N_8302);
nand U10311 (N_10311,N_8975,N_7854);
and U10312 (N_10312,N_7649,N_7681);
and U10313 (N_10313,N_7829,N_8894);
or U10314 (N_10314,N_8853,N_8207);
nor U10315 (N_10315,N_8658,N_8273);
or U10316 (N_10316,N_7752,N_8108);
nand U10317 (N_10317,N_8188,N_8221);
or U10318 (N_10318,N_8376,N_7765);
or U10319 (N_10319,N_7993,N_8686);
nor U10320 (N_10320,N_8096,N_8255);
or U10321 (N_10321,N_8912,N_8067);
or U10322 (N_10322,N_8829,N_8059);
or U10323 (N_10323,N_8841,N_8879);
xnor U10324 (N_10324,N_8739,N_8863);
and U10325 (N_10325,N_7916,N_8659);
or U10326 (N_10326,N_7710,N_8872);
nand U10327 (N_10327,N_8676,N_8868);
nand U10328 (N_10328,N_8469,N_7523);
nand U10329 (N_10329,N_7706,N_8880);
and U10330 (N_10330,N_8999,N_8605);
xnor U10331 (N_10331,N_8922,N_8415);
xnor U10332 (N_10332,N_7697,N_8629);
nand U10333 (N_10333,N_7945,N_7782);
and U10334 (N_10334,N_8542,N_8331);
nand U10335 (N_10335,N_8774,N_8356);
and U10336 (N_10336,N_8578,N_8593);
or U10337 (N_10337,N_7647,N_8965);
xor U10338 (N_10338,N_8531,N_7865);
and U10339 (N_10339,N_8092,N_8679);
nor U10340 (N_10340,N_8046,N_7567);
nand U10341 (N_10341,N_8096,N_8891);
nor U10342 (N_10342,N_8729,N_8815);
nor U10343 (N_10343,N_7966,N_8607);
nand U10344 (N_10344,N_8369,N_7581);
nand U10345 (N_10345,N_8949,N_8904);
nand U10346 (N_10346,N_7633,N_8057);
and U10347 (N_10347,N_8586,N_8904);
nor U10348 (N_10348,N_7670,N_7553);
nand U10349 (N_10349,N_8468,N_7811);
nand U10350 (N_10350,N_7810,N_8685);
xnor U10351 (N_10351,N_7780,N_8248);
xnor U10352 (N_10352,N_7948,N_7803);
nand U10353 (N_10353,N_7503,N_7753);
and U10354 (N_10354,N_8783,N_8420);
or U10355 (N_10355,N_8138,N_8444);
or U10356 (N_10356,N_8131,N_8636);
nor U10357 (N_10357,N_8920,N_8077);
nor U10358 (N_10358,N_8331,N_8635);
nand U10359 (N_10359,N_8769,N_8001);
and U10360 (N_10360,N_8898,N_7585);
nand U10361 (N_10361,N_8451,N_8798);
and U10362 (N_10362,N_7552,N_8012);
xnor U10363 (N_10363,N_8852,N_7584);
nand U10364 (N_10364,N_7784,N_7543);
and U10365 (N_10365,N_7573,N_8527);
xnor U10366 (N_10366,N_8892,N_8234);
nor U10367 (N_10367,N_8416,N_8926);
nor U10368 (N_10368,N_8531,N_8908);
or U10369 (N_10369,N_7754,N_8540);
or U10370 (N_10370,N_8682,N_8790);
and U10371 (N_10371,N_7834,N_7850);
xor U10372 (N_10372,N_8528,N_7758);
and U10373 (N_10373,N_8098,N_8907);
nand U10374 (N_10374,N_8772,N_8007);
nand U10375 (N_10375,N_8318,N_8631);
nor U10376 (N_10376,N_8397,N_8049);
xor U10377 (N_10377,N_8894,N_8814);
and U10378 (N_10378,N_8751,N_8712);
and U10379 (N_10379,N_8838,N_8432);
or U10380 (N_10380,N_8072,N_8907);
nand U10381 (N_10381,N_8588,N_7977);
nor U10382 (N_10382,N_8755,N_8388);
or U10383 (N_10383,N_7968,N_7625);
and U10384 (N_10384,N_7877,N_8870);
xor U10385 (N_10385,N_8727,N_7739);
nand U10386 (N_10386,N_7599,N_8265);
or U10387 (N_10387,N_7934,N_8586);
or U10388 (N_10388,N_8491,N_8172);
nor U10389 (N_10389,N_8600,N_8810);
nor U10390 (N_10390,N_8022,N_8849);
and U10391 (N_10391,N_8028,N_8732);
xor U10392 (N_10392,N_8405,N_8410);
and U10393 (N_10393,N_8235,N_8822);
nand U10394 (N_10394,N_8390,N_8068);
nor U10395 (N_10395,N_8139,N_7691);
and U10396 (N_10396,N_7558,N_8264);
nand U10397 (N_10397,N_8219,N_8117);
nand U10398 (N_10398,N_8960,N_8615);
or U10399 (N_10399,N_8959,N_7907);
or U10400 (N_10400,N_7892,N_8717);
and U10401 (N_10401,N_7560,N_7907);
nor U10402 (N_10402,N_8976,N_7998);
or U10403 (N_10403,N_7722,N_8083);
nor U10404 (N_10404,N_8419,N_8364);
xor U10405 (N_10405,N_8488,N_7949);
xor U10406 (N_10406,N_7631,N_8057);
nor U10407 (N_10407,N_8301,N_7774);
and U10408 (N_10408,N_8200,N_8468);
or U10409 (N_10409,N_7580,N_7806);
nand U10410 (N_10410,N_7532,N_7704);
and U10411 (N_10411,N_8405,N_7541);
and U10412 (N_10412,N_8562,N_7890);
xnor U10413 (N_10413,N_8576,N_7640);
nor U10414 (N_10414,N_8780,N_8662);
nand U10415 (N_10415,N_8230,N_8497);
or U10416 (N_10416,N_7542,N_8648);
or U10417 (N_10417,N_8671,N_8966);
and U10418 (N_10418,N_7952,N_8682);
and U10419 (N_10419,N_7969,N_7623);
nor U10420 (N_10420,N_8961,N_8689);
and U10421 (N_10421,N_7977,N_7578);
or U10422 (N_10422,N_8889,N_7946);
or U10423 (N_10423,N_8453,N_8168);
nand U10424 (N_10424,N_8315,N_7772);
xnor U10425 (N_10425,N_8249,N_8222);
and U10426 (N_10426,N_7564,N_8004);
and U10427 (N_10427,N_8792,N_7945);
nand U10428 (N_10428,N_8039,N_8660);
nand U10429 (N_10429,N_7899,N_8824);
or U10430 (N_10430,N_8674,N_8513);
or U10431 (N_10431,N_8845,N_7847);
xor U10432 (N_10432,N_7895,N_7902);
and U10433 (N_10433,N_7692,N_7812);
nand U10434 (N_10434,N_7595,N_8394);
xnor U10435 (N_10435,N_7804,N_8035);
xor U10436 (N_10436,N_8216,N_8641);
nor U10437 (N_10437,N_8019,N_7968);
or U10438 (N_10438,N_7792,N_7740);
nand U10439 (N_10439,N_8794,N_8968);
nand U10440 (N_10440,N_7830,N_8709);
nor U10441 (N_10441,N_7641,N_7885);
or U10442 (N_10442,N_7674,N_8064);
and U10443 (N_10443,N_8947,N_7774);
nor U10444 (N_10444,N_8577,N_8051);
or U10445 (N_10445,N_8982,N_7656);
and U10446 (N_10446,N_8319,N_8951);
nand U10447 (N_10447,N_8230,N_8149);
nand U10448 (N_10448,N_7858,N_8074);
and U10449 (N_10449,N_8748,N_7581);
or U10450 (N_10450,N_8541,N_8406);
nor U10451 (N_10451,N_8738,N_8640);
and U10452 (N_10452,N_8909,N_8380);
nand U10453 (N_10453,N_8918,N_8357);
nand U10454 (N_10454,N_8729,N_8027);
nand U10455 (N_10455,N_8066,N_8269);
nor U10456 (N_10456,N_7527,N_8030);
nor U10457 (N_10457,N_7877,N_8305);
and U10458 (N_10458,N_7849,N_8305);
xnor U10459 (N_10459,N_8151,N_8873);
nor U10460 (N_10460,N_8435,N_8156);
and U10461 (N_10461,N_8791,N_8939);
or U10462 (N_10462,N_7598,N_8540);
nand U10463 (N_10463,N_7581,N_8066);
xnor U10464 (N_10464,N_7884,N_8565);
nand U10465 (N_10465,N_8470,N_7885);
nor U10466 (N_10466,N_7833,N_7711);
nand U10467 (N_10467,N_8278,N_8405);
nor U10468 (N_10468,N_8740,N_7828);
nand U10469 (N_10469,N_7926,N_8483);
nand U10470 (N_10470,N_7636,N_7878);
xnor U10471 (N_10471,N_7794,N_8520);
and U10472 (N_10472,N_8979,N_8874);
nand U10473 (N_10473,N_8461,N_8251);
and U10474 (N_10474,N_7605,N_7834);
nor U10475 (N_10475,N_8843,N_7600);
nor U10476 (N_10476,N_7690,N_7609);
or U10477 (N_10477,N_8352,N_7521);
xnor U10478 (N_10478,N_8699,N_8720);
nand U10479 (N_10479,N_8007,N_8276);
nand U10480 (N_10480,N_8635,N_8586);
or U10481 (N_10481,N_7665,N_8982);
nand U10482 (N_10482,N_8954,N_7861);
and U10483 (N_10483,N_8599,N_8743);
and U10484 (N_10484,N_8028,N_8374);
and U10485 (N_10485,N_8091,N_8754);
and U10486 (N_10486,N_7636,N_8893);
nor U10487 (N_10487,N_8224,N_7816);
nand U10488 (N_10488,N_7913,N_7857);
and U10489 (N_10489,N_8987,N_7614);
or U10490 (N_10490,N_8472,N_8567);
nand U10491 (N_10491,N_7564,N_7976);
nand U10492 (N_10492,N_7565,N_7642);
nor U10493 (N_10493,N_8603,N_8893);
nand U10494 (N_10494,N_8551,N_8668);
and U10495 (N_10495,N_8807,N_8646);
nand U10496 (N_10496,N_8190,N_8637);
and U10497 (N_10497,N_8093,N_8567);
xor U10498 (N_10498,N_8639,N_7591);
or U10499 (N_10499,N_7965,N_8432);
nor U10500 (N_10500,N_9265,N_9735);
nand U10501 (N_10501,N_9172,N_9697);
nand U10502 (N_10502,N_9853,N_9141);
nand U10503 (N_10503,N_9540,N_9405);
nor U10504 (N_10504,N_9271,N_10401);
and U10505 (N_10505,N_9279,N_9469);
nand U10506 (N_10506,N_9218,N_9794);
or U10507 (N_10507,N_9505,N_9968);
nand U10508 (N_10508,N_10149,N_9413);
nor U10509 (N_10509,N_9064,N_9013);
xor U10510 (N_10510,N_10183,N_10467);
nor U10511 (N_10511,N_9841,N_10296);
or U10512 (N_10512,N_9459,N_9401);
xor U10513 (N_10513,N_9016,N_10313);
xor U10514 (N_10514,N_10394,N_9896);
xnor U10515 (N_10515,N_9925,N_9617);
nor U10516 (N_10516,N_10103,N_10203);
and U10517 (N_10517,N_9456,N_10021);
or U10518 (N_10518,N_10282,N_9494);
and U10519 (N_10519,N_9024,N_9913);
nand U10520 (N_10520,N_10457,N_9009);
or U10521 (N_10521,N_9408,N_9254);
or U10522 (N_10522,N_9890,N_10327);
nand U10523 (N_10523,N_10381,N_9670);
xnor U10524 (N_10524,N_9879,N_10274);
and U10525 (N_10525,N_9883,N_9067);
nor U10526 (N_10526,N_9430,N_9035);
xor U10527 (N_10527,N_9870,N_9900);
nand U10528 (N_10528,N_9221,N_9875);
nand U10529 (N_10529,N_9575,N_10452);
nand U10530 (N_10530,N_9981,N_9777);
or U10531 (N_10531,N_9814,N_9287);
nand U10532 (N_10532,N_10321,N_9483);
or U10533 (N_10533,N_10148,N_9418);
and U10534 (N_10534,N_9306,N_9346);
nor U10535 (N_10535,N_9121,N_9641);
xnor U10536 (N_10536,N_10017,N_9757);
and U10537 (N_10537,N_9305,N_9344);
and U10538 (N_10538,N_10458,N_10308);
xnor U10539 (N_10539,N_9688,N_9703);
and U10540 (N_10540,N_9582,N_9257);
and U10541 (N_10541,N_9911,N_10189);
or U10542 (N_10542,N_9281,N_9343);
and U10543 (N_10543,N_10406,N_9127);
nor U10544 (N_10544,N_9770,N_9200);
xor U10545 (N_10545,N_9391,N_10291);
xor U10546 (N_10546,N_10034,N_9043);
xnor U10547 (N_10547,N_9165,N_9188);
nor U10548 (N_10548,N_10253,N_9719);
xnor U10549 (N_10549,N_9440,N_10358);
nand U10550 (N_10550,N_9213,N_9982);
or U10551 (N_10551,N_9274,N_10191);
xor U10552 (N_10552,N_9050,N_9086);
and U10553 (N_10553,N_9518,N_10319);
nor U10554 (N_10554,N_9732,N_10429);
xnor U10555 (N_10555,N_9721,N_9349);
nor U10556 (N_10556,N_10047,N_9962);
and U10557 (N_10557,N_9821,N_9302);
xor U10558 (N_10558,N_9198,N_9537);
and U10559 (N_10559,N_9155,N_9951);
nand U10560 (N_10560,N_9991,N_9810);
xor U10561 (N_10561,N_9149,N_10414);
nand U10562 (N_10562,N_9796,N_10153);
and U10563 (N_10563,N_9065,N_9194);
and U10564 (N_10564,N_10366,N_10051);
nand U10565 (N_10565,N_10426,N_9517);
and U10566 (N_10566,N_9795,N_10045);
or U10567 (N_10567,N_9601,N_9618);
xor U10568 (N_10568,N_9380,N_9292);
xor U10569 (N_10569,N_10079,N_9565);
xnor U10570 (N_10570,N_10307,N_10386);
xor U10571 (N_10571,N_9269,N_10081);
and U10572 (N_10572,N_9402,N_9362);
or U10573 (N_10573,N_10114,N_10015);
or U10574 (N_10574,N_9659,N_10065);
xnor U10575 (N_10575,N_9264,N_9579);
nand U10576 (N_10576,N_9529,N_9135);
nor U10577 (N_10577,N_10447,N_9247);
and U10578 (N_10578,N_9359,N_9376);
xor U10579 (N_10579,N_9929,N_10338);
xnor U10580 (N_10580,N_10198,N_10258);
or U10581 (N_10581,N_9410,N_9416);
nand U10582 (N_10582,N_9633,N_10354);
xnor U10583 (N_10583,N_10231,N_9476);
and U10584 (N_10584,N_10437,N_10279);
or U10585 (N_10585,N_9230,N_9316);
nand U10586 (N_10586,N_10001,N_10434);
nor U10587 (N_10587,N_9032,N_9764);
and U10588 (N_10588,N_10074,N_9867);
or U10589 (N_10589,N_9513,N_9078);
or U10590 (N_10590,N_9304,N_9425);
xnor U10591 (N_10591,N_9125,N_10295);
xnor U10592 (N_10592,N_10350,N_9710);
xnor U10593 (N_10593,N_9873,N_10263);
nand U10594 (N_10594,N_10475,N_9387);
xnor U10595 (N_10595,N_9415,N_9698);
nand U10596 (N_10596,N_10133,N_9174);
xor U10597 (N_10597,N_9115,N_9328);
xor U10598 (N_10598,N_9566,N_9436);
or U10599 (N_10599,N_10109,N_9948);
nor U10600 (N_10600,N_10388,N_9338);
nor U10601 (N_10601,N_10112,N_10091);
and U10602 (N_10602,N_10123,N_10052);
nor U10603 (N_10603,N_9379,N_9352);
nor U10604 (N_10604,N_10344,N_9630);
xnor U10605 (N_10605,N_9224,N_9222);
nor U10606 (N_10606,N_9515,N_9945);
and U10607 (N_10607,N_10325,N_10478);
or U10608 (N_10608,N_9322,N_10352);
nand U10609 (N_10609,N_9830,N_9140);
xor U10610 (N_10610,N_9453,N_9095);
nand U10611 (N_10611,N_9191,N_9649);
nor U10612 (N_10612,N_9594,N_9591);
nand U10613 (N_10613,N_9817,N_9446);
nand U10614 (N_10614,N_9278,N_10206);
xnor U10615 (N_10615,N_10069,N_9008);
xnor U10616 (N_10616,N_10407,N_10187);
xnor U10617 (N_10617,N_9826,N_10225);
xor U10618 (N_10618,N_9943,N_9286);
nand U10619 (N_10619,N_9984,N_9258);
and U10620 (N_10620,N_9743,N_10362);
nor U10621 (N_10621,N_9134,N_10041);
or U10622 (N_10622,N_9574,N_9573);
or U10623 (N_10623,N_10442,N_10353);
or U10624 (N_10624,N_10404,N_9122);
and U10625 (N_10625,N_9248,N_9809);
nand U10626 (N_10626,N_9604,N_9685);
and U10627 (N_10627,N_10010,N_10210);
and U10628 (N_10628,N_10373,N_10004);
or U10629 (N_10629,N_10300,N_10097);
and U10630 (N_10630,N_10339,N_9484);
nand U10631 (N_10631,N_10066,N_9069);
and U10632 (N_10632,N_10427,N_10056);
nand U10633 (N_10633,N_9836,N_9980);
nor U10634 (N_10634,N_9592,N_10312);
xnor U10635 (N_10635,N_9154,N_9812);
nor U10636 (N_10636,N_9746,N_10385);
or U10637 (N_10637,N_9301,N_9329);
nand U10638 (N_10638,N_9860,N_9936);
nor U10639 (N_10639,N_10193,N_9974);
or U10640 (N_10640,N_9040,N_10044);
nand U10641 (N_10641,N_9861,N_10455);
nand U10642 (N_10642,N_10374,N_9527);
nand U10643 (N_10643,N_9905,N_9458);
xnor U10644 (N_10644,N_9106,N_9838);
nor U10645 (N_10645,N_9805,N_10113);
xnor U10646 (N_10646,N_9335,N_9038);
nor U10647 (N_10647,N_9935,N_9481);
and U10648 (N_10648,N_10244,N_9912);
or U10649 (N_10649,N_9157,N_10417);
nand U10650 (N_10650,N_9827,N_9243);
nand U10651 (N_10651,N_10345,N_9152);
or U10652 (N_10652,N_10342,N_9110);
and U10653 (N_10653,N_9775,N_10042);
nor U10654 (N_10654,N_9028,N_9502);
and U10655 (N_10655,N_9276,N_9747);
nand U10656 (N_10656,N_10043,N_10317);
or U10657 (N_10657,N_10267,N_10461);
xor U10658 (N_10658,N_10039,N_9046);
nand U10659 (N_10659,N_10125,N_9855);
nand U10660 (N_10660,N_9293,N_9022);
xor U10661 (N_10661,N_10190,N_9748);
nand U10662 (N_10662,N_9741,N_9216);
and U10663 (N_10663,N_10375,N_9284);
nand U10664 (N_10664,N_9108,N_9461);
or U10665 (N_10665,N_9899,N_9037);
xor U10666 (N_10666,N_10389,N_10294);
nand U10667 (N_10667,N_9220,N_10402);
and U10668 (N_10668,N_10139,N_9350);
nand U10669 (N_10669,N_9431,N_9275);
xnor U10670 (N_10670,N_9282,N_9137);
xnor U10671 (N_10671,N_9175,N_9428);
nor U10672 (N_10672,N_10077,N_9498);
and U10673 (N_10673,N_10222,N_9311);
or U10674 (N_10674,N_10424,N_9160);
or U10675 (N_10675,N_9189,N_9300);
nand U10676 (N_10676,N_10260,N_9345);
nand U10677 (N_10677,N_9854,N_10326);
xnor U10678 (N_10678,N_9631,N_9092);
or U10679 (N_10679,N_9104,N_10235);
nor U10680 (N_10680,N_9412,N_9183);
nor U10681 (N_10681,N_10172,N_10161);
or U10682 (N_10682,N_10384,N_9435);
nand U10683 (N_10683,N_9180,N_10242);
nor U10684 (N_10684,N_10055,N_9534);
nor U10685 (N_10685,N_9307,N_9686);
or U10686 (N_10686,N_9718,N_10217);
xnor U10687 (N_10687,N_10273,N_9680);
nand U10688 (N_10688,N_9560,N_9313);
and U10689 (N_10689,N_9823,N_9298);
nand U10690 (N_10690,N_9767,N_9755);
nor U10691 (N_10691,N_10068,N_9705);
nand U10692 (N_10692,N_9950,N_10162);
nor U10693 (N_10693,N_10140,N_10158);
nor U10694 (N_10694,N_9385,N_9118);
nor U10695 (N_10695,N_9166,N_9934);
nand U10696 (N_10696,N_9876,N_9903);
nand U10697 (N_10697,N_10130,N_10151);
nand U10698 (N_10698,N_9558,N_9246);
xor U10699 (N_10699,N_10208,N_10164);
or U10700 (N_10700,N_9859,N_9760);
nor U10701 (N_10701,N_9820,N_10270);
xor U10702 (N_10702,N_9580,N_10092);
or U10703 (N_10703,N_10209,N_9319);
and U10704 (N_10704,N_9632,N_9620);
nand U10705 (N_10705,N_9370,N_9520);
nor U10706 (N_10706,N_9627,N_9672);
nor U10707 (N_10707,N_9716,N_10477);
nor U10708 (N_10708,N_9207,N_9522);
nor U10709 (N_10709,N_9400,N_10322);
or U10710 (N_10710,N_10062,N_9372);
nand U10711 (N_10711,N_10281,N_10144);
and U10712 (N_10712,N_9399,N_10119);
or U10713 (N_10713,N_9964,N_10059);
nand U10714 (N_10714,N_9897,N_10329);
xnor U10715 (N_10715,N_9671,N_9953);
xnor U10716 (N_10716,N_9355,N_10292);
nand U10717 (N_10717,N_10205,N_9506);
and U10718 (N_10718,N_10432,N_9158);
and U10719 (N_10719,N_9182,N_9126);
nand U10720 (N_10720,N_9947,N_9759);
nand U10721 (N_10721,N_9280,N_9098);
or U10722 (N_10722,N_10016,N_9708);
nand U10723 (N_10723,N_10013,N_10423);
or U10724 (N_10724,N_10498,N_9310);
or U10725 (N_10725,N_9419,N_10096);
xor U10726 (N_10726,N_10129,N_9321);
xnor U10727 (N_10727,N_10028,N_9800);
nor U10728 (N_10728,N_9363,N_9332);
nand U10729 (N_10729,N_10201,N_9331);
or U10730 (N_10730,N_9695,N_9162);
nor U10731 (N_10731,N_9614,N_10224);
nor U10732 (N_10732,N_9012,N_9051);
nor U10733 (N_10733,N_9116,N_9993);
and U10734 (N_10734,N_9482,N_9087);
xor U10735 (N_10735,N_10029,N_9524);
and U10736 (N_10736,N_9988,N_9845);
or U10737 (N_10737,N_9740,N_9366);
or U10738 (N_10738,N_9195,N_9113);
nand U10739 (N_10739,N_9569,N_9117);
and U10740 (N_10740,N_9779,N_9958);
or U10741 (N_10741,N_9930,N_10464);
xnor U10742 (N_10742,N_9815,N_9217);
nor U10743 (N_10743,N_9285,N_9295);
xor U10744 (N_10744,N_10247,N_10037);
xnor U10745 (N_10745,N_9598,N_10323);
and U10746 (N_10746,N_9957,N_9895);
nand U10747 (N_10747,N_10122,N_10080);
and U10748 (N_10748,N_10440,N_9383);
nand U10749 (N_10749,N_10473,N_9423);
xor U10750 (N_10750,N_10438,N_9798);
nor U10751 (N_10751,N_9597,N_9554);
or U10752 (N_10752,N_9365,N_9915);
xor U10753 (N_10753,N_9864,N_9268);
xor U10754 (N_10754,N_9062,N_9831);
nand U10755 (N_10755,N_9151,N_9625);
or U10756 (N_10756,N_10487,N_9025);
or U10757 (N_10757,N_9786,N_10003);
nand U10758 (N_10758,N_9309,N_10431);
nor U10759 (N_10759,N_9789,N_9645);
or U10760 (N_10760,N_9568,N_9992);
nor U10761 (N_10761,N_9877,N_10076);
nor U10762 (N_10762,N_10262,N_10484);
and U10763 (N_10763,N_9555,N_9865);
or U10764 (N_10764,N_9758,N_9595);
and U10765 (N_10765,N_9681,N_10233);
xor U10766 (N_10766,N_10428,N_9393);
nor U10767 (N_10767,N_9003,N_9496);
and U10768 (N_10768,N_10040,N_9512);
nor U10769 (N_10769,N_9082,N_10390);
xnor U10770 (N_10770,N_9939,N_10018);
or U10771 (N_10771,N_9738,N_9572);
nor U10772 (N_10772,N_10173,N_9531);
nand U10773 (N_10773,N_9563,N_10421);
xor U10774 (N_10774,N_9612,N_9130);
or U10775 (N_10775,N_9467,N_9186);
and U10776 (N_10776,N_10240,N_9253);
xnor U10777 (N_10777,N_9226,N_10476);
xor U10778 (N_10778,N_10182,N_10124);
xor U10779 (N_10779,N_9752,N_9105);
nor U10780 (N_10780,N_9168,N_9600);
nor U10781 (N_10781,N_10071,N_9602);
nor U10782 (N_10782,N_9530,N_9111);
xor U10783 (N_10783,N_10328,N_9143);
nand U10784 (N_10784,N_9414,N_9634);
xor U10785 (N_10785,N_9150,N_9843);
nand U10786 (N_10786,N_9825,N_9792);
xor U10787 (N_10787,N_10035,N_9128);
nor U10788 (N_10788,N_9214,N_9756);
nand U10789 (N_10789,N_9990,N_10286);
and U10790 (N_10790,N_9267,N_10272);
nand U10791 (N_10791,N_10171,N_10460);
nand U10792 (N_10792,N_10234,N_9369);
and U10793 (N_10793,N_10372,N_9337);
and U10794 (N_10794,N_9771,N_9209);
nand U10795 (N_10795,N_10002,N_9395);
and U10796 (N_10796,N_9424,N_9358);
or U10797 (N_10797,N_9479,N_9544);
nor U10798 (N_10798,N_10492,N_9442);
or U10799 (N_10799,N_9977,N_9159);
or U10800 (N_10800,N_9987,N_10254);
nand U10801 (N_10801,N_9657,N_10269);
or U10802 (N_10802,N_9176,N_10443);
xor U10803 (N_10803,N_9463,N_9259);
or U10804 (N_10804,N_10023,N_9869);
and U10805 (N_10805,N_9546,N_9486);
nand U10806 (N_10806,N_10365,N_9840);
nand U10807 (N_10807,N_9723,N_9891);
xor U10808 (N_10808,N_9510,N_10207);
nor U10809 (N_10809,N_9768,N_9525);
xnor U10810 (N_10810,N_10166,N_10493);
nand U10811 (N_10811,N_10073,N_10121);
and U10812 (N_10812,N_9398,N_9937);
and U10813 (N_10813,N_9054,N_9788);
or U10814 (N_10814,N_9711,N_10022);
and U10815 (N_10815,N_9171,N_9228);
nor U10816 (N_10816,N_9661,N_10499);
xor U10817 (N_10817,N_9227,N_9808);
nand U10818 (N_10818,N_9559,N_9384);
and U10819 (N_10819,N_9924,N_9689);
xor U10820 (N_10820,N_10064,N_9761);
xnor U10821 (N_10821,N_9596,N_9251);
and U10822 (N_10822,N_10318,N_9263);
nand U10823 (N_10823,N_9133,N_9577);
nor U10824 (N_10824,N_9570,N_10251);
xnor U10825 (N_10825,N_9109,N_9707);
and U10826 (N_10826,N_9644,N_9970);
xnor U10827 (N_10827,N_9717,N_10072);
or U10828 (N_10828,N_9438,N_10006);
nand U10829 (N_10829,N_9683,N_10093);
or U10830 (N_10830,N_9539,N_9403);
and U10831 (N_10831,N_10104,N_9375);
xnor U10832 (N_10832,N_9197,N_9535);
or U10833 (N_10833,N_9439,N_9033);
nor U10834 (N_10834,N_10216,N_9858);
nand U10835 (N_10835,N_10090,N_10367);
or U10836 (N_10836,N_9273,N_9377);
nor U10837 (N_10837,N_9235,N_9262);
nor U10838 (N_10838,N_10060,N_9781);
or U10839 (N_10839,N_10186,N_10194);
xnor U10840 (N_10840,N_9093,N_9324);
nand U10841 (N_10841,N_9392,N_10131);
nand U10842 (N_10842,N_9107,N_9099);
or U10843 (N_10843,N_9312,N_10061);
nand U10844 (N_10844,N_9536,N_9356);
nor U10845 (N_10845,N_9881,N_9629);
xnor U10846 (N_10846,N_10058,N_9720);
nor U10847 (N_10847,N_9842,N_9927);
and U10848 (N_10848,N_10252,N_9932);
nor U10849 (N_10849,N_10157,N_9029);
or U10850 (N_10850,N_9581,N_10310);
or U10851 (N_10851,N_9824,N_10361);
nand U10852 (N_10852,N_9908,N_9204);
or U10853 (N_10853,N_9206,N_10287);
and U10854 (N_10854,N_9411,N_10398);
and U10855 (N_10855,N_9240,N_10368);
or U10856 (N_10856,N_9804,N_9255);
and U10857 (N_10857,N_9849,N_9452);
nor U10858 (N_10858,N_9007,N_9561);
and U10859 (N_10859,N_9822,N_9916);
and U10860 (N_10860,N_10330,N_10168);
and U10861 (N_10861,N_9341,N_9079);
nor U10862 (N_10862,N_9521,N_9852);
nand U10863 (N_10863,N_9998,N_9739);
or U10864 (N_10864,N_9910,N_9640);
nand U10865 (N_10865,N_9089,N_9734);
and U10866 (N_10866,N_9289,N_9211);
nor U10867 (N_10867,N_9123,N_10453);
or U10868 (N_10868,N_9210,N_9138);
xor U10869 (N_10869,N_9762,N_9851);
nand U10870 (N_10870,N_9669,N_9325);
and U10871 (N_10871,N_9704,N_10446);
or U10872 (N_10872,N_9066,N_9499);
xor U10873 (N_10873,N_10070,N_10057);
xnor U10874 (N_10874,N_10019,N_9421);
or U10875 (N_10875,N_9959,N_10048);
nor U10876 (N_10876,N_9085,N_10202);
nor U10877 (N_10877,N_9074,N_10177);
nand U10878 (N_10878,N_10356,N_10215);
and U10879 (N_10879,N_9557,N_10142);
xnor U10880 (N_10880,N_9509,N_9696);
nand U10881 (N_10881,N_9485,N_10471);
nand U10882 (N_10882,N_9797,N_9765);
nand U10883 (N_10883,N_9238,N_9966);
nand U10884 (N_10884,N_9793,N_9407);
and U10885 (N_10885,N_9058,N_10200);
and U10886 (N_10886,N_10221,N_9063);
xor U10887 (N_10887,N_9010,N_10435);
or U10888 (N_10888,N_9893,N_9941);
or U10889 (N_10889,N_10433,N_10419);
xor U10890 (N_10890,N_10441,N_9241);
or U10891 (N_10891,N_9989,N_9381);
nand U10892 (N_10892,N_10204,N_9653);
xnor U10893 (N_10893,N_9516,N_10430);
nor U10894 (N_10894,N_9702,N_9769);
or U10895 (N_10895,N_10462,N_9406);
or U10896 (N_10896,N_10246,N_9196);
or U10897 (N_10897,N_10243,N_9480);
nand U10898 (N_10898,N_9684,N_9100);
and U10899 (N_10899,N_9173,N_10400);
or U10900 (N_10900,N_10335,N_9744);
and U10901 (N_10901,N_9260,N_9208);
and U10902 (N_10902,N_10181,N_9909);
nor U10903 (N_10903,N_9234,N_10049);
or U10904 (N_10904,N_9886,N_10012);
nand U10905 (N_10905,N_9465,N_10110);
or U10906 (N_10906,N_9503,N_9219);
nand U10907 (N_10907,N_10275,N_9889);
nor U10908 (N_10908,N_9039,N_10214);
nand U10909 (N_10909,N_9652,N_10152);
nor U10910 (N_10910,N_10343,N_9148);
or U10911 (N_10911,N_10036,N_9715);
xor U10912 (N_10912,N_10314,N_9474);
or U10913 (N_10913,N_10232,N_10094);
nand U10914 (N_10914,N_9700,N_10351);
xnor U10915 (N_10915,N_10087,N_9933);
and U10916 (N_10916,N_9621,N_9120);
or U10917 (N_10917,N_9663,N_9420);
or U10918 (N_10918,N_9464,N_9250);
and U10919 (N_10919,N_9662,N_10132);
nor U10920 (N_10920,N_9139,N_10155);
or U10921 (N_10921,N_9541,N_9807);
xnor U10922 (N_10922,N_10086,N_9894);
nand U10923 (N_10923,N_9832,N_10369);
or U10924 (N_10924,N_9315,N_10285);
xor U10925 (N_10925,N_9547,N_9986);
nand U10926 (N_10926,N_9564,N_10305);
xor U10927 (N_10927,N_10211,N_9187);
or U10928 (N_10928,N_9511,N_9952);
nor U10929 (N_10929,N_9972,N_10415);
nand U10930 (N_10930,N_9588,N_9960);
xnor U10931 (N_10931,N_9205,N_9487);
nand U10932 (N_10932,N_9094,N_9587);
nand U10933 (N_10933,N_9448,N_9971);
or U10934 (N_10934,N_10000,N_9979);
or U10935 (N_10935,N_10409,N_9144);
or U10936 (N_10936,N_10212,N_9665);
or U10937 (N_10937,N_9996,N_9203);
xnor U10938 (N_10938,N_9283,N_10309);
nand U10939 (N_10939,N_9553,N_10280);
nand U10940 (N_10940,N_9156,N_10485);
or U10941 (N_10941,N_9586,N_9178);
and U10942 (N_10942,N_9942,N_10337);
nand U10943 (N_10943,N_10357,N_10259);
and U10944 (N_10944,N_9837,N_9327);
or U10945 (N_10945,N_9725,N_9863);
xnor U10946 (N_10946,N_9682,N_9584);
nor U10947 (N_10947,N_9455,N_9426);
nor U10948 (N_10948,N_9919,N_10289);
or U10949 (N_10949,N_10333,N_9468);
or U10950 (N_10950,N_9272,N_10392);
and U10951 (N_10951,N_9846,N_10320);
nand U10952 (N_10952,N_9928,N_9611);
and U10953 (N_10953,N_9847,N_9164);
nand U10954 (N_10954,N_9556,N_9101);
and U10955 (N_10955,N_10245,N_10391);
xnor U10956 (N_10956,N_9607,N_9599);
and U10957 (N_10957,N_9277,N_9585);
nor U10958 (N_10958,N_9296,N_9623);
and U10959 (N_10959,N_10449,N_9252);
or U10960 (N_10960,N_9396,N_9887);
nand U10961 (N_10961,N_9776,N_9288);
nor U10962 (N_10962,N_10380,N_10085);
and U10963 (N_10963,N_9462,N_9031);
nand U10964 (N_10964,N_10118,N_9005);
xnor U10965 (N_10965,N_9857,N_10377);
xnor U10966 (N_10966,N_9351,N_10228);
or U10967 (N_10967,N_9097,N_10180);
or U10968 (N_10968,N_10256,N_9583);
or U10969 (N_10969,N_9457,N_9334);
xor U10970 (N_10970,N_10469,N_10027);
nand U10971 (N_10971,N_10347,N_10025);
or U10972 (N_10972,N_9081,N_9199);
nand U10973 (N_10973,N_9048,N_10436);
or U10974 (N_10974,N_10032,N_9112);
xor U10975 (N_10975,N_9034,N_10276);
xnor U10976 (N_10976,N_9878,N_9364);
nor U10977 (N_10977,N_10218,N_9353);
or U10978 (N_10978,N_9027,N_9567);
and U10979 (N_10979,N_9729,N_9961);
nor U10980 (N_10980,N_9643,N_9997);
nand U10981 (N_10981,N_9488,N_9639);
nor U10982 (N_10982,N_9361,N_9080);
or U10983 (N_10983,N_10128,N_10174);
or U10984 (N_10984,N_10226,N_9922);
and U10985 (N_10985,N_9880,N_10306);
nor U10986 (N_10986,N_10179,N_9437);
nand U10987 (N_10987,N_9654,N_10156);
nand U10988 (N_10988,N_10283,N_10364);
nor U10989 (N_10989,N_10084,N_9340);
nand U10990 (N_10990,N_9026,N_9811);
and U10991 (N_10991,N_10116,N_9994);
nor U10992 (N_10992,N_9828,N_9806);
xor U10993 (N_10993,N_9545,N_10489);
and U10994 (N_10994,N_9619,N_9742);
xor U10995 (N_10995,N_9637,N_10230);
and U10996 (N_10996,N_10020,N_9898);
and U10997 (N_10997,N_9850,N_9103);
nor U10998 (N_10998,N_10150,N_10236);
xor U10999 (N_10999,N_9626,N_9507);
and U11000 (N_11000,N_9733,N_9006);
or U11001 (N_11001,N_10451,N_9354);
or U11002 (N_11002,N_9023,N_9871);
or U11003 (N_11003,N_9675,N_9433);
nor U11004 (N_11004,N_10147,N_9646);
nor U11005 (N_11005,N_9589,N_10298);
nor U11006 (N_11006,N_10399,N_9904);
and U11007 (N_11007,N_10418,N_9018);
or U11008 (N_11008,N_9699,N_10106);
nor U11009 (N_11009,N_10229,N_10411);
nor U11010 (N_11010,N_10220,N_9750);
nor U11011 (N_11011,N_9677,N_9215);
and U11012 (N_11012,N_9914,N_10468);
nand U11013 (N_11013,N_10188,N_10376);
or U11014 (N_11014,N_9374,N_9429);
nor U11015 (N_11015,N_9330,N_9232);
and U11016 (N_11016,N_10038,N_10175);
nand U11017 (N_11017,N_9642,N_9136);
nand U11018 (N_11018,N_10494,N_9651);
and U11019 (N_11019,N_9212,N_9514);
nor U11020 (N_11020,N_10141,N_9417);
or U11021 (N_11021,N_10278,N_9833);
and U11022 (N_11022,N_9318,N_9070);
nand U11023 (N_11023,N_9042,N_9475);
xnor U11024 (N_11024,N_9441,N_9347);
and U11025 (N_11025,N_10102,N_9976);
or U11026 (N_11026,N_9477,N_10336);
nor U11027 (N_11027,N_9057,N_9713);
or U11028 (N_11028,N_9073,N_9443);
nand U11029 (N_11029,N_10223,N_9147);
and U11030 (N_11030,N_9709,N_10459);
or U11031 (N_11031,N_9975,N_10227);
xnor U11032 (N_11032,N_9844,N_9021);
or U11033 (N_11033,N_9049,N_9790);
nand U11034 (N_11034,N_10349,N_9386);
and U11035 (N_11035,N_9114,N_9382);
xor U11036 (N_11036,N_9676,N_9142);
or U11037 (N_11037,N_10138,N_10495);
or U11038 (N_11038,N_10135,N_9550);
or U11039 (N_11039,N_10334,N_10111);
and U11040 (N_11040,N_9799,N_9882);
or U11041 (N_11041,N_9648,N_9427);
nor U11042 (N_11042,N_10444,N_9470);
nor U11043 (N_11043,N_9730,N_9868);
xnor U11044 (N_11044,N_9606,N_9161);
or U11045 (N_11045,N_10143,N_9466);
xor U11046 (N_11046,N_9169,N_9145);
and U11047 (N_11047,N_10371,N_9233);
or U11048 (N_11048,N_9508,N_10160);
xor U11049 (N_11049,N_9985,N_9552);
or U11050 (N_11050,N_9236,N_10359);
nor U11051 (N_11051,N_10063,N_9060);
nor U11052 (N_11052,N_9674,N_9290);
xor U11053 (N_11053,N_10466,N_10098);
or U11054 (N_11054,N_9727,N_9803);
nand U11055 (N_11055,N_9874,N_10410);
xor U11056 (N_11056,N_10331,N_10005);
xor U11057 (N_11057,N_9266,N_10030);
or U11058 (N_11058,N_10115,N_9917);
xnor U11059 (N_11059,N_9059,N_9132);
and U11060 (N_11060,N_10363,N_9004);
or U11061 (N_11061,N_9249,N_9170);
nor U11062 (N_11062,N_9963,N_10403);
nand U11063 (N_11063,N_9862,N_10184);
nand U11064 (N_11064,N_10192,N_10324);
or U11065 (N_11065,N_9002,N_9237);
xnor U11066 (N_11066,N_9726,N_10483);
nand U11067 (N_11067,N_9177,N_10117);
nor U11068 (N_11068,N_10382,N_10340);
xor U11069 (N_11069,N_9839,N_9445);
xnor U11070 (N_11070,N_9872,N_9519);
and U11071 (N_11071,N_9816,N_9967);
or U11072 (N_11072,N_9562,N_9819);
nand U11073 (N_11073,N_9088,N_9679);
nand U11074 (N_11074,N_9014,N_9036);
nand U11075 (N_11075,N_10031,N_9017);
or U11076 (N_11076,N_10379,N_10439);
nor U11077 (N_11077,N_9239,N_10332);
or U11078 (N_11078,N_9076,N_10082);
xor U11079 (N_11079,N_9668,N_9472);
or U11080 (N_11080,N_9749,N_9636);
or U11081 (N_11081,N_10265,N_9954);
or U11082 (N_11082,N_9202,N_10304);
or U11083 (N_11083,N_10213,N_9432);
and U11084 (N_11084,N_9052,N_9270);
nor U11085 (N_11085,N_9694,N_10100);
and U11086 (N_11086,N_10241,N_10299);
or U11087 (N_11087,N_9528,N_9444);
nor U11088 (N_11088,N_9818,N_10136);
xor U11089 (N_11089,N_9763,N_10293);
nor U11090 (N_11090,N_10033,N_9691);
xor U11091 (N_11091,N_9451,N_9965);
nand U11092 (N_11092,N_9722,N_10303);
or U11093 (N_11093,N_10450,N_9478);
xor U11094 (N_11094,N_10355,N_9231);
nor U11095 (N_11095,N_9084,N_9163);
xnor U11096 (N_11096,N_10348,N_10405);
or U11097 (N_11097,N_9001,N_10395);
or U11098 (N_11098,N_10120,N_10266);
and U11099 (N_11099,N_9542,N_9501);
and U11100 (N_11100,N_10008,N_9973);
nand U11101 (N_11101,N_10238,N_9902);
xnor U11102 (N_11102,N_9603,N_10250);
nor U11103 (N_11103,N_9242,N_9667);
or U11104 (N_11104,N_9551,N_9693);
xnor U11105 (N_11105,N_10456,N_10316);
or U11106 (N_11106,N_9782,N_10099);
nor U11107 (N_11107,N_10146,N_9728);
xor U11108 (N_11108,N_9075,N_10249);
nor U11109 (N_11109,N_10195,N_9124);
and U11110 (N_11110,N_10346,N_9339);
nor U11111 (N_11111,N_10383,N_9090);
nand U11112 (N_11112,N_10261,N_9778);
xor U11113 (N_11113,N_10075,N_9787);
and U11114 (N_11114,N_9373,N_9785);
nor U11115 (N_11115,N_9673,N_9449);
and U11116 (N_11116,N_9613,N_9737);
nor U11117 (N_11117,N_9549,N_9129);
nand U11118 (N_11118,N_9856,N_10054);
xnor U11119 (N_11119,N_9179,N_9802);
nor U11120 (N_11120,N_9303,N_9225);
and U11121 (N_11121,N_9348,N_9342);
xnor U11122 (N_11122,N_9692,N_9724);
nor U11123 (N_11123,N_10154,N_9834);
and U11124 (N_11124,N_9576,N_10176);
nor U11125 (N_11125,N_10089,N_9714);
or U11126 (N_11126,N_9772,N_9801);
or U11127 (N_11127,N_10178,N_10024);
nor U11128 (N_11128,N_9367,N_9690);
xor U11129 (N_11129,N_10271,N_9297);
or U11130 (N_11130,N_9624,N_9314);
or U11131 (N_11131,N_9096,N_9884);
nor U11132 (N_11132,N_9615,N_10078);
nand U11133 (N_11133,N_10496,N_10067);
nand U11134 (N_11134,N_10445,N_10378);
nand U11135 (N_11135,N_9999,N_10416);
or U11136 (N_11136,N_9783,N_10101);
nor U11137 (N_11137,N_9185,N_9192);
and U11138 (N_11138,N_10408,N_9532);
or U11139 (N_11139,N_9647,N_10185);
and U11140 (N_11140,N_10126,N_9969);
nand U11141 (N_11141,N_9923,N_9394);
nand U11142 (N_11142,N_9946,N_9533);
and U11143 (N_11143,N_10393,N_9921);
xor U11144 (N_11144,N_10219,N_10341);
and U11145 (N_11145,N_9523,N_10083);
or U11146 (N_11146,N_9491,N_9578);
or U11147 (N_11147,N_9000,N_9745);
or U11148 (N_11148,N_9995,N_9678);
nand U11149 (N_11149,N_9434,N_10053);
xor U11150 (N_11150,N_9299,N_9020);
nor U11151 (N_11151,N_9072,N_10277);
nand U11152 (N_11152,N_10007,N_9885);
nand U11153 (N_11153,N_10479,N_10046);
nor U11154 (N_11154,N_10095,N_10422);
or U11155 (N_11155,N_9944,N_10257);
or U11156 (N_11156,N_9320,N_10009);
xnor U11157 (N_11157,N_10448,N_9460);
or U11158 (N_11158,N_9791,N_9256);
and U11159 (N_11159,N_9835,N_9153);
and U11160 (N_11160,N_9083,N_9077);
nand U11161 (N_11161,N_9616,N_10167);
or U11162 (N_11162,N_9422,N_9829);
nand U11163 (N_11163,N_9390,N_9931);
xnor U11164 (N_11164,N_9404,N_9495);
nand U11165 (N_11165,N_9223,N_10465);
and U11166 (N_11166,N_10387,N_9047);
xor U11167 (N_11167,N_9548,N_9201);
xor U11168 (N_11168,N_9368,N_10412);
or U11169 (N_11169,N_10288,N_9706);
or U11170 (N_11170,N_9492,N_9041);
nor U11171 (N_11171,N_9053,N_9650);
nand U11172 (N_11172,N_9888,N_9091);
nand U11173 (N_11173,N_10137,N_9901);
or U11174 (N_11174,N_9543,N_9055);
or U11175 (N_11175,N_9773,N_10425);
nand U11176 (N_11176,N_10360,N_10026);
xnor U11177 (N_11177,N_9056,N_10397);
and U11178 (N_11178,N_9751,N_9609);
xor U11179 (N_11179,N_9938,N_9473);
nor U11180 (N_11180,N_9493,N_9918);
and U11181 (N_11181,N_10284,N_10134);
and U11182 (N_11182,N_9622,N_9848);
xnor U11183 (N_11183,N_9590,N_9190);
nand U11184 (N_11184,N_10197,N_10268);
or U11185 (N_11185,N_9409,N_10497);
xor U11186 (N_11186,N_9712,N_9538);
and U11187 (N_11187,N_10302,N_9471);
xnor U11188 (N_11188,N_10088,N_9317);
or U11189 (N_11189,N_9605,N_9774);
and U11190 (N_11190,N_10491,N_10315);
nand U11191 (N_11191,N_10165,N_10014);
or U11192 (N_11192,N_9181,N_9011);
and U11193 (N_11193,N_9628,N_10011);
and U11194 (N_11194,N_9571,N_9244);
nor U11195 (N_11195,N_10199,N_9019);
nor U11196 (N_11196,N_10481,N_10050);
nand U11197 (N_11197,N_9489,N_9378);
or U11198 (N_11198,N_10127,N_9955);
nand U11199 (N_11199,N_9593,N_10108);
nand U11200 (N_11200,N_10301,N_9956);
or U11201 (N_11201,N_9608,N_10255);
nor U11202 (N_11202,N_9371,N_9736);
or U11203 (N_11203,N_10482,N_10170);
and U11204 (N_11204,N_10237,N_9184);
and U11205 (N_11205,N_9068,N_9920);
nor U11206 (N_11206,N_9389,N_10420);
and U11207 (N_11207,N_10488,N_9926);
xnor U11208 (N_11208,N_9638,N_10159);
nand U11209 (N_11209,N_9907,N_10490);
nand U11210 (N_11210,N_9635,N_9892);
or U11211 (N_11211,N_9655,N_9813);
nand U11212 (N_11212,N_9866,N_9753);
nand U11213 (N_11213,N_9660,N_10196);
xor U11214 (N_11214,N_9701,N_10470);
xor U11215 (N_11215,N_9308,N_10297);
nand U11216 (N_11216,N_9261,N_9526);
and U11217 (N_11217,N_9447,N_9336);
nor U11218 (N_11218,N_9978,N_9397);
xor U11219 (N_11219,N_9497,N_9454);
xnor U11220 (N_11220,N_10413,N_9780);
xnor U11221 (N_11221,N_10480,N_9071);
xnor U11222 (N_11222,N_10264,N_9687);
and U11223 (N_11223,N_9146,N_10474);
or U11224 (N_11224,N_9193,N_10145);
nor U11225 (N_11225,N_9500,N_9504);
xnor U11226 (N_11226,N_9490,N_10107);
or U11227 (N_11227,N_9245,N_10454);
nand U11228 (N_11228,N_9229,N_10472);
nand U11229 (N_11229,N_9983,N_9291);
and U11230 (N_11230,N_9333,N_9940);
or U11231 (N_11231,N_9323,N_9045);
or U11232 (N_11232,N_9610,N_9044);
xor U11233 (N_11233,N_9731,N_9015);
nor U11234 (N_11234,N_10163,N_9784);
or U11235 (N_11235,N_10311,N_9666);
xor U11236 (N_11236,N_9754,N_9388);
or U11237 (N_11237,N_10486,N_9664);
or U11238 (N_11238,N_9658,N_10396);
xnor U11239 (N_11239,N_9766,N_10370);
nor U11240 (N_11240,N_10169,N_9102);
xor U11241 (N_11241,N_9030,N_9906);
nor U11242 (N_11242,N_9119,N_9131);
xnor U11243 (N_11243,N_9656,N_10290);
nor U11244 (N_11244,N_9949,N_10239);
or U11245 (N_11245,N_10248,N_9450);
nor U11246 (N_11246,N_9360,N_10463);
nand U11247 (N_11247,N_9326,N_9294);
and U11248 (N_11248,N_10105,N_9167);
nor U11249 (N_11249,N_9061,N_9357);
or U11250 (N_11250,N_10403,N_9347);
and U11251 (N_11251,N_10355,N_10118);
nor U11252 (N_11252,N_10251,N_9145);
xor U11253 (N_11253,N_10059,N_10340);
xor U11254 (N_11254,N_9660,N_9935);
nand U11255 (N_11255,N_9144,N_9401);
xor U11256 (N_11256,N_10476,N_10445);
nor U11257 (N_11257,N_9999,N_10446);
nor U11258 (N_11258,N_9780,N_9257);
nor U11259 (N_11259,N_9154,N_9650);
nand U11260 (N_11260,N_10335,N_9850);
xor U11261 (N_11261,N_9164,N_9061);
nor U11262 (N_11262,N_9856,N_10271);
and U11263 (N_11263,N_9701,N_9984);
and U11264 (N_11264,N_9260,N_10084);
nand U11265 (N_11265,N_9520,N_9432);
nor U11266 (N_11266,N_9926,N_9475);
nand U11267 (N_11267,N_10096,N_10494);
and U11268 (N_11268,N_9954,N_9429);
or U11269 (N_11269,N_9316,N_9608);
nand U11270 (N_11270,N_9327,N_9399);
nand U11271 (N_11271,N_10386,N_9994);
xor U11272 (N_11272,N_9941,N_9092);
and U11273 (N_11273,N_10158,N_9659);
nor U11274 (N_11274,N_9304,N_9269);
or U11275 (N_11275,N_9010,N_9659);
nand U11276 (N_11276,N_9858,N_9599);
xnor U11277 (N_11277,N_10098,N_9630);
xnor U11278 (N_11278,N_9300,N_9109);
or U11279 (N_11279,N_9941,N_9651);
or U11280 (N_11280,N_10450,N_9111);
nor U11281 (N_11281,N_9916,N_9776);
and U11282 (N_11282,N_10093,N_9017);
and U11283 (N_11283,N_9468,N_9774);
or U11284 (N_11284,N_9143,N_9831);
xor U11285 (N_11285,N_10210,N_9303);
nand U11286 (N_11286,N_9266,N_9158);
nand U11287 (N_11287,N_10467,N_9237);
or U11288 (N_11288,N_9333,N_9570);
nor U11289 (N_11289,N_9693,N_9665);
nand U11290 (N_11290,N_9779,N_9099);
nand U11291 (N_11291,N_9987,N_10393);
and U11292 (N_11292,N_9842,N_9682);
xnor U11293 (N_11293,N_9763,N_10299);
or U11294 (N_11294,N_9839,N_10339);
xor U11295 (N_11295,N_9433,N_9597);
nand U11296 (N_11296,N_10224,N_10312);
nand U11297 (N_11297,N_9884,N_10310);
nor U11298 (N_11298,N_10422,N_10447);
and U11299 (N_11299,N_10468,N_10077);
and U11300 (N_11300,N_10026,N_10284);
and U11301 (N_11301,N_9257,N_9812);
and U11302 (N_11302,N_9561,N_9591);
and U11303 (N_11303,N_10346,N_10120);
and U11304 (N_11304,N_10013,N_9106);
nand U11305 (N_11305,N_10304,N_10142);
nor U11306 (N_11306,N_9548,N_9419);
nand U11307 (N_11307,N_9991,N_9921);
or U11308 (N_11308,N_9455,N_9201);
or U11309 (N_11309,N_9726,N_10358);
nand U11310 (N_11310,N_9000,N_9853);
or U11311 (N_11311,N_10097,N_9693);
xor U11312 (N_11312,N_10364,N_9456);
nand U11313 (N_11313,N_10495,N_9203);
or U11314 (N_11314,N_9266,N_9606);
xnor U11315 (N_11315,N_9158,N_10373);
nor U11316 (N_11316,N_10179,N_9732);
nand U11317 (N_11317,N_9278,N_9413);
xnor U11318 (N_11318,N_9962,N_9572);
or U11319 (N_11319,N_9953,N_10023);
nand U11320 (N_11320,N_10354,N_9277);
or U11321 (N_11321,N_9584,N_9799);
xor U11322 (N_11322,N_10113,N_9730);
nor U11323 (N_11323,N_9674,N_10280);
and U11324 (N_11324,N_9557,N_10037);
or U11325 (N_11325,N_9570,N_9761);
and U11326 (N_11326,N_9711,N_9480);
or U11327 (N_11327,N_9245,N_9640);
nand U11328 (N_11328,N_9793,N_10036);
nand U11329 (N_11329,N_10243,N_10365);
and U11330 (N_11330,N_9618,N_9342);
or U11331 (N_11331,N_9764,N_9976);
nand U11332 (N_11332,N_9763,N_9090);
or U11333 (N_11333,N_9427,N_9528);
and U11334 (N_11334,N_10433,N_9797);
xnor U11335 (N_11335,N_9328,N_9760);
nor U11336 (N_11336,N_9971,N_10245);
xnor U11337 (N_11337,N_10225,N_9978);
nor U11338 (N_11338,N_10085,N_10411);
nor U11339 (N_11339,N_9304,N_9511);
or U11340 (N_11340,N_9702,N_10056);
or U11341 (N_11341,N_9420,N_9697);
or U11342 (N_11342,N_10384,N_10278);
xor U11343 (N_11343,N_10161,N_9807);
nor U11344 (N_11344,N_9630,N_9879);
or U11345 (N_11345,N_9148,N_10313);
nand U11346 (N_11346,N_10159,N_10296);
xnor U11347 (N_11347,N_9476,N_9454);
xnor U11348 (N_11348,N_9981,N_10014);
or U11349 (N_11349,N_10052,N_9425);
and U11350 (N_11350,N_9638,N_9100);
nor U11351 (N_11351,N_9601,N_9704);
nand U11352 (N_11352,N_9687,N_9584);
and U11353 (N_11353,N_9850,N_9610);
nand U11354 (N_11354,N_9804,N_9954);
and U11355 (N_11355,N_10164,N_10182);
nand U11356 (N_11356,N_9925,N_9240);
nor U11357 (N_11357,N_9536,N_9955);
xnor U11358 (N_11358,N_9490,N_10119);
nand U11359 (N_11359,N_9576,N_10461);
and U11360 (N_11360,N_9530,N_10446);
nor U11361 (N_11361,N_9096,N_9082);
nand U11362 (N_11362,N_9894,N_9785);
and U11363 (N_11363,N_9129,N_10056);
xnor U11364 (N_11364,N_10435,N_9354);
xor U11365 (N_11365,N_9816,N_9203);
nor U11366 (N_11366,N_9789,N_9021);
or U11367 (N_11367,N_9097,N_10069);
nor U11368 (N_11368,N_9156,N_9248);
xor U11369 (N_11369,N_9087,N_9440);
xor U11370 (N_11370,N_10456,N_10421);
or U11371 (N_11371,N_9080,N_10290);
and U11372 (N_11372,N_9994,N_9729);
xor U11373 (N_11373,N_9696,N_9058);
or U11374 (N_11374,N_9396,N_9744);
or U11375 (N_11375,N_10483,N_10475);
xnor U11376 (N_11376,N_10091,N_9935);
nand U11377 (N_11377,N_9345,N_9950);
and U11378 (N_11378,N_9789,N_9653);
xnor U11379 (N_11379,N_9398,N_9926);
and U11380 (N_11380,N_9708,N_9002);
nor U11381 (N_11381,N_10319,N_9618);
nor U11382 (N_11382,N_9713,N_10190);
xnor U11383 (N_11383,N_9672,N_9874);
xnor U11384 (N_11384,N_10014,N_10101);
or U11385 (N_11385,N_10414,N_9030);
and U11386 (N_11386,N_9747,N_9756);
nor U11387 (N_11387,N_10084,N_9589);
nor U11388 (N_11388,N_10096,N_9649);
nor U11389 (N_11389,N_10023,N_10251);
nand U11390 (N_11390,N_10427,N_10086);
and U11391 (N_11391,N_9081,N_10356);
or U11392 (N_11392,N_9029,N_10214);
nor U11393 (N_11393,N_9732,N_10320);
and U11394 (N_11394,N_10299,N_9708);
nand U11395 (N_11395,N_9281,N_10039);
xor U11396 (N_11396,N_9658,N_10145);
nand U11397 (N_11397,N_9654,N_10333);
nand U11398 (N_11398,N_9515,N_9453);
and U11399 (N_11399,N_9276,N_9119);
and U11400 (N_11400,N_9695,N_9870);
nand U11401 (N_11401,N_9974,N_9507);
or U11402 (N_11402,N_10499,N_10052);
and U11403 (N_11403,N_10055,N_9280);
nor U11404 (N_11404,N_9638,N_10477);
nand U11405 (N_11405,N_9586,N_10449);
and U11406 (N_11406,N_9356,N_9892);
or U11407 (N_11407,N_10498,N_9192);
xnor U11408 (N_11408,N_9891,N_10265);
and U11409 (N_11409,N_9900,N_9474);
nand U11410 (N_11410,N_9359,N_9370);
nand U11411 (N_11411,N_10421,N_10199);
and U11412 (N_11412,N_9464,N_9902);
nor U11413 (N_11413,N_9411,N_9390);
nor U11414 (N_11414,N_9691,N_9994);
or U11415 (N_11415,N_9650,N_9638);
nor U11416 (N_11416,N_10312,N_9223);
nor U11417 (N_11417,N_9643,N_9844);
nor U11418 (N_11418,N_10007,N_9344);
nor U11419 (N_11419,N_9779,N_9074);
xor U11420 (N_11420,N_10289,N_9992);
xnor U11421 (N_11421,N_9457,N_10462);
xnor U11422 (N_11422,N_9954,N_10462);
xnor U11423 (N_11423,N_10090,N_9181);
or U11424 (N_11424,N_9581,N_10219);
xnor U11425 (N_11425,N_9341,N_9744);
xnor U11426 (N_11426,N_9873,N_9911);
xnor U11427 (N_11427,N_10073,N_10307);
and U11428 (N_11428,N_9070,N_9390);
or U11429 (N_11429,N_9566,N_9739);
and U11430 (N_11430,N_9312,N_10222);
or U11431 (N_11431,N_9419,N_9708);
xnor U11432 (N_11432,N_9491,N_9854);
and U11433 (N_11433,N_9988,N_9528);
xnor U11434 (N_11434,N_9567,N_9285);
nor U11435 (N_11435,N_10026,N_9182);
nand U11436 (N_11436,N_9107,N_10471);
xor U11437 (N_11437,N_9585,N_10363);
xor U11438 (N_11438,N_9539,N_9184);
and U11439 (N_11439,N_9671,N_9906);
nor U11440 (N_11440,N_9388,N_10360);
nor U11441 (N_11441,N_10322,N_10372);
xnor U11442 (N_11442,N_10391,N_9064);
nand U11443 (N_11443,N_10258,N_9581);
or U11444 (N_11444,N_10156,N_9863);
nand U11445 (N_11445,N_10290,N_9365);
and U11446 (N_11446,N_9062,N_9371);
nor U11447 (N_11447,N_10424,N_9706);
nor U11448 (N_11448,N_9883,N_10031);
xnor U11449 (N_11449,N_9408,N_10084);
or U11450 (N_11450,N_10187,N_10133);
or U11451 (N_11451,N_9905,N_9239);
nor U11452 (N_11452,N_9343,N_9183);
and U11453 (N_11453,N_9055,N_10296);
xnor U11454 (N_11454,N_10436,N_9255);
nor U11455 (N_11455,N_9773,N_9541);
or U11456 (N_11456,N_9368,N_9330);
xor U11457 (N_11457,N_9371,N_9679);
or U11458 (N_11458,N_9225,N_10358);
nand U11459 (N_11459,N_9499,N_9372);
and U11460 (N_11460,N_10281,N_10087);
xor U11461 (N_11461,N_9258,N_9248);
xnor U11462 (N_11462,N_9328,N_10145);
xnor U11463 (N_11463,N_9347,N_10228);
nor U11464 (N_11464,N_9029,N_9172);
xnor U11465 (N_11465,N_9213,N_10267);
nand U11466 (N_11466,N_9656,N_10131);
and U11467 (N_11467,N_9236,N_10033);
nor U11468 (N_11468,N_9163,N_9849);
and U11469 (N_11469,N_9079,N_9821);
or U11470 (N_11470,N_9402,N_10363);
or U11471 (N_11471,N_9370,N_9092);
nor U11472 (N_11472,N_10103,N_9005);
nand U11473 (N_11473,N_10295,N_9485);
or U11474 (N_11474,N_9520,N_9871);
nor U11475 (N_11475,N_10237,N_9655);
or U11476 (N_11476,N_10044,N_9704);
nand U11477 (N_11477,N_10401,N_9546);
nor U11478 (N_11478,N_9762,N_10421);
nand U11479 (N_11479,N_9111,N_9712);
nor U11480 (N_11480,N_10120,N_10151);
xnor U11481 (N_11481,N_9748,N_9476);
nor U11482 (N_11482,N_9847,N_9350);
or U11483 (N_11483,N_9390,N_10154);
nor U11484 (N_11484,N_9273,N_10394);
xor U11485 (N_11485,N_9059,N_9573);
nor U11486 (N_11486,N_10044,N_10278);
nor U11487 (N_11487,N_9649,N_9316);
xnor U11488 (N_11488,N_9183,N_10073);
or U11489 (N_11489,N_9718,N_9455);
or U11490 (N_11490,N_9531,N_9937);
and U11491 (N_11491,N_10104,N_9043);
xor U11492 (N_11492,N_9211,N_9286);
or U11493 (N_11493,N_9400,N_10057);
nand U11494 (N_11494,N_10124,N_9802);
and U11495 (N_11495,N_10480,N_10391);
or U11496 (N_11496,N_9049,N_9432);
or U11497 (N_11497,N_10467,N_9625);
nand U11498 (N_11498,N_9356,N_9690);
xnor U11499 (N_11499,N_9198,N_10016);
nand U11500 (N_11500,N_9047,N_9582);
and U11501 (N_11501,N_9464,N_9859);
or U11502 (N_11502,N_9340,N_10386);
nand U11503 (N_11503,N_9814,N_10168);
or U11504 (N_11504,N_9110,N_9046);
and U11505 (N_11505,N_9506,N_10359);
or U11506 (N_11506,N_9903,N_9772);
nor U11507 (N_11507,N_9826,N_9424);
nand U11508 (N_11508,N_9548,N_10448);
and U11509 (N_11509,N_10256,N_9776);
and U11510 (N_11510,N_10468,N_9208);
or U11511 (N_11511,N_10008,N_9399);
or U11512 (N_11512,N_10306,N_9710);
nor U11513 (N_11513,N_9328,N_9344);
nor U11514 (N_11514,N_10399,N_10234);
xor U11515 (N_11515,N_9683,N_9853);
or U11516 (N_11516,N_10046,N_9118);
or U11517 (N_11517,N_10094,N_10373);
nand U11518 (N_11518,N_9078,N_9224);
xnor U11519 (N_11519,N_9117,N_10436);
nor U11520 (N_11520,N_9427,N_9661);
and U11521 (N_11521,N_9532,N_9541);
or U11522 (N_11522,N_9168,N_10318);
nor U11523 (N_11523,N_9775,N_10094);
nor U11524 (N_11524,N_9131,N_10289);
xnor U11525 (N_11525,N_9955,N_9804);
and U11526 (N_11526,N_9254,N_10264);
or U11527 (N_11527,N_10369,N_10414);
nand U11528 (N_11528,N_10337,N_9188);
nand U11529 (N_11529,N_9863,N_9232);
and U11530 (N_11530,N_9419,N_9490);
and U11531 (N_11531,N_10022,N_9121);
and U11532 (N_11532,N_9241,N_9195);
or U11533 (N_11533,N_10098,N_10028);
and U11534 (N_11534,N_9213,N_10485);
nand U11535 (N_11535,N_9866,N_9623);
xnor U11536 (N_11536,N_9084,N_9304);
and U11537 (N_11537,N_10419,N_9548);
nor U11538 (N_11538,N_9277,N_9194);
nand U11539 (N_11539,N_10470,N_9611);
nand U11540 (N_11540,N_9287,N_9705);
or U11541 (N_11541,N_9614,N_9098);
or U11542 (N_11542,N_9151,N_10462);
xor U11543 (N_11543,N_10438,N_10015);
xnor U11544 (N_11544,N_9561,N_10066);
nor U11545 (N_11545,N_10310,N_9589);
xor U11546 (N_11546,N_9575,N_10308);
xor U11547 (N_11547,N_10022,N_9017);
xnor U11548 (N_11548,N_9898,N_9926);
nand U11549 (N_11549,N_9991,N_9757);
and U11550 (N_11550,N_9405,N_9137);
or U11551 (N_11551,N_10004,N_10145);
and U11552 (N_11552,N_10189,N_10287);
nand U11553 (N_11553,N_9827,N_9256);
and U11554 (N_11554,N_9677,N_9991);
and U11555 (N_11555,N_10447,N_10366);
nor U11556 (N_11556,N_9238,N_9096);
xor U11557 (N_11557,N_9776,N_9068);
nor U11558 (N_11558,N_9048,N_9618);
nor U11559 (N_11559,N_9120,N_10176);
or U11560 (N_11560,N_9253,N_9455);
nand U11561 (N_11561,N_9078,N_10063);
xnor U11562 (N_11562,N_10475,N_10332);
nor U11563 (N_11563,N_10229,N_9488);
nor U11564 (N_11564,N_9169,N_10293);
nand U11565 (N_11565,N_10381,N_9373);
nor U11566 (N_11566,N_10051,N_9504);
or U11567 (N_11567,N_10479,N_9420);
nand U11568 (N_11568,N_10203,N_9292);
and U11569 (N_11569,N_9464,N_10061);
nand U11570 (N_11570,N_9615,N_9032);
nand U11571 (N_11571,N_10253,N_10483);
nor U11572 (N_11572,N_10233,N_9736);
or U11573 (N_11573,N_9476,N_10000);
xor U11574 (N_11574,N_9388,N_9891);
nor U11575 (N_11575,N_9719,N_10344);
nor U11576 (N_11576,N_10006,N_9021);
xor U11577 (N_11577,N_9189,N_9681);
xnor U11578 (N_11578,N_9030,N_9546);
and U11579 (N_11579,N_9575,N_9702);
or U11580 (N_11580,N_10437,N_9959);
nand U11581 (N_11581,N_10204,N_10276);
or U11582 (N_11582,N_10151,N_9314);
nand U11583 (N_11583,N_9344,N_10478);
xnor U11584 (N_11584,N_10388,N_10371);
nand U11585 (N_11585,N_9715,N_9858);
nand U11586 (N_11586,N_9936,N_9118);
or U11587 (N_11587,N_9899,N_10003);
and U11588 (N_11588,N_9918,N_9590);
and U11589 (N_11589,N_9176,N_9312);
xnor U11590 (N_11590,N_9942,N_9499);
and U11591 (N_11591,N_10332,N_9097);
nand U11592 (N_11592,N_9110,N_9359);
and U11593 (N_11593,N_9600,N_9118);
or U11594 (N_11594,N_10494,N_10361);
nor U11595 (N_11595,N_10268,N_9134);
or U11596 (N_11596,N_10028,N_9880);
and U11597 (N_11597,N_9131,N_10071);
nor U11598 (N_11598,N_9247,N_10167);
and U11599 (N_11599,N_9538,N_9989);
nand U11600 (N_11600,N_9914,N_9577);
nand U11601 (N_11601,N_9335,N_9219);
nand U11602 (N_11602,N_9232,N_10473);
nand U11603 (N_11603,N_10191,N_10126);
xnor U11604 (N_11604,N_9956,N_9303);
or U11605 (N_11605,N_9118,N_9026);
or U11606 (N_11606,N_9173,N_9745);
nand U11607 (N_11607,N_10302,N_10153);
or U11608 (N_11608,N_10399,N_10251);
and U11609 (N_11609,N_9603,N_9387);
and U11610 (N_11610,N_10054,N_9767);
nor U11611 (N_11611,N_10273,N_10051);
nand U11612 (N_11612,N_9762,N_9363);
nor U11613 (N_11613,N_9199,N_9894);
or U11614 (N_11614,N_10229,N_9365);
and U11615 (N_11615,N_10101,N_9260);
nand U11616 (N_11616,N_9856,N_10280);
or U11617 (N_11617,N_10385,N_10035);
and U11618 (N_11618,N_10399,N_9933);
nand U11619 (N_11619,N_10476,N_9518);
xor U11620 (N_11620,N_9589,N_9605);
nor U11621 (N_11621,N_9749,N_9665);
xnor U11622 (N_11622,N_10233,N_9443);
or U11623 (N_11623,N_10082,N_10170);
nand U11624 (N_11624,N_9729,N_10039);
xnor U11625 (N_11625,N_9337,N_9318);
xnor U11626 (N_11626,N_9380,N_9996);
or U11627 (N_11627,N_10448,N_9015);
nand U11628 (N_11628,N_10228,N_9080);
xnor U11629 (N_11629,N_9935,N_9542);
or U11630 (N_11630,N_9229,N_10099);
xnor U11631 (N_11631,N_9543,N_10226);
and U11632 (N_11632,N_10124,N_9590);
nand U11633 (N_11633,N_9446,N_9806);
xnor U11634 (N_11634,N_9514,N_9001);
or U11635 (N_11635,N_10440,N_10486);
nor U11636 (N_11636,N_9235,N_9797);
nor U11637 (N_11637,N_9554,N_9289);
nor U11638 (N_11638,N_10086,N_9875);
xor U11639 (N_11639,N_9047,N_9636);
nor U11640 (N_11640,N_10087,N_9117);
or U11641 (N_11641,N_10075,N_10166);
nor U11642 (N_11642,N_10018,N_9993);
nor U11643 (N_11643,N_9016,N_9937);
xor U11644 (N_11644,N_9085,N_9258);
nor U11645 (N_11645,N_9698,N_10235);
and U11646 (N_11646,N_9515,N_9120);
nand U11647 (N_11647,N_10125,N_10197);
xor U11648 (N_11648,N_9695,N_9909);
xnor U11649 (N_11649,N_9345,N_10488);
nand U11650 (N_11650,N_9912,N_10018);
xnor U11651 (N_11651,N_9538,N_9958);
nor U11652 (N_11652,N_9788,N_10443);
or U11653 (N_11653,N_9734,N_9206);
or U11654 (N_11654,N_10038,N_10191);
nand U11655 (N_11655,N_9319,N_9526);
nand U11656 (N_11656,N_9176,N_9514);
xnor U11657 (N_11657,N_10058,N_9447);
or U11658 (N_11658,N_9208,N_9067);
and U11659 (N_11659,N_9755,N_9651);
and U11660 (N_11660,N_10134,N_10205);
or U11661 (N_11661,N_9549,N_9783);
nor U11662 (N_11662,N_10382,N_9685);
nand U11663 (N_11663,N_10121,N_9259);
nor U11664 (N_11664,N_9129,N_10423);
and U11665 (N_11665,N_10116,N_10055);
nand U11666 (N_11666,N_9814,N_9726);
xnor U11667 (N_11667,N_9744,N_9702);
and U11668 (N_11668,N_9268,N_9532);
xor U11669 (N_11669,N_10439,N_9577);
nor U11670 (N_11670,N_9769,N_9176);
nor U11671 (N_11671,N_9132,N_10048);
and U11672 (N_11672,N_9473,N_9200);
and U11673 (N_11673,N_9608,N_9022);
nor U11674 (N_11674,N_9163,N_10308);
or U11675 (N_11675,N_10021,N_10455);
nor U11676 (N_11676,N_10001,N_9013);
and U11677 (N_11677,N_9458,N_9496);
xnor U11678 (N_11678,N_9287,N_9455);
or U11679 (N_11679,N_9148,N_9938);
xnor U11680 (N_11680,N_10036,N_10023);
and U11681 (N_11681,N_9997,N_9199);
or U11682 (N_11682,N_9630,N_10263);
and U11683 (N_11683,N_9407,N_9774);
and U11684 (N_11684,N_9377,N_9985);
xor U11685 (N_11685,N_9843,N_10306);
or U11686 (N_11686,N_9930,N_9276);
and U11687 (N_11687,N_10375,N_9459);
or U11688 (N_11688,N_10390,N_9538);
and U11689 (N_11689,N_10402,N_10457);
or U11690 (N_11690,N_10346,N_9177);
nor U11691 (N_11691,N_10423,N_9804);
xor U11692 (N_11692,N_9797,N_10280);
nand U11693 (N_11693,N_10415,N_9643);
and U11694 (N_11694,N_9589,N_10067);
nor U11695 (N_11695,N_9428,N_9744);
and U11696 (N_11696,N_9673,N_10162);
and U11697 (N_11697,N_9121,N_9265);
nand U11698 (N_11698,N_10175,N_9676);
and U11699 (N_11699,N_9190,N_9648);
or U11700 (N_11700,N_9811,N_9119);
xor U11701 (N_11701,N_9786,N_9896);
nor U11702 (N_11702,N_10298,N_9973);
xor U11703 (N_11703,N_9603,N_9743);
xnor U11704 (N_11704,N_9481,N_10175);
and U11705 (N_11705,N_9332,N_9371);
xnor U11706 (N_11706,N_10160,N_9256);
nor U11707 (N_11707,N_10459,N_9755);
or U11708 (N_11708,N_10488,N_9965);
nor U11709 (N_11709,N_9476,N_10061);
and U11710 (N_11710,N_9606,N_9198);
or U11711 (N_11711,N_10053,N_9632);
or U11712 (N_11712,N_9174,N_9643);
nor U11713 (N_11713,N_10206,N_9958);
xnor U11714 (N_11714,N_10033,N_9349);
and U11715 (N_11715,N_9732,N_10284);
nor U11716 (N_11716,N_10359,N_9951);
nand U11717 (N_11717,N_10049,N_9807);
and U11718 (N_11718,N_9740,N_9484);
nor U11719 (N_11719,N_9358,N_10014);
or U11720 (N_11720,N_9930,N_9298);
nand U11721 (N_11721,N_9894,N_10359);
or U11722 (N_11722,N_9280,N_10377);
nor U11723 (N_11723,N_10453,N_10495);
and U11724 (N_11724,N_10458,N_9638);
xnor U11725 (N_11725,N_9364,N_9525);
nor U11726 (N_11726,N_9283,N_9713);
or U11727 (N_11727,N_9472,N_9264);
xor U11728 (N_11728,N_10424,N_9929);
or U11729 (N_11729,N_9764,N_9186);
nand U11730 (N_11730,N_9463,N_9333);
and U11731 (N_11731,N_9096,N_9553);
xor U11732 (N_11732,N_10378,N_9016);
nand U11733 (N_11733,N_10347,N_9985);
xnor U11734 (N_11734,N_9299,N_10272);
or U11735 (N_11735,N_9719,N_9052);
and U11736 (N_11736,N_9386,N_10346);
nand U11737 (N_11737,N_9861,N_10287);
nand U11738 (N_11738,N_10378,N_9540);
and U11739 (N_11739,N_9600,N_9583);
or U11740 (N_11740,N_9703,N_9990);
nor U11741 (N_11741,N_9831,N_10112);
and U11742 (N_11742,N_9639,N_10409);
and U11743 (N_11743,N_9062,N_9710);
and U11744 (N_11744,N_9544,N_9985);
and U11745 (N_11745,N_10104,N_9384);
xor U11746 (N_11746,N_9349,N_9412);
nand U11747 (N_11747,N_9588,N_10470);
nand U11748 (N_11748,N_9679,N_9043);
nand U11749 (N_11749,N_9848,N_9813);
xnor U11750 (N_11750,N_10247,N_10260);
nor U11751 (N_11751,N_10283,N_9908);
nand U11752 (N_11752,N_10239,N_10333);
or U11753 (N_11753,N_10422,N_10298);
xnor U11754 (N_11754,N_10037,N_10432);
nand U11755 (N_11755,N_10356,N_9416);
and U11756 (N_11756,N_9524,N_9955);
nand U11757 (N_11757,N_9001,N_9375);
xor U11758 (N_11758,N_10002,N_9106);
nor U11759 (N_11759,N_9599,N_9725);
nor U11760 (N_11760,N_9805,N_10147);
and U11761 (N_11761,N_9870,N_9474);
and U11762 (N_11762,N_9848,N_10166);
xnor U11763 (N_11763,N_9385,N_10032);
or U11764 (N_11764,N_10166,N_10197);
or U11765 (N_11765,N_10202,N_10066);
xor U11766 (N_11766,N_9472,N_10481);
nand U11767 (N_11767,N_9166,N_9359);
and U11768 (N_11768,N_9477,N_10048);
xor U11769 (N_11769,N_9487,N_9701);
nand U11770 (N_11770,N_9171,N_10182);
or U11771 (N_11771,N_9486,N_9875);
nor U11772 (N_11772,N_9210,N_9850);
or U11773 (N_11773,N_10412,N_9091);
and U11774 (N_11774,N_9662,N_9236);
nand U11775 (N_11775,N_9033,N_9362);
nor U11776 (N_11776,N_9384,N_10401);
nor U11777 (N_11777,N_9010,N_10381);
nand U11778 (N_11778,N_10209,N_9819);
or U11779 (N_11779,N_9523,N_10230);
and U11780 (N_11780,N_10195,N_10183);
nand U11781 (N_11781,N_9424,N_9244);
xnor U11782 (N_11782,N_9057,N_10283);
and U11783 (N_11783,N_9408,N_9992);
nor U11784 (N_11784,N_9460,N_10090);
xnor U11785 (N_11785,N_9973,N_9632);
and U11786 (N_11786,N_9539,N_9373);
nand U11787 (N_11787,N_10064,N_9462);
nand U11788 (N_11788,N_9279,N_9001);
or U11789 (N_11789,N_9089,N_9354);
nor U11790 (N_11790,N_9416,N_9812);
and U11791 (N_11791,N_10354,N_10375);
xor U11792 (N_11792,N_9190,N_10070);
nor U11793 (N_11793,N_10442,N_9796);
nor U11794 (N_11794,N_9852,N_9820);
nor U11795 (N_11795,N_9452,N_9216);
xor U11796 (N_11796,N_9919,N_9236);
or U11797 (N_11797,N_10260,N_9803);
and U11798 (N_11798,N_9783,N_10170);
xor U11799 (N_11799,N_10454,N_9780);
and U11800 (N_11800,N_9648,N_9756);
and U11801 (N_11801,N_9766,N_9943);
nor U11802 (N_11802,N_9129,N_9051);
nor U11803 (N_11803,N_9964,N_9656);
nor U11804 (N_11804,N_10282,N_9708);
or U11805 (N_11805,N_9037,N_10093);
nand U11806 (N_11806,N_10318,N_10269);
nor U11807 (N_11807,N_10188,N_9619);
or U11808 (N_11808,N_9459,N_9220);
nand U11809 (N_11809,N_9998,N_9908);
and U11810 (N_11810,N_10292,N_10062);
nor U11811 (N_11811,N_9834,N_10361);
nor U11812 (N_11812,N_9856,N_9588);
nand U11813 (N_11813,N_10372,N_9368);
or U11814 (N_11814,N_10344,N_10161);
or U11815 (N_11815,N_10050,N_10168);
and U11816 (N_11816,N_9666,N_9463);
and U11817 (N_11817,N_10293,N_9997);
nor U11818 (N_11818,N_9185,N_9302);
nor U11819 (N_11819,N_9699,N_10218);
xor U11820 (N_11820,N_9726,N_9522);
nand U11821 (N_11821,N_10057,N_9541);
xor U11822 (N_11822,N_9992,N_10480);
nor U11823 (N_11823,N_10366,N_10227);
xor U11824 (N_11824,N_10382,N_9801);
or U11825 (N_11825,N_9821,N_10111);
xnor U11826 (N_11826,N_10371,N_9373);
nand U11827 (N_11827,N_9673,N_9086);
xor U11828 (N_11828,N_9828,N_9054);
nor U11829 (N_11829,N_9986,N_9627);
xnor U11830 (N_11830,N_9243,N_10258);
nor U11831 (N_11831,N_10117,N_10293);
and U11832 (N_11832,N_9529,N_9961);
or U11833 (N_11833,N_10081,N_9745);
nor U11834 (N_11834,N_9559,N_9616);
and U11835 (N_11835,N_9848,N_9874);
and U11836 (N_11836,N_9235,N_9009);
and U11837 (N_11837,N_9930,N_9540);
and U11838 (N_11838,N_9984,N_9334);
nor U11839 (N_11839,N_9260,N_9597);
xor U11840 (N_11840,N_9589,N_10433);
or U11841 (N_11841,N_9677,N_9966);
nand U11842 (N_11842,N_9916,N_9204);
nand U11843 (N_11843,N_9429,N_9526);
or U11844 (N_11844,N_9506,N_10334);
nand U11845 (N_11845,N_9695,N_9235);
nand U11846 (N_11846,N_10408,N_10438);
xor U11847 (N_11847,N_10143,N_9333);
and U11848 (N_11848,N_9199,N_9326);
and U11849 (N_11849,N_9468,N_9126);
nand U11850 (N_11850,N_10021,N_10227);
xor U11851 (N_11851,N_10255,N_9740);
or U11852 (N_11852,N_10033,N_10205);
or U11853 (N_11853,N_10250,N_9111);
nor U11854 (N_11854,N_9772,N_9991);
or U11855 (N_11855,N_9183,N_10169);
xor U11856 (N_11856,N_9296,N_9146);
nor U11857 (N_11857,N_9658,N_9723);
or U11858 (N_11858,N_9755,N_10249);
xor U11859 (N_11859,N_9295,N_9832);
nand U11860 (N_11860,N_10023,N_9472);
nand U11861 (N_11861,N_9334,N_9588);
xnor U11862 (N_11862,N_9716,N_10201);
nor U11863 (N_11863,N_9689,N_10350);
or U11864 (N_11864,N_9162,N_10007);
nand U11865 (N_11865,N_9915,N_10080);
and U11866 (N_11866,N_10282,N_9872);
nand U11867 (N_11867,N_9329,N_9112);
or U11868 (N_11868,N_9036,N_9447);
and U11869 (N_11869,N_10485,N_9395);
nor U11870 (N_11870,N_9060,N_10442);
or U11871 (N_11871,N_9930,N_9401);
or U11872 (N_11872,N_9574,N_9152);
or U11873 (N_11873,N_10199,N_9951);
and U11874 (N_11874,N_9611,N_9868);
nor U11875 (N_11875,N_9178,N_9770);
xor U11876 (N_11876,N_9060,N_9994);
or U11877 (N_11877,N_10081,N_9378);
nor U11878 (N_11878,N_9430,N_9758);
or U11879 (N_11879,N_9719,N_10070);
or U11880 (N_11880,N_9755,N_9436);
or U11881 (N_11881,N_10322,N_9993);
nor U11882 (N_11882,N_10102,N_10375);
nand U11883 (N_11883,N_9243,N_10219);
xor U11884 (N_11884,N_10202,N_9019);
nand U11885 (N_11885,N_10064,N_9607);
or U11886 (N_11886,N_10213,N_10097);
and U11887 (N_11887,N_10401,N_9196);
nor U11888 (N_11888,N_10390,N_9897);
or U11889 (N_11889,N_9752,N_9919);
nand U11890 (N_11890,N_9709,N_10368);
or U11891 (N_11891,N_9802,N_9760);
or U11892 (N_11892,N_9259,N_9768);
xnor U11893 (N_11893,N_9999,N_9291);
xor U11894 (N_11894,N_9786,N_10161);
nand U11895 (N_11895,N_9279,N_10394);
nand U11896 (N_11896,N_9839,N_10305);
nor U11897 (N_11897,N_10058,N_9803);
xor U11898 (N_11898,N_9731,N_9296);
nor U11899 (N_11899,N_9900,N_9525);
xnor U11900 (N_11900,N_9574,N_9993);
nand U11901 (N_11901,N_10098,N_10072);
and U11902 (N_11902,N_10020,N_9936);
nand U11903 (N_11903,N_9424,N_9560);
or U11904 (N_11904,N_9145,N_9223);
or U11905 (N_11905,N_10366,N_9477);
or U11906 (N_11906,N_9274,N_10410);
nor U11907 (N_11907,N_9975,N_9733);
nand U11908 (N_11908,N_9795,N_9056);
nand U11909 (N_11909,N_9328,N_9005);
or U11910 (N_11910,N_10057,N_9566);
xor U11911 (N_11911,N_10001,N_9728);
nor U11912 (N_11912,N_10290,N_10449);
nor U11913 (N_11913,N_9342,N_9739);
or U11914 (N_11914,N_9244,N_9877);
or U11915 (N_11915,N_9817,N_9069);
nand U11916 (N_11916,N_9644,N_10067);
and U11917 (N_11917,N_10139,N_9504);
xnor U11918 (N_11918,N_9305,N_9589);
and U11919 (N_11919,N_9199,N_10441);
and U11920 (N_11920,N_10190,N_10443);
and U11921 (N_11921,N_10313,N_9139);
xor U11922 (N_11922,N_9772,N_10147);
nor U11923 (N_11923,N_10421,N_9519);
and U11924 (N_11924,N_9213,N_9901);
nand U11925 (N_11925,N_10213,N_10352);
xor U11926 (N_11926,N_9188,N_9229);
xnor U11927 (N_11927,N_10495,N_9392);
xor U11928 (N_11928,N_9989,N_10100);
or U11929 (N_11929,N_9953,N_9727);
nor U11930 (N_11930,N_9331,N_10296);
or U11931 (N_11931,N_10325,N_9677);
and U11932 (N_11932,N_10356,N_9796);
xnor U11933 (N_11933,N_10045,N_9936);
nor U11934 (N_11934,N_9585,N_9131);
and U11935 (N_11935,N_9364,N_9089);
nand U11936 (N_11936,N_10223,N_10046);
nand U11937 (N_11937,N_10182,N_10359);
nor U11938 (N_11938,N_10253,N_9077);
nand U11939 (N_11939,N_9113,N_10454);
nand U11940 (N_11940,N_9484,N_9730);
or U11941 (N_11941,N_10246,N_9461);
or U11942 (N_11942,N_9020,N_9635);
nand U11943 (N_11943,N_10040,N_9628);
or U11944 (N_11944,N_10351,N_9795);
nor U11945 (N_11945,N_9951,N_10410);
nor U11946 (N_11946,N_9457,N_9384);
and U11947 (N_11947,N_10094,N_9055);
and U11948 (N_11948,N_10338,N_9080);
nand U11949 (N_11949,N_10469,N_10075);
nand U11950 (N_11950,N_9254,N_9618);
xnor U11951 (N_11951,N_9089,N_10225);
nand U11952 (N_11952,N_9701,N_10091);
or U11953 (N_11953,N_10430,N_10384);
and U11954 (N_11954,N_9646,N_9688);
and U11955 (N_11955,N_9447,N_9237);
xor U11956 (N_11956,N_10489,N_10143);
nor U11957 (N_11957,N_10175,N_9099);
or U11958 (N_11958,N_10300,N_10390);
or U11959 (N_11959,N_9686,N_10093);
nor U11960 (N_11960,N_9359,N_9622);
or U11961 (N_11961,N_9734,N_9934);
xnor U11962 (N_11962,N_9960,N_9874);
xor U11963 (N_11963,N_9900,N_9752);
nor U11964 (N_11964,N_10357,N_9108);
and U11965 (N_11965,N_9383,N_9884);
or U11966 (N_11966,N_9108,N_10398);
nor U11967 (N_11967,N_10066,N_9248);
and U11968 (N_11968,N_9200,N_9322);
or U11969 (N_11969,N_10032,N_9748);
nand U11970 (N_11970,N_9219,N_9882);
xor U11971 (N_11971,N_9389,N_9320);
or U11972 (N_11972,N_10298,N_9526);
nand U11973 (N_11973,N_10403,N_9283);
nand U11974 (N_11974,N_10181,N_9924);
xor U11975 (N_11975,N_9260,N_9344);
nand U11976 (N_11976,N_9144,N_9527);
and U11977 (N_11977,N_9671,N_9078);
and U11978 (N_11978,N_9361,N_9460);
and U11979 (N_11979,N_10062,N_9725);
nor U11980 (N_11980,N_9743,N_9199);
and U11981 (N_11981,N_9308,N_9188);
nand U11982 (N_11982,N_10073,N_9997);
or U11983 (N_11983,N_9894,N_9726);
and U11984 (N_11984,N_9894,N_9055);
xor U11985 (N_11985,N_9181,N_10212);
xnor U11986 (N_11986,N_9038,N_9219);
nand U11987 (N_11987,N_10459,N_10483);
and U11988 (N_11988,N_9136,N_9895);
xor U11989 (N_11989,N_10394,N_10404);
and U11990 (N_11990,N_10264,N_10460);
nor U11991 (N_11991,N_9337,N_10015);
nand U11992 (N_11992,N_9391,N_10304);
nand U11993 (N_11993,N_10403,N_10411);
and U11994 (N_11994,N_9600,N_9661);
or U11995 (N_11995,N_10161,N_10341);
nor U11996 (N_11996,N_9081,N_9829);
or U11997 (N_11997,N_10445,N_9589);
nor U11998 (N_11998,N_10430,N_9251);
or U11999 (N_11999,N_10064,N_9565);
nor U12000 (N_12000,N_10906,N_11425);
nand U12001 (N_12001,N_11895,N_10501);
and U12002 (N_12002,N_11161,N_11344);
nor U12003 (N_12003,N_11866,N_10712);
and U12004 (N_12004,N_10972,N_10996);
nand U12005 (N_12005,N_10647,N_10587);
xor U12006 (N_12006,N_10739,N_11351);
xor U12007 (N_12007,N_10576,N_10646);
nand U12008 (N_12008,N_11239,N_11499);
nand U12009 (N_12009,N_11748,N_11525);
and U12010 (N_12010,N_11500,N_11578);
nand U12011 (N_12011,N_11032,N_10849);
nand U12012 (N_12012,N_11126,N_11698);
nor U12013 (N_12013,N_11002,N_11579);
nand U12014 (N_12014,N_10567,N_11462);
xnor U12015 (N_12015,N_11106,N_11865);
and U12016 (N_12016,N_10971,N_11876);
xor U12017 (N_12017,N_10905,N_10948);
and U12018 (N_12018,N_11268,N_11181);
xnor U12019 (N_12019,N_11538,N_11175);
nor U12020 (N_12020,N_10880,N_10591);
and U12021 (N_12021,N_11202,N_11927);
nor U12022 (N_12022,N_11911,N_11632);
nand U12023 (N_12023,N_11154,N_11037);
nand U12024 (N_12024,N_11460,N_11364);
or U12025 (N_12025,N_10541,N_11017);
and U12026 (N_12026,N_11329,N_11281);
and U12027 (N_12027,N_10653,N_11055);
nor U12028 (N_12028,N_11070,N_11832);
nand U12029 (N_12029,N_11681,N_11254);
or U12030 (N_12030,N_11324,N_11881);
nand U12031 (N_12031,N_11802,N_11136);
nor U12032 (N_12032,N_11687,N_11516);
or U12033 (N_12033,N_11296,N_10584);
nor U12034 (N_12034,N_10837,N_11269);
nand U12035 (N_12035,N_10518,N_11323);
nand U12036 (N_12036,N_11609,N_10812);
xnor U12037 (N_12037,N_11200,N_11192);
and U12038 (N_12038,N_10525,N_10774);
nor U12039 (N_12039,N_11741,N_11084);
or U12040 (N_12040,N_11233,N_11640);
xnor U12041 (N_12041,N_11003,N_10984);
or U12042 (N_12042,N_11835,N_10630);
nand U12043 (N_12043,N_10607,N_11733);
nand U12044 (N_12044,N_11999,N_11820);
or U12045 (N_12045,N_11496,N_10960);
nor U12046 (N_12046,N_10750,N_11488);
and U12047 (N_12047,N_11121,N_11085);
and U12048 (N_12048,N_11814,N_11857);
and U12049 (N_12049,N_10519,N_11582);
xnor U12050 (N_12050,N_11886,N_10830);
nor U12051 (N_12051,N_11913,N_11683);
and U12052 (N_12052,N_11893,N_10779);
xnor U12053 (N_12053,N_11731,N_11091);
or U12054 (N_12054,N_11561,N_11197);
or U12055 (N_12055,N_11937,N_11674);
xor U12056 (N_12056,N_11860,N_11135);
and U12057 (N_12057,N_11479,N_11367);
nand U12058 (N_12058,N_10895,N_10717);
nand U12059 (N_12059,N_11259,N_10896);
or U12060 (N_12060,N_11973,N_11387);
nand U12061 (N_12061,N_11747,N_10556);
xor U12062 (N_12062,N_11558,N_11921);
or U12063 (N_12063,N_11401,N_11427);
nand U12064 (N_12064,N_11374,N_11332);
nor U12065 (N_12065,N_10531,N_10565);
and U12066 (N_12066,N_11095,N_11792);
nand U12067 (N_12067,N_11215,N_11616);
or U12068 (N_12068,N_10593,N_11411);
nor U12069 (N_12069,N_11724,N_10543);
xor U12070 (N_12070,N_10737,N_11679);
xor U12071 (N_12071,N_11313,N_11133);
nor U12072 (N_12072,N_10511,N_10904);
nand U12073 (N_12073,N_11399,N_10809);
or U12074 (N_12074,N_11097,N_11512);
nor U12075 (N_12075,N_11203,N_10752);
xnor U12076 (N_12076,N_11406,N_10644);
xnor U12077 (N_12077,N_10638,N_11027);
xnor U12078 (N_12078,N_11656,N_11416);
nand U12079 (N_12079,N_11436,N_10705);
or U12080 (N_12080,N_11537,N_11607);
or U12081 (N_12081,N_11306,N_11507);
and U12082 (N_12082,N_11584,N_10635);
nor U12083 (N_12083,N_10631,N_11829);
and U12084 (N_12084,N_11263,N_11847);
nor U12085 (N_12085,N_11685,N_11328);
xor U12086 (N_12086,N_11934,N_10754);
xnor U12087 (N_12087,N_11942,N_10934);
nor U12088 (N_12088,N_11129,N_11535);
and U12089 (N_12089,N_11874,N_11447);
nor U12090 (N_12090,N_10911,N_11429);
nand U12091 (N_12091,N_10965,N_11806);
or U12092 (N_12092,N_11041,N_11583);
nand U12093 (N_12093,N_10711,N_10862);
or U12094 (N_12094,N_11849,N_10944);
nor U12095 (N_12095,N_11896,N_11676);
nand U12096 (N_12096,N_11532,N_10522);
nor U12097 (N_12097,N_11998,N_11498);
and U12098 (N_12098,N_10695,N_11264);
nor U12099 (N_12099,N_11072,N_11255);
xnor U12100 (N_12100,N_11803,N_10514);
nand U12101 (N_12101,N_11650,N_10552);
nor U12102 (N_12102,N_11751,N_11932);
nand U12103 (N_12103,N_11780,N_11689);
nand U12104 (N_12104,N_10975,N_10852);
or U12105 (N_12105,N_11018,N_11625);
nor U12106 (N_12106,N_10732,N_10879);
nor U12107 (N_12107,N_10530,N_11164);
nand U12108 (N_12108,N_11162,N_11707);
and U12109 (N_12109,N_11840,N_10982);
or U12110 (N_12110,N_11050,N_11702);
and U12111 (N_12111,N_10561,N_10840);
and U12112 (N_12112,N_11441,N_11527);
and U12113 (N_12113,N_11450,N_11004);
and U12114 (N_12114,N_11423,N_11760);
and U12115 (N_12115,N_10641,N_10677);
or U12116 (N_12116,N_11524,N_11229);
or U12117 (N_12117,N_11530,N_11603);
nor U12118 (N_12118,N_11275,N_11856);
xor U12119 (N_12119,N_11930,N_11598);
xnor U12120 (N_12120,N_11761,N_10560);
xnor U12121 (N_12121,N_11504,N_11173);
or U12122 (N_12122,N_10835,N_10838);
or U12123 (N_12123,N_11737,N_11636);
and U12124 (N_12124,N_11972,N_11667);
nor U12125 (N_12125,N_11790,N_11920);
nor U12126 (N_12126,N_10990,N_11186);
or U12127 (N_12127,N_11428,N_10938);
xor U12128 (N_12128,N_10598,N_10819);
nand U12129 (N_12129,N_10824,N_11143);
nor U12130 (N_12130,N_11025,N_10997);
nand U12131 (N_12131,N_10640,N_11614);
nor U12132 (N_12132,N_10861,N_11333);
and U12133 (N_12133,N_10932,N_11812);
xnor U12134 (N_12134,N_11390,N_10766);
nor U12135 (N_12135,N_11246,N_11388);
nand U12136 (N_12136,N_11119,N_11049);
xnor U12137 (N_12137,N_11178,N_10691);
xor U12138 (N_12138,N_11848,N_11888);
and U12139 (N_12139,N_10998,N_11536);
nor U12140 (N_12140,N_11109,N_10915);
nor U12141 (N_12141,N_11916,N_11613);
nor U12142 (N_12142,N_10933,N_11809);
nand U12143 (N_12143,N_10509,N_11659);
or U12144 (N_12144,N_11470,N_10921);
xor U12145 (N_12145,N_11023,N_11120);
nor U12146 (N_12146,N_11997,N_11312);
xnor U12147 (N_12147,N_11398,N_11182);
and U12148 (N_12148,N_10860,N_11720);
or U12149 (N_12149,N_11692,N_10864);
xnor U12150 (N_12150,N_11563,N_11574);
or U12151 (N_12151,N_10970,N_10540);
xnor U12152 (N_12152,N_11377,N_11956);
nor U12153 (N_12153,N_11321,N_11690);
nand U12154 (N_12154,N_11189,N_11863);
or U12155 (N_12155,N_10558,N_10757);
nor U12156 (N_12156,N_10592,N_10622);
nand U12157 (N_12157,N_10871,N_10697);
nor U12158 (N_12158,N_11838,N_11458);
nand U12159 (N_12159,N_11358,N_11252);
xnor U12160 (N_12160,N_11483,N_11206);
and U12161 (N_12161,N_11785,N_10882);
nor U12162 (N_12162,N_11216,N_11648);
or U12163 (N_12163,N_10856,N_10987);
nor U12164 (N_12164,N_10920,N_11174);
or U12165 (N_12165,N_11871,N_11623);
nor U12166 (N_12166,N_11034,N_11278);
nand U12167 (N_12167,N_11240,N_11249);
nand U12168 (N_12168,N_10666,N_10648);
or U12169 (N_12169,N_11279,N_11311);
or U12170 (N_12170,N_10950,N_11082);
xor U12171 (N_12171,N_10733,N_10834);
or U12172 (N_12172,N_10555,N_11782);
and U12173 (N_12173,N_10942,N_10553);
nand U12174 (N_12174,N_11503,N_11058);
and U12175 (N_12175,N_11048,N_10801);
xnor U12176 (N_12176,N_10650,N_11123);
and U12177 (N_12177,N_10642,N_11836);
nor U12178 (N_12178,N_11984,N_11370);
or U12179 (N_12179,N_11457,N_11092);
and U12180 (N_12180,N_11317,N_10981);
and U12181 (N_12181,N_11381,N_10577);
and U12182 (N_12182,N_11168,N_11211);
xor U12183 (N_12183,N_10749,N_11982);
or U12184 (N_12184,N_11918,N_11601);
xnor U12185 (N_12185,N_11697,N_10776);
nand U12186 (N_12186,N_10758,N_10597);
nor U12187 (N_12187,N_11187,N_11993);
and U12188 (N_12188,N_11062,N_11088);
and U12189 (N_12189,N_11759,N_10545);
xnor U12190 (N_12190,N_11469,N_11908);
nor U12191 (N_12191,N_11622,N_11967);
or U12192 (N_12192,N_10741,N_10742);
or U12193 (N_12193,N_11083,N_11285);
xnor U12194 (N_12194,N_11585,N_11334);
nor U12195 (N_12195,N_10913,N_10544);
and U12196 (N_12196,N_10788,N_11686);
nand U12197 (N_12197,N_10993,N_10829);
or U12198 (N_12198,N_10925,N_11804);
nor U12199 (N_12199,N_10964,N_10989);
and U12200 (N_12200,N_11455,N_10775);
and U12201 (N_12201,N_10863,N_10656);
nor U12202 (N_12202,N_11850,N_11020);
or U12203 (N_12203,N_11319,N_11675);
nand U12204 (N_12204,N_11740,N_11193);
nand U12205 (N_12205,N_11734,N_10582);
and U12206 (N_12206,N_11854,N_11652);
xnor U12207 (N_12207,N_10515,N_11708);
or U12208 (N_12208,N_11823,N_11253);
or U12209 (N_12209,N_11201,N_11996);
and U12210 (N_12210,N_10782,N_11047);
and U12211 (N_12211,N_11494,N_11115);
nor U12212 (N_12212,N_10927,N_11872);
and U12213 (N_12213,N_10804,N_10557);
and U12214 (N_12214,N_11420,N_10872);
or U12215 (N_12215,N_11277,N_10969);
nand U12216 (N_12216,N_11672,N_11439);
xor U12217 (N_12217,N_11354,N_11506);
or U12218 (N_12218,N_11968,N_11940);
xor U12219 (N_12219,N_11900,N_11459);
nand U12220 (N_12220,N_10743,N_10894);
nand U12221 (N_12221,N_11959,N_11985);
or U12222 (N_12222,N_10551,N_11087);
and U12223 (N_12223,N_11620,N_10575);
nor U12224 (N_12224,N_11326,N_11565);
nand U12225 (N_12225,N_10976,N_11099);
nand U12226 (N_12226,N_10632,N_11188);
and U12227 (N_12227,N_10899,N_10727);
xnor U12228 (N_12228,N_11360,N_10859);
or U12229 (N_12229,N_11426,N_10523);
xor U12230 (N_12230,N_10818,N_10817);
or U12231 (N_12231,N_11247,N_11798);
nor U12232 (N_12232,N_11597,N_10667);
nand U12233 (N_12233,N_11012,N_11067);
or U12234 (N_12234,N_11361,N_11757);
and U12235 (N_12235,N_11052,N_11610);
xor U12236 (N_12236,N_11163,N_11774);
or U12237 (N_12237,N_11477,N_11978);
nand U12238 (N_12238,N_10617,N_11341);
and U12239 (N_12239,N_11534,N_10586);
nor U12240 (N_12240,N_11242,N_10759);
and U12241 (N_12241,N_11980,N_11631);
and U12242 (N_12242,N_11957,N_11555);
xor U12243 (N_12243,N_11294,N_11432);
nor U12244 (N_12244,N_11080,N_11238);
and U12245 (N_12245,N_10926,N_11693);
and U12246 (N_12246,N_11293,N_11875);
and U12247 (N_12247,N_10764,N_11299);
and U12248 (N_12248,N_11327,N_10596);
xor U12249 (N_12249,N_11094,N_11618);
xor U12250 (N_12250,N_11570,N_10985);
xnor U12251 (N_12251,N_11343,N_11624);
nor U12252 (N_12252,N_11413,N_11827);
or U12253 (N_12253,N_11042,N_11699);
and U12254 (N_12254,N_11237,N_11830);
xnor U12255 (N_12255,N_10763,N_10908);
nor U12256 (N_12256,N_10901,N_11864);
and U12257 (N_12257,N_11743,N_11873);
xnor U12258 (N_12258,N_10928,N_11262);
nand U12259 (N_12259,N_10686,N_11657);
xnor U12260 (N_12260,N_11190,N_10594);
xnor U12261 (N_12261,N_11437,N_10892);
xor U12262 (N_12262,N_11302,N_10671);
or U12263 (N_12263,N_11222,N_11396);
or U12264 (N_12264,N_10684,N_11663);
nor U12265 (N_12265,N_11726,N_10858);
and U12266 (N_12266,N_10947,N_11521);
or U12267 (N_12267,N_11762,N_10968);
or U12268 (N_12268,N_11209,N_10790);
xor U12269 (N_12269,N_10943,N_10747);
nand U12270 (N_12270,N_11635,N_11606);
xnor U12271 (N_12271,N_11588,N_11405);
and U12272 (N_12272,N_11495,N_11779);
nand U12273 (N_12273,N_10564,N_10799);
and U12274 (N_12274,N_11752,N_11770);
or U12275 (N_12275,N_11227,N_11764);
xnor U12276 (N_12276,N_11668,N_11904);
or U12277 (N_12277,N_10922,N_11452);
or U12278 (N_12278,N_10841,N_10923);
or U12279 (N_12279,N_11195,N_10599);
and U12280 (N_12280,N_10687,N_11905);
xnor U12281 (N_12281,N_11149,N_11038);
nand U12282 (N_12282,N_11591,N_11449);
nand U12283 (N_12283,N_11219,N_10959);
xnor U12284 (N_12284,N_11990,N_10548);
and U12285 (N_12285,N_11853,N_11571);
and U12286 (N_12286,N_11292,N_11412);
and U12287 (N_12287,N_10706,N_11977);
xor U12288 (N_12288,N_11270,N_11717);
and U12289 (N_12289,N_10612,N_10729);
nand U12290 (N_12290,N_11608,N_11128);
nor U12291 (N_12291,N_11898,N_11371);
nor U12292 (N_12292,N_10792,N_10581);
and U12293 (N_12293,N_11511,N_11156);
nand U12294 (N_12294,N_11950,N_11236);
nand U12295 (N_12295,N_10725,N_10713);
nor U12296 (N_12296,N_10603,N_11564);
nand U12297 (N_12297,N_11662,N_11706);
and U12298 (N_12298,N_11960,N_10798);
and U12299 (N_12299,N_10738,N_10736);
xor U12300 (N_12300,N_10977,N_10827);
or U12301 (N_12301,N_11651,N_11039);
or U12302 (N_12302,N_10869,N_11710);
and U12303 (N_12303,N_10655,N_10602);
and U12304 (N_12304,N_11011,N_11112);
xnor U12305 (N_12305,N_11947,N_11643);
and U12306 (N_12306,N_10802,N_11653);
nand U12307 (N_12307,N_11513,N_11595);
or U12308 (N_12308,N_11291,N_11304);
nor U12309 (N_12309,N_10888,N_10781);
and U12310 (N_12310,N_11079,N_10504);
or U12311 (N_12311,N_11783,N_10589);
xor U12312 (N_12312,N_11604,N_10506);
nor U12313 (N_12313,N_11348,N_11443);
nand U12314 (N_12314,N_11258,N_11475);
nor U12315 (N_12315,N_10626,N_11152);
nand U12316 (N_12316,N_10953,N_11124);
and U12317 (N_12317,N_11907,N_11446);
and U12318 (N_12318,N_10930,N_10949);
or U12319 (N_12319,N_11402,N_11251);
and U12320 (N_12320,N_11705,N_11111);
nand U12321 (N_12321,N_11194,N_10780);
or U12322 (N_12322,N_11283,N_10615);
nand U12323 (N_12323,N_11965,N_11014);
and U12324 (N_12324,N_10855,N_10857);
nand U12325 (N_12325,N_11403,N_10669);
nand U12326 (N_12326,N_10562,N_11397);
nand U12327 (N_12327,N_11979,N_11533);
xnor U12328 (N_12328,N_11592,N_10878);
and U12329 (N_12329,N_11922,N_10848);
nand U12330 (N_12330,N_11260,N_11562);
and U12331 (N_12331,N_10570,N_10625);
or U12332 (N_12332,N_10580,N_11223);
xnor U12333 (N_12333,N_11101,N_11081);
nand U12334 (N_12334,N_11515,N_10751);
and U12335 (N_12335,N_10778,N_11725);
and U12336 (N_12336,N_10865,N_11666);
xor U12337 (N_12337,N_11815,N_11290);
nor U12338 (N_12338,N_11243,N_10786);
and U12339 (N_12339,N_11822,N_10728);
nor U12340 (N_12340,N_10692,N_10924);
nand U12341 (N_12341,N_10973,N_10636);
nand U12342 (N_12342,N_10867,N_11730);
nand U12343 (N_12343,N_11870,N_11303);
and U12344 (N_12344,N_11655,N_11357);
xnor U12345 (N_12345,N_10701,N_11917);
xnor U12346 (N_12346,N_11395,N_10670);
and U12347 (N_12347,N_11590,N_11064);
and U12348 (N_12348,N_11821,N_11071);
nor U12349 (N_12349,N_11104,N_10508);
xnor U12350 (N_12350,N_11245,N_10874);
and U12351 (N_12351,N_10868,N_10681);
nand U12352 (N_12352,N_11518,N_11946);
nand U12353 (N_12353,N_10931,N_10688);
xor U12354 (N_12354,N_10843,N_11867);
and U12355 (N_12355,N_10682,N_11573);
xor U12356 (N_12356,N_11713,N_11224);
or U12357 (N_12357,N_11941,N_11150);
nand U12358 (N_12358,N_10994,N_11819);
and U12359 (N_12359,N_11755,N_11198);
xnor U12360 (N_12360,N_11502,N_10715);
xor U12361 (N_12361,N_11786,N_11673);
or U12362 (N_12362,N_11409,N_11926);
and U12363 (N_12363,N_11811,N_10574);
nor U12364 (N_12364,N_11523,N_11093);
nor U12365 (N_12365,N_10929,N_10995);
xor U12366 (N_12366,N_10816,N_10621);
or U12367 (N_12367,N_11028,N_11468);
or U12368 (N_12368,N_11943,N_10619);
nand U12369 (N_12369,N_11953,N_11061);
nand U12370 (N_12370,N_11176,N_11077);
nor U12371 (N_12371,N_11378,N_11885);
and U12372 (N_12372,N_11880,N_11694);
nand U12373 (N_12373,N_11484,N_11744);
xnor U12374 (N_12374,N_11955,N_11805);
or U12375 (N_12375,N_11424,N_11289);
and U12376 (N_12376,N_10572,N_11817);
or U12377 (N_12377,N_11855,N_10955);
nor U12378 (N_12378,N_11529,N_10524);
xor U12379 (N_12379,N_11665,N_11975);
nor U12380 (N_12380,N_10588,N_11700);
nor U12381 (N_12381,N_11753,N_10900);
xor U12382 (N_12382,N_11218,N_10726);
or U12383 (N_12383,N_11497,N_11400);
or U12384 (N_12384,N_10794,N_10730);
nor U12385 (N_12385,N_11501,N_10696);
xnor U12386 (N_12386,N_11221,N_10919);
nor U12387 (N_12387,N_10777,N_10634);
and U12388 (N_12388,N_11031,N_11723);
or U12389 (N_12389,N_10645,N_11248);
xnor U12390 (N_12390,N_11954,N_11105);
and U12391 (N_12391,N_11711,N_11630);
or U12392 (N_12392,N_10673,N_11330);
or U12393 (N_12393,N_11989,N_11266);
nor U12394 (N_12394,N_11474,N_10623);
xnor U12395 (N_12395,N_11988,N_11777);
nand U12396 (N_12396,N_11345,N_11491);
nor U12397 (N_12397,N_11791,N_11056);
or U12398 (N_12398,N_10568,N_11756);
nor U12399 (N_12399,N_11362,N_11580);
xnor U12400 (N_12400,N_11046,N_11137);
nor U12401 (N_12401,N_11554,N_11615);
or U12402 (N_12402,N_10643,N_11931);
nor U12403 (N_12403,N_10909,N_10611);
nand U12404 (N_12404,N_11828,N_10633);
xor U12405 (N_12405,N_10753,N_11465);
nor U12406 (N_12406,N_11519,N_11925);
and U12407 (N_12407,N_10585,N_11671);
and U12408 (N_12408,N_11379,N_11271);
nand U12409 (N_12409,N_11001,N_11964);
or U12410 (N_12410,N_11076,N_11131);
and U12411 (N_12411,N_10952,N_11546);
xnor U12412 (N_12412,N_11750,N_11818);
and U12413 (N_12413,N_10527,N_10659);
nand U12414 (N_12414,N_11540,N_11295);
and U12415 (N_12415,N_10748,N_11634);
and U12416 (N_12416,N_10590,N_11600);
nor U12417 (N_12417,N_11172,N_11602);
nor U12418 (N_12418,N_11763,N_11102);
nor U12419 (N_12419,N_11138,N_11440);
nor U12420 (N_12420,N_11421,N_10986);
nor U12421 (N_12421,N_11408,N_11765);
nand U12422 (N_12422,N_11183,N_11909);
xor U12423 (N_12423,N_10559,N_11471);
xor U12424 (N_12424,N_11727,N_10898);
xnor U12425 (N_12425,N_10660,N_10566);
nand U12426 (N_12426,N_11781,N_10658);
nor U12427 (N_12427,N_10958,N_10604);
or U12428 (N_12428,N_11257,N_11331);
and U12429 (N_12429,N_11297,N_10844);
nor U12430 (N_12430,N_10999,N_10704);
xnor U12431 (N_12431,N_11349,N_11526);
and U12432 (N_12432,N_11619,N_11912);
nor U12433 (N_12433,N_11068,N_10912);
nand U12434 (N_12434,N_11030,N_11180);
nand U12435 (N_12435,N_11766,N_11235);
or U12436 (N_12436,N_10845,N_11134);
nand U12437 (N_12437,N_10839,N_11418);
or U12438 (N_12438,N_11844,N_11810);
nand U12439 (N_12439,N_11974,N_11721);
xor U12440 (N_12440,N_11122,N_10500);
xnor U12441 (N_12441,N_11899,N_11894);
nand U12442 (N_12442,N_10698,N_11575);
or U12443 (N_12443,N_11026,N_10502);
and U12444 (N_12444,N_11641,N_11029);
nand U12445 (N_12445,N_11688,N_11280);
nor U12446 (N_12446,N_11794,N_11318);
xnor U12447 (N_12447,N_11214,N_11910);
nor U12448 (N_12448,N_10886,N_11678);
and U12449 (N_12449,N_11556,N_11576);
or U12450 (N_12450,N_11649,N_10966);
and U12451 (N_12451,N_11435,N_11664);
nand U12452 (N_12452,N_11843,N_11165);
nor U12453 (N_12453,N_11628,N_11605);
xor U12454 (N_12454,N_11308,N_11557);
nand U12455 (N_12455,N_11098,N_11928);
nor U12456 (N_12456,N_10690,N_11919);
nand U12457 (N_12457,N_10520,N_11417);
or U12458 (N_12458,N_10785,N_10517);
nor U12459 (N_12459,N_10674,N_11581);
xor U12460 (N_12460,N_10866,N_10988);
xor U12461 (N_12461,N_11878,N_11670);
xnor U12462 (N_12462,N_11626,N_10967);
xnor U12463 (N_12463,N_10979,N_10808);
or U12464 (N_12464,N_11144,N_11044);
or U12465 (N_12465,N_11191,N_11482);
xnor U12466 (N_12466,N_10639,N_11695);
nand U12467 (N_12467,N_11914,N_10832);
or U12468 (N_12468,N_11113,N_11852);
and U12469 (N_12469,N_11593,N_11480);
or U12470 (N_12470,N_10569,N_11903);
or U12471 (N_12471,N_11566,N_10980);
xnor U12472 (N_12472,N_11244,N_11572);
or U12473 (N_12473,N_11463,N_11948);
xnor U12474 (N_12474,N_11066,N_10722);
nor U12475 (N_12475,N_11587,N_10554);
nand U12476 (N_12476,N_11991,N_11445);
nand U12477 (N_12477,N_11808,N_10710);
nor U12478 (N_12478,N_10770,N_11793);
or U12479 (N_12479,N_10700,N_11212);
nand U12480 (N_12480,N_11736,N_11551);
nor U12481 (N_12481,N_11315,N_10618);
or U12482 (N_12482,N_11594,N_11718);
or U12483 (N_12483,N_11735,N_11489);
nor U12484 (N_12484,N_11325,N_10825);
nor U12485 (N_12485,N_11386,N_10836);
or U12486 (N_12486,N_10795,N_11684);
nand U12487 (N_12487,N_11231,N_11701);
or U12488 (N_12488,N_10610,N_11282);
or U12489 (N_12489,N_11745,N_11320);
nand U12490 (N_12490,N_11544,N_11531);
and U12491 (N_12491,N_11359,N_11185);
xor U12492 (N_12492,N_10893,N_11966);
xnor U12493 (N_12493,N_10534,N_10870);
xor U12494 (N_12494,N_11207,N_10961);
nor U12495 (N_12495,N_11448,N_11069);
nor U12496 (N_12496,N_10884,N_11891);
or U12497 (N_12497,N_10745,N_11797);
or U12498 (N_12498,N_11276,N_11310);
and U12499 (N_12499,N_11116,N_10744);
or U12500 (N_12500,N_11589,N_10516);
and U12501 (N_12501,N_11936,N_10724);
xnor U12502 (N_12502,N_11958,N_10689);
nand U12503 (N_12503,N_11472,N_10546);
xor U12504 (N_12504,N_10873,N_11890);
xor U12505 (N_12505,N_11442,N_11250);
nand U12506 (N_12506,N_11043,N_10628);
xnor U12507 (N_12507,N_11868,N_10579);
nand U12508 (N_12508,N_11179,N_11438);
nor U12509 (N_12509,N_11073,N_11145);
and U12510 (N_12510,N_10627,N_10956);
or U12511 (N_12511,N_10936,N_11778);
or U12512 (N_12512,N_10772,N_11389);
or U12513 (N_12513,N_10897,N_10721);
and U12514 (N_12514,N_11125,N_10784);
xnor U12515 (N_12515,N_11944,N_11226);
or U12516 (N_12516,N_11419,N_11035);
nor U12517 (N_12517,N_11464,N_11009);
nand U12518 (N_12518,N_10536,N_10538);
or U12519 (N_12519,N_10914,N_10796);
or U12520 (N_12520,N_11430,N_11159);
nand U12521 (N_12521,N_10791,N_10963);
and U12522 (N_12522,N_10746,N_10854);
xnor U12523 (N_12523,N_10815,N_10851);
nor U12524 (N_12524,N_11383,N_10760);
nand U12525 (N_12525,N_11141,N_11771);
and U12526 (N_12526,N_10537,N_11611);
xor U12527 (N_12527,N_11256,N_11510);
or U12528 (N_12528,N_11205,N_11008);
nand U12529 (N_12529,N_11013,N_11007);
nand U12530 (N_12530,N_11487,N_11380);
and U12531 (N_12531,N_11644,N_11709);
or U12532 (N_12532,N_10654,N_11100);
or U12533 (N_12533,N_11177,N_11935);
and U12534 (N_12534,N_11772,N_10693);
and U12535 (N_12535,N_11669,N_11824);
nand U12536 (N_12536,N_11040,N_11274);
or U12537 (N_12537,N_10842,N_11542);
xnor U12538 (N_12538,N_11170,N_11393);
nand U12539 (N_12539,N_10797,N_11261);
or U12540 (N_12540,N_11340,N_11879);
xor U12541 (N_12541,N_10761,N_10992);
xnor U12542 (N_12542,N_10740,N_11410);
xor U12543 (N_12543,N_11691,N_11356);
xor U12544 (N_12544,N_11451,N_11375);
nand U12545 (N_12545,N_11833,N_11807);
and U12546 (N_12546,N_10821,N_11166);
xnor U12547 (N_12547,N_10941,N_11831);
or U12548 (N_12548,N_11660,N_11627);
xnor U12549 (N_12549,N_11729,N_10573);
nor U12550 (N_12550,N_11075,N_11638);
nand U12551 (N_12551,N_11716,N_11902);
xor U12552 (N_12552,N_10716,N_11090);
or U12553 (N_12553,N_10547,N_11033);
nand U12554 (N_12554,N_11799,N_10793);
nor U12555 (N_12555,N_11987,N_11148);
xor U12556 (N_12556,N_11858,N_11712);
nand U12557 (N_12557,N_10767,N_10510);
xnor U12558 (N_12558,N_11859,N_11924);
nand U12559 (N_12559,N_11976,N_11877);
or U12560 (N_12560,N_11434,N_10755);
nand U12561 (N_12561,N_11316,N_11146);
nand U12562 (N_12562,N_11637,N_11784);
nand U12563 (N_12563,N_11365,N_10629);
nand U12564 (N_12564,N_11995,N_11127);
or U12565 (N_12565,N_10890,N_11739);
and U12566 (N_12566,N_11951,N_11599);
nand U12567 (N_12567,N_10850,N_11407);
nand U12568 (N_12568,N_11517,N_10550);
and U12569 (N_12569,N_11228,N_11719);
nand U12570 (N_12570,N_11971,N_11476);
nand U12571 (N_12571,N_10946,N_11220);
xnor U12572 (N_12572,N_11338,N_11816);
xnor U12573 (N_12573,N_10651,N_11915);
nand U12574 (N_12574,N_11103,N_11742);
nor U12575 (N_12575,N_11961,N_11204);
nand U12576 (N_12576,N_11086,N_10664);
nor U12577 (N_12577,N_11298,N_11633);
or U12578 (N_12578,N_11963,N_11454);
or U12579 (N_12579,N_11906,N_10678);
or U12580 (N_12580,N_11107,N_11654);
xnor U12581 (N_12581,N_10803,N_11994);
xnor U12582 (N_12582,N_11549,N_11490);
nand U12583 (N_12583,N_10846,N_10652);
xor U12584 (N_12584,N_11461,N_10608);
or U12585 (N_12585,N_10614,N_10823);
or U12586 (N_12586,N_11481,N_11108);
nand U12587 (N_12587,N_11834,N_10807);
xnor U12588 (N_12588,N_11057,N_10902);
nand U12589 (N_12589,N_11983,N_11225);
nand U12590 (N_12590,N_11514,N_11063);
nand U12591 (N_12591,N_10661,N_11142);
nand U12592 (N_12592,N_10595,N_10613);
xor U12593 (N_12593,N_11749,N_11157);
nand U12594 (N_12594,N_11147,N_10578);
nand U12595 (N_12595,N_10683,N_11884);
nor U12596 (N_12596,N_11682,N_11139);
or U12597 (N_12597,N_10800,N_11728);
nand U12598 (N_12598,N_11006,N_11078);
or U12599 (N_12599,N_11796,N_10983);
or U12600 (N_12600,N_11897,N_11234);
nor U12601 (N_12601,N_11862,N_11369);
nor U12602 (N_12602,N_11586,N_11130);
or U12603 (N_12603,N_10820,N_11933);
nor U12604 (N_12604,N_11629,N_11000);
or U12605 (N_12605,N_10789,N_11769);
and U12606 (N_12606,N_11869,N_10907);
nand U12607 (N_12607,N_11775,N_11232);
or U12608 (N_12608,N_10549,N_10676);
and U12609 (N_12609,N_10680,N_11846);
or U12610 (N_12610,N_10771,N_11677);
and U12611 (N_12611,N_11962,N_11553);
and U12612 (N_12612,N_11284,N_11569);
and U12613 (N_12613,N_10539,N_10571);
nand U12614 (N_12614,N_11732,N_11547);
or U12615 (N_12615,N_11153,N_11696);
xor U12616 (N_12616,N_10535,N_11617);
xor U12617 (N_12617,N_11704,N_10814);
xor U12618 (N_12618,N_11845,N_11404);
nand U12619 (N_12619,N_11074,N_10723);
and U12620 (N_12620,N_11372,N_11520);
xor U12621 (N_12621,N_11355,N_10765);
nor U12622 (N_12622,N_10624,N_10605);
xor U12623 (N_12623,N_11051,N_10877);
nor U12624 (N_12624,N_10945,N_10910);
xor U12625 (N_12625,N_10526,N_11199);
or U12626 (N_12626,N_10917,N_11171);
and U12627 (N_12627,N_11339,N_10806);
xor U12628 (N_12628,N_11473,N_10885);
nor U12629 (N_12629,N_10935,N_11889);
and U12630 (N_12630,N_11680,N_11612);
nand U12631 (N_12631,N_11768,N_11923);
xor U12632 (N_12632,N_11350,N_11314);
xnor U12633 (N_12633,N_11167,N_11505);
or U12634 (N_12634,N_11347,N_10620);
and U12635 (N_12635,N_11486,N_11132);
nor U12636 (N_12636,N_11053,N_11839);
xnor U12637 (N_12637,N_11813,N_11342);
or U12638 (N_12638,N_10811,N_11528);
and U12639 (N_12639,N_11060,N_11970);
or U12640 (N_12640,N_10606,N_11639);
nor U12641 (N_12641,N_10563,N_10637);
xnor U12642 (N_12642,N_11883,N_11015);
nand U12643 (N_12643,N_11552,N_10718);
xor U12644 (N_12644,N_11621,N_11160);
nand U12645 (N_12645,N_11022,N_10918);
xor U12646 (N_12646,N_11433,N_11096);
xor U12647 (N_12647,N_11305,N_11208);
and U12648 (N_12648,N_11826,N_10507);
and U12649 (N_12649,N_11522,N_11336);
nand U12650 (N_12650,N_10954,N_10665);
and U12651 (N_12651,N_11478,N_10609);
nor U12652 (N_12652,N_10903,N_11010);
nand U12653 (N_12653,N_11089,N_10672);
or U12654 (N_12654,N_11415,N_11887);
or U12655 (N_12655,N_11841,N_11352);
and U12656 (N_12656,N_11938,N_11114);
and U12657 (N_12657,N_10978,N_11414);
nand U12658 (N_12658,N_11541,N_11661);
and U12659 (N_12659,N_11543,N_10735);
nand U12660 (N_12660,N_10769,N_11596);
and U12661 (N_12661,N_10876,N_11882);
xor U12662 (N_12662,N_10601,N_11939);
and U12663 (N_12663,N_11485,N_11776);
or U12664 (N_12664,N_11754,N_11337);
or U12665 (N_12665,N_10685,N_11385);
or U12666 (N_12666,N_11568,N_11059);
xnor U12667 (N_12667,N_11851,N_10708);
xnor U12668 (N_12668,N_11353,N_11322);
and U12669 (N_12669,N_11265,N_11548);
xnor U12670 (N_12670,N_11508,N_10957);
nor U12671 (N_12671,N_11384,N_11065);
and U12672 (N_12672,N_11493,N_11738);
nor U12673 (N_12673,N_11492,N_10731);
nor U12674 (N_12674,N_11422,N_10937);
xor U12675 (N_12675,N_10756,N_11301);
nor U12676 (N_12676,N_11758,N_11949);
and U12677 (N_12677,N_10962,N_10694);
xor U12678 (N_12678,N_11158,N_10887);
xor U12679 (N_12679,N_11658,N_11795);
and U12680 (N_12680,N_10810,N_11210);
and U12681 (N_12681,N_10503,N_10881);
nand U12682 (N_12682,N_11453,N_10702);
xnor U12683 (N_12683,N_11550,N_11024);
nor U12684 (N_12684,N_10831,N_11288);
xor U12685 (N_12685,N_11929,N_11184);
nor U12686 (N_12686,N_11560,N_11267);
and U12687 (N_12687,N_11901,N_11789);
nand U12688 (N_12688,N_10891,N_11307);
nand U12689 (N_12689,N_10528,N_10826);
xnor U12690 (N_12690,N_10853,N_10521);
and U12691 (N_12691,N_11969,N_11773);
nor U12692 (N_12692,N_10822,N_10663);
nand U12693 (N_12693,N_10916,N_10720);
or U12694 (N_12694,N_10773,N_11545);
xor U12695 (N_12695,N_11992,N_10707);
and U12696 (N_12696,N_11016,N_10512);
or U12697 (N_12697,N_10662,N_10533);
nor U12698 (N_12698,N_10709,N_11054);
nor U12699 (N_12699,N_10833,N_11788);
or U12700 (N_12700,N_10734,N_11366);
xor U12701 (N_12701,N_11036,N_11952);
and U12702 (N_12702,N_11825,N_10951);
and U12703 (N_12703,N_10649,N_11431);
or U12704 (N_12704,N_11273,N_11703);
or U12705 (N_12705,N_11241,N_11456);
and U12706 (N_12706,N_11981,N_11986);
or U12707 (N_12707,N_11300,N_10883);
xnor U12708 (N_12708,N_10940,N_10542);
or U12709 (N_12709,N_10768,N_11230);
and U12710 (N_12710,N_11892,N_10668);
xor U12711 (N_12711,N_11376,N_10828);
xor U12712 (N_12712,N_11110,N_11151);
or U12713 (N_12713,N_11715,N_10813);
nand U12714 (N_12714,N_11287,N_11767);
xnor U12715 (N_12715,N_11140,N_11005);
or U12716 (N_12716,N_10529,N_10783);
nand U12717 (N_12717,N_11019,N_10714);
and U12718 (N_12718,N_10679,N_11722);
nand U12719 (N_12719,N_10875,N_11382);
nand U12720 (N_12720,N_11272,N_11309);
xor U12721 (N_12721,N_10974,N_10805);
or U12722 (N_12722,N_10699,N_11645);
nand U12723 (N_12723,N_11021,N_10616);
nor U12724 (N_12724,N_10532,N_11577);
and U12725 (N_12725,N_10762,N_11444);
or U12726 (N_12726,N_11800,N_11714);
nand U12727 (N_12727,N_11213,N_11567);
and U12728 (N_12728,N_10505,N_11394);
or U12729 (N_12729,N_11155,N_11509);
or U12730 (N_12730,N_10787,N_11392);
xnor U12731 (N_12731,N_11801,N_11363);
nor U12732 (N_12732,N_11559,N_11945);
nor U12733 (N_12733,N_10719,N_11837);
nor U12734 (N_12734,N_11746,N_11861);
or U12735 (N_12735,N_10583,N_10991);
or U12736 (N_12736,N_11346,N_11335);
xnor U12737 (N_12737,N_11286,N_11196);
xor U12738 (N_12738,N_11391,N_11368);
and U12739 (N_12739,N_11539,N_10600);
and U12740 (N_12740,N_11373,N_11647);
or U12741 (N_12741,N_10889,N_11842);
nand U12742 (N_12742,N_11045,N_11217);
nand U12743 (N_12743,N_10703,N_10657);
or U12744 (N_12744,N_10847,N_10939);
xnor U12745 (N_12745,N_11646,N_10675);
and U12746 (N_12746,N_11466,N_11117);
and U12747 (N_12747,N_11169,N_11118);
nor U12748 (N_12748,N_10513,N_11787);
nor U12749 (N_12749,N_11642,N_11467);
nand U12750 (N_12750,N_11086,N_11242);
or U12751 (N_12751,N_10523,N_11262);
or U12752 (N_12752,N_11249,N_11557);
nand U12753 (N_12753,N_11020,N_11589);
and U12754 (N_12754,N_11121,N_11211);
xnor U12755 (N_12755,N_11068,N_10611);
nand U12756 (N_12756,N_11796,N_11777);
or U12757 (N_12757,N_10959,N_10516);
nand U12758 (N_12758,N_10996,N_11166);
nor U12759 (N_12759,N_11520,N_10975);
nand U12760 (N_12760,N_10637,N_10521);
nand U12761 (N_12761,N_11430,N_10528);
xor U12762 (N_12762,N_11312,N_11357);
nand U12763 (N_12763,N_11911,N_10535);
nand U12764 (N_12764,N_11542,N_11085);
and U12765 (N_12765,N_11610,N_11653);
nor U12766 (N_12766,N_11041,N_11414);
xor U12767 (N_12767,N_11075,N_11135);
nor U12768 (N_12768,N_11282,N_11430);
nand U12769 (N_12769,N_10706,N_11642);
xor U12770 (N_12770,N_11618,N_10601);
and U12771 (N_12771,N_10876,N_11635);
xnor U12772 (N_12772,N_10981,N_11161);
and U12773 (N_12773,N_11994,N_11989);
and U12774 (N_12774,N_10596,N_11814);
and U12775 (N_12775,N_11611,N_11164);
nor U12776 (N_12776,N_11858,N_10684);
nor U12777 (N_12777,N_11358,N_10886);
nor U12778 (N_12778,N_10568,N_11833);
nand U12779 (N_12779,N_11058,N_11453);
and U12780 (N_12780,N_11975,N_11698);
nand U12781 (N_12781,N_11652,N_11404);
nor U12782 (N_12782,N_11951,N_10731);
xnor U12783 (N_12783,N_10581,N_11285);
nand U12784 (N_12784,N_10676,N_11874);
nor U12785 (N_12785,N_11567,N_11212);
xnor U12786 (N_12786,N_10628,N_11493);
nor U12787 (N_12787,N_10666,N_11726);
or U12788 (N_12788,N_10990,N_10707);
nor U12789 (N_12789,N_10699,N_11186);
nor U12790 (N_12790,N_11494,N_10744);
or U12791 (N_12791,N_10912,N_10932);
xnor U12792 (N_12792,N_11766,N_10821);
nor U12793 (N_12793,N_11879,N_11814);
or U12794 (N_12794,N_10779,N_10658);
and U12795 (N_12795,N_11052,N_10869);
nor U12796 (N_12796,N_11003,N_10556);
nand U12797 (N_12797,N_11664,N_11057);
xnor U12798 (N_12798,N_10604,N_11093);
nor U12799 (N_12799,N_10853,N_11079);
and U12800 (N_12800,N_11392,N_10790);
or U12801 (N_12801,N_10858,N_11891);
nor U12802 (N_12802,N_10985,N_11332);
or U12803 (N_12803,N_10981,N_10512);
and U12804 (N_12804,N_11914,N_10770);
nand U12805 (N_12805,N_11423,N_11798);
or U12806 (N_12806,N_11062,N_11355);
or U12807 (N_12807,N_10984,N_11001);
nor U12808 (N_12808,N_11693,N_11821);
xnor U12809 (N_12809,N_10855,N_11208);
nor U12810 (N_12810,N_11087,N_11421);
nor U12811 (N_12811,N_11373,N_11649);
xor U12812 (N_12812,N_11334,N_11214);
nand U12813 (N_12813,N_11092,N_10686);
and U12814 (N_12814,N_11428,N_11128);
or U12815 (N_12815,N_10568,N_11572);
nand U12816 (N_12816,N_11444,N_11362);
and U12817 (N_12817,N_11799,N_11605);
nor U12818 (N_12818,N_10842,N_11112);
xnor U12819 (N_12819,N_11901,N_11077);
xnor U12820 (N_12820,N_10639,N_11867);
xor U12821 (N_12821,N_10727,N_11986);
or U12822 (N_12822,N_10703,N_11640);
and U12823 (N_12823,N_11420,N_11277);
nand U12824 (N_12824,N_11430,N_11656);
xnor U12825 (N_12825,N_11763,N_10544);
nand U12826 (N_12826,N_10547,N_11212);
xnor U12827 (N_12827,N_11354,N_11355);
nand U12828 (N_12828,N_10760,N_10774);
nand U12829 (N_12829,N_11961,N_10757);
xnor U12830 (N_12830,N_11346,N_10766);
or U12831 (N_12831,N_10609,N_11741);
and U12832 (N_12832,N_11249,N_10844);
xnor U12833 (N_12833,N_11509,N_11419);
and U12834 (N_12834,N_11627,N_11366);
or U12835 (N_12835,N_11834,N_11064);
nor U12836 (N_12836,N_11447,N_11161);
and U12837 (N_12837,N_10559,N_10698);
nor U12838 (N_12838,N_11574,N_11498);
and U12839 (N_12839,N_11501,N_11908);
xor U12840 (N_12840,N_11586,N_11770);
xor U12841 (N_12841,N_10796,N_11233);
xnor U12842 (N_12842,N_11682,N_10902);
nor U12843 (N_12843,N_10974,N_11307);
xnor U12844 (N_12844,N_11111,N_10589);
nand U12845 (N_12845,N_10812,N_10642);
and U12846 (N_12846,N_11114,N_11294);
xnor U12847 (N_12847,N_11533,N_11143);
nand U12848 (N_12848,N_11442,N_11812);
nand U12849 (N_12849,N_11080,N_10806);
and U12850 (N_12850,N_11933,N_11467);
nand U12851 (N_12851,N_11091,N_11039);
or U12852 (N_12852,N_11083,N_11576);
nand U12853 (N_12853,N_11088,N_11026);
xnor U12854 (N_12854,N_10599,N_10692);
nand U12855 (N_12855,N_10769,N_11830);
or U12856 (N_12856,N_11629,N_11468);
nor U12857 (N_12857,N_10565,N_11249);
xnor U12858 (N_12858,N_10766,N_10658);
or U12859 (N_12859,N_11668,N_11002);
xor U12860 (N_12860,N_11532,N_11154);
nor U12861 (N_12861,N_10657,N_11216);
nand U12862 (N_12862,N_10709,N_11016);
nor U12863 (N_12863,N_11677,N_11729);
nor U12864 (N_12864,N_10547,N_10651);
nor U12865 (N_12865,N_10792,N_10644);
or U12866 (N_12866,N_10969,N_11978);
xnor U12867 (N_12867,N_11741,N_11682);
nor U12868 (N_12868,N_11289,N_11388);
and U12869 (N_12869,N_11720,N_11873);
and U12870 (N_12870,N_10884,N_10526);
nor U12871 (N_12871,N_10873,N_11589);
or U12872 (N_12872,N_11101,N_10858);
and U12873 (N_12873,N_10736,N_11594);
nand U12874 (N_12874,N_11893,N_10724);
nor U12875 (N_12875,N_11634,N_10502);
and U12876 (N_12876,N_10959,N_10803);
nor U12877 (N_12877,N_11011,N_10873);
nand U12878 (N_12878,N_10850,N_11920);
nand U12879 (N_12879,N_11535,N_11568);
nor U12880 (N_12880,N_10874,N_11585);
nand U12881 (N_12881,N_10751,N_11108);
xor U12882 (N_12882,N_11363,N_11235);
nor U12883 (N_12883,N_10914,N_11486);
and U12884 (N_12884,N_11441,N_10972);
xor U12885 (N_12885,N_11258,N_11498);
and U12886 (N_12886,N_11429,N_11383);
nand U12887 (N_12887,N_11814,N_11974);
xnor U12888 (N_12888,N_11527,N_11274);
and U12889 (N_12889,N_11034,N_11174);
or U12890 (N_12890,N_11337,N_11012);
and U12891 (N_12891,N_10515,N_10937);
and U12892 (N_12892,N_11476,N_10646);
or U12893 (N_12893,N_11368,N_10882);
xor U12894 (N_12894,N_10623,N_11580);
or U12895 (N_12895,N_11494,N_10906);
xor U12896 (N_12896,N_10502,N_10712);
nand U12897 (N_12897,N_11597,N_11724);
xnor U12898 (N_12898,N_11136,N_11323);
nand U12899 (N_12899,N_11696,N_11908);
xnor U12900 (N_12900,N_11239,N_11609);
nor U12901 (N_12901,N_11789,N_10927);
nor U12902 (N_12902,N_10768,N_11493);
nor U12903 (N_12903,N_10679,N_11822);
nor U12904 (N_12904,N_10513,N_11044);
xor U12905 (N_12905,N_11747,N_11820);
nor U12906 (N_12906,N_11364,N_11903);
nand U12907 (N_12907,N_11112,N_11727);
nor U12908 (N_12908,N_10541,N_11555);
nand U12909 (N_12909,N_10716,N_11120);
nor U12910 (N_12910,N_11077,N_10604);
nor U12911 (N_12911,N_10532,N_11373);
or U12912 (N_12912,N_10992,N_10699);
nor U12913 (N_12913,N_10912,N_11305);
nor U12914 (N_12914,N_11209,N_11310);
or U12915 (N_12915,N_11742,N_10587);
or U12916 (N_12916,N_11585,N_11888);
or U12917 (N_12917,N_11337,N_11324);
nand U12918 (N_12918,N_11565,N_11497);
xnor U12919 (N_12919,N_11269,N_11180);
nand U12920 (N_12920,N_11490,N_11827);
nor U12921 (N_12921,N_10522,N_11679);
nand U12922 (N_12922,N_11792,N_11785);
nand U12923 (N_12923,N_11830,N_11772);
nand U12924 (N_12924,N_11604,N_10896);
and U12925 (N_12925,N_11941,N_11383);
nand U12926 (N_12926,N_10505,N_10998);
nor U12927 (N_12927,N_11108,N_10690);
xor U12928 (N_12928,N_11423,N_11334);
nor U12929 (N_12929,N_11573,N_10780);
xnor U12930 (N_12930,N_10667,N_11942);
xor U12931 (N_12931,N_11794,N_11135);
or U12932 (N_12932,N_10863,N_10581);
nor U12933 (N_12933,N_10793,N_11043);
xnor U12934 (N_12934,N_10943,N_11706);
or U12935 (N_12935,N_11174,N_11802);
xnor U12936 (N_12936,N_11036,N_10933);
and U12937 (N_12937,N_10774,N_11961);
and U12938 (N_12938,N_11128,N_10661);
or U12939 (N_12939,N_11193,N_11877);
or U12940 (N_12940,N_11514,N_11027);
nor U12941 (N_12941,N_10552,N_11341);
nor U12942 (N_12942,N_11346,N_10519);
and U12943 (N_12943,N_11604,N_11613);
xor U12944 (N_12944,N_11550,N_11127);
nand U12945 (N_12945,N_11741,N_11599);
xor U12946 (N_12946,N_10995,N_10732);
or U12947 (N_12947,N_11870,N_11012);
nand U12948 (N_12948,N_10823,N_10763);
nand U12949 (N_12949,N_11800,N_11708);
xor U12950 (N_12950,N_10658,N_11928);
nor U12951 (N_12951,N_11636,N_10678);
xnor U12952 (N_12952,N_11488,N_11661);
or U12953 (N_12953,N_11102,N_10735);
xor U12954 (N_12954,N_11047,N_11569);
nor U12955 (N_12955,N_11427,N_11267);
nor U12956 (N_12956,N_10827,N_10892);
nand U12957 (N_12957,N_11818,N_11243);
or U12958 (N_12958,N_11279,N_10695);
and U12959 (N_12959,N_11108,N_11010);
nand U12960 (N_12960,N_11886,N_11347);
and U12961 (N_12961,N_10851,N_11812);
and U12962 (N_12962,N_11779,N_11220);
xnor U12963 (N_12963,N_10795,N_10583);
nor U12964 (N_12964,N_11005,N_11118);
nor U12965 (N_12965,N_11019,N_10632);
and U12966 (N_12966,N_11547,N_11371);
nor U12967 (N_12967,N_11862,N_10967);
or U12968 (N_12968,N_11390,N_10816);
nand U12969 (N_12969,N_11811,N_11229);
nor U12970 (N_12970,N_11781,N_11352);
and U12971 (N_12971,N_11947,N_10574);
xnor U12972 (N_12972,N_10692,N_10933);
xor U12973 (N_12973,N_10990,N_11239);
nor U12974 (N_12974,N_11893,N_11801);
nor U12975 (N_12975,N_11997,N_11406);
nor U12976 (N_12976,N_10621,N_10774);
nor U12977 (N_12977,N_10940,N_10547);
nor U12978 (N_12978,N_10981,N_11854);
nand U12979 (N_12979,N_11742,N_10588);
xor U12980 (N_12980,N_10996,N_11366);
and U12981 (N_12981,N_11636,N_11519);
or U12982 (N_12982,N_11992,N_11945);
nand U12983 (N_12983,N_10671,N_10517);
and U12984 (N_12984,N_11124,N_10558);
and U12985 (N_12985,N_10753,N_11629);
xnor U12986 (N_12986,N_11674,N_11640);
xnor U12987 (N_12987,N_11841,N_10676);
nand U12988 (N_12988,N_10548,N_11679);
nand U12989 (N_12989,N_11459,N_10677);
and U12990 (N_12990,N_10655,N_11494);
or U12991 (N_12991,N_11618,N_10617);
or U12992 (N_12992,N_10805,N_11712);
xor U12993 (N_12993,N_10669,N_10784);
nand U12994 (N_12994,N_10907,N_10943);
nand U12995 (N_12995,N_11892,N_10672);
nor U12996 (N_12996,N_11839,N_10712);
or U12997 (N_12997,N_11726,N_11014);
xnor U12998 (N_12998,N_11914,N_10658);
nor U12999 (N_12999,N_11380,N_11562);
xnor U13000 (N_13000,N_11759,N_11768);
nor U13001 (N_13001,N_11871,N_11272);
or U13002 (N_13002,N_10831,N_11044);
nand U13003 (N_13003,N_11895,N_11020);
nand U13004 (N_13004,N_11752,N_10622);
nor U13005 (N_13005,N_11429,N_11822);
or U13006 (N_13006,N_10635,N_11719);
nor U13007 (N_13007,N_10547,N_11629);
nor U13008 (N_13008,N_11012,N_11898);
or U13009 (N_13009,N_10582,N_11316);
xnor U13010 (N_13010,N_11450,N_11381);
or U13011 (N_13011,N_11543,N_10982);
nor U13012 (N_13012,N_11307,N_10938);
and U13013 (N_13013,N_10691,N_11527);
xor U13014 (N_13014,N_10576,N_10651);
and U13015 (N_13015,N_10747,N_11584);
or U13016 (N_13016,N_11959,N_11287);
nand U13017 (N_13017,N_11374,N_10690);
or U13018 (N_13018,N_10749,N_11798);
and U13019 (N_13019,N_10550,N_11652);
xnor U13020 (N_13020,N_11201,N_10933);
nor U13021 (N_13021,N_11507,N_10575);
or U13022 (N_13022,N_11500,N_11781);
xor U13023 (N_13023,N_11741,N_11832);
xnor U13024 (N_13024,N_11197,N_11880);
and U13025 (N_13025,N_10661,N_11846);
nor U13026 (N_13026,N_11357,N_11517);
or U13027 (N_13027,N_11835,N_11546);
and U13028 (N_13028,N_11444,N_11382);
nand U13029 (N_13029,N_11242,N_11817);
nor U13030 (N_13030,N_11037,N_11316);
nor U13031 (N_13031,N_11110,N_11862);
nand U13032 (N_13032,N_11143,N_11552);
and U13033 (N_13033,N_11192,N_10528);
nand U13034 (N_13034,N_10740,N_11409);
or U13035 (N_13035,N_10963,N_10602);
and U13036 (N_13036,N_10918,N_11255);
nand U13037 (N_13037,N_10862,N_10883);
nand U13038 (N_13038,N_11910,N_10957);
nand U13039 (N_13039,N_10684,N_11722);
xor U13040 (N_13040,N_11571,N_11390);
xnor U13041 (N_13041,N_10773,N_11661);
or U13042 (N_13042,N_10813,N_11143);
and U13043 (N_13043,N_10768,N_11679);
or U13044 (N_13044,N_11189,N_10971);
xor U13045 (N_13045,N_11243,N_10601);
xor U13046 (N_13046,N_11806,N_11166);
or U13047 (N_13047,N_10823,N_11918);
nand U13048 (N_13048,N_10931,N_11690);
or U13049 (N_13049,N_11855,N_11880);
or U13050 (N_13050,N_11342,N_11375);
nand U13051 (N_13051,N_11226,N_10751);
nand U13052 (N_13052,N_10812,N_10811);
xnor U13053 (N_13053,N_11745,N_11188);
nand U13054 (N_13054,N_10642,N_10595);
and U13055 (N_13055,N_11510,N_10878);
nand U13056 (N_13056,N_10765,N_11305);
and U13057 (N_13057,N_11359,N_11367);
nor U13058 (N_13058,N_11435,N_10614);
and U13059 (N_13059,N_11608,N_11124);
xor U13060 (N_13060,N_11716,N_11821);
or U13061 (N_13061,N_11737,N_11893);
nor U13062 (N_13062,N_10852,N_11444);
and U13063 (N_13063,N_11936,N_11534);
and U13064 (N_13064,N_11165,N_11871);
and U13065 (N_13065,N_11847,N_11478);
nor U13066 (N_13066,N_11940,N_11154);
nand U13067 (N_13067,N_11752,N_11824);
nor U13068 (N_13068,N_11692,N_11839);
xnor U13069 (N_13069,N_11914,N_11756);
xnor U13070 (N_13070,N_11072,N_11343);
xor U13071 (N_13071,N_11624,N_10695);
nand U13072 (N_13072,N_11157,N_11811);
nor U13073 (N_13073,N_11909,N_11362);
and U13074 (N_13074,N_11043,N_11680);
xor U13075 (N_13075,N_10723,N_11300);
nand U13076 (N_13076,N_11220,N_11851);
xor U13077 (N_13077,N_10575,N_11649);
nor U13078 (N_13078,N_10580,N_11667);
or U13079 (N_13079,N_10915,N_11042);
nand U13080 (N_13080,N_11081,N_11365);
xor U13081 (N_13081,N_11724,N_10637);
nand U13082 (N_13082,N_10810,N_10864);
xnor U13083 (N_13083,N_11673,N_10844);
or U13084 (N_13084,N_11996,N_11648);
nand U13085 (N_13085,N_10568,N_10534);
nand U13086 (N_13086,N_11826,N_11621);
nand U13087 (N_13087,N_10796,N_11220);
xor U13088 (N_13088,N_11177,N_11042);
xnor U13089 (N_13089,N_11052,N_11725);
and U13090 (N_13090,N_10896,N_10990);
xnor U13091 (N_13091,N_11057,N_10947);
nor U13092 (N_13092,N_11554,N_10576);
and U13093 (N_13093,N_10558,N_10848);
nand U13094 (N_13094,N_10565,N_10568);
and U13095 (N_13095,N_11880,N_11259);
nor U13096 (N_13096,N_11012,N_11152);
xor U13097 (N_13097,N_11355,N_11587);
xnor U13098 (N_13098,N_11057,N_10787);
or U13099 (N_13099,N_11685,N_11107);
xor U13100 (N_13100,N_11573,N_10666);
nor U13101 (N_13101,N_11211,N_10654);
nand U13102 (N_13102,N_10989,N_11836);
xor U13103 (N_13103,N_11384,N_10719);
nand U13104 (N_13104,N_11702,N_10958);
and U13105 (N_13105,N_11487,N_11328);
nand U13106 (N_13106,N_11804,N_11484);
nor U13107 (N_13107,N_11419,N_11954);
nand U13108 (N_13108,N_10785,N_11997);
xnor U13109 (N_13109,N_10527,N_11700);
nand U13110 (N_13110,N_10629,N_11389);
or U13111 (N_13111,N_11720,N_11537);
and U13112 (N_13112,N_10780,N_10845);
or U13113 (N_13113,N_11061,N_10547);
xor U13114 (N_13114,N_11847,N_11124);
xnor U13115 (N_13115,N_11320,N_11018);
nor U13116 (N_13116,N_10532,N_11705);
nor U13117 (N_13117,N_11216,N_10501);
and U13118 (N_13118,N_11233,N_11511);
nand U13119 (N_13119,N_10616,N_11884);
nand U13120 (N_13120,N_11812,N_11063);
nand U13121 (N_13121,N_11714,N_11370);
nand U13122 (N_13122,N_11249,N_10922);
nor U13123 (N_13123,N_11247,N_11472);
and U13124 (N_13124,N_11995,N_11317);
xor U13125 (N_13125,N_11193,N_11848);
nand U13126 (N_13126,N_11002,N_11049);
nor U13127 (N_13127,N_11481,N_11534);
xor U13128 (N_13128,N_10566,N_11988);
xnor U13129 (N_13129,N_10911,N_10807);
xnor U13130 (N_13130,N_11040,N_11156);
xor U13131 (N_13131,N_11332,N_11344);
xor U13132 (N_13132,N_11118,N_11157);
or U13133 (N_13133,N_11841,N_11680);
nand U13134 (N_13134,N_11599,N_10698);
xor U13135 (N_13135,N_10675,N_11630);
nor U13136 (N_13136,N_11165,N_11620);
nand U13137 (N_13137,N_10598,N_10517);
or U13138 (N_13138,N_10815,N_10677);
xor U13139 (N_13139,N_11308,N_10728);
or U13140 (N_13140,N_11841,N_10659);
nand U13141 (N_13141,N_11304,N_10664);
nand U13142 (N_13142,N_10924,N_10948);
and U13143 (N_13143,N_10905,N_10862);
and U13144 (N_13144,N_11875,N_10608);
and U13145 (N_13145,N_11906,N_11449);
and U13146 (N_13146,N_11218,N_11088);
xor U13147 (N_13147,N_11526,N_11859);
or U13148 (N_13148,N_10982,N_11005);
and U13149 (N_13149,N_11043,N_11685);
nor U13150 (N_13150,N_11450,N_10881);
xnor U13151 (N_13151,N_11234,N_11075);
nand U13152 (N_13152,N_11051,N_11863);
xnor U13153 (N_13153,N_11980,N_11668);
nor U13154 (N_13154,N_10820,N_10882);
nor U13155 (N_13155,N_11445,N_11813);
nor U13156 (N_13156,N_11781,N_11822);
or U13157 (N_13157,N_11801,N_10754);
xor U13158 (N_13158,N_11973,N_10987);
and U13159 (N_13159,N_11744,N_11541);
or U13160 (N_13160,N_11851,N_10869);
xor U13161 (N_13161,N_10710,N_10953);
or U13162 (N_13162,N_10531,N_10700);
and U13163 (N_13163,N_11942,N_11340);
nor U13164 (N_13164,N_11843,N_11415);
and U13165 (N_13165,N_11809,N_10859);
or U13166 (N_13166,N_11261,N_11234);
xor U13167 (N_13167,N_11568,N_11617);
nor U13168 (N_13168,N_11923,N_11330);
nand U13169 (N_13169,N_11951,N_11097);
or U13170 (N_13170,N_11589,N_11912);
nand U13171 (N_13171,N_11108,N_11136);
nand U13172 (N_13172,N_11482,N_11651);
nor U13173 (N_13173,N_11143,N_11576);
or U13174 (N_13174,N_11707,N_11366);
and U13175 (N_13175,N_11588,N_10832);
nand U13176 (N_13176,N_10898,N_10859);
nand U13177 (N_13177,N_10878,N_11166);
and U13178 (N_13178,N_10745,N_11195);
xnor U13179 (N_13179,N_11672,N_10576);
nor U13180 (N_13180,N_11493,N_11009);
nand U13181 (N_13181,N_11525,N_11450);
xnor U13182 (N_13182,N_11304,N_10788);
and U13183 (N_13183,N_11007,N_11343);
nand U13184 (N_13184,N_11999,N_10899);
and U13185 (N_13185,N_11920,N_11534);
and U13186 (N_13186,N_11454,N_11978);
or U13187 (N_13187,N_11503,N_11197);
nand U13188 (N_13188,N_11754,N_11247);
xor U13189 (N_13189,N_11926,N_10956);
xor U13190 (N_13190,N_10975,N_10954);
or U13191 (N_13191,N_11288,N_11381);
and U13192 (N_13192,N_11243,N_10920);
nand U13193 (N_13193,N_11755,N_11920);
nand U13194 (N_13194,N_11921,N_11632);
xor U13195 (N_13195,N_11323,N_10943);
nand U13196 (N_13196,N_10693,N_10615);
and U13197 (N_13197,N_10754,N_11340);
nand U13198 (N_13198,N_10937,N_10890);
nor U13199 (N_13199,N_11537,N_10776);
nand U13200 (N_13200,N_10677,N_11707);
nand U13201 (N_13201,N_11932,N_11148);
nor U13202 (N_13202,N_10579,N_10748);
nand U13203 (N_13203,N_11897,N_10611);
or U13204 (N_13204,N_10975,N_11979);
nor U13205 (N_13205,N_11415,N_10501);
nand U13206 (N_13206,N_10633,N_11376);
and U13207 (N_13207,N_11322,N_11206);
xnor U13208 (N_13208,N_11055,N_11529);
xnor U13209 (N_13209,N_11041,N_11205);
and U13210 (N_13210,N_10931,N_10865);
xnor U13211 (N_13211,N_11196,N_11389);
nor U13212 (N_13212,N_10543,N_11459);
nor U13213 (N_13213,N_11454,N_11148);
nand U13214 (N_13214,N_10566,N_11127);
and U13215 (N_13215,N_10737,N_10952);
nor U13216 (N_13216,N_10985,N_10640);
nor U13217 (N_13217,N_11809,N_11730);
nor U13218 (N_13218,N_11103,N_10916);
xor U13219 (N_13219,N_11503,N_11775);
nor U13220 (N_13220,N_11938,N_11181);
nor U13221 (N_13221,N_11495,N_10967);
xor U13222 (N_13222,N_10562,N_11720);
nor U13223 (N_13223,N_11455,N_11483);
or U13224 (N_13224,N_10941,N_10658);
xnor U13225 (N_13225,N_11768,N_11283);
and U13226 (N_13226,N_10893,N_11671);
xnor U13227 (N_13227,N_11109,N_11108);
nor U13228 (N_13228,N_11049,N_11227);
nor U13229 (N_13229,N_11296,N_11246);
or U13230 (N_13230,N_10635,N_11531);
xor U13231 (N_13231,N_10987,N_11875);
or U13232 (N_13232,N_11788,N_11049);
and U13233 (N_13233,N_10841,N_11284);
nand U13234 (N_13234,N_11908,N_11147);
nor U13235 (N_13235,N_11432,N_11399);
nor U13236 (N_13236,N_11548,N_11945);
nor U13237 (N_13237,N_11012,N_11527);
nor U13238 (N_13238,N_10919,N_11758);
nand U13239 (N_13239,N_11870,N_11032);
xor U13240 (N_13240,N_10563,N_11941);
nor U13241 (N_13241,N_11022,N_11321);
and U13242 (N_13242,N_11054,N_11707);
nor U13243 (N_13243,N_11697,N_11133);
xnor U13244 (N_13244,N_11154,N_11256);
nand U13245 (N_13245,N_11584,N_11573);
nor U13246 (N_13246,N_11606,N_11656);
nand U13247 (N_13247,N_11111,N_11910);
nor U13248 (N_13248,N_10588,N_11425);
or U13249 (N_13249,N_11021,N_11436);
xnor U13250 (N_13250,N_11523,N_10804);
nand U13251 (N_13251,N_11192,N_10783);
and U13252 (N_13252,N_11950,N_11468);
xnor U13253 (N_13253,N_11066,N_10732);
nand U13254 (N_13254,N_11191,N_11352);
and U13255 (N_13255,N_11555,N_11043);
nor U13256 (N_13256,N_11563,N_11320);
or U13257 (N_13257,N_11542,N_11659);
xor U13258 (N_13258,N_10574,N_11968);
xnor U13259 (N_13259,N_11095,N_11661);
xor U13260 (N_13260,N_11901,N_11053);
or U13261 (N_13261,N_11808,N_10751);
or U13262 (N_13262,N_11994,N_11833);
and U13263 (N_13263,N_11685,N_10549);
nand U13264 (N_13264,N_11427,N_11358);
xnor U13265 (N_13265,N_10954,N_10503);
xor U13266 (N_13266,N_11627,N_11339);
nand U13267 (N_13267,N_11798,N_11085);
nand U13268 (N_13268,N_11120,N_11788);
or U13269 (N_13269,N_10792,N_10790);
or U13270 (N_13270,N_11304,N_10821);
and U13271 (N_13271,N_11488,N_11195);
nor U13272 (N_13272,N_11858,N_10667);
nand U13273 (N_13273,N_11811,N_11498);
nand U13274 (N_13274,N_11415,N_11478);
or U13275 (N_13275,N_10886,N_11273);
and U13276 (N_13276,N_10947,N_11188);
xnor U13277 (N_13277,N_10748,N_11231);
nand U13278 (N_13278,N_11651,N_10576);
nand U13279 (N_13279,N_11104,N_11149);
or U13280 (N_13280,N_10746,N_11192);
and U13281 (N_13281,N_11407,N_11144);
and U13282 (N_13282,N_11769,N_11732);
or U13283 (N_13283,N_11795,N_10602);
and U13284 (N_13284,N_11663,N_10772);
xor U13285 (N_13285,N_11685,N_11806);
xor U13286 (N_13286,N_11493,N_11715);
or U13287 (N_13287,N_11900,N_11297);
nand U13288 (N_13288,N_11678,N_10859);
nand U13289 (N_13289,N_11402,N_10829);
and U13290 (N_13290,N_10906,N_10864);
nand U13291 (N_13291,N_11172,N_11092);
nand U13292 (N_13292,N_11336,N_11207);
xnor U13293 (N_13293,N_11123,N_11663);
or U13294 (N_13294,N_11182,N_11697);
and U13295 (N_13295,N_11541,N_11828);
and U13296 (N_13296,N_10872,N_11276);
and U13297 (N_13297,N_11142,N_11777);
nor U13298 (N_13298,N_11480,N_10682);
nand U13299 (N_13299,N_11706,N_11432);
or U13300 (N_13300,N_11837,N_11918);
xnor U13301 (N_13301,N_11376,N_11065);
xnor U13302 (N_13302,N_10860,N_10896);
or U13303 (N_13303,N_11912,N_11031);
or U13304 (N_13304,N_10818,N_10514);
xnor U13305 (N_13305,N_11067,N_10837);
nor U13306 (N_13306,N_11362,N_10790);
or U13307 (N_13307,N_10994,N_11328);
and U13308 (N_13308,N_10641,N_11541);
nor U13309 (N_13309,N_11921,N_11989);
nor U13310 (N_13310,N_10913,N_11534);
nand U13311 (N_13311,N_11410,N_10791);
nor U13312 (N_13312,N_10913,N_10931);
nor U13313 (N_13313,N_10555,N_11339);
or U13314 (N_13314,N_10665,N_11075);
or U13315 (N_13315,N_11564,N_11862);
nor U13316 (N_13316,N_11991,N_11457);
xnor U13317 (N_13317,N_11400,N_11165);
and U13318 (N_13318,N_10677,N_11397);
and U13319 (N_13319,N_11022,N_10569);
nor U13320 (N_13320,N_10769,N_11874);
nor U13321 (N_13321,N_11759,N_10877);
nor U13322 (N_13322,N_10883,N_11386);
or U13323 (N_13323,N_10595,N_11407);
nor U13324 (N_13324,N_11382,N_11793);
nor U13325 (N_13325,N_11392,N_11623);
xor U13326 (N_13326,N_11397,N_11468);
nand U13327 (N_13327,N_10617,N_11815);
xor U13328 (N_13328,N_10608,N_10590);
or U13329 (N_13329,N_11390,N_11634);
and U13330 (N_13330,N_11491,N_11433);
nor U13331 (N_13331,N_11591,N_11932);
or U13332 (N_13332,N_11267,N_11841);
nand U13333 (N_13333,N_11244,N_10988);
or U13334 (N_13334,N_11175,N_11904);
nor U13335 (N_13335,N_10941,N_10587);
nor U13336 (N_13336,N_10711,N_11285);
xnor U13337 (N_13337,N_10879,N_11099);
nand U13338 (N_13338,N_10912,N_11714);
nor U13339 (N_13339,N_11928,N_10516);
and U13340 (N_13340,N_10903,N_11701);
nor U13341 (N_13341,N_11692,N_10537);
or U13342 (N_13342,N_10867,N_10984);
xor U13343 (N_13343,N_11069,N_11000);
or U13344 (N_13344,N_11573,N_11404);
and U13345 (N_13345,N_10518,N_11010);
nor U13346 (N_13346,N_10614,N_10584);
nor U13347 (N_13347,N_10520,N_10538);
xor U13348 (N_13348,N_11011,N_10998);
nor U13349 (N_13349,N_11859,N_10684);
nor U13350 (N_13350,N_11943,N_11945);
or U13351 (N_13351,N_10713,N_11884);
nor U13352 (N_13352,N_11370,N_10620);
xor U13353 (N_13353,N_10784,N_11384);
nand U13354 (N_13354,N_11093,N_11220);
nor U13355 (N_13355,N_10729,N_11696);
nand U13356 (N_13356,N_11101,N_10588);
and U13357 (N_13357,N_11883,N_11230);
nand U13358 (N_13358,N_11260,N_11055);
nand U13359 (N_13359,N_11196,N_11425);
xor U13360 (N_13360,N_11428,N_11205);
nor U13361 (N_13361,N_10730,N_11795);
and U13362 (N_13362,N_10913,N_11871);
nor U13363 (N_13363,N_11790,N_11597);
xor U13364 (N_13364,N_11540,N_10652);
xor U13365 (N_13365,N_10975,N_11198);
xnor U13366 (N_13366,N_11426,N_11922);
or U13367 (N_13367,N_11417,N_11244);
nand U13368 (N_13368,N_11172,N_11502);
or U13369 (N_13369,N_10825,N_10694);
nor U13370 (N_13370,N_10810,N_10515);
nor U13371 (N_13371,N_10777,N_11212);
xnor U13372 (N_13372,N_10743,N_11487);
xnor U13373 (N_13373,N_11312,N_11307);
nor U13374 (N_13374,N_11202,N_10631);
xnor U13375 (N_13375,N_10709,N_11827);
nor U13376 (N_13376,N_11170,N_10540);
and U13377 (N_13377,N_11497,N_10946);
nor U13378 (N_13378,N_10690,N_10663);
xnor U13379 (N_13379,N_11871,N_11720);
and U13380 (N_13380,N_11778,N_11905);
nor U13381 (N_13381,N_11590,N_10919);
xnor U13382 (N_13382,N_11551,N_11117);
nor U13383 (N_13383,N_11016,N_11208);
xnor U13384 (N_13384,N_11671,N_11155);
nor U13385 (N_13385,N_11699,N_11295);
and U13386 (N_13386,N_10531,N_11949);
nand U13387 (N_13387,N_11444,N_11187);
nor U13388 (N_13388,N_10653,N_11142);
or U13389 (N_13389,N_10696,N_10961);
and U13390 (N_13390,N_11504,N_10687);
xor U13391 (N_13391,N_11596,N_11289);
nand U13392 (N_13392,N_10950,N_11833);
and U13393 (N_13393,N_10974,N_10976);
or U13394 (N_13394,N_10508,N_10588);
xnor U13395 (N_13395,N_10554,N_11877);
or U13396 (N_13396,N_10888,N_11390);
and U13397 (N_13397,N_11180,N_10556);
xor U13398 (N_13398,N_11003,N_11675);
and U13399 (N_13399,N_11039,N_10984);
or U13400 (N_13400,N_11177,N_10740);
nor U13401 (N_13401,N_11237,N_11053);
or U13402 (N_13402,N_11252,N_11540);
nor U13403 (N_13403,N_10516,N_10532);
xnor U13404 (N_13404,N_10879,N_11073);
nor U13405 (N_13405,N_11671,N_11079);
xor U13406 (N_13406,N_11312,N_11869);
nor U13407 (N_13407,N_10838,N_10677);
xor U13408 (N_13408,N_11187,N_11327);
and U13409 (N_13409,N_10848,N_10573);
nand U13410 (N_13410,N_10607,N_11654);
or U13411 (N_13411,N_11630,N_11857);
or U13412 (N_13412,N_11314,N_11339);
or U13413 (N_13413,N_10897,N_11563);
nor U13414 (N_13414,N_11129,N_11435);
nor U13415 (N_13415,N_10561,N_11576);
xnor U13416 (N_13416,N_10621,N_10833);
and U13417 (N_13417,N_11337,N_11150);
nor U13418 (N_13418,N_11392,N_11291);
xor U13419 (N_13419,N_10993,N_10641);
xor U13420 (N_13420,N_10626,N_11461);
or U13421 (N_13421,N_11646,N_11043);
and U13422 (N_13422,N_11808,N_11358);
or U13423 (N_13423,N_11176,N_11673);
or U13424 (N_13424,N_11161,N_11133);
and U13425 (N_13425,N_11091,N_10571);
or U13426 (N_13426,N_10990,N_11454);
nand U13427 (N_13427,N_10722,N_11754);
nor U13428 (N_13428,N_11078,N_10513);
or U13429 (N_13429,N_10920,N_10878);
or U13430 (N_13430,N_10559,N_10897);
or U13431 (N_13431,N_11732,N_11054);
nand U13432 (N_13432,N_11025,N_10968);
or U13433 (N_13433,N_11251,N_10757);
and U13434 (N_13434,N_11674,N_10853);
xor U13435 (N_13435,N_11805,N_11425);
and U13436 (N_13436,N_11775,N_10548);
xor U13437 (N_13437,N_10890,N_10919);
xor U13438 (N_13438,N_10659,N_10918);
nand U13439 (N_13439,N_10953,N_11024);
nor U13440 (N_13440,N_11392,N_11463);
nand U13441 (N_13441,N_10546,N_11403);
and U13442 (N_13442,N_10717,N_10522);
xor U13443 (N_13443,N_10698,N_11417);
or U13444 (N_13444,N_10990,N_10941);
and U13445 (N_13445,N_10798,N_10840);
and U13446 (N_13446,N_10652,N_11346);
nand U13447 (N_13447,N_10949,N_10975);
nor U13448 (N_13448,N_11238,N_11861);
or U13449 (N_13449,N_11444,N_11857);
and U13450 (N_13450,N_11844,N_10960);
and U13451 (N_13451,N_11776,N_11315);
or U13452 (N_13452,N_11638,N_10693);
nor U13453 (N_13453,N_11494,N_10661);
and U13454 (N_13454,N_10652,N_11902);
nand U13455 (N_13455,N_11179,N_10920);
and U13456 (N_13456,N_11225,N_10961);
nor U13457 (N_13457,N_10912,N_11609);
or U13458 (N_13458,N_10837,N_10836);
nor U13459 (N_13459,N_11073,N_11297);
or U13460 (N_13460,N_11008,N_11495);
nand U13461 (N_13461,N_11576,N_10908);
xor U13462 (N_13462,N_11485,N_10846);
nor U13463 (N_13463,N_11153,N_11072);
or U13464 (N_13464,N_11857,N_11668);
and U13465 (N_13465,N_11640,N_10772);
xnor U13466 (N_13466,N_10835,N_11094);
and U13467 (N_13467,N_11488,N_11375);
and U13468 (N_13468,N_11115,N_11790);
and U13469 (N_13469,N_11127,N_10733);
nor U13470 (N_13470,N_10530,N_11444);
and U13471 (N_13471,N_11294,N_11180);
nor U13472 (N_13472,N_11355,N_10945);
and U13473 (N_13473,N_11535,N_11926);
nand U13474 (N_13474,N_10937,N_11816);
and U13475 (N_13475,N_10504,N_11366);
or U13476 (N_13476,N_10796,N_10577);
and U13477 (N_13477,N_10688,N_10848);
or U13478 (N_13478,N_11913,N_11004);
nor U13479 (N_13479,N_11163,N_11583);
nand U13480 (N_13480,N_11720,N_10591);
xnor U13481 (N_13481,N_11221,N_11102);
nand U13482 (N_13482,N_11209,N_11870);
xnor U13483 (N_13483,N_11837,N_10915);
and U13484 (N_13484,N_10704,N_11228);
xor U13485 (N_13485,N_11716,N_11322);
and U13486 (N_13486,N_11787,N_11650);
nand U13487 (N_13487,N_11017,N_11960);
xnor U13488 (N_13488,N_10944,N_11791);
or U13489 (N_13489,N_11555,N_10847);
nor U13490 (N_13490,N_10780,N_10621);
xor U13491 (N_13491,N_10580,N_10514);
and U13492 (N_13492,N_10857,N_11118);
xor U13493 (N_13493,N_10777,N_11997);
nand U13494 (N_13494,N_11366,N_11984);
xnor U13495 (N_13495,N_11896,N_10640);
and U13496 (N_13496,N_10534,N_10698);
and U13497 (N_13497,N_11406,N_11044);
xor U13498 (N_13498,N_10718,N_11580);
xnor U13499 (N_13499,N_10530,N_11343);
or U13500 (N_13500,N_13264,N_12083);
xor U13501 (N_13501,N_12274,N_12381);
or U13502 (N_13502,N_12774,N_12717);
or U13503 (N_13503,N_12510,N_12435);
nor U13504 (N_13504,N_13328,N_12447);
nand U13505 (N_13505,N_13291,N_12764);
nor U13506 (N_13506,N_13426,N_12310);
and U13507 (N_13507,N_12414,N_13229);
nand U13508 (N_13508,N_12626,N_12410);
xnor U13509 (N_13509,N_12289,N_13466);
nand U13510 (N_13510,N_13339,N_13020);
nand U13511 (N_13511,N_13434,N_12632);
nor U13512 (N_13512,N_12538,N_12411);
and U13513 (N_13513,N_12944,N_13416);
nor U13514 (N_13514,N_13216,N_12400);
and U13515 (N_13515,N_12174,N_12208);
and U13516 (N_13516,N_13159,N_12919);
xor U13517 (N_13517,N_12317,N_12228);
nor U13518 (N_13518,N_13385,N_13178);
xnor U13519 (N_13519,N_13032,N_13236);
xor U13520 (N_13520,N_12288,N_13322);
and U13521 (N_13521,N_13183,N_12389);
xor U13522 (N_13522,N_12280,N_12456);
xnor U13523 (N_13523,N_12111,N_12459);
and U13524 (N_13524,N_12155,N_12143);
nor U13525 (N_13525,N_12494,N_12258);
xnor U13526 (N_13526,N_12725,N_12253);
nor U13527 (N_13527,N_12245,N_12238);
or U13528 (N_13528,N_13153,N_12776);
and U13529 (N_13529,N_12360,N_13070);
nor U13530 (N_13530,N_13030,N_13366);
xor U13531 (N_13531,N_13173,N_12067);
or U13532 (N_13532,N_12606,N_12285);
or U13533 (N_13533,N_12800,N_12276);
xor U13534 (N_13534,N_13319,N_13223);
xor U13535 (N_13535,N_12221,N_13083);
xor U13536 (N_13536,N_12858,N_13053);
nand U13537 (N_13537,N_12380,N_12949);
nand U13538 (N_13538,N_12209,N_12295);
nor U13539 (N_13539,N_13448,N_12882);
nand U13540 (N_13540,N_12860,N_12145);
nand U13541 (N_13541,N_13078,N_12242);
or U13542 (N_13542,N_13072,N_13330);
nand U13543 (N_13543,N_13482,N_12893);
and U13544 (N_13544,N_12149,N_13082);
nand U13545 (N_13545,N_12779,N_13058);
and U13546 (N_13546,N_12850,N_12146);
xor U13547 (N_13547,N_12994,N_13429);
nand U13548 (N_13548,N_13498,N_13338);
nand U13549 (N_13549,N_13002,N_12681);
and U13550 (N_13550,N_12403,N_12487);
or U13551 (N_13551,N_12361,N_12333);
nor U13552 (N_13552,N_13294,N_12399);
or U13553 (N_13553,N_12071,N_12402);
nor U13554 (N_13554,N_12485,N_12051);
nor U13555 (N_13555,N_12337,N_12202);
nor U13556 (N_13556,N_12785,N_12345);
xnor U13557 (N_13557,N_12767,N_13023);
nor U13558 (N_13558,N_12680,N_13104);
nor U13559 (N_13559,N_13101,N_12152);
nor U13560 (N_13560,N_13077,N_12637);
and U13561 (N_13561,N_12002,N_12303);
nor U13562 (N_13562,N_12819,N_12495);
nand U13563 (N_13563,N_12147,N_12124);
xor U13564 (N_13564,N_13048,N_12529);
and U13565 (N_13565,N_12598,N_12840);
and U13566 (N_13566,N_12019,N_13487);
xnor U13567 (N_13567,N_12406,N_12112);
nor U13568 (N_13568,N_13379,N_12913);
xor U13569 (N_13569,N_12079,N_12206);
or U13570 (N_13570,N_13421,N_12102);
nand U13571 (N_13571,N_13103,N_12896);
nor U13572 (N_13572,N_12237,N_12169);
nand U13573 (N_13573,N_12477,N_12788);
and U13574 (N_13574,N_12772,N_12533);
nor U13575 (N_13575,N_12607,N_12682);
or U13576 (N_13576,N_12951,N_12508);
nand U13577 (N_13577,N_13118,N_12679);
and U13578 (N_13578,N_12687,N_12325);
xnor U13579 (N_13579,N_12297,N_12318);
or U13580 (N_13580,N_13222,N_12883);
nand U13581 (N_13581,N_12105,N_12639);
nor U13582 (N_13582,N_12790,N_13239);
nor U13583 (N_13583,N_12877,N_12178);
and U13584 (N_13584,N_13261,N_13478);
nand U13585 (N_13585,N_12960,N_13361);
nor U13586 (N_13586,N_13389,N_12955);
and U13587 (N_13587,N_12287,N_12600);
xnor U13588 (N_13588,N_12300,N_12664);
nand U13589 (N_13589,N_12195,N_12012);
nor U13590 (N_13590,N_13255,N_12670);
or U13591 (N_13591,N_12186,N_13475);
nor U13592 (N_13592,N_13213,N_13484);
or U13593 (N_13593,N_12476,N_12142);
xnor U13594 (N_13594,N_13189,N_12007);
or U13595 (N_13595,N_12873,N_12677);
nand U13596 (N_13596,N_13408,N_13022);
nand U13597 (N_13597,N_13457,N_12044);
nand U13598 (N_13598,N_13311,N_12291);
nor U13599 (N_13599,N_12685,N_12610);
nand U13600 (N_13600,N_13370,N_12552);
nand U13601 (N_13601,N_12698,N_13026);
xor U13602 (N_13602,N_12507,N_12353);
and U13603 (N_13603,N_12379,N_13432);
nand U13604 (N_13604,N_13157,N_13374);
nand U13605 (N_13605,N_12842,N_12290);
and U13606 (N_13606,N_13332,N_13262);
xor U13607 (N_13607,N_13209,N_12281);
and U13608 (N_13608,N_13350,N_13220);
nand U13609 (N_13609,N_13211,N_13152);
nor U13610 (N_13610,N_13035,N_12128);
xnor U13611 (N_13611,N_13177,N_12993);
and U13612 (N_13612,N_13165,N_12780);
or U13613 (N_13613,N_13259,N_12879);
xor U13614 (N_13614,N_12423,N_12009);
nand U13615 (N_13615,N_12967,N_12453);
nor U13616 (N_13616,N_13176,N_12176);
nand U13617 (N_13617,N_13451,N_12702);
nor U13618 (N_13618,N_12961,N_12984);
and U13619 (N_13619,N_12871,N_13256);
nor U13620 (N_13620,N_12455,N_13212);
or U13621 (N_13621,N_12348,N_12557);
xnor U13622 (N_13622,N_13100,N_13201);
or U13623 (N_13623,N_12065,N_12577);
nand U13624 (N_13624,N_13453,N_12405);
or U13625 (N_13625,N_12084,N_12123);
nor U13626 (N_13626,N_12052,N_13156);
and U13627 (N_13627,N_12540,N_12060);
nor U13628 (N_13628,N_12544,N_12746);
and U13629 (N_13629,N_12366,N_12829);
or U13630 (N_13630,N_12415,N_13476);
nor U13631 (N_13631,N_12104,N_12101);
nand U13632 (N_13632,N_13348,N_12810);
and U13633 (N_13633,N_12900,N_13033);
nor U13634 (N_13634,N_12426,N_12865);
xnor U13635 (N_13635,N_12099,N_12575);
or U13636 (N_13636,N_13192,N_12103);
xnor U13637 (N_13637,N_13489,N_12728);
nand U13638 (N_13638,N_12620,N_12897);
xnor U13639 (N_13639,N_12642,N_12196);
xor U13640 (N_13640,N_12587,N_12975);
nand U13641 (N_13641,N_13093,N_12823);
nor U13642 (N_13642,N_13198,N_12046);
nand U13643 (N_13643,N_12266,N_13166);
or U13644 (N_13644,N_12981,N_13283);
xor U13645 (N_13645,N_12581,N_12255);
nand U13646 (N_13646,N_13321,N_12837);
or U13647 (N_13647,N_13135,N_12923);
nand U13648 (N_13648,N_12753,N_13267);
nand U13649 (N_13649,N_13123,N_13195);
nor U13650 (N_13650,N_12458,N_12054);
and U13651 (N_13651,N_12811,N_13430);
nand U13652 (N_13652,N_12501,N_12603);
nand U13653 (N_13653,N_12938,N_12653);
xor U13654 (N_13654,N_13386,N_12230);
xor U13655 (N_13655,N_12576,N_12484);
nor U13656 (N_13656,N_12601,N_13074);
and U13657 (N_13657,N_12787,N_12250);
or U13658 (N_13658,N_12945,N_12356);
or U13659 (N_13659,N_13175,N_13092);
or U13660 (N_13660,N_12542,N_13493);
nor U13661 (N_13661,N_12828,N_13016);
nand U13662 (N_13662,N_12489,N_13240);
nor U13663 (N_13663,N_12541,N_12891);
nor U13664 (N_13664,N_12995,N_12008);
and U13665 (N_13665,N_12134,N_12931);
nand U13666 (N_13666,N_13019,N_12590);
or U13667 (N_13667,N_13293,N_12889);
and U13668 (N_13668,N_13280,N_13237);
nor U13669 (N_13669,N_12856,N_13423);
xor U13670 (N_13670,N_12796,N_12969);
nand U13671 (N_13671,N_12109,N_12032);
nand U13672 (N_13672,N_12985,N_13233);
xor U13673 (N_13673,N_12806,N_12370);
or U13674 (N_13674,N_12964,N_12049);
xnor U13675 (N_13675,N_12390,N_12699);
nand U13676 (N_13676,N_13433,N_12661);
nand U13677 (N_13677,N_12409,N_12886);
nor U13678 (N_13678,N_13472,N_13396);
xor U13679 (N_13679,N_13214,N_12132);
and U13680 (N_13680,N_12096,N_12383);
nor U13681 (N_13681,N_13288,N_12346);
xnor U13682 (N_13682,N_12254,N_12205);
or U13683 (N_13683,N_13308,N_13431);
nor U13684 (N_13684,N_12768,N_12910);
and U13685 (N_13685,N_12907,N_13499);
xnor U13686 (N_13686,N_12497,N_12652);
nor U13687 (N_13687,N_12614,N_12732);
nand U13688 (N_13688,N_13226,N_12398);
nor U13689 (N_13689,N_12983,N_12619);
nor U13690 (N_13690,N_12941,N_13044);
or U13691 (N_13691,N_13064,N_12222);
nand U13692 (N_13692,N_12125,N_13090);
and U13693 (N_13693,N_13352,N_12420);
or U13694 (N_13694,N_12773,N_13008);
xor U13695 (N_13695,N_12150,N_12613);
nand U13696 (N_13696,N_13485,N_12988);
and U13697 (N_13697,N_12180,N_12665);
xnor U13698 (N_13698,N_13184,N_12056);
nor U13699 (N_13699,N_12277,N_13272);
nor U13700 (N_13700,N_12997,N_13474);
nor U13701 (N_13701,N_12836,N_12211);
or U13702 (N_13702,N_12734,N_12674);
or U13703 (N_13703,N_12043,N_12956);
or U13704 (N_13704,N_12093,N_13113);
nand U13705 (N_13705,N_12880,N_12121);
and U13706 (N_13706,N_12094,N_13479);
xnor U13707 (N_13707,N_13425,N_12513);
nand U13708 (N_13708,N_13012,N_12991);
or U13709 (N_13709,N_12187,N_12010);
xnor U13710 (N_13710,N_12654,N_13017);
xor U13711 (N_13711,N_13144,N_12504);
or U13712 (N_13712,N_13084,N_12352);
nand U13713 (N_13713,N_12689,N_12364);
nand U13714 (N_13714,N_13463,N_12271);
nand U13715 (N_13715,N_12678,N_13038);
nand U13716 (N_13716,N_13327,N_12531);
and U13717 (N_13717,N_13377,N_12530);
nor U13718 (N_13718,N_12996,N_13407);
xnor U13719 (N_13719,N_12025,N_13378);
nand U13720 (N_13720,N_12135,N_12551);
nor U13721 (N_13721,N_12016,N_12210);
nand U13722 (N_13722,N_13371,N_12260);
xnor U13723 (N_13723,N_12901,N_12387);
xor U13724 (N_13724,N_12080,N_12257);
or U13725 (N_13725,N_13120,N_13372);
nand U13726 (N_13726,N_12166,N_12091);
nor U13727 (N_13727,N_13124,N_13341);
nor U13728 (N_13728,N_12926,N_12092);
xor U13729 (N_13729,N_12377,N_12133);
nand U13730 (N_13730,N_12499,N_12616);
nor U13731 (N_13731,N_12704,N_13029);
nor U13732 (N_13732,N_12292,N_12562);
nor U13733 (N_13733,N_13337,N_12857);
nand U13734 (N_13734,N_12082,N_12673);
nand U13735 (N_13735,N_13164,N_13042);
xor U13736 (N_13736,N_13050,N_13461);
or U13737 (N_13737,N_12920,N_12408);
xnor U13738 (N_13738,N_12048,N_12797);
nor U13739 (N_13739,N_12468,N_12434);
nand U13740 (N_13740,N_12520,N_12752);
nand U13741 (N_13741,N_12866,N_12701);
xnor U13742 (N_13742,N_13143,N_12436);
xor U13743 (N_13743,N_12845,N_12739);
xor U13744 (N_13744,N_12469,N_12730);
xor U13745 (N_13745,N_12256,N_12457);
nand U13746 (N_13746,N_12462,N_12475);
or U13747 (N_13747,N_12430,N_12618);
and U13748 (N_13748,N_12812,N_13422);
xnor U13749 (N_13749,N_13305,N_12251);
nand U13750 (N_13750,N_12193,N_12020);
or U13751 (N_13751,N_13174,N_12332);
nor U13752 (N_13752,N_12167,N_12761);
or U13753 (N_13753,N_12001,N_13249);
nor U13754 (N_13754,N_12904,N_13024);
nor U13755 (N_13755,N_13115,N_12201);
or U13756 (N_13756,N_13238,N_13284);
nand U13757 (N_13757,N_12488,N_12267);
nor U13758 (N_13758,N_12355,N_13186);
nor U13759 (N_13759,N_12026,N_13447);
xor U13760 (N_13760,N_12737,N_12902);
or U13761 (N_13761,N_12688,N_13041);
nand U13762 (N_13762,N_13155,N_12425);
nor U13763 (N_13763,N_12793,N_13483);
and U13764 (N_13764,N_12077,N_12813);
or U13765 (N_13765,N_12608,N_13162);
nor U13766 (N_13766,N_13219,N_12733);
or U13767 (N_13767,N_12214,N_12358);
nand U13768 (N_13768,N_12264,N_13215);
xnor U13769 (N_13769,N_13496,N_13119);
or U13770 (N_13770,N_12869,N_13403);
and U13771 (N_13771,N_13139,N_13227);
xor U13772 (N_13772,N_12179,N_12185);
and U13773 (N_13773,N_13442,N_13376);
xor U13774 (N_13774,N_13336,N_13441);
nand U13775 (N_13775,N_13318,N_12129);
and U13776 (N_13776,N_12262,N_12073);
or U13777 (N_13777,N_12921,N_12825);
or U13778 (N_13778,N_12535,N_12395);
nor U13779 (N_13779,N_12980,N_13252);
and U13780 (N_13780,N_12404,N_12261);
or U13781 (N_13781,N_13464,N_12885);
xor U13782 (N_13782,N_13490,N_12736);
nand U13783 (N_13783,N_12041,N_12731);
and U13784 (N_13784,N_12782,N_13025);
xnor U13785 (N_13785,N_12153,N_12331);
nor U13786 (N_13786,N_12175,N_13140);
or U13787 (N_13787,N_13460,N_12072);
or U13788 (N_13788,N_12036,N_13069);
nor U13789 (N_13789,N_12861,N_12478);
nand U13790 (N_13790,N_12014,N_12461);
nor U13791 (N_13791,N_12493,N_12374);
or U13792 (N_13792,N_12748,N_12522);
nand U13793 (N_13793,N_12867,N_12470);
nor U13794 (N_13794,N_12948,N_12013);
and U13795 (N_13795,N_13170,N_13185);
xor U13796 (N_13796,N_13208,N_12959);
and U13797 (N_13797,N_12321,N_12713);
nor U13798 (N_13798,N_12933,N_12066);
and U13799 (N_13799,N_12759,N_12097);
xnor U13800 (N_13800,N_13117,N_13231);
nor U13801 (N_13801,N_12799,N_13197);
nor U13802 (N_13802,N_13302,N_12064);
or U13803 (N_13803,N_13193,N_12536);
and U13804 (N_13804,N_13459,N_12846);
nor U13805 (N_13805,N_12638,N_13251);
and U13806 (N_13806,N_13365,N_12669);
nor U13807 (N_13807,N_12464,N_13128);
nand U13808 (N_13808,N_12572,N_13000);
nand U13809 (N_13809,N_12597,N_12848);
nor U13810 (N_13810,N_13182,N_12668);
xor U13811 (N_13811,N_12301,N_12627);
and U13812 (N_13812,N_12643,N_13027);
and U13813 (N_13813,N_12357,N_12074);
nor U13814 (N_13814,N_12421,N_13269);
and U13815 (N_13815,N_13415,N_13218);
or U13816 (N_13816,N_13187,N_12200);
xnor U13817 (N_13817,N_13456,N_12584);
nor U13818 (N_13818,N_12446,N_12227);
xor U13819 (N_13819,N_12235,N_12419);
nand U13820 (N_13820,N_13329,N_12037);
nand U13821 (N_13821,N_12525,N_13351);
and U13822 (N_13822,N_12662,N_12293);
or U13823 (N_13823,N_12986,N_12031);
xor U13824 (N_13824,N_13061,N_12363);
and U13825 (N_13825,N_12131,N_13194);
or U13826 (N_13826,N_12527,N_12362);
or U13827 (N_13827,N_13354,N_13056);
nor U13828 (N_13828,N_13362,N_12946);
or U13829 (N_13829,N_13036,N_12862);
or U13830 (N_13830,N_12624,N_12107);
nor U13831 (N_13831,N_12830,N_13458);
xor U13832 (N_13832,N_13404,N_12438);
nand U13833 (N_13833,N_13492,N_12786);
xor U13834 (N_13834,N_13413,N_13047);
nand U13835 (N_13835,N_12473,N_13467);
xnor U13836 (N_13836,N_12809,N_12514);
nand U13837 (N_13837,N_13011,N_12947);
nor U13838 (N_13838,N_12549,N_12777);
nand U13839 (N_13839,N_13381,N_13205);
and U13840 (N_13840,N_13109,N_12448);
or U13841 (N_13841,N_12151,N_13275);
or U13842 (N_13842,N_12047,N_12903);
nand U13843 (N_13843,N_12069,N_12750);
nor U13844 (N_13844,N_12335,N_13449);
xor U13845 (N_13845,N_12296,N_12385);
xor U13846 (N_13846,N_13346,N_12022);
and U13847 (N_13847,N_13263,N_13224);
xor U13848 (N_13848,N_13419,N_13465);
xor U13849 (N_13849,N_12231,N_13411);
or U13850 (N_13850,N_12059,N_13126);
xnor U13851 (N_13851,N_13247,N_13129);
and U13852 (N_13852,N_12220,N_12480);
nand U13853 (N_13853,N_12573,N_12791);
and U13854 (N_13854,N_13323,N_13316);
or U13855 (N_13855,N_12173,N_12483);
and U13856 (N_13856,N_12068,N_12213);
and U13857 (N_13857,N_12471,N_13266);
xnor U13858 (N_13858,N_12141,N_13052);
and U13859 (N_13859,N_12629,N_12905);
nor U13860 (N_13860,N_12249,N_12328);
nand U13861 (N_13861,N_13160,N_13488);
xnor U13862 (N_13862,N_12417,N_12429);
nand U13863 (N_13863,N_13018,N_12755);
xor U13864 (N_13864,N_12843,N_13246);
nand U13865 (N_13865,N_12263,N_13297);
and U13866 (N_13866,N_12623,N_12098);
and U13867 (N_13867,N_12934,N_13473);
or U13868 (N_13868,N_12343,N_12106);
and U13869 (N_13869,N_12694,N_12824);
or U13870 (N_13870,N_12892,N_12952);
or U13871 (N_13871,N_12798,N_13169);
and U13872 (N_13872,N_13087,N_12878);
and U13873 (N_13873,N_12087,N_13309);
nand U13874 (N_13874,N_12006,N_12864);
or U13875 (N_13875,N_12838,N_12894);
xor U13876 (N_13876,N_12968,N_13342);
nand U13877 (N_13877,N_12868,N_12609);
and U13878 (N_13878,N_12412,N_13045);
xor U13879 (N_13879,N_12286,N_12351);
xnor U13880 (N_13880,N_12496,N_12617);
nor U13881 (N_13881,N_12751,N_12962);
nor U13882 (N_13882,N_12524,N_12226);
xnor U13883 (N_13883,N_13145,N_12992);
xnor U13884 (N_13884,N_12939,N_12088);
and U13885 (N_13885,N_12413,N_12863);
xor U13886 (N_13886,N_12721,N_12817);
nor U13887 (N_13887,N_12816,N_12712);
nand U13888 (N_13888,N_13388,N_13138);
and U13889 (N_13889,N_12376,N_12081);
and U13890 (N_13890,N_12030,N_12181);
or U13891 (N_13891,N_12971,N_13481);
or U13892 (N_13892,N_13244,N_13300);
or U13893 (N_13893,N_12467,N_12298);
xnor U13894 (N_13894,N_12183,N_12275);
and U13895 (N_13895,N_12528,N_12028);
and U13896 (N_13896,N_12309,N_13307);
xor U13897 (N_13897,N_12686,N_12334);
nor U13898 (N_13898,N_12646,N_12943);
nor U13899 (N_13899,N_12592,N_12466);
or U13900 (N_13900,N_12749,N_12729);
xor U13901 (N_13901,N_12693,N_13439);
nor U13902 (N_13902,N_13395,N_12272);
nor U13903 (N_13903,N_12396,N_12519);
nand U13904 (N_13904,N_12416,N_12397);
and U13905 (N_13905,N_12159,N_13171);
or U13906 (N_13906,N_13110,N_12070);
and U13907 (N_13907,N_12936,N_12116);
nor U13908 (N_13908,N_12930,N_12954);
nand U13909 (N_13909,N_12763,N_12239);
nand U13910 (N_13910,N_12229,N_13142);
or U13911 (N_13911,N_12341,N_13279);
xor U13912 (N_13912,N_13007,N_12611);
xnor U13913 (N_13913,N_12567,N_12442);
nand U13914 (N_13914,N_12929,N_13037);
and U13915 (N_13915,N_12038,N_13452);
nand U13916 (N_13916,N_12979,N_12320);
nand U13917 (N_13917,N_13014,N_12168);
and U13918 (N_13918,N_12906,N_12391);
and U13919 (N_13919,N_12989,N_12795);
xor U13920 (N_13920,N_12122,N_12095);
nor U13921 (N_13921,N_13276,N_13282);
nand U13922 (N_13922,N_13418,N_12369);
nor U13923 (N_13923,N_13063,N_13394);
xnor U13924 (N_13924,N_13257,N_13060);
or U13925 (N_13925,N_12170,N_12526);
nand U13926 (N_13926,N_13368,N_13204);
nand U13927 (N_13927,N_13438,N_12808);
nand U13928 (N_13928,N_12615,N_12695);
and U13929 (N_13929,N_13331,N_13131);
or U13930 (N_13930,N_12509,N_13235);
and U13931 (N_13931,N_12784,N_12963);
or U13932 (N_13932,N_13270,N_12648);
or U13933 (N_13933,N_12870,N_12973);
nand U13934 (N_13934,N_13340,N_12647);
nor U13935 (N_13935,N_12696,N_12024);
xnor U13936 (N_13936,N_12735,N_12085);
nor U13937 (N_13937,N_12718,N_13073);
nand U13938 (N_13938,N_12240,N_12970);
and U13939 (N_13939,N_12223,N_12876);
or U13940 (N_13940,N_12350,N_12801);
xor U13941 (N_13941,N_12117,N_13491);
nand U13942 (N_13942,N_12518,N_12898);
xnor U13943 (N_13943,N_12783,N_12241);
and U13944 (N_13944,N_12625,N_12667);
xor U13945 (N_13945,N_13301,N_13040);
or U13946 (N_13946,N_12633,N_12062);
nor U13947 (N_13947,N_12781,N_13364);
or U13948 (N_13948,N_12506,N_12110);
xnor U13949 (N_13949,N_13363,N_12766);
nand U13950 (N_13950,N_12742,N_12724);
or U13951 (N_13951,N_13250,N_12977);
or U13952 (N_13952,N_12437,N_12382);
nand U13953 (N_13953,N_12283,N_13241);
xor U13954 (N_13954,N_13405,N_12957);
nand U13955 (N_13955,N_12449,N_13296);
nand U13956 (N_13956,N_12741,N_12427);
xnor U13957 (N_13957,N_13277,N_12454);
and U13958 (N_13958,N_13325,N_12268);
or U13959 (N_13959,N_13188,N_12378);
nor U13960 (N_13960,N_12057,N_12854);
and U13961 (N_13961,N_12928,N_12663);
or U13962 (N_13962,N_12177,N_12657);
or U13963 (N_13963,N_13179,N_13290);
and U13964 (N_13964,N_12822,N_12491);
and U13965 (N_13965,N_12844,N_13310);
xor U13966 (N_13966,N_12017,N_12553);
nor U13967 (N_13967,N_12743,N_12053);
and U13968 (N_13968,N_12517,N_12820);
nand U13969 (N_13969,N_12965,N_12762);
nor U13970 (N_13970,N_12004,N_13373);
nand U13971 (N_13971,N_12953,N_12561);
xnor U13972 (N_13972,N_12708,N_12197);
xor U13973 (N_13973,N_12547,N_12302);
or U13974 (N_13974,N_12697,N_12778);
or U13975 (N_13975,N_13470,N_12826);
nor U13976 (N_13976,N_12940,N_13102);
nor U13977 (N_13977,N_13134,N_12063);
nand U13978 (N_13978,N_12566,N_13414);
or U13979 (N_13979,N_12148,N_13043);
nand U13980 (N_13980,N_13347,N_12212);
nor U13981 (N_13981,N_12216,N_12612);
and U13982 (N_13982,N_12246,N_12218);
and U13983 (N_13983,N_12852,N_13021);
nand U13984 (N_13984,N_12683,N_12503);
and U13985 (N_13985,N_13136,N_13105);
nand U13986 (N_13986,N_12120,N_13089);
and U13987 (N_13987,N_12998,N_12847);
nor U13988 (N_13988,N_13444,N_12347);
nand U13989 (N_13989,N_13133,N_12723);
nor U13990 (N_13990,N_12486,N_13149);
nand U13991 (N_13991,N_12086,N_13245);
xor U13992 (N_13992,N_12666,N_12671);
and U13993 (N_13993,N_13497,N_12874);
and U13994 (N_13994,N_12537,N_12716);
xor U13995 (N_13995,N_13440,N_12171);
nor U13996 (N_13996,N_12775,N_12534);
nor U13997 (N_13997,N_13137,N_12888);
or U13998 (N_13998,N_12198,N_13477);
nand U13999 (N_13999,N_12252,N_12559);
and U14000 (N_14000,N_12265,N_13001);
xor U14001 (N_14001,N_12859,N_12814);
and U14002 (N_14002,N_12340,N_12583);
xor U14003 (N_14003,N_13357,N_12418);
and U14004 (N_14004,N_12184,N_13443);
nor U14005 (N_14005,N_13367,N_13401);
nand U14006 (N_14006,N_13141,N_12916);
nand U14007 (N_14007,N_12978,N_13450);
and U14008 (N_14008,N_12744,N_13049);
xor U14009 (N_14009,N_13398,N_13387);
nand U14010 (N_14010,N_13446,N_13468);
and U14011 (N_14011,N_12021,N_12911);
and U14012 (N_14012,N_12672,N_13004);
or U14013 (N_14013,N_12760,N_13010);
xor U14014 (N_14014,N_13299,N_12189);
and U14015 (N_14015,N_12912,N_12675);
nand U14016 (N_14016,N_13260,N_12443);
nor U14017 (N_14017,N_13312,N_12720);
or U14018 (N_14018,N_12545,N_12359);
nor U14019 (N_14019,N_12539,N_12807);
or U14020 (N_14020,N_12881,N_13172);
or U14021 (N_14021,N_13076,N_12336);
nor U14022 (N_14022,N_13292,N_13424);
nand U14023 (N_14023,N_13151,N_13108);
and U14024 (N_14024,N_13314,N_13079);
and U14025 (N_14025,N_12108,N_12884);
and U14026 (N_14026,N_13278,N_12909);
or U14027 (N_14027,N_12324,N_13034);
or U14028 (N_14028,N_13015,N_13130);
nand U14029 (N_14029,N_12029,N_12388);
and U14030 (N_14030,N_12569,N_13248);
nor U14031 (N_14031,N_12015,N_12191);
nor U14032 (N_14032,N_13360,N_12234);
or U14033 (N_14033,N_12444,N_13031);
or U14034 (N_14034,N_12574,N_13003);
nor U14035 (N_14035,N_13005,N_12203);
or U14036 (N_14036,N_12719,N_12605);
xor U14037 (N_14037,N_12312,N_13285);
nand U14038 (N_14038,N_13281,N_12375);
or U14039 (N_14039,N_12532,N_13271);
and U14040 (N_14040,N_12521,N_12407);
nand U14041 (N_14041,N_13402,N_12139);
and U14042 (N_14042,N_12690,N_12076);
xnor U14043 (N_14043,N_12851,N_12543);
nand U14044 (N_14044,N_12450,N_12684);
nor U14045 (N_14045,N_12114,N_12855);
or U14046 (N_14046,N_12803,N_13268);
nand U14047 (N_14047,N_13163,N_13295);
nand U14048 (N_14048,N_12371,N_13304);
nor U14049 (N_14049,N_13071,N_13333);
xor U14050 (N_14050,N_12327,N_12492);
or U14051 (N_14051,N_13427,N_13306);
xor U14052 (N_14052,N_13343,N_13200);
nor U14053 (N_14053,N_12279,N_12621);
nor U14054 (N_14054,N_13486,N_13454);
and U14055 (N_14055,N_13068,N_12232);
or U14056 (N_14056,N_13289,N_12472);
or U14057 (N_14057,N_12394,N_12215);
or U14058 (N_14058,N_12313,N_12225);
xor U14059 (N_14059,N_13344,N_12563);
nor U14060 (N_14060,N_13154,N_12315);
nor U14061 (N_14061,N_12119,N_13382);
nand U14062 (N_14062,N_12792,N_12329);
or U14063 (N_14063,N_12972,N_12839);
nor U14064 (N_14064,N_13420,N_13062);
xnor U14065 (N_14065,N_12144,N_12634);
and U14066 (N_14066,N_12207,N_12452);
or U14067 (N_14067,N_13258,N_12589);
or U14068 (N_14068,N_12401,N_12727);
and U14069 (N_14069,N_13298,N_13355);
and U14070 (N_14070,N_13335,N_13400);
nand U14071 (N_14071,N_12349,N_13096);
xor U14072 (N_14072,N_12003,N_13075);
nand U14073 (N_14073,N_13116,N_13054);
and U14074 (N_14074,N_12588,N_12722);
and U14075 (N_14075,N_13203,N_12367);
nor U14076 (N_14076,N_12384,N_12516);
or U14077 (N_14077,N_12278,N_12596);
nand U14078 (N_14078,N_12922,N_12089);
nor U14079 (N_14079,N_12011,N_12428);
or U14080 (N_14080,N_12630,N_12802);
nor U14081 (N_14081,N_12754,N_13409);
and U14082 (N_14082,N_12154,N_12163);
nand U14083 (N_14083,N_13273,N_12319);
nor U14084 (N_14084,N_12747,N_13232);
or U14085 (N_14085,N_12714,N_12126);
nand U14086 (N_14086,N_12570,N_12805);
nand U14087 (N_14087,N_13480,N_13006);
nor U14088 (N_14088,N_13180,N_12344);
nand U14089 (N_14089,N_13202,N_12034);
or U14090 (N_14090,N_12445,N_13392);
nand U14091 (N_14091,N_12342,N_12460);
or U14092 (N_14092,N_12075,N_13326);
xor U14093 (N_14093,N_12976,N_12935);
xor U14094 (N_14094,N_12927,N_12705);
xnor U14095 (N_14095,N_12190,N_13397);
xnor U14096 (N_14096,N_13099,N_13383);
nor U14097 (N_14097,N_13207,N_13435);
nor U14098 (N_14098,N_12918,N_12756);
nand U14099 (N_14099,N_12635,N_13125);
and U14100 (N_14100,N_12311,N_12033);
xnor U14101 (N_14101,N_12316,N_12571);
and U14102 (N_14102,N_12308,N_12259);
xor U14103 (N_14103,N_13057,N_12433);
nand U14104 (N_14104,N_12832,N_13181);
nor U14105 (N_14105,N_12247,N_12113);
or U14106 (N_14106,N_12932,N_12925);
nand U14107 (N_14107,N_12770,N_12990);
xnor U14108 (N_14108,N_12330,N_12604);
or U14109 (N_14109,N_12511,N_12050);
nor U14110 (N_14110,N_13112,N_12127);
nand U14111 (N_14111,N_12000,N_12512);
xnor U14112 (N_14112,N_12555,N_12550);
or U14113 (N_14113,N_13315,N_13230);
nand U14114 (N_14114,N_12745,N_12236);
xnor U14115 (N_14115,N_12546,N_12322);
or U14116 (N_14116,N_12039,N_12849);
nand U14117 (N_14117,N_12831,N_12649);
and U14118 (N_14118,N_13028,N_12269);
and U14119 (N_14119,N_12365,N_13254);
and U14120 (N_14120,N_12061,N_12474);
and U14121 (N_14121,N_12515,N_13013);
xnor U14122 (N_14122,N_13274,N_12023);
nor U14123 (N_14123,N_13455,N_12659);
and U14124 (N_14124,N_12982,N_13462);
nor U14125 (N_14125,N_12700,N_12224);
nand U14126 (N_14126,N_12270,N_12548);
nor U14127 (N_14127,N_12595,N_12490);
nor U14128 (N_14128,N_12987,N_12726);
and U14129 (N_14129,N_13349,N_12160);
xor U14130 (N_14130,N_12393,N_12233);
or U14131 (N_14131,N_12294,N_13471);
or U14132 (N_14132,N_13399,N_12042);
nand U14133 (N_14133,N_12479,N_12999);
xor U14134 (N_14134,N_13225,N_12890);
or U14135 (N_14135,N_12658,N_13393);
and U14136 (N_14136,N_13234,N_13359);
nand U14137 (N_14137,N_13147,N_12192);
xor U14138 (N_14138,N_13085,N_13406);
nor U14139 (N_14139,N_12580,N_12482);
nor U14140 (N_14140,N_13080,N_13106);
and U14141 (N_14141,N_12500,N_12641);
and U14142 (N_14142,N_12655,N_12711);
nor U14143 (N_14143,N_12498,N_12915);
xor U14144 (N_14144,N_12827,N_12554);
xnor U14145 (N_14145,N_12771,N_12182);
or U14146 (N_14146,N_12386,N_12899);
nor U14147 (N_14147,N_12703,N_12631);
or U14148 (N_14148,N_13428,N_12305);
nand U14149 (N_14149,N_12821,N_12908);
or U14150 (N_14150,N_12137,N_12284);
xor U14151 (N_14151,N_13097,N_12676);
xnor U14152 (N_14152,N_12942,N_12027);
or U14153 (N_14153,N_13317,N_12556);
or U14154 (N_14154,N_12660,N_12651);
or U14155 (N_14155,N_12656,N_13098);
nor U14156 (N_14156,N_12585,N_13320);
and U14157 (N_14157,N_13358,N_12424);
xor U14158 (N_14158,N_12431,N_12818);
or U14159 (N_14159,N_12194,N_13345);
xnor U14160 (N_14160,N_13051,N_12765);
nor U14161 (N_14161,N_12560,N_12339);
nand U14162 (N_14162,N_12924,N_13243);
xor U14163 (N_14163,N_13469,N_12018);
xor U14164 (N_14164,N_12917,N_13380);
nor U14165 (N_14165,N_13146,N_12306);
and U14166 (N_14166,N_13391,N_12579);
nor U14167 (N_14167,N_12523,N_13122);
nand U14168 (N_14168,N_12372,N_12958);
or U14169 (N_14169,N_13161,N_12966);
xnor U14170 (N_14170,N_12640,N_12243);
nand U14171 (N_14171,N_12323,N_12691);
and U14172 (N_14172,N_13039,N_13091);
nor U14173 (N_14173,N_13088,N_12273);
nor U14174 (N_14174,N_13253,N_12055);
and U14175 (N_14175,N_12692,N_12594);
nor U14176 (N_14176,N_12282,N_13066);
xor U14177 (N_14177,N_12040,N_12115);
or U14178 (N_14178,N_12578,N_12758);
nand U14179 (N_14179,N_12833,N_13191);
xor U14180 (N_14180,N_13132,N_13217);
or U14181 (N_14181,N_12045,N_12599);
xnor U14182 (N_14182,N_13353,N_13111);
or U14183 (N_14183,N_13148,N_13286);
and U14184 (N_14184,N_12439,N_13081);
or U14185 (N_14185,N_13437,N_12368);
nand U14186 (N_14186,N_13107,N_13324);
nor U14187 (N_14187,N_13303,N_12794);
xor U14188 (N_14188,N_12769,N_12757);
nand U14189 (N_14189,N_12834,N_13059);
nand U14190 (N_14190,N_12373,N_13417);
xnor U14191 (N_14191,N_12422,N_12853);
and U14192 (N_14192,N_12841,N_12158);
or U14193 (N_14193,N_13384,N_13046);
and U14194 (N_14194,N_12914,N_13094);
or U14195 (N_14195,N_12804,N_12090);
nand U14196 (N_14196,N_12304,N_12100);
nor U14197 (N_14197,N_12974,N_12887);
nand U14198 (N_14198,N_12338,N_12432);
and U14199 (N_14199,N_12005,N_13445);
or U14200 (N_14200,N_12299,N_13190);
xor U14201 (N_14201,N_13221,N_13206);
and U14202 (N_14202,N_12118,N_13065);
or U14203 (N_14203,N_13168,N_12710);
or U14204 (N_14204,N_12157,N_13167);
or U14205 (N_14205,N_12709,N_13095);
or U14206 (N_14206,N_12465,N_12451);
or U14207 (N_14207,N_13369,N_13375);
nor U14208 (N_14208,N_12565,N_12650);
and U14209 (N_14209,N_13196,N_12622);
and U14210 (N_14210,N_13067,N_12156);
nor U14211 (N_14211,N_13265,N_12481);
nand U14212 (N_14212,N_13158,N_12314);
xor U14213 (N_14213,N_13334,N_12248);
nand U14214 (N_14214,N_13210,N_13086);
nand U14215 (N_14215,N_12199,N_13494);
and U14216 (N_14216,N_12895,N_12204);
nand U14217 (N_14217,N_12035,N_13412);
nor U14218 (N_14218,N_12165,N_12564);
or U14219 (N_14219,N_12789,N_13356);
nand U14220 (N_14220,N_13114,N_12244);
nand U14221 (N_14221,N_12740,N_13436);
and U14222 (N_14222,N_12392,N_12715);
nand U14223 (N_14223,N_12502,N_12162);
and U14224 (N_14224,N_12591,N_12568);
nand U14225 (N_14225,N_12937,N_12138);
and U14226 (N_14226,N_12219,N_12161);
xor U14227 (N_14227,N_12505,N_12586);
nor U14228 (N_14228,N_12440,N_13150);
and U14229 (N_14229,N_13121,N_12602);
xor U14230 (N_14230,N_12950,N_12354);
nand U14231 (N_14231,N_13127,N_13228);
and U14232 (N_14232,N_12644,N_13390);
nor U14233 (N_14233,N_12738,N_12172);
xnor U14234 (N_14234,N_12835,N_13495);
and U14235 (N_14235,N_12140,N_12130);
nor U14236 (N_14236,N_12628,N_12326);
nor U14237 (N_14237,N_13009,N_12707);
xnor U14238 (N_14238,N_12078,N_12875);
nor U14239 (N_14239,N_13199,N_12441);
or U14240 (N_14240,N_13242,N_13410);
or U14241 (N_14241,N_13055,N_12307);
xnor U14242 (N_14242,N_12188,N_12645);
xor U14243 (N_14243,N_12136,N_12593);
or U14244 (N_14244,N_13287,N_12558);
nor U14245 (N_14245,N_12815,N_13313);
nor U14246 (N_14246,N_12872,N_12582);
nor U14247 (N_14247,N_12463,N_12217);
and U14248 (N_14248,N_12058,N_12706);
nor U14249 (N_14249,N_12164,N_12636);
and U14250 (N_14250,N_13481,N_12706);
or U14251 (N_14251,N_12389,N_12429);
nand U14252 (N_14252,N_13147,N_12819);
and U14253 (N_14253,N_12053,N_13305);
nand U14254 (N_14254,N_12366,N_12801);
nor U14255 (N_14255,N_12576,N_12142);
or U14256 (N_14256,N_12885,N_13117);
xnor U14257 (N_14257,N_13470,N_12996);
xnor U14258 (N_14258,N_13449,N_13116);
nand U14259 (N_14259,N_12022,N_12089);
xor U14260 (N_14260,N_13377,N_12685);
and U14261 (N_14261,N_13333,N_13381);
nor U14262 (N_14262,N_12329,N_13259);
or U14263 (N_14263,N_13245,N_13314);
xor U14264 (N_14264,N_12264,N_12066);
nand U14265 (N_14265,N_13325,N_12095);
xnor U14266 (N_14266,N_13273,N_12414);
nor U14267 (N_14267,N_12796,N_12747);
or U14268 (N_14268,N_12328,N_13166);
nor U14269 (N_14269,N_12666,N_12644);
xor U14270 (N_14270,N_12565,N_13337);
nand U14271 (N_14271,N_13293,N_12567);
and U14272 (N_14272,N_12124,N_13354);
xor U14273 (N_14273,N_12391,N_13370);
nor U14274 (N_14274,N_12022,N_12730);
xor U14275 (N_14275,N_12501,N_13157);
nand U14276 (N_14276,N_12397,N_12596);
and U14277 (N_14277,N_12249,N_12811);
and U14278 (N_14278,N_12176,N_13104);
nand U14279 (N_14279,N_12045,N_12612);
and U14280 (N_14280,N_12937,N_12223);
xnor U14281 (N_14281,N_13348,N_12764);
nor U14282 (N_14282,N_13361,N_12367);
or U14283 (N_14283,N_13489,N_12028);
xnor U14284 (N_14284,N_12084,N_12537);
or U14285 (N_14285,N_13304,N_13051);
or U14286 (N_14286,N_13442,N_12994);
or U14287 (N_14287,N_12042,N_13147);
nor U14288 (N_14288,N_12816,N_12723);
or U14289 (N_14289,N_12170,N_13397);
and U14290 (N_14290,N_12626,N_12126);
xnor U14291 (N_14291,N_12132,N_13175);
xor U14292 (N_14292,N_13484,N_12685);
and U14293 (N_14293,N_12418,N_13280);
or U14294 (N_14294,N_12493,N_12440);
xnor U14295 (N_14295,N_12849,N_13226);
or U14296 (N_14296,N_12169,N_12122);
nor U14297 (N_14297,N_13349,N_13290);
nor U14298 (N_14298,N_12257,N_13149);
xor U14299 (N_14299,N_12621,N_12549);
and U14300 (N_14300,N_12536,N_12362);
xor U14301 (N_14301,N_12511,N_13164);
nand U14302 (N_14302,N_12844,N_13069);
nand U14303 (N_14303,N_12046,N_12603);
nor U14304 (N_14304,N_12610,N_12239);
xor U14305 (N_14305,N_13302,N_13100);
and U14306 (N_14306,N_12730,N_12969);
or U14307 (N_14307,N_12639,N_12171);
or U14308 (N_14308,N_13416,N_12978);
and U14309 (N_14309,N_12008,N_12293);
and U14310 (N_14310,N_12679,N_12465);
xor U14311 (N_14311,N_12237,N_12397);
and U14312 (N_14312,N_13089,N_13043);
xnor U14313 (N_14313,N_13164,N_12780);
xnor U14314 (N_14314,N_12247,N_12655);
nor U14315 (N_14315,N_13216,N_13233);
nor U14316 (N_14316,N_12815,N_13266);
and U14317 (N_14317,N_12729,N_12332);
xnor U14318 (N_14318,N_12988,N_13494);
nor U14319 (N_14319,N_13236,N_13211);
nor U14320 (N_14320,N_12847,N_13223);
nand U14321 (N_14321,N_13228,N_12482);
nor U14322 (N_14322,N_13092,N_13477);
or U14323 (N_14323,N_13240,N_13250);
nor U14324 (N_14324,N_12200,N_12814);
xor U14325 (N_14325,N_12700,N_12583);
nor U14326 (N_14326,N_13197,N_12074);
nand U14327 (N_14327,N_12228,N_12879);
nand U14328 (N_14328,N_13043,N_12842);
and U14329 (N_14329,N_13002,N_13266);
nand U14330 (N_14330,N_12046,N_13221);
nand U14331 (N_14331,N_12684,N_12800);
and U14332 (N_14332,N_12426,N_12141);
nor U14333 (N_14333,N_12072,N_12726);
and U14334 (N_14334,N_12640,N_13483);
and U14335 (N_14335,N_13208,N_13282);
or U14336 (N_14336,N_12864,N_13242);
nor U14337 (N_14337,N_12017,N_13013);
and U14338 (N_14338,N_12679,N_13282);
or U14339 (N_14339,N_13022,N_12939);
or U14340 (N_14340,N_12614,N_12792);
xnor U14341 (N_14341,N_12915,N_13028);
nand U14342 (N_14342,N_12678,N_13349);
nor U14343 (N_14343,N_13267,N_12903);
nand U14344 (N_14344,N_12070,N_12859);
or U14345 (N_14345,N_13105,N_12885);
and U14346 (N_14346,N_13335,N_12615);
and U14347 (N_14347,N_13164,N_12076);
xor U14348 (N_14348,N_13003,N_13485);
or U14349 (N_14349,N_13374,N_13260);
nor U14350 (N_14350,N_12556,N_12624);
nor U14351 (N_14351,N_12865,N_12102);
and U14352 (N_14352,N_12020,N_12884);
and U14353 (N_14353,N_12837,N_12496);
xor U14354 (N_14354,N_13201,N_12914);
nor U14355 (N_14355,N_13059,N_13187);
nand U14356 (N_14356,N_12269,N_12723);
nor U14357 (N_14357,N_12618,N_12035);
xor U14358 (N_14358,N_12303,N_13166);
nor U14359 (N_14359,N_13128,N_13126);
nor U14360 (N_14360,N_12436,N_12739);
or U14361 (N_14361,N_12559,N_12139);
xnor U14362 (N_14362,N_13161,N_13382);
xor U14363 (N_14363,N_12817,N_12621);
nor U14364 (N_14364,N_12258,N_13322);
nor U14365 (N_14365,N_13208,N_12570);
and U14366 (N_14366,N_13437,N_12450);
nand U14367 (N_14367,N_13268,N_13437);
or U14368 (N_14368,N_12426,N_13133);
nand U14369 (N_14369,N_13348,N_12078);
nor U14370 (N_14370,N_12685,N_13139);
and U14371 (N_14371,N_12974,N_12324);
or U14372 (N_14372,N_12534,N_12908);
xor U14373 (N_14373,N_12714,N_13347);
xnor U14374 (N_14374,N_13038,N_12471);
nor U14375 (N_14375,N_13230,N_12726);
xor U14376 (N_14376,N_12023,N_12150);
xnor U14377 (N_14377,N_12892,N_12389);
or U14378 (N_14378,N_12214,N_13026);
xnor U14379 (N_14379,N_12772,N_12309);
and U14380 (N_14380,N_13242,N_12469);
nand U14381 (N_14381,N_12851,N_13049);
xor U14382 (N_14382,N_13276,N_13154);
or U14383 (N_14383,N_13038,N_12133);
xor U14384 (N_14384,N_12484,N_12775);
and U14385 (N_14385,N_12047,N_12659);
and U14386 (N_14386,N_12352,N_12136);
nand U14387 (N_14387,N_12633,N_12136);
and U14388 (N_14388,N_12313,N_13031);
nor U14389 (N_14389,N_13032,N_13192);
nand U14390 (N_14390,N_12494,N_12748);
nand U14391 (N_14391,N_13358,N_12301);
nor U14392 (N_14392,N_13169,N_13404);
nand U14393 (N_14393,N_12732,N_12895);
nand U14394 (N_14394,N_12569,N_12693);
nand U14395 (N_14395,N_12291,N_12263);
nand U14396 (N_14396,N_12598,N_12984);
nor U14397 (N_14397,N_12939,N_13343);
nand U14398 (N_14398,N_12927,N_13389);
xnor U14399 (N_14399,N_13425,N_12177);
or U14400 (N_14400,N_13145,N_12471);
nand U14401 (N_14401,N_12480,N_12846);
nand U14402 (N_14402,N_12009,N_13188);
nor U14403 (N_14403,N_13064,N_12394);
nand U14404 (N_14404,N_12763,N_12704);
nand U14405 (N_14405,N_13157,N_13203);
and U14406 (N_14406,N_12438,N_12096);
and U14407 (N_14407,N_12591,N_13221);
or U14408 (N_14408,N_12548,N_12772);
xor U14409 (N_14409,N_12064,N_13068);
or U14410 (N_14410,N_12745,N_13281);
nor U14411 (N_14411,N_13036,N_13039);
nand U14412 (N_14412,N_12322,N_12654);
or U14413 (N_14413,N_13057,N_13365);
xor U14414 (N_14414,N_12434,N_12746);
or U14415 (N_14415,N_12339,N_12314);
or U14416 (N_14416,N_12095,N_12245);
nor U14417 (N_14417,N_12835,N_12103);
nor U14418 (N_14418,N_13435,N_12275);
and U14419 (N_14419,N_13240,N_12141);
xnor U14420 (N_14420,N_12423,N_13379);
and U14421 (N_14421,N_12934,N_13067);
and U14422 (N_14422,N_13343,N_12968);
or U14423 (N_14423,N_13078,N_13127);
or U14424 (N_14424,N_12987,N_12468);
nor U14425 (N_14425,N_12687,N_13468);
xnor U14426 (N_14426,N_12875,N_12066);
nor U14427 (N_14427,N_13104,N_12343);
or U14428 (N_14428,N_13370,N_12049);
xor U14429 (N_14429,N_13313,N_12633);
nor U14430 (N_14430,N_13415,N_12977);
nor U14431 (N_14431,N_13273,N_12796);
or U14432 (N_14432,N_13158,N_12173);
nor U14433 (N_14433,N_13470,N_13153);
nand U14434 (N_14434,N_12583,N_13355);
xnor U14435 (N_14435,N_12861,N_12505);
and U14436 (N_14436,N_12437,N_12669);
or U14437 (N_14437,N_12923,N_13319);
nand U14438 (N_14438,N_12569,N_12828);
or U14439 (N_14439,N_12809,N_13442);
xor U14440 (N_14440,N_13496,N_13105);
xor U14441 (N_14441,N_12309,N_13443);
nor U14442 (N_14442,N_12894,N_13154);
nor U14443 (N_14443,N_12345,N_12082);
xor U14444 (N_14444,N_12071,N_13221);
and U14445 (N_14445,N_13076,N_12982);
xnor U14446 (N_14446,N_13451,N_13430);
nor U14447 (N_14447,N_13008,N_12102);
nand U14448 (N_14448,N_12227,N_13199);
nand U14449 (N_14449,N_13308,N_12127);
and U14450 (N_14450,N_13337,N_12413);
or U14451 (N_14451,N_12698,N_12148);
xnor U14452 (N_14452,N_13269,N_12091);
nand U14453 (N_14453,N_12054,N_12557);
or U14454 (N_14454,N_12064,N_12151);
and U14455 (N_14455,N_12813,N_12183);
nand U14456 (N_14456,N_13148,N_13199);
nor U14457 (N_14457,N_13133,N_12851);
nand U14458 (N_14458,N_13150,N_13465);
nor U14459 (N_14459,N_12575,N_13116);
xor U14460 (N_14460,N_12699,N_12984);
or U14461 (N_14461,N_13371,N_13413);
or U14462 (N_14462,N_13405,N_13398);
or U14463 (N_14463,N_12169,N_12969);
nor U14464 (N_14464,N_13128,N_12465);
or U14465 (N_14465,N_13169,N_12737);
nand U14466 (N_14466,N_12136,N_12411);
nand U14467 (N_14467,N_12207,N_12653);
xnor U14468 (N_14468,N_12293,N_12168);
nor U14469 (N_14469,N_13015,N_13280);
or U14470 (N_14470,N_13029,N_12759);
nor U14471 (N_14471,N_13100,N_13127);
nor U14472 (N_14472,N_12799,N_13377);
xnor U14473 (N_14473,N_12992,N_12307);
or U14474 (N_14474,N_12091,N_13460);
nand U14475 (N_14475,N_13389,N_12529);
and U14476 (N_14476,N_12619,N_13358);
xor U14477 (N_14477,N_12699,N_13016);
nand U14478 (N_14478,N_12803,N_13183);
nand U14479 (N_14479,N_12080,N_12709);
xor U14480 (N_14480,N_13441,N_12473);
nand U14481 (N_14481,N_13270,N_13391);
xor U14482 (N_14482,N_12569,N_12472);
nand U14483 (N_14483,N_12262,N_13196);
nand U14484 (N_14484,N_12152,N_13022);
and U14485 (N_14485,N_13125,N_13362);
nor U14486 (N_14486,N_12757,N_13494);
xnor U14487 (N_14487,N_13363,N_12359);
or U14488 (N_14488,N_12510,N_13152);
and U14489 (N_14489,N_12794,N_12219);
xnor U14490 (N_14490,N_12261,N_13028);
nand U14491 (N_14491,N_12086,N_12141);
nand U14492 (N_14492,N_12568,N_12328);
nor U14493 (N_14493,N_12295,N_13287);
xnor U14494 (N_14494,N_12036,N_12607);
xnor U14495 (N_14495,N_12238,N_13313);
or U14496 (N_14496,N_12511,N_13150);
nor U14497 (N_14497,N_12360,N_12536);
and U14498 (N_14498,N_12886,N_12107);
nor U14499 (N_14499,N_13385,N_12689);
xor U14500 (N_14500,N_12742,N_12660);
and U14501 (N_14501,N_12793,N_13331);
nand U14502 (N_14502,N_12280,N_12715);
or U14503 (N_14503,N_13178,N_12656);
and U14504 (N_14504,N_13356,N_12988);
and U14505 (N_14505,N_12609,N_12071);
xnor U14506 (N_14506,N_12424,N_12698);
and U14507 (N_14507,N_12512,N_13367);
or U14508 (N_14508,N_12677,N_12105);
and U14509 (N_14509,N_12472,N_12691);
and U14510 (N_14510,N_13248,N_12413);
and U14511 (N_14511,N_12727,N_12742);
xor U14512 (N_14512,N_12539,N_12534);
xnor U14513 (N_14513,N_12469,N_12933);
xor U14514 (N_14514,N_12751,N_12040);
and U14515 (N_14515,N_12743,N_12111);
and U14516 (N_14516,N_12012,N_12194);
nor U14517 (N_14517,N_12450,N_12504);
nor U14518 (N_14518,N_13069,N_13056);
and U14519 (N_14519,N_12016,N_13350);
nand U14520 (N_14520,N_12036,N_13440);
nor U14521 (N_14521,N_12261,N_12841);
nor U14522 (N_14522,N_12173,N_13007);
and U14523 (N_14523,N_12000,N_13110);
xnor U14524 (N_14524,N_12167,N_12886);
nand U14525 (N_14525,N_13196,N_12358);
nor U14526 (N_14526,N_12637,N_12572);
nand U14527 (N_14527,N_12609,N_13057);
nand U14528 (N_14528,N_12909,N_13422);
nor U14529 (N_14529,N_13125,N_12306);
or U14530 (N_14530,N_13359,N_13427);
and U14531 (N_14531,N_12802,N_13116);
xnor U14532 (N_14532,N_13335,N_12113);
or U14533 (N_14533,N_12570,N_13116);
nand U14534 (N_14534,N_13396,N_12272);
nor U14535 (N_14535,N_12307,N_13042);
xnor U14536 (N_14536,N_12861,N_12866);
or U14537 (N_14537,N_13464,N_12576);
nand U14538 (N_14538,N_12975,N_12204);
xor U14539 (N_14539,N_12889,N_12692);
and U14540 (N_14540,N_13424,N_12591);
and U14541 (N_14541,N_12101,N_13361);
nor U14542 (N_14542,N_12548,N_12817);
or U14543 (N_14543,N_13175,N_12238);
and U14544 (N_14544,N_12979,N_12183);
nor U14545 (N_14545,N_13498,N_13377);
xor U14546 (N_14546,N_13282,N_13335);
nor U14547 (N_14547,N_13444,N_12872);
nand U14548 (N_14548,N_12599,N_13129);
or U14549 (N_14549,N_12520,N_12899);
nor U14550 (N_14550,N_12161,N_13132);
nand U14551 (N_14551,N_12238,N_12736);
xor U14552 (N_14552,N_12495,N_12618);
nor U14553 (N_14553,N_12597,N_13092);
xnor U14554 (N_14554,N_13306,N_13171);
or U14555 (N_14555,N_13186,N_12765);
nand U14556 (N_14556,N_12466,N_12860);
nand U14557 (N_14557,N_12056,N_12283);
and U14558 (N_14558,N_12487,N_13338);
and U14559 (N_14559,N_12394,N_12971);
nand U14560 (N_14560,N_12769,N_12351);
nand U14561 (N_14561,N_13026,N_12992);
nand U14562 (N_14562,N_12522,N_13112);
xnor U14563 (N_14563,N_12757,N_13237);
nor U14564 (N_14564,N_12882,N_12402);
xor U14565 (N_14565,N_12132,N_12867);
and U14566 (N_14566,N_12587,N_12158);
nand U14567 (N_14567,N_12881,N_12811);
xnor U14568 (N_14568,N_12274,N_13087);
or U14569 (N_14569,N_13107,N_13485);
xor U14570 (N_14570,N_12059,N_13401);
xor U14571 (N_14571,N_12201,N_13367);
or U14572 (N_14572,N_12260,N_12613);
xnor U14573 (N_14573,N_12418,N_12938);
or U14574 (N_14574,N_12120,N_12551);
nand U14575 (N_14575,N_12622,N_13267);
or U14576 (N_14576,N_12816,N_13027);
nand U14577 (N_14577,N_12471,N_12444);
and U14578 (N_14578,N_12085,N_12058);
nand U14579 (N_14579,N_12666,N_12099);
nand U14580 (N_14580,N_13256,N_12774);
xor U14581 (N_14581,N_13388,N_12337);
nand U14582 (N_14582,N_12659,N_12594);
nor U14583 (N_14583,N_12301,N_12168);
and U14584 (N_14584,N_13282,N_12355);
and U14585 (N_14585,N_13374,N_13493);
nand U14586 (N_14586,N_13224,N_13489);
nor U14587 (N_14587,N_12192,N_12891);
or U14588 (N_14588,N_12431,N_12900);
and U14589 (N_14589,N_13282,N_12745);
and U14590 (N_14590,N_12641,N_13393);
xor U14591 (N_14591,N_12533,N_12899);
xnor U14592 (N_14592,N_12481,N_12059);
nand U14593 (N_14593,N_13304,N_12885);
nand U14594 (N_14594,N_12373,N_13021);
nor U14595 (N_14595,N_12785,N_13143);
nor U14596 (N_14596,N_12293,N_13110);
or U14597 (N_14597,N_12799,N_12977);
and U14598 (N_14598,N_12513,N_12963);
nand U14599 (N_14599,N_12311,N_12129);
and U14600 (N_14600,N_12262,N_13366);
xor U14601 (N_14601,N_13227,N_12660);
xnor U14602 (N_14602,N_13424,N_12512);
xnor U14603 (N_14603,N_12240,N_12376);
nand U14604 (N_14604,N_13414,N_13101);
nand U14605 (N_14605,N_12597,N_12026);
nor U14606 (N_14606,N_12316,N_12966);
xor U14607 (N_14607,N_12214,N_12774);
nand U14608 (N_14608,N_13301,N_13183);
nor U14609 (N_14609,N_12436,N_12897);
nor U14610 (N_14610,N_12040,N_13406);
and U14611 (N_14611,N_12497,N_12163);
and U14612 (N_14612,N_12544,N_12754);
or U14613 (N_14613,N_12834,N_13324);
nor U14614 (N_14614,N_12553,N_13106);
or U14615 (N_14615,N_12215,N_12488);
nor U14616 (N_14616,N_13359,N_12291);
nand U14617 (N_14617,N_12208,N_12402);
and U14618 (N_14618,N_12086,N_12303);
or U14619 (N_14619,N_12438,N_12199);
or U14620 (N_14620,N_12497,N_12266);
nor U14621 (N_14621,N_12798,N_12926);
or U14622 (N_14622,N_13035,N_13154);
nand U14623 (N_14623,N_12418,N_13452);
nand U14624 (N_14624,N_12112,N_13013);
or U14625 (N_14625,N_12541,N_12316);
and U14626 (N_14626,N_13407,N_13195);
nor U14627 (N_14627,N_12113,N_13396);
or U14628 (N_14628,N_12519,N_12559);
xnor U14629 (N_14629,N_13137,N_12540);
nor U14630 (N_14630,N_13327,N_12029);
nor U14631 (N_14631,N_12684,N_12819);
xnor U14632 (N_14632,N_12313,N_12106);
or U14633 (N_14633,N_12740,N_12593);
nor U14634 (N_14634,N_13028,N_13108);
or U14635 (N_14635,N_12232,N_13471);
nor U14636 (N_14636,N_12814,N_12035);
and U14637 (N_14637,N_13272,N_13182);
nand U14638 (N_14638,N_12300,N_12950);
and U14639 (N_14639,N_13102,N_12413);
nor U14640 (N_14640,N_12189,N_12604);
nor U14641 (N_14641,N_12488,N_12318);
xnor U14642 (N_14642,N_13001,N_13237);
nor U14643 (N_14643,N_12903,N_13027);
xor U14644 (N_14644,N_12046,N_12714);
or U14645 (N_14645,N_12767,N_12897);
nor U14646 (N_14646,N_13493,N_12102);
nand U14647 (N_14647,N_13424,N_12197);
nand U14648 (N_14648,N_13153,N_13163);
xnor U14649 (N_14649,N_12868,N_12857);
xnor U14650 (N_14650,N_12754,N_12293);
nand U14651 (N_14651,N_12673,N_12776);
nand U14652 (N_14652,N_13373,N_12920);
nor U14653 (N_14653,N_13053,N_12771);
and U14654 (N_14654,N_12846,N_13263);
nor U14655 (N_14655,N_12530,N_12170);
or U14656 (N_14656,N_12594,N_12301);
xor U14657 (N_14657,N_13056,N_13495);
or U14658 (N_14658,N_12751,N_12950);
nand U14659 (N_14659,N_13180,N_12688);
and U14660 (N_14660,N_12689,N_12019);
and U14661 (N_14661,N_12911,N_12608);
and U14662 (N_14662,N_13153,N_12053);
xnor U14663 (N_14663,N_12801,N_13299);
xnor U14664 (N_14664,N_13244,N_12128);
nand U14665 (N_14665,N_12040,N_13482);
or U14666 (N_14666,N_12854,N_12203);
nor U14667 (N_14667,N_13077,N_13268);
nor U14668 (N_14668,N_12890,N_12748);
nor U14669 (N_14669,N_12714,N_12923);
xor U14670 (N_14670,N_12698,N_12686);
xnor U14671 (N_14671,N_12289,N_12823);
nand U14672 (N_14672,N_12382,N_12274);
nand U14673 (N_14673,N_13229,N_12889);
xor U14674 (N_14674,N_12901,N_12962);
xnor U14675 (N_14675,N_12134,N_12462);
or U14676 (N_14676,N_13490,N_12429);
nand U14677 (N_14677,N_13216,N_12540);
nand U14678 (N_14678,N_13363,N_12260);
xor U14679 (N_14679,N_13271,N_13263);
or U14680 (N_14680,N_12261,N_12178);
nand U14681 (N_14681,N_12203,N_12523);
or U14682 (N_14682,N_12731,N_12032);
nor U14683 (N_14683,N_13123,N_13083);
nor U14684 (N_14684,N_12803,N_13202);
nand U14685 (N_14685,N_12439,N_12447);
nand U14686 (N_14686,N_12690,N_12345);
or U14687 (N_14687,N_12185,N_12655);
or U14688 (N_14688,N_13323,N_12201);
xor U14689 (N_14689,N_13321,N_13417);
or U14690 (N_14690,N_12723,N_12740);
or U14691 (N_14691,N_13199,N_12222);
and U14692 (N_14692,N_13151,N_12133);
nor U14693 (N_14693,N_13232,N_12283);
xnor U14694 (N_14694,N_12901,N_13216);
nor U14695 (N_14695,N_13271,N_12664);
and U14696 (N_14696,N_13493,N_13081);
xnor U14697 (N_14697,N_13443,N_12117);
xor U14698 (N_14698,N_12355,N_12511);
and U14699 (N_14699,N_13186,N_12614);
nor U14700 (N_14700,N_12680,N_12422);
nor U14701 (N_14701,N_12856,N_13277);
and U14702 (N_14702,N_12817,N_13170);
and U14703 (N_14703,N_12489,N_13016);
and U14704 (N_14704,N_13182,N_12265);
or U14705 (N_14705,N_12352,N_13167);
xnor U14706 (N_14706,N_13143,N_12998);
xor U14707 (N_14707,N_12638,N_12797);
nor U14708 (N_14708,N_12466,N_12166);
or U14709 (N_14709,N_12868,N_13343);
or U14710 (N_14710,N_13326,N_13343);
or U14711 (N_14711,N_13131,N_13156);
and U14712 (N_14712,N_13214,N_13405);
and U14713 (N_14713,N_12181,N_13228);
nor U14714 (N_14714,N_12950,N_13188);
xor U14715 (N_14715,N_13135,N_12893);
nor U14716 (N_14716,N_12923,N_13182);
and U14717 (N_14717,N_13414,N_12918);
or U14718 (N_14718,N_12088,N_12085);
xor U14719 (N_14719,N_13280,N_12499);
nor U14720 (N_14720,N_13180,N_13075);
nand U14721 (N_14721,N_12414,N_12682);
or U14722 (N_14722,N_12158,N_12733);
xor U14723 (N_14723,N_12644,N_12189);
nand U14724 (N_14724,N_12918,N_12639);
nor U14725 (N_14725,N_13265,N_13441);
xor U14726 (N_14726,N_12974,N_13273);
nor U14727 (N_14727,N_12798,N_12004);
or U14728 (N_14728,N_12370,N_13338);
or U14729 (N_14729,N_12840,N_12368);
xnor U14730 (N_14730,N_13324,N_12674);
xor U14731 (N_14731,N_12925,N_12539);
nand U14732 (N_14732,N_13205,N_13307);
and U14733 (N_14733,N_13080,N_12116);
nand U14734 (N_14734,N_12470,N_12427);
xor U14735 (N_14735,N_12803,N_13403);
or U14736 (N_14736,N_12821,N_12532);
or U14737 (N_14737,N_12931,N_12476);
nand U14738 (N_14738,N_12321,N_12198);
or U14739 (N_14739,N_12080,N_12446);
nand U14740 (N_14740,N_12519,N_12663);
nor U14741 (N_14741,N_12339,N_13206);
xnor U14742 (N_14742,N_12105,N_13274);
nor U14743 (N_14743,N_12260,N_12241);
and U14744 (N_14744,N_13436,N_12977);
and U14745 (N_14745,N_13177,N_12950);
nand U14746 (N_14746,N_12139,N_13396);
nand U14747 (N_14747,N_12912,N_12685);
or U14748 (N_14748,N_12670,N_12730);
xor U14749 (N_14749,N_12146,N_12312);
nor U14750 (N_14750,N_12391,N_12087);
or U14751 (N_14751,N_12302,N_13226);
xor U14752 (N_14752,N_13175,N_12617);
xor U14753 (N_14753,N_12003,N_12485);
and U14754 (N_14754,N_12410,N_12288);
or U14755 (N_14755,N_12858,N_12837);
nor U14756 (N_14756,N_12939,N_12696);
nand U14757 (N_14757,N_12246,N_13057);
or U14758 (N_14758,N_13049,N_12192);
or U14759 (N_14759,N_12454,N_12847);
nor U14760 (N_14760,N_12811,N_12439);
xnor U14761 (N_14761,N_12879,N_13141);
nor U14762 (N_14762,N_12706,N_12498);
nand U14763 (N_14763,N_12934,N_13387);
and U14764 (N_14764,N_12677,N_12893);
and U14765 (N_14765,N_12070,N_12069);
nand U14766 (N_14766,N_12209,N_13102);
nand U14767 (N_14767,N_12859,N_13011);
xor U14768 (N_14768,N_12813,N_12788);
nand U14769 (N_14769,N_13180,N_13476);
and U14770 (N_14770,N_12098,N_13108);
xor U14771 (N_14771,N_13207,N_12038);
nand U14772 (N_14772,N_12693,N_12527);
or U14773 (N_14773,N_12249,N_13328);
nand U14774 (N_14774,N_12436,N_12074);
nor U14775 (N_14775,N_12095,N_12468);
and U14776 (N_14776,N_12545,N_13225);
nand U14777 (N_14777,N_13025,N_12432);
nand U14778 (N_14778,N_12116,N_13444);
xnor U14779 (N_14779,N_12749,N_13075);
and U14780 (N_14780,N_12414,N_12907);
nand U14781 (N_14781,N_13463,N_12966);
and U14782 (N_14782,N_12229,N_12227);
nor U14783 (N_14783,N_12996,N_12241);
nor U14784 (N_14784,N_12760,N_12851);
and U14785 (N_14785,N_12250,N_12667);
xor U14786 (N_14786,N_12223,N_12351);
xor U14787 (N_14787,N_12800,N_12707);
xnor U14788 (N_14788,N_12040,N_12527);
and U14789 (N_14789,N_13245,N_12994);
and U14790 (N_14790,N_13341,N_13264);
nand U14791 (N_14791,N_13463,N_13130);
xor U14792 (N_14792,N_12212,N_12215);
or U14793 (N_14793,N_12698,N_12881);
and U14794 (N_14794,N_13215,N_12218);
or U14795 (N_14795,N_13225,N_13197);
or U14796 (N_14796,N_12224,N_12053);
nor U14797 (N_14797,N_12507,N_12865);
nand U14798 (N_14798,N_12124,N_12610);
and U14799 (N_14799,N_12258,N_12780);
nor U14800 (N_14800,N_12106,N_12810);
or U14801 (N_14801,N_12277,N_13336);
nand U14802 (N_14802,N_12723,N_13385);
nor U14803 (N_14803,N_13153,N_12829);
xnor U14804 (N_14804,N_12843,N_13093);
nand U14805 (N_14805,N_13364,N_12795);
nor U14806 (N_14806,N_13093,N_13003);
nor U14807 (N_14807,N_13184,N_12975);
and U14808 (N_14808,N_12469,N_12950);
xor U14809 (N_14809,N_12859,N_12697);
or U14810 (N_14810,N_12505,N_13001);
nor U14811 (N_14811,N_12408,N_12318);
and U14812 (N_14812,N_12729,N_12287);
nand U14813 (N_14813,N_12835,N_12090);
xor U14814 (N_14814,N_12841,N_12725);
xnor U14815 (N_14815,N_12012,N_13144);
and U14816 (N_14816,N_12278,N_12834);
nor U14817 (N_14817,N_12855,N_12618);
nor U14818 (N_14818,N_12492,N_12663);
or U14819 (N_14819,N_12827,N_13279);
nor U14820 (N_14820,N_13263,N_12788);
xor U14821 (N_14821,N_12643,N_13384);
and U14822 (N_14822,N_13120,N_13228);
xor U14823 (N_14823,N_12861,N_13019);
nor U14824 (N_14824,N_12588,N_12604);
or U14825 (N_14825,N_13017,N_12058);
and U14826 (N_14826,N_12337,N_12331);
or U14827 (N_14827,N_12323,N_13248);
nor U14828 (N_14828,N_12896,N_13494);
and U14829 (N_14829,N_13058,N_13013);
nand U14830 (N_14830,N_12084,N_13195);
xor U14831 (N_14831,N_13027,N_12893);
or U14832 (N_14832,N_12534,N_13467);
nand U14833 (N_14833,N_13046,N_13187);
nor U14834 (N_14834,N_12536,N_12668);
nand U14835 (N_14835,N_13329,N_12130);
and U14836 (N_14836,N_12026,N_12802);
and U14837 (N_14837,N_12045,N_13419);
and U14838 (N_14838,N_12804,N_13407);
nor U14839 (N_14839,N_13347,N_12704);
or U14840 (N_14840,N_13466,N_12994);
or U14841 (N_14841,N_12051,N_12493);
nand U14842 (N_14842,N_13125,N_12721);
nor U14843 (N_14843,N_13020,N_12552);
nor U14844 (N_14844,N_12341,N_13316);
xor U14845 (N_14845,N_13209,N_12806);
nand U14846 (N_14846,N_12234,N_13448);
nor U14847 (N_14847,N_12505,N_12879);
and U14848 (N_14848,N_13011,N_12581);
or U14849 (N_14849,N_13347,N_12564);
xor U14850 (N_14850,N_13367,N_13070);
nor U14851 (N_14851,N_12437,N_12660);
or U14852 (N_14852,N_12131,N_12192);
or U14853 (N_14853,N_12402,N_13034);
nor U14854 (N_14854,N_12667,N_12641);
or U14855 (N_14855,N_12257,N_12276);
xor U14856 (N_14856,N_13205,N_12838);
or U14857 (N_14857,N_12584,N_12064);
nand U14858 (N_14858,N_13040,N_13374);
nand U14859 (N_14859,N_13476,N_13319);
and U14860 (N_14860,N_13465,N_12153);
nand U14861 (N_14861,N_12352,N_12555);
nor U14862 (N_14862,N_12264,N_12535);
nand U14863 (N_14863,N_12562,N_12256);
xor U14864 (N_14864,N_13019,N_12164);
nor U14865 (N_14865,N_12180,N_12045);
nor U14866 (N_14866,N_12384,N_12333);
and U14867 (N_14867,N_12915,N_12851);
xnor U14868 (N_14868,N_13354,N_13005);
nand U14869 (N_14869,N_12135,N_13139);
or U14870 (N_14870,N_13447,N_12650);
xor U14871 (N_14871,N_13222,N_12983);
nand U14872 (N_14872,N_12661,N_12672);
and U14873 (N_14873,N_13361,N_13284);
nand U14874 (N_14874,N_12634,N_12385);
nor U14875 (N_14875,N_12508,N_13321);
or U14876 (N_14876,N_12197,N_12912);
xor U14877 (N_14877,N_12498,N_13009);
and U14878 (N_14878,N_12325,N_12050);
or U14879 (N_14879,N_12734,N_12864);
nand U14880 (N_14880,N_12359,N_13276);
nor U14881 (N_14881,N_12118,N_12850);
xor U14882 (N_14882,N_12701,N_12895);
or U14883 (N_14883,N_13015,N_12036);
or U14884 (N_14884,N_12795,N_12937);
xor U14885 (N_14885,N_12934,N_12833);
nand U14886 (N_14886,N_12373,N_13408);
nor U14887 (N_14887,N_13072,N_13152);
nand U14888 (N_14888,N_12145,N_13134);
xor U14889 (N_14889,N_12875,N_13219);
or U14890 (N_14890,N_13192,N_13235);
nand U14891 (N_14891,N_13252,N_12677);
nor U14892 (N_14892,N_12433,N_12154);
xnor U14893 (N_14893,N_13006,N_13303);
or U14894 (N_14894,N_13043,N_12229);
and U14895 (N_14895,N_12839,N_12635);
or U14896 (N_14896,N_12639,N_12251);
xor U14897 (N_14897,N_13217,N_12390);
nand U14898 (N_14898,N_12308,N_12187);
nor U14899 (N_14899,N_12299,N_12965);
or U14900 (N_14900,N_12894,N_13441);
nand U14901 (N_14901,N_12518,N_12058);
and U14902 (N_14902,N_12808,N_13491);
nor U14903 (N_14903,N_13356,N_12184);
nand U14904 (N_14904,N_12932,N_12698);
nand U14905 (N_14905,N_13471,N_12997);
xnor U14906 (N_14906,N_13243,N_13149);
or U14907 (N_14907,N_12904,N_13041);
and U14908 (N_14908,N_12629,N_12162);
and U14909 (N_14909,N_12412,N_13065);
nor U14910 (N_14910,N_12939,N_13245);
nand U14911 (N_14911,N_12535,N_13169);
nand U14912 (N_14912,N_12651,N_12256);
nand U14913 (N_14913,N_13116,N_12336);
xnor U14914 (N_14914,N_13343,N_13247);
or U14915 (N_14915,N_12588,N_12475);
and U14916 (N_14916,N_12048,N_13233);
xnor U14917 (N_14917,N_13032,N_13364);
and U14918 (N_14918,N_13067,N_12090);
or U14919 (N_14919,N_13121,N_12462);
nand U14920 (N_14920,N_12022,N_13301);
nand U14921 (N_14921,N_12369,N_13292);
or U14922 (N_14922,N_13460,N_13338);
xor U14923 (N_14923,N_12860,N_12002);
nand U14924 (N_14924,N_12499,N_13408);
xnor U14925 (N_14925,N_13026,N_12978);
nor U14926 (N_14926,N_12062,N_12626);
or U14927 (N_14927,N_12733,N_12663);
nand U14928 (N_14928,N_13006,N_12460);
xnor U14929 (N_14929,N_12458,N_12423);
xnor U14930 (N_14930,N_12573,N_13210);
nand U14931 (N_14931,N_12935,N_13026);
xnor U14932 (N_14932,N_13371,N_12228);
or U14933 (N_14933,N_13094,N_12019);
xor U14934 (N_14934,N_12866,N_12833);
xor U14935 (N_14935,N_12957,N_12339);
nand U14936 (N_14936,N_12376,N_13390);
nand U14937 (N_14937,N_13046,N_12252);
or U14938 (N_14938,N_12473,N_12105);
xnor U14939 (N_14939,N_13216,N_12602);
nand U14940 (N_14940,N_13396,N_12353);
or U14941 (N_14941,N_13240,N_12129);
nor U14942 (N_14942,N_12928,N_12628);
or U14943 (N_14943,N_12833,N_12666);
nor U14944 (N_14944,N_12370,N_12721);
and U14945 (N_14945,N_12605,N_13436);
or U14946 (N_14946,N_13427,N_12888);
or U14947 (N_14947,N_13117,N_12292);
or U14948 (N_14948,N_12458,N_13373);
and U14949 (N_14949,N_12779,N_12002);
or U14950 (N_14950,N_12041,N_12669);
or U14951 (N_14951,N_13005,N_13194);
nand U14952 (N_14952,N_13227,N_13494);
and U14953 (N_14953,N_12058,N_13268);
or U14954 (N_14954,N_12097,N_12728);
and U14955 (N_14955,N_12177,N_13322);
nor U14956 (N_14956,N_12975,N_12182);
xor U14957 (N_14957,N_13197,N_12542);
nand U14958 (N_14958,N_12935,N_12900);
or U14959 (N_14959,N_12301,N_12240);
or U14960 (N_14960,N_13366,N_12749);
nand U14961 (N_14961,N_13403,N_13098);
and U14962 (N_14962,N_13010,N_13315);
nor U14963 (N_14963,N_12389,N_13031);
or U14964 (N_14964,N_12020,N_12108);
nor U14965 (N_14965,N_12730,N_13119);
or U14966 (N_14966,N_12399,N_12003);
xor U14967 (N_14967,N_12028,N_12768);
nor U14968 (N_14968,N_13321,N_12986);
nand U14969 (N_14969,N_12408,N_12353);
or U14970 (N_14970,N_13419,N_12994);
nand U14971 (N_14971,N_13156,N_12185);
nand U14972 (N_14972,N_12689,N_12280);
nand U14973 (N_14973,N_12087,N_12224);
nor U14974 (N_14974,N_13338,N_12040);
nand U14975 (N_14975,N_12024,N_13291);
xnor U14976 (N_14976,N_12633,N_13468);
nand U14977 (N_14977,N_13018,N_12440);
xnor U14978 (N_14978,N_13049,N_12969);
xnor U14979 (N_14979,N_12142,N_12448);
or U14980 (N_14980,N_12442,N_13337);
nand U14981 (N_14981,N_12527,N_12240);
and U14982 (N_14982,N_13488,N_12341);
or U14983 (N_14983,N_12739,N_12053);
nor U14984 (N_14984,N_12790,N_12676);
and U14985 (N_14985,N_12116,N_12824);
and U14986 (N_14986,N_13425,N_12367);
xor U14987 (N_14987,N_13099,N_12506);
nor U14988 (N_14988,N_12372,N_13317);
xnor U14989 (N_14989,N_12684,N_12302);
and U14990 (N_14990,N_13078,N_12086);
nor U14991 (N_14991,N_13292,N_12616);
nand U14992 (N_14992,N_12381,N_12170);
or U14993 (N_14993,N_12035,N_12044);
nand U14994 (N_14994,N_12051,N_13237);
nand U14995 (N_14995,N_13362,N_12006);
or U14996 (N_14996,N_12866,N_12948);
and U14997 (N_14997,N_12977,N_12651);
xor U14998 (N_14998,N_13303,N_12115);
nor U14999 (N_14999,N_12407,N_12633);
nand UO_0 (O_0,N_14982,N_14842);
and UO_1 (O_1,N_14456,N_14552);
nand UO_2 (O_2,N_14774,N_13704);
nor UO_3 (O_3,N_13895,N_14018);
and UO_4 (O_4,N_14191,N_13852);
or UO_5 (O_5,N_13606,N_13943);
and UO_6 (O_6,N_14492,N_14983);
xor UO_7 (O_7,N_14036,N_14439);
or UO_8 (O_8,N_13619,N_14912);
xor UO_9 (O_9,N_14985,N_13514);
xor UO_10 (O_10,N_14940,N_14825);
nor UO_11 (O_11,N_13611,N_13995);
nor UO_12 (O_12,N_13787,N_13925);
or UO_13 (O_13,N_13693,N_14088);
nor UO_14 (O_14,N_13939,N_14909);
or UO_15 (O_15,N_14617,N_14645);
nor UO_16 (O_16,N_14213,N_13894);
or UO_17 (O_17,N_14103,N_13622);
xor UO_18 (O_18,N_14901,N_14202);
xnor UO_19 (O_19,N_14053,N_14276);
nor UO_20 (O_20,N_14206,N_14557);
or UO_21 (O_21,N_14768,N_13518);
and UO_22 (O_22,N_14190,N_13836);
or UO_23 (O_23,N_14111,N_14736);
nand UO_24 (O_24,N_14179,N_14833);
and UO_25 (O_25,N_13569,N_14859);
or UO_26 (O_26,N_14561,N_13978);
nor UO_27 (O_27,N_14042,N_14091);
nor UO_28 (O_28,N_14619,N_13535);
nor UO_29 (O_29,N_14291,N_14586);
or UO_30 (O_30,N_14994,N_14177);
nand UO_31 (O_31,N_13557,N_13631);
and UO_32 (O_32,N_14851,N_14393);
nor UO_33 (O_33,N_14476,N_14612);
or UO_34 (O_34,N_14641,N_14563);
nand UO_35 (O_35,N_13809,N_13563);
nor UO_36 (O_36,N_13603,N_14565);
nand UO_37 (O_37,N_13769,N_14237);
xnor UO_38 (O_38,N_13820,N_13792);
nor UO_39 (O_39,N_14231,N_13899);
or UO_40 (O_40,N_13979,N_14220);
nand UO_41 (O_41,N_14418,N_14265);
and UO_42 (O_42,N_14693,N_13878);
xor UO_43 (O_43,N_14654,N_14081);
nor UO_44 (O_44,N_14322,N_13758);
and UO_45 (O_45,N_14482,N_14333);
nor UO_46 (O_46,N_14382,N_13813);
or UO_47 (O_47,N_14343,N_14584);
xnor UO_48 (O_48,N_14351,N_13969);
xnor UO_49 (O_49,N_14970,N_14942);
nand UO_50 (O_50,N_13972,N_14678);
xnor UO_51 (O_51,N_13691,N_14757);
xnor UO_52 (O_52,N_14426,N_13613);
nand UO_53 (O_53,N_14271,N_13651);
xor UO_54 (O_54,N_14717,N_13519);
nand UO_55 (O_55,N_14871,N_14251);
nor UO_56 (O_56,N_13621,N_14246);
or UO_57 (O_57,N_13729,N_14958);
xor UO_58 (O_58,N_14181,N_13749);
and UO_59 (O_59,N_14010,N_14473);
and UO_60 (O_60,N_14372,N_14708);
nor UO_61 (O_61,N_14498,N_14039);
and UO_62 (O_62,N_13774,N_14315);
nand UO_63 (O_63,N_13879,N_14420);
nor UO_64 (O_64,N_13529,N_14437);
nor UO_65 (O_65,N_13964,N_14021);
or UO_66 (O_66,N_13703,N_14793);
or UO_67 (O_67,N_13659,N_14258);
nor UO_68 (O_68,N_14361,N_14579);
or UO_69 (O_69,N_13928,N_13791);
xor UO_70 (O_70,N_14688,N_13949);
or UO_71 (O_71,N_14150,N_14178);
nor UO_72 (O_72,N_14417,N_14301);
nor UO_73 (O_73,N_14935,N_14822);
nor UO_74 (O_74,N_14628,N_13628);
nand UO_75 (O_75,N_14542,N_14978);
and UO_76 (O_76,N_14357,N_14742);
nand UO_77 (O_77,N_14622,N_14256);
and UO_78 (O_78,N_14931,N_14033);
nor UO_79 (O_79,N_14120,N_13762);
xnor UO_80 (O_80,N_13892,N_14187);
xor UO_81 (O_81,N_13641,N_14288);
and UO_82 (O_82,N_14649,N_14588);
and UO_83 (O_83,N_13881,N_14199);
nor UO_84 (O_84,N_14997,N_13980);
xor UO_85 (O_85,N_13540,N_14795);
xnor UO_86 (O_86,N_14841,N_14151);
nor UO_87 (O_87,N_14594,N_13745);
nor UO_88 (O_88,N_14124,N_14041);
nand UO_89 (O_89,N_14723,N_13847);
nand UO_90 (O_90,N_13977,N_14433);
nor UO_91 (O_91,N_14303,N_13545);
nor UO_92 (O_92,N_14149,N_14950);
nor UO_93 (O_93,N_13757,N_14380);
or UO_94 (O_94,N_13629,N_14434);
nand UO_95 (O_95,N_14758,N_14442);
xnor UO_96 (O_96,N_14059,N_13921);
and UO_97 (O_97,N_14674,N_14672);
and UO_98 (O_98,N_13526,N_14268);
nand UO_99 (O_99,N_14530,N_14536);
nor UO_100 (O_100,N_14740,N_14196);
or UO_101 (O_101,N_13826,N_13929);
and UO_102 (O_102,N_14703,N_14129);
and UO_103 (O_103,N_14142,N_13576);
or UO_104 (O_104,N_14948,N_14496);
nand UO_105 (O_105,N_14786,N_13864);
xnor UO_106 (O_106,N_14780,N_14014);
and UO_107 (O_107,N_13827,N_14153);
xor UO_108 (O_108,N_14429,N_14131);
xnor UO_109 (O_109,N_14720,N_14847);
or UO_110 (O_110,N_14567,N_14082);
or UO_111 (O_111,N_14028,N_14828);
or UO_112 (O_112,N_13633,N_14020);
xnor UO_113 (O_113,N_14309,N_14943);
nand UO_114 (O_114,N_14304,N_13687);
and UO_115 (O_115,N_14779,N_13642);
nand UO_116 (O_116,N_14870,N_14646);
and UO_117 (O_117,N_14696,N_14218);
nor UO_118 (O_118,N_14527,N_14173);
nor UO_119 (O_119,N_14174,N_13962);
nand UO_120 (O_120,N_14752,N_14918);
or UO_121 (O_121,N_14419,N_14585);
and UO_122 (O_122,N_13866,N_14085);
or UO_123 (O_123,N_14972,N_14069);
or UO_124 (O_124,N_14478,N_13507);
or UO_125 (O_125,N_14394,N_13688);
xnor UO_126 (O_126,N_13844,N_14171);
or UO_127 (O_127,N_14182,N_14423);
nand UO_128 (O_128,N_14250,N_13912);
and UO_129 (O_129,N_14753,N_14575);
and UO_130 (O_130,N_13503,N_14548);
nor UO_131 (O_131,N_14876,N_13671);
and UO_132 (O_132,N_13824,N_13948);
or UO_133 (O_133,N_14805,N_14262);
or UO_134 (O_134,N_14000,N_14656);
xnor UO_135 (O_135,N_14049,N_13920);
or UO_136 (O_136,N_13586,N_13654);
xnor UO_137 (O_137,N_13875,N_13889);
and UO_138 (O_138,N_14440,N_13931);
nor UO_139 (O_139,N_14247,N_14381);
nor UO_140 (O_140,N_13910,N_13656);
xor UO_141 (O_141,N_13989,N_14292);
xor UO_142 (O_142,N_14311,N_14454);
and UO_143 (O_143,N_13635,N_14992);
nor UO_144 (O_144,N_14733,N_13560);
nor UO_145 (O_145,N_14669,N_14580);
nand UO_146 (O_146,N_14308,N_14705);
or UO_147 (O_147,N_13616,N_13763);
and UO_148 (O_148,N_13793,N_14624);
nor UO_149 (O_149,N_14186,N_14868);
or UO_150 (O_150,N_13788,N_13686);
or UO_151 (O_151,N_13950,N_14812);
nand UO_152 (O_152,N_14759,N_14260);
nor UO_153 (O_153,N_14813,N_14274);
and UO_154 (O_154,N_14852,N_14684);
nor UO_155 (O_155,N_13823,N_14406);
xnor UO_156 (O_156,N_14501,N_14694);
or UO_157 (O_157,N_14378,N_14883);
xnor UO_158 (O_158,N_14620,N_13834);
or UO_159 (O_159,N_14517,N_14508);
xor UO_160 (O_160,N_14076,N_14254);
nand UO_161 (O_161,N_14269,N_14286);
xnor UO_162 (O_162,N_14031,N_14718);
xor UO_163 (O_163,N_14449,N_14494);
or UO_164 (O_164,N_13802,N_13850);
nor UO_165 (O_165,N_13590,N_14067);
nor UO_166 (O_166,N_14762,N_14407);
nand UO_167 (O_167,N_14928,N_14077);
and UO_168 (O_168,N_14468,N_14116);
xor UO_169 (O_169,N_14354,N_14306);
and UO_170 (O_170,N_14167,N_14305);
xnor UO_171 (O_171,N_14615,N_14648);
xnor UO_172 (O_172,N_14377,N_13551);
nor UO_173 (O_173,N_14763,N_14092);
or UO_174 (O_174,N_14959,N_14317);
nor UO_175 (O_175,N_13500,N_14232);
and UO_176 (O_176,N_14829,N_14865);
xnor UO_177 (O_177,N_13799,N_13644);
and UO_178 (O_178,N_13668,N_14836);
and UO_179 (O_179,N_14906,N_13754);
nand UO_180 (O_180,N_14112,N_13807);
nand UO_181 (O_181,N_13991,N_13942);
nand UO_182 (O_182,N_13657,N_13814);
nor UO_183 (O_183,N_13821,N_14110);
xor UO_184 (O_184,N_14373,N_13672);
or UO_185 (O_185,N_13940,N_13731);
nand UO_186 (O_186,N_14511,N_13832);
xnor UO_187 (O_187,N_14332,N_13679);
nor UO_188 (O_188,N_13699,N_14556);
nand UO_189 (O_189,N_13601,N_13845);
nor UO_190 (O_190,N_14801,N_14485);
and UO_191 (O_191,N_14491,N_13857);
and UO_192 (O_192,N_13747,N_14045);
or UO_193 (O_193,N_14570,N_14070);
or UO_194 (O_194,N_14566,N_14510);
xor UO_195 (O_195,N_14529,N_14497);
or UO_196 (O_196,N_14375,N_14991);
and UO_197 (O_197,N_14690,N_14706);
xor UO_198 (O_198,N_13626,N_14714);
xor UO_199 (O_199,N_14798,N_14143);
and UO_200 (O_200,N_13843,N_14969);
nand UO_201 (O_201,N_13573,N_14209);
or UO_202 (O_202,N_14610,N_14412);
nor UO_203 (O_203,N_14119,N_14760);
or UO_204 (O_204,N_14259,N_14233);
nor UO_205 (O_205,N_13682,N_14858);
and UO_206 (O_206,N_14105,N_14387);
xnor UO_207 (O_207,N_14152,N_14633);
nor UO_208 (O_208,N_14154,N_13968);
nor UO_209 (O_209,N_13930,N_14904);
nor UO_210 (O_210,N_14545,N_13524);
or UO_211 (O_211,N_14810,N_14503);
xor UO_212 (O_212,N_13527,N_14936);
nor UO_213 (O_213,N_14448,N_13959);
or UO_214 (O_214,N_14896,N_13795);
and UO_215 (O_215,N_14724,N_14789);
nand UO_216 (O_216,N_14242,N_14058);
and UO_217 (O_217,N_13963,N_13650);
nor UO_218 (O_218,N_14682,N_13746);
and UO_219 (O_219,N_14846,N_14138);
nand UO_220 (O_220,N_14574,N_14653);
and UO_221 (O_221,N_14791,N_14629);
or UO_222 (O_222,N_14804,N_14219);
nand UO_223 (O_223,N_14626,N_14095);
xnor UO_224 (O_224,N_13708,N_14662);
and UO_225 (O_225,N_13860,N_14834);
nor UO_226 (O_226,N_13753,N_14692);
or UO_227 (O_227,N_13781,N_14782);
xnor UO_228 (O_228,N_14344,N_14438);
nand UO_229 (O_229,N_14908,N_13865);
nand UO_230 (O_230,N_14012,N_13984);
xor UO_231 (O_231,N_14287,N_14115);
and UO_232 (O_232,N_14686,N_14083);
nand UO_233 (O_233,N_14593,N_13610);
or UO_234 (O_234,N_14026,N_13734);
or UO_235 (O_235,N_14680,N_13805);
nand UO_236 (O_236,N_13591,N_14880);
or UO_237 (O_237,N_14401,N_13579);
nand UO_238 (O_238,N_14605,N_14980);
nand UO_239 (O_239,N_14981,N_13660);
nor UO_240 (O_240,N_14356,N_13662);
nor UO_241 (O_241,N_13596,N_13649);
nand UO_242 (O_242,N_14873,N_14374);
nand UO_243 (O_243,N_13508,N_14891);
nor UO_244 (O_244,N_14100,N_14872);
and UO_245 (O_245,N_14974,N_14685);
or UO_246 (O_246,N_13770,N_13897);
xor UO_247 (O_247,N_14389,N_14596);
nand UO_248 (O_248,N_14683,N_13741);
or UO_249 (O_249,N_14734,N_13869);
nor UO_250 (O_250,N_13789,N_13967);
and UO_251 (O_251,N_14318,N_14073);
xnor UO_252 (O_252,N_14408,N_13760);
xnor UO_253 (O_253,N_14272,N_14721);
nor UO_254 (O_254,N_13880,N_14535);
or UO_255 (O_255,N_14197,N_14400);
or UO_256 (O_256,N_14993,N_14790);
and UO_257 (O_257,N_13882,N_14651);
and UO_258 (O_258,N_14298,N_13550);
xnor UO_259 (O_259,N_14634,N_14043);
and UO_260 (O_260,N_14544,N_13504);
nor UO_261 (O_261,N_14207,N_13811);
nor UO_262 (O_262,N_13988,N_13740);
or UO_263 (O_263,N_13511,N_14074);
xnor UO_264 (O_264,N_14471,N_14062);
nor UO_265 (O_265,N_14821,N_14409);
xnor UO_266 (O_266,N_13521,N_14513);
xor UO_267 (O_267,N_13785,N_14702);
nor UO_268 (O_268,N_13572,N_14032);
and UO_269 (O_269,N_14211,N_13965);
or UO_270 (O_270,N_14583,N_14236);
nor UO_271 (O_271,N_14384,N_14848);
nand UO_272 (O_272,N_13893,N_14787);
xor UO_273 (O_273,N_14297,N_13604);
nand UO_274 (O_274,N_13825,N_14845);
and UO_275 (O_275,N_13607,N_14314);
nand UO_276 (O_276,N_13822,N_13851);
xor UO_277 (O_277,N_13808,N_14888);
xnor UO_278 (O_278,N_14338,N_14413);
xnor UO_279 (O_279,N_14360,N_14118);
and UO_280 (O_280,N_13653,N_14457);
or UO_281 (O_281,N_13539,N_14358);
nor UO_282 (O_282,N_13743,N_13849);
or UO_283 (O_283,N_13568,N_14516);
and UO_284 (O_284,N_13618,N_14266);
xnor UO_285 (O_285,N_13970,N_14145);
or UO_286 (O_286,N_14961,N_14097);
or UO_287 (O_287,N_13830,N_13617);
nor UO_288 (O_288,N_14144,N_14163);
or UO_289 (O_289,N_14553,N_13971);
nor UO_290 (O_290,N_13531,N_14331);
nand UO_291 (O_291,N_14212,N_13625);
or UO_292 (O_292,N_13800,N_14486);
and UO_293 (O_293,N_14743,N_14345);
nor UO_294 (O_294,N_13537,N_13755);
xnor UO_295 (O_295,N_13523,N_13509);
nand UO_296 (O_296,N_13707,N_14293);
or UO_297 (O_297,N_14956,N_13870);
xor UO_298 (O_298,N_14860,N_13914);
and UO_299 (O_299,N_14296,N_14528);
and UO_300 (O_300,N_14355,N_13839);
nor UO_301 (O_301,N_14899,N_13953);
or UO_302 (O_302,N_14534,N_14493);
and UO_303 (O_303,N_14507,N_14295);
xnor UO_304 (O_304,N_14136,N_13666);
nor UO_305 (O_305,N_13555,N_14953);
or UO_306 (O_306,N_14745,N_14934);
nand UO_307 (O_307,N_14932,N_14630);
and UO_308 (O_308,N_14521,N_14679);
nand UO_309 (O_309,N_13549,N_14160);
nor UO_310 (O_310,N_13876,N_14455);
or UO_311 (O_311,N_14270,N_14965);
nand UO_312 (O_312,N_13713,N_14595);
xnor UO_313 (O_313,N_13567,N_13501);
nand UO_314 (O_314,N_14427,N_13609);
xor UO_315 (O_315,N_14328,N_14764);
and UO_316 (O_316,N_14807,N_14464);
xor UO_317 (O_317,N_14778,N_14551);
and UO_318 (O_318,N_14506,N_13934);
nand UO_319 (O_319,N_13623,N_14664);
and UO_320 (O_320,N_14363,N_13717);
xor UO_321 (O_321,N_14255,N_13548);
nand UO_322 (O_322,N_14892,N_14435);
or UO_323 (O_323,N_14155,N_13883);
xor UO_324 (O_324,N_13946,N_14558);
nor UO_325 (O_325,N_14346,N_13999);
nand UO_326 (O_326,N_14016,N_14830);
and UO_327 (O_327,N_14184,N_14359);
nand UO_328 (O_328,N_14897,N_13938);
nand UO_329 (O_329,N_14336,N_13571);
or UO_330 (O_330,N_14707,N_13715);
and UO_331 (O_331,N_14907,N_13846);
xnor UO_332 (O_332,N_14227,N_14766);
xnor UO_333 (O_333,N_13562,N_13855);
and UO_334 (O_334,N_13896,N_13819);
and UO_335 (O_335,N_14243,N_14137);
nor UO_336 (O_336,N_14792,N_13801);
nor UO_337 (O_337,N_14302,N_13775);
nand UO_338 (O_338,N_14108,N_14221);
nor UO_339 (O_339,N_14424,N_14564);
or UO_340 (O_340,N_14712,N_13605);
or UO_341 (O_341,N_14923,N_13905);
xor UO_342 (O_342,N_13552,N_14771);
and UO_343 (O_343,N_14979,N_14023);
xor UO_344 (O_344,N_14660,N_14327);
or UO_345 (O_345,N_14546,N_13690);
nor UO_346 (O_346,N_14422,N_14109);
and UO_347 (O_347,N_14446,N_13574);
nand UO_348 (O_348,N_13887,N_14189);
nor UO_349 (O_349,N_14550,N_14093);
and UO_350 (O_350,N_14937,N_14921);
nand UO_351 (O_351,N_14616,N_14253);
nor UO_352 (O_352,N_14040,N_14903);
or UO_353 (O_353,N_14863,N_14898);
nor UO_354 (O_354,N_14307,N_14135);
nor UO_355 (O_355,N_14554,N_14035);
nor UO_356 (O_356,N_14915,N_14671);
or UO_357 (O_357,N_14540,N_14484);
nor UO_358 (O_358,N_14938,N_13673);
nor UO_359 (O_359,N_13646,N_14451);
nor UO_360 (O_360,N_13674,N_14738);
xor UO_361 (O_361,N_13522,N_13599);
nor UO_362 (O_362,N_14371,N_14240);
nor UO_363 (O_363,N_13890,N_14668);
nand UO_364 (O_364,N_13675,N_13685);
or UO_365 (O_365,N_14902,N_13658);
xnor UO_366 (O_366,N_14465,N_13541);
nor UO_367 (O_367,N_14663,N_14239);
or UO_368 (O_368,N_14725,N_14224);
nor UO_369 (O_369,N_14831,N_14495);
and UO_370 (O_370,N_14019,N_14323);
nand UO_371 (O_371,N_13737,N_14955);
or UO_372 (O_372,N_14391,N_14541);
and UO_373 (O_373,N_14447,N_14827);
and UO_374 (O_374,N_13561,N_14319);
nand UO_375 (O_375,N_14749,N_14816);
or UO_376 (O_376,N_14509,N_14500);
nand UO_377 (O_377,N_14106,N_13833);
or UO_378 (O_378,N_14430,N_14261);
nor UO_379 (O_379,N_14013,N_13724);
nor UO_380 (O_380,N_13736,N_13692);
or UO_381 (O_381,N_13994,N_14367);
nand UO_382 (O_382,N_14230,N_13877);
nand UO_383 (O_383,N_13922,N_13652);
or UO_384 (O_384,N_14800,N_14676);
xor UO_385 (O_385,N_13790,N_14263);
or UO_386 (O_386,N_14123,N_14125);
and UO_387 (O_387,N_14056,N_14647);
or UO_388 (O_388,N_13764,N_14655);
xor UO_389 (O_389,N_14887,N_13584);
xnor UO_390 (O_390,N_13945,N_14637);
nor UO_391 (O_391,N_13676,N_14329);
or UO_392 (O_392,N_14882,N_14364);
and UO_393 (O_393,N_14783,N_14857);
and UO_394 (O_394,N_14313,N_14603);
or UO_395 (O_395,N_14889,N_14470);
nand UO_396 (O_396,N_13702,N_14954);
xnor UO_397 (O_397,N_13992,N_14576);
nand UO_398 (O_398,N_14957,N_14927);
and UO_399 (O_399,N_14735,N_14537);
xnor UO_400 (O_400,N_14525,N_14582);
or UO_401 (O_401,N_14397,N_14117);
and UO_402 (O_402,N_13638,N_13798);
and UO_403 (O_403,N_13806,N_13716);
nor UO_404 (O_404,N_14555,N_14238);
xnor UO_405 (O_405,N_14611,N_14754);
nand UO_406 (O_406,N_14055,N_14919);
xor UO_407 (O_407,N_14063,N_14988);
or UO_408 (O_408,N_13547,N_13722);
nand UO_409 (O_409,N_14689,N_14627);
and UO_410 (O_410,N_14729,N_14017);
or UO_411 (O_411,N_13816,N_13543);
xor UO_412 (O_412,N_14638,N_14002);
and UO_413 (O_413,N_14716,N_14929);
nor UO_414 (O_414,N_14518,N_14569);
nand UO_415 (O_415,N_14414,N_14597);
or UO_416 (O_416,N_14463,N_14573);
nor UO_417 (O_417,N_14078,N_13927);
nand UO_418 (O_418,N_13553,N_13612);
and UO_419 (O_419,N_14879,N_13782);
nor UO_420 (O_420,N_14472,N_14445);
xor UO_421 (O_421,N_14670,N_14282);
and UO_422 (O_422,N_14425,N_14699);
and UO_423 (O_423,N_13771,N_13528);
or UO_424 (O_424,N_13947,N_14205);
nor UO_425 (O_425,N_13854,N_14549);
nor UO_426 (O_426,N_13624,N_14204);
or UO_427 (O_427,N_14046,N_13630);
or UO_428 (O_428,N_14850,N_14966);
and UO_429 (O_429,N_14312,N_14913);
nand UO_430 (O_430,N_13648,N_14607);
nand UO_431 (O_431,N_14411,N_14175);
xor UO_432 (O_432,N_14875,N_14975);
xor UO_433 (O_433,N_14223,N_13780);
xnor UO_434 (O_434,N_13502,N_14784);
or UO_435 (O_435,N_14681,N_14608);
nand UO_436 (O_436,N_14618,N_14215);
nor UO_437 (O_437,N_14794,N_14390);
xor UO_438 (O_438,N_14170,N_14458);
xnor UO_439 (O_439,N_13935,N_14949);
xor UO_440 (O_440,N_14443,N_13564);
nand UO_441 (O_441,N_14996,N_14631);
nor UO_442 (O_442,N_13768,N_14166);
and UO_443 (O_443,N_13706,N_13918);
xnor UO_444 (O_444,N_14700,N_13570);
nor UO_445 (O_445,N_13634,N_13627);
and UO_446 (O_446,N_13554,N_14941);
xnor UO_447 (O_447,N_13538,N_14973);
nand UO_448 (O_448,N_14107,N_14987);
xor UO_449 (O_449,N_14838,N_13990);
and UO_450 (O_450,N_14330,N_14487);
and UO_451 (O_451,N_13739,N_13585);
and UO_452 (O_452,N_14962,N_14599);
nand UO_453 (O_453,N_14697,N_14005);
nand UO_454 (O_454,N_14862,N_14526);
or UO_455 (O_455,N_13664,N_14057);
nor UO_456 (O_456,N_14064,N_14300);
nor UO_457 (O_457,N_14376,N_14096);
or UO_458 (O_458,N_14715,N_13505);
xnor UO_459 (O_459,N_14543,N_13678);
and UO_460 (O_460,N_14855,N_13861);
and UO_461 (O_461,N_13901,N_14890);
and UO_462 (O_462,N_14808,N_14480);
and UO_463 (O_463,N_13862,N_13544);
nand UO_464 (O_464,N_14713,N_14824);
or UO_465 (O_465,N_14977,N_14460);
or UO_466 (O_466,N_13615,N_14141);
nand UO_467 (O_467,N_14369,N_13923);
nor UO_468 (O_468,N_13898,N_14691);
nand UO_469 (O_469,N_14968,N_14130);
and UO_470 (O_470,N_14415,N_14775);
or UO_471 (O_471,N_14844,N_13996);
and UO_472 (O_472,N_13718,N_14737);
or UO_473 (O_473,N_14826,N_13683);
and UO_474 (O_474,N_13982,N_14416);
xor UO_475 (O_475,N_14450,N_13751);
or UO_476 (O_476,N_13714,N_13513);
nor UO_477 (O_477,N_14806,N_14481);
and UO_478 (O_478,N_14711,N_14132);
or UO_479 (O_479,N_13725,N_13902);
nor UO_480 (O_480,N_14235,N_13784);
xor UO_481 (O_481,N_14477,N_14933);
xor UO_482 (O_482,N_14572,N_14722);
or UO_483 (O_483,N_14642,N_14951);
and UO_484 (O_484,N_14281,N_13933);
and UO_485 (O_485,N_14037,N_13695);
nand UO_486 (O_486,N_14652,N_14164);
xnor UO_487 (O_487,N_13907,N_14193);
nand UO_488 (O_488,N_13677,N_14161);
and UO_489 (O_489,N_14431,N_14479);
and UO_490 (O_490,N_14185,N_14094);
nor UO_491 (O_491,N_14229,N_14180);
or UO_492 (O_492,N_14198,N_13856);
and UO_493 (O_493,N_14632,N_13998);
nand UO_494 (O_494,N_13661,N_14337);
nor UO_495 (O_495,N_14050,N_14823);
and UO_496 (O_496,N_13643,N_14701);
nor UO_497 (O_497,N_13993,N_14644);
nand UO_498 (O_498,N_14591,N_14386);
or UO_499 (O_499,N_13694,N_14340);
and UO_500 (O_500,N_13828,N_14625);
nand UO_501 (O_501,N_14886,N_13587);
nor UO_502 (O_502,N_14025,N_14519);
nor UO_503 (O_503,N_14623,N_14324);
xor UO_504 (O_504,N_14283,N_14370);
xor UO_505 (O_505,N_13932,N_14796);
or UO_506 (O_506,N_14201,N_13709);
and UO_507 (O_507,N_14788,N_14090);
or UO_508 (O_508,N_13867,N_14818);
or UO_509 (O_509,N_14169,N_14578);
nor UO_510 (O_510,N_14009,N_13696);
and UO_511 (O_511,N_13614,N_13730);
nor UO_512 (O_512,N_13888,N_14075);
nand UO_513 (O_513,N_13689,N_14421);
xor UO_514 (O_514,N_13700,N_14126);
and UO_515 (O_515,N_13595,N_14522);
and UO_516 (O_516,N_13794,N_14194);
and UO_517 (O_517,N_14210,N_14884);
nand UO_518 (O_518,N_13796,N_13759);
nor UO_519 (O_519,N_14731,N_14392);
nor UO_520 (O_520,N_13600,N_14395);
nand UO_521 (O_521,N_14864,N_14727);
or UO_522 (O_522,N_14947,N_14533);
or UO_523 (O_523,N_14113,N_14349);
or UO_524 (O_524,N_14052,N_14071);
or UO_525 (O_525,N_14849,N_14128);
nor UO_526 (O_526,N_14547,N_14101);
or UO_527 (O_527,N_13951,N_14441);
or UO_528 (O_528,N_14203,N_13701);
and UO_529 (O_529,N_14278,N_14399);
xor UO_530 (O_530,N_13580,N_14589);
nand UO_531 (O_531,N_13726,N_13669);
xnor UO_532 (O_532,N_13558,N_14072);
xor UO_533 (O_533,N_14614,N_14853);
and UO_534 (O_534,N_14741,N_14065);
or UO_535 (O_535,N_14960,N_14746);
nand UO_536 (O_536,N_13733,N_13944);
nor UO_537 (O_537,N_13728,N_14208);
or UO_538 (O_538,N_14244,N_14462);
nor UO_539 (O_539,N_14428,N_13533);
or UO_540 (O_540,N_13637,N_14121);
nor UO_541 (O_541,N_13909,N_14636);
or UO_542 (O_542,N_13961,N_14122);
nor UO_543 (O_543,N_14080,N_14134);
xnor UO_544 (O_544,N_14772,N_14695);
nor UO_545 (O_545,N_14732,N_14245);
xor UO_546 (O_546,N_13536,N_13838);
or UO_547 (O_547,N_14279,N_14104);
and UO_548 (O_548,N_14661,N_14867);
nor UO_549 (O_549,N_14140,N_13903);
or UO_550 (O_550,N_13987,N_14604);
xor UO_551 (O_551,N_14639,N_13681);
and UO_552 (O_552,N_14650,N_13917);
xnor UO_553 (O_553,N_13546,N_14432);
nand UO_554 (O_554,N_13582,N_13958);
nor UO_555 (O_555,N_14007,N_14362);
xnor UO_556 (O_556,N_13742,N_13840);
nor UO_557 (O_557,N_14765,N_13756);
nand UO_558 (O_558,N_14048,N_13773);
and UO_559 (O_559,N_14922,N_14228);
nand UO_560 (O_560,N_14761,N_13885);
xnor UO_561 (O_561,N_13698,N_14592);
nor UO_562 (O_562,N_14524,N_14514);
and UO_563 (O_563,N_14881,N_14587);
and UO_564 (O_564,N_14967,N_13981);
or UO_565 (O_565,N_14832,N_13778);
nor UO_566 (O_566,N_13723,N_14139);
nor UO_567 (O_567,N_14459,N_13911);
nor UO_568 (O_568,N_13772,N_13732);
and UO_569 (O_569,N_14325,N_14767);
and UO_570 (O_570,N_13520,N_14505);
and UO_571 (O_571,N_13916,N_13602);
nand UO_572 (O_572,N_14776,N_14347);
and UO_573 (O_573,N_13667,N_14515);
xor UO_574 (O_574,N_14341,N_14248);
xnor UO_575 (O_575,N_13727,N_13906);
xor UO_576 (O_576,N_13597,N_14840);
nor UO_577 (O_577,N_14299,N_14917);
nand UO_578 (O_578,N_14755,N_13665);
nand UO_579 (O_579,N_14963,N_13744);
and UO_580 (O_580,N_14285,N_14606);
nor UO_581 (O_581,N_14030,N_14234);
and UO_582 (O_582,N_13941,N_14027);
nand UO_583 (O_583,N_13960,N_14011);
xor UO_584 (O_584,N_14709,N_13803);
nor UO_585 (O_585,N_14133,N_14188);
and UO_586 (O_586,N_14837,N_13530);
or UO_587 (O_587,N_13915,N_14079);
nor UO_588 (O_588,N_14335,N_13697);
xnor UO_589 (O_589,N_14157,N_14719);
or UO_590 (O_590,N_14008,N_14159);
or UO_591 (O_591,N_13936,N_14986);
and UO_592 (O_592,N_14869,N_14635);
nand UO_593 (O_593,N_13868,N_14944);
nand UO_594 (O_594,N_13783,N_14726);
nand UO_595 (O_595,N_13684,N_14339);
and UO_596 (O_596,N_14084,N_13884);
nor UO_597 (O_597,N_14945,N_13565);
nand UO_598 (O_598,N_13594,N_14267);
or UO_599 (O_599,N_14924,N_13956);
or UO_600 (O_600,N_14581,N_13542);
or UO_601 (O_601,N_14819,N_14216);
and UO_602 (O_602,N_14621,N_13750);
nand UO_603 (O_603,N_14665,N_14984);
and UO_604 (O_604,N_13738,N_14910);
nand UO_605 (O_605,N_14461,N_14326);
xor UO_606 (O_606,N_13720,N_14061);
nand UO_607 (O_607,N_14168,N_14466);
and UO_608 (O_608,N_14114,N_14368);
and UO_609 (O_609,N_14257,N_13829);
nor UO_610 (O_610,N_14905,N_13871);
or UO_611 (O_611,N_13767,N_13812);
nor UO_612 (O_612,N_14029,N_14971);
and UO_613 (O_613,N_14930,N_14952);
nand UO_614 (O_614,N_14571,N_14047);
or UO_615 (O_615,N_13786,N_14352);
nand UO_616 (O_616,N_13598,N_14559);
nor UO_617 (O_617,N_13919,N_14577);
or UO_618 (O_618,N_14490,N_13712);
nand UO_619 (O_619,N_13886,N_14797);
or UO_620 (O_620,N_13636,N_14060);
nor UO_621 (O_621,N_13985,N_13873);
nand UO_622 (O_622,N_13577,N_14148);
nand UO_623 (O_623,N_14402,N_14004);
xnor UO_624 (O_624,N_13592,N_14404);
and UO_625 (O_625,N_14747,N_14222);
and UO_626 (O_626,N_14383,N_14264);
and UO_627 (O_627,N_14677,N_13779);
nand UO_628 (O_628,N_14280,N_13632);
or UO_629 (O_629,N_13581,N_14353);
nand UO_630 (O_630,N_13966,N_14499);
nand UO_631 (O_631,N_14348,N_14099);
nor UO_632 (O_632,N_14659,N_14809);
nand UO_633 (O_633,N_13954,N_14874);
or UO_634 (O_634,N_14916,N_13766);
xnor UO_635 (O_635,N_14728,N_13810);
nor UO_636 (O_636,N_14249,N_14086);
or UO_637 (O_637,N_14502,N_14531);
and UO_638 (O_638,N_13837,N_13639);
or UO_639 (O_639,N_14398,N_14539);
and UO_640 (O_640,N_14568,N_14044);
and UO_641 (O_641,N_13957,N_13556);
nor UO_642 (O_642,N_14241,N_14165);
xnor UO_643 (O_643,N_14102,N_13817);
nor UO_644 (O_644,N_13516,N_14146);
nand UO_645 (O_645,N_14158,N_13842);
xor UO_646 (O_646,N_14925,N_13955);
xor UO_647 (O_647,N_14799,N_14773);
nor UO_648 (O_648,N_14814,N_14900);
xor UO_649 (O_649,N_14856,N_14673);
nand UO_650 (O_650,N_13924,N_14022);
or UO_651 (O_651,N_14275,N_13512);
nand UO_652 (O_652,N_14704,N_14038);
nor UO_653 (O_653,N_14687,N_14290);
or UO_654 (O_654,N_14946,N_13986);
xnor UO_655 (O_655,N_14284,N_13797);
nor UO_656 (O_656,N_13777,N_13663);
nor UO_657 (O_657,N_14388,N_14006);
xnor UO_658 (O_658,N_14200,N_14835);
and UO_659 (O_659,N_14710,N_14751);
nand UO_660 (O_660,N_14895,N_14976);
or UO_661 (O_661,N_14452,N_14469);
and UO_662 (O_662,N_14667,N_13711);
xnor UO_663 (O_663,N_14273,N_13710);
or UO_664 (O_664,N_14811,N_14467);
xnor UO_665 (O_665,N_14878,N_14613);
nand UO_666 (O_666,N_14675,N_14602);
nand UO_667 (O_667,N_13515,N_13680);
nor UO_668 (O_668,N_13973,N_14730);
or UO_669 (O_669,N_14520,N_13620);
nor UO_670 (O_670,N_13566,N_13997);
xnor UO_671 (O_671,N_13752,N_13976);
or UO_672 (O_672,N_14127,N_14385);
nand UO_673 (O_673,N_13608,N_13748);
nand UO_674 (O_674,N_13908,N_14643);
nand UO_675 (O_675,N_14815,N_13848);
nor UO_676 (O_676,N_14504,N_14001);
and UO_677 (O_677,N_13721,N_13872);
nor UO_678 (O_678,N_13525,N_14839);
nand UO_679 (O_679,N_14474,N_14666);
nor UO_680 (O_680,N_13765,N_13815);
and UO_681 (O_681,N_14172,N_14176);
nand UO_682 (O_682,N_14403,N_13655);
nor UO_683 (O_683,N_14366,N_13853);
xor UO_684 (O_684,N_14003,N_14861);
or UO_685 (O_685,N_14316,N_14488);
and UO_686 (O_686,N_14914,N_14098);
nor UO_687 (O_687,N_14192,N_14854);
or UO_688 (O_688,N_14739,N_14744);
xnor UO_689 (O_689,N_13761,N_14989);
and UO_690 (O_690,N_14939,N_13874);
nand UO_691 (O_691,N_14024,N_14156);
xor UO_692 (O_692,N_13593,N_14964);
and UO_693 (O_693,N_14920,N_13863);
nand UO_694 (O_694,N_14217,N_13926);
xor UO_695 (O_695,N_14289,N_14877);
or UO_696 (O_696,N_14396,N_14277);
and UO_697 (O_697,N_14781,N_14802);
and UO_698 (O_698,N_13913,N_14453);
nor UO_699 (O_699,N_14598,N_14893);
and UO_700 (O_700,N_14770,N_13583);
xor UO_701 (O_701,N_13735,N_13532);
xnor UO_702 (O_702,N_14147,N_13647);
nand UO_703 (O_703,N_14087,N_13589);
or UO_704 (O_704,N_13575,N_13719);
nand UO_705 (O_705,N_13891,N_13900);
xor UO_706 (O_706,N_14885,N_14756);
and UO_707 (O_707,N_13804,N_13559);
nor UO_708 (O_708,N_13645,N_14601);
and UO_709 (O_709,N_14995,N_14034);
and UO_710 (O_710,N_14183,N_13670);
and UO_711 (O_711,N_14054,N_13859);
xor UO_712 (O_712,N_14334,N_13831);
and UO_713 (O_713,N_14379,N_14483);
nand UO_714 (O_714,N_13974,N_14475);
xor UO_715 (O_715,N_13975,N_14698);
xnor UO_716 (O_716,N_14410,N_14609);
xnor UO_717 (O_717,N_14590,N_13517);
xnor UO_718 (O_718,N_14748,N_14321);
nand UO_719 (O_719,N_14294,N_14444);
or UO_720 (O_720,N_14405,N_14999);
nor UO_721 (O_721,N_13858,N_14310);
nand UO_722 (O_722,N_14512,N_13534);
and UO_723 (O_723,N_14803,N_14769);
nand UO_724 (O_724,N_13904,N_13506);
and UO_725 (O_725,N_13835,N_14560);
nor UO_726 (O_726,N_14365,N_14350);
or UO_727 (O_727,N_14226,N_13818);
nand UO_728 (O_728,N_13705,N_14068);
nor UO_729 (O_729,N_13841,N_13983);
nand UO_730 (O_730,N_14820,N_14926);
nand UO_731 (O_731,N_14015,N_14866);
nor UO_732 (O_732,N_14195,N_14600);
xor UO_733 (O_733,N_14489,N_13776);
and UO_734 (O_734,N_14657,N_14843);
or UO_735 (O_735,N_14990,N_14320);
nor UO_736 (O_736,N_14911,N_14436);
xnor UO_737 (O_737,N_14658,N_14089);
nand UO_738 (O_738,N_13510,N_14640);
nand UO_739 (O_739,N_14750,N_14562);
nor UO_740 (O_740,N_14998,N_14252);
nand UO_741 (O_741,N_14066,N_14051);
or UO_742 (O_742,N_13937,N_14894);
nor UO_743 (O_743,N_14777,N_14785);
nand UO_744 (O_744,N_14225,N_14342);
and UO_745 (O_745,N_13640,N_14162);
nand UO_746 (O_746,N_14523,N_13588);
nor UO_747 (O_747,N_14538,N_13952);
xor UO_748 (O_748,N_14817,N_13578);
and UO_749 (O_749,N_14214,N_14532);
and UO_750 (O_750,N_14218,N_14419);
nand UO_751 (O_751,N_14650,N_14460);
nor UO_752 (O_752,N_14555,N_13597);
nor UO_753 (O_753,N_14909,N_13504);
or UO_754 (O_754,N_14571,N_14391);
or UO_755 (O_755,N_14761,N_13688);
nor UO_756 (O_756,N_13800,N_14439);
nor UO_757 (O_757,N_13716,N_14811);
or UO_758 (O_758,N_14230,N_14100);
or UO_759 (O_759,N_14067,N_14223);
nand UO_760 (O_760,N_14776,N_13833);
or UO_761 (O_761,N_14774,N_14135);
nor UO_762 (O_762,N_14960,N_14157);
and UO_763 (O_763,N_13753,N_14891);
or UO_764 (O_764,N_13716,N_14306);
xor UO_765 (O_765,N_14690,N_14314);
xnor UO_766 (O_766,N_14437,N_14164);
nand UO_767 (O_767,N_14984,N_13926);
and UO_768 (O_768,N_13980,N_14904);
and UO_769 (O_769,N_13902,N_13537);
and UO_770 (O_770,N_14521,N_14060);
nand UO_771 (O_771,N_14023,N_14865);
and UO_772 (O_772,N_14658,N_14499);
xor UO_773 (O_773,N_14459,N_13675);
nor UO_774 (O_774,N_14254,N_14051);
nand UO_775 (O_775,N_14184,N_14573);
and UO_776 (O_776,N_13826,N_13907);
and UO_777 (O_777,N_14169,N_14106);
nand UO_778 (O_778,N_14741,N_13848);
nand UO_779 (O_779,N_14419,N_14326);
or UO_780 (O_780,N_14427,N_14231);
nor UO_781 (O_781,N_13700,N_14038);
nor UO_782 (O_782,N_13676,N_14953);
or UO_783 (O_783,N_13605,N_14375);
nor UO_784 (O_784,N_14369,N_13861);
xnor UO_785 (O_785,N_13916,N_13936);
nand UO_786 (O_786,N_14280,N_13615);
nand UO_787 (O_787,N_13978,N_14616);
and UO_788 (O_788,N_14367,N_13915);
nand UO_789 (O_789,N_14097,N_14587);
or UO_790 (O_790,N_14227,N_13669);
nand UO_791 (O_791,N_14311,N_14606);
nand UO_792 (O_792,N_13870,N_14231);
or UO_793 (O_793,N_14205,N_14253);
xnor UO_794 (O_794,N_14312,N_14613);
nand UO_795 (O_795,N_14468,N_13894);
xor UO_796 (O_796,N_13875,N_14563);
and UO_797 (O_797,N_14614,N_14434);
nand UO_798 (O_798,N_14687,N_14881);
and UO_799 (O_799,N_14576,N_13782);
and UO_800 (O_800,N_14597,N_13869);
nor UO_801 (O_801,N_14538,N_13772);
nand UO_802 (O_802,N_14610,N_14519);
or UO_803 (O_803,N_14734,N_14311);
and UO_804 (O_804,N_13765,N_14671);
or UO_805 (O_805,N_14008,N_13794);
nor UO_806 (O_806,N_14369,N_14986);
nor UO_807 (O_807,N_14461,N_14354);
and UO_808 (O_808,N_14020,N_13553);
or UO_809 (O_809,N_14872,N_14659);
nor UO_810 (O_810,N_14759,N_14883);
and UO_811 (O_811,N_14415,N_14778);
xor UO_812 (O_812,N_14068,N_14197);
nor UO_813 (O_813,N_13746,N_14925);
and UO_814 (O_814,N_14624,N_13597);
nor UO_815 (O_815,N_13728,N_14141);
or UO_816 (O_816,N_14347,N_14411);
or UO_817 (O_817,N_14540,N_13902);
nand UO_818 (O_818,N_14873,N_14202);
and UO_819 (O_819,N_14604,N_14533);
xnor UO_820 (O_820,N_14135,N_13593);
or UO_821 (O_821,N_13602,N_14851);
nor UO_822 (O_822,N_14894,N_14270);
and UO_823 (O_823,N_14629,N_14803);
and UO_824 (O_824,N_14506,N_14603);
xor UO_825 (O_825,N_14296,N_14038);
and UO_826 (O_826,N_13819,N_14386);
nand UO_827 (O_827,N_14802,N_14965);
and UO_828 (O_828,N_14218,N_14799);
xnor UO_829 (O_829,N_14154,N_13889);
and UO_830 (O_830,N_14020,N_14922);
and UO_831 (O_831,N_13562,N_14992);
nor UO_832 (O_832,N_14055,N_14035);
nand UO_833 (O_833,N_13600,N_13725);
nor UO_834 (O_834,N_14478,N_13997);
nor UO_835 (O_835,N_14261,N_14507);
nand UO_836 (O_836,N_14444,N_14248);
xor UO_837 (O_837,N_14605,N_13820);
nand UO_838 (O_838,N_14481,N_14501);
nor UO_839 (O_839,N_14636,N_14986);
or UO_840 (O_840,N_14806,N_13601);
xor UO_841 (O_841,N_13629,N_14180);
nand UO_842 (O_842,N_13688,N_14574);
and UO_843 (O_843,N_14234,N_13563);
nor UO_844 (O_844,N_14507,N_14898);
xnor UO_845 (O_845,N_14043,N_14075);
nor UO_846 (O_846,N_14572,N_13762);
or UO_847 (O_847,N_13663,N_14774);
and UO_848 (O_848,N_13635,N_14751);
xor UO_849 (O_849,N_14435,N_14451);
nand UO_850 (O_850,N_14213,N_13843);
nor UO_851 (O_851,N_14700,N_13849);
or UO_852 (O_852,N_14481,N_13990);
nand UO_853 (O_853,N_13507,N_14224);
and UO_854 (O_854,N_14925,N_13946);
or UO_855 (O_855,N_13545,N_14090);
xor UO_856 (O_856,N_13633,N_13710);
nor UO_857 (O_857,N_14678,N_14180);
and UO_858 (O_858,N_14268,N_14693);
nand UO_859 (O_859,N_14210,N_14873);
nor UO_860 (O_860,N_14854,N_14102);
or UO_861 (O_861,N_14017,N_13523);
xor UO_862 (O_862,N_13748,N_14972);
and UO_863 (O_863,N_14718,N_14675);
nand UO_864 (O_864,N_14767,N_13940);
nor UO_865 (O_865,N_13606,N_14607);
nor UO_866 (O_866,N_14275,N_13681);
nand UO_867 (O_867,N_14591,N_14717);
or UO_868 (O_868,N_14182,N_14532);
nor UO_869 (O_869,N_13767,N_13735);
and UO_870 (O_870,N_14265,N_13758);
and UO_871 (O_871,N_14952,N_13765);
xor UO_872 (O_872,N_13586,N_13824);
or UO_873 (O_873,N_13609,N_14159);
or UO_874 (O_874,N_14545,N_14749);
nand UO_875 (O_875,N_13670,N_14728);
and UO_876 (O_876,N_13631,N_13626);
xor UO_877 (O_877,N_14940,N_14867);
xor UO_878 (O_878,N_13771,N_13684);
or UO_879 (O_879,N_14544,N_14313);
or UO_880 (O_880,N_14361,N_14334);
or UO_881 (O_881,N_13965,N_14287);
nand UO_882 (O_882,N_14182,N_14553);
nand UO_883 (O_883,N_13580,N_13625);
and UO_884 (O_884,N_14286,N_14433);
nand UO_885 (O_885,N_14488,N_14952);
or UO_886 (O_886,N_14923,N_13693);
or UO_887 (O_887,N_14644,N_13773);
and UO_888 (O_888,N_13647,N_14804);
xnor UO_889 (O_889,N_14116,N_14871);
nand UO_890 (O_890,N_14768,N_14013);
xnor UO_891 (O_891,N_14886,N_14329);
nor UO_892 (O_892,N_14207,N_13676);
and UO_893 (O_893,N_14539,N_14112);
and UO_894 (O_894,N_14046,N_14763);
nor UO_895 (O_895,N_14149,N_14288);
nor UO_896 (O_896,N_14659,N_13638);
nor UO_897 (O_897,N_14928,N_14241);
and UO_898 (O_898,N_14309,N_13999);
xnor UO_899 (O_899,N_14037,N_14949);
and UO_900 (O_900,N_14539,N_14533);
nand UO_901 (O_901,N_13535,N_13574);
or UO_902 (O_902,N_14250,N_13733);
or UO_903 (O_903,N_14601,N_14416);
or UO_904 (O_904,N_14904,N_13554);
nor UO_905 (O_905,N_14486,N_13929);
xnor UO_906 (O_906,N_14455,N_14046);
nand UO_907 (O_907,N_13827,N_13537);
nand UO_908 (O_908,N_14434,N_13570);
nand UO_909 (O_909,N_14968,N_13523);
and UO_910 (O_910,N_14565,N_14095);
nand UO_911 (O_911,N_14954,N_14470);
nor UO_912 (O_912,N_13946,N_13698);
or UO_913 (O_913,N_14085,N_14127);
nor UO_914 (O_914,N_14123,N_13722);
nand UO_915 (O_915,N_13732,N_14159);
nand UO_916 (O_916,N_14462,N_14970);
xor UO_917 (O_917,N_14059,N_14244);
nor UO_918 (O_918,N_13731,N_14135);
xnor UO_919 (O_919,N_14960,N_13805);
and UO_920 (O_920,N_14738,N_14869);
nor UO_921 (O_921,N_14800,N_14814);
and UO_922 (O_922,N_14006,N_14142);
and UO_923 (O_923,N_13944,N_13739);
nor UO_924 (O_924,N_13864,N_13828);
nand UO_925 (O_925,N_14421,N_13579);
or UO_926 (O_926,N_14099,N_14533);
or UO_927 (O_927,N_13743,N_14753);
or UO_928 (O_928,N_14304,N_14793);
xnor UO_929 (O_929,N_14544,N_14524);
or UO_930 (O_930,N_14463,N_13561);
nand UO_931 (O_931,N_14960,N_14726);
and UO_932 (O_932,N_13875,N_13947);
nor UO_933 (O_933,N_14554,N_13513);
xor UO_934 (O_934,N_14492,N_13950);
or UO_935 (O_935,N_14359,N_14446);
nand UO_936 (O_936,N_14191,N_14831);
and UO_937 (O_937,N_14819,N_14626);
and UO_938 (O_938,N_14257,N_14989);
or UO_939 (O_939,N_14974,N_14195);
and UO_940 (O_940,N_13903,N_13964);
nand UO_941 (O_941,N_13799,N_14652);
nor UO_942 (O_942,N_13648,N_14808);
or UO_943 (O_943,N_14448,N_13646);
xnor UO_944 (O_944,N_14578,N_14350);
nand UO_945 (O_945,N_14516,N_14278);
xnor UO_946 (O_946,N_14945,N_13622);
xnor UO_947 (O_947,N_13650,N_13948);
nor UO_948 (O_948,N_13576,N_13657);
nand UO_949 (O_949,N_13987,N_14591);
xor UO_950 (O_950,N_14062,N_14805);
nor UO_951 (O_951,N_14182,N_13583);
nor UO_952 (O_952,N_14471,N_13508);
nand UO_953 (O_953,N_14269,N_13514);
or UO_954 (O_954,N_13882,N_14683);
or UO_955 (O_955,N_14555,N_13927);
and UO_956 (O_956,N_14343,N_14197);
nand UO_957 (O_957,N_14111,N_13569);
nor UO_958 (O_958,N_14631,N_14815);
nand UO_959 (O_959,N_14817,N_14888);
nand UO_960 (O_960,N_13987,N_13759);
xor UO_961 (O_961,N_13889,N_14791);
nor UO_962 (O_962,N_14376,N_14706);
or UO_963 (O_963,N_13964,N_14821);
nand UO_964 (O_964,N_13519,N_14656);
or UO_965 (O_965,N_13670,N_14566);
xnor UO_966 (O_966,N_13943,N_13830);
xnor UO_967 (O_967,N_14529,N_14453);
nor UO_968 (O_968,N_14630,N_14216);
nand UO_969 (O_969,N_13598,N_13676);
nor UO_970 (O_970,N_14606,N_14806);
or UO_971 (O_971,N_14516,N_14927);
nor UO_972 (O_972,N_13579,N_14708);
nand UO_973 (O_973,N_13741,N_14257);
nor UO_974 (O_974,N_13541,N_14126);
and UO_975 (O_975,N_14686,N_14148);
nor UO_976 (O_976,N_14794,N_14343);
xor UO_977 (O_977,N_14581,N_14849);
nand UO_978 (O_978,N_14998,N_14867);
or UO_979 (O_979,N_13552,N_14707);
nand UO_980 (O_980,N_13612,N_13575);
xnor UO_981 (O_981,N_14284,N_14231);
nand UO_982 (O_982,N_13818,N_13883);
xor UO_983 (O_983,N_14826,N_14865);
or UO_984 (O_984,N_13940,N_14886);
xor UO_985 (O_985,N_14947,N_14106);
or UO_986 (O_986,N_14503,N_13761);
and UO_987 (O_987,N_14912,N_14909);
or UO_988 (O_988,N_14872,N_14952);
and UO_989 (O_989,N_14786,N_14563);
nor UO_990 (O_990,N_13789,N_13545);
or UO_991 (O_991,N_14076,N_14448);
xor UO_992 (O_992,N_14640,N_14843);
and UO_993 (O_993,N_14200,N_14688);
and UO_994 (O_994,N_14513,N_14479);
xor UO_995 (O_995,N_13850,N_14037);
nor UO_996 (O_996,N_14700,N_13555);
nand UO_997 (O_997,N_14515,N_13972);
xor UO_998 (O_998,N_13911,N_13667);
and UO_999 (O_999,N_14622,N_14930);
or UO_1000 (O_1000,N_14847,N_13685);
or UO_1001 (O_1001,N_13987,N_14891);
and UO_1002 (O_1002,N_14074,N_13601);
nor UO_1003 (O_1003,N_13789,N_14380);
xnor UO_1004 (O_1004,N_14587,N_14116);
and UO_1005 (O_1005,N_14443,N_14599);
nor UO_1006 (O_1006,N_13963,N_14712);
nor UO_1007 (O_1007,N_14940,N_13924);
nand UO_1008 (O_1008,N_14552,N_13977);
nand UO_1009 (O_1009,N_14541,N_14681);
nor UO_1010 (O_1010,N_13900,N_14550);
xor UO_1011 (O_1011,N_13875,N_13873);
and UO_1012 (O_1012,N_13965,N_14589);
xor UO_1013 (O_1013,N_13880,N_14547);
nor UO_1014 (O_1014,N_13879,N_14518);
xor UO_1015 (O_1015,N_14960,N_14360);
nand UO_1016 (O_1016,N_14010,N_13887);
xor UO_1017 (O_1017,N_14826,N_14599);
or UO_1018 (O_1018,N_14035,N_14319);
nor UO_1019 (O_1019,N_14820,N_13998);
nor UO_1020 (O_1020,N_13628,N_13509);
and UO_1021 (O_1021,N_13814,N_14909);
and UO_1022 (O_1022,N_13596,N_14109);
nand UO_1023 (O_1023,N_14865,N_13885);
and UO_1024 (O_1024,N_13925,N_13710);
nor UO_1025 (O_1025,N_14306,N_13834);
and UO_1026 (O_1026,N_13781,N_14119);
nand UO_1027 (O_1027,N_13768,N_14533);
and UO_1028 (O_1028,N_13720,N_14296);
nor UO_1029 (O_1029,N_14248,N_14442);
nand UO_1030 (O_1030,N_14118,N_13584);
and UO_1031 (O_1031,N_13545,N_13703);
nand UO_1032 (O_1032,N_14226,N_14127);
or UO_1033 (O_1033,N_14076,N_13844);
nand UO_1034 (O_1034,N_13988,N_14566);
nor UO_1035 (O_1035,N_14619,N_14324);
and UO_1036 (O_1036,N_13865,N_14610);
xor UO_1037 (O_1037,N_14704,N_14209);
and UO_1038 (O_1038,N_14070,N_14323);
or UO_1039 (O_1039,N_14532,N_14873);
nor UO_1040 (O_1040,N_14804,N_14671);
or UO_1041 (O_1041,N_13626,N_14399);
or UO_1042 (O_1042,N_14281,N_13730);
nor UO_1043 (O_1043,N_13587,N_13570);
or UO_1044 (O_1044,N_14931,N_14872);
nand UO_1045 (O_1045,N_14562,N_13855);
nor UO_1046 (O_1046,N_13982,N_14706);
nand UO_1047 (O_1047,N_14722,N_14340);
and UO_1048 (O_1048,N_13841,N_13753);
and UO_1049 (O_1049,N_13995,N_13541);
and UO_1050 (O_1050,N_14545,N_14070);
nand UO_1051 (O_1051,N_14997,N_13720);
xor UO_1052 (O_1052,N_14237,N_13849);
and UO_1053 (O_1053,N_14630,N_14544);
or UO_1054 (O_1054,N_13532,N_14030);
xor UO_1055 (O_1055,N_14220,N_14471);
and UO_1056 (O_1056,N_13702,N_13827);
nor UO_1057 (O_1057,N_14007,N_14433);
xnor UO_1058 (O_1058,N_14245,N_13670);
xnor UO_1059 (O_1059,N_14015,N_14532);
nor UO_1060 (O_1060,N_14968,N_14709);
xnor UO_1061 (O_1061,N_13673,N_14695);
and UO_1062 (O_1062,N_14805,N_14903);
nand UO_1063 (O_1063,N_14103,N_13748);
xnor UO_1064 (O_1064,N_13689,N_14049);
and UO_1065 (O_1065,N_14018,N_13609);
nor UO_1066 (O_1066,N_14828,N_13602);
or UO_1067 (O_1067,N_14550,N_13808);
xor UO_1068 (O_1068,N_14826,N_14499);
xnor UO_1069 (O_1069,N_13692,N_14360);
nor UO_1070 (O_1070,N_14407,N_14963);
and UO_1071 (O_1071,N_13695,N_13764);
or UO_1072 (O_1072,N_14298,N_13794);
nor UO_1073 (O_1073,N_14168,N_14308);
and UO_1074 (O_1074,N_14906,N_14740);
nor UO_1075 (O_1075,N_13601,N_13752);
nand UO_1076 (O_1076,N_14683,N_13765);
nand UO_1077 (O_1077,N_14657,N_14640);
and UO_1078 (O_1078,N_13885,N_14601);
xor UO_1079 (O_1079,N_14312,N_13528);
or UO_1080 (O_1080,N_14949,N_13535);
or UO_1081 (O_1081,N_14129,N_14491);
and UO_1082 (O_1082,N_14570,N_13767);
nor UO_1083 (O_1083,N_14691,N_13928);
xor UO_1084 (O_1084,N_14724,N_14992);
nand UO_1085 (O_1085,N_13917,N_14996);
and UO_1086 (O_1086,N_14627,N_14941);
xor UO_1087 (O_1087,N_14136,N_14743);
and UO_1088 (O_1088,N_14854,N_14144);
and UO_1089 (O_1089,N_14495,N_13850);
xnor UO_1090 (O_1090,N_14264,N_14913);
or UO_1091 (O_1091,N_14726,N_13653);
and UO_1092 (O_1092,N_14633,N_14628);
xor UO_1093 (O_1093,N_13745,N_14564);
or UO_1094 (O_1094,N_14955,N_14194);
xor UO_1095 (O_1095,N_14837,N_13756);
or UO_1096 (O_1096,N_13531,N_13671);
xor UO_1097 (O_1097,N_14275,N_14851);
and UO_1098 (O_1098,N_13748,N_14911);
and UO_1099 (O_1099,N_14430,N_14435);
or UO_1100 (O_1100,N_14656,N_13867);
xor UO_1101 (O_1101,N_14710,N_14103);
xnor UO_1102 (O_1102,N_14947,N_13619);
nand UO_1103 (O_1103,N_14504,N_14604);
or UO_1104 (O_1104,N_13671,N_13625);
and UO_1105 (O_1105,N_13655,N_13931);
and UO_1106 (O_1106,N_14665,N_14602);
and UO_1107 (O_1107,N_14114,N_13543);
nand UO_1108 (O_1108,N_13714,N_14700);
and UO_1109 (O_1109,N_14792,N_13973);
or UO_1110 (O_1110,N_13718,N_14459);
nand UO_1111 (O_1111,N_13629,N_14749);
nand UO_1112 (O_1112,N_13757,N_14596);
xnor UO_1113 (O_1113,N_14608,N_13759);
nor UO_1114 (O_1114,N_13847,N_14130);
xor UO_1115 (O_1115,N_14368,N_13760);
nor UO_1116 (O_1116,N_14234,N_13882);
nand UO_1117 (O_1117,N_14913,N_13543);
nor UO_1118 (O_1118,N_13754,N_14191);
xnor UO_1119 (O_1119,N_13977,N_13684);
nor UO_1120 (O_1120,N_13857,N_14187);
nand UO_1121 (O_1121,N_14923,N_14733);
xor UO_1122 (O_1122,N_14309,N_13594);
xor UO_1123 (O_1123,N_14212,N_13712);
xnor UO_1124 (O_1124,N_13776,N_14181);
and UO_1125 (O_1125,N_14582,N_14938);
xnor UO_1126 (O_1126,N_14822,N_13622);
nor UO_1127 (O_1127,N_14693,N_14210);
nand UO_1128 (O_1128,N_13636,N_13731);
nor UO_1129 (O_1129,N_14398,N_13677);
nand UO_1130 (O_1130,N_13995,N_14048);
xor UO_1131 (O_1131,N_14345,N_14724);
or UO_1132 (O_1132,N_14464,N_14898);
nor UO_1133 (O_1133,N_14174,N_14092);
or UO_1134 (O_1134,N_13824,N_13929);
nor UO_1135 (O_1135,N_13576,N_14932);
and UO_1136 (O_1136,N_14282,N_13970);
and UO_1137 (O_1137,N_14287,N_14758);
nand UO_1138 (O_1138,N_14965,N_13660);
nor UO_1139 (O_1139,N_14315,N_14401);
nor UO_1140 (O_1140,N_14519,N_14991);
nor UO_1141 (O_1141,N_14016,N_13586);
xnor UO_1142 (O_1142,N_14866,N_14337);
and UO_1143 (O_1143,N_13808,N_14333);
and UO_1144 (O_1144,N_13622,N_14177);
or UO_1145 (O_1145,N_14899,N_14845);
nor UO_1146 (O_1146,N_13723,N_13938);
nor UO_1147 (O_1147,N_14268,N_14641);
nor UO_1148 (O_1148,N_14447,N_13775);
or UO_1149 (O_1149,N_14752,N_13537);
nor UO_1150 (O_1150,N_14906,N_14183);
nand UO_1151 (O_1151,N_14781,N_14426);
nand UO_1152 (O_1152,N_14691,N_14240);
and UO_1153 (O_1153,N_13795,N_14134);
nand UO_1154 (O_1154,N_14098,N_14924);
xor UO_1155 (O_1155,N_14582,N_14239);
nand UO_1156 (O_1156,N_13525,N_14907);
xnor UO_1157 (O_1157,N_14060,N_14780);
xor UO_1158 (O_1158,N_14315,N_13871);
or UO_1159 (O_1159,N_13984,N_14874);
or UO_1160 (O_1160,N_14210,N_14967);
nand UO_1161 (O_1161,N_14996,N_14568);
and UO_1162 (O_1162,N_14476,N_14985);
and UO_1163 (O_1163,N_14115,N_14788);
xnor UO_1164 (O_1164,N_13670,N_14609);
nor UO_1165 (O_1165,N_14844,N_13726);
nand UO_1166 (O_1166,N_13976,N_13537);
or UO_1167 (O_1167,N_13888,N_14906);
and UO_1168 (O_1168,N_14504,N_14722);
or UO_1169 (O_1169,N_14798,N_14004);
and UO_1170 (O_1170,N_13652,N_13868);
or UO_1171 (O_1171,N_14418,N_13937);
xnor UO_1172 (O_1172,N_14327,N_13661);
or UO_1173 (O_1173,N_13563,N_14085);
or UO_1174 (O_1174,N_14962,N_13596);
nor UO_1175 (O_1175,N_14881,N_14041);
or UO_1176 (O_1176,N_14337,N_14706);
nand UO_1177 (O_1177,N_14232,N_14272);
xor UO_1178 (O_1178,N_13652,N_14783);
xnor UO_1179 (O_1179,N_13548,N_13991);
xor UO_1180 (O_1180,N_14690,N_14402);
nor UO_1181 (O_1181,N_13728,N_14535);
xor UO_1182 (O_1182,N_13791,N_13578);
xor UO_1183 (O_1183,N_14602,N_13622);
nand UO_1184 (O_1184,N_13768,N_13942);
nor UO_1185 (O_1185,N_14681,N_14678);
nand UO_1186 (O_1186,N_13906,N_13720);
nor UO_1187 (O_1187,N_14742,N_13888);
nor UO_1188 (O_1188,N_14062,N_14423);
nand UO_1189 (O_1189,N_14683,N_13740);
and UO_1190 (O_1190,N_13956,N_14206);
and UO_1191 (O_1191,N_13658,N_14235);
nor UO_1192 (O_1192,N_14521,N_13742);
nand UO_1193 (O_1193,N_13861,N_14348);
xnor UO_1194 (O_1194,N_14124,N_14660);
nor UO_1195 (O_1195,N_14845,N_14309);
or UO_1196 (O_1196,N_13759,N_13971);
nor UO_1197 (O_1197,N_13918,N_13891);
or UO_1198 (O_1198,N_14963,N_14989);
nor UO_1199 (O_1199,N_14851,N_14263);
nand UO_1200 (O_1200,N_14104,N_13511);
nor UO_1201 (O_1201,N_13836,N_13903);
xor UO_1202 (O_1202,N_13614,N_13959);
or UO_1203 (O_1203,N_13699,N_13752);
or UO_1204 (O_1204,N_14859,N_14175);
nand UO_1205 (O_1205,N_14454,N_13714);
or UO_1206 (O_1206,N_13507,N_14607);
nand UO_1207 (O_1207,N_14669,N_14952);
nand UO_1208 (O_1208,N_13619,N_13975);
nand UO_1209 (O_1209,N_14007,N_14948);
nor UO_1210 (O_1210,N_14390,N_14496);
xor UO_1211 (O_1211,N_14372,N_14997);
nand UO_1212 (O_1212,N_13552,N_13968);
xor UO_1213 (O_1213,N_14579,N_14053);
or UO_1214 (O_1214,N_14499,N_13536);
nor UO_1215 (O_1215,N_13576,N_13556);
nand UO_1216 (O_1216,N_13829,N_14489);
xor UO_1217 (O_1217,N_13612,N_14437);
or UO_1218 (O_1218,N_14966,N_14132);
nor UO_1219 (O_1219,N_14703,N_14373);
nor UO_1220 (O_1220,N_14335,N_14448);
and UO_1221 (O_1221,N_14192,N_14426);
and UO_1222 (O_1222,N_13830,N_14188);
or UO_1223 (O_1223,N_14988,N_14257);
nor UO_1224 (O_1224,N_13977,N_14651);
nand UO_1225 (O_1225,N_14834,N_14670);
nand UO_1226 (O_1226,N_14396,N_14742);
and UO_1227 (O_1227,N_13754,N_14617);
nor UO_1228 (O_1228,N_14389,N_14024);
xor UO_1229 (O_1229,N_14571,N_14187);
nand UO_1230 (O_1230,N_14966,N_14274);
xor UO_1231 (O_1231,N_14830,N_14361);
nor UO_1232 (O_1232,N_14776,N_14832);
nand UO_1233 (O_1233,N_14092,N_13584);
nor UO_1234 (O_1234,N_14068,N_14647);
nand UO_1235 (O_1235,N_13968,N_14824);
or UO_1236 (O_1236,N_14219,N_14188);
or UO_1237 (O_1237,N_13580,N_13948);
xnor UO_1238 (O_1238,N_13625,N_14275);
nor UO_1239 (O_1239,N_14886,N_13850);
or UO_1240 (O_1240,N_14934,N_13950);
xor UO_1241 (O_1241,N_14769,N_14859);
nor UO_1242 (O_1242,N_14904,N_14243);
and UO_1243 (O_1243,N_14649,N_14413);
and UO_1244 (O_1244,N_13785,N_13584);
nor UO_1245 (O_1245,N_14298,N_14675);
and UO_1246 (O_1246,N_13620,N_13882);
xor UO_1247 (O_1247,N_14978,N_13700);
nand UO_1248 (O_1248,N_14652,N_13830);
xor UO_1249 (O_1249,N_14553,N_14201);
nand UO_1250 (O_1250,N_14810,N_14350);
xnor UO_1251 (O_1251,N_13533,N_13781);
and UO_1252 (O_1252,N_13831,N_14854);
or UO_1253 (O_1253,N_13596,N_14394);
or UO_1254 (O_1254,N_14959,N_13588);
nand UO_1255 (O_1255,N_13765,N_14385);
nor UO_1256 (O_1256,N_13826,N_14184);
and UO_1257 (O_1257,N_13541,N_14443);
nand UO_1258 (O_1258,N_14395,N_14876);
or UO_1259 (O_1259,N_14873,N_14975);
nand UO_1260 (O_1260,N_14709,N_14679);
and UO_1261 (O_1261,N_14491,N_13860);
or UO_1262 (O_1262,N_14198,N_14832);
and UO_1263 (O_1263,N_14071,N_14446);
and UO_1264 (O_1264,N_13655,N_14317);
nor UO_1265 (O_1265,N_14993,N_13508);
nor UO_1266 (O_1266,N_14366,N_14155);
nand UO_1267 (O_1267,N_14623,N_13971);
xnor UO_1268 (O_1268,N_13529,N_13932);
and UO_1269 (O_1269,N_14657,N_13502);
or UO_1270 (O_1270,N_13530,N_14835);
or UO_1271 (O_1271,N_13537,N_13505);
nand UO_1272 (O_1272,N_14692,N_14067);
and UO_1273 (O_1273,N_13913,N_14597);
nand UO_1274 (O_1274,N_13919,N_14455);
xor UO_1275 (O_1275,N_14983,N_13668);
and UO_1276 (O_1276,N_13560,N_14435);
or UO_1277 (O_1277,N_14056,N_14981);
xnor UO_1278 (O_1278,N_13715,N_14421);
nand UO_1279 (O_1279,N_13607,N_14886);
or UO_1280 (O_1280,N_14470,N_14510);
or UO_1281 (O_1281,N_14649,N_14037);
nand UO_1282 (O_1282,N_14088,N_13929);
nand UO_1283 (O_1283,N_14612,N_14103);
xnor UO_1284 (O_1284,N_14065,N_14640);
xnor UO_1285 (O_1285,N_14054,N_14202);
and UO_1286 (O_1286,N_14979,N_14236);
xor UO_1287 (O_1287,N_14110,N_13689);
nand UO_1288 (O_1288,N_13878,N_13631);
xor UO_1289 (O_1289,N_13617,N_14550);
or UO_1290 (O_1290,N_13815,N_13776);
and UO_1291 (O_1291,N_13936,N_14037);
and UO_1292 (O_1292,N_14212,N_13950);
and UO_1293 (O_1293,N_14241,N_14081);
nand UO_1294 (O_1294,N_13588,N_13967);
xnor UO_1295 (O_1295,N_13734,N_13772);
nand UO_1296 (O_1296,N_14260,N_14288);
and UO_1297 (O_1297,N_13503,N_14505);
nand UO_1298 (O_1298,N_14757,N_14306);
xnor UO_1299 (O_1299,N_14738,N_14857);
xnor UO_1300 (O_1300,N_13889,N_13540);
xor UO_1301 (O_1301,N_14116,N_13923);
nand UO_1302 (O_1302,N_14171,N_14555);
nor UO_1303 (O_1303,N_14029,N_14445);
or UO_1304 (O_1304,N_14134,N_14217);
and UO_1305 (O_1305,N_13817,N_14346);
xnor UO_1306 (O_1306,N_14930,N_14774);
nor UO_1307 (O_1307,N_14151,N_14242);
nor UO_1308 (O_1308,N_13741,N_13555);
xnor UO_1309 (O_1309,N_13574,N_13993);
xor UO_1310 (O_1310,N_13926,N_13857);
xnor UO_1311 (O_1311,N_14937,N_14689);
xnor UO_1312 (O_1312,N_14933,N_14188);
and UO_1313 (O_1313,N_14861,N_14167);
nand UO_1314 (O_1314,N_14349,N_13785);
or UO_1315 (O_1315,N_14412,N_14271);
xor UO_1316 (O_1316,N_13757,N_14742);
nor UO_1317 (O_1317,N_13827,N_14296);
nand UO_1318 (O_1318,N_14564,N_13979);
or UO_1319 (O_1319,N_14193,N_13670);
or UO_1320 (O_1320,N_14515,N_14562);
and UO_1321 (O_1321,N_14714,N_14331);
nor UO_1322 (O_1322,N_14744,N_14697);
nor UO_1323 (O_1323,N_13781,N_13760);
and UO_1324 (O_1324,N_14497,N_14727);
and UO_1325 (O_1325,N_14009,N_14631);
and UO_1326 (O_1326,N_14679,N_13642);
or UO_1327 (O_1327,N_14141,N_14166);
or UO_1328 (O_1328,N_14423,N_13986);
xnor UO_1329 (O_1329,N_13966,N_13522);
nor UO_1330 (O_1330,N_14680,N_14532);
xor UO_1331 (O_1331,N_13537,N_14856);
nand UO_1332 (O_1332,N_13643,N_14491);
nand UO_1333 (O_1333,N_14871,N_14002);
nand UO_1334 (O_1334,N_14513,N_14046);
and UO_1335 (O_1335,N_14716,N_14447);
xnor UO_1336 (O_1336,N_14327,N_14259);
nor UO_1337 (O_1337,N_13859,N_14430);
nor UO_1338 (O_1338,N_13759,N_14814);
and UO_1339 (O_1339,N_14780,N_14462);
xor UO_1340 (O_1340,N_14392,N_14979);
and UO_1341 (O_1341,N_14331,N_14098);
nand UO_1342 (O_1342,N_14071,N_14570);
nor UO_1343 (O_1343,N_13713,N_14943);
nor UO_1344 (O_1344,N_14603,N_13586);
xor UO_1345 (O_1345,N_14254,N_13885);
xnor UO_1346 (O_1346,N_14583,N_14874);
or UO_1347 (O_1347,N_14573,N_14366);
xor UO_1348 (O_1348,N_13533,N_14078);
xor UO_1349 (O_1349,N_14284,N_13889);
or UO_1350 (O_1350,N_13632,N_14757);
and UO_1351 (O_1351,N_14337,N_14804);
and UO_1352 (O_1352,N_14699,N_13805);
xor UO_1353 (O_1353,N_14696,N_14142);
and UO_1354 (O_1354,N_14416,N_14683);
xor UO_1355 (O_1355,N_13923,N_14821);
nor UO_1356 (O_1356,N_13510,N_14589);
nor UO_1357 (O_1357,N_14612,N_13595);
and UO_1358 (O_1358,N_14092,N_14673);
nor UO_1359 (O_1359,N_13813,N_14219);
or UO_1360 (O_1360,N_14861,N_14942);
nand UO_1361 (O_1361,N_14276,N_14729);
nand UO_1362 (O_1362,N_14973,N_14592);
and UO_1363 (O_1363,N_13509,N_13681);
nor UO_1364 (O_1364,N_14854,N_14496);
or UO_1365 (O_1365,N_14958,N_13705);
nor UO_1366 (O_1366,N_13527,N_14697);
and UO_1367 (O_1367,N_14453,N_14897);
or UO_1368 (O_1368,N_14354,N_14626);
nand UO_1369 (O_1369,N_13827,N_14006);
xor UO_1370 (O_1370,N_13532,N_14527);
xor UO_1371 (O_1371,N_14761,N_14212);
and UO_1372 (O_1372,N_13962,N_14532);
nand UO_1373 (O_1373,N_13723,N_14933);
xnor UO_1374 (O_1374,N_13999,N_13919);
nor UO_1375 (O_1375,N_14509,N_14937);
xnor UO_1376 (O_1376,N_14288,N_14557);
xnor UO_1377 (O_1377,N_14777,N_14012);
xnor UO_1378 (O_1378,N_13528,N_14489);
nand UO_1379 (O_1379,N_13691,N_13623);
nand UO_1380 (O_1380,N_14336,N_14880);
xnor UO_1381 (O_1381,N_14648,N_13785);
xnor UO_1382 (O_1382,N_14029,N_14672);
xor UO_1383 (O_1383,N_13801,N_14136);
nand UO_1384 (O_1384,N_14174,N_14712);
or UO_1385 (O_1385,N_14215,N_14084);
nor UO_1386 (O_1386,N_14762,N_14802);
and UO_1387 (O_1387,N_13986,N_14176);
and UO_1388 (O_1388,N_14193,N_14823);
or UO_1389 (O_1389,N_13815,N_14020);
and UO_1390 (O_1390,N_14781,N_14562);
nor UO_1391 (O_1391,N_13652,N_13844);
and UO_1392 (O_1392,N_14022,N_14479);
nor UO_1393 (O_1393,N_14063,N_14024);
nor UO_1394 (O_1394,N_13791,N_14710);
nor UO_1395 (O_1395,N_13757,N_14969);
nor UO_1396 (O_1396,N_13695,N_14317);
nand UO_1397 (O_1397,N_14769,N_14710);
or UO_1398 (O_1398,N_14387,N_14264);
nor UO_1399 (O_1399,N_13945,N_14078);
nor UO_1400 (O_1400,N_13816,N_14841);
and UO_1401 (O_1401,N_14958,N_13739);
nor UO_1402 (O_1402,N_14339,N_14544);
or UO_1403 (O_1403,N_13944,N_14545);
nand UO_1404 (O_1404,N_14185,N_13574);
xnor UO_1405 (O_1405,N_14435,N_13957);
nor UO_1406 (O_1406,N_14784,N_14922);
nor UO_1407 (O_1407,N_13568,N_14765);
nor UO_1408 (O_1408,N_14841,N_13583);
or UO_1409 (O_1409,N_14660,N_14129);
or UO_1410 (O_1410,N_13599,N_14992);
or UO_1411 (O_1411,N_14067,N_13849);
or UO_1412 (O_1412,N_14699,N_13889);
xor UO_1413 (O_1413,N_14993,N_14569);
nor UO_1414 (O_1414,N_13718,N_14498);
or UO_1415 (O_1415,N_14785,N_13650);
and UO_1416 (O_1416,N_14482,N_14585);
xor UO_1417 (O_1417,N_13859,N_14166);
nand UO_1418 (O_1418,N_14873,N_14213);
or UO_1419 (O_1419,N_14807,N_14469);
nor UO_1420 (O_1420,N_14381,N_14081);
nand UO_1421 (O_1421,N_13535,N_14107);
and UO_1422 (O_1422,N_13652,N_13978);
nand UO_1423 (O_1423,N_13935,N_13740);
xnor UO_1424 (O_1424,N_14686,N_14062);
or UO_1425 (O_1425,N_14087,N_14157);
or UO_1426 (O_1426,N_14023,N_13671);
or UO_1427 (O_1427,N_14396,N_14205);
xor UO_1428 (O_1428,N_14019,N_13687);
and UO_1429 (O_1429,N_13867,N_14201);
nor UO_1430 (O_1430,N_13714,N_14041);
and UO_1431 (O_1431,N_14621,N_14641);
nor UO_1432 (O_1432,N_13600,N_13733);
or UO_1433 (O_1433,N_13619,N_14033);
and UO_1434 (O_1434,N_14570,N_14044);
xnor UO_1435 (O_1435,N_14709,N_14068);
nor UO_1436 (O_1436,N_14876,N_14940);
or UO_1437 (O_1437,N_14111,N_14562);
xnor UO_1438 (O_1438,N_14128,N_14990);
nand UO_1439 (O_1439,N_14353,N_13547);
nand UO_1440 (O_1440,N_14862,N_14375);
nand UO_1441 (O_1441,N_13618,N_13725);
or UO_1442 (O_1442,N_14800,N_14283);
nor UO_1443 (O_1443,N_13966,N_13509);
nand UO_1444 (O_1444,N_14629,N_14502);
and UO_1445 (O_1445,N_13894,N_14201);
and UO_1446 (O_1446,N_13705,N_14984);
or UO_1447 (O_1447,N_14279,N_14573);
xor UO_1448 (O_1448,N_14133,N_13642);
and UO_1449 (O_1449,N_14224,N_14433);
or UO_1450 (O_1450,N_13951,N_14561);
and UO_1451 (O_1451,N_14658,N_13570);
nor UO_1452 (O_1452,N_14288,N_14327);
nand UO_1453 (O_1453,N_14844,N_14490);
xnor UO_1454 (O_1454,N_14865,N_13612);
nand UO_1455 (O_1455,N_14379,N_13561);
nand UO_1456 (O_1456,N_14694,N_13788);
nand UO_1457 (O_1457,N_14391,N_14828);
and UO_1458 (O_1458,N_14380,N_14584);
or UO_1459 (O_1459,N_14674,N_14934);
nand UO_1460 (O_1460,N_13727,N_14637);
and UO_1461 (O_1461,N_14276,N_14230);
or UO_1462 (O_1462,N_13837,N_14640);
nor UO_1463 (O_1463,N_14524,N_14163);
nor UO_1464 (O_1464,N_14443,N_13881);
and UO_1465 (O_1465,N_13658,N_14672);
nand UO_1466 (O_1466,N_13727,N_14558);
and UO_1467 (O_1467,N_14132,N_14272);
nand UO_1468 (O_1468,N_13886,N_14235);
or UO_1469 (O_1469,N_13551,N_13839);
and UO_1470 (O_1470,N_14848,N_13969);
and UO_1471 (O_1471,N_14443,N_14863);
nor UO_1472 (O_1472,N_14699,N_13595);
nand UO_1473 (O_1473,N_14627,N_13631);
nand UO_1474 (O_1474,N_14429,N_13953);
nor UO_1475 (O_1475,N_13500,N_14627);
nor UO_1476 (O_1476,N_13846,N_14362);
xnor UO_1477 (O_1477,N_14882,N_14247);
nor UO_1478 (O_1478,N_14405,N_14138);
xor UO_1479 (O_1479,N_14532,N_14445);
nand UO_1480 (O_1480,N_13757,N_13792);
or UO_1481 (O_1481,N_13521,N_14252);
xnor UO_1482 (O_1482,N_14312,N_13865);
xnor UO_1483 (O_1483,N_13545,N_14515);
nor UO_1484 (O_1484,N_13738,N_14719);
nor UO_1485 (O_1485,N_14622,N_13869);
and UO_1486 (O_1486,N_14276,N_14115);
nor UO_1487 (O_1487,N_14139,N_14995);
nand UO_1488 (O_1488,N_14363,N_14293);
xor UO_1489 (O_1489,N_14596,N_13887);
and UO_1490 (O_1490,N_14410,N_14066);
and UO_1491 (O_1491,N_14746,N_14759);
and UO_1492 (O_1492,N_13548,N_14987);
and UO_1493 (O_1493,N_14028,N_14173);
and UO_1494 (O_1494,N_14658,N_13824);
nand UO_1495 (O_1495,N_14351,N_13804);
nor UO_1496 (O_1496,N_14240,N_14083);
and UO_1497 (O_1497,N_14843,N_14962);
nor UO_1498 (O_1498,N_14974,N_13781);
and UO_1499 (O_1499,N_14393,N_14187);
xnor UO_1500 (O_1500,N_14977,N_13768);
nand UO_1501 (O_1501,N_14170,N_13921);
nand UO_1502 (O_1502,N_14143,N_13915);
nand UO_1503 (O_1503,N_13557,N_13980);
or UO_1504 (O_1504,N_14824,N_14973);
xnor UO_1505 (O_1505,N_14998,N_13792);
nand UO_1506 (O_1506,N_13917,N_14081);
and UO_1507 (O_1507,N_14845,N_14229);
nor UO_1508 (O_1508,N_13608,N_14718);
nand UO_1509 (O_1509,N_13574,N_13907);
nor UO_1510 (O_1510,N_14297,N_14803);
and UO_1511 (O_1511,N_13902,N_14734);
and UO_1512 (O_1512,N_14595,N_13742);
nor UO_1513 (O_1513,N_14917,N_14100);
or UO_1514 (O_1514,N_14236,N_14636);
and UO_1515 (O_1515,N_14431,N_14274);
or UO_1516 (O_1516,N_14826,N_14245);
or UO_1517 (O_1517,N_14781,N_14776);
or UO_1518 (O_1518,N_14323,N_14805);
nand UO_1519 (O_1519,N_13623,N_13661);
xnor UO_1520 (O_1520,N_14320,N_14938);
and UO_1521 (O_1521,N_14266,N_14279);
or UO_1522 (O_1522,N_14806,N_13835);
xor UO_1523 (O_1523,N_13507,N_14809);
nand UO_1524 (O_1524,N_14251,N_14092);
or UO_1525 (O_1525,N_13798,N_14029);
and UO_1526 (O_1526,N_13754,N_14506);
or UO_1527 (O_1527,N_14259,N_13874);
xnor UO_1528 (O_1528,N_14955,N_14123);
nand UO_1529 (O_1529,N_14090,N_13683);
and UO_1530 (O_1530,N_13841,N_14541);
and UO_1531 (O_1531,N_14747,N_14234);
nor UO_1532 (O_1532,N_13958,N_13783);
xor UO_1533 (O_1533,N_14495,N_14892);
nand UO_1534 (O_1534,N_14365,N_14510);
and UO_1535 (O_1535,N_13873,N_13690);
xnor UO_1536 (O_1536,N_14590,N_13726);
and UO_1537 (O_1537,N_13956,N_14748);
nand UO_1538 (O_1538,N_13905,N_14768);
or UO_1539 (O_1539,N_13889,N_14285);
or UO_1540 (O_1540,N_13688,N_14426);
xor UO_1541 (O_1541,N_14979,N_13539);
or UO_1542 (O_1542,N_13609,N_13523);
and UO_1543 (O_1543,N_14997,N_14177);
and UO_1544 (O_1544,N_13684,N_13623);
and UO_1545 (O_1545,N_14495,N_14760);
and UO_1546 (O_1546,N_14805,N_13732);
nor UO_1547 (O_1547,N_13744,N_14401);
nor UO_1548 (O_1548,N_14157,N_14418);
and UO_1549 (O_1549,N_14845,N_13840);
xnor UO_1550 (O_1550,N_13742,N_13778);
and UO_1551 (O_1551,N_14456,N_13667);
or UO_1552 (O_1552,N_14955,N_14784);
or UO_1553 (O_1553,N_14114,N_14759);
xnor UO_1554 (O_1554,N_13674,N_14976);
nand UO_1555 (O_1555,N_13896,N_13511);
and UO_1556 (O_1556,N_14134,N_14484);
or UO_1557 (O_1557,N_14734,N_13815);
nand UO_1558 (O_1558,N_14002,N_14251);
or UO_1559 (O_1559,N_14991,N_14369);
nand UO_1560 (O_1560,N_14799,N_14276);
or UO_1561 (O_1561,N_13940,N_14258);
nor UO_1562 (O_1562,N_13915,N_14078);
nand UO_1563 (O_1563,N_14688,N_14642);
or UO_1564 (O_1564,N_13912,N_14855);
or UO_1565 (O_1565,N_14617,N_14933);
nand UO_1566 (O_1566,N_14941,N_14783);
or UO_1567 (O_1567,N_14469,N_13647);
nor UO_1568 (O_1568,N_14134,N_14705);
or UO_1569 (O_1569,N_14323,N_14917);
nand UO_1570 (O_1570,N_14813,N_14778);
nand UO_1571 (O_1571,N_13925,N_13996);
and UO_1572 (O_1572,N_13939,N_14807);
nor UO_1573 (O_1573,N_14929,N_14314);
or UO_1574 (O_1574,N_14074,N_14790);
nor UO_1575 (O_1575,N_14382,N_14227);
xnor UO_1576 (O_1576,N_14951,N_14489);
xor UO_1577 (O_1577,N_13840,N_14728);
or UO_1578 (O_1578,N_14504,N_14776);
or UO_1579 (O_1579,N_13626,N_14556);
nand UO_1580 (O_1580,N_14778,N_14265);
nand UO_1581 (O_1581,N_14143,N_14998);
nand UO_1582 (O_1582,N_14680,N_14473);
and UO_1583 (O_1583,N_13810,N_13538);
and UO_1584 (O_1584,N_14817,N_13813);
nand UO_1585 (O_1585,N_14169,N_14281);
xor UO_1586 (O_1586,N_14221,N_14931);
xnor UO_1587 (O_1587,N_13763,N_13725);
xnor UO_1588 (O_1588,N_14644,N_13523);
or UO_1589 (O_1589,N_14181,N_14471);
nand UO_1590 (O_1590,N_13991,N_14064);
or UO_1591 (O_1591,N_14456,N_14766);
nand UO_1592 (O_1592,N_14359,N_14681);
xnor UO_1593 (O_1593,N_13833,N_13741);
and UO_1594 (O_1594,N_14592,N_14186);
nand UO_1595 (O_1595,N_13898,N_13787);
nand UO_1596 (O_1596,N_14350,N_13784);
nand UO_1597 (O_1597,N_13976,N_14314);
nand UO_1598 (O_1598,N_13704,N_13681);
nand UO_1599 (O_1599,N_13777,N_14120);
or UO_1600 (O_1600,N_13879,N_13510);
and UO_1601 (O_1601,N_14881,N_14459);
xnor UO_1602 (O_1602,N_13701,N_13931);
nor UO_1603 (O_1603,N_13765,N_13835);
nand UO_1604 (O_1604,N_14911,N_14331);
and UO_1605 (O_1605,N_13830,N_13878);
nor UO_1606 (O_1606,N_14316,N_13829);
xor UO_1607 (O_1607,N_13827,N_14184);
or UO_1608 (O_1608,N_14326,N_14999);
nor UO_1609 (O_1609,N_14634,N_14009);
or UO_1610 (O_1610,N_14170,N_13697);
nor UO_1611 (O_1611,N_14341,N_14455);
xor UO_1612 (O_1612,N_14712,N_13542);
nand UO_1613 (O_1613,N_14768,N_14748);
or UO_1614 (O_1614,N_13512,N_14799);
and UO_1615 (O_1615,N_13669,N_13882);
or UO_1616 (O_1616,N_13921,N_14997);
or UO_1617 (O_1617,N_14035,N_14606);
or UO_1618 (O_1618,N_14672,N_14197);
xnor UO_1619 (O_1619,N_13763,N_13633);
or UO_1620 (O_1620,N_14600,N_14993);
nand UO_1621 (O_1621,N_14511,N_14707);
xnor UO_1622 (O_1622,N_14605,N_14222);
nand UO_1623 (O_1623,N_13545,N_13539);
or UO_1624 (O_1624,N_14160,N_13695);
or UO_1625 (O_1625,N_13565,N_13558);
or UO_1626 (O_1626,N_14294,N_13620);
or UO_1627 (O_1627,N_14959,N_14099);
nand UO_1628 (O_1628,N_13862,N_14767);
nor UO_1629 (O_1629,N_14355,N_14938);
and UO_1630 (O_1630,N_13864,N_14201);
nor UO_1631 (O_1631,N_13714,N_14251);
nor UO_1632 (O_1632,N_14283,N_14409);
xor UO_1633 (O_1633,N_13519,N_13933);
and UO_1634 (O_1634,N_14977,N_13621);
or UO_1635 (O_1635,N_14515,N_14049);
xnor UO_1636 (O_1636,N_14264,N_13958);
and UO_1637 (O_1637,N_14741,N_13669);
and UO_1638 (O_1638,N_13547,N_14366);
xor UO_1639 (O_1639,N_14070,N_14444);
nor UO_1640 (O_1640,N_14788,N_13887);
and UO_1641 (O_1641,N_14875,N_14471);
nor UO_1642 (O_1642,N_14856,N_14410);
and UO_1643 (O_1643,N_14176,N_14600);
xnor UO_1644 (O_1644,N_13831,N_14574);
nor UO_1645 (O_1645,N_14025,N_13886);
xor UO_1646 (O_1646,N_14656,N_14358);
or UO_1647 (O_1647,N_14837,N_14822);
and UO_1648 (O_1648,N_14509,N_14617);
or UO_1649 (O_1649,N_14027,N_14138);
xnor UO_1650 (O_1650,N_13851,N_13938);
xor UO_1651 (O_1651,N_14219,N_14921);
nand UO_1652 (O_1652,N_14084,N_13793);
and UO_1653 (O_1653,N_14040,N_13696);
xor UO_1654 (O_1654,N_14268,N_13654);
or UO_1655 (O_1655,N_14016,N_13726);
xnor UO_1656 (O_1656,N_14066,N_14949);
nor UO_1657 (O_1657,N_14603,N_13938);
and UO_1658 (O_1658,N_14113,N_13664);
nand UO_1659 (O_1659,N_14253,N_13987);
nor UO_1660 (O_1660,N_13603,N_14258);
or UO_1661 (O_1661,N_14573,N_13715);
nor UO_1662 (O_1662,N_14147,N_14152);
and UO_1663 (O_1663,N_14124,N_13759);
xor UO_1664 (O_1664,N_13807,N_14019);
and UO_1665 (O_1665,N_14039,N_14309);
nor UO_1666 (O_1666,N_14088,N_14133);
nand UO_1667 (O_1667,N_13675,N_14346);
nand UO_1668 (O_1668,N_14227,N_14886);
or UO_1669 (O_1669,N_14791,N_14379);
or UO_1670 (O_1670,N_14612,N_14781);
xor UO_1671 (O_1671,N_13610,N_14377);
nor UO_1672 (O_1672,N_14525,N_14326);
xnor UO_1673 (O_1673,N_14951,N_13515);
and UO_1674 (O_1674,N_14341,N_14683);
or UO_1675 (O_1675,N_14492,N_14915);
or UO_1676 (O_1676,N_14941,N_14427);
and UO_1677 (O_1677,N_14731,N_14140);
xnor UO_1678 (O_1678,N_13722,N_13735);
and UO_1679 (O_1679,N_14579,N_14250);
nor UO_1680 (O_1680,N_14529,N_14700);
nand UO_1681 (O_1681,N_14745,N_13965);
and UO_1682 (O_1682,N_14769,N_14806);
or UO_1683 (O_1683,N_14225,N_14297);
nand UO_1684 (O_1684,N_14530,N_14152);
nor UO_1685 (O_1685,N_13776,N_14753);
xnor UO_1686 (O_1686,N_13545,N_13585);
nand UO_1687 (O_1687,N_13680,N_14488);
and UO_1688 (O_1688,N_14773,N_13917);
xnor UO_1689 (O_1689,N_14510,N_14952);
and UO_1690 (O_1690,N_14997,N_13576);
xnor UO_1691 (O_1691,N_13895,N_13869);
xnor UO_1692 (O_1692,N_14749,N_14293);
nand UO_1693 (O_1693,N_14997,N_14260);
nor UO_1694 (O_1694,N_14515,N_14022);
nor UO_1695 (O_1695,N_14111,N_14291);
nand UO_1696 (O_1696,N_14343,N_13863);
nor UO_1697 (O_1697,N_14705,N_14901);
nand UO_1698 (O_1698,N_14597,N_13963);
xnor UO_1699 (O_1699,N_14192,N_14008);
and UO_1700 (O_1700,N_14674,N_13693);
and UO_1701 (O_1701,N_13696,N_14088);
or UO_1702 (O_1702,N_14539,N_14439);
or UO_1703 (O_1703,N_14031,N_13955);
or UO_1704 (O_1704,N_13650,N_14648);
nor UO_1705 (O_1705,N_14329,N_14850);
nor UO_1706 (O_1706,N_13905,N_14749);
nand UO_1707 (O_1707,N_13786,N_14368);
and UO_1708 (O_1708,N_14162,N_13908);
and UO_1709 (O_1709,N_14902,N_14260);
nor UO_1710 (O_1710,N_14213,N_14967);
or UO_1711 (O_1711,N_13872,N_14432);
nor UO_1712 (O_1712,N_14055,N_14169);
and UO_1713 (O_1713,N_14515,N_14363);
xor UO_1714 (O_1714,N_14342,N_14627);
or UO_1715 (O_1715,N_14654,N_13784);
and UO_1716 (O_1716,N_13655,N_13981);
and UO_1717 (O_1717,N_14577,N_13920);
nand UO_1718 (O_1718,N_14345,N_14251);
xor UO_1719 (O_1719,N_13872,N_14940);
nor UO_1720 (O_1720,N_13650,N_13649);
or UO_1721 (O_1721,N_14702,N_14041);
and UO_1722 (O_1722,N_14769,N_13900);
nor UO_1723 (O_1723,N_13646,N_14166);
xor UO_1724 (O_1724,N_14451,N_14977);
xnor UO_1725 (O_1725,N_13761,N_14263);
nand UO_1726 (O_1726,N_14926,N_14373);
nand UO_1727 (O_1727,N_13586,N_13637);
and UO_1728 (O_1728,N_14873,N_14054);
nor UO_1729 (O_1729,N_14007,N_13546);
and UO_1730 (O_1730,N_14347,N_14999);
or UO_1731 (O_1731,N_14618,N_13746);
or UO_1732 (O_1732,N_13942,N_13817);
xor UO_1733 (O_1733,N_13744,N_13996);
or UO_1734 (O_1734,N_13605,N_14615);
and UO_1735 (O_1735,N_13500,N_14091);
and UO_1736 (O_1736,N_13532,N_14171);
and UO_1737 (O_1737,N_13527,N_13523);
and UO_1738 (O_1738,N_14840,N_14864);
and UO_1739 (O_1739,N_14823,N_14086);
xnor UO_1740 (O_1740,N_14174,N_14306);
xnor UO_1741 (O_1741,N_13544,N_14656);
and UO_1742 (O_1742,N_14534,N_13658);
nor UO_1743 (O_1743,N_14436,N_14097);
nand UO_1744 (O_1744,N_14967,N_13873);
and UO_1745 (O_1745,N_14402,N_13616);
and UO_1746 (O_1746,N_14689,N_14926);
and UO_1747 (O_1747,N_14653,N_13655);
nand UO_1748 (O_1748,N_13587,N_14284);
or UO_1749 (O_1749,N_14623,N_13763);
xnor UO_1750 (O_1750,N_14615,N_14384);
nand UO_1751 (O_1751,N_13692,N_13726);
nor UO_1752 (O_1752,N_13654,N_14147);
or UO_1753 (O_1753,N_14208,N_14299);
or UO_1754 (O_1754,N_14823,N_14433);
and UO_1755 (O_1755,N_14535,N_13673);
and UO_1756 (O_1756,N_14568,N_14355);
nand UO_1757 (O_1757,N_13632,N_14668);
nand UO_1758 (O_1758,N_13937,N_14344);
or UO_1759 (O_1759,N_14916,N_14790);
and UO_1760 (O_1760,N_14738,N_14536);
or UO_1761 (O_1761,N_14698,N_13623);
xnor UO_1762 (O_1762,N_14008,N_14438);
nor UO_1763 (O_1763,N_14809,N_13651);
nand UO_1764 (O_1764,N_14324,N_14182);
or UO_1765 (O_1765,N_13748,N_14730);
nor UO_1766 (O_1766,N_14057,N_14352);
and UO_1767 (O_1767,N_14590,N_14644);
or UO_1768 (O_1768,N_14921,N_13787);
nor UO_1769 (O_1769,N_13548,N_14828);
or UO_1770 (O_1770,N_13795,N_14967);
xnor UO_1771 (O_1771,N_13941,N_14339);
nor UO_1772 (O_1772,N_13918,N_14148);
xor UO_1773 (O_1773,N_13947,N_14631);
and UO_1774 (O_1774,N_13751,N_14740);
xor UO_1775 (O_1775,N_14625,N_14978);
or UO_1776 (O_1776,N_13666,N_13552);
or UO_1777 (O_1777,N_13834,N_13702);
nor UO_1778 (O_1778,N_14515,N_13784);
nand UO_1779 (O_1779,N_14695,N_14196);
or UO_1780 (O_1780,N_14234,N_13640);
nor UO_1781 (O_1781,N_14160,N_14992);
xor UO_1782 (O_1782,N_13684,N_14253);
and UO_1783 (O_1783,N_13845,N_14310);
or UO_1784 (O_1784,N_14832,N_13527);
nor UO_1785 (O_1785,N_14412,N_14847);
and UO_1786 (O_1786,N_13654,N_13848);
and UO_1787 (O_1787,N_14884,N_14482);
and UO_1788 (O_1788,N_13872,N_13570);
nand UO_1789 (O_1789,N_14249,N_14834);
and UO_1790 (O_1790,N_14293,N_14473);
nand UO_1791 (O_1791,N_14513,N_14786);
xnor UO_1792 (O_1792,N_14248,N_14015);
nor UO_1793 (O_1793,N_13552,N_14150);
nor UO_1794 (O_1794,N_14193,N_13744);
and UO_1795 (O_1795,N_13656,N_13716);
and UO_1796 (O_1796,N_14535,N_14873);
or UO_1797 (O_1797,N_13746,N_13827);
nor UO_1798 (O_1798,N_14041,N_14289);
nor UO_1799 (O_1799,N_14858,N_14170);
and UO_1800 (O_1800,N_14260,N_14521);
nand UO_1801 (O_1801,N_14006,N_14670);
nand UO_1802 (O_1802,N_14406,N_14148);
and UO_1803 (O_1803,N_14021,N_14323);
nand UO_1804 (O_1804,N_14598,N_13925);
nor UO_1805 (O_1805,N_13691,N_14379);
xnor UO_1806 (O_1806,N_14897,N_13960);
and UO_1807 (O_1807,N_13560,N_13739);
nor UO_1808 (O_1808,N_14215,N_14691);
and UO_1809 (O_1809,N_13697,N_13783);
or UO_1810 (O_1810,N_14674,N_13751);
nor UO_1811 (O_1811,N_14576,N_13982);
and UO_1812 (O_1812,N_14392,N_14458);
or UO_1813 (O_1813,N_14161,N_14033);
nor UO_1814 (O_1814,N_14156,N_14201);
nor UO_1815 (O_1815,N_14673,N_14501);
and UO_1816 (O_1816,N_13910,N_14554);
nor UO_1817 (O_1817,N_14691,N_13956);
nor UO_1818 (O_1818,N_14602,N_13942);
or UO_1819 (O_1819,N_13776,N_13981);
xor UO_1820 (O_1820,N_13774,N_14250);
nand UO_1821 (O_1821,N_14934,N_14981);
nand UO_1822 (O_1822,N_13597,N_14219);
nor UO_1823 (O_1823,N_14158,N_14320);
nand UO_1824 (O_1824,N_14032,N_13595);
nand UO_1825 (O_1825,N_14285,N_14195);
xnor UO_1826 (O_1826,N_14154,N_14746);
nor UO_1827 (O_1827,N_14375,N_13921);
or UO_1828 (O_1828,N_14005,N_13857);
or UO_1829 (O_1829,N_14499,N_14958);
and UO_1830 (O_1830,N_13902,N_14568);
and UO_1831 (O_1831,N_14299,N_13714);
and UO_1832 (O_1832,N_14942,N_13598);
nand UO_1833 (O_1833,N_14777,N_14262);
nand UO_1834 (O_1834,N_14168,N_13698);
nor UO_1835 (O_1835,N_14159,N_14652);
and UO_1836 (O_1836,N_14335,N_14785);
or UO_1837 (O_1837,N_14637,N_13618);
nand UO_1838 (O_1838,N_13697,N_13709);
nor UO_1839 (O_1839,N_14931,N_13685);
nand UO_1840 (O_1840,N_14295,N_14145);
xnor UO_1841 (O_1841,N_14944,N_14813);
nor UO_1842 (O_1842,N_13649,N_14996);
xnor UO_1843 (O_1843,N_13771,N_14558);
xor UO_1844 (O_1844,N_14220,N_13759);
and UO_1845 (O_1845,N_14923,N_14884);
or UO_1846 (O_1846,N_14525,N_14846);
xnor UO_1847 (O_1847,N_14968,N_14071);
xor UO_1848 (O_1848,N_13932,N_14595);
or UO_1849 (O_1849,N_14900,N_14746);
or UO_1850 (O_1850,N_13976,N_13610);
nor UO_1851 (O_1851,N_14843,N_14421);
xnor UO_1852 (O_1852,N_14583,N_13850);
nor UO_1853 (O_1853,N_14395,N_14190);
or UO_1854 (O_1854,N_14788,N_14694);
nor UO_1855 (O_1855,N_14794,N_13886);
xor UO_1856 (O_1856,N_14820,N_14906);
nand UO_1857 (O_1857,N_14950,N_14830);
xor UO_1858 (O_1858,N_13830,N_14276);
and UO_1859 (O_1859,N_14095,N_14058);
nand UO_1860 (O_1860,N_14301,N_14312);
nand UO_1861 (O_1861,N_14826,N_13986);
nand UO_1862 (O_1862,N_13726,N_14610);
or UO_1863 (O_1863,N_14305,N_14331);
and UO_1864 (O_1864,N_13628,N_14159);
xor UO_1865 (O_1865,N_14621,N_14567);
and UO_1866 (O_1866,N_14357,N_14643);
and UO_1867 (O_1867,N_14860,N_13938);
nand UO_1868 (O_1868,N_13568,N_13992);
and UO_1869 (O_1869,N_13609,N_14957);
nor UO_1870 (O_1870,N_14821,N_13994);
and UO_1871 (O_1871,N_13580,N_14614);
xor UO_1872 (O_1872,N_14031,N_14378);
or UO_1873 (O_1873,N_13637,N_14823);
nor UO_1874 (O_1874,N_13878,N_14673);
or UO_1875 (O_1875,N_14534,N_13896);
or UO_1876 (O_1876,N_14509,N_14341);
or UO_1877 (O_1877,N_14048,N_14964);
and UO_1878 (O_1878,N_14965,N_13595);
and UO_1879 (O_1879,N_14861,N_13964);
xnor UO_1880 (O_1880,N_14168,N_13805);
nand UO_1881 (O_1881,N_14159,N_14722);
nand UO_1882 (O_1882,N_14789,N_13673);
nand UO_1883 (O_1883,N_13671,N_14257);
and UO_1884 (O_1884,N_14841,N_13640);
and UO_1885 (O_1885,N_14886,N_13954);
and UO_1886 (O_1886,N_14556,N_14625);
xor UO_1887 (O_1887,N_14230,N_14890);
xor UO_1888 (O_1888,N_14844,N_14578);
nor UO_1889 (O_1889,N_14368,N_14989);
nand UO_1890 (O_1890,N_14434,N_14789);
nand UO_1891 (O_1891,N_13724,N_14472);
and UO_1892 (O_1892,N_14499,N_13504);
and UO_1893 (O_1893,N_14147,N_14078);
nor UO_1894 (O_1894,N_13803,N_14665);
nor UO_1895 (O_1895,N_13570,N_14173);
nor UO_1896 (O_1896,N_14887,N_13621);
nor UO_1897 (O_1897,N_13981,N_13618);
and UO_1898 (O_1898,N_14282,N_14354);
or UO_1899 (O_1899,N_13521,N_14244);
or UO_1900 (O_1900,N_14259,N_13647);
nand UO_1901 (O_1901,N_14206,N_14181);
xor UO_1902 (O_1902,N_13787,N_14077);
or UO_1903 (O_1903,N_13618,N_13875);
nor UO_1904 (O_1904,N_13556,N_14485);
nand UO_1905 (O_1905,N_14264,N_14424);
nand UO_1906 (O_1906,N_14959,N_13614);
or UO_1907 (O_1907,N_13532,N_13885);
and UO_1908 (O_1908,N_14012,N_14119);
or UO_1909 (O_1909,N_14376,N_14250);
nand UO_1910 (O_1910,N_13555,N_14420);
or UO_1911 (O_1911,N_14226,N_13667);
or UO_1912 (O_1912,N_14363,N_14586);
or UO_1913 (O_1913,N_13527,N_13560);
nor UO_1914 (O_1914,N_13827,N_13909);
and UO_1915 (O_1915,N_13557,N_13846);
or UO_1916 (O_1916,N_13760,N_13955);
nor UO_1917 (O_1917,N_13754,N_13653);
xnor UO_1918 (O_1918,N_14670,N_14169);
nand UO_1919 (O_1919,N_14708,N_13625);
and UO_1920 (O_1920,N_14571,N_14539);
and UO_1921 (O_1921,N_13658,N_13999);
and UO_1922 (O_1922,N_14720,N_14489);
or UO_1923 (O_1923,N_14280,N_14513);
nand UO_1924 (O_1924,N_14009,N_14472);
nand UO_1925 (O_1925,N_14241,N_14393);
nor UO_1926 (O_1926,N_14356,N_14346);
xnor UO_1927 (O_1927,N_13624,N_13816);
nand UO_1928 (O_1928,N_13517,N_13691);
and UO_1929 (O_1929,N_14032,N_13833);
nor UO_1930 (O_1930,N_13545,N_14318);
nor UO_1931 (O_1931,N_13626,N_14511);
xnor UO_1932 (O_1932,N_14926,N_14013);
and UO_1933 (O_1933,N_13691,N_13858);
and UO_1934 (O_1934,N_14546,N_14620);
and UO_1935 (O_1935,N_14142,N_14914);
and UO_1936 (O_1936,N_13884,N_13846);
nand UO_1937 (O_1937,N_14181,N_14674);
or UO_1938 (O_1938,N_13520,N_13886);
nor UO_1939 (O_1939,N_13854,N_14134);
or UO_1940 (O_1940,N_14945,N_13884);
xnor UO_1941 (O_1941,N_13936,N_13944);
nor UO_1942 (O_1942,N_14340,N_13889);
and UO_1943 (O_1943,N_13941,N_14465);
and UO_1944 (O_1944,N_14103,N_14248);
nor UO_1945 (O_1945,N_13662,N_14012);
or UO_1946 (O_1946,N_14343,N_14433);
xnor UO_1947 (O_1947,N_13505,N_13653);
and UO_1948 (O_1948,N_13844,N_14726);
or UO_1949 (O_1949,N_14876,N_14802);
xor UO_1950 (O_1950,N_14629,N_14863);
nand UO_1951 (O_1951,N_13629,N_14371);
or UO_1952 (O_1952,N_14341,N_13615);
xnor UO_1953 (O_1953,N_13896,N_14504);
and UO_1954 (O_1954,N_14875,N_14310);
or UO_1955 (O_1955,N_14277,N_14911);
nand UO_1956 (O_1956,N_14944,N_14003);
or UO_1957 (O_1957,N_13747,N_14660);
nand UO_1958 (O_1958,N_14940,N_14570);
and UO_1959 (O_1959,N_14026,N_14394);
nor UO_1960 (O_1960,N_14557,N_14220);
or UO_1961 (O_1961,N_14196,N_13777);
or UO_1962 (O_1962,N_14482,N_14669);
xor UO_1963 (O_1963,N_13964,N_13791);
nor UO_1964 (O_1964,N_13730,N_13631);
nor UO_1965 (O_1965,N_13621,N_14428);
and UO_1966 (O_1966,N_14192,N_13641);
or UO_1967 (O_1967,N_14275,N_13928);
and UO_1968 (O_1968,N_13675,N_14300);
nand UO_1969 (O_1969,N_13979,N_14950);
xnor UO_1970 (O_1970,N_14250,N_14410);
nor UO_1971 (O_1971,N_13892,N_14889);
nand UO_1972 (O_1972,N_13816,N_14261);
nand UO_1973 (O_1973,N_13830,N_13915);
nor UO_1974 (O_1974,N_14238,N_13940);
nor UO_1975 (O_1975,N_14520,N_14333);
or UO_1976 (O_1976,N_13733,N_14097);
nand UO_1977 (O_1977,N_14960,N_14678);
nor UO_1978 (O_1978,N_14130,N_14886);
and UO_1979 (O_1979,N_14444,N_13851);
xnor UO_1980 (O_1980,N_14897,N_14247);
or UO_1981 (O_1981,N_14549,N_14403);
xnor UO_1982 (O_1982,N_14639,N_13849);
nor UO_1983 (O_1983,N_13645,N_13846);
nor UO_1984 (O_1984,N_14305,N_14148);
xor UO_1985 (O_1985,N_14619,N_14076);
and UO_1986 (O_1986,N_14154,N_14038);
nand UO_1987 (O_1987,N_14574,N_13958);
nor UO_1988 (O_1988,N_14513,N_14099);
xnor UO_1989 (O_1989,N_14504,N_14738);
nand UO_1990 (O_1990,N_14102,N_13902);
and UO_1991 (O_1991,N_13815,N_14426);
nor UO_1992 (O_1992,N_14874,N_13644);
nor UO_1993 (O_1993,N_13984,N_13537);
or UO_1994 (O_1994,N_14541,N_13601);
nor UO_1995 (O_1995,N_14353,N_14309);
or UO_1996 (O_1996,N_14696,N_13953);
nor UO_1997 (O_1997,N_13881,N_14779);
or UO_1998 (O_1998,N_14501,N_13880);
nand UO_1999 (O_1999,N_14163,N_13853);
endmodule